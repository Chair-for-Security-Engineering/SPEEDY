
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_SPEEDY_Top is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_SPEEDY_Top;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Rounds7_0 is

   port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : out
         std_logic_vector (191 downto 0));

end SPEEDY_Rounds7_0;

architecture SYN_Behavioral of SPEEDY_Rounds7_0 is

   component INV_X2
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( I0, I1, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X4
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X12
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X8
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X8
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n7, n10, n11, n12, n13, n17, n19, n21, n25, n26, n28,
      n29, n32, n35, n36, n37, n40, n42, n43, n45, n46, n50, n52, n53, n54, n56
      , n57, n59, n61, n62, n63, n64, n70, n71, n76, n81, n85, n89, n94, n98, 
      n99, n104, n105, n106, n109, n110, n113, n114, n118, n119, n121, n122, 
      n123, n124, n126, n129, n130, n133, n135, n137, n138, n139, n140, n142, 
      n149, n154, n155, n156, n157, n158, n159, n160, n161, n164, n167, n170, 
      n171, n178, n180, n182, n183, n184, n187, n190, n193, n195, n196, n197, 
      n198, n199, n200, n205, n207, n208, n209, n212, n214, n215, n217, n219, 
      n220, n224, n229, n230, n231, n232, n233, n237, n238, n242, n248, n250, 
      n251, n252, n253, n254, n257, n259, n260, n261, n263, n266, n269, n272, 
      n274, n275, n277, n278, n280, n281, n282, n284, n287, n288, n291, n293, 
      n295, n296, n298, n299, n301, n302, n305, n306, n307, n309, n310, n311, 
      n314, n317, n318, n319, n320, n321, n326, n327, n331, n334, n336, n342, 
      n343, n344, n345, n346, n347, n353, n354, n355, n357, n359, n360, n362, 
      n364, n365, n367, n370, n371, n372, n378, n379, n382, n383, n384, n385, 
      n386, n387, n388, n391, n396, n399, n400, n404, n406, n407, n411, n412, 
      n416, n422, n423, n424, n425, n427, n430, n431, n434, n436, n437, n438, 
      n439, n440, n441, n442, n443, n445, n446, n447, n449, n450, n451, n452, 
      n454, n455, n457, n459, n462, n465, n467, n471, n474, n476, n479, n481, 
      n482, n484, n485, n487, n489, n491, n494, n495, n496, n502, n505, n507, 
      n509, n514, n515, n517, n518, n523, n524, n525, n526, n528, n529, n530, 
      n531, n532, n533, n538, n540, n541, n542, n543, n545, n547, n548, n550, 
      n551, n552, n554, n556, n557, n560, n562, n566, n576, n579, n580, n583, 
      n584, n585, n586, n587, n588, n589, n591, n596, n598, n599, n601, n603, 
      n605, n606, n608, n609, n611, n614, n615, n616, n619, n621, n626, n628, 
      n629, n632, n633, n635, n636, n637, n638, n639, n640, n642, n644, n646, 
      n648, n649, n650, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n672, n673, n674, n675, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n688, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n704, 
      n705, n706, n707, n708, n709, n710, n711, n713, n714, n718, n719, n720, 
      n721, n722, n723, n724, n727, n728, n729, n730, n731, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n754, n755, n756, n759, n760, n761, n762, n763, 
      n764, n765, n767, n769, n770, n771, n772, n773, n774, n775, n777, n778, 
      n779, n780, n781, n782, n783, n784, n787, n788, n789, n790, n791, n792, 
      n794, n798, n800, n801, n802, n807, n808, n810, n812, n813, n814, n815, 
      n816, n817, n819, n820, n821, n823, n824, n825, n826, n828, n830, n831, 
      n832, n833, n834, n835, n837, n838, n839, n840, n841, n844, n845, n846, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n865, n866, n867, n869, n870, n871, n873, n875, 
      n876, n877, n878, n879, n881, n882, n883, n885, n886, n888, n889, n892, 
      n893, n894, n896, n898, n900, n902, n903, n906, n907, n910, n911, n914, 
      n915, n916, n917, n918, n919, n920, n921, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n933, n934, n935, n936, n937, n938, n939, n941, 
      n943, n944, n945, n946, n948, n949, n950, n951, n952, n953, n954, n955, 
      n957, n958, n959, n960, n961, n962, n963, n965, n966, n967, n968, n969, 
      n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, 
      n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, 
      n995, n997, n998, n999, n1000, n1002, n1003, n1006, n1008, n1009, n1010, 
      n1011, n1012, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, 
      n1022, n1024, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1038, n1039, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1065, n1066, n1068, 
      n1069, n1070, n1071, n1072, n1073, n1074, n1076, n1077, n1079, n1080, 
      n1081, n1082, n1084, n1085, n1086, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1112, n1113, n1115, 
      n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, 
      n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, 
      n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, 
      n1146, n1147, n1148, n1149, n1151, n1152, n1154, n1155, n1156, n1157, 
      n1158, n1159, n1160, n1161, n1162, n1163, n1165, n1167, n1169, n1170, 
      n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1181, 
      n1182, n1183, n1184, n1186, n1187, n1189, n1190, n1192, n1193, n1194, 
      n1195, n1196, n1197, n1198, n1200, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1211, n1212, n1214, n1215, n1217, n1218, n1220, 
      n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1229, n1230, n1231, 
      n1232, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1242, n1243, 
      n1244, n1245, n1249, n1252, n1253, n1254, n1255, n1256, n1257, n1258, 
      n1259, n1260, n1261, n1262, n1263, n1265, n1267, n1268, n1269, n1270, 
      n1271, n1273, n1274, n1275, n1276, n1279, n1280, n1282, n1283, n1284, 
      n1285, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1297, 
      n1298, n1299, n1300, n1301, n1302, n1304, n1306, n1307, n1308, n1310, 
      n1312, n1313, n1314, n1315, n1316, n1318, n1319, n1320, n1322, n1323, 
      n1324, n1326, n1327, n1328, n1329, n1331, n1332, n1333, n1334, n1335, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1344, n1345, n1346, n1348, 
      n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1361, n1362, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1374, n1375, n1377, n1378, n1379, n1380, n1382, n1383, n1385, n1387, 
      n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1396, n1397, n1398, 
      n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, 
      n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, 
      n1419, n1420, n1424, n1425, n1426, n1427, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1444, n1445, n1446, n1447, n1448, n1450, n1451, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1477, 
      n1478, n1480, n1481, n1483, n1484, n1486, n1487, n1489, n1490, n1491, 
      n1492, n1493, n1494, n1495, n1497, n1500, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1509, n1510, n1511, n1512, n1514, n1515, n1518, n1519, 
      n1520, n1521, n1522, n1523, n1524, n1527, n1528, n1529, n1530, n1531, 
      n1532, n1534, n1535, n1536, n1537, n1539, n1541, n1543, n1545, n1546, 
      n1547, n1548, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1563, n1564, n1565, n1566, n1567, n1570, n1573, 
      n1574, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1586, 
      n1587, n1588, n1589, n1591, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1612, n1613, n1614, n1616, n1617, n1618, n1619, n1620, n1621, 
      n1622, n1623, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1666, n1667, 
      n1668, n1669, n1670, n1671, n1672, n1673, n1675, n1676, n1678, n1679, 
      n1680, n1681, n1683, n1684, n1686, n1687, n1688, n1689, n1690, n1692, 
      n1693, n1694, n1695, n1697, n1698, n1699, n1700, n1702, n1703, n1704, 
      n1706, n1707, n1708, n1710, n1711, n1713, n1714, n1717, n1718, n1719, 
      n1722, n1723, n1724, n1725, n1726, n1727, n1730, n1733, n1734, n1735, 
      n1737, n1738, n1740, n1741, n1742, n1743, n1745, n1746, n1752, n1753, 
      n1755, n1757, n1758, n1759, n1760, n1763, n1765, n1766, n1769, n1771, 
      n1775, n1777, n1778, n1781, n1782, n1783, n1784, n1785, n1786, n1787, 
      n1788, n1790, n1791, n1792, n1793, n1794, n1796, n1797, n1798, n1799, 
      n1802, n1805, n1807, n1808, n1809, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1827, n1829, 
      n1830, n1831, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1842, 
      n1843, n1844, n1845, n1847, n1849, n1850, n1851, n1852, n1855, n1859, 
      n1861, n1862, n1864, n1865, n1866, n1867, n1868, n1872, n1873, n1874, 
      n1875, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, 
      n1886, n1890, n1891, n1893, n1894, n1895, n1896, n1897, n1898, n1902, 
      n1904, n1906, n1907, n1909, n1911, n1912, n1913, n1914, n1915, n1917, 
      n1918, n1919, n1921, n1923, n1929, n1930, n1932, n1933, n1934, n1936, 
      n1938, n1939, n1940, n1944, n1945, n1946, n1947, n1948, n1949, n1951, 
      n1953, n1954, n1956, n1961, n1962, n1965, n1966, n1969, n1971, n1978, 
      n1980, n1984, n1986, n1989, n1990, n1991, n1992, n1993, n1995, n1996, 
      n1997, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2008, n2009, 
      n2012, n2013, n2016, n2017, n2018, n2022, n2023, n2025, n2028, n2029, 
      n2030, n2031, n2032, n2035, n2036, n2041, n2042, n2044, n2045, n2046, 
      n2047, n2049, n2050, n2052, n2055, n2057, n2058, n2059, n2060, n2062, 
      n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2073, n2075, n2076, 
      n2077, n2078, n2079, n2081, n2082, n2084, n2085, n2086, n2087, n2088, 
      n2089, n2091, n2092, n2094, n2096, n2097, n2100, n2101, n2102, n2104, 
      n2105, n2106, n2107, n2110, n2111, n2112, n2113, n2114, n2116, n2117, 
      n2119, n2120, n2121, n2122, n2124, n2125, n2126, n2127, n2128, n2129, 
      n2130, n2132, n2134, n2135, n2136, n2138, n2139, n2140, n2142, n2145, 
      n2147, n2148, n2149, n2150, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2166, n2167, n2168, 
      n2170, n2175, n2176, n2177, n2178, n2182, n2184, n2185, n2186, n2187, 
      n2189, n2190, n2191, n2192, n2193, n2195, n2196, n2198, n2199, n2200, 
      n2202, n2203, n2205, n2207, n2208, n2209, n2211, n2214, n2215, n2216, 
      n2217, n2218, n2220, n2221, n2222, n2223, n2226, n2229, n2231, n2233, 
      n2234, n2235, n2236, n2237, n2238, n2239, n2242, n2243, n2246, n2247, 
      n2248, n2250, n2253, n2254, n2257, n2258, n2259, n2260, n2262, n2263, 
      n2264, n2268, n2269, n2270, n2272, n2273, n2274, n2276, n2277, n2278, 
      n2279, n2280, n2281, n2283, n2284, n2285, n2288, n2292, n2294, n2296, 
      n2297, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2309, n2310, 
      n2311, n2316, n2317, n2318, n2319, n2321, n2322, n2326, n2327, n2328, 
      n2330, n2331, n2333, n2334, n2335, n2336, n2338, n2339, n2340, n2341, 
      n2342, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2354, n2356, 
      n2362, n2363, n2364, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2386, n2387, 
      n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2398, 
      n2400, n2402, n2403, n2404, n2405, n2410, n2413, n2416, n2417, n2418, 
      n2421, n2423, n2424, n2428, n2429, n2430, n2431, n2434, n2435, n2436, 
      n2437, n2439, n2443, n2445, n2446, n2448, n2449, n2450, n2451, n2453, 
      n2454, n2456, n2457, n2458, n2461, n2462, n2464, n2465, n2466, n2467, 
      n2469, n2471, n2473, n2474, n2475, n2476, n2478, n2479, n2480, n2481, 
      n2482, n2484, n2485, n2487, n2488, n2489, n2490, n2491, n2493, n2495, 
      n2496, n2498, n2500, n2502, n2503, n2505, n2506, n2507, n2510, n2511, 
      n2512, n2515, n2518, n2519, n2520, n2522, n2524, n2525, n2526, n2527, 
      n2529, n2530, n2531, n2532, n2533, n2534, n2537, n2541, n2542, n2543, 
      n2544, n2545, n2546, n2547, n2549, n2553, n2554, n2555, n2557, n2559, 
      n2560, n2561, n2563, n2566, n2569, n2572, n2573, n2574, n2576, n2579, 
      n2580, n2581, n2582, n2585, n2586, n2587, n2588, n2589, n2590, n2592, 
      n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2603, n2604, 
      n2607, n2608, n2610, n2613, n2614, n2615, n2616, n2618, n2621, n2622, 
      n2623, n2625, n2626, n2627, n2628, n2629, n2630, n2632, n2633, n2634, 
      n2635, n2637, n2639, n2643, n2644, n2645, n2646, n2647, n2648, n2649, 
      n2650, n2651, n2653, n2654, n2656, n2657, n2658, n2660, n2662, n2663, 
      n2664, n2666, n2667, n2668, n2671, n2674, n2675, n2677, n2678, n2679, 
      n2681, n2682, n2683, n2684, n2685, n2688, n2690, n2692, n2695, n2696, 
      n2697, n2698, n2701, n2703, n2704, n2705, n2707, n2709, n2711, n2712, 
      n2713, n2714, n2716, n2717, n2721, n2722, n2725, n2726, n2727, n2728, 
      n2730, n2731, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, 
      n2743, n2745, n2746, n2747, n2751, n2752, n2753, n2754, n2757, n2758, 
      n2759, n2760, n2761, n2765, n2766, n2767, n2768, n2769, n2771, n2772, 
      n2774, n2778, n2780, n2781, n2782, n2784, n2785, n2788, n2789, n2790, 
      n2792, n2794, n2795, n2796, n2798, n2799, n2800, n2801, n2802, n2803, 
      n2805, n2806, n2808, n2812, n2813, n2814, n2815, n2816, n2818, n2819, 
      n2822, n2823, n2824, n2825, n2830, n2832, n2833, n2835, n2837, n2838, 
      n2839, n2840, n2841, n2842, n2846, n2847, n2848, n2850, n2853, n2856, 
      n2858, n2859, n2860, n2861, n2864, n2865, n2866, n2867, n2868, n2870, 
      n2872, n2873, n2874, n2876, n2877, n2878, n2880, n2881, n2882, n2883, 
      n2886, n2888, n2889, n2891, n2892, n2895, n2896, n2898, n2899, n2900, 
      n2903, n2904, n2905, n2906, n2907, n2909, n2910, n2914, n2915, n2919, 
      n2920, n2921, n2922, n2923, n2927, n2928, n2929, n2930, n2931, n2932, 
      n2933, n2935, n2937, n2940, n2941, n2942, n2943, n2944, n2945, n2946, 
      n2947, n2949, n2950, n2953, n2954, n2955, n2957, n2958, n2959, n2960, 
      n2961, n2962, n2965, n2966, n2967, n2968, n2969, n2971, n2972, n2974, 
      n2975, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2985, n2986, 
      n2987, n2988, n2989, n2990, n2991, n2995, n2996, n2997, n2998, n3001, 
      n3002, n3003, n3004, n3005, n3006, n3010, n3011, n3012, n3013, n3014, 
      n3015, n3016, n3018, n3019, n3021, n3022, n3023, n3024, n3025, n3027, 
      n3028, n3029, n3031, n3032, n3035, n3036, n3037, n3039, n3040, n3041, 
      n3044, n3045, n3046, n3047, n3048, n3050, n3052, n3053, n3055, n3056, 
      n3057, n3058, n3059, n3060, n3065, n3066, n3067, n3069, n3070, n3071, 
      n3072, n3076, n3077, n3081, n3082, n3083, n3085, n3086, n3088, n3090, 
      n3091, n3092, n3093, n3095, n3096, n3097, n3098, n3099, n3100, n3101, 
      n3102, n3103, n3105, n3106, n3107, n3109, n3110, n3111, n3112, n3114, 
      n3116, n3117, n3118, n3119, n3120, n3122, n3124, n3125, n3126, n3127, 
      n3128, n3129, n3133, n3134, n3135, n3136, n3137, n3140, n3141, n3142, 
      n3145, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, 
      n3159, n3161, n3163, n3164, n3166, n3167, n3169, n3170, n3172, n3174, 
      n3175, n3181, n3185, n3186, n3187, n3188, n3190, n3191, n3192, n3193, 
      n3194, n3195, n3198, n3199, n3200, n3203, n3206, n3207, n3213, n3214, 
      n3215, n3217, n3218, n3219, n3221, n3223, n3224, n3226, n3227, n3228, 
      n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3239, 
      n3240, n3241, n3242, n3244, n3245, n3246, n3247, n3248, n3250, n3252, 
      n3253, n3255, n3256, n3257, n3258, n3261, n3262, n3263, n3264, n3265, 
      n3266, n3267, n3268, n3269, n3270, n3271, n3273, n3274, n3275, n3276, 
      n3277, n3278, n3280, n3282, n3283, n3284, n3285, n3287, n3288, n3289, 
      n3290, n3292, n3293, n3294, n3295, n3297, n3299, n3301, n3303, n3304, 
      n3305, n3307, n3309, n3310, n3312, n3313, n3316, n3317, n3319, n3320, 
      n3323, n3325, n3326, n3327, n3328, n3330, n3331, n3332, n3333, n3336, 
      n3337, n3342, n3343, n3345, n3346, n3348, n3349, n3350, n3351, n3352, 
      n3356, n3359, n3360, n3361, n3363, n3364, n3365, n3366, n3368, n3369, 
      n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3382, 
      n3383, n3386, n3387, n3388, n3389, n3390, n3392, n3393, n3395, n3398, 
      n3399, n3402, n3404, n3409, n3410, n3411, n3412, n3413, n3415, n3417, 
      n3422, n3424, n3426, n3427, n3429, n3430, n3433, n3434, n3435, n3437, 
      n3438, n3441, n3443, n3445, n3446, n3447, n3448, n3449, n3450, n3451, 
      n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3461, n3462, 
      n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
      n3473, n3474, n3475, n3476, n3478, n3480, n3484, n3486, n3487, n3488, 
      n3489, n3490, n3493, n3495, n3496, n3497, n3498, n3499, n3501, n3503, 
      n3506, n3507, n3509, n3510, n3511, n3513, n3514, n3515, n3516, n3517, 
      n3518, n3519, n3521, n3522, n3523, n3525, n3526, n3527, n3528, n3529, 
      n3530, n3531, n3532, n3533, n3534, n3535, n3538, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3557, n3559, n3560, n3561, n3562, n3564, n3568, 
      n3571, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3581, n3583, 
      n3584, n3585, n3589, n3593, n3598, n3599, n3600, n3601, n3602, n3603, 
      n3604, n3605, n3606, n3609, n3610, n3611, n3612, n3614, n3616, n3618, 
      n3619, n3620, n3621, n3622, n3623, n3624, n3626, n3627, n3628, n3629, 
      n3630, n3631, n3632, n3633, n3634, n3637, n3638, n3639, n3641, n3642, 
      n3644, n3645, n3647, n3649, n3650, n3651, n3652, n3653, n3654, n3655, 
      n3656, n3657, n3659, n3662, n3663, n3664, n3665, n3666, n3668, n3669, 
      n3670, n3671, n3672, n3674, n3675, n3676, n3677, n3678, n3679, n3680, 
      n3681, n3682, n3683, n3685, n3687, n3690, n3691, n3692, n3693, n3694, 
      n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3703, n3705, n3707, 
      n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, 
      n3718, n3722, n3723, n3725, n3726, n3727, n3731, n3732, n3733, n3734, 
      n3735, n3736, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, 
      n3750, n3751, n3760, n3761, n3769, n3770, n3771, n3773, n3776, n3777, 
      n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3787, n3790, 
      n3791, n3792, n3793, n3794, n3795, n3798, n3799, n3800, n3801, n3802, 
      n3803, n3804, n3806, n3807, n3809, n3811, n3813, n3815, n3818, n3819, 
      n3820, n3821, n3823, n3824, n3825, n3826, n3827, n3832, n3833, n3835, 
      n3837, n3838, n3839, n3840, n3843, n3844, n3845, n3846, n3849, n3850, 
      n3851, n3852, n3855, n3857, n3858, n3860, n3861, n3862, n3863, n3864, 
      n3865, n3867, n3868, n3869, n3872, n3873, n3874, n3877, n3878, n3879, 
      n3884, n3885, n3886, n3887, n3889, n3890, n3891, n3893, n3894, n3895, 
      n3896, n3897, n3898, n3899, n3900, n3903, n3904, n3906, n3907, n3909, 
      n3912, n3913, n3914, n3916, n3917, n3918, n3919, n3920, n3921, n3923, 
      n3926, n3927, n3928, n3929, n3930, n3932, n3935, n3937, n3938, n3941, 
      n3943, n3944, n3945, n3947, n3949, n3951, n3952, n3953, n3954, n3956, 
      n3958, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3969, n3971, 
      n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3981, n3983, 
      n3985, n3986, n3988, n3989, n3990, n3992, n3993, n3995, n3996, n3998, 
      n3999, n4000, n4001, n4002, n4005, n4007, n4008, n4009, n4010, n4011, 
      n4013, n4014, n4015, n4016, n4018, n4021, n4022, n4023, n4024, n4025, 
      n4028, n4033, n4034, n4037, n4038, n4039, n4041, n4045, n4046, n4047, 
      n4048, n4050, n4051, n4053, n4056, n4057, n4058, n4059, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4070, n4072, n4073, n4075, n4076, n4077, 
      n4079, n4080, n4081, n4083, n4084, n4085, n4086, n4089, n4090, n4091, 
      n4092, n4093, n4094, n4095, n4098, n4099, n4100, n4102, n4104, n4105, 
      n4107, n4108, n4109, n4110, n4111, n4114, n4116, n4117, n4118, n4119, 
      n4120, n4121, n4122, n4123, n4126, n4127, n4128, n4129, n4131, n4132, 
      n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4147, 
      n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4159, n4160, 
      n4161, n4162, n4163, n4168, n4169, n4171, n4172, n4173, n4176, n4177, 
      n4178, n4179, n4182, n4183, n4184, n4188, n4189, n4190, n4191, n4192, 
      n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4204, 
      n4205, n4207, n4209, n4210, n4211, n4214, n4215, n4216, n4217, n4218, 
      n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4231, 
      n4232, n4235, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, 
      n4246, n4247, n4248, n4251, n4253, n4254, n4255, n4256, n4257, n4258, 
      n4266, n4268, n4269, n4270, n4271, n4272, n4273, n4277, n4278, n4279, 
      n4280, n4282, n4283, n4284, n4286, n4287, n4288, n4290, n4291, n4292, 
      n4293, n4294, n4296, n4297, n4298, n4300, n4301, n4302, n4305, n4306, 
      n4308, n4313, n4314, n4315, n4316, n4317, n4318, n4321, n4322, n4323, 
      n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4332, n4333, n4334, 
      n4335, n4336, n4337, n4339, n4340, n4341, n4342, n4345, n4346, n4347, 
      n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, 
      n4359, n4360, n4361, n4362, n4364, n4366, n4367, n4368, n4369, n4371, 
      n4372, n4373, n4375, n4377, n4378, n4379, n4381, n4382, n4384, n4385, 
      n4386, n4387, n4388, n4391, n4392, n4393, n4396, n4397, n4398, n4399, 
      n4400, n4401, n4409, n4410, n4411, n4412, n4413, n4415, n4416, n4417, 
      n4419, n4423, n4424, n4427, n4428, n4429, n4430, n4431, n4433, n4434, 
      n4436, n4438, n4439, n4440, n4441, n4442, n4443, n4445, n4447, n4448, 
      n4449, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, 
      n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4472, 
      n4473, n4475, n4476, n4477, n4479, n4483, n4484, n4485, n4486, n4489, 
      n4490, n4492, n4493, n4494, n4495, n4497, n4498, n4499, n4500, n4501, 
      n4502, n4503, n4504, n4506, n4507, n4508, n4511, n4512, n4515, n4516, 
      n4518, n4519, n4520, n4523, n4524, n4525, n4526, n4527, n4528, n4529, 
      n4531, n4534, n4536, n4538, n4540, n4542, n4543, n4549, n4550, n4551, 
      n4552, n4553, n4556, n4558, n4559, n4560, n4561, n4562, n4563, n4564, 
      n4565, n4566, n4568, n4570, n4572, n4573, n4574, n4576, n4578, n4579, 
      n4580, n4581, n4582, n4583, n4584, n4587, n4588, n4589, n4591, n4592, 
      n4595, n4597, n4599, n4600, n4601, n4602, n4603, n4604, n4606, n4608, 
      n4610, n4611, n4612, n4613, n4616, n4618, n4619, n4620, n4621, n4622, 
      n4624, n4625, n4627, n4629, n4630, n4631, n4632, n4633, n4634, n4636, 
      n4637, n4638, n4640, n4641, n4642, n4644, n4646, n4647, n4649, n4651, 
      n4655, n4656, n4658, n4660, n4661, n4662, n4664, n4665, n4666, n4667, 
      n4668, n4669, n4670, n4671, n4673, n4674, n4677, n4682, n4686, n4687, 
      n4688, n4689, n4690, n4694, n4697, n4698, n4699, n4700, n4702, n4703, 
      n4704, n4707, n4709, n4713, n4714, n4715, n4716, n4720, n4724, n4726, 
      n4729, n4730, n4734, n4736, n4737, n4738, n4739, n4741, n4743, n4745, 
      n4746, n4748, n4750, n4752, n4754, n4755, n4756, n4759, n4760, n4761, 
      n4765, n4766, n4767, n4768, n4769, n4771, n4772, n4773, n4775, n4776, 
      n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4788, n4790, n4791, 
      n4792, n4794, n4796, n4799, n4800, n4801, n4803, n4805, n4807, n4808, 
      n4809, n4815, n4816, n4819, n4821, n4823, n4824, n4825, n4827, n4828, 
      n4829, n4832, n4833, n4834, n4840, n4841, n4845, n4846, n4847, n4849, 
      n4850, n4851, n4852, n4853, n4854, n4856, n4857, n4858, n4859, n4862, 
      n4864, n4865, n4866, n4867, n4868, n4869, n4871, n4874, n4875, n4876, 
      n4878, n4879, n4880, n4882, n4883, n4884, n4885, n4886, n4887, n4888, 
      n4889, n4890, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, 
      n4901, n4902, n4903, n4905, n4908, n4909, n4910, n4913, n4914, n4915, 
      n4916, n4917, n4918, n4919, n4924, n4925, n4926, n4927, n4929, n4931, 
      n4932, n4934, n4935, n4936, n4937, n4938, n4941, n4945, n4946, n4947, 
      n4948, n4949, n4950, n4952, n4956, n4957, n4958, n4959, n4960, n4963, 
      n4964, n4967, n4968, n4969, n4970, n4972, n4973, n4975, n4976, n4977, 
      n4978, n4980, n4982, n4986, n4987, n4988, n4989, n4990, n4991, n4992, 
      n4993, n4997, n4999, n5001, n5002, n5003, n5005, n5006, n5009, n5010, 
      n5011, n5012, n5014, n5015, n5018, n5019, n5020, n5021, n5022, n5023, 
      n5024, n5026, n5027, n5028, n5030, n5031, n5033, n5034, n5035, n5037, 
      n5038, n5039, n5041, n5042, n5044, n5047, n5048, n5049, n5050, n5051, 
      n5053, n5054, n5055, n5056, n5058, n5059, n5061, n5062, n5063, n5065, 
      n5066, n5067, n5070, n5071, n5073, n5075, n5077, n5078, n5080, n5082, 
      n5083, n5084, n5085, n5086, n5088, n5089, n5090, n5091, n5093, n5094, 
      n5096, n5098, n5100, n5101, n5103, n5104, n5107, n5108, n5110, n5111, 
      n5112, n5114, n5115, n5116, n5118, n5119, n5120, n5122, n5123, n5124, 
      n5126, n5127, n5129, n5130, n5131, n5132, n5137, n5138, n5139, n5140, 
      n5142, n5143, n5144, n5145, n5146, n5147, n5149, n5150, n5151, n5152, 
      n5153, n5154, n5156, n5158, n5160, n5161, n5162, n5164, n5166, n5167, 
      n5171, n5172, n5174, n5176, n5177, n5179, n5181, n5183, n5184, n5185, 
      n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, 
      n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5214, 
      n5215, n5218, n5219, n5220, n5221, n5223, n5224, n5225, n5226, n5227, 
      n5228, n5229, n5231, n5232, n5233, n5235, n5236, n5237, n5238, n5239, 
      n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5251, 
      n5252, n5253, n5254, n5255, n5258, n5261, n5263, n5264, n5266, n5270, 
      n5271, n5274, n5276, n5277, n5279, n5282, n5283, n5284, n5285, n5286, 
      n5287, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5297, n5299, 
      n5300, n5302, n5303, n5304, n5305, n5306, n5308, n5309, n5311, n5312, 
      n5314, n5315, n5316, n5317, n5318, n5320, n5322, n5323, n5325, n5326, 
      n5327, n5330, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5342, 
      n5343, n5344, n5345, n5347, n5348, n5350, n5351, n5352, n5354, n5355, 
      n5356, n5357, n5358, n5359, n5360, n5361, n5363, n5365, n5366, n5367, 
      n5369, n5370, n5371, n5374, n5377, n5380, n5381, n5382, n5383, n5384, 
      n5385, n5387, n5388, n5389, n5390, n5391, n5392, n5394, n5395, n5396, 
      n5397, n5398, n5399, n5401, n5402, n5403, n5405, n5407, n5408, n5410, 
      n5412, n5413, n5414, n5415, n5417, n5418, n5422, n5423, n5424, n5427, 
      n5430, n5431, n5432, n5433, n5434, n5436, n5437, n5438, n5439, n5441, 
      n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, 
      n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5461, n5462, 
      n5463, n5464, n5465, n5467, n5468, n5469, n5470, n5471, n5472, n5473, 
      n5474, n5475, n5477, n5479, n5480, n5481, n5483, n5484, n5486, n5487, 
      n5488, n5490, n5491, n5492, n5494, n5495, n5496, n5497, n5498, n5500, 
      n5501, n5503, n5504, n5505, n5508, n5509, n5510, n5511, n5514, n5515, 
      n5516, n5517, n5518, n5519, n5520, n5522, n5524, n5525, n5527, n5530, 
      n5531, n5533, n5534, n5535, n5537, n5538, n5539, n5540, n5541, n5542, 
      n5543, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, 
      n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5569, n5570, n5571, 
      n5572, n5576, n5577, n5579, n5580, n5581, n5582, n5583, n5584, n5586, 
      n5587, n5588, n5589, n5590, n5591, n5592, n5596, n5597, n5598, n5599, 
      n5600, n5601, n5603, n5607, n5609, n5610, n5613, n5616, n5617, n5618, 
      n5619, n5621, n5622, n5623, n5625, n5628, n5629, n5630, n5632, n5634, 
      n5635, n5636, n5637, n5638, n5639, n5641, n5642, n5645, n5646, n5647, 
      n5648, n5649, n5650, n5651, n5652, n5653, n5655, n5656, n5657, n5658, 
      n5662, n5664, n5665, n5667, n5669, n5670, n5671, n5672, n5674, n5675, 
      n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5686, n5687, 
      n5688, n5690, n5691, n5692, n5693, n5694, n5695, n5697, n5698, n5699, 
      n5702, n5703, n5705, n5706, n5707, n5709, n5710, n5711, n5712, n5713, 
      n5714, n5716, n5717, n5719, n5720, n5721, n5722, n5723, n5724, n5725, 
      n5726, n5728, n5730, n5731, n5732, n5733, n5734, n5736, n5737, n5738, 
      n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, 
      n5750, n5751, n5753, n5755, n5757, n5758, n5759, n5760, n5761, n5762, 
      n5763, n5764, n5765, n5766, n5768, n5769, n5770, n5771, n5772, n5773, 
      n5774, n5775, n5776, n5777, n5778, n5779, n5781, n5782, n5785, n5786, 
      n5787, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5798, 
      n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5810, n5811, 
      n5813, n5814, n5815, n5816, n5817, n5819, n5820, n5821, n5822, n5823, 
      n5825, n5829, n5830, n5831, n5834, n5835, n5836, n5837, n5838, n5839, 
      n5841, n5842, n5843, n5844, n5845, n5848, n5849, n5851, n5853, n5854, 
      n5855, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5866, 
      n5867, n5869, n5871, n5873, n5874, n5876, n5877, n5878, n5880, n5881, 
      n5882, n5883, n5884, n5885, n5886, n5888, n5889, n5890, n5891, n5892, 
      n5894, n5895, n5896, n5897, n5899, n5900, n5901, n5902, n5905, n5906, 
      n5907, n5908, n5910, n5913, n5914, n5915, n5917, n5918, n5919, n5920, 
      n5921, n5923, n5924, n5926, n5927, n5928, n5929, n5930, n5931, n5932, 
      n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, 
      n5943, n5944, n5945, n5946, n5949, n5951, n5953, n5954, n5955, n5956, 
      n5957, n5959, n5960, n5963, n5965, n5966, n5968, n5969, n5970, n5971, 
      n5972, n5973, n5974, n5975, n5976, n5977, n5979, n5980, n5981, n5982, 
      n5983, n5985, n5986, n5988, n5991, n5992, n5993, n5994, n5997, n5998, 
      n5999, n6000, n6001, n6002, n6005, n6007, n6008, n6009, n6010, n6012, 
      n6013, n6014, n6015, n6017, n6018, n6019, n6023, n6026, n6027, n6029, 
      n6030, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, 
      n6041, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, 
      n6052, n6053, n6054, n6056, n6057, n6058, n6062, n6064, n6065, n6066, 
      n6067, n6068, n6071, n6075, n6077, n6078, n6081, n6083, n6087, n6088, 
      n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6097, n6098, n6099, 
      n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, 
      n6112, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6124, 
      n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6133, n6134, n6136, 
      n6137, n6139, n6141, n6142, n6145, n6147, n6148, n6149, n6150, n6152, 
      n6153, n6154, n6156, n6158, n6159, n6160, n6161, n6163, n6164, n6165, 
      n6169, n6170, n6171, n6172, n6173, n6175, n6176, n6177, n6178, n6179, 
      n6180, n6181, n6183, n6184, n6185, n6186, n6187, n6189, n6190, n6191, 
      n6192, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, 
      n6204, n6205, n6206, n6207, n6208, n6211, n6212, n6213, n6214, n6215, 
      n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, 
      n6226, n6227, n6228, n6229, n6231, n6232, n6233, n6234, n6235, n6236, 
      n6241, n6243, n6244, n6245, n6246, n6248, n6252, n6253, n6254, n6257, 
      n6261, n6262, n6263, n6264, n6269, n6270, n6271, n6273, n6274, n6277, 
      n6281, n6282, n6283, n6285, n6286, n6287, n6289, n6291, n6293, n6294, 
      n6295, n6297, n6298, n6300, n6301, n6302, n6303, n6304, n6305, n6306, 
      n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6316, n6317, 
      n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6327, n6328, 
      n6329, n6331, n6332, n6335, n6336, n6337, n6339, n6340, n6341, n6342, 
      n6343, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, 
      n6355, n6357, n6360, n6361, n6363, n6365, n6366, n6368, n6369, n6370, 
      n6371, n6372, n6373, n6374, n6375, n6376, n6379, n6381, n6383, n6384, 
      n6385, n6387, n6388, n6389, n6390, n6392, n6393, n6394, n6395, n6396, 
      n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6405, n6408, n6409, 
      n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, 
      n6420, n6421, n6423, n6424, n6426, n6427, n6428, n6429, n6430, n6431, 
      n6432, n6433, n6435, n6436, n6438, n6440, n6441, n6443, n6445, n6446, 
      n6447, n6448, n6449, n6450, n6451, n6453, n6454, n6455, n6456, n6457, 
      n6458, n6460, n6461, n6462, n6463, n6465, n6466, n6467, n6468, n6469, 
      n6470, n6471, n6472, n6473, n6474, n6475, n6477, n6478, n6479, n6480, 
      n6481, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, 
      n6492, n6493, n6496, n6497, n6498, n6499, n6500, n6501, n6503, n6504, 
      n6505, n6506, n6507, n6508, n6509, n6511, n6512, n6513, n6514, n6515, 
      n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6525, n6526, 
      n6527, n6528, n6530, n6531, n6533, n6534, n6535, n6536, n6537, n6539, 
      n6540, n6541, n6542, n6543, n6544, n6546, n6548, n6549, n6550, n6554, 
      n6555, n6556, n6557, n6559, n6560, n6561, n6562, n6563, n6564, n6567, 
      n6569, n6570, n6571, n6572, n6573, n6574, n6576, n6578, n6579, n6580, 
      n6581, n6582, n6583, n6585, n6586, n6587, n6588, n6589, n6590, n6591, 
      n6592, n6593, n6595, n6596, n6598, n6599, n6600, n6601, n6602, n6604, 
      n6605, n6606, n6608, n6609, n6610, n6611, n6615, n6619, n6622, n6623, 
      n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6632, n6633, n6634, 
      n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, 
      n6645, n6646, n6647, n6648, n6649, n6650, n6652, n6654, n6656, n6657, 
      n6658, n6661, n6668, n6669, n6670, n6671, n6672, n6674, n6675, n6676, 
      n6677, n6681, n6684, n6686, n6687, n6688, n6689, n6690, n6691, n6692, 
      n6693, n6694, n6696, n6697, n6698, n6703, n6706, n6707, n6709, n6710, 
      n6711, n6712, n6713, n6714, n6715, n6717, n6719, n6720, n6721, n6722, 
      n6723, n6724, n6727, n6728, n6729, n6731, n6732, n6733, n6734, n6739, 
      n6741, n6744, n6746, n6747, n6748, n6749, n6751, n6752, n6753, n6756, 
      n6757, n6758, n6759, n6762, n6763, n6764, n6765, n6768, n6770, n6771, 
      n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6780, n6781, n6782, 
      n6783, n6784, n6785, n6786, n6788, n6789, n6790, n6791, n6795, n6796, 
      n6797, n6799, n6800, n6801, n6802, n6803, n6807, n6808, n6809, n6810, 
      n6817, n6818, n6819, n6822, n6825, n6826, n6827, n6830, n6831, n6834, 
      n6835, n6836, n6837, n6838, n6839, n6841, n6842, n6843, n6844, n6845, 
      n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6860, 
      n6862, n6863, n6864, n6865, n6866, n6874, n6875, n6876, n6877, n6878, 
      n6879, n6880, n6881, n6883, n6885, n6886, n6887, n6891, n6892, n6893, 
      n6894, n6895, n6896, n6898, n6900, n6901, n6902, n6903, n6904, n6905, 
      n6906, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6916, n6917, 
      n6919, n6920, n6921, n6922, n6923, n6924, n6926, n6927, n6930, n6932, 
      n6933, n6934, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, 
      n6946, n6947, n6948, n6949, n6951, n6952, n6953, n6954, n6955, n6956, 
      n6957, n6960, n6963, n6965, n6969, n6970, n6972, n6975, n6977, n6978, 
      n6980, n6981, n6982, n6984, n6985, n6986, n6987, n6988, n6989, n6990, 
      n6991, n6992, n6993, n6994, n6996, n6997, n6998, n6999, n7000, n7001, 
      n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, 
      n7012, n7013, n7014, n7015, n7017, n7018, n7022, n7023, n7024, n7025, 
      n7026, n7028, n7030, n7031, n7032, n7033, n7034, n7036, n7037, n7038, 
      n7039, n7040, n7041, n7042, n7044, n7046, n7047, n7048, n7049, n7052, 
      n7055, n7056, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, 
      n7066, n7067, n7068, n7069, n7070, n7071, n7075, n7076, n7079, n7080, 
      n7081, n7082, n7083, n7084, n7085, n7086, n7088, n7089, n7090, n7093, 
      n7096, n7097, n7099, n7100, n7101, n7102, n7104, n7105, n7106, n7107, 
      n7108, n7110, n7111, n7112, n7113, n7114, n7115, n7118, n7119, n7120, 
      n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, 
      n7133, n7134, n7135, n7136, n7137, n7140, n7141, n7144, n7145, n7146, 
      n7148, n7149, n7150, n7152, n7153, n7154, n7158, n7160, n7161, n7162, 
      n7163, n7164, n7166, n7167, n7168, n7170, n7171, n7173, n7175, n7176, 
      n7177, n7179, n7180, n7182, n7183, n7185, n7186, n7190, n7191, n7193, 
      n7194, n7195, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7206, 
      n7207, n7208, n7209, n7210, n7212, n7216, n7219, n7220, n7221, n7223, 
      n7224, n7225, n7227, n7230, n7231, n7232, n7234, n7235, n7236, n7237, 
      n7238, n7239, n7240, n7241, n7242, n7243, n7245, n7247, n7248, n7250, 
      n7251, n7252, n7253, n7255, n7256, n7257, n7258, n7260, n7261, n7263, 
      n7265, n7266, n7267, n7270, n7271, n7273, n7275, n7276, n7277, n7278, 
      n7279, n7281, n7282, n7284, n7286, n7287, n7288, n7291, n7292, n7293, 
      n7294, n7295, n7296, n7300, n7302, n7303, n7304, n7305, n7309, n7310, 
      n7312, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7323, n7324, 
      n7325, n7326, n7327, n7328, n7329, n7333, n7335, n7337, n7339, n7341, 
      n7342, n7344, n7345, n7346, n7349, n7350, n7352, n7353, n7355, n7357, 
      n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, 
      n7369, n7370, n7371, n7373, n7374, n7376, n7377, n7379, n7380, n7382, 
      n7384, n7387, n7389, n7391, n7392, n7393, n7396, n7397, n7399, n7402, 
      n7403, n7404, n7406, n7409, n7414, n7415, n7416, n7418, n7423, n7424, 
      n7425, n7426, n7427, n7428, n7429, n7431, n7432, n7434, n7435, n7436, 
      n7437, n7439, n7440, n7443, n7445, n7448, n7451, n7454, n7457, n7459, 
      n7460, n7462, n7464, n7466, n7467, n7468, n7469, n7471, n7472, n7474, 
      n7475, n7478, n7479, n7480, n7481, n7482, n7483, n7485, n7486, n7487, 
      n7488, n7489, n7490, n7491, n7492, n7494, n7495, n7496, n7497, n7498, 
      n7499, n7500, n7502, n7504, n7506, n7507, n7510, n7511, n7512, n7513, 
      n7515, n7516, n7517, n7518, n7520, n7523, n7526, n7527, n7528, n7529, 
      n7530, n7534, n7535, n7536, n7537, n7539, n7540, n7541, n7542, n7543, 
      n7544, n7546, n7547, n7548, n7549, n7551, n7552, n7553, n7555, n7558, 
      n7560, n7564, n7565, n7569, n7570, n7571, n7572, n7573, n7575, n7577, 
      n7578, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, 
      n7591, n7593, n7595, n7596, n7598, n7600, n7601, n7602, n7603, n7606, 
      n7607, n7608, n7610, n7611, n7612, n7613, n7614, n7615, n7619, n7620, 
      n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, 
      n7635, n7636, n7637, n7639, n7640, n7643, n7644, n7647, n7651, n7654, 
      n7657, n7658, n7659, n7660, n7661, n7663, n7664, n7665, n7666, n7667, 
      n7673, n7674, n7676, n7677, n7678, n7680, n7681, n7683, n7689, n7690, 
      n7691, n7693, n7694, n7695, n7696, n7698, n7699, n7703, n7705, n7706, 
      n7708, n7710, n7712, n7714, n7716, n7717, n7718, n7719, n7720, n7722, 
      n7724, n7725, n7726, n7728, n7729, n7730, n7732, n7733, n7734, n7737, 
      n7741, n7742, n7744, n7745, n7749, n7751, n7752, n7755, n7757, n7759, 
      n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, 
      n7772, n7773, n7778, n7779, n7780, n7781, n7783, n7785, n7786, n7787, 
      n7789, n7790, n7792, n7795, n7796, n7797, n7799, n7800, n7801, n7802, 
      n7804, n7805, n7806, n7808, n7810, n7811, n7812, n7813, n7814, n7815, 
      n7816, n7817, n7818, n7819, n7820, n7825, n7828, n7829, n7830, n7831, 
      n7832, n7833, n7834, n7835, n7839, n7840, n7843, n7845, n7846, n7847, 
      n7848, n7849, n7851, n7852, n7853, n7854, n7855, n7859, n7861, n7862, 
      n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7874, 
      n7875, n7876, n7877, n7878, n7880, n7882, n7883, n7884, n7885, n7886, 
      n7888, n7890, n7892, n7893, n7894, n7895, n7896, n7897, n7899, n7900, 
      n7901, n7902, n7904, n7905, n7907, n7908, n7910, n7911, n7912, n7913, 
      n7914, n7915, n7916, n7917, n7919, n7920, n7921, n7922, n7923, n7924, 
      n7926, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7938, 
      n7939, n7941, n7942, n7944, n7945, n7946, n7949, n7950, n7954, n7955, 
      n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, 
      n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, 
      n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7986, n7987, n7989, 
      n7990, n7992, n7993, n7998, n7999, n8000, n8002, n8003, n8005, n8006, 
      n8008, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8019, 
      n8020, n8021, n8023, n8026, n8027, n8028, n8029, n8030, n8031, n8032, 
      n8033, n8034, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8045, 
      n8046, n8048, n8050, n8052, n8053, n8054, n8056, n8057, n8058, n8059, 
      n8060, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, 
      n8071, n8073, n8074, n8075, n8076, n8078, n8080, n8082, n8083, n8085, 
      n8087, n8089, n8090, n8092, n8093, n8094, n8096, n8100, n8101, n8103, 
      n8105, n8106, n8107, n8108, n8109, n8110, n8112, n8113, n8116, n8118, 
      n8119, n8120, n8121, n8122, n8123, n8125, n8127, n8128, n8131, n8132, 
      n8133, n8135, n8136, n8137, n8138, n8139, n8141, n8142, n8143, n8144, 
      n8145, n8146, n8147, n8148, n8149, n8151, n8154, n8155, n8156, n8157, 
      n8158, n8159, n8160, n8161, n8163, n8165, n8166, n8168, n8169, n8171, 
      n8172, n8173, n8174, n8175, n8176, n8177, n8180, n8181, n8182, n8183, 
      n8184, n8186, n8187, n8188, n8189, n8190, n8193, n8194, n8196, n8197, 
      n8199, n8200, n8201, n8202, n8204, n8205, n8206, n8207, n8208, n8210, 
      n8211, n8212, n8213, n8214, n8216, n8217, n8218, n8219, n8221, n8222, 
      n8223, n8228, n8229, n8231, n8232, n8233, n8234, n8235, n8236, n8238, 
      n8239, n8240, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, 
      n8250, n8251, n8252, n8253, n8255, n8257, n8260, n8261, n8262, n8263, 
      n8264, n8265, n8267, n8268, n8269, n8272, n8275, n8276, n8277, n8280, 
      n8281, n8283, n8284, n8285, n8286, n8287, n8289, n8290, n8291, n8293, 
      n8294, n8295, n8296, n8298, n8299, n8300, n8301, n8302, n8303, n8304, 
      n8305, n8307, n8308, n8310, n8311, n8312, n8313, n8314, n8315, n8316, 
      n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, 
      n8327, n8328, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, 
      n8339, n8340, n8342, n8343, n8345, n8346, n8347, n8348, n8349, n8350, 
      n8351, n8355, n8358, n8359, n8360, n8361, n8362, n8364, n8365, n8366, 
      n8368, n8369, n8370, n8371, n8372, n8375, n8376, n8377, n8380, n8381, 
      n8382, n8383, n8384, n8385, n8386, n8388, n8389, n8390, n8392, n8393, 
      n8395, n8396, n8397, n8399, n8400, n8401, n8402, n8403, n8404, n8406, 
      n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8415, n8416, n8419, 
      n8423, n8424, n8425, n8426, n8428, n8430, n8431, n8432, n8434, n8436, 
      n8438, n8439, n8440, n8441, n8442, n8443, n8445, n8446, n8447, n8449, 
      n8452, n8453, n8454, n8458, n8459, n8460, n8461, n8462, n8463, n8465, 
      n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, 
      n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8485, n8486, 
      n8491, n8493, n8494, n8495, n8496, n8498, n8499, n8500, n8501, n8502, 
      n8503, n8504, n8505, n8506, n8507, n8508, n8511, n8512, n8514, n8515, 
      n8516, n8517, n8518, n8519, n8520, n8522, n8523, n8524, n8525, n8526, 
      n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8537, 
      n8538, n8539, n8540, n8542, n8543, n8544, n8546, n8547, n8549, n8552, 
      n8553, n8554, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, 
      n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8574, n8575, n8576, 
      n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, 
      n8590, n8591, n8592, n8593, n8594, n8595, n8597, n8598, n8599, n8600, 
      n8601, n8602, n8604, n8605, n8606, n8607, n8608, n8618, n8621, n8622, 
      n8623, n8625, n8626, n8627, n8628, n8629, n8631, n8632, n8634, n8635, 
      n8637, n8640, n8641, n8642, n8644, n8645, n8646, n8647, n8648, n8649, 
      n8650, n8651, n8652, n8653, n8654, n8656, n8657, n8658, n8659, n8660, 
      n8662, n8666, n8668, n8670, n8671, n8673, n8674, n8676, n8677, n8678, 
      n8679, n8680, n8681, n8682, n8683, n8685, n8686, n8687, n8688, n8689, 
      n8690, n8691, n8692, n8693, n8694, n8696, n8697, n8698, n8699, n8700, 
      n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, 
      n8711, n8713, n8714, n8716, n8717, n8719, n8720, n8721, n8723, n8726, 
      n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, 
      n8737, n8738, n8739, n8741, n8742, n8743, n8744, n8745, n8746, n8747, 
      n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8757, n8758, 
      n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8769, n8770, 
      n8771, n8773, n8774, n8775, n8776, n8780, n8781, n8782, n8784, n8785, 
      n8787, n8788, n8792, n8793, n8794, n8796, n8798, n8799, n8800, n8801, 
      n8803, n8804, n8805, n8806, n8809, n8812, n8814, n8815, n8816, n8817, 
      n8818, n8819, n8820, n8822, n8824, n8825, n8826, n8830, n8833, n8839, 
      n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8849, n8850, 
      n8852, n8853, n8854, n8856, n8858, n8860, n8863, n8865, n8869, n8873, 
      n8874, n8875, n8878, n8879, n8880, n8882, n8883, n8884, n8885, n8887, 
      n8888, n8889, n8890, n8891, n8892, n8894, n8896, n8897, n8898, n8899, 
      n8900, n8901, n8902, n8904, n8905, n8906, n8907, n8908, n8909, n8910, 
      n8911, n8913, n8914, n8916, n8917, n8918, n8919, n8920, n8922, n8923, 
      n8924, n8925, n8927, n8928, n8929, n8931, n8932, n8933, n8934, n8936, 
      n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8946, n8947, 
      n8948, n8949, n8950, n8951, n8952, n8954, n8955, n8957, n8958, n8960, 
      n8961, n8963, n8964, n8965, n8966, n8968, n8969, n8970, n8971, n8972, 
      n8974, n8975, n8977, n8978, n8979, n8980, n8982, n8983, n8985, n8986, 
      n8987, n8988, n8989, n8990, n8993, n8996, n8999, n9000, n9001, n9003, 
      n9005, n9007, n9008, n9009, n9010, n9011, n9013, n9014, n9015, n9016, 
      n9017, n9018, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, 
      n9028, n9029, n9030, n9031, n9032, n9033, n9035, n9036, n9037, n9038, 
      n9039, n9040, n9041, n9043, n9044, n9045, n9046, n9047, n9048, n9049, 
      n9050, n9053, n9054, n9056, n9058, n9059, n9060, n9061, n9062, n9063, 
      n9064, n9066, n9068, n9071, n9073, n9074, n9075, n9077, n9078, n9080, 
      n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9089, n9091, n9092, 
      n9093, n9094, n9095, n9098, n9099, n9101, n9102, n9103, n9104, n9105, 
      n9106, n9107, n9108, n9109, n9111, n9112, n9113, n9114, n9115, n9116, 
      n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, 
      n9127, n9129, n9131, n9132, n9133, n9135, n9137, n9139, n9140, n9141, 
      n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9151, n9152, 
      n9153, n9154, n9155, n9156, n9159, n9160, n9161, n9162, n9164, n9165, 
      n9166, n9168, n9169, n9170, n9173, n9174, n9175, n9176, n9177, n9178, 
      n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9187, n9188, n9190, 
      n9192, n9193, n9195, n9196, n9197, n9198, n9200, n9201, n9202, n9203, 
      n9204, n9205, n9206, n9207, n9209, n9211, n9212, n9213, n9214, n9217, 
      n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, 
      n9228, n9230, n9231, n9233, n9235, n9236, n9237, n9238, n9239, n9240, 
      n9241, n9242, n9243, n9244, n9246, n9247, n9248, n9249, n9250, n9251, 
      n9252, n9253, n9255, n9256, n9257, n9261, n9263, n9264, n9265, n9266, 
      n9267, n9268, n9269, n9270, n9271, n9272, n9274, n9275, n9276, n9277, 
      n9278, n9280, n9286, n9287, n9288, n9290, n9292, n9293, n9294, n9295, 
      n9297, n9298, n9299, n9300, n9301, n9303, n9305, n9308, n9309, n9310, 
      n9312, n9313, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, 
      n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9333, n9334, 
      n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, 
      n9346, n9347, n9349, n9350, n9352, n9353, n9355, n9357, n9360, n9362, 
      n9363, n9364, n9366, n9367, n9369, n9370, n9371, n9373, n9374, n9375, 
      n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, 
      n9387, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9398, n9400, 
      n9401, n9404, n9405, n9408, n9409, n9410, n9411, n9412, n9413, n9415, 
      n9416, n9417, n9418, n9420, n9422, n9423, n9424, n9425, n9427, n9429, 
      n9430, n9431, n9435, n9436, n9438, n9439, n9440, n9441, n9442, n9443, 
      n9444, n9445, n9446, n9448, n9449, n9452, n9454, n9456, n9457, n9458, 
      n9459, n9460, n9461, n9466, n9468, n9469, n9470, n9472, n9474, n9478, 
      n9479, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, 
      n9490, n9491, n9493, n9495, n9496, n9497, n9499, n9500, n9501, n9503, 
      n9504, n9506, n9507, n9508, n9509, n9511, n9512, n9513, n9514, n9516, 
      n9518, n9519, n9520, n9521, n9523, n9524, n9526, n9528, n9529, n9530, 
      n9534, n9535, n9539, n9540, n9541, n9543, n9546, n9547, n9548, n9549, 
      n9550, n9552, n9553, n9554, n9555, n9557, n9559, n9563, n9564, n9565, 
      n9567, n9568, n9569, n9570, n9572, n9573, n9575, n9576, n9577, n9578, 
      n9579, n9580, n9581, n9583, n9584, n9585, n9586, n9587, n9588, n9589, 
      n9590, n9591, n9592, n9593, n9594, n9595, n9597, n9598, n9599, n9602, 
      n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9614, 
      n9616, n9618, n9619, n9621, n9624, n9625, n9626, n9627, n9632, n9633, 
      n9634, n9636, n9638, n9639, n9642, n9643, n9646, n9648, n9649, n9650, 
      n9651, n9654, n9655, n9656, n9658, n9660, n9663, n9667, n9668, n9669, 
      n9670, n9672, n9673, n9674, n9676, n9677, n9680, n9682, n9683, n9684, 
      n9685, n9686, n9687, n9688, n9690, n9692, n9694, n9695, n9698, n9699, 
      n9700, n9701, n9702, n9703, n9705, n9707, n9708, n9711, n9712, n9714, 
      n9715, n9716, n9719, n9721, n9722, n9723, n9725, n9726, n9727, n9731, 
      n9732, n9733, n9734, n9735, n9736, n9737, n9739, n9740, n9743, n9745, 
      n9746, n9748, n9751, n9756, n9757, n9758, n9759, n9762, n9763, n9764, 
      n9766, n9768, n9769, n9770, n9772, n9775, n9776, n9777, n9780, n9781, 
      n9783, n9786, n9787, n9788, n9790, n9791, n9794, n9795, n9796, n9797, 
      n9798, n9799, n9800, n9801, n9802, n9803, n9805, n9806, n9807, n9808, 
      n9809, n9811, n9813, n9815, n9816, n9817, n9818, n9821, n9822, n9823, 
      n9824, n9825, n9826, n9828, n9829, n9833, n9835, n9836, n9837, n9838, 
      n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, 
      n9849, n9850, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, 
      n9861, n9862, n9863, n9865, n9868, n9869, n9870, n9872, n9873, n9874, 
      n9875, n9876, n9878, n9880, n9882, n9883, n9884, n9885, n9886, n9887, 
      n9888, n9889, n9891, n9892, n9893, n9894, n9895, n9897, n9899, n9900, 
      n9903, n9904, n9907, n9909, n9911, n9912, n9913, n9914, n9915, n9916, 
      n9917, n9918, n9920, n9921, n9922, n9923, n9924, n9926, n9928, n9930, 
      n9931, n9932, n9935, n9937, n9938, n9939, n9941, n9942, n9943, n9944, 
      n9945, n9947, n9948, n9951, n9952, n9953, n9954, n9955, n9956, n9957, 
      n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9967, n9968, n9969, 
      n9970, n9971, n9972, n9973, n9975, n9976, n9977, n9979, n9980, n9981, 
      n9982, n9983, n9984, n9986, n9987, n9988, n9989, n9990, n9991, n9992, 
      n9993, n9994, n9996, n9997, n9999, n10001, n10002, n10003, n10004, n10006
      , n10008, n10009, n10012, n10013, n10014, n10015, n10016, n10018, n10019,
      n10023, n10024, n10025, n10026, n10027, n10029, n10030, n10031, n10032, 
      n10034, n10036, n10037, n10038, n10039, n10040, n10041, n10044, n10046, 
      n10047, n10048, n10050, n10051, n10052, n10054, n10055, n10056, n10057, 
      n10058, n10059, n10061, n10062, n10065, n10066, n10069, n10070, n10071, 
      n10073, n10074, n10076, n10078, n10079, n10080, n10081, n10082, n10083, 
      n10084, n10085, n10087, n10089, n10092, n10096, n10097, n10098, n10100, 
      n10101, n10104, n10107, n10109, n10110, n10111, n10112, n10113, n10114, 
      n10115, n10116, n10117, n10118, n10120, n10122, n10123, n10125, n10126, 
      n10127, n10128, n10129, n10131, n10132, n10134, n10136, n10137, n10138, 
      n10139, n10140, n10141, n10143, n10144, n10146, n10147, n10148, n10150, 
      n10151, n10152, n10153, n10154, n10155, n10156, n10158, n10159, n10160, 
      n10161, n10162, n10163, n10166, n10167, n10168, n10169, n10171, n10174, 
      n10176, n10177, n10179, n10180, n10181, n10182, n10183, n10185, n10186, 
      n10187, n10189, n10190, n10193, n10195, n10196, n10197, n10199, n10200, 
      n10201, n10202, n10203, n10204, n10205, n10207, n10208, n10209, n10210, 
      n10211, n10212, n10213, n10214, n10215, n10216, n10219, n10220, n10221, 
      n10223, n10224, n10225, n10226, n10228, n10230, n10231, n10233, n10234, 
      n10236, n10237, n10239, n10240, n10242, n10243, n10244, n10245, n10246, 
      n10247, n10248, n10250, n10251, n10252, n10253, n10254, n10255, n10256, 
      n10258, n10259, n10261, n10263, n10266, n10267, n10268, n10269, n10270, 
      n10272, n10273, n10275, n10276, n10278, n10279, n10282, n10284, n10287, 
      n10288, n10289, n10290, n10292, n10293, n10294, n10295, n10296, n10297, 
      n10299, n10301, n10302, n10303, n10304, n10305, n10309, n10312, n10313, 
      n10314, n10315, n10316, n10317, n10318, n10319, n10321, n10323, n10324, 
      n10325, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10336, 
      n10337, n10338, n10340, n10342, n10343, n10345, n10346, n10349, n10351, 
      n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10361, 
      n10364, n10365, n10366, n10369, n10370, n10371, n10373, n10374, n10375, 
      n10377, n10378, n10379, n10380, n10382, n10383, n10384, n10385, n10386, 
      n10387, n10388, n10389, n10390, n10391, n10393, n10394, n10396, n10399, 
      n10400, n10401, n10402, n10403, n10404, n10406, n10407, n10408, n10409, 
      n10410, n10412, n10413, n10414, n10417, n10418, n10419, n10420, n10421, 
      n10422, n10424, n10426, n10427, n10428, n10429, n10430, n10431, n10432, 
      n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, 
      n10442, n10443, n10444, n10447, n10451, n10452, n10455, n10457, n10458, 
      n10461, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, 
      n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, 
      n10480, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10491, 
      n10492, n10493, n10494, n10495, n10498, n10501, n10502, n10507, n10508, 
      n10509, n10510, n10511, n10513, n10515, n10516, n10518, n10519, n10520, 
      n10521, n10523, n10524, n10525, n10526, n10530, n10532, n10534, n10535, 
      n10536, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10546, 
      n10548, n10549, n10551, n10552, n10553, n10555, n10556, n10558, n10559, 
      n10560, n10561, n10562, n10563, n10564, n10565, n10567, n10568, n10569, 
      n10570, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, 
      n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10589, n10590, 
      n10592, n10593, n10595, n10596, n10597, n10598, n10599, n10605, n10606, 
      n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, 
      n10619, n10620, n10621, n10622, n10623, n10626, n10628, n10629, n10630, 
      n10631, n10632, n10633, n10634, n10635, n10636, n10638, n10640, n10642, 
      n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, 
      n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10662, n10663, 
      n10665, n10667, n10668, n10670, n10671, n10673, n10674, n10676, n10677, 
      n10678, n10679, n10680, n10681, n10683, n10684, n10685, n10686, n10689, 
      n10690, n10691, n10693, n10694, n10695, n10697, n10698, n10699, n10702, 
      n10703, n10705, n10706, n10707, n10708, n10709, n10711, n10712, n10713, 
      n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, 
      n10723, n10724, n10729, n10731, n10733, n10734, n10735, n10736, n10737, 
      n10739, n10742, n10743, n10744, n10746, n10747, n10748, n10751, n10753, 
      n10754, n10755, n10756, n10757, n10758, n10762, n10763, n10764, n10765, 
      n10766, n10767, n10769, n10770, n10771, n10773, n10774, n10775, n10776, 
      n10777, n10779, n10782, n10783, n10784, n10785, n10786, n10787, n10788, 
      n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, 
      n10800, n10801, n10803, n10806, n10807, n10810, n10811, n10812, n10813, 
      n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, 
      n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, 
      n10832, n10834, n10835, n10836, n10837, n10839, n10840, n10841, n10842, 
      n10845, n10846, n10847, n10848, n10850, n10853, n10854, n10855, n10856, 
      n10857, n10858, n10859, n10860, n10862, n10863, n10864, n10866, n10867, 
      n10868, n10869, n10870, n10872, n10874, n10875, n10876, n10878, n10882, 
      n10883, n10884, n10885, n10887, n10888, n10889, n10890, n10891, n10893, 
      n10894, n10896, n10897, n10898, n10899, n10901, n10902, n10903, n10904, 
      n10905, n10906, n10907, n10908, n10910, n10913, n10914, n10915, n10918, 
      n10920, n10924, n10925, n10926, n10928, n10929, n10930, n10931, n10935, 
      n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10946, 
      n10949, n10953, n10955, n10957, n10959, n10961, n10962, n10963, n10965, 
      n10966, n10967, n10969, n10970, n10971, n10972, n10973, n10974, n10976, 
      n10977, n10978, n10979, n10980, n10982, n10983, n10984, n10986, n10987, 
      n10988, n10989, n10992, n10996, n10997, n10998, n10999, n11001, n11003, 
      n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11012, n11013, 
      n11015, n11016, n11017, n11018, n11020, n11022, n11024, n11025, n11026, 
      n11028, n11030, n11031, n11032, n11033, n11034, n11036, n11037, n11038, 
      n11039, n11040, n11041, n11042, n11043, n11044, n11046, n11047, n11048, 
      n11050, n11053, n11054, n11055, n11056, n11057, n11059, n11060, n11061, 
      n11062, n11063, n11064, n11065, n11066, n11067, n11072, n11074, n11075, 
      n11076, n11077, n11081, n11082, n11083, n11084, n11087, n11088, n11089, 
      n11090, n11091, n11092, n11094, n11095, n11097, n11098, n11099, n11102, 
      n11103, n11104, n11105, n11108, n11111, n11114, n11115, n11116, n11117, 
      n11118, n11119, n11120, n11121, n11124, n11125, n11126, n11127, n11128, 
      n11129, n11130, n11131, n11132, n11133, n11134, n11136, n11137, n11138, 
      n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, 
      n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, 
      n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, 
      n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11180, n11181, 
      n11182, n11183, n11185, n11186, n11187, n11188, n11189, n11190, n11192, 
      n11194, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11207, 
      n11208, n11210, n11211, n11213, n11214, n11215, n11217, n11218, n11219, 
      n11220, n11222, n11224, n11225, n11226, n11227, n11230, n11233, n11234, 
      n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11243, n11245, 
      n11247, n11248, n11250, n11251, n11252, n11253, n11254, n11255, n11256, 
      n11257, n11258, n11260, n11261, n11263, n11264, n11265, n11266, n11267, 
      n11268, n11269, n11270, n11271, n11274, n11275, n11276, n11277, n11278, 
      n11279, n11280, n11283, n11284, n11286, n11288, n11289, n11290, n11291, 
      n11292, n11293, n11295, n11296, n11297, n11298, n11299, n11300, n11301, 
      n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, 
      n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, 
      n11321, n11322, n11323, n11325, n11327, n11328, n11329, n11330, n11331, 
      n11332, n11333, n11334, n11335, n11336, n11337, n11339, n11342, n11344, 
      n11345, n11346, n11347, n11348, n11349, n11350, n11353, n11354, n11355, 
      n11356, n11358, n11361, n11363, n11364, n11365, n11366, n11367, n11368, 
      n11369, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, 
      n11382, n11383, n11384, n11386, n11387, n11388, n11389, n11390, n11391, 
      n11392, n11394, n11395, n11397, n11398, n11399, n11401, n11402, n11404, 
      n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, 
      n11415, n11416, n11417, n11418, n11419, n11421, n11423, n11424, n11425, 
      n11428, n11429, n11431, n11432, n11433, n11434, n11435, n11436, n11437, 
      n11438, n11439, n11440, n11441, n11442, n11443, n11446, n11448, n11449, 
      n11451, n11452, n11453, n11455, n11456, n11458, n11459, n11461, n11462, 
      n11463, n11464, n11465, n11467, n11468, n11469, n11470, n11472, n11473, 
      n11474, n11475, n11476, n11477, n11479, n11481, n11482, n11484, n11485, 
      n11486, n11487, n11488, n11490, n11491, n11492, n11494, n11495, n11496, 
      n11497, n11498, n11500, n11501, n11502, n11503, n11506, n11507, n11508, 
      n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, 
      n11520, n11521, n11522, n11523, n11525, n11526, n11528, n11529, n11530, 
      n11533, n11534, n11536, n11541, n11542, n11543, n11544, n11547, n11548, 
      n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, 
      n11558, n11559, n11560, n11562, n11563, n11564, n11567, n11568, n11569, 
      n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11581, 
      n11582, n11583, n11584, n11585, n11586, n11588, n11589, n11590, n11591, 
      n11594, n11595, n11596, n11597, n11598, n11600, n11601, n11602, n11603, 
      n11605, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, 
      n11617, n11620, n11621, n11622, n11623, n11624, n11625, n11627, n11628, 
      n11630, n11631, n11633, n11634, n11635, n11636, n11637, n11638, n11639, 
      n11641, n11642, n11643, n11644, n11646, n11647, n11648, n11649, n11650, 
      n11651, n11652, n11653, n11657, n11658, n11659, n11661, n11663, n11664, 
      n11665, n11667, n11668, n11669, n11671, n11672, n11673, n11674, n11676, 
      n11677, n11678, n11679, n11680, n11682, n11683, n11684, n11687, n11688, 
      n11689, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, 
      n11702, n11703, n11704, n11705, n11707, n11708, n11709, n11710, n11711, 
      n11712, n11713, n11714, n11717, n11718, n11719, n11721, n11722, n11723, 
      n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11732, n11734, 
      n11735, n11736, n11737, n11738, n11739, n11740, n11742, n11743, n11746, 
      n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, 
      n11756, n11757, n11758, n11759, n11760, n11762, n11763, n11764, n11765, 
      n11767, n11768, n11769, n11770, n11771, n11773, n11776, n11777, n11778, 
      n11779, n11780, n11782, n11783, n11784, n11785, n11787, n11788, n11789, 
      n11790, n11791, n11793, n11794, n11795, n11796, n11797, n11800, n11803, 
      n11805, n11806, n11807, n11809, n11810, n11814, n11818, n11820, n11822, 
      n11823, n11826, n11828, n11830, n11831, n11833, n11834, n11835, n11838, 
      n11842, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, 
      n11853, n11854, n11855, n11856, n11858, n11859, n11860, n11861, n11864, 
      n11866, n11867, n11868, n11869, n11870, n11871, n11873, n11874, n11875, 
      n11876, n11877, n11878, n11880, n11881, n11882, n11883, n11885, n11886, 
      n11887, n11888, n11889, n11890, n11891, n11893, n11895, n11896, n11897, 
      n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, 
      n11907, n11908, n11910, n11911, n11912, n11913, n11914, n11916, n11917, 
      n11918, n11919, n11921, n11922, n11923, n11924, n11925, n11926, n11927, 
      n11935, n11937, n11938, n11939, n11940, n11942, n11943, n11944, n11945, 
      n11946, n11947, n11948, n11950, n11951, n11952, n11954, n11956, n11957, 
      n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, 
      n11969, n11970, n11972, n11973, n11974, n11975, n11976, n11977, n11980, 
      n11981, n11984, n11985, n11986, n11987, n11989, n11994, n11996, n11997, 
      n11998, n11999, n12000, n12001, n12002, n12003, n12008, n12009, n12011, 
      n12012, n12014, n12015, n12016, n12017, n12018, n12020, n12022, n12023, 
      n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, 
      n12033, n12036, n12038, n12039, n12040, n12044, n12045, n12046, n12049, 
      n12050, n12053, n12054, n12055, n12056, n12060, n12061, n12062, n12063, 
      n12064, n12065, n12066, n12067, n12069, n12072, n12073, n12074, n12075, 
      n12076, n12077, n12078, n12079, n12080, n12081, n12083, n12084, n12085, 
      n12086, n12090, n12091, n12093, n12094, n12096, n12097, n12100, n12101, 
      n12102, n12103, n12104, n12105, n12107, n12108, n12109, n12111, n12112, 
      n12113, n12114, n12115, n12118, n12119, n12120, n12121, n12122, n12123, 
      n12124, n12125, n12130, n12131, n12132, n12133, n12138, n12139, n12141, 
      n12142, n12144, n12145, n12146, n12148, n12150, n12151, n12152, n12153, 
      n12154, n12155, n12156, n12157, n12159, n12160, n12161, n12162, n12163, 
      n12165, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, 
      n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12183, n12184, 
      n12185, n12187, n12189, n12191, n12192, n12194, n12195, n12196, n12197, 
      n12198, n12199, n12200, n12202, n12203, n12204, n12205, n12206, n12207, 
      n12208, n12212, n12213, n12214, n12215, n12218, n12220, n12221, n12225, 
      n12227, n12228, n12230, n12231, n12232, n12233, n12234, n12235, n12236, 
      n12237, n12238, n12239, n12240, n12242, n12243, n12244, n12245, n12246, 
      n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12257, 
      n12258, n12259, n12260, n12261, n12262, n12263, n12265, n12266, n12267, 
      n12268, n12269, n12272, n12273, n12275, n12276, n12277, n12279, n12282, 
      n12283, n12286, n12287, n12288, n12289, n12290, n12293, n12296, n12297, 
      n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12306, n12307, 
      n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, 
      n12318, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, 
      n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12336, n12337, 
      n12339, n12340, n12341, n12342, n12343, n12345, n12349, n12350, n12351, 
      n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12360, n12362, 
      n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, 
      n12372, n12373, n12374, n12375, n12377, n12378, n12379, n12381, n12382, 
      n12383, n12385, n12387, n12388, n12391, n12392, n12393, n12394, n12396, 
      n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, 
      n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, 
      n12416, n12417, n12418, n12420, n12422, n12423, n12424, n12425, n12426, 
      n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12435, n12437, 
      n12438, n12439, n12441, n12442, n12443, n12446, n12447, n12448, n12449, 
      n12450, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12460, 
      n12461, n12462, n12463, n12464, n12466, n12468, n12469, n12470, n12471, 
      n12472, n12473, n12475, n12477, n12478, n12479, n12480, n12481, n12485, 
      n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, 
      n12495, n12497, n12498, n12499, n12500, n12503, n12504, n12505, n12507, 
      n12508, n12509, n12510, n12511, n12512, n12513, n12515, n12516, n12517, 
      n12518, n12519, n12520, n12522, n12523, n12524, n12525, n12526, n12527, 
      n12529, n12531, n12533, n12534, n12535, n12537, n12538, n12539, n12540, 
      n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, 
      n12551, n12552, n12553, n12556, n12557, n12558, n12560, n12561, n12562, 
      n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12572, 
      n12574, n12575, n12576, n12578, n12579, n12580, n12586, n12587, n12588, 
      n12590, n12592, n12593, n12594, n12597, n12598, n12599, n12601, n12604, 
      n12605, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12616, 
      n12617, n12618, n12620, n12621, n12622, n12623, n12624, n12625, n12626, 
      n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12638, n12639, 
      n12641, n12642, n12643, n12644, n12646, n12649, n12650, n12651, n12653, 
      n12654, n12655, n12657, n12659, n12660, n12661, n12663, n12664, n12665, 
      n12667, n12669, n12670, n12671, n12672, n12673, n12675, n12676, n12680, 
      n12681, n12682, n12683, n12684, n12685, n12686, n12689, n12690, n12691, 
      n12692, n12694, n12696, n12697, n12698, n12699, n12702, n12703, n12704, 
      n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, 
      n12714, n12715, n12717, n12718, n12721, n12722, n12723, n12726, n12727, 
      n12728, n12729, n12730, n12732, n12733, n12735, n12736, n12737, n12738, 
      n12741, n12744, n12745, n12746, n12748, n12749, n12751, n12752, n12754, 
      n12755, n12756, n12758, n12759, n12760, n12762, n12763, n12765, n12766, 
      n12767, n12768, n12769, n12770, n12771, n12772, n12775, n12776, n12778, 
      n12779, n12780, n12782, n12784, n12785, n12787, n12788, n12790, n12793, 
      n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, 
      n12804, n12805, n12806, n12807, n12808, n12809, n12812, n12813, n12814, 
      n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12824, 
      n12825, n12826, n12828, n12829, n12830, n12832, n12833, n12834, n12835, 
      n12836, n12838, n12839, n12840, n12842, n12844, n12846, n12847, n12848, 
      n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, 
      n12859, n12860, n12861, n12862, n12863, n12865, n12866, n12869, n12870, 
      n12871, n12876, n12878, n12879, n12880, n12882, n12883, n12884, n12885, 
      n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12895, n12896, 
      n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12908, n12909, 
      n12910, n12912, n12914, n12915, n12916, n12918, n12919, n12920, n12921, 
      n12922, n12923, n12924, n12925, n12926, n12927, n12930, n12931, n12933, 
      n12934, n12935, n12936, n12939, n12940, n12941, n12942, n12943, n12944, 
      n12946, n12947, n12950, n12951, n12952, n12953, n12954, n12955, n12960, 
      n12961, n12964, n12966, n12969, n12970, n12971, n12972, n12973, n12974, 
      n12975, n12976, n12978, n12979, n12982, n12983, n12984, n12985, n12986, 
      n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, 
      n12996, n12997, n12999, n13000, n13001, n13002, n13004, n13005, n13006, 
      n13008, n13009, n13010, n13012, n13013, n13014, n13015, n13016, n13018, 
      n13019, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, 
      n13030, n13033, n13034, n13035, n13036, n13038, n13039, n13040, n13042, 
      n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13052, n13053, 
      n13054, n13055, n13056, n13059, n13060, n13061, n13062, n13064, n13065, 
      n13066, n13067, n13068, n13069, n13070, n13072, n13073, n13074, n13075, 
      n13076, n13077, n13078, n13081, n13082, n13083, n13085, n13087, n13088, 
      n13090, n13091, n13093, n13094, n13095, n13096, n13097, n13098, n13099, 
      n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13110, 
      n13111, n13112, n13113, n13114, n13115, n13116, n13118, n13119, n13121, 
      n13123, n13124, n13127, n13128, n13129, n13131, n13132, n13133, n13134, 
      n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, 
      n13147, n13149, n13150, n13151, n13153, n13154, n13155, n13156, n13157, 
      n13158, n13159, n13161, n13163, n13164, n13165, n13166, n13167, n13168, 
      n13170, n13171, n13172, n13174, n13176, n13177, n13178, n13179, n13181, 
      n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, 
      n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13199, n13200, 
      n13201, n13202, n13205, n13206, n13207, n13208, n13210, n13211, n13212, 
      n13213, n13214, n13215, n13217, n13218, n13219, n13220, n13221, n13222, 
      n13223, n13224, n13226, n13227, n13228, n13229, n13231, n13232, n13233, 
      n13234, n13235, n13236, n13237, n13239, n13240, n13241, n13242, n13243, 
      n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, 
      n13254, n13255, n13257, n13258, n13259, n13260, n13261, n13262, n13263, 
      n13264, n13266, n13267, n13268, n13270, n13273, n13274, n13275, n13277, 
      n13278, n13279, n13280, n13281, n13282, n13283, n13285, n13286, n13287, 
      n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, 
      n13298, n13300, n13301, n13302, n13304, n13305, n13306, n13308, n13310, 
      n13311, n13312, n13313, n13315, n13316, n13317, n13318, n13320, n13321, 
      n13322, n13323, n13324, n13326, n13327, n13329, n13332, n13333, n13334, 
      n13335, n13336, n13337, n13339, n13340, n13342, n13345, n13348, n13349, 
      n13350, n13351, n13352, n13354, n13356, n13358, n13359, n13361, n13362, 
      n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, 
      n13372, n13373, n13374, n13375, n13378, n13379, n13381, n13383, n13384, 
      n13386, n13387, n13388, n13389, n13391, n13392, n13393, n13395, n13397, 
      n13398, n13400, n13401, n13403, n13404, n13406, n13407, n13408, n13409, 
      n13410, n13411, n13412, n13413, n13414, n13415, n13417, n13419, n13420, 
      n13421, n13422, n13424, n13425, n13426, n13427, n13428, n13429, n13430, 
      n13431, n13432, n13433, n13437, n13438, n13439, n13440, n13441, n13442, 
      n13443, n13444, n13445, n13446, n13448, n13450, n13451, n13453, n13454, 
      n13455, n13457, n13458, n13460, n13461, n13462, n13465, n13466, n13467, 
      n13468, n13469, n13471, n13472, n13473, n13475, n13476, n13477, n13478, 
      n13479, n13480, n13481, n13483, n13484, n13485, n13487, n13488, n13489, 
      n13491, n13492, n13494, n13495, n13496, n13497, n13498, n13499, n13500, 
      n13501, n13502, n13503, n13504, n13508, n13510, n13512, n13513, n13514, 
      n13515, n13516, n13518, n13519, n13521, n13522, n13523, n13524, n13525, 
      n13526, n13527, n13528, n13530, n13531, n13533, n13534, n13535, n13536, 
      n13537, n13538, n13539, n13540, n13542, n13543, n13544, n13545, n13547, 
      n13548, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, 
      n13558, n13559, n13560, n13561, n13563, n13564, n13565, n13566, n13568, 
      n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13578, n13579, 
      n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, 
      n13589, n13591, n13592, n13593, n13594, n13595, n13596, n13598, n13599, 
      n13600, n13601, n13602, n13603, n13605, n13606, n13607, n13608, n13609, 
      n13610, n13614, n13615, n13616, n13617, n13618, n13620, n13621, n13623, 
      n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, 
      n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, 
      n13642, n13644, n13645, n13646, n13649, n13650, n13652, n13653, n13654, 
      n13656, n13657, n13658, n13663, n13664, n13665, n13666, n13667, n13668, 
      n13669, n13670, n13671, n13672, n13673, n13674, n13677, n13678, n13679, 
      n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13688, n13689, 
      n13690, n13691, n13692, n13694, n13695, n13696, n13697, n13698, n13699, 
      n13700, n13701, n13703, n13704, n13705, n13706, n13707, n13708, n13709, 
      n13710, n13711, n13712, n13713, n13714, n13716, n13717, n13718, n13719, 
      n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, 
      n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13738, n13739, 
      n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, 
      n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, 
      n13759, n13761, n13762, n13763, n13765, n13766, n13767, n13768, n13769, 
      n13770, n13771, n13774, n13775, n13776, n13777, n13778, n13779, n13780, 
      n13782, n13784, n13785, n13786, n13787, n13788, n13789, n13791, n13792, 
      n13793, n13794, n13797, n13799, n13800, n13801, n13802, n13803, n13804, 
      n13805, n13806, n13807, n13808, n13809, n13811, n13814, n13815, n13817, 
      n13818, n13820, n13823, n13824, n13825, n13826, n13827, n13829, n13830, 
      n13831, n13832, n13833, n13834, n13837, n13839, n13840, n13842, n13843, 
      n13844, n13845, n13846, n13847, n13849, n13850, n13851, n13852, n13853, 
      n13854, n13855, n13856, n13858, n13859, n13860, n13861, n13862, n13869, 
      n13870, n13871, n13872, n13873, n13875, n13876, n13877, n13878, n13879, 
      n13880, n13881, n13883, n13884, n13885, n13886, n13890, n13891, n13892, 
      n13893, n13894, n13895, n13896, n13897, n13899, n13900, n13901, n13903, 
      n13904, n13905, n13906, n13907, n13909, n13910, n13911, n13912, n13913, 
      n13914, n13917, n13918, n13919, n13920, n13922, n13926, n13927, n13928, 
      n13931, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13942, 
      n13943, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, 
      n13954, n13955, n13956, n13959, n13961, n13962, n13963, n13964, n13965, 
      n13966, n13967, n13969, n13970, n13971, n13973, n13976, n13977, n13978, 
      n13980, n13981, n13982, n13983, n13984, n13986, n13988, n13989, n13990, 
      n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n14000, 
      n14001, n14002, n14003, n14004, n14006, n14007, n14008, n14009, n14011, 
      n14012, n14015, n14016, n14017, n14020, n14022, n14023, n14024, n14025, 
      n14027, n14028, n14030, n14031, n14034, n14035, n14036, n14037, n14038, 
      n14039, n14041, n14043, n14045, n14046, n14049, n14050, n14051, n14052, 
      n14053, n14056, n14057, n14058, n14060, n14061, n14062, n14063, n14064, 
      n14065, n14066, n14069, n14072, n14073, n14075, n14076, n14079, n14080, 
      n14081, n14082, n14083, n14084, n14085, n14086, n14088, n14089, n14091, 
      n14093, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, 
      n14105, n14106, n14107, n14109, n14110, n14112, n14113, n14115, n14116, 
      n14117, n14118, n14121, n14122, n14123, n14124, n14125, n14126, n14127, 
      n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, 
      n14139, n14140, n14143, n14144, n14145, n14146, n14147, n14148, n14150, 
      n14151, n14152, n14153, n14154, n14156, n14157, n14158, n14160, n14163, 
      n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14173, 
      n14174, n14176, n14178, n14179, n14181, n14183, n14184, n14186, n14187, 
      n14188, n14189, n14191, n14192, n14193, n14194, n14195, n14196, n14197, 
      n14198, n14199, n14200, n14201, n14203, n14205, n14206, n14209, n14211, 
      n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, 
      n14221, n14222, n14224, n14226, n14228, n14229, n14230, n14231, n14232, 
      n14233, n14234, n14235, n14237, n14239, n14241, n14244, n14245, n14248, 
      n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14257, n14258, 
      n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14269, 
      n14270, n14271, n14272, n14273, n14275, n14276, n14277, n14278, n14280, 
      n14281, n14282, n14283, n14285, n14286, n14287, n14289, n14290, n14291, 
      n14292, n14293, n14294, n14295, n14297, n14300, n14302, n14303, n14304, 
      n14305, n14306, n14307, n14309, n14311, n14312, n14316, n14318, n14319, 
      n14322, n14323, n14325, n14326, n14327, n14330, n14331, n14332, n14333, 
      n14337, n14338, n14339, n14343, n14345, n14346, n14347, n14349, n14350, 
      n14351, n14352, n14353, n14354, n14355, n14359, n14361, n14362, n14363, 
      n14364, n14365, n14367, n14369, n14371, n14373, n14374, n14375, n14376, 
      n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14385, n14386, 
      n14387, n14388, n14389, n14390, n14392, n14393, n14394, n14395, n14396, 
      n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, 
      n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, 
      n14417, n14418, n14420, n14421, n14422, n14423, n14424, n14425, n14426, 
      n14427, n14428, n14429, n14431, n14432, n14433, n14435, n14436, n14437, 
      n14438, n14439, n14440, n14442, n14443, n14444, n14448, n14449, n14450, 
      n14451, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, 
      n14461, n14462, n14463, n14469, n14471, n14472, n14473, n14474, n14475, 
      n14476, n14477, n14478, n14480, n14481, n14482, n14483, n14484, n14485, 
      n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, 
      n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, 
      n14504, n14505, n14506, n14507, n14508, n14509, n14511, n14512, n14513, 
      n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, 
      n14524, n14525, n14526, n14527, n14529, n14530, n14532, n14533, n14534, 
      n14535, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14546, 
      n14548, n14549, n14551, n14553, n14556, n14557, n14558, n14559, n14560, 
      n14561, n14562, n14563, n14564, n14565, n14566, n14568, n14569, n14571, 
      n14572, n14573, n14576, n14577, n14578, n14579, n14581, n14582, n14583, 
      n14585, n14586, n14587, n14588, n14589, n14590, n14592, n14593, n14594, 
      n14596, n14597, n14600, n14601, n14602, n14603, n14604, n14605, n14606, 
      n14608, n14609, n14610, n14613, n14614, n14615, n14617, n14618, n14619, 
      n14621, n14622, n14623, n14625, n14626, n14628, n14630, n14631, n14632, 
      n14634, n14635, n14636, n14638, n14639, n14640, n14641, n14642, n14643, 
      n14644, n14645, n14646, n14648, n14649, n14650, n14651, n14652, n14654, 
      n14655, n14656, n14657, n14658, n14659, n14660, n14662, n14664, n14665, 
      n14666, n14667, n14668, n14669, n14670, n14672, n14673, n14675, n14677, 
      n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, 
      n14689, n14691, n14692, n14693, n14694, n14695, n14696, n14699, n14701, 
      n14703, n14704, n14705, n14708, n14709, n14712, n14713, n14715, n14716, 
      n14717, n14718, n14719, n14720, n14721, n14722, n14724, n14725, n14729, 
      n14732, n14734, n14735, n14736, n14737, n14738, n14739, n14742, n14743, 
      n14744, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14754, 
      n14755, n14756, n14757, n14758, n14759, n14760, n14762, n14764, n14765, 
      n14766, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14777, 
      n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14787, n14788, 
      n14789, n14790, n14791, n14793, n14794, n14795, n14796, n14797, n14798, 
      n14800, n14801, n14802, n14804, n14805, n14807, n14808, n14810, n14811, 
      n14813, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, 
      n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14833, 
      n14834, n14835, n14837, n14838, n14839, n14840, n14843, n14844, n14845, 
      n14846, n14848, n14850, n14851, n14854, n14855, n14856, n14857, n14858, 
      n14859, n14861, n14862, n14866, n14867, n14868, n14869, n14872, n14873, 
      n14874, n14875, n14876, n14877, n14879, n14880, n14881, n14882, n14887, 
      n14888, n14890, n14891, n14892, n14894, n14895, n14896, n14897, n14898, 
      n14899, n14900, n14901, n14902, n14903, n14904, n14907, n14908, n14909, 
      n14910, n14911, n14912, n14914, n14915, n14916, n14919, n14920, n14921, 
      n14922, n14924, n14925, n14926, n14927, n14928, n14929, n14931, n14933, 
      n14934, n14935, n14936, n14939, n14940, n14941, n14945, n14946, n14947, 
      n14949, n14952, n14953, n14955, n14956, n14957, n14962, n14966, n14967, 
      n14968, n14969, n14970, n14971, n14974, n14977, n14978, n14979, n14980, 
      n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, 
      n14990, n14991, n14993, n14994, n14995, n14997, n14998, n14999, n15001, 
      n15003, n15004, n15005, n15006, n15007, n15009, n15010, n15011, n15012, 
      n15013, n15014, n15015, n15017, n15018, n15019, n15020, n15021, n15022, 
      n15023, n15024, n15026, n15027, n15028, n15029, n15030, n15031, n15032, 
      n15033, n15034, n15036, n15037, n15038, n15039, n15040, n15041, n15042, 
      n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, 
      n15052, n15053, n15056, n15058, n15062, n15063, n15068, n15069, n15071, 
      n15072, n15073, n15074, n15075, n15077, n15078, n15079, n15080, n15081, 
      n15082, n15084, n15085, n15087, n15089, n15090, n15091, n15093, n15094, 
      n15096, n15097, n15099, n15102, n15109, n15110, n15112, n15113, n15114, 
      n15115, n15118, n15120, n15121, n15122, n15123, n15124, n15125, n15126, 
      n15127, n15128, n15131, n15132, n15134, n15135, n15136, n15137, n15138, 
      n15139, n15140, n15141, n15142, n15143, n15145, n15146, n15148, n15149, 
      n15151, n15152, n15153, n15155, n15156, n15157, n15158, n15159, n15160, 
      n15162, n15163, n15164, n15165, n15168, n15169, n15171, n15172, n15173, 
      n15174, n15175, n15176, n15177, n15178, n15180, n15181, n15183, n15184, 
      n15186, n15187, n15189, n15193, n15194, n15195, n15196, n15197, n15199, 
      n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15208, n15209, 
      n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15218, n15219, 
      n15220, n15222, n15223, n15224, n15226, n15227, n15229, n15230, n15232, 
      n15233, n15235, n15237, n15238, n15239, n15240, n15242, n15243, n15245, 
      n15246, n15248, n15249, n15250, n15251, n15254, n15256, n15257, n15258, 
      n15259, n15261, n15265, n15266, n15267, n15268, n15269, n15270, n15271, 
      n15272, n15273, n15274, n15275, n15276, n15277, n15280, n15281, n15282, 
      n15283, n15284, n15286, n15287, n15288, n15289, n15290, n15292, n15293, 
      n15294, n15295, n15296, n15298, n15299, n15301, n15303, n15304, n15305, 
      n15307, n15308, n15310, n15311, n15312, n15313, n15314, n15315, n15316, 
      n15317, n15319, n15320, n15321, n15323, n15324, n15325, n15327, n15328, 
      n15329, n15330, n15331, n15332, n15333, n15334, n15336, n15337, n15338, 
      n15339, n15340, n15341, n15343, n15344, n15345, n15346, n15347, n15348, 
      n15349, n15350, n15352, n15353, n15354, n15355, n15356, n15357, n15358, 
      n15359, n15360, n15361, n15364, n15365, n15368, n15369, n15370, n15371, 
      n15372, n15373, n15375, n15376, n15377, n15378, n15380, n15381, n15382, 
      n15384, n15385, n15386, n15388, n15389, n15391, n15393, n15394, n15395, 
      n15398, n15400, n15401, n15404, n15405, n15406, n15410, n15411, n15412, 
      n15413, n15414, n15419, n15420, n15421, n15422, n15423, n15424, n15426, 
      n15427, n15429, n15430, n15432, n15433, n15434, n15435, n15436, n15437, 
      n15439, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, 
      n15449, n15450, n15451, n15452, n15453, n15455, n15456, n15457, n15458, 
      n15459, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, 
      n15471, n15473, n15476, n15477, n15480, n15481, n15482, n15483, n15485, 
      n15487, n15488, n15490, n15491, n15492, n15493, n15495, n15496, n15497, 
      n15499, n15500, n15502, n15503, n15507, n15508, n15509, n15512, n15513, 
      n15514, n15515, n15516, n15517, n15518, n15519, n15521, n15522, n15523, 
      n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, 
      n15534, n15535, n15540, n15541, n15542, n15543, n15545, n15546, n15547, 
      n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15558, 
      n15559, n15560, n15562, n15564, n15565, n15566, n15568, n15569, n15570, 
      n15571, n15572, n15573, n15575, n15577, n15579, n15580, n15581, n15583, 
      n15584, n15585, n15586, n15588, n15589, n15591, n15592, n15594, n15595, 
      n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, 
      n15607, n15608, n15609, n15610, n15613, n15614, n15615, n15616, n15617, 
      n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, 
      n15627, n15629, n15630, n15631, n15633, n15634, n15635, n15638, n15641, 
      n15642, n15643, n15644, n15647, n15648, n15649, n15650, n15651, n15652, 
      n15653, n15654, n15656, n15660, n15663, n15664, n15667, n15668, n15669, 
      n15670, n15671, n15672, n15673, n15674, n15676, n15677, n15678, n15679, 
      n15681, n15682, n15684, n15685, n15686, n15688, n15689, n15691, n15692, 
      n15693, n15694, n15695, n15696, n15697, n15700, n15701, n15702, n15703, 
      n15704, n15706, n15707, n15708, n15709, n15710, n15712, n15713, n15715, 
      n15716, n15717, n15718, n15719, n15721, n15722, n15723, n15726, n15727, 
      n15728, n15729, n15730, n15733, n15735, n15736, n15737, n15738, n15739, 
      n15740, n15741, n15742, n15743, n15745, n15748, n15750, n15751, n15752, 
      n15753, n15754, n15755, n15757, n15758, n15761, n15762, n15763, n15765, 
      n15767, n15768, n15770, n15771, n15772, n15773, n15774, n15775, n15776, 
      n15777, n15779, n15780, n15782, n15785, n15787, n15788, n15789, n15790, 
      n15791, n15792, n15794, n15795, n15796, n15797, n15798, n15799, n15800, 
      n15801, n15802, n15803, n15804, n15805, n15806, n15808, n15809, n15810, 
      n15811, n15812, n15814, n15816, n15817, n15818, n15819, n15821, n15822, 
      n15823, n15824, n15825, n15826, n15828, n15829, n15831, n15832, n15834, 
      n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15844, 
      n15846, n15848, n15849, n15850, n15852, n15853, n15854, n15855, n15857, 
      n15858, n15859, n15860, n15861, n15862, n15864, n15865, n15867, n15868, 
      n15869, n15870, n15871, n15872, n15873, n15876, n15877, n15878, n15879, 
      n15880, n15881, n15882, n15883, n15884, n15885, n15888, n15890, n15891, 
      n15892, n15893, n15894, n15896, n15897, n15898, n15899, n15903, n15904, 
      n15907, n15909, n15910, n15911, n15912, n15913, n15915, n15916, n15917, 
      n15918, n15919, n15922, n15924, n15925, n15926, n15928, n15929, n15930, 
      n15932, n15933, n15935, n15936, n15937, n15938, n15940, n15941, n15943, 
      n15945, n15946, n15947, n15949, n15951, n15952, n15953, n15955, n15956, 
      n15957, n15958, n15959, n15960, n15963, n15964, n15966, n15967, n15968, 
      n15969, n15971, n15972, n15973, n15974, n15975, n15978, n15979, n15980, 
      n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, 
      n15991, n15992, n15993, n15994, n15995, n15996, n15998, n15999, n16000, 
      n16004, n16006, n16007, n16009, n16010, n16013, n16014, n16015, n16016, 
      n16017, n16019, n16021, n16022, n16024, n16026, n16027, n16028, n16029, 
      n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16038, n16039, 
      n16040, n16041, n16042, n16043, n16045, n16046, n16047, n16048, n16049, 
      n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, 
      n16059, n16060, n16061, n16062, n16063, n16065, n16066, n16067, n16068, 
      n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, 
      n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, 
      n16091, n16093, n16094, n16095, n16096, n16097, n16098, n16101, n16102, 
      n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16113, 
      n16114, n16115, n16116, n16117, n16118, n16121, n16123, n16124, n16126, 
      n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, 
      n16137, n16138, n16140, n16141, n16144, n16146, n16147, n16149, n16150, 
      n16151, n16153, n16154, n16158, n16159, n16160, n16161, n16162, n16163, 
      n16165, n16167, n16168, n16169, n16170, n16171, n16173, n16174, n16175, 
      n16177, n16179, n16180, n16181, n16182, n16183, n16184, n16186, n16187, 
      n16190, n16191, n16192, n16193, n16195, n16196, n16197, n16198, n16199, 
      n16200, n16201, n16202, n16203, n16206, n16208, n16209, n16210, n16211, 
      n16213, n16216, n16217, n16218, n16220, n16221, n16222, n16224, n16225, 
      n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, 
      n16235, n16236, n16237, n16238, n16239, n16240, n16243, n16244, n16245, 
      n16246, n16247, n16248, n16249, n16250, n16252, n16254, n16255, n16256, 
      n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, 
      n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16275, n16277, 
      n16278, n16281, n16282, n16283, n16284, n16287, n16288, n16289, n16290, 
      n16291, n16292, n16293, n16294, n16295, n16296, n16298, n16299, n16301, 
      n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, 
      n16311, n16312, n16313, n16315, n16316, n16317, n16318, n16320, n16321, 
      n16324, n16325, n16327, n16328, n16332, n16333, n16334, n16336, n16337, 
      n16338, n16339, n16342, n16343, n16344, n16345, n16346, n16347, n16348, 
      n16350, n16351, n16353, n16355, n16356, n16357, n16358, n16359, n16360, 
      n16362, n16363, n16364, n16366, n16367, n16368, n16369, n16370, n16371, 
      n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, 
      n16381, n16382, n16385, n16388, n16389, n16390, n16391, n16392, n16393, 
      n16394, n16395, n16397, n16398, n16400, n16401, n16402, n16403, n16406, 
      n16407, n16410, n16411, n16412, n16416, n16417, n16419, n16420, n16421, 
      n16422, n16423, n16424, n16425, n16427, n16428, n16430, n16431, n16432, 
      n16435, n16439, n16440, n16443, n16444, n16445, n16446, n16447, n16448, 
      n16449, n16450, n16452, n16453, n16454, n16455, n16456, n16458, n16459, 
      n16460, n16461, n16463, n16466, n16467, n16468, n16469, n16470, n16471, 
      n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, 
      n16482, n16484, n16487, n16488, n16489, n16490, n16492, n16494, n16495, 
      n16496, n16497, n16498, n16499, n16500, n16502, n16503, n16505, n16508, 
      n16510, n16511, n16513, n16514, n16516, n16517, n16520, n16522, n16523, 
      n16524, n16525, n16526, n16528, n16529, n16530, n16531, n16532, n16533, 
      n16534, n16535, n16536, n16537, n16539, n16540, n16541, n16542, n16543, 
      n16544, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, 
      n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, 
      n16565, n16566, n16567, n16569, n16570, n16573, n16575, n16576, n16577, 
      n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16587, 
      n16589, n16590, n16591, n16593, n16595, n16596, n16597, n16598, n16599, 
      n16601, n16604, n16605, n16606, n16607, n16610, n16612, n16613, n16615, 
      n16617, n16618, n16619, n16621, n16623, n16624, n16625, n16627, n16628, 
      n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16638, 
      n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16647, n16648, 
      n16650, n16651, n16653, n16654, n16655, n16656, n16657, n16658, n16659, 
      n16660, n16663, n16665, n16666, n16667, n16668, n16669, n16670, n16671, 
      n16672, n16673, n16674, n16676, n16677, n16678, n16679, n16682, n16683, 
      n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, 
      n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16704, n16705, 
      n16706, n16707, n16708, n16709, n16712, n16713, n16715, n16716, n16720, 
      n16721, n16722, n16723, n16726, n16728, n16729, n16731, n16732, n16733, 
      n16735, n16736, n16737, n16739, n16740, n16741, n16742, n16743, n16744, 
      n16745, n16746, n16747, n16749, n16750, n16751, n16753, n16755, n16757, 
      n16758, n16759, n16760, n16762, n16763, n16765, n16766, n16767, n16771, 
      n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16781, 
      n16782, n16783, n16785, n16786, n16787, n16790, n16791, n16792, n16793, 
      n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, 
      n16803, n16804, n16805, n16806, n16809, n16810, n16813, n16814, n16815, 
      n16816, n16819, n16820, n16825, n16828, n16829, n16830, n16832, n16833, 
      n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, 
      n16843, n16845, n16847, n16848, n16849, n16851, n16853, n16854, n16855, 
      n16856, n16857, n16858, n16859, n16860, n16861, n16863, n16864, n16867, 
      n16868, n16869, n16871, n16873, n16874, n16876, n16877, n16878, n16879, 
      n16880, n16881, n16882, n16883, n16884, n16886, n16887, n16888, n16889, 
      n16890, n16892, n16893, n16896, n16897, n16898, n16900, n16901, n16902, 
      n16903, n16904, n16905, n16907, n16908, n16911, n16912, n16917, n16918, 
      n16919, n16920, n16921, n16922, n16924, n16929, n16930, n16931, n16932, 
      n16933, n16934, n16935, n16936, n16939, n16941, n16942, n16945, n16946, 
      n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, 
      n16957, n16960, n16961, n16962, n16963, n16964, n16966, n16967, n16968, 
      n16970, n16971, n16972, n16975, n16976, n16977, n16982, n16985, n16987, 
      n16988, n16989, n16990, n16992, n16993, n16994, n16996, n16997, n16998, 
      n16999, n17000, n17001, n17002, n17003, n17006, n17007, n17008, n17009, 
      n17013, n17017, n17018, n17020, n17021, n17022, n17023, n17024, n17025, 
      n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, 
      n17037, n17038, n17039, n17040, n17041, n17043, n17045, n17047, n17048, 
      n17051, n17055, n17057, n17058, n17060, n17062, n17063, n17064, n17066, 
      n17067, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17080, 
      n17081, n17083, n17084, n17085, n17086, n17087, n17089, n17090, n17091, 
      n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, 
      n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17110, n17112, 
      n17113, n17114, n17115, n17117, n17118, n17119, n17120, n17121, n17122, 
      n17124, n17125, n17126, n17127, n17128, n17129, n17131, n17132, n17134, 
      n17136, n17137, n17138, n17139, n17140, n17142, n17143, n17144, n17145, 
      n17147, n17148, n17150, n17151, n17152, n17153, n17154, n17155, n17156, 
      n17158, n17159, n17160, n17161, n17163, n17166, n17167, n17168, n17169, 
      n17171, n17172, n17173, n17176, n17177, n17178, n17179, n17180, n17182, 
      n17183, n17184, n17187, n17188, n17189, n17190, n17191, n17192, n17193, 
      n17194, n17195, n17197, n17198, n17201, n17202, n17205, n17207, n17209, 
      n17210, n17211, n17212, n17213, n17214, n17217, n17219, n17220, n17221, 
      n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17231, n17232, 
      n17233, n17234, n17236, n17237, n17238, n17240, n17242, n17243, n17245, 
      n17246, n17248, n17249, n17250, n17252, n17253, n17254, n17255, n17256, 
      n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, 
      n17266, n17267, n17269, n17270, n17271, n17272, n17273, n17274, n17275, 
      n17276, n17277, n17278, n17279, n17281, n17282, n17283, n17284, n17285, 
      n17286, n17287, n17288, n17292, n17293, n17294, n17295, n17296, n17297, 
      n17298, n17299, n17301, n17302, n17303, n17304, n17305, n17307, n17308, 
      n17309, n17310, n17311, n17312, n17313, n17314, n17316, n17317, n17318, 
      n17319, n17320, n17321, n17322, n17323, n17325, n17326, n17328, n17329, 
      n17331, n17332, n17333, n17334, n17335, n17338, n17339, n17340, n17341, 
      n17342, n17343, n17344, n17346, n17347, n17348, n17349, n17350, n17351, 
      n17353, n17354, n17356, n17357, n17358, n17359, n17360, n17361, n17363, 
      n17364, n17365, n17366, n17368, n17369, n17371, n17372, n17373, n17374, 
      n17377, n17378, n17381, n17382, n17383, n17388, n17390, n17391, n17392, 
      n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17402, 
      n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, 
      n17412, n17413, n17415, n17416, n17417, n17418, n17420, n17422, n17423, 
      n17424, n17425, n17426, n17428, n17429, n17430, n17433, n17435, n17436, 
      n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17447, n17448, 
      n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, 
      n17458, n17459, n17461, n17462, n17463, n17464, n17465, n17466, n17467, 
      n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, 
      n17478, n17480, n17482, n17483, n17484, n17485, n17486, n17487, n17489, 
      n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, 
      n17499, n17500, n17501, n17502, n17508, n17509, n17511, n17513, n17514, 
      n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, 
      n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, 
      n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, 
      n17542, n17544, n17546, n17551, n17552, n17553, n17554, n17555, n17556, 
      n17557, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17573, 
      n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17583, 
      n17584, n17586, n17591, n17592, n17593, n17594, n17595, n17596, n17597, 
      n17598, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, 
      n17612, n17613, n17615, n17616, n17617, n17618, n17621, n17623, n17624, 
      n17627, n17628, n17630, n17632, n17633, n17634, n17635, n17636, n17637, 
      n17638, n17639, n17642, n17643, n17644, n17645, n17646, n17647, n17648, 
      n17650, n17651, n17653, n17655, n17657, n17658, n17659, n17660, n17661, 
      n17662, n17663, n17664, n17665, n17668, n17669, n17673, n17674, n17677, 
      n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, 
      n17687, n17688, n17691, n17692, n17693, n17696, n17697, n17698, n17699, 
      n17700, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, 
      n17711, n17712, n17714, n17715, n17716, n17717, n17718, n17719, n17720, 
      n17721, n17723, n17724, n17725, n17726, n17727, n17730, n17731, n17732, 
      n17735, n17737, n17738, n17739, n17740, n17742, n17744, n17745, n17747, 
      n17748, n17750, n17751, n17753, n17754, n17755, n17756, n17757, n17758, 
      n17759, n17760, n17763, n17764, n17765, n17767, n17768, n17770, n17771, 
      n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17781, n17782, 
      n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, 
      n17793, n17794, n17795, n17797, n17798, n17799, n17800, n17801, n17803, 
      n17804, n17806, n17810, n17811, n17812, n17813, n17815, n17816, n17817, 
      n17818, n17819, n17820, n17821, n17823, n17824, n17826, n17829, n17830, 
      n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, 
      n17841, n17842, n17844, n17847, n17848, n17849, n17850, n17852, n17853, 
      n17854, n17855, n17856, n17857, n17858, n17859, n17861, n17862, n17863, 
      n17864, n17865, n17866, n17867, n17868, n17869, n17871, n17872, n17874, 
      n17875, n17876, n17877, n17878, n17879, n17880, n17882, n17884, n17885, 
      n17886, n17887, n17888, n17890, n17891, n17893, n17894, n17896, n17897, 
      n17898, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, 
      n17908, n17909, n17910, n17911, n17912, n17915, n17916, n17917, n17918, 
      n17920, n17921, n17922, n17923, n17925, n17926, n17927, n17928, n17929, 
      n17930, n17931, n17934, n17935, n17936, n17937, n17938, n17939, n17940, 
      n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17951, n17952, 
      n17954, n17955, n17957, n17958, n17959, n17960, n17961, n17962, n17963, 
      n17964, n17965, n17966, n17967, n17968, n17970, n17971, n17972, n17973, 
      n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17982, n17983, 
      n17984, n17985, n17986, n17987, n17988, n17989, n17991, n17992, n17993, 
      n17994, n17995, n17996, n17997, n17998, n17999, n18001, n18002, n18003, 
      n18004, n18005, n18006, n18007, n18012, n18013, n18014, n18015, n18017, 
      n18018, n18019, n18020, n18023, n18024, n18025, n18026, n18027, n18028, 
      n18029, n18031, n18032, n18034, n18035, n18036, n18037, n18038, n18039, 
      n18041, n18042, n18043, n18044, n18047, n18048, n18049, n18050, n18051, 
      n18054, n18055, n18056, n18058, n18059, n18060, n18061, n18062, n18063, 
      n18064, n18065, n18066, n18070, n18071, n18072, n18073, n18074, n18075, 
      n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, 
      n18086, n18087, n18088, n18089, n18090, n18094, n18095, n18096, n18098, 
      n18101, n18103, n18104, n18106, n18107, n18108, n18109, n18110, n18112, 
      n18113, n18114, n18115, n18116, n18120, n18121, n18122, n18123, n18124, 
      n18125, n18127, n18129, n18131, n18133, n18134, n18135, n18137, n18140, 
      n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, 
      n18150, n18152, n18153, n18155, n18156, n18157, n18159, n18160, n18162, 
      n18163, n18164, n18166, n18168, n18170, n18171, n18172, n18174, n18175, 
      n18176, n18178, n18179, n18180, n18182, n18183, n18184, n18186, n18187, 
      n18188, n18189, n18190, n18191, n18192, n18193, n18195, n18196, n18197, 
      n18198, n18199, n18200, n18201, n18202, n18204, n18205, n18207, n18208, 
      n18209, n18210, n18211, n18213, n18214, n18215, n18216, n18217, n18218, 
      n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, 
      n18228, n18229, n18231, n18232, n18233, n18234, n18235, n18236, n18237, 
      n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18246, n18249, 
      n18250, n18251, n18253, n18255, n18256, n18257, n18259, n18261, n18263, 
      n18264, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, 
      n18274, n18276, n18277, n18278, n18279, n18281, n18282, n18283, n18284, 
      n18288, n18289, n18290, n18291, n18293, n18294, n18295, n18296, n18298, 
      n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18308, n18309, 
      n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18319, 
      n18320, n18322, n18324, n18325, n18326, n18327, n18328, n18329, n18330, 
      n18331, n18335, n18338, n18339, n18340, n18341, n18342, n18345, n18346, 
      n18347, n18348, n18349, n18350, n18352, n18353, n18354, n18357, n18359, 
      n18360, n18362, n18363, n18364, n18365, n18366, n18367, n18369, n18370, 
      n18371, n18372, n18374, n18375, n18376, n18377, n18378, n18379, n18380, 
      n18381, n18382, n18383, n18384, n18386, n18388, n18389, n18390, n18391, 
      n18392, n18393, n18394, n18395, n18398, n18399, n18401, n18402, n18403, 
      n18404, n18405, n18406, n18407, n18408, n18410, n18412, n18413, n18415, 
      n18416, n18417, n18420, n18421, n18422, n18423, n18424, n18425, n18426, 
      n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18436, 
      n18438, n18439, n18440, n18445, n18446, n18447, n18449, n18450, n18451, 
      n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, 
      n18461, n18462, n18463, n18464, n18466, n18467, n18468, n18469, n18470, 
      n18471, n18472, n18473, n18474, n18475, n18477, n18478, n18479, n18480, 
      n18481, n18482, n18483, n18484, n18485, n18487, n18488, n18489, n18490, 
      n18491, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, 
      n18501, n18502, n18504, n18505, n18506, n18507, n18508, n18509, n18510, 
      n18511, n18512, n18515, n18516, n18518, n18519, n18520, n18522, n18523, 
      n18524, n18525, n18526, n18527, n18529, n18530, n18532, n18534, n18536, 
      n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, 
      n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18554, n18556, 
      n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, 
      n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, 
      n18575, n18576, n18577, n18578, n18579, n18580, n18582, n18584, n18585, 
      n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, 
      n18595, n18597, n18599, n18600, n18601, n18602, n18603, n18604, n18605, 
      n18606, n18608, n18609, n18610, n18611, n18612, n18615, n18616, n18617, 
      n18618, n18619, n18620, n18622, n18623, n18624, n18625, n18626, n18628, 
      n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18640, 
      n18641, n18642, n18643, n18645, n18647, n18650, n18651, n18652, n18653, 
      n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, 
      n18663, n18665, n18667, n18668, n18669, n18670, n18671, n18673, n18674, 
      n18675, n18679, n18680, n18681, n18682, n18683, n18685, n18686, n18687, 
      n18688, n18689, n18690, n18691, n18692, n18694, n18696, n18697, n18698, 
      n18699, n18700, n18701, n18702, n18704, n18705, n18706, n18707, n18708, 
      n18709, n18710, n18711, n18712, n18715, n18716, n18717, n18718, n18719, 
      n18720, n18721, n18722, n18723, n18725, n18726, n18728, n18729, n18730, 
      n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18741, 
      n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, 
      n18751, n18752, n18755, n18757, n18758, n18759, n18762, n18763, n18764, 
      n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18773, n18774, 
      n18776, n18777, n18778, n18780, n18782, n18783, n18784, n18785, n18786, 
      n18787, n18788, n18790, n18792, n18793, n18794, n18795, n18796, n18797, 
      n18800, n18801, n18803, n18804, n18806, n18807, n18808, n18809, n18810, 
      n18811, n18813, n18814, n18815, n18816, n18817, n18819, n18822, n18825, 
      n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18836, 
      n18837, n18838, n18841, n18842, n18843, n18844, n18845, n18846, n18847, 
      n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, 
      n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, 
      n18867, n18869, n18870, n18871, n18872, n18873, n18875, n18876, n18877, 
      n18879, n18880, n18883, n18884, n18886, n18887, n18888, n18889, n18890, 
      n18891, n18893, n18894, n18896, n18897, n18898, n18900, n18901, n18902, 
      n18903, n18904, n18905, n18907, n18908, n18909, n18910, n18911, n18912, 
      n18913, n18914, n18915, n18917, n18918, n18920, n18921, n18922, n18923, 
      n18924, n18926, n18927, n18928, n18929, n18930, n18931, n18933, n18934, 
      n18935, n18936, n18937, n18938, n18939, n18941, n18942, n18943, n18944, 
      n18945, n18946, n18947, n18948, n18950, n18951, n18952, n18953, n18954, 
      n18956, n18958, n18959, n18960, n18961, n18962, n18966, n18967, n18968, 
      n18969, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18979, 
      n18980, n18981, n18983, n18984, n18985, n18986, n18987, n18988, n18989, 
      n18990, n18991, n18992, n18993, n18994, n18996, n18997, n18998, n18999, 
      n19000, n19001, n19002, n19003, n19005, n19006, n19007, n19008, n19009, 
      n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, 
      n19020, n19021, n19022, n19024, n19025, n19026, n19027, n19028, n19030, 
      n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, 
      n19041, n19042, n19043, n19045, n19047, n19048, n19050, n19051, n19052, 
      n19053, n19054, n19055, n19059, n19060, n19061, n19062, n19064, n19065, 
      n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, 
      n19075, n19077, n19078, n19080, n19081, n19082, n19083, n19084, n19085, 
      n19088, n19089, n19090, n19091, n19093, n19094, n19095, n19096, n19097, 
      n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19108, 
      n19109, n19111, n19112, n19113, n19115, n19118, n19119, n19120, n19121, 
      n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, 
      n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, 
      n19142, n19143, n19145, n19146, n19147, n19151, n19152, n19153, n19154, 
      n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, 
      n19164, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19175, 
      n19177, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, 
      n19187, n19188, n19191, n19193, n19194, n19195, n19196, n19197, n19198, 
      n19200, n19201, n19202, n19203, n19204, n19206, n19207, n19209, n19210, 
      n19211, n19213, n19214, n19215, n19216, n19217, n19218, n19220, n19221, 
      n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19231, 
      n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19240, n19241, 
      n19242, n19244, n19246, n19249, n19250, n19252, n19253, n19254, n19255, 
      n19257, n19258, n19259, n19260, n19261, n19262, n19264, n19266, n19268, 
      n19270, n19271, n19272, n19274, n19276, n19277, n19278, n19279, n19280, 
      n19281, n19283, n19284, n19285, n19287, n19288, n19289, n19290, n19292, 
      n19293, n19294, n19295, n19296, n19297, n19298, n19300, n19302, n19303, 
      n19304, n19305, n19307, n19308, n19309, n19310, n19311, n19312, n19313, 
      n19316, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, 
      n19326, n19327, n19328, n19329, n19331, n19332, n19334, n19335, n19336, 
      n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19347, 
      n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, 
      n19358, n19359, n19360, n19361, n19362, n19364, n19366, n19367, n19368, 
      n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, 
      n19379, n19380, n19381, n19382, n19384, n19385, n19387, n19388, n19389, 
      n19391, n19392, n19393, n19395, n19396, n19397, n19398, n19400, n19401, 
      n19402, n19403, n19404, n19405, n19407, n19408, n19409, n19410, n19411, 
      n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19420, n19421, 
      n19422, n19423, n19424, n19425, n19426, n19428, n19430, n19431, n19432, 
      n19433, n19434, n19435, n19436, n19438, n19439, n19440, n19442, n19443, 
      n19444, n19445, n19446, n19448, n19449, n19450, n19452, n19453, n19454, 
      n19455, n19456, n19458, n19459, n19460, n19463, n19464, n19465, n19466, 
      n19467, n19469, n19470, n19471, n19472, n19473, n19475, n19476, n19477, 
      n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19486, n19488, 
      n19490, n19492, n19493, n19495, n19496, n19497, n19498, n19499, n19501, 
      n19503, n19504, n19505, n19507, n19508, n19511, n19513, n19514, n19515, 
      n19516, n19517, n19518, n19521, n19524, n19525, n19527, n19528, n19529, 
      n19530, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, 
      n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19548, n19549, 
      n19550, n19551, n19552, n19553, n19554, n19557, n19559, n19560, n19561, 
      n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, 
      n19572, n19573, n19574, n19575, n19576, n19577, n19579, n19580, n19581, 
      n19582, n19583, n19584, n19586, n19587, n19588, n19589, n19590, n19591, 
      n19592, n19593, n19594, n19595, n19596, n19597, n19599, n19600, n19601, 
      n19604, n19605, n19606, n19608, n19609, n19610, n19612, n19613, n19614, 
      n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, 
      n19624, n19627, n19629, n19630, n19631, n19632, n19633, n19636, n19637, 
      n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, 
      n19648, n19649, n19650, n19652, n19653, n19654, n19655, n19656, n19657, 
      n19658, n19659, n19660, n19661, n19662, n19663, n19665, n19666, n19667, 
      n19668, n19669, n19670, n19671, n19673, n19674, n19675, n19676, n19677, 
      n19678, n19679, n19680, n19681, n19682, n19683, n19685, n19686, n19687, 
      n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19696, n19697, 
      n19698, n19699, n19700, n19701, n19702, n19704, n19706, n19707, n19708, 
      n19709, n19712, n19713, n19714, n19716, n19717, n19718, n19719, n19720, 
      n19721, n19722, n19724, n19725, n19726, n19727, n19728, n19729, n19730, 
      n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, 
      n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, 
      n19749, n19750, n19751, n19754, n19755, n19756, n19758, n19759, n19760, 
      n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, 
      n19770, n19771, n19772, n19773, n19774, n19775, n19777, n19778, n19780, 
      n19781, n19782, n19783, n19784, n19785, n19786, n19788, n19791, n19792, 
      n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, 
      n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, 
      n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, 
      n19821, n19822, n19823, n19824, n19825, n19827, n19828, n19829, n19830, 
      n19831, n19833, n19835, n19836, n19837, n19838, n19839, n19840, n19843, 
      n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, 
      n19855, n19856, n19857, n19859, n19860, n19862, n19863, n19864, n19865, 
      n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, 
      n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, 
      n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, 
      n19893, n19894, n19895, n19896, n19897, n19898, n19900, n19901, n19902, 
      n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, 
      n19913, n19914, n19915, n19918, n19919, n19920, n19921, n19922, n19923, 
      n19924, n19925, n19927, n19928, n19929, n19930, n19931, n19932, n19933, 
      n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, 
      n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, 
      n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19962, n19963, 
      n19964, n19965, n19966, n19967, n19968, n19969, n19971, n19972, n19973, 
      n19975, n19976, n19978, n19979, n19980, n19982, n19983, n19984, n19985, 
      n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, 
      n19995, n19996, n19997, n19998, n19999, n20000, n20002, n20003, n20004, 
      n20006, n20007, n20008, n20010, n20013, n20016, n20018, n20019, n20020, 
      n20021, n20022, n20024, n20025, n20026, n20027, n20028, n20029, n20030, 
      n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, 
      n20041, n20042, n20043, n20044, n20045, n20047, n20048, n20049, n20050, 
      n20051, n20052, n20053, n20056, n20057, n20058, n20059, n20061, n20062, 
      n20063, n20064, n20065, n20066, n20068, n20069, n20070, n20074, n20076, 
      n20077, n20078, n20080, n20082, n20083, n20084, n20085, n20087, n20088, 
      n20089, n20090, n20092, n20093, n20094, n20095, n20096, n20097, n20098, 
      n20099, n20100, n20101, n20102, n20103, n20105, n20107, n20108, n20109, 
      n20111, n20112, n20113, n20116, n20117, n20118, n20119, n20120, n20121, 
      n20122, n20123, n20125, n20126, n20128, n20129, n20131, n20132, n20133, 
      n20134, n20135, n20136, n20137, n20139, n20140, n20143, n20145, n20146, 
      n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, 
      n20156, n20157, n20158, n20159, n20160, n20164, n20166, n20167, n20168, 
      n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, 
      n20180, n20184, n20185, n20186, n20187, n20188, n20190, n20191, n20194, 
      n20196, n20197, n20198, n20199, n20200, n20201, n20203, n20205, n20206, 
      n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20216, 
      n20217, n20219, n20221, n20222, n20223, n20225, n20226, n20227, n20229, 
      n20230, n20232, n20234, n20235, n20236, n20237, n20238, n20239, n20241, 
      n20242, n20243, n20244, n20245, n20250, n20251, n20254, n20255, n20256, 
      n20257, n20260, n20261, n20262, n20263, n20264, n20266, n20267, n20268, 
      n20270, n20274, n20276, n20277, n20278, n20279, n20280, n20282, n20284, 
      n20286, n20287, n20288, n20289, n20290, n20294, n20295, n20296, n20297, 
      n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, 
      n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20316, 
      n20317, n20319, n20321, n20322, n20323, n20324, n20325, n20326, n20328, 
      n20329, n20330, n20331, n20332, n20333, n20335, n20336, n20337, n20339, 
      n20340, n20341, n20342, n20343, n20344, n20346, n20347, n20348, n20350, 
      n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, 
      n20361, n20362, n20363, n20364, n20365, n20367, n20368, n20369, n20370, 
      n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20381, 
      n20384, n20386, n20387, n20388, n20389, n20391, n20392, n20394, n20395, 
      n20396, n20397, n20398, n20399, n20400, n20402, n20403, n20404, n20405, 
      n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20414, n20416, 
      n20418, n20419, n20420, n20421, n20423, n20424, n20425, n20426, n20427, 
      n20429, n20430, n20431, n20433, n20434, n20435, n20436, n20437, n20438, 
      n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, 
      n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, 
      n20457, n20458, n20460, n20462, n20463, n20464, n20465, n20468, n20469, 
      n20470, n20472, n20473, n20474, n20476, n20479, n20480, n20481, n20482, 
      n20483, n20484, n20485, n20486, n20487, n20489, n20490, n20491, n20492, 
      n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, 
      n20502, n20503, n20504, n20505, n20507, n20508, n20509, n20510, n20511, 
      n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20522, 
      n20524, n20525, n20526, n20528, n20530, n20531, n20533, n20535, n20536, 
      n20537, n20538, n20539, n20540, n20541, n20544, n20545, n20546, n20547, 
      n20549, n20550, n20551, n20554, n20555, n20559, n20560, n20561, n20562, 
      n20564, n20565, n20566, n20570, n20571, n20572, n20573, n20574, n20575, 
      n20576, n20577, n20578, n20579, n20580, n20581, n20583, n20584, n20585, 
      n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, 
      n20595, n20596, n20597, n20600, n20601, n20602, n20604, n20605, n20607, 
      n20608, n20609, n20611, n20612, n20613, n20614, n20615, n20616, n20618, 
      n20619, n20620, n20621, n20622, n20623, n20625, n20626, n20627, n20628, 
      n20629, n20632, n20634, n20635, n20636, n20637, n20638, n20639, n20641, 
      n20642, n20643, n20644, n20646, n20648, n20649, n20651, n20653, n20654, 
      n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, 
      n20665, n20666, n20668, n20669, n20670, n20671, n20672, n20673, n20674, 
      n20675, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, 
      n20685, n20686, n20687, n20689, n20690, n20691, n20692, n20693, n20694, 
      n20695, n20696, n20697, n20698, n20699, n20701, n20702, n20703, n20704, 
      n20706, n20707, n20708, n20709, n20713, n20715, n20716, n20717, n20718, 
      n20719, n20720, n20721, n20723, n20724, n20725, n20726, n20727, n20728, 
      n20730, n20731, n20732, n20734, n20735, n20736, n20737, n20738, n20739, 
      n20740, n20741, n20743, n20744, n20746, n20747, n20748, n20749, n20750, 
      n20751, n20752, n20753, n20754, n20756, n20758, n20759, n20761, n20762, 
      n20764, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, 
      n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20787, 
      n20788, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, 
      n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, 
      n20807, n20808, n20809, n20810, n20811, n20813, n20815, n20816, n20817, 
      n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20827, 
      n20828, n20829, n20830, n20831, n20832, n20833, n20835, n20836, n20838, 
      n20839, n20840, n20841, n20843, n20844, n20845, n20846, n20849, n20850, 
      n20851, n20852, n20855, n20856, n20858, n20859, n20860, n20862, n20863, 
      n20864, n20865, n20866, n20867, n20869, n20870, n20871, n20872, n20873, 
      n20874, n20875, n20876, n20877, n20878, n20879, n20881, n20882, n20883, 
      n20884, n20885, n20886, n20887, n20888, n20889, n20891, n20892, n20893, 
      n20894, n20895, n20896, n20897, n20898, n20901, n20903, n20907, n20910, 
      n20911, n20912, n20914, n20915, n20919, n20920, n20921, n20922, n20923, 
      n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20936, 
      n20939, n20941, n20943, n20944, n20945, n20946, n20947, n20948, n20949, 
      n20951, n20952, n20954, n20955, n20956, n20957, n20958, n20959, n20960, 
      n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, 
      n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, 
      n20980, n20981, n20982, n20984, n20986, n20987, n20988, n20989, n20991, 
      n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, 
      n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, 
      n21010, n21011, n21012, n21013, n21014, n21017, n21018, n21019, n21020, 
      n21021, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, 
      n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, 
      n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, 
      n21049, n21050, n21051, n21052, n21053, n21055, n21056, n21057, n21058, 
      n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, 
      n21068, n21069, n21071, n21072, n21073, n21074, n21076, n21077, n21079, 
      n21080, n21081, n21084, n21085, n21086, n21087, n21090, n21091, n21093, 
      n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21103, 
      n21104, n21105, n21108, n21109, n21110, n21111, n21114, n21116, n21117, 
      n21118, n21119, n21120, n21121, n21124, n21125, n21126, n21127, n21128, 
      n21130, n21132, n21133, n21134, n21135, n21136, n21137, n21139, n21140, 
      n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, 
      n21150, n21152, n21154, n21156, n21157, n21158, n21159, n21160, n21161, 
      n21162, n21163, n21164, n21166, n21167, n21168, n21169, n21170, n21171, 
      n21172, n21174, n21176, n21177, n21181, n21182, n21184, n21186, n21187, 
      n21188, n21190, n21191, n21192, n21195, n21196, n21197, n21198, n21201, 
      n21202, n21204, n21206, n21207, n21208, n21211, n21212, n21213, n21214, 
      n21215, n21216, n21217, n21218, n21219, n21220, n21223, n21224, n21225, 
      n21226, n21227, n21229, n21231, n21232, n21233, n21234, n21235, n21236, 
      n21238, n21239, n21241, n21242, n21245, n21246, n21247, n21248, n21249, 
      n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21259, 
      n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, 
      n21269, n21270, n21271, n21272, n21274, n21277, n21278, n21279, n21280, 
      n21282, n21283, n21284, n21285, n21287, n21288, n21289, n21290, n21291, 
      n21292, n21293, n21294, n21296, n21297, n21298, n21299, n21300, n21301, 
      n21302, n21305, n21306, n21307, n21308, n21309, n21310, n21316, n21317, 
      n21318, n21319, n21322, n21323, n21324, n21326, n21327, n21328, n21329, 
      n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, 
      n21339, n21340, n21341, n21342, n21343, n21345, n21346, n21347, n21349, 
      n21350, n21351, n21352, n21354, n21356, n21357, n21358, n21359, n21360, 
      n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, 
      n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, 
      n21379, n21380, n21381, n21382, n21383, n21384, n21386, n21387, n21388, 
      n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21397, n21398, 
      n21399, n21401, n21402, n21403, n21405, n21406, n21407, n21408, n21409, 
      n21410, n21412, n21413, n21414, n21415, n21416, n21417, n21419, n21420, 
      n21421, n21422, n21423, n21424, n21426, n21428, n21429, n21431, n21432, 
      n21433, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, 
      n21443, n21445, n21446, n21448, n21449, n21450, n21451, n21452, n21453, 
      n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, 
      n21463, n21464, n21465, n21467, n21468, n21469, n21472, n21475, n21476, 
      n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, 
      n21486, n21488, n21489, n21491, n21492, n21493, n21494, n21496, n21497, 
      n21498, n21499, n21501, n21503, n21504, n21505, n21506, n21507, n21508, 
      n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, 
      n21518, n21519, n21520, n21521, n21522, n21524, n21527, n21528, n21529, 
      n21531, n21532, n21533, n21534, n21535, n21536, n21539, n21540, n21541, 
      n21542, n21543, n21545, n21546, n21547, n21548, n21549, n21550, n21551, 
      n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, 
      n21561, n21562, n21564, n21565, n21566, n21567, n21568, n21569, n21570, 
      n21571, n21573, n21574, n21575, n21576, n21577, n21579, n21580, n21581, 
      n21582, n21583, n21584, n21586, n21587, n21588, n21589, n21590, n21591, 
      n21592, n21593, n21594, n21596, n21597, n21598, n21599, n21601, n21602, 
      n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21612, n21614, 
      n21616, n21617, n21618, n21620, n21621, n21622, n21623, n21624, n21625, 
      n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, 
      n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21644, 
      n21645, n21646, n21647, n21648, n21649, n21652, n21653, n21654, n21655, 
      n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, 
      n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, 
      n21674, n21675, n21676, n21678, n21679, n21681, n21682, n21683, n21684, 
      n21685, n21686, n21687, n21688, n21690, n21691, n21692, n21693, n21694, 
      n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, 
      n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, 
      n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, 
      n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21730, n21731, 
      n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, 
      n21741, n21742, n21743, n21745, n21747, n21748, n21749, n21750, n21751, 
      n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, 
      n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21770, 
      n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, 
      n21780, n21782, n21783, n21784, n21786, n21787, n21788, n21789, n21790, 
      n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21799, n21800, 
      n21801, n21802, n21803, n21804, n21805, n21806, n21808, n21809, n21810, 
      n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21820, n21821, 
      n21822, n21823, n21825, n21826, n21827, n21828, n21829, n21830, n21831, 
      n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, 
      n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, 
      n21850, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, 
      n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, 
      n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, 
      n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, 
      n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, 
      n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, 
      n21905, n21906, n21908, n21909, n21910, n21911, n21912, n21913, n21914, 
      n21915, n21916, n21917, n21919, n21920, n21921, n21923, n21924, n21925, 
      n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, 
      n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, 
      n21944, n21945, n21946, n21947, n21949, n21950, n21951, n21952, n21953, 
      n21954, n21956, n21957, n21958, n21959, n21960, n21961, n21963, n21964, 
      n21965, n21966, n21967, n21968, n21969, n21971, n21972, n21973, n21974, 
      n21975, n21976, n21977, n21978, n21979, n21980, n21982, n21983, n21984, 
      n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, 
      n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, 
      n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22012, 
      n22013, n22014, n22015, n22017, n22018, n22019, n22020, n22021, n22022, 
      n22023, n22024, n22025, n22026, n22027, n22029, n22030, n22032, n22034, 
      n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, 
      n22044, n22045, n22047, n22048, n22050, n22051, n22055, n22056, n22057, 
      n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, 
      n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22075, n22076, 
      n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, 
      n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, 
      n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, 
      n22104, n22105, n22106, n22107, n22108, n22110, n22111, n22113, n22114, 
      n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, 
      n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, 
      n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22143, 
      n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, 
      n22153, n22154, n22155, n22156, n22157, n22159, n22160, n22161, n22162, 
      n22163, n22165, n22166, n22167, n22168, n22170, n22171, n22172, n22173, 
      n22174, n22176, n22177, n22178, n22181, n22182, n22183, n22184, n22186, 
      n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, 
      n22196, n22197, n22198, n22199, n22200, n22201, n22203, n22204, n22205, 
      n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, 
      n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, 
      n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, 
      n22233, n22234, n22235, n22236, n22238, n22239, n22240, n22241, n22242, 
      n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22252, 
      n22253, n22254, n22255, n22256, n22258, n22259, n22261, n22262, n22263, 
      n22264, n22265, n22266, n22267, n22268, n22270, n22271, n22272, n22274, 
      n22275, n22277, n22278, n22279, n22280, n22281, n22282, n22284, n22285, 
      n22286, n22287, n22288, n22289, n22291, n22292, n22293, n22294, n22295, 
      n22296, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, 
      n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, 
      n22315, n22316, n22317, n22319, n22320, n22321, n22322, n22323, n22324, 
      n22325, n22326, n22327, n22328, n22329, n22330, n22332, n22333, n22334, 
      n22335, n22337, n22340, n22341, n22342, n22343, n22344, n22345, n22346, 
      n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22356, 
      n22358, n22359, n22360, n22361, n22362, n22364, n22365, n22366, n22367, 
      n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, 
      n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, 
      n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22396, 
      n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, 
      n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, 
      n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22424, n22425, 
      n22426, n22427, n22429, n22430, n22431, n22432, n22433, n22435, n22436, 
      n22438, n22439, n22441, n22442, n22443, n22444, n22445, n22446, n22447, 
      n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22456, n22457, 
      n22458, n22459, n22462, n22463, n22464, n22465, n22466, n22467, n22468, 
      n22469, n22470, n22473, n22474, n22475, n22476, n22478, n22479, n22482, 
      n22483, n22484, n22485, n22486, n22487, n22488, n22490, n22491, n22492, 
      n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, 
      n22503, n22505, n22506, n22508, n22509, n22510, n22511, n22512, n22513, 
      n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, 
      n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, 
      n22532, n22533, n22534, n22536, n22537, n22538, n22541, n22542, n22543, 
      n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, 
      n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562, 
      n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, 
      n22572, n22573, n22574, n22575, n22576, n22579, n22580, n22581, n22582, 
      n22583, n22584, n22586, n22587, n22588, n22590, n22592, n22594, n22595, 
      n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, 
      n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22613, n22614, 
      n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, 
      n22624, n22625, n22627, n22628, n22629, n22630, n22633, n22634, n22635, 
      n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, 
      n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, 
      n22654, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, 
      n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, 
      n22673, n22674, n22675, n22676, n22677, n22678, n22680, n22681, n22682, 
      n22683, n22684, n22686, n22687, n22688, n22689, n22690, n22693, n22694, 
      n22695, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, 
      n22705, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, 
      n22716, n22717, n22718, n22719, n22720, n22722, n22723, n22724, n22725, 
      n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, 
      n22735, n22736, n22737, n22740, n22741, n22742, n22743, n22744, n22745, 
      n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, 
      n22755, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, 
      n22765, n22766, n22767, n22768, n22769, n22771, n22772, n22773, n22774, 
      n22775, n22776, n22778, n22780, n22781, n22782, n22783, n22784, n22787, 
      n22789, n22790, n22791, n22792, n22793, n22795, n22796, n22797, n22798, 
      n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, 
      n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, 
      n22818, n22819, n22820, n22822, n22823, n22824, n22825, n22826, n22828, 
      n22829, n22830, n22831, n22833, n22834, n22836, n22837, n22838, n22839, 
      n22840, n22841, n22842, n22843, n22845, n22846, n22849, n22850, n22851, 
      n22852, n22853, n22854, n22856, n22857, n22858, n22859, n22860, n22861, 
      n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, 
      n22871, n22872, n22873, n22875, n22876, n22877, n22878, n22879, n22880, 
      n22881, n22882, n22884, n22885, n22886, n22887, n22889, n22890, n22891, 
      n22892, n22893, n22894, n22895, n22896, n22897, n22899, n22900, n22901, 
      n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, 
      n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, 
      n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, 
      n22929, n22931, n22932, n22934, n22935, n22937, n22939, n22940, n22942, 
      n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, 
      n22952, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22962, 
      n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, 
      n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22982, n22983, 
      n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, 
      n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23003, 
      n23004, n23005, n23006, n23007, n23009, n23010, n23011, n23012, n23013, 
      n23015, n23016, n23017, n23018, n23019, n23020, n23022, n23023, n23024, 
      n23025, n23026, n23027, n23028, n23030, n23031, n23032, n23033, n23034, 
      n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23044, 
      n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, 
      n23054, n23055, n23056, n23057, n23058, n23060, n23061, n23062, n23063, 
      n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, 
      n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, 
      n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, 
      n23091, n23093, n23094, n23095, n23096, n23098, n23099, n23100, n23101, 
      n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23110, n23111, 
      n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120, 
      n23121, n23122, n23123, n23124, n23125, n23127, n23128, n23129, n23131, 
      n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23140, n23141, 
      n23142, n23143, n23145, n23146, n23147, n23148, n23149, n23151, n23152, 
      n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, 
      n23163, n23164, n23165, n23166, n23167, n23169, n23171, n23172, n23173, 
      n23174, n23175, n23177, n23178, n23180, n23181, n23182, n23183, n23184, 
      n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, 
      n23194, n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23206, 
      n23207, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, 
      n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, 
      n23226, n23227, n23228, n23229, n23232, n23234, n23237, n23238, n23239, 
      n23240, n23241, n23242, n23243, n23244, n23245, n23247, n23248, n23249, 
      n23250, n23251, n23252, n23253, n23255, n23256, n23257, n23259, n23262, 
      n23263, n23264, n23265, n23266, n23267, n23270, n23271, n23272, n23274, 
      n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, 
      n23284, n23286, n23289, n23290, n23291, n23292, n23293, n23294, n23295, 
      n23296, n23297, n23298, n23299, n23301, n23302, n23303, n23305, n23306, 
      n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, 
      n23316, n23317, n23318, n23320, n23321, n23322, n23324, n23325, n23328, 
      n23329, n23330, n23331, n23333, n23334, n23335, n23337, n23338, n23340, 
      n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23349, n23350, 
      n23351, n23352, n23354, n23355, n23356, n23357, n23358, n23359, n23360, 
      n23361, n23362, n23363, n23364, n23365, n23367, n23368, n23369, n23370, 
      n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, 
      n23381, n23382, n23383, n23385, n23386, n23387, n23389, n23390, n23391, 
      n23392, n23393, n23394, n23396, n23397, n23399, n23400, n23401, n23403, 
      n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23412, n23413, 
      n23414, n23416, n23418, n23419, n23420, n23421, n23422, n23423, n23425, 
      n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, 
      n23435, n23439, n23440, n23441, n23442, n23444, n23447, n23450, n23452, 
      n23453, n23455, n23456, n23458, n23459, n23460, n23461, n23462, n23464, 
      n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473, 
      n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23482, n23483, 
      n23484, n23485, n23487, n23488, n23489, n23493, n23494, n23496, n23500, 
      n23502, n23504, n23505, n23506, n23508, n23509, n23510, n23511, n23512, 
      n23513, n23515, n23516, n23517, n23518, n23520, n23521, n23522, n23523, 
      n23525, n23526, n23528, n23529, n23530, n23531, n23532, n23533, n23534, 
      n23535, n23537, n23538, n23539, n23540, n23542, n23543, n23544, n23545, 
      n23546, n23547, n23548, n23549, n23550, n23552, n23553, n23554, n23555, 
      n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23565, 
      n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23574, n23575, 
      n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, 
      n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, 
      n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, 
      n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23613, 
      n23614, n23616, n23617, n23619, n23620, n23621, n23622, n23623, n23624, 
      n23625, n23627, n23630, n23631, n23632, n23633, n23634, n23635, n23636, 
      n23637, n23638, n23639, n23640, n23641, n23645, n23648, n23649, n23652, 
      n23653, n23654, n23655, n23656, n23658, n23659, n23660, n23661, n23662, 
      n23663, n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, 
      n23674, n23675, n23676, n23677, n23680, n23681, n23682, n23683, n23684, 
      n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, 
      n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23702, n23704, 
      n23705, n23707, n23709, n23710, n23711, n23712, n23713, n23714, n23715, 
      n23716, n23717, n23719, n23720, n23722, n23723, n23724, n23725, n23727, 
      n23728, n23729, n23730, n23732, n23733, n23734, n23736, n23737, n23738, 
      n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, 
      n23748, n23749, n23750, n23751, n23752, n23754, n23755, n23756, n23757, 
      n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, 
      n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, 
      n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, 
      n23785, n23786, n23787, n23788, n23789, n23790, n23792, n23793, n23794, 
      n23795, n23796, n23797, n23799, n23800, n23801, n23802, n23803, n23804, 
      n23805, n23806, n23807, n23808, n23809, n23812, n23813, n23814, n23816, 
      n23817, n23818, n23819, n23820, n23821, n23822, n23824, n23825, n23826, 
      n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, 
      n23836, n23838, n23839, n23841, n23842, n23843, n23844, n23845, n23846, 
      n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23855, n23857, 
      n23858, n23859, n23861, n23862, n23863, n23864, n23865, n23866, n23867, 
      n23868, n23869, n23870, n23871, n23873, n23874, n23876, n23878, n23879, 
      n23880, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, 
      n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, 
      n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, 
      n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23917, 
      n23918, n23919, n23920, n23921, n23922, n23924, n23925, n23926, n23927, 
      n23928, n23929, n23930, n23931, n23933, n23934, n23936, n23937, n23938, 
      n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, 
      n23948, n23949, n23950, n23952, n23953, n23954, n23955, n23957, n23958, 
      n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, 
      n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, 
      n23977, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23987, 
      n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, 
      n23997, n24000, n24001, n24002, n24005, n24006, n24007, n24009, n24011, 
      n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020, 
      n24022, n24023, n24024, n24025, n24026, n24028, n24029, n24030, n24031, 
      n24032, n24033, n24034, n24036, n24037, n24038, n24039, n24040, n24042, 
      n24043, n24045, n24047, n24048, n24049, n24050, n24051, n24052, n24053, 
      n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062, 
      n24063, n24064, n24065, n24067, n24068, n24069, n24070, n24071, n24072, 
      n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24081, n24082, 
      n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, 
      n24094, n24095, n24096, n24098, n24100, n24101, n24102, n24104, n24105, 
      n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, 
      n24116, n24117, n24118, n24119, n24120, n24121, n24123, n24125, n24126, 
      n24127, n24128, n24129, n24131, n24132, n24133, n24134, n24135, n24136, 
      n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24145, n24146, 
      n24147, n24148, n24149, n24150, n24152, n24153, n24154, n24155, n24156, 
      n24157, n24158, n24159, n24161, n24162, n24163, n24164, n24165, n24166, 
      n24167, n24168, n24169, n24170, n24172, n24173, n24174, n24175, n24176, 
      n24177, n24178, n24180, n24181, n24182, n24184, n24185, n24187, n24191, 
      n24192, n24193, n24194, n24195, n24196, n24198, n24199, n24202, n24203, 
      n24205, n24206, n24207, n24208, n24209, n24210, n24214, n24216, n24217, 
      n24218, n24219, n24221, n24222, n24223, n24224, n24225, n24226, n24227, 
      n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24238, 
      n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24250, 
      n24251, n24253, n24254, n24257, n24258, n24261, n24263, n24265, n24266, 
      n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275, 
      n24276, n24277, n24278, n24279, n24280, n24282, n24283, n24284, n24285, 
      n24287, n24290, n24292, n24293, n24294, n24295, n24296, n24297, n24298, 
      n24300, n24301, n24302, n24303, n24304, n24305, n24307, n24308, n24309, 
      n24310, n24311, n24312, n24313, n24314, n24316, n24317, n24318, n24323, 
      n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332, 
      n24333, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, 
      n24343, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24353, 
      n24355, n24357, n24359, n24360, n24363, n24364, n24365, n24366, n24369, 
      n24370, n24371, n24372, n24373, n24374, n24377, n24378, n24380, n24381, 
      n24382, n24383, n24386, n24387, n24388, n24389, n24390, n24391, n24392, 
      n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401, 
      n24402, n24403, n24404, n24406, n24407, n24408, n24410, n24411, n24412, 
      n24413, n24414, n24415, n24416, n24417, n24419, n24420, n24421, n24424, 
      n24425, n24426, n24427, n24429, n24430, n24431, n24432, n24433, n24434, 
      n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, 
      n24445, n24446, n24447, n24448, n24449, n24451, n24452, n24453, n24455, 
      n24456, n24457, n24458, n24459, n24460, n24461, n24463, n24464, n24465, 
      n24466, n24467, n24469, n24470, n24471, n24472, n24473, n24474, n24475, 
      n24476, n24477, n24478, n24479, n24481, n24483, n24484, n24485, n24490, 
      n24491, n24492, n24493, n24494, n24495, n24496, n24498, n24499, n24500, 
      n24502, n24504, n24506, n24507, n24509, n24510, n24511, n24514, n24515, 
      n24516, n24517, n24518, n24524, n24525, n24526, n24527, n24528, n24529, 
      n24530, n24531, n24532, n24534, n24535, n24536, n24538, n24539, n24540, 
      n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24550, n24551, 
      n24552, n24553, n24554, n24556, n24557, n24558, n24560, n24561, n24563, 
      n24565, n24566, n24568, n24569, n24571, n24572, n24573, n24574, n24575, 
      n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584, 
      n24585, n24586, n24588, n24589, n24590, n24591, n24592, n24593, n24595, 
      n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24605, 
      n24606, n24607, n24608, n24609, n24610, n24612, n24613, n24614, n24615, 
      n24616, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, 
      n24626, n24627, n24629, n24630, n24631, n24632, n24633, n24634, n24635, 
      n24637, n24638, n24639, n24641, n24643, n24644, n24646, n24647, n24648, 
      n24649, n24650, n24651, n24652, n24655, n24656, n24657, n24658, n24659, 
      n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24668, n24669, 
      n24670, n24671, n24672, n24673, n24674, n24676, n24678, n24679, n24680, 
      n24681, n24683, n24685, n24686, n24687, n24689, n24690, n24691, n24692, 
      n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, 
      n24702, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, 
      n24712, n24713, n24715, n24716, n24717, n24719, n24720, n24721, n24723, 
      n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, 
      n24733, n24734, n24735, n24736, n24737, n24738, n24740, n24741, n24743, 
      n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752, 
      n24753, n24754, n24755, n24757, n24759, n24761, n24762, n24763, n24764, 
      n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24774, 
      n24775, n24776, n24777, n24778, n24779, n24780, n24782, n24783, n24784, 
      n24785, n24786, n24787, n24788, n24789, n24792, n24793, n24794, n24795, 
      n24798, n24799, n24800, n24801, n24802, n24804, n24805, n24806, n24810, 
      n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, 
      n24820, n24821, n24822, n24823, n24824, n24826, n24827, n24828, n24829, 
      n24832, n24833, n24834, n24836, n24838, n24839, n24840, n24841, n24842, 
      n24843, n24844, n24845, n24847, n24849, n24850, n24852, n24853, n24854, 
      n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863, 
      n24864, n24866, n24868, n24869, n24871, n24872, n24873, n24874, n24875, 
      n24876, n24877, n24878, n24879, n24882, n24883, n24884, n24885, n24886, 
      n24887, n24891, n24892, n24894, n24895, n24896, n24897, n24898, n24899, 
      n24900, n24902, n24903, n24904, n24905, n24906, n24907, n24909, n24910, 
      n24912, n24913, n24914, n24915, n24917, n24918, n24919, n24920, n24921, 
      n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, 
      n24931, n24932, n24933, n24935, n24936, n24937, n24938, n24940, n24941, 
      n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950, 
      n24952, n24953, n24954, n24955, n24957, n24958, n24959, n24960, n24961, 
      n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24970, n24971, 
      n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24981, n24982, 
      n24984, n24985, n24987, n24988, n24989, n24990, n24991, n24992, n24994, 
      n24997, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006, 
      n25007, n25008, n25009, n25010, n25011, n25012, n25014, n25015, n25016, 
      n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, 
      n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, 
      n25036, n25037, n25039, n25040, n25041, n25042, n25043, n25044, n25045, 
      n25046, n25047, n25048, n25049, n25051, n25052, n25053, n25054, n25055, 
      n25056, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066, 
      n25067, n25068, n25070, n25071, n25072, n25073, n25074, n25075, n25076, 
      n25077, n25078, n25079, n25080, n25081, n25083, n25085, n25086, n25087, 
      n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, 
      n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, 
      n25106, n25108, n25110, n25111, n25112, n25113, n25114, n25115, n25116, 
      n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, 
      n25127, n25128, n25129, n25132, n25133, n25134, n25135, n25136, n25137, 
      n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, 
      n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, 
      n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, 
      n25166, n25167, n25170, n25171, n25172, n25173, n25174, n25175, n25176, 
      n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, 
      n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, 
      n25195, n25196, n25197, n25198, n25200, n25201, n25202, n25203, n25204, 
      n25206, n25207, n25208, n25210, n25211, n25213, n25214, n25215, n25216, 
      n25217, n25218, n25219, n25220, n25221, n25222, n25224, n25225, n25226, 
      n25229, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, 
      n25239, n25240, n25241, n25242, n25243, n25245, n25246, n25247, n25248, 
      n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, 
      n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, 
      n25267, n25268, n25269, n25270, n25271, n25272, n25274, n25275, n25276, 
      n25277, n25278, n25279, n25280, n25281, n25283, n25284, n25285, n25286, 
      n25288, n25289, n25290, n25291, n25292, n25293, n25295, n25296, n25298, 
      n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25307, n25309, 
      n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318, 
      n25319, n25320, n25322, n25323, n25324, n25326, n25327, n25328, n25329, 
      n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25339, 
      n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349, 
      n25351, n25352, n25353, n25354, n25355, n25358, n25359, n25360, n25361, 
      n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370, 
      n25371, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, 
      n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, 
      n25390, n25392, n25393, n25394, n25395, n25396, n25397, n25399, n25400, 
      n25401, n25402, n25404, n25405, n25406, n25407, n25408, n25409, n25410, 
      n25412, n25416, n25418, n25420, n25421, n25422, n25424, n25425, n25427, 
      n25428, n25429, n25430, n25431, n25433, n25434, n25435, n25436, n25437, 
      n25438, n25439, n25440, n25441, n25443, n25444, n25445, n25447, n25448, 
      n25449, n25450, n25451, n25452, n25454, n25455, n25456, n25457, n25458, 
      n25459, n25460, n25462, n25464, n25466, n25467, n25468, n25469, n25470, 
      n25471, n25472, n25473, n25474, n25476, n25477, n25478, n25479, n25480, 
      n25481, n25482, n25483, n25484, n25486, n25487, n25488, n25489, n25490, 
      n25491, n25495, n25497, n25498, n25499, n25501, n25502, n25503, n25506, 
      n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, 
      n25516, n25517, n25519, n25525, n25526, n25527, n25528, n25529, n25530, 
      n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539, 
      n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, 
      n25549, n25550, n25552, n25553, n25554, n25555, n25556, n25557, n25558, 
      n25559, n25560, n25562, n25563, n25564, n25566, n25567, n25568, n25569, 
      n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25581, n25582, 
      n25583, n25584, n25585, n25586, n25587, n25592, n25593, n25594, n25595, 
      n25596, n25597, n25598, n25600, n25601, n25602, n25603, n25604, n25605, 
      n25606, n25608, n25609, n25611, n25612, n25613, n25614, n25615, n25616, 
      n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25625, n25627, 
      n25628, n25630, n25631, n25633, n25634, n25635, n25636, n25637, n25638, 
      n25639, n25641, n25642, n25643, n25644, n25645, n25647, n25649, n25650, 
      n25651, n25655, n25657, n25658, n25659, n25660, n25661, n25662, n25665, 
      n25666, n25667, n25669, n25670, n25674, n25675, n25676, n25677, n25678, 
      n25679, n25680, n25681, n25682, n25683, n25685, n25686, n25687, n25688, 
      n25689, n25690, n25691, n25692, n25694, n25695, n25696, n25697, n25698, 
      n25699, n25700, n25702, n25705, n25706, n25707, n25708, n25712, n25713, 
      n25714, n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723, 
      n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732, 
      n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742, 
      n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25751, n25753, 
      n25754, n25755, n25756, n25758, n25759, n25760, n25761, n25762, n25764, 
      n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25774, n25775, 
      n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784, 
      n25785, n25787, n25788, n25790, n25792, n25793, n25794, n25795, n25796, 
      n25797, n25798, n25799, n25800, n25801, n25803, n25804, n25805, n25807, 
      n25808, n25809, n25810, n25812, n25813, n25814, n25815, n25817, n25818, 
      n25819, n25820, n25821, n25822, n25825, n25826, n25827, n25828, n25829, 
      n25830, n25831, n25833, n25834, n25835, n25836, n25837, n25838, n25840, 
      n25841, n25842, n25844, n25845, n25846, n25847, n25848, n25849, n25850, 
      n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25860, 
      n25861, n25862, n25865, n25866, n25867, n25868, n25869, n25870, n25871, 
      n25872, n25874, n25875, n25876, n25877, n25878, n25879, n25882, n25883, 
      n25886, n25887, n25888, n25889, n25891, n25892, n25894, n25896, n25897, 
      n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25907, 
      n25910, n25911, n25912, n25914, n25915, n25916, n25917, n25918, n25919, 
      n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928, 
      n25930, n25931, n25933, n25934, n25936, n25937, n25938, n25939, n25940, 
      n25941, n25942, n25943, n25945, n25946, n25947, n25949, n25950, n25951, 
      n25954, n25955, n25956, n25957, n25958, n25959, n25961, n25962, n25964, 
      n25965, n25966, n25967, n25970, n25971, n25972, n25975, n25977, n25978, 
      n25979, n25981, n25982, n25983, n25984, n25985, n25986, n25988, n25989, 
      n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25998, n25999, 
      n26000, n26001, n26003, n26004, n26005, n26006, n26008, n26009, n26010, 
      n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, 
      n26020, n26021, n26022, n26023, n26024, n26026, n26027, n26028, n26029, 
      n26030, n26031, n26032, n26034, n26035, n26036, n26037, n26038, n26039, 
      n26041, n26042, n26045, n26048, n26050, n26051, n26052, n26053, n26054, 
      n26055, n26056, n26058, n26059, n26060, n26061, n26063, n26065, n26066, 
      n26067, n26068, n26070, n26071, n26072, n26073, n26074, n26075, n26076, 
      n26077, n26078, n26079, n26081, n26083, n26084, n26085, n26086, n26088, 
      n26089, n26090, n26092, n26093, n26094, n26095, n26096, n26097, n26098, 
      n26099, n26101, n26103, n26104, n26105, n26106, n26107, n26108, n26109, 
      n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, 
      n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26128, 
      n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26137, n26138, 
      n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, 
      n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157, 
      n26158, n26160, n26161, n26162, n26163, n26165, n26166, n26167, n26168, 
      n26169, n26171, n26172, n26173, n26176, n26177, n26178, n26179, n26180, 
      n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26190, 
      n26191, n26192, n26194, n26195, n26196, n26197, n26198, n26200, n26201, 
      n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, 
      n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221, 
      n26222, n26223, n26224, n26225, n26227, n26228, n26229, n26230, n26231, 
      n26232, n26233, n26234, n26236, n26237, n26238, n26239, n26240, n26241, 
      n26242, n26243, n26244, n26245, n26246, n26247, n26249, n26250, n26251, 
      n26252, n26253, n26254, n26255, n26257, n26258, n26259, n26260, n26261, 
      n26262, n26263, n26264, n26265, n26266, n26268, n26269, n26270, n26272, 
      n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281, 
      n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290, 
      n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26299, n26301, 
      n26302, n26303, n26304, n26305, n26307, n26308, n26309, n26310, n26311, 
      n26312, n26313, n26314, n26316, n26317, n26318, n26319, n26320, n26321, 
      n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331, 
      n26332, n26333, n26334, n26335, n26336, n26338, n26339, n26340, n26341, 
      n26342, n26343, n26344, n26346, n26347, n26348, n26349, n26350, n26352, 
      n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, 
      n26363, n26364, n26365, n26366, n26368, n26369, n26370, n26371, n26372, 
      n26373, n26374, n26375, n26376, n26377, n26379, n26380, n26381, n26382, 
      n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, 
      n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400, 
      n26401, n26402, n26403, n26404, n26405, n26407, n26408, n26409, n26410, 
      n26411, n26412, n26413, n26415, n26417, n26418, n26419, n26420, n26421, 
      n26422, n26424, n26425, n26426, n26427, n26428, n26429, n26431, n26432, 
      n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441, 
      n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450, 
      n26451, n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, 
      n26461, n26462, n26463, n26464, n26465, n26466, n26468, n26470, n26471, 
      n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26480, n26481, 
      n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, 
      n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499, 
      n26500, n26502, n26503, n26504, n26508, n26509, n26510, n26511, n26512, 
      n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, 
      n26522, n26523, n26525, n26526, n26527, n26528, n26529, n26530, n26531, 
      n26532, n26536, n26537, n26538, n26539, n26541, n26542, n26544, n26545, 
      n26547, n26548, n26550, n26551, n26553, n26554, n26555, n26556, n26557, 
      n26558, n26559, n26560, n26561, n26562, n26564, n26565, n26566, n26567, 
      n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26577, 
      n26578, n26579, n26580, n26581, n26582, n26584, n26585, n26587, n26588, 
      n26590, n26591, n26593, n26594, n26595, n26596, n26597, n26598, n26599, 
      n26600, n26601, n26602, n26605, n26606, n26607, n26608, n26609, n26610, 
      n26612, n26614, n26618, n26619, n26621, n26622, n26623, n26624, n26625, 
      n26626, n26627, n26628, n26630, n26632, n26634, n26635, n26636, n26637, 
      n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26647, 
      n26648, n26650, n26651, n26652, n26653, n26655, n26657, n26659, n26660, 
      n26661, n26662, n26663, n26665, n26666, n26667, n26668, n26670, n26671, 
      n26672, n26674, n26675, n26678, n26679, n26682, n26684, n26686, n26687, 
      n26688, n26689, n26691, n26692, n26694, n26695, n26696, n26697, n26698, 
      n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707, 
      n26708, n26709, n26710, n26713, n26717, n26718, n26719, n26720, n26721, 
      n26722, n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731, 
      n26732, n26733, n26734, n26737, n26738, n26740, n26741, n26743, n26744, 
      n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26754, 
      n26755, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, 
      n26766, n26767, n26768, n26769, n26770, n26772, n26773, n26774, n26775, 
      n26776, n26777, n26778, n26779, n26780, n26783, n26784, n26785, n26786, 
      n26787, n26788, n26789, n26790, n26791, n26793, n26794, n26795, n26796, 
      n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, 
      n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26815, 
      n26816, n26817, n26818, n26819, n26822, n26823, n26824, n26825, n26826, 
      n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, 
      n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, 
      n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26856, 
      n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, 
      n26866, n26868, n26869, n26870, n26871, n26872, n26876, n26877, n26878, 
      n26879, n26882, n26885, n26887, n26888, n26889, n26890, n26892, n26893, 
      n26895, n26897, n26898, n26899, n26901, n26902, n26903, n26905, n26906, 
      n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915, 
      n26916, n26918, n26919, n26920, n26921, n26922, n26923, n26926, n26927, 
      n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936, 
      n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945, 
      n26946, n26948, n26950, n26951, n26952, n26953, n26954, n26955, n26956, 
      n26957, n26958, n26959, n26961, n26962, n26963, n26964, n26965, n26966, 
      n26967, n26968, n26970, n26972, n26973, n26974, n26975, n26976, n26977, 
      n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, 
      n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, 
      n26996, n26998, n26999, n27000, n27001, n27004, n27006, n27007, n27009, 
      n27010, n27011, n27013, n27014, n27015, n27017, n27018, n27020, n27021, 
      n27023, n27024, n27026, n27027, n27028, n27029, n27030, n27031, n27032, 
      n27033, n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042, 
      n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27051, n27052, 
      n27053, n27054, n27055, n27056, n27057, n27059, n27060, n27061, n27062, 
      n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071, 
      n27072, n27073, n27076, n27078, n27079, n27080, n27081, n27083, n27084, 
      n27085, n27087, n27088, n27089, n27090, n27092, n27093, n27094, n27095, 
      n27096, n27097, n27098, n27099, n27102, n27103, n27106, n27107, n27108, 
      n27109, n27110, n27111, n27113, n27114, n27115, n27116, n27118, n27119, 
      n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, 
      n27130, n27131, n27133, n27135, n27137, n27138, n27139, n27140, n27141, 
      n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, 
      n27151, n27152, n27153, n27154, n27155, n27158, n27159, n27161, n27163, 
      n27164, n27165, n27166, n27167, n27169, n27170, n27171, n27172, n27174, 
      n27175, n27176, n27178, n27180, n27181, n27182, n27184, n27185, n27187, 
      n27189, n27192, n27193, n27194, n27196, n27197, n27198, n27199, n27200, 
      n27201, n27203, n27204, n27205, n27206, n27207, n27211, n27213, n27214, 
      n27215, n27218, n27220, n27221, n27224, n27225, n27226, n27228, n27229, 
      n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, 
      n27240, n27242, n27244, n27245, n27247, n27248, n27249, n27250, n27251, 
      n27252, n27253, n27255, n27256, n27257, n27258, n27259, n27263, n27265, 
      n27266, n27267, n27269, n27270, n27271, n27272, n27273, n27274, n27275, 
      n27276, n27278, n27279, n27282, n27283, n27284, n27285, n27286, n27287, 
      n27288, n27289, n27291, n27292, n27295, n27296, n27297, n27298, n27299, 
      n27300, n27302, n27304, n27305, n27306, n27307, n27310, n27311, n27312, 
      n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27324, 
      n27325, n27326, n27328, n27329, n27331, n27332, n27333, n27334, n27335, 
      n27336, n27337, n27338, n27341, n27342, n27343, n27344, n27345, n27346, 
      n27347, n27348, n27349, n27350, n27351, n27353, n27354, n27356, n27357, 
      n27358, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27368, 
      n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377, 
      n27378, n27379, n27381, n27382, n27383, n27384, n27385, n27386, n27387, 
      n27388, n27389, n27390, n27391, n27392, n27393, n27395, n27397, n27398, 
      n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407, 
      n27408, n27409, n27410, n27411, n27412, n27413, n27415, n27416, n27417, 
      n27419, n27420, n27421, n27422, n27424, n27426, n27428, n27429, n27430, 
      n27431, n27433, n27434, n27435, n27436, n27438, n27440, n27441, n27444, 
      n27445, n27446, n27447, n27448, n27449, n27451, n27452, n27453, n27455, 
      n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464, 
      n27465, n27466, n27467, n27469, n27470, n27471, n27472, n27473, n27474, 
      n27475, n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, 
      n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493, 
      n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, 
      n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27511, n27513, 
      n27514, n27515, n27516, n27517, n27518, n27520, n27521, n27522, n27523, 
      n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532, 
      n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541, 
      n27542, n27543, n27546, n27547, n27548, n27549, n27550, n27551, n27552, 
      n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561, 
      n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570, 
      n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579, 
      n27580, n27581, n27583, n27584, n27585, n27586, n27587, n27588, n27589, 
      n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598, 
      n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, 
      n27609, n27611, n27612, n27613, n27614, n27615, n27617, n27618, n27619, 
      n27620, n27621, n27622, n27624, n27626, n27627, n27628, n27630, n27631, 
      n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640, 
      n27641, n27642, n27643, n27645, n27646, n27647, n27648, n27649, n27650, 
      n27651, n27652, n27653, n27654, n27655, n27657, n27658, n27659, n27661, 
      n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27671, 
      n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680, 
      n27681, n27683, n27685, n27686, n27687, n27688, n27689, n27690, n27692, 
      n27695, n27696, n27697, n27698, n27700, n27701, n27703, n27704, n27705, 
      n27706, n27707, n27709, n27710, n27711, n27712, n27713, n27714, n27715, 
      n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724, 
      n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733, 
      n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743, 
      n27745, n27746, n27748, n27749, n27750, n27751, n27753, n27754, n27755, 
      n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764, 
      n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773, 
      n27774, n27776, n27777, n27778, n27779, n27781, n27782, n27784, n27785, 
      n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794, 
      n27795, n27796, n27797, n27798, n27799, n27800, n27802, n27803, n27804, 
      n27805, n27806, n27807, n27808, n27809, n27810, n27812, n27813, n27815, 
      n27816, n27817, n27818, n27819, n27820, n27822, n27823, n27825, n27826, 
      n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, 
      n27836, n27837, n27839, n27840, n27841, n27842, n27843, n27844, n27845, 
      n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855, 
      n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864, 
      n27865, n27866, n27867, n27868, n27870, n27871, n27872, n27873, n27874, 
      n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883, 
      n27884, n27885, n27887, n27888, n27889, n27890, n27891, n27892, n27893, 
      n27894, n27895, n27896, n27897, n27898, n27900, n27901, n27902, n27903, 
      n27904, n27906, n27907, n27908, n27909, n27910, n27911, n27913, n27914, 
      n27915, n27917, n27918, n27919, n27920, n27921, n27925, n27926, n27927, 
      n27928, n27929, n27930, n27932, n27934, n27935, n27936, n27938, n27940, 
      n27941, n27942, n27943, n27944, n27946, n27948, n27951, n27955, n27956, 
      n27957, n27958, n27959, n27962, n27963, n27964, n27966, n27967, n27969, 
      n27970, n27972, n27973, n27974, n27976, n27978, n27979, n27980, n27981, 
      n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990, 
      n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998, n28001, 
      n28002, n28004, n28006, n28007, n28008, n28009, n28010, n28011, n28012, 
      n28013, n28014, n28015, n28017, n28021, n28022, n28023, n28024, n28025, 
      n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034, 
      n28035, n28036, n28038, n28039, n28040, n28041, n28042, n28043, n28045, 
      n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28056, 
      n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065, 
      n28066, n28067, n28068, n28069, n28073, n28074, n28075, n28079, n28080, 
      n28081, n28082, n28083, n28085, n28086, n28087, n28089, n28091, n28093, 
      n28095, n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105, 
      n28106, n28107, n28108, n28109, n28111, n28112, n28113, n28114, n28115, 
      n28117, n28118, n28119, n28122, n28123, n28124, n28125, n28126, n28127, 
      n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28137, n28138, 
      n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147, 
      n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156, 
      n28157, n28159, n28161, n28162, n28163, n28164, n28165, n28167, n28168, 
      n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178, 
      n28179, n28180, n28181, n28182, n28184, n28185, n28186, n28187, n28188, 
      n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28197, n28199, 
      n28200, n28202, n28203, n28204, n28205, n28206, n28207, n28209, n28210, 
      n28212, n28213, n28214, n28215, n28216, n28217, n28219, n28220, n28221, 
      n28222, n28223, n28224, n28226, n28227, n28228, n28229, n28230, n28231, 
      n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28240, n28242, 
      n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251, 
      n28255, n28256, n28257, n28258, n28259, n28260, n28262, n28263, n28264, 
      n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273, 
      n28274, n28276, n28278, n28279, n28281, n28282, n28283, n28284, n28285, 
      n28286, n28287, n28288, n28289, n28290, n28291, n28293, n28297, n28298, 
      n28299, n28301, n28302, n28304, n28305, n28306, n28307, n28308, n28309, 
      n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318, 
      n28319, n28320, n28322, n28323, n28324, n28325, n28326, n28327, n28328, 
      n28330, n28331, n28332, n28333, n28335, n28336, n28337, n28338, n28339, 
      n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348, 
      n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357, 
      n28358, n28359, n28360, n28361, n28362, n28364, n28365, n28366, n28368, 
      n28369, n28370, n28372, n28373, n28375, n28376, n28377, n28378, n28380, 
      n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28389, n28390, 
      n28391, n28392, n28394, n28395, n28396, n28398, n28399, n28400, n28401, 
      n28402, n28403, n28406, n28408, n28409, n28410, n28411, n28412, n28414, 
      n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423, 
      n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28433, 
      n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28442, n28443, 
      n28444, n28445, n28448, n28450, n28452, n28453, n28454, n28455, n28456, 
      n28457, n28458, n28460, n28463, n28464, n28465, n28466, n28467, n28468, 
      n28470, n28471, n28473, n28475, n28477, n28478, n28479, n28480, n28483, 
      n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, 
      n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, 
      n28502, n28503, n28504, n28505, n28507, n28508, n28509, n28510, n28513, 
      n28514, n28515, n28516, n28518, n28520, n28521, n28522, n28523, n28524, 
      n28525, n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535, 
      n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545, 
      n28546, n28547, n28548, n28549, n28550, n28551, n28553, n28554, n28555, 
      n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, 
      n28565, n28568, n28569, n28570, n28571, n28573, n28574, n28575, n28576, 
      n28577, n28578, n28579, n28580, n28583, n28584, n28585, n28586, n28587, 
      n28589, n28590, n28591, n28592, n28594, n28595, n28596, n28598, n28601, 
      n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611, 
      n28612, n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621, 
      n28622, n28623, n28625, n28626, n28627, n28630, n28631, n28632, n28633, 
      n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28643, 
      n28644, n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, 
      n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28664, 
      n28665, n28666, n28669, n28670, n28671, n28673, n28674, n28675, n28676, 
      n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28685, n28686, 
      n28689, n28690, n28691, n28692, n28693, n28695, n28696, n28697, n28698, 
      n28699, n28700, n28704, n28705, n28707, n28708, n28709, n28710, n28712, 
      n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721, 
      n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730, 
      n28732, n28733, n28735, n28736, n28738, n28739, n28740, n28742, n28743, 
      n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752, 
      n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28761, n28762, 
      n28763, n28764, n28765, n28767, n28768, n28769, n28770, n28771, n28772, 
      n28773, n28775, n28776, n28777, n28778, n28779, n28780, n28782, n28783, 
      n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28793, n28794, 
      n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803, 
      n28804, n28805, n28806, n28807, n28808, n28811, n28812, n28813, n28814, 
      n28815, n28817, n28819, n28820, n28821, n28822, n28823, n28824, n28825, 
      n28826, n28827, n28828, n28829, n28830, n28831, n28834, n28835, n28836, 
      n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845, 
      n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28857, 
      n28858, n28859, n28860, n28862, n28863, n28864, n28865, n28866, n28867, 
      n28868, n28869, n28870, n28871, n28873, n28874, n28876, n28878, n28880, 
      n28882, n28883, n28885, n28886, n28887, n28888, n28889, n28891, n28892, 
      n28893, n28894, n28895, n28896, n28898, n28899, n28900, n28901, n28902, 
      n28903, n28904, n28905, n28906, n28907, n28909, n28910, n28912, n28913, 
      n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28923, n28924, 
      n28925, n28927, n28928, n28930, n28931, n28933, n28934, n28935, n28940, 
      n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951, 
      n28953, n28954, n28955, n28957, n28958, n28959, n28960, n28961, n28962, 
      n28963, n28964, n28966, n28967, n28968, n28969, n28970, n28971, n28972, 
      n28973, n28975, n28976, n28977, n28978, n28979, n28980, n28982, n28983, 
      n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992, 
      n28993, n28994, n28996, n28997, n28998, n28999, n29000, n29001, n29002, 
      n29003, n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012, 
      n29014, n29015, n29016, n29017, n29019, n29021, n29022, n29023, n29024, 
      n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29033, n29034, 
      n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043, 
      n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, 
      n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29063, 
      n29064, n29065, n29066, n29067, n29068, n29070, n29071, n29072, n29073, 
      n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082, 
      n29083, n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092, 
      n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29102, 
      n29103, n29104, n29105, n29107, n29108, n29109, n29110, n29111, n29113, 
      n29114, n29115, n29119, n29120, n29121, n29122, n29123, n29124, n29125, 
      n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134, 
      n29135, n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144, 
      n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153, 
      n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163, 
      n29164, n29165, n29166, n29167, n29168, n29169, n29171, n29173, n29174, 
      n29175, n29176, n29180, n29181, n29182, n29183, n29184, n29185, n29187, 
      n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196, 
      n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205, 
      n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29214, n29217, 
      n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29226, n29228, 
      n29229, n29230, n29231, n29232, n29233, n29234, n29236, n29237, n29238, 
      n29239, n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248, 
      n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29257, n29258, 
      n29260, n29262, n29263, n29265, n29266, n29267, n29268, n29269, n29270, 
      n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279, 
      n29280, n29281, n29282, n29284, n29285, n29286, n29287, n29289, n29290, 
      n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299, 
      n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29309, 
      n29310, n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319, 
      n29320, n29321, n29323, n29324, n29325, n29326, n29327, n29328, n29329, 
      n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338, 
      n29339, n29340, n29341, n29342, n29344, n29345, n29346, n29347, n29348, 
      n29349, n29350, n29351, n29353, n29354, n29355, n29356, n29357, n29358, 
      n29359, n29360, n29361, n29362, n29363, n29365, n29367, n29368, n29369, 
      n29370, n29371, n29372, n29373, n29375, n29377, n29378, n29379, n29380, 
      n29381, n29382, n29383, n29384, n29385, n29389, n29390, n29391, n29392, 
      n29393, n29394, n29396, n29397, n29398, n29399, n29400, n29401, n29402, 
      n29403, n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, 
      n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, 
      n29422, n29423, n29424, n29425, n29426, n29427, n29430, n29431, n29432, 
      n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441, 
      n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450, 
      n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459, 
      n29461, n29462, n29463, n29464, n29466, n29467, n29468, n29469, n29470, 
      n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480, 
      n29481, n29482, n29483, n29485, n29486, n29488, n29489, n29490, n29491, 
      n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501, 
      n29502, n29503, n29504, n29505, n29506, n29509, n29510, n29511, n29512, 
      n29513, n29514, n29515, n29516, n29517, n29519, n29520, n29521, n29522, 
      n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531, 
      n29532, n29533, n29534, n29535, n29536, n29538, n29539, n29540, n29541, 
      n29542, n29543, n29546, n29547, n29548, n29549, n29550, n29551, n29552, 
      n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29562, 
      n29563, n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572, 
      n29573, n29574, n29575, n29577, n29578, n29579, n29580, n29581, n29583, 
      n29586, n29587, n29591, n29592, n29593, n29595, n29596, n29597, n29598, 
      n29599, n29600, n29601, n29602, n29604, n29605, n29607, n29608, n29610, 
      n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, 
      n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629, 
      n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638, 
      n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648, 
      n29649, n29652, n29654, n29656, n29657, n29658, n29659, n29660, n29661, 
      n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670, 
      n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679, 
      n29680, n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689, 
      n29690, n29692, n29693, n29694, n29696, n29697, n29698, n29699, n29700, 
      n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, 
      n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, 
      n29719, n29720, n29721, n29722, n29723, n29725, n29726, n29727, n29728, 
      n29729, n29730, n29731, n29732, n29733, n29735, n29736, n29737, n29739, 
      n29740, n29741, n29747, n29749, n29750, n29751, n29752, n29753, n29754, 
      n29755, n29756, n29758, n29759, n29760, n29761, n29762, n29763, n29764, 
      n29767, n29768, n29769, n29770, n29771, n29774, n29775, n29776, n29777, 
      n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29787, n29788, 
      n29789, n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797, 
      n29798, n29799, n29800, n29801, n29802, n29803, n29805, n29806, n29807, 
      n29808, n29809, n29810, n29811, n29812, n29813, n29815, n29816, n29817, 
      n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29827, 
      n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836, 
      n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845, 
      n29846, n29847, n29849, n29851, n29852, n29854, n29855, n29856, n29857, 
      n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866, 
      n29867, n29869, n29870, n29871, n29873, n29874, n29875, n29876, n29877, 
      n29879, n29880, n29881, n29883, n29884, n29885, n29887, n29888, n29889, 
      n29890, n29892, n29895, n29896, n29897, n29898, n29899, n29900, n29901, 
      n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910, 
      n29911, n29912, n29913, n29914, n29915, n29916, n29918, n29919, n29920, 
      n29922, n29923, n29924, n29925, n29927, n29928, n29929, n29930, n29931, 
      n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939, n29940, 
      n29941, n29942, n29943, n29946, n29947, n29948, n29949, n29951, n29952, 
      n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961, 
      n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29970, n29971, 
      n29973, n29974, n29975, n29977, n29978, n29979, n29980, n29981, n29982, 
      n29983, n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992, 
      n29993, n29994, n29996, n29997, n29998, n30000, n30001, n30002, n30003, 
      n30004, n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013, 
      n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022, 
      n30023, n30024, n30025, n30026, n30027, n30028, n30030, n30031, n30032, 
      n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041, 
      n30042, n30043, n30045, n30046, n30047, n30048, n30049, n30051, n30052, 
      n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30062, 
      n30063, n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072, 
      n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081, 
      n30083, n30084, n30085, n30086, n30087, n30089, n30090, n30091, n30092, 
      n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101, 
      n30102, n30104, n30105, n30106, n30107, n30109, n30110, n30111, n30112, 
      n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30122, 
      n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134, 
      n30135, n30136, n30138, n30139, n30140, n30141, n30143, n30144, n30145, 
      n30146, n30147, n30150, n30152, n30153, n30154, n30155, n30156, n30158, 
      n30159, n30160, n30161, n30162, n30163, n30165, n30166, n30168, n30169, 
      n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178, 
      n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187, 
      n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198, 
      n30199, n30201, n30203, n30204, n30205, n30206, n30207, n30210, n30211, 
      n30212, n30213, n30214, n30215, n30216, n30217, n30220, n30221, n30222, 
      n30223, n30225, n30228, n30229, n30230, n30231, n30232, n30233, n30237, 
      n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246, 
      n30247, n30248, n30249, n30250, n30252, n30253, n30255, n30256, n30257, 
      n30258, n30259, n30260, n30261, n30262, n30263, n30272, n30274, n30275, 
      n30276, n30279, n30280, n30282, n30283, n30284, n30285, n30288, n30290, 
      n30292, n30293, n30295, n30299, n30302, n30304, n30306, n30311, n30315, 
      n30317, n30318, n30320, n30321, n30322, n30323, n30324, n30326, n30329, 
      n30330, n30333, n30334, n30335, n30336, n30338, n30339, n30340, n30342, 
      n30345, n30347, n30348, n30350, n30352, n30353, n30354, n30355, n30356, 
      n30357, n30358, n30360, n30363, n30364, n30365, n30366, n30368, n30369, 
      n30370, n30371, n30372, n30373, n30377, n30378, n30379, n30380, n30381, 
      n30384, n30385, n30386, n30388, n30389, n30391, n30392, n30393, n30394, 
      n30396, n30397, n30399, n30400, n30401, n30402, n30403, n30404, n30405, 
      n30406, n30408, n30409, n30410, n30412, n30413, n30414, n30416, n30417, 
      n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30427, n30429, 
      n30431, n30432, n30433, n30434, n30435, n30436, n30440, n30442, n30443, 
      n30444, n30445, n30446, n30447, n30448, n30450, n30451, n30452, n30453, 
      n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30463, 
      n30464, n30465, n30468, n30469, n30470, n30471, n30473, n30475, n30478, 
      n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487, 
      n30488, n30489, n30494, n30496, n30499, n30500, n30502, n30503, n30504, 
      n30506, n30507, n30509, n30512, n30519, n30520, n30524, n30526, n30528, 
      n30529, n30530, n30534, n30539, n30541, n30542, n30544, n30546, n30547, 
      n30548, n30550, n30551, n30554, n30555, n30556, n30558, n30560, n30561, 
      n30562, n30565, n30568, n30571, n30572, n30574, n30577, n30578, n30580, 
      n30581, n30582, n30584, n30585, n30587, n30588, n30594, n30595, n30596, 
      n30597, n30598, n30599, n30602, n30603, n30607, n30608, n30609, n30610, 
      n30611, n30612, n30613, n30615, n30616, n30617, n30619, n30621, n30623, 
      n30625, n30626, n30629, n30631, n30632, n30633, n30635, n30636, n30642, 
      n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30651, n30652, 
      n30653, n30655, n30656, n30657, n30659, n30661, n30663, n30664, n30665, 
      n30667, n30668, n30671, n30674, n30675, n30676, n30677, n30678, n30680, 
      n30682, n30684, n30687, n30688, n30689, n30694, n30695, n30696, n30698, 
      n30699, n30700, n30701, n30702, n30704, n30705, n30706, n30709, n30711, 
      n30712, n30714, n30715, n30716, n30720, n30722, n30724, n30725, n30726, 
      n30727, n30728, n30730, n30731, n30732, n30733, n30734, n30736, n30738, 
      n30740, n30741, n30745, n30746, n30747, n30748, n30756, n30757, n30758, 
      n30761, n30764, n30766, n30768, n30771, n30773, n30775, n30776, n30778, 
      n30780, n30781, n30785, n30786, n30788, n30789, n30793, n30794, n30795, 
      n30796, n30798, n30799, n30800, n30803, n30805, n30806, n30808, n30811, 
      n30813, n30815, n30817, n30818, n30819, n30822, n30824, n30825, n30826, 
      n30828, n30831, n30833, n30835, n30837, n30838, n30839, n30840, n30842, 
      n30843, n30844, n30845, n30846, n30847, n30849, n30850, n30851, n30853, 
      n30854, n30856, n30857, n30858, n30859, n30862, n30863, n30865, n30871, 
      n30872, n30874, n30877, n30878, n30881, n30883, n30886, n30888, n30890, 
      n30891, n30893, n30894, n30895, n30897, n30898, n30900, n30905, n30907, 
      n30908, n30910, n30913, n30914, n30915, n30917, n30925, n30927, n30928, 
      n30929, n30930, n30931, n30933, n30934, n30936, n30937, n30938, n30939, 
      n30941, n30942, n30944, n30945, n30946, n30947, n30948, n30949, n30950, 
      n30951, n30952, n30953, n30955, n30956, n30957, n30958, n30959, n30960, 
      n30962, n30963, n30964, n30965, n30966, n30967, n30971, n30972, n30973, 
      n30974, n30976, n30980, n30981, n30982, n30983, n30986, n30988, n30989, 
      n30990, n30991, n30993, n30994, n30995, n30996, n31000, n31001, n31002, 
      n31003, n31004, n31005, n31006, n31010, n31012, n31014, n31015, n31016, 
      n31017, n31018, n31019, n31020, n31022, n31023, n31025, n31027, n31028, 
      n31030, n31031, n31034, n31035, n31036, n31037, n31038, n31042, n31043, 
      n31044, n31045, n31046, n31047, n31048, n31049, n31052, n31055, n31059, 
      n31060, n31061, n31062, n31065, n31070, n31073, n31074, n31075, n31077, 
      n31078, n31079, n31080, n31081, n31082, n31086, n31087, n31088, n31089, 
      n31090, n31091, n31092, n31093, n31094, n31095, n31098, n31102, n31103, 
      n31107, n31108, n31110, n31112, n31114, n31115, n31116, n31118, n31119, 
      n31120, n31121, n31122, n31123, n31124, n31125, n31127, n31129, n31130, 
      n31131, n31132, n31133, n31137, n31138, n31139, n31143, n31144, n31146, 
      n31147, n31149, n31150, n31151, n31152, n31154, n31156, n31157, n31158, 
      n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31168, n31170, 
      n31173, n31175, n31177, n31178, n31179, n31180, n31181, n31183, n31184, 
      n31185, n31191, n31192, n31194, n31196, n31197, n31198, n31199, n31200, 
      n31202, n31204, n31205, n31206, n31207, n31211, n31212, n31213, n31214, 
      n31215, n31218, n31220, n31222, n31223, n31225, n31226, n31227, n31230, 
      n31231, n31233, n31234, n31235, n31236, n31237, n31238, n31240, n31242, 
      n31245, n31247, n31248, n31249, n31250, n31252, n31253, n31254, n31257, 
      n31258, n31261, n31263, n31264, n31267, n31268, n31269, n31270, n31271, 
      n31272, n31273, n31274, n31275, n31277, n31278, n31279, n31280, n31281, 
      n31283, n31284, n31287, n31289, n31290, n31292, n31293, n31294, n31295, 
      n31296, n31298, n31299, n31300, n31302, n31304, n31305, n31307, n31310, 
      n31311, n31312, n31313, n31314, n31318, n31319, n31320, n31321, n31322, 
      n31325, n31326, n31327, n31328, n31329, n31331, n31332, n31334, n31335, 
      n31339, n31340, n31341, n31343, n31345, n31346, n31347, n31348, n31349, 
      n31350, n31351, n31352, n31353, n31355, n31356, n31357, n31358, n31359, 
      n31360, n31361, n31362, n31364, n31365, n31366, n31367, n31369, n31370, 
      n31371, n31374, n31375, n31376, n31377, n31378, n31379, n31381, n31383, 
      n31385, n31386, n31388, n31389, n31390, n31393, n31396, n31398, n31399, 
      n31400, n31401, n31403, n31404, n31406, n31407, n31410, n31412, n31414, 
      n31416, n31418, n31421, n31424, n31425, n31426, n31427, n31428, n31430, 
      n31432, n31433, n31437, n31438, n31441, n31442, n31443, n31444, n31445, 
      n31446, n31447, n31452, n31453, n31455, n31457, n31458, n31459, n31461, 
      n31464, n31465, n31466, n31470, n31471, n31473, n31474, n31475, n31476, 
      n31477, n31480, n31481, n31483, n31484, n31485, n31486, n31488, n31490, 
      n31492, n31494, n31495, n31496, n31498, n31499, n31500, n31502, n31504, 
      n31505, n31507, n31508, n31509, n31511, n31512, n31513, n31515, n31516, 
      n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525, 
      n31526, n31527, n31528, n31529, n31530, n31532, n31533, n31534, n31535, 
      n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31545, n31546, 
      n31547, n31548, n31549, n31550, n31551, n31552, n31554, n31555, n31557, 
      n31558, n31559, n31562, n31563, n31564, n31565, n31566, n31568, n31569, 
      n31570, n31571, n31573, n31574, n31575, n31576, n31579, n31580, n31581, 
      n31582, n31583, n31584, n31585, n31586, n31587, n31591, n31594, n31595, 
      n31596, n31597, n31598, n31599, n31601, n31602, n31603, n31604, n31605, 
      n31606, n31607, n31608, n31611, n31612, n31615, n31616, n31617, n31618, 
      n31619, n31620, n31621, n31622, n31624, n31625, n31626, n31627, n31628, 
      n31629, n31630, n31633, n31634, n31636, n31637, n31638, n31640, n31643, 
      n31644, n31647, n31648, n31649, n31650, n31651, n31652, n31654, n31655, 
      n31656, n31657, n31660, n31661, n31662, n31663, n31664, n31665, n31667, 
      n31668, n31669, n31670, n31672, n31673, n31678, n31679, n31680, n31682, 
      n31683, n31684, n31685, n31688, n31689, n31692, n31693, n31695, n31696, 
      n31697, n31698, n31699, n31701, n31702, n31704, n31705, n31707, n31708, 
      n31710, n31711, n31712, n31713, n31714, n31716, n31717, n31718, n31719, 
      n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31731, 
      n31734, n31735, n31736, n31737, n31739, n31743, n31744, n31745, n31748, 
      n31749, n31751, n31752, n31755, n31759, n31760, n31762, n31764, n31765, 
      n31766, n31767, n31769, n31771, n31772, n31773, n31774, n31775, n31777, 
      n31778, n31779, n31780, n31781, n31782, n31784, n31785, n31786, n31787, 
      n31788, n31790, n31791, n31794, n31795, n31796, n31797, n31798, n31799, 
      n31801, n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812, 
      n31815, n31816, n31820, n31821, n31822, n31823, n31824, n31825, n31827, 
      n31829, n31830, n31831, n31832, n31835, n31836, n31838, n31840, n31841, 
      n31842, n31843, n31845, n31846, n31847, n31848, n31849, n31851, n31852, 
      n31854, n31855, n31857, n31859, n31860, n31861, n31862, n31863, n31867, 
      n31869, n31871, n31872, n31875, n31876, n31880, n31882, n31883, n31887, 
      n31888, n31889, n31891, n31893, n31895, n31897, n31898, n31899, n31900, 
      n31904, n31906, n31908, n31909, n31911, n31912, n31913, n31914, n31916, 
      n31917, n31918, n31919, n31920, n31921, n31924, n31925, n31926, n31927, 
      n31931, n31932, n31933, n31934, n31937, n31939, n31940, n31941, n31942, 
      n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31951, n31953, 
      n31954, n31955, n31958, n31959, n31960, n31963, n31964, n31965, n31966, 
      n31967, n31968, n31971, n31972, n31975, n31976, n31978, n31980, n31982, 
      n31983, n31984, n31985, n31986, n31987, n31994, n31996, n31997, n31999, 
      n32001, n32002, n32003, n32004, n32005, n32006, n32009, n32010, n32011, 
      n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020, 
      n32021, n32022, n32024, n32025, n32026, n32032, n32033, n32035, n32036, 
      n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32049, 
      n32050, n32051, n32052, n32053, n32054, n32056, n32057, n32059, n32060, 
      n32061, n32062, n32063, n32064, n32068, n32069, n32071, n32072, n32073, 
      n32075, n32076, n32077, n32079, n32080, n32081, n32083, n32084, n32085, 
      n32087, n32089, n32090, n32091, n32092, n32093, n32095, n32096, n32097, 
      n32099, n32101, n32103, n32105, n32106, n32107, n32109, n32110, n32111, 
      n32113, n32114, n32118, n32120, n32122, n32123, n32125, n32126, n32127, 
      n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136, 
      n32137, n32138, n32141, n32142, n32146, n32149, n32150, n32151, n32152, 
      n32153, n32154, n32156, n32157, n32158, n32159, n32160, n32161, n32162, 
      n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32172, 
      n32174, n32175, n32176, n32178, n32181, n32182, n32183, n32184, n32185, 
      n32186, n32188, n32189, n32190, n32191, n32192, n32193, n32195, n32196, 
      n32197, n32200, n32202, n32203, n32204, n32205, n32206, n32207, n32208, 
      n32209, n32210, n32211, n32215, n32216, n32217, n32218, n32219, n32221, 
      n32223, n32226, n32227, n32228, n32230, n32232, n32233, n32234, n32235, 
      n32236, n32239, n32243, n32245, n32246, n32247, n32248, n32250, n32251, 
      n32253, n32255, n32256, n32258, n32259, n32260, n32261, n32262, n32263, 
      n32266, n32267, n32268, n32270, n32273, n32274, n32275, n32276, n32278, 
      n32279, n32280, n32282, n32283, n32284, n32286, n32288, n32290, n32291, 
      n32292, n32293, n32294, n32297, n32298, n32301, n32302, n32303, n32304, 
      n32306, n32308, n32309, n32310, n32312, n32313, n32314, n32315, n32317, 
      n32318, n32319, n32322, n32324, n32325, n32326, n32327, n32331, n32332, 
      n32333, n32335, n32337, n32338, n32339, n32340, n32343, n32344, n32345, 
      n32346, n32347, n32348, n32349, n32351, n32352, n32353, n32354, n32355, 
      n32358, n32359, n32360, n32361, n32362, n32363, n32365, n32366, n32367, 
      n32368, n32369, n32370, n32372, n32374, n32375, n32376, n32377, n32380, 
      n32382, n32383, n32385, n32386, n32387, n32388, n32389, n32390, n32391, 
      n32394, n32396, n32397, n32398, n32400, n32401, n32402, n32403, n32404, 
      n32406, n32407, n32408, n32410, n32411, n32412, n32413, n32415, n32418, 
      n32419, n32420, n32423, n32424, n32425, n32427, n32430, n32431, n32432, 
      n32433, n32434, n32436, n32440, n32441, n32442, n32443, n32444, n32446, 
      n32447, n32448, n32449, n32450, n32452, n32456, n32457, n32460, n32462, 
      n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471, 
      n32472, n32474, n32477, n32478, n32479, n32480, n32481, n32482, n32483, 
      n32484, n32485, n32486, n32487, n32488, n32490, n32491, n32492, n32494, 
      n32495, n32497, n32498, n32499, n32504, n32505, n32506, n32507, n32508, 
      n32510, n32512, n32515, n32516, n32518, n32519, n32520, n32524, n32525, 
      n32526, n32527, n32528, n32531, n32532, n32534, n32535, n32536, n32537, 
      n32539, n32540, n32542, n32543, n32544, n32545, n32546, n32548, n32549, 
      n32551, n32552, n32555, n32556, n32557, n32558, n32559, n32562, n32563, 
      n32566, n32567, n32570, n32571, n32572, n32573, n32574, n32575, n32577, 
      n32579, n32580, n32581, n32583, n32584, n32585, n32586, n32588, n32590, 
      n32594, n32595, n32596, n32598, n32599, n32601, n32602, n32604, n32607, 
      n32608, n32609, n32610, n32613, n32614, n32615, n32616, n32617, n32618, 
      n32619, n32620, n32621, n32622, n32623, n32625, n32626, n32628, n32630, 
      n32631, n32633, n32634, n32636, n32637, n32638, n32639, n32640, n32641, 
      n32643, n32644, n32646, n32647, n32648, n32649, n32650, n32651, n32654, 
      n32657, n32658, n32660, n32661, n32662, n32663, n32664, n32666, n32667, 
      n32668, n32669, n32670, n32671, n32675, n32676, n32677, n32678, n32681, 
      n32682, n32683, n32684, n32685, n32686, n32689, n32690, n32691, n32693, 
      n32695, n32696, n32697, n32698, n32699, n32702, n32703, n32704, n32705, 
      n32706, n32708, n32712, n32714, n32718, n32719, n32720, n32721, n32722, 
      n32725, n32727, n32728, n32734, n32740, n32741, n32742, n32743, n32745, 
      n32746, n32747, n32748, n32750, n32752, n32753, n32755, n32756, n32757, 
      n32758, n32759, n32760, n32761, n32762, n32763, n32765, n32766, n32767, 
      n32768, n32769, n32771, n32773, n32775, n32776, n32777, n32778, n32779, 
      n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32789, n32790, 
      n32791, n32795, n32796, n32797, n32798, n32799, n32800, n32802, n32803, 
      n32805, n32806, n32807, n32808, n32811, n32813, n32814, n32815, n32817, 
      n32818, n32820, n32821, n32822, n32825, n32826, n32827, n32829, n32831, 
      n32832, n32833, n32836, n32837, n32838, n32839, n32842, n32843, n32844, 
      n32847, n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856, 
      n32857, n32858, n32860, n32861, n32863, n32865, n32866, n32867, n32868, 
      n32869, n32870, n32871, n32872, n32873, n32877, n32878, n32879, n32881, 
      n32882, n32883, n32884, n32885, n32886, n32889, n32890, n32891, n32892, 
      n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32902, n32903, 
      n32904, n32906, n32909, n32910, n32911, n32913, n32915, n32916, n32917, 
      n32918, n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931, 
      n32932, n32933, n32934, n32937, n32938, n32940, n32941, n32942, n32943, 
      n32944, n32945, n32946, n32948, n32950, n32951, n32952, n32953, n32954, 
      n32955, n32956, n32958, n32959, n32960, n32961, n32962, n32963, n32971, 
      n32972, n32973, n32974, n32976, n32977, n32979, n32980, n32981, n32983, 
      n32984, n32985, n32986, n32987, n32989, n32993, n32994, n32999, n33001, 
      n33002, n33004, n33005, n33006, n33007, n33008, n33010, n33011, n33012, 
      n33013, n33015, n33016, n33017, n33020, n33022, n33023, n33025, n33026, 
      n33027, n33028, n33029, n33030, n33032, n33034, n33036, n33037, n33038, 
      n33039, n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048, 
      n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057, 
      n33058, n33059, n33061, n33062, n33063, n33067, n33070, n33071, n33072, 
      n33073, n33074, n33075, n33077, n33080, n33081, n33082, n33083, n33085, 
      n33086, n33087, n33088, n33091, n33092, n33093, n33094, n33097, n33098, 
      n33100, n33101, n33102, n33104, n33106, n33107, n33108, n33109, n33111, 
      n33112, n33113, n33114, n33115, n33116, n33118, n33120, n33121, n33123, 
      n33125, n33128, n33129, n33130, n33131, n33132, n33133, n33135, n33138, 
      n33139, n33140, n33141, n33142, n33144, n33145, n33146, n33147, n33148, 
      n33151, n33152, n33153, n33154, n33155, n33156, n33158, n33160, n33161, 
      n33163, n33165, n33166, n33168, n33170, n33176, n33177, n33178, n33179, 
      n33180, n33182, n33183, n33184, n33185, n33186, n33187, n33188, n33190, 
      n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200, 
      n33201, n33202, n33203, n33204, n33206, n33207, n33208, n33209, n33215, 
      n33216, n33217, n33218, n33219, n33220, n33223, n33224, n33226, n33227, 
      n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33237, 
      n33239, n33240, n33242, n33243, n33244, n33246, n33247, n33248, n33249, 
      n33250, n33251, n33252, n33254, n33255, n33256, n33257, n33258, n33261, 
      n33262, n33263, n33264, n33266, n33267, n33268, n33270, n33271, n33272, 
      n33273, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283, 
      n33284, n33285, n33286, n33287, n33288, n33289, n33291, n33292, n33293, 
      n33295, n33296, n33297, n33299, n33300, n33301, n33302, n33303, n33304, 
      n33307, n33308, n33309, n33310, n33311, n33313, n33314, n33315, n33316, 
      n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325, 
      n33326, n33327, n33328, n33331, n33333, n33334, n33335, n33336, n33337, 
      n33340, n33344, n33346, n33347, n33348, n33349, n33350, n33352, n33353, 
      n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362, 
      n33363, n33364, n33365, n33366, n33368, n33369, n33370, n33371, n33372, 
      n33373, n33375, n33376, n33379, n33380, n33383, n33384, n33385, n33387, 
      n33388, n33389, n33392, n33393, n33394, n33395, n33396, n33398, n33399, 
      n33400, n33401, n33402, n33403, n33404, n33405, n33407, n33409, n33410, 
      n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420, 
      n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33431, 
      n33433, n33434, n33436, n33437, n33438, n33439, n33440, n33442, n33446, 
      n33449, n33450, n33452, n33453, n33455, n33456, n33457, n33459, n33460, 
      n33461, n33462, n33463, n33464, n33465, n33466, n33468, n33470, n33472, 
      n33473, n33474, n33476, n33478, n33479, n33480, n33481, n33482, n33483, 
      n33484, n33485, n33486, n33487, n33488, n33489, n33491, n33493, n33495, 
      n33496, n33498, n33500, n33503, n33504, n33505, n33506, n33509, n33510, 
      n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33519, n33520, 
      n33521, n33522, n33524, n33526, n33527, n33528, n33529, n33530, n33531, 
      n33532, n33533, n33534, n33535, n33538, n33539, n33541, n33544, n33546, 
      n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555, 
      n33557, n33558, n33559, n33561, n33563, n33565, n33566, n33567, n33568, 
      n33569, n33571, n33572, n33573, n33574, n33576, n33577, n33578, n33579, 
      n33580, n33581, n33582, n33584, n33585, n33586, n33587, n33591, n33593, 
      n33594, n33595, n33597, n33598, n33599, n33601, n33603, n33604, n33607, 
      n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33616, n33619, 
      n33620, n33621, n33622, n33623, n33625, n33628, n33629, n33630, n33631, 
      n33633, n33636, n33638, n33640, n33642, n33643, n33644, n33645, n33646, 
      n33647, n33648, n33649, n33650, n33651, n33653, n33655, n33656, n33659, 
      n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668, 
      n33669, n33671, n33672, n33674, n33675, n33676, n33677, n33678, n33679, 
      n33686, n33687, n33689, n33690, n33693, n33694, n33695, n33696, n33697, 
      n33698, n33700, n33701, n33702, n33703, n33705, n33706, n33707, n33708, 
      n33709, n33712, n33713, n33715, n33716, n33717, n33718, n33719, n33720, 
      n33721, n33722, n33724, n33725, n33726, n33727, n33730, n33731, n33733, 
      n33734, n33735, n33736, n33737, n33738, n33743, n33745, n33746, n33747, 
      n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756, 
      n33757, n33758, n33759, n33760, n33763, n33764, n33765, n33766, n33767, 
      n33771, n33773, n33775, n33776, n33777, n33780, n33781, n33782, n33784, 
      n33785, n33786, n33788, n33789, n33792, n33793, n33795, n33799, n33802, 
      n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811, 
      n33812, n33813, n33815, n33816, n33817, n33818, n33821, n33824, n33825, 
      n33826, n33829, n33831, n33832, n33833, n33834, n33837, n33839, n33840, 
      n33841, n33842, n33843, n33844, n33845, n33847, n33848, n33849, n33850, 
      n33851, n33852, n33853, n33855, n33856, n33858, n33859, n33860, n33861, 
      n33862, n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870, 
      n33871, n33876, n33879, n33883, n33885, n33886, n33887, n33888, n33890, 
      n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33899, n33902, 
      n33904, n33905, n33906, n33908, n33909, n33910, n33911, n33912, n33913, 
      n33916, n33919, n33921, n33924, n33925, n33926, n33928, n33929, n33931, 
      n33933, n33934, n33935, n33936, n33937, n33939, n33944, n33945, n33946, 
      n33947, n33948, n33949, n33950, n33952, n33954, n33955, n33956, n33957, 
      n33958, n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966, 
      n33967, n33968, n33969, n33972, n33973, n33976, n33978, n33979, n33980, 
      n33981, n33986, n33987, n33990, n33993, n33995, n33996, n33997, n33999, 
      n34000, n34001, n34003, n34004, n34005, n34006, n34007, n34008, n34009, 
      n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018, 
      n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34027, n34028, 
      n34030, n34031, n34032, n34033, n34034, n34036, n34037, n34038, n34039, 
      n34040, n34041, n34042, n34043, n34044, n34046, n34047, n34048, n34049, 
      n34050, n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059, 
      n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068, 
      n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076, n34077, 
      n34078, n34080, n34081, n34082, n34083, n34085, n34086, n34087, n34088, 
      n34089, n34090, n34091, n34092, n34094, n34096, n34097, n34099, n34103, 
      n34104, n34105, n34108, n34111, n34112, n34113, n34114, n34115, n34116, 
      n34117, n34120, n34121, n34122, n34123, n34124, n34126, n34128, n34129, 
      n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139, 
      n34141, n34142, n34143, n34144, n34145, n34147, n34148, n34149, n34150, 
      n34151, n34152, n34153, n34154, n34156, n34157, n34160, n34161, n34162, 
      n34163, n34165, n34166, n34167, n34170, n34171, n34172, n34173, n34175, 
      n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183, n34184, 
      n34185, n34186, n34188, n34189, n34190, n34192, n34193, n34194, n34195, 
      n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34205, 
      n34206, n34208, n34210, n34212, n34213, n34214, n34215, n34216, n34217, 
      n34218, n34220, n34221, n34223, n34224, n34225, n34226, n34227, n34228, 
      n34231, n34233, n34235, n34237, n34238, n34239, n34244, n34245, n34246, 
      n34247, n34249, n34250, n34251, n34252, n34254, n34256, n34257, n34259, 
      n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268, 
      n34269, n34270, n34272, n34274, n34275, n34276, n34277, n34279, n34282, 
      n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291, 
      n34292, n34296, n34297, n34298, n34299, n34301, n34303, n34305, n34306, 
      n34307, n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34317, 
      n34319, n34323, n34324, n34325, n34326, n34329, n34330, n34332, n34335, 
      n34336, n34337, n34339, n34340, n34342, n34343, n34344, n34345, n34347, 
      n34350, n34351, n34352, n34354, n34357, n34358, n34359, n34360, n34365, 
      n34366, n34368, n34370, n34371, n34372, n34373, n34374, n34375, n34377, 
      n34378, n34379, n34382, n34383, n34384, n34386, n34387, n34389, n34391, 
      n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34401, 
      n34402, n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411, 
      n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421, 
      n34422, n34424, n34426, n34427, n34428, n34430, n34433, n34435, n34436, 
      n34437, n34438, n34439, n34440, n34441, n34442, n34446, n34447, n34448, 
      n34450, n34451, n34452, n34453, n34454, n34457, n34458, n34459, n34460, 
      n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468, n34469, 
      n34470, n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479, 
      n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488, 
      n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497, 
      n34498, n34499, n34501, n34503, n34504, n34506, n34510, n34512, n34513, 
      n34514, n34515, n34516, n34518, n34519, n34520, n34521, n34522, n34524, 
      n34525, n34526, n34531, n34532, n34533, n34534, n34535, n34538, n34539, 
      n34540, n34541, n34544, n34545, n34546, n34547, n34549, n34552, n34553, 
      n34554, n34557, n34558, n34559, n34561, n34562, n34564, n34565, n34567, 
      n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576, 
      n34577, n34579, n34580, n34581, n34583, n34585, n34586, n34587, n34589, 
      n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599, n34601, 
      n34602, n34603, n34604, n34606, n34608, n34609, n34610, n34611, n34613, 
      n34615, n34616, n34618, n34619, n34620, n34621, n34622, n34627, n34630, 
      n34632, n34634, n34635, n34636, n34637, n34638, n34639, n34641, n34642, 
      n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651, 
      n34652, n34653, n34654, n34655, n34656, n34658, n34660, n34662, n34663, 
      n34664, n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673, 
      n34678, n34680, n34681, n34682, n34683, n34685, n34686, n34688, n34689, 
      n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697, n34698, 
      n34699, n34702, n34703, n34704, n34705, n34706, n34707, n34708, n34709, 
      n34711, n34712, n34713, n34715, n34716, n34717, n34718, n34719, n34720, 
      n34722, n34723, n34724, n34726, n34727, n34728, n34733, n34737, n34738, 
      n34739, n34740, n34742, n34743, n34745, n34746, n34747, n34750, n34751, 
      n34752, n34753, n34755, n34757, n34758, n34760, n34761, n34762, n34763, 
      n34764, n34766, n34767, n34768, n34769, n34770, n34772, n34773, n34774, 
      n34776, n34777, n34778, n34780, n34781, n34783, n34785, n34786, n34787, 
      n34788, n34789, n34790, n34793, n34794, n34795, n34796, n34799, n34800, 
      n34801, n34802, n34804, n34805, n34806, n34808, n34809, n34811, n34812, 
      n34813, n34814, n34815, n34817, n34819, n34820, n34821, n34822, n34823, 
      n34825, n34826, n34828, n34829, n34830, n34832, n34836, n34837, n34838, 
      n34840, n34841, n34842, n34843, n34844, n34846, n34847, n34848, n34849, 
      n34850, n34851, n34853, n34854, n34855, n34856, n34857, n34858, n34861, 
      n34863, n34866, n34867, n34868, n34869, n34870, n34871, n34876, n34877, 
      n34878, n34881, n34882, n34883, n34884, n34885, n34886, n34889, n34890, 
      n34891, n34892, n34893, n34894, n34895, n34897, n34898, n34899, n34900, 
      n34901, n34902, n34903, n34904, n34905, n34906, n34908, n34909, n34911, 
      n34912, n34913, n34914, n34915, n34918, n34920, n34922, n34923, n34924, 
      n34925, n34926, n34930, n34931, n34932, n34933, n34934, n34935, n34938, 
      n34939, n34940, n34942, n34943, n34944, n34945, n34947, n34948, n34949, 
      n34952, n34953, n34955, n34956, n34957, n34958, n34959, n34961, n34962, 
      n34963, n34964, n34965, n34966, n34967, n34969, n34972, n34973, n34974, 
      n34977, n34979, n34981, n34982, n34983, n34984, n34985, n34986, n34987, 
      n34989, n34990, n34993, n34995, n34996, n34997, n34998, n34999, n35000, 
      n35001, n35003, n35004, n35005, n35006, n35007, n35010, n35012, n35013, 
      n35014, n35015, n35016, n35017, n35018, n35019, n35021, n35022, n35023, 
      n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033, 
      n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35042, n35043, 
      n35045, n35046, n35047, n35048, n35049, n35051, n35053, n35054, n35055, 
      n35056, n35057, n35059, n35060, n35061, n35062, n35063, n35064, n35065, 
      n35067, n35068, n35070, n35071, n35072, n35073, n35075, n35076, n35077, 
      n35078, n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086, 
      n35087, n35088, n35089, n35092, n35093, n35095, n35096, n35097, n35098, 
      n35099, n35102, n35103, n35105, n35107, n35108, n35109, n35112, n35113, 
      n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122, 
      n35123, n35124, n35128, n35129, n35130, n35134, n35135, n35137, n35138, 
      n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147, 
      n35148, n35149, n35150, n35151, n35153, n35155, n35156, n35157, n35158, 
      n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35168, n35169, 
      n35170, n35171, n35172, n35173, n35175, n35176, n35177, n35178, n35179, 
      n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188, 
      n35189, n35190, n35191, n35192, n35193, n35194, n35196, n35197, n35198, 
      n35199, n35200, n35202, n35203, n35207, n35208, n35209, n35210, n35211, 
      n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220, 
      n35221, n35222, n35224, n35225, n35227, n35228, n35229, n35230, n35231, 
      n35232, n35233, n35234, n35235, n35237, n35238, n35239, n35240, n35241, 
      n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250, 
      n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259, 
      n35260, n35262, n35264, n35265, n35266, n35267, n35268, n35269, n35270, 
      n35271, n35272, n35273, n35274, n35278, n35279, n35280, n35281, n35282, 
      n35285, n35286, n35287, n35288, n35290, n35293, n35294, n35295, n35296, 
      n35297, n35299, n35300, n35301, n35302, n35303, n35309, n35310, n35311, 
      n35312, n35313, n35314, n35315, n35317, n35318, n35320, n35321, n35322, 
      n35323, n35324, n35326, n35327, n35329, n35330, n35331, n35332, n35333, 
      n35334, n35335, n35336, n35339, n35340, n35342, n35343, n35344, n35345, 
      n35347, n35348, n35349, n35350, n35351, n35353, n35355, n35357, n35359, 
      n35360, n35361, n35362, n35363, n35367, n35368, n35369, n35370, n35371, 
      n35373, n35374, n35376, n35377, n35379, n35380, n35381, n35384, n35386, 
      n35387, n35389, n35390, n35391, n35392, n35394, n35395, n35397, n35398, 
      n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35407, n35409, 
      n35410, n35414, n35415, n35417, n35419, n35420, n35421, n35422, n35423, 
      n35424, n35425, n35427, n35429, n35431, n35434, n35435, n35436, n35437, 
      n35438, n35439, n35440, n35441, n35442, n35443, n35445, n35446, n35447, 
      n35448, n35449, n35450, n35452, n35453, n35454, n35455, n35457, n35462, 
      n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471, 
      n35472, n35473, n35474, n35476, n35477, n35478, n35479, n35480, n35481, 
      n35483, n35485, n35487, n35489, n35490, n35491, n35492, n35494, n35495, 
      n35496, n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505, 
      n35506, n35507, n35508, n35510, n35511, n35513, n35514, n35517, n35519, 
      n35520, n35521, n35523, n35525, n35526, n35528, n35529, n35532, n35534, 
      n35535, n35536, n35537, n35541, n35542, n35543, n35544, n35545, n35547, 
      n35548, n35549, n35550, n35551, n35553, n35554, n35556, n35559, n35560, 
      n35561, n35563, n35564, n35566, n35567, n35568, n35569, n35570, n35571, 
      n35572, n35573, n35574, n35576, n35577, n35578, n35579, n35580, n35583, 
      n35584, n35585, n35586, n35588, n35590, n35591, n35594, n35595, n35596, 
      n35598, n35599, n35600, n35601, n35603, n35604, n35607, n35608, n35610, 
      n35611, n35612, n35613, n35614, n35616, n35617, n35618, n35619, n35621, 
      n35622, n35623, n35624, n35625, n35626, n35627, n35629, n35630, n35631, 
      n35632, n35633, n35636, n35637, n35639, n35640, n35642, n35644, n35645, 
      n35646, n35647, n35648, n35649, n35651, n35652, n35653, n35654, n35655, 
      n35656, n35657, n35658, n35659, n35660, n35663, n35664, n35665, n35666, 
      n35667, n35668, n35670, n35671, n35673, n35675, n35676, n35677, n35678, 
      n35679, n35681, n35684, n35685, n35686, n35687, n35688, n35689, n35690, 
      n35693, n35694, n35695, n35696, n35697, n35699, n35702, n35704, n35705, 
      n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35715, n35718, 
      n35720, n35721, n35722, n35723, n35724, n35726, n35727, n35728, n35729, 
      n35730, n35731, n35732, n35733, n35734, n35735, n35737, n35741, n35743, 
      n35744, n35745, n35746, n35747, n35748, n35749, n35750, n35752, n35753, 
      n35754, n35755, n35756, n35757, n35758, n35760, n35761, n35762, n35763, 
      n35764, n35765, n35766, n35767, n35768, n35769, n35771, n35772, n35774, 
      n35776, n35777, n35779, n35780, n35781, n35782, n35784, n35785, n35786, 
      n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795, 
      n35796, n35801, n35802, n35803, n35804, n35805, n35806, n35808, n35809, 
      n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35818, n35819, 
      n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828, 
      n35830, n35832, n35833, n35834, n35835, n35836, n35837, n35839, n35840, 
      n35841, n35842, n35843, n35844, n35846, n35847, n35848, n35849, n35851, 
      n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860, 
      n35862, n35863, n35864, n35867, n35868, n35869, n35870, n35871, n35872, 
      n35873, n35874, n35875, n35877, n35878, n35879, n35880, n35881, n35882, 
      n35883, n35885, n35886, n35887, n35888, n35889, n35890, n35891, n35892, 
      n35893, n35894, n35895, n35896, n35897, n35899, n35900, n35901, n35902, 
      n35903, n35904, n35905, n35906, n35908, n35909, n35910, n35911, n35912, 
      n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35923, 
      n35924, n35925, n35926, n35928, n35931, n35932, n35935, n35936, n35938, 
      n35939, n35941, n35942, n35943, n35944, n35947, n35948, n35950, n35952, 
      n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961, 
      n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970, 
      n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979, 
      n35981, n35983, n35984, n35985, n35986, n35987, n35988, n35990, n35992, 
      n35993, n35994, n35996, n35997, n35998, n35999, n36000, n36001, n36002, 
      n36003, n36004, n36005, n36006, n36007, n36008, n36011, n36013, n36016, 
      n36017, n36019, n36020, n36021, n36022, n36023, n36024, n36026, n36027, 
      n36029, n36030, n36031, n36032, n36034, n36035, n36036, n36038, n36039, 
      n36040, n36041, n36043, n36044, n36046, n36048, n36050, n36051, n36052, 
      n36053, n36055, n36057, n36058, n36059, n36060, n36062, n36063, n36064, 
      n36065, n36066, n36067, n36068, n36069, n36071, n36072, n36073, n36074, 
      n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083, 
      n36084, n36085, n36086, n36087, n36090, n36091, n36092, n36094, n36095, 
      n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104, 
      n36105, n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36117, 
      n36119, n36120, n36123, n36124, n36125, n36126, n36127, n36128, n36129, 
      n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138, 
      n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147, 
      n36150, n36151, n36152, n36154, n36157, n36159, n36160, n36162, n36163, 
      n36164, n36165, n36166, n36167, n36168, n36170, n36171, n36172, n36173, 
      n36175, n36176, n36177, n36180, n36181, n36182, n36183, n36184, n36185, 
      n36186, n36187, n36188, n36190, n36191, n36193, n36194, n36195, n36196, 
      n36197, n36199, n36200, n36201, n36203, n36204, n36205, n36206, n36207, 
      n36209, n36210, n36211, n36212, n36214, n36216, n36217, n36218, n36219, 
      n36222, n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230, 
      n36231, n36232, n36233, n36234, n36236, n36237, n36238, n36239, n36240, 
      n36241, n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250, 
      n36251, n36253, n36254, n36255, n36257, n36258, n36259, n36260, n36261, 
      n36262, n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270, 
      n36271, n36272, n36273, n36275, n36277, n36279, n36280, n36281, n36283, 
      n36284, n36286, n36287, n36289, n36290, n36291, n36292, n36293, n36295, 
      n36296, n36297, n36300, n36301, n36302, n36303, n36304, n36305, n36306, 
      n36307, n36308, n36309, n36310, n36311, n36313, n36314, n36317, n36320, 
      n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329, 
      n36333, n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36341, 
      n36342, n36343, n36344, n36345, n36346, n36348, n36349, n36351, n36352, 
      n36353, n36354, n36355, n36357, n36358, n36360, n36361, n36362, n36363, 
      n36364, n36365, n36366, n36368, n36369, n36371, n36372, n36373, n36374, 
      n36375, n36376, n36377, n36378, n36379, n36380, n36382, n36383, n36384, 
      n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393, 
      n36394, n36395, n36396, n36397, n36400, n36402, n36403, n36404, n36406, 
      n36407, n36408, n36410, n36411, n36412, n36413, n36414, n36415, n36416, 
      n36418, n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36428, 
      n36429, n36430, n36431, n36433, n36434, n36435, n36436, n36441, n36442, 
      n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451, 
      n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459, n36460, 
      n36461, n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470, 
      n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478, n36480, 
      n36481, n36483, n36485, n36486, n36487, n36488, n36490, n36491, n36492, 
      n36493, n36494, n36496, n36497, n36498, n36499, n36500, n36501, n36502, 
      n36506, n36507, n36508, n36509, n36510, n36511, n36513, n36514, n36515, 
      n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523, n36524, 
      n36525, n36526, n36527, n36528, n36529, n36530, n36532, n36535, n36537, 
      n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546, 
      n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556, 
      n36558, n36559, n36560, n36561, n36563, n36564, n36566, n36567, n36568, 
      n36569, n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578, 
      n36579, n36581, n36582, n36583, n36584, n36585, n36587, n36588, n36589, 
      n36590, n36591, n36592, n36593, n36594, n36595, n36596, n36598, n36601, 
      n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36611, 
      n36612, n36613, n36615, n36616, n36617, n36618, n36620, n36621, n36622, 
      n36623, n36624, n36626, n36627, n36628, n36629, n36630, n36631, n36632, 
      n36633, n36634, n36635, n36637, n36638, n36639, n36640, n36641, n36643, 
      n36644, n36645, n36646, n36647, n36649, n36651, n36654, n36655, n36656, 
      n36658, n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36668, 
      n36669, n36671, n36672, n36673, n36674, n36676, n36677, n36678, n36679, 
      n36680, n36682, n36683, n36685, n36686, n36687, n36689, n36690, n36691, 
      n36692, n36693, n36694, n36696, n36697, n36698, n36699, n36700, n36701, 
      n36702, n36703, n36705, n36706, n36707, n36708, n36709, n36711, n36712, 
      n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724, 
      n36725, n36726, n36727, n36728, n36729, n36730, n36731, n36734, n36735, 
      n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743, n36744, 
      n36745, n36746, n36748, n36750, n36751, n36752, n36753, n36754, n36755, 
      n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764, 
      n36765, n36766, n36767, n36769, n36772, n36773, n36774, n36775, n36776, 
      n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36785, n36786, 
      n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795, 
      n36796, n36797, n36798, n36799, n36800, n36801, n36803, n36804, n36805, 
      n36806, n36807, n36808, n36809, n36810, n36812, n36814, n36815, n36816, 
      n36817, n36818, n36819, n36821, n36822, n36824, n36827, n36828, n36829, 
      n36830, n36831, n36832, n36833, n36834, n36835, n36837, n36838, n36839, 
      n36840, n36842, n36843, n36844, n36846, n36847, n36848, n36849, n36850, 
      n36851, n36852, n36853, n36854, n36856, n36857, n36858, n36859, n36860, 
      n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869, 
      n36871, n36872, n36873, n36876, n36877, n36878, n36880, n36882, n36884, 
      n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892, n36893, 
      n36894, n36895, n36896, n36897, n36899, n36900, n36902, n36903, n36905, 
      n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914, 
      n36915, n36916, n36918, n36919, n36920, n36922, n36923, n36924, n36925, 
      n36926, n36927, n36928, n36929, n36930, n36931, n36932, n36935, n36936, 
      n36938, n36939, n36940, n36941, n36942, n36944, n36945, n36946, n36947, 
      n36949, n36951, n36952, n36953, n36954, n36955, n36957, n36958, n36959, 
      n36960, n36961, n36962, n36964, n36965, n36966, n36967, n36968, n36969, 
      n36970, n36971, n36972, n36974, n36976, n36977, n36979, n36980, n36981, 
      n36984, n36985, n36986, n36988, n36989, n36990, n36991, n36992, n36993, 
      n36994, n36995, n36996, n36997, n36998, n36999, n37001, n37002, n37003, 
      n37005, n37006, n37007, n37008, n37010, n37011, n37012, n37013, n37014, 
      n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37023, n37024, 
      n37025, n37026, n37027, n37028, n37030, n37031, n37032, n37033, n37034, 
      n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043, 
      n37044, n37045, n37047, n37048, n37049, n37050, n37051, n37052, n37053, 
      n37054, n37055, n37056, n37057, n37059, n37060, n37061, n37062, n37063, 
      n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072, 
      n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081, 
      n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37092, 
      n37093, n37094, n37095, n37096, n37097, n37098, n37099, n37100, n37101, 
      n37102, n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110, 
      n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119, 
      n37120, n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128, 
      n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137, 
      n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146, 
      n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155, 
      n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163, n37164, 
      n37165, n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173, 
      n37174, n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182, 
      n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191, 
      n37192, n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200, 
      n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209, 
      n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218, 
      n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227, 
      n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236, 
      n37237, n37238, n37239, n37240, n37241, n37242, n37243, n37244, n37245, 
      n37246, n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254, 
      n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263, 
      n37264, n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272, 
      n37273, n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281, 
      n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290, 
      n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299, 
      n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307, n37308, 
      n37309, n37310, n37311, n37312, n37313, n37314, n37315, n37316, n37317, 
      n37318, n37319, n37320, n37321, n37322, n37324, n37325, n37326, n37327, 
      n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336, 
      n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345, 
      n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354, 
      n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363, 
      n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372, 
      n37373, n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381, 
      n37382, n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390, 
      n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399, 
      n37400, n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408, 
      n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417, 
      n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426, 
      n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435, 
      n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444, 
      n37445, n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453, 
      n37454, n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462, 
      n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471, 
      n37472, n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480, 
      n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37489, n37490, 
      n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499, 
      n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508, 
      n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517, 
      n37518, n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526, 
      n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535, 
      n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544, 
      n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553, 
      n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562, 
      n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571, 
      n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580, 
      n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588, n37589, 
      n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598, 
      n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607, 
      n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616, 
      n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625, 
      n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634, 
      n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643, 
      n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652, 
      n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660, n37661, 
      n37662, n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670, 
      n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678, n37679, 
      n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688, 
      n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697, 
      n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706, 
      n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715, 
      n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724, 
      n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732, n37733, 
      n37734, n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742, 
      n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750, n37751, 
      n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760, 
      n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769, 
      n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778, 
      n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787, 
      n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796, 
      n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804, n37805, 
      n37806, n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814, 
      n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822, n37823, 
      n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832, 
      n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841, 
      n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850, 
      n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859, 
      n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867, n37868, 
      n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876, n37877, 
      n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886, 
      n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895, 
      n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904, 
      n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913, 
      n37914, n37915, n37916, n37918, n37919, n37920, n37921, n37922, n37923, 
      n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931, n37932, 
      n37933, n37934, n37935, n37936, n37937, n37938, n37939, n37940, n37941, 
      n37942, n37943, n37944, n37945, n37946, n37947, n37948, n37949, n37950, 
      n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958, n37959, 
      n37960, n37961, n37962, n37963, n37964, n37965, n37966, n37967, n37968, 
      n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977, 
      n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985, n37986, 
      n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994, n37995, 
      n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003, n38004, 
      n38005, n38006, n38007, n38008, n38009, n38010, n38011, n38012, n38013, 
      n38014, n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022, 
      n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030, n38031, 
      n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040, 
      n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049, 
      n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058, 
      n38059, n38060, n38061, n38062, n38063, n38064, n38065, n38066, n38067, 
      n38068, n38069, n38070, n38071, n38072, n38073, n38074, n38075, n38076, 
      n38077, n38078, n38079, n38080, n38081, n38082, n38083, n38084, n38085, 
      n38086, n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094, 
      n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102, n38103, 
      n38104, n38105, n38106, n38107, n38108, n38109, n38110, n38111, n38112, 
      n38113, n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121, 
      n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129, n38130, 
      n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138, n38139, 
      n38140, n38141, n38142, n38143, n38144, n38145, n38146, n38147, n38148, 
      n38149, n38150, n38151, n38152, n38153, n38154, n38155, n38156, n38157, 
      n38158, n38159, n38160, n38161, n38162, n38163, n38164, n38165, n38166, 
      n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174, n38175, 
      n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184, 
      n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193, 
      n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202, 
      n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210, n38211, 
      n38212, n38213, n38214, n38215, n38216, n38217, n38218, n38219, n38220, 
      n38221, n38222, n38223, n38224, n38225, n38226, n38227, n38228, n38229, 
      n38230, n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238, 
      n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246, n38247, 
      n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256, 
      n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265, 
      n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274, 
      n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282, n38283, 
      n38284, n38285, n38286, n38287, n38288, n38289, n38290, n38291, n38292, 
      n38293, n38294, n38295, n38296, n38297, n38298, n38299, n38300, n38301, 
      n38302, n38303, n38305, n38306, n38307, n38308, n38309, n38310, n38311, 
      n38312, n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320, 
      n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329, 
      n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338, 
      n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347, 
      n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355, n38356, 
      n38357, n38358, n38359, n38360, n38361, n38362, n38363, n38364, n38365, 
      n38366, n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374, 
      n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383, 
      n38384, n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392, 
      n38393, n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401, 
      n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410, 
      n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419, 
      n38420, n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428, 
      n38429, n38430, n38431, n38432, n38433, n38434, n38435, n38436, n38437, 
      n38438, n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446, 
      n38448, n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457, 
      n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466, 
      n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475, 
      n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484, 
      n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493, 
      n38494, n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502, 
      n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511, 
      n38512, n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520, 
      n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529, 
      n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538, 
      n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547, 
      n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556, 
      n38557, n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565, 
      n38566, n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574, 
      n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583, 
      n38584, n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592, 
      n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601, 
      n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610, 
      n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619, 
      n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628, 
      n38629, n38630, n38631, n38632, n38633, n38634, n38635, n38636, n38637, 
      n38638, n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646, 
      n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655, 
      n38656, n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664, 
      n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673, 
      n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682, 
      n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691, 
      n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699, n38700, 
      n38701, n38702, n38703, n38704, n38705, n38706, n38707, n38708, n38709, 
      n38710, n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718, 
      n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727, 
      n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736, 
      n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745, 
      n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754, 
      n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763, 
      n38764, n38765, n38766, n38767, n38768, n38769, n38770, n38771, n38772, 
      n38773, n38774, n38775, n38776, n38777, n38778, n38779, n38780, n38781, 
      n38782, n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790, 
      n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799, 
      n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808, 
      n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817, 
      n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826, 
      n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835, 
      n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843, n38844, 
      n38845, n38846, n38847, n38848, n38849, n38850, n38851, n38852, n38853, 
      n38854, n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862, 
      n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870, n38871, 
      n38872, n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880, 
      n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889, 
      n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898, 
      n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907, 
      n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915, n38916, 
      n38917, n38918, n38919, n38920, n38921, n38922, n38923, n38924, n38925, 
      n38926, n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934, 
      n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942, n38943, 
      n38944, n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952, 
      n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961, 
      n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970, 
      n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979, 
      n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987, n38988, 
      n38989, n38990, n38991, n38992, n38993, n38994, n38995, n38996, n38997, 
      n38998, n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006, 
      n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015, 
      n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024, 
      n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033, 
      n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042, 
      n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051, 
      n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059, n39060, 
      n39061, n39062, n39063, n39064, n39065, n39066, n39067, n39068, n39069, 
      n39070, n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078, 
      n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086, n39087, 
      n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096, 
      n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105, 
      n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114, 
      n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123, 
      n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131, n39132, 
      n39133, n39134, n39135, n39136, n39137, n39138, n39139, n39140, n39141, 
      n39142, n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150, 
      n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158, n39159, 
      n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168, 
      n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177, 
      n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186, 
      n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195, 
      n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203, n39204, 
      n39205, n39206, n39207, n39208, n39209, n39210, n39211, n39212, n39213, 
      n39214, n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222, 
      n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231, 
      n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240, 
      n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249, 
      n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258, 
      n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266, n39267, 
      n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275, n39276, 
      n39277, n39278, n39279, n39280, n39281, n39282, n39283, n39284, n39285, 
      n39286, n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294, 
      n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303, 
      n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312, 
      n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321, 
      n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330, 
      n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338, n39339, 
      n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347, n39348, 
      n39349, n39350, n39351, n39352, n39353, n39354, n39355, n39356, n39357, 
      n39358, n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366, 
      n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374, n39375, 
      n39376, n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384, 
      n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393, 
      n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402, 
      n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410, n39411, 
      n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419, n39420, 
      n39421, n39422, n39423, n39424, n39425, n39426, n39427, n39428, n39429, 
      n39430, n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438, 
      n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446, n39447, 
      n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456, 
      n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465, 
      n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474, 
      n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483, 
      n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491, n39492, 
      n39493, n39494, n39495, n39496, n39497, n39498, n39499, n39500, n39501, 
      n39502, n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510, 
      n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518, n39519, 
      n39520, n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528, 
      n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537, 
      n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546, 
      n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555, 
      n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563, n39564, 
      n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39572, n39573, 
      n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582, 
      n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590, n39591, 
      n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600, 
      n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609, 
      n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618, 
      n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627, 
      n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635, n39636, 
      n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644, n39645, 
      n39646, n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39654, 
      n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662, n39663, 
      n39664, n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672, 
      n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681, 
      n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690, 
      n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699, 
      n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708, 
      n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716, n39717, 
      n39718, n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726, 
      n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734, n39735, 
      n39736, n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744, 
      n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753, 
      n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762, 
      n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770, n39771, 
      n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779, n39780, 
      n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788, n39789, 
      n39790, n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798, 
      n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806, n39807, 
      n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816, 
      n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825, 
      n39826, n39827, n39828, n39829, n39830 : std_logic;

begin
   
   U42 : INV_X1 port map( I => n29438, ZN => n1383);
   U65 : NAND2_X1 port map( A1 => n17238, A2 => n30229, ZN => n18043);
   U73 : NOR2_X1 port map( A1 => n29491, A2 => n37099, ZN => n28649);
   U108 : INV_X1 port map( I => n32304, ZN => n30187);
   U115 : AND2_X1 port map( A1 => n15153, A2 => n9393, Z => n15605);
   U117 : NOR2_X1 port map( A1 => n30232, A2 => n29263, ZN => n19310);
   U150 : INV_X1 port map( I => n19910, ZN => n29614);
   U153 : INV_X1 port map( I => n29045, ZN => n5741);
   U157 : INV_X1 port map( I => n19833, ZN => n20329);
   U231 : NOR2_X1 port map( A1 => n9686, A2 => n14278, ZN => n450);
   U234 : AOI21_X1 port map( A1 => n36814, A2 => n39664, B => n37460, ZN => 
                           n15110);
   U268 : INV_X2 port map( I => n28689, ZN => n17771);
   U293 : NAND2_X1 port map( A1 => n11283, A2 => n7690, ZN => n76);
   U361 : INV_X1 port map( I => n27671, ZN => n14828);
   U375 : INV_X1 port map( I => n30101, ZN => n1703);
   U376 : INV_X1 port map( I => n19774, ZN => n29854);
   U377 : INV_X1 port map( I => n19947, ZN => n17275);
   U378 : INV_X1 port map( I => n29538, ZN => n1698);
   U384 : INV_X1 port map( I => n29838, ZN => n1702);
   U385 : INV_X1 port map( I => n19751, ZN => n21226);
   U403 : INV_X1 port map( I => n19877, ZN => n27465);
   U419 : NAND2_X1 port map( A1 => n27455, A2 => n5101, ZN => n19030);
   U449 : INV_X1 port map( I => n27108, ZN => n27230);
   U459 : INV_X1 port map( I => n37075, ZN => n943);
   U471 : NAND2_X1 port map( A1 => n1079, A2 => n995, ZN => n1797);
   U487 : NOR2_X1 port map( A1 => n998, A2 => n27508, ZN => n27421);
   U518 : INV_X1 port map( I => n26784, ZN => n3);
   U527 : OAI22_X1 port map( A1 => n36873, A2 => n925, B1 => n9147, B2 => 
                           n17034, ZN => n7006);
   U533 : NAND3_X1 port map( A1 => n2292, A2 => n33858, A3 => n8651, ZN => 
                           n27125);
   U538 : NOR3_X1 port map( A1 => n32168, A2 => n13181, A3 => n38483, ZN => 
                           n17573);
   U540 : NAND2_X1 port map( A1 => n9654, A2 => n925, ZN => n81);
   U546 : OAI22_X1 port map( A1 => n17823, A2 => n32797, B1 => n26284, B2 => 
                           n1229, ZN => n5221);
   U552 : INV_X1 port map( I => n19615, ZN => n20021);
   U560 : OR2_X1 port map( A1 => n14455, A2 => n26876, Z => n13184);
   U629 : INV_X1 port map( I => n28968, ZN => n15046);
   U633 : INV_X1 port map( I => n26587, ZN => n12383);
   U641 : INV_X1 port map( I => n28910, ZN => n1730);
   U642 : INV_X1 port map( I => n19952, ZN => n19799);
   U643 : INV_X1 port map( I => n19887, ZN => n16498);
   U644 : INV_X1 port map( I => n29671, ZN => n19432);
   U781 : AOI21_X1 port map( A1 => n6300, A2 => n34010, B => n18837, ZN => 
                           n13533);
   U783 : AOI21_X1 port map( A1 => n1535, A2 => n2581, B => n25466, ZN => n1933
                           );
   U794 : INV_X1 port map( I => n579, ZN => n25443);
   U822 : AOI21_X1 port map( A1 => n25681, A2 => n7705, B => n24536, ZN => n242
                           );
   U827 : NOR3_X1 port map( A1 => n18810, A2 => n14436, A3 => n1543, ZN => 
                           n5710);
   U830 : NAND2_X1 port map( A1 => n20052, A2 => n31809, ZN => n25554);
   U852 : NAND2_X1 port map( A1 => n36105, A2 => n34427, ZN => n25519);
   U892 : INV_X1 port map( I => n19729, ZN => n1733);
   U893 : INV_X1 port map( I => n29319, ZN => n14969);
   U900 : INV_X1 port map( I => n19851, ZN => n1719);
   U903 : INV_X1 port map( I => n29707, ZN => n21280);
   U904 : INV_X1 port map( I => n19885, ZN => n1735);
   U905 : INV_X1 port map( I => n29801, ZN => n20781);
   U906 : INV_X1 port map( I => n19913, ZN => n18993);
   U912 : INV_X1 port map( I => n29298, ZN => n17646);
   U913 : INV_X1 port map( I => n30207, ZN => n20804);
   U922 : INV_X1 port map( I => n19649, ZN => n20748);
   U925 : OR2_X1 port map( A1 => n25184, A2 => n7967, Z => n817);
   U933 : NAND2_X1 port map( A1 => n39817, A2 => n18845, ZN => n24754);
   U938 : NAND2_X1 port map( A1 => n35560, A2 => n1580, ZN => n24490);
   U939 : NAND3_X1 port map( A1 => n9921, A2 => n24685, A3 => n24686, ZN => 
                           n7969);
   U985 : INV_X1 port map( I => n24795, ZN => n7177);
   U1004 : NAND2_X1 port map( A1 => n24734, A2 => n5390, ZN => n5389);
   U1020 : INV_X1 port map( I => n18983, ZN => n24614);
   U1041 : INV_X1 port map( I => n37227, ZN => n24275);
   U1052 : NOR2_X1 port map( A1 => n14686, A2 => n37994, ZN => n12);
   U1117 : NAND2_X1 port map( A1 => n15892, A2 => n9383, ZN => n3398);
   U1143 : INV_X1 port map( I => n23846, ZN => n20594);
   U1168 : NAND2_X1 port map( A1 => n1861, A2 => n1632, ZN => n530);
   U1171 : OR2_X1 port map( A1 => n23567, A2 => n1643, Z => n788);
   U1181 : INV_X1 port map( I => n23484, ZN => n23364);
   U1189 : INV_X1 port map( I => n38704, ZN => n98);
   U1218 : INV_X1 port map( I => n7644, ZN => n16729);
   U1284 : NAND2_X1 port map( A1 => n18415, A2 => n22859, ZN => n5110);
   U1288 : INV_X1 port map( I => n19440, ZN => n14188);
   U1294 : NOR2_X1 port map( A1 => n19698, A2 => n23103, ZN => n23105);
   U1304 : INV_X1 port map( I => n36453, ZN => n19769);
   U1309 : OAI21_X1 port map( A1 => n22860, A2 => n22861, B => n22859, ZN => 
                           n4760);
   U1311 : NOR2_X1 port map( A1 => n23032, A2 => n22958, ZN => n22954);
   U1331 : INV_X1 port map( I => n407, ZN => n8809);
   U1341 : INV_X1 port map( I => n19167, ZN => n22875);
   U1351 : INV_X1 port map( I => n22879, ZN => n5892);
   U1362 : INV_X1 port map( I => n11778, ZN => n22900);
   U1369 : BUF_X2 port map( I => n17628, Z => n906);
   U1388 : NAND2_X1 port map( A1 => n9546, A2 => n64, ZN => n9521);
   U1390 : INV_X1 port map( I => n6014, ZN => n1808);
   U1409 : NAND2_X1 port map( A1 => n35193, A2 => n4497, ZN => n367);
   U1453 : INV_X2 port map( I => n16760, ZN => n22310);
   U1470 : AOI21_X1 port map( A1 => n21524, A2 => n21478, B => n533, ZN => n532
                           );
   U1484 : OR2_X1 port map( A1 => n21688, A2 => n21339, Z => n5047);
   U1490 : NOR2_X1 port map( A1 => n19470, A2 => n13472, ZN => n3943);
   U1499 : INV_X1 port map( I => n21750, ZN => n21029);
   U1504 : NOR2_X1 port map( A1 => n19545, A2 => n7536, ZN => n10918);
   U1508 : NAND2_X1 port map( A1 => n37200, A2 => n18576, ZN => n18699);
   U1529 : INV_X1 port map( I => n17964, ZN => n15338);
   U1532 : AND2_X1 port map( A1 => n21722, A2 => n20685, Z => n12738);
   U1541 : INV_X1 port map( I => n688, ZN => n1348);
   U1571 : INV_X2 port map( I => n1897, ZN => n4734);
   U1572 : INV_X2 port map( I => n10004, ZN => n14635);
   U1587 : OAI22_X2 port map( A1 => n6542, A2 => n24576, B1 => n958, B2 => 
                           n24723, ZN => n6541);
   U1608 : OAI21_X2 port map( A1 => n4636, A2 => n17353, B => n5355, ZN => 
                           n25567);
   U1611 : INV_X2 port map( I => n28054, ZN => n6788);
   U1638 : INV_X4 port map( I => n27235, ZN => n945);
   U1640 : AND2_X1 port map( A1 => n27314, A2 => n33417, Z => n18436);
   U1646 : INV_X4 port map( I => n26839, ZN => n1092);
   U1682 : NAND2_X2 port map( A1 => n10140, A2 => n26107, ZN => n10139);
   U1722 : OAI21_X2 port map( A1 => n5022, A2 => n7431, B => n27215, ZN => 
                           n28350);
   U1761 : INV_X2 port map( I => n6657, ZN => n21042);
   U1792 : AOI21_X2 port map( A1 => n14541, A2 => n18143, B => n17866, ZN => 
                           n17865);
   U1827 : OAI21_X2 port map( A1 => n22230, A2 => n17156, B => n36237, ZN => 
                           n17155);
   U1830 : INV_X4 port map( I => n22160, ZN => n1333);
   U1831 : AOI21_X2 port map( A1 => n24599, A2 => n24597, B => n1563, ZN => 
                           n7443);
   U1846 : BUF_X2 port map( I => n37043, Z => n4714);
   U1860 : INV_X2 port map( I => n30464, ZN => n11846);
   U1871 : INV_X2 port map( I => n29574, ZN => n1393);
   U1873 : BUF_X4 port map( I => n17696, Z => n603);
   U1876 : OAI21_X2 port map( A1 => n26003, A2 => n603, B => n26005, ZN => 
                           n9667);
   U1883 : INV_X4 port map( I => n17712, ZN => n1236);
   U1884 : NOR2_X2 port map( A1 => n37106, A2 => n259, ZN => n9217);
   U1912 : AOI21_X2 port map( A1 => n15585, A2 => n24695, B => n38777, ZN => 
                           n12504);
   U1913 : NOR2_X1 port map( A1 => n13036, A2 => n17824, ZN => n207);
   U1922 : AOI21_X2 port map( A1 => n21836, A2 => n21837, B => n14911, ZN => 
                           n14910);
   U1927 : INV_X2 port map( I => n882, ZN => n1202);
   U1942 : AOI21_X2 port map( A1 => n16353, A2 => n20102, B => n37021, ZN => 
                           n8446);
   U1966 : OAI21_X2 port map( A1 => n7972, A2 => n7966, B => n3655, ZN => n3654
                           );
   U1967 : AOI21_X2 port map( A1 => n25388, A2 => n25389, B => n25582, ZN => 
                           n4827);
   U1973 : INV_X2 port map( I => n30465, ZN => n1545);
   U2044 : INV_X2 port map( I => n27253, ZN => n27115);
   U2057 : INV_X2 port map( I => n20858, ZN => n17712);
   U2066 : OAI21_X2 port map( A1 => n37151, A2 => n26005, B => n26004, ZN => 
                           n20050);
   U2079 : INV_X2 port map( I => n19223, ZN => n25677);
   U2093 : OAI21_X2 port map( A1 => n39446, A2 => n23095, B => n8594, ZN => 
                           n14305);
   U2111 : OAI21_X2 port map( A1 => n15737, A2 => n35224, B => n1424, ZN => 
                           n8008);
   U2132 : NAND2_X2 port map( A1 => n23391, A2 => n37093, ZN => n15642);
   U2152 : INV_X2 port map( I => n7364, ZN => n15385);
   U2194 : INV_X4 port map( I => n13758, ZN => n1494);
   U2222 : NAND2_X1 port map( A1 => n31527, A2 => n17469, ZN => n4768);
   U2228 : NOR2_X1 port map( A1 => n15768, A2 => n37096, ZN => n29358);
   U2274 : NAND2_X2 port map( A1 => n6257, A2 => n17348, ZN => n17347);
   U2291 : NOR3_X1 port map( A1 => n23110, A2 => n20782, A3 => n12392, ZN => 
                           n16132);
   U2295 : AND2_X1 port map( A1 => n9725, A2 => n22920, Z => n22858);
   U2304 : INV_X1 port map( I => n9516, ZN => n7904);
   U2307 : INV_X1 port map( I => n22571, ZN => n629);
   U2352 : NOR2_X1 port map( A1 => n33966, A2 => n5579, ZN => n633);
   U2357 : INV_X2 port map( I => n24247, ZN => n1130);
   U2393 : INV_X1 port map( I => n28940, ZN => n110);
   U2403 : INV_X2 port map( I => n8519, ZN => n8518);
   U2423 : INV_X1 port map( I => n28204, ZN => n1208);
   U2424 : NAND2_X1 port map( A1 => n8583, A2 => n29924, ZN => n8582);
   U2426 : OR2_X2 port map( A1 => n13425, A2 => n26177, Z => n26655);
   U2428 : NOR2_X1 port map( A1 => n5089, A2 => n27284, ZN => n4716);
   U2442 : AND2_X2 port map( A1 => n21567, A2 => n3294, Z => n3821);
   U2455 : AOI21_X1 port map( A1 => n11067, A2 => n13981, B => n37096, ZN => 
                           n13273);
   U2469 : OAI21_X2 port map( A1 => n11773, A2 => n14774, B => n11771, ZN => 
                           n2546);
   U2483 : INV_X2 port map( I => n853, ZN => n19712);
   U2504 : INV_X2 port map( I => n33966, ZN => n2347);
   U2515 : AND2_X1 port map( A1 => n27910, A2 => n33845, Z => n15372);
   U2519 : XOR2_X1 port map( A1 => n9205, A2 => n22382, Z => n2781);
   U2522 : NAND2_X2 port map( A1 => n2607, A2 => n2610, ZN => n9701);
   U2544 : OAI21_X2 port map( A1 => n37124, A2 => n7590, B => n21094, ZN => n10
                           );
   U2545 : INV_X2 port map( I => n11, ZN => n6163);
   U2559 : AOI22_X2 port map( A1 => n22193, A2 => n22194, B1 => n22191, B2 => 
                           n22192, ZN => n9982);
   U2560 : INV_X2 port map( I => n25307, ZN => n18837);
   U2587 : NAND3_X1 port map( A1 => n21063, A2 => n21062, A3 => n13352, ZN => 
                           n21061);
   U2597 : INV_X2 port map( I => n22904, ZN => n4862);
   U2613 : OAI21_X2 port map( A1 => n28190, A2 => n28191, B => n7310, ZN => 
                           n14030);
   U2641 : NAND2_X2 port map( A1 => n8053, A2 => n8052, ZN => n23609);
   U2643 : NOR2_X2 port map( A1 => n1821, A2 => n29078, ZN => n16839);
   U2646 : NOR2_X2 port map( A1 => n20112, A2 => n27315, ZN => n20111);
   U2660 : XOR2_X1 port map( A1 => n507, A2 => n30324, Z => n2446);
   U2688 : AOI21_X2 port map( A1 => n37069, A2 => n25512, B => n36486, ZN => 
                           n46);
   U2727 : NAND2_X2 port map( A1 => n13624, A2 => n13636, ZN => n15332);
   U2730 : INV_X2 port map( I => n63, ZN => n21285);
   U2788 : INV_X1 port map( I => n9616, ZN => n19089);
   U2802 : OR2_X1 port map( A1 => n24902, A2 => n20158, Z => n812);
   U2812 : INV_X1 port map( I => n20207, ZN => n24146);
   U2815 : NAND2_X2 port map( A1 => n27967, A2 => n27966, ZN => n28559);
   U2821 : NAND2_X1 port map( A1 => n170, A2 => n4095, ZN => n29991);
   U2828 : NOR3_X2 port map( A1 => n29448, A2 => n19791, A3 => n29447, ZN => 
                           n85);
   U2831 : OAI21_X2 port map( A1 => n19579, A2 => n3821, B => n3295, ZN => 
                           n3327);
   U2869 : AOI21_X2 port map( A1 => n5972, A2 => n5973, B => n5971, ZN => n5579
                           );
   U2877 : XOR2_X1 port map( A1 => n15671, A2 => n2352, Z => n2351);
   U2893 : NAND2_X2 port map( A1 => n12030, A2 => n22161, ZN => n22162);
   U2897 : NAND2_X2 port map( A1 => n2413, A2 => n109, ZN => n13217);
   U2900 : XOR2_X1 port map( A1 => n110, A2 => n5755, Z => n5889);
   U2918 : XOR2_X1 port map( A1 => n22639, A2 => n6329, Z => n8313);
   U2940 : NAND2_X2 port map( A1 => n19963, A2 => n25587, ZN => n6448);
   U2941 : INV_X2 port map( I => n118, ZN => n759);
   U2942 : XOR2_X1 port map( A1 => n5096, A2 => n12919, Z => n118);
   U2971 : XOR2_X1 port map( A1 => n5031, A2 => n19910, Z => n11881);
   U2994 : XOR2_X1 port map( A1 => n22640, A2 => n22551, Z => n12102);
   U3023 : OAI21_X2 port map( A1 => n6043, A2 => n8800, B => n1194, ZN => n137)
                           ;
   U3044 : XOR2_X1 port map( A1 => n15336, A2 => n39073, Z => n16270);
   U3058 : XOR2_X1 port map( A1 => n8015, A2 => n8016, Z => n16271);
   U3094 : XOR2_X1 port map( A1 => n1458, A2 => n27776, Z => n27675);
   U3099 : OR2_X1 port map( A1 => n25772, A2 => n25939, Z => n155);
   U3105 : AOI21_X2 port map( A1 => n2405, A2 => n21924, B => n8076, ZN => 
                           n2404);
   U3107 : INV_X2 port map( I => n157, ZN => n8000);
   U3115 : XOR2_X1 port map( A1 => n158, A2 => n2592, Z => n11335);
   U3116 : XOR2_X1 port map( A1 => n159, A2 => n31605, Z => n158);
   U3119 : NAND2_X2 port map( A1 => n6263, A2 => n17094, ZN => n8249);
   U3140 : INV_X2 port map( I => n170, ZN => n775);
   U3150 : XOR2_X1 port map( A1 => n27831, A2 => n20796, Z => n18663);
   U3152 : AOI21_X2 port map( A1 => n20209, A2 => n16074, B => n14151, ZN => 
                           n14150);
   U3153 : NAND2_X2 port map( A1 => n171, A2 => n24498, ZN => n25266);
   U3163 : XOR2_X1 port map( A1 => n22757, A2 => n15753, Z => n3530);
   U3201 : OR2_X1 port map( A1 => n26116, A2 => n30302, Z => n187);
   U3211 : NAND4_X2 port map( A1 => n26426, A2 => n26425, A3 => n26427, A4 => 
                           n26674, ZN => n19135);
   U3213 : XOR2_X1 port map( A1 => n18512, A2 => n190, Z => n27671);
   U3214 : XOR2_X1 port map( A1 => n18510, A2 => n18511, Z => n190);
   U3224 : XOR2_X1 port map( A1 => n30322, A2 => n12437, Z => n13235);
   U3225 : NOR2_X2 port map( A1 => n11275, A2 => n4619, ZN => n22465);
   U3228 : INV_X2 port map( I => n37678, ZN => n21410);
   U3253 : NAND3_X2 port map( A1 => n10774, A2 => n17961, A3 => n24757, ZN => 
                           n25197);
   U3260 : CLKBUF_X2 port map( I => Key(63), Z => n19953);
   U3261 : BUF_X2 port map( I => Key(74), Z => n30150);
   U3266 : NAND2_X1 port map( A1 => n16692, A2 => n34073, ZN => n19013);
   U3269 : INV_X2 port map( I => n25203, ZN => n3655);
   U3288 : AOI21_X1 port map( A1 => n263, A2 => n10152, B => n1603, ZN => n7813
                           );
   U3294 : AOI21_X2 port map( A1 => n37201, A2 => n20981, B => n19569, ZN => 
                           n17829);
   U3295 : XOR2_X1 port map( A1 => n35463, A2 => n26573, Z => n5447);
   U3308 : NOR2_X2 port map( A1 => n207, A2 => n5221, ZN => n27385);
   U3323 : OR2_X1 port map( A1 => n11375, A2 => n28286, Z => n6714);
   U3330 : NOR2_X2 port map( A1 => n13111, A2 => n13110, ZN => n26996);
   U3331 : INV_X2 port map( I => n20613, ZN => n13110);
   U3334 : NAND2_X1 port map( A1 => n33703, A2 => n23399, ZN => n214);
   U3371 : NOR2_X1 port map( A1 => n230, A2 => n10050, ZN => n10190);
   U3372 : NOR2_X1 port map( A1 => n3415, A2 => n32209, ZN => n230);
   U3379 : XOR2_X1 port map( A1 => n33736, A2 => n9981, Z => n13001);
   U3382 : INV_X2 port map( I => n15337, ZN => n21571);
   U3390 : XNOR2_X1 port map( A1 => n23670, A2 => n19890, ZN => n540);
   U3398 : NAND2_X2 port map( A1 => n23826, A2 => n23825, ZN => n25040);
   U3399 : INV_X4 port map( I => n19718, ZN => n20376);
   U3401 : NAND2_X2 port map( A1 => n2276, A2 => n237, ZN => n22239);
   U3423 : AND2_X1 port map( A1 => n37157, A2 => n19085, Z => n5825);
   U3425 : OAI21_X1 port map( A1 => n18298, A2 => n25681, B => n242, ZN => 
                           n19503);
   U3443 : NOR2_X1 port map( A1 => n251, A2 => n30845, ZN => n11957);
   U3452 : XOR2_X1 port map( A1 => n19472, A2 => n26158, Z => n254);
   U3457 : XOR2_X1 port map( A1 => n15912, A2 => n16498, Z => n648);
   U3481 : XOR2_X1 port map( A1 => n27794, A2 => n1214, Z => n27497);
   U3498 : XOR2_X1 port map( A1 => n266, A2 => n17737, Z => n29450);
   U3503 : OR2_X1 port map( A1 => n13637, A2 => n13638, Z => n13019);
   U3514 : XNOR2_X1 port map( A1 => n16359, A2 => n16358, ZN => n523);
   U3522 : NAND3_X2 port map( A1 => n23818, A2 => n24184, A3 => n39703, ZN => 
                           n13782);
   U3532 : XOR2_X1 port map( A1 => n27737, A2 => n20479, Z => n27483);
   U3545 : OAI21_X2 port map( A1 => n27391, A2 => n14881, B => n37246, ZN => 
                           n26869);
   U3552 : OAI22_X1 port map( A1 => n11939, A2 => n15601, B1 => n280, B2 => 
                           n3462, ZN => n5811);
   U3555 : OAI21_X2 port map( A1 => n24700, A2 => n6791, B => n6490, ZN => 
                           n8388);
   U3568 : XOR2_X1 port map( A1 => n22703, A2 => n4493, Z => n22571);
   U3570 : NAND2_X2 port map( A1 => n15787, A2 => n23560, ZN => n23340);
   U3574 : AOI22_X2 port map( A1 => n11517, A2 => n14377, B1 => n26759, B2 => 
                           n6891, ZN => n11516);
   U3581 : XOR2_X1 port map( A1 => n17342, A2 => n1162, Z => n5692);
   U3590 : INV_X2 port map( I => n18829, ZN => n30109);
   U3606 : NAND2_X2 port map( A1 => n6898, A2 => n13252, ZN => n5218);
   U3613 : INV_X1 port map( I => n26818, ZN => n26990);
   U3648 : BUF_X2 port map( I => n12961, Z => n301);
   U3653 : XOR2_X1 port map( A1 => n476, A2 => n36065, Z => n23793);
   U3660 : BUF_X2 port map( I => n28673, Z => n306);
   U3661 : XOR2_X1 port map( A1 => n35654, A2 => n26532, Z => n6879);
   U3663 : NAND2_X1 port map( A1 => n12150, A2 => n12547, ZN => n307);
   U3666 : INV_X2 port map( I => n26919, ZN => n3606);
   U3674 : INV_X4 port map( I => n14379, ZN => n24390);
   U3715 : XOR2_X1 port map( A1 => n320, A2 => n9563, Z => n15159);
   U3747 : NAND2_X2 port map( A1 => n24646, A2 => n36321, ZN => n24599);
   U3758 : XOR2_X1 port map( A1 => n23723, A2 => n9153, Z => n6516);
   U3762 : XOR2_X1 port map( A1 => n331, A2 => n9003, Z => n14290);
   U3776 : OR2_X1 port map( A1 => n31518, A2 => n27424, Z => n336);
   U3807 : XOR2_X1 port map( A1 => n7022, A2 => n342, Z => n19888);
   U3813 : AND2_X1 port map( A1 => n21023, A2 => n344, Z => n8761);
   U3816 : NAND2_X2 port map( A1 => n346, A2 => n24485, ZN => n24874);
   U3826 : AOI21_X2 port map( A1 => n37165, A2 => n11243, B => n11241, ZN => 
                           n26124);
   U3838 : NOR2_X2 port map( A1 => n5098, A2 => n4516, ZN => n4515);
   U3853 : XOR2_X1 port map( A1 => n353, A2 => n6223, Z => n5656);
   U3856 : XOR2_X1 port map( A1 => n6033, A2 => n19355, Z => n27194);
   U3857 : OAI21_X2 port map( A1 => n37, A2 => n7872, B => n28215, ZN => n3928)
                           ;
   U3880 : NAND2_X2 port map( A1 => n21231, A2 => n24735, ZN => n24620);
   U3882 : XOR2_X1 port map( A1 => n2615, A2 => n6436, Z => n13207);
   U3884 : AOI22_X2 port map( A1 => n9461, A2 => n37837, B1 => n15298, B2 => 
                           n36819, ZN => n26163);
   U3945 : INV_X2 port map( I => n27798, ZN => n379);
   U3958 : NAND2_X2 port map( A1 => n1289, A2 => n1596, ZN => n23983);
   U3961 : INV_X2 port map( I => n29923, ZN => n29924);
   U3966 : INV_X4 port map( I => n11120, ZN => n12543);
   U3974 : AOI21_X2 port map( A1 => n21362, A2 => n21361, B => n21360, ZN => 
                           n19718);
   U3981 : NOR2_X2 port map( A1 => n21847, A2 => n21672, ZN => n20469);
   U3985 : INV_X2 port map( I => n23083, ZN => n23188);
   U3991 : XOR2_X1 port map( A1 => n387, A2 => n18416, Z => n9176);
   U4002 : XOR2_X1 port map( A1 => n15656, A2 => n15660, Z => n391);
   U4010 : NAND3_X2 port map( A1 => n25707, A2 => n25706, A3 => n25705, ZN => 
                           n26602);
   U4011 : OR2_X1 port map( A1 => n20776, A2 => n32471, Z => n12642);
   U4012 : NAND2_X2 port map( A1 => n24353, A2 => n24477, ZN => n1898);
   U4023 : NAND2_X1 port map( A1 => n36552, A2 => n8193, ZN => n4761);
   U4025 : INV_X2 port map( I => n9942, ZN => n21902);
   U4029 : BUF_X2 port map( I => n7757, Z => n6445);
   U4033 : INV_X4 port map( I => n17307, ZN => n22265);
   U4039 : NAND2_X2 port map( A1 => n13986, A2 => n2792, ZN => n13606);
   U4041 : OAI21_X1 port map( A1 => n20474, A2 => n29704, B => n29581, ZN => 
                           n20473);
   U4044 : OAI21_X1 port map( A1 => n28699, A2 => n16295, B => n28696, ZN => 
                           n10303);
   U4052 : XOR2_X1 port map( A1 => n2317, A2 => n16133, Z => n10026);
   U4054 : BUF_X2 port map( I => Key(109), Z => n19825);
   U4060 : XOR2_X1 port map( A1 => n27724, A2 => n27640, Z => n27798);
   U4070 : INV_X2 port map( I => n22665, ZN => n1324);
   U4079 : NAND2_X2 port map( A1 => n13293, A2 => n13292, ZN => n13289);
   U4093 : NOR2_X2 port map( A1 => n21416, A2 => n21415, ZN => n21982);
   U4100 : XOR2_X1 port map( A1 => n412, A2 => n851, Z => n3486);
   U4106 : XOR2_X1 port map( A1 => n416, A2 => n17642, Z => n20702);
   U4107 : XOR2_X1 port map( A1 => n29148, A2 => n14221, Z => n416);
   U4123 : NAND2_X1 port map( A1 => n16158, A2 => n34783, ZN => n422);
   U4127 : AND2_X1 port map( A1 => n7536, A2 => n21410, Z => n10915);
   U4138 : XOR2_X1 port map( A1 => n2473, A2 => n427, Z => n3027);
   U4139 : XOR2_X1 port map( A1 => n2471, A2 => n22654, Z => n427);
   U4147 : XOR2_X1 port map( A1 => n431, A2 => n33965, Z => n15854);
   U4156 : AOI21_X1 port map( A1 => n29918, A2 => n29919, B => n434, ZN => 
                           n16992);
   U4194 : INV_X1 port map( I => n10144, ZN => n440);
   U4197 : XOR2_X1 port map( A1 => n29085, A2 => n28826, Z => n4141);
   U4213 : XOR2_X1 port map( A1 => n16523, A2 => n5370, Z => n3709);
   U4220 : INV_X2 port map( I => n18959, ZN => n21730);
   U4225 : AOI21_X2 port map( A1 => n16578, A2 => n12793, B => n5147, ZN => 
                           n5146);
   U4230 : AOI22_X1 port map( A1 => n9907, A2 => n13108, B1 => n13106, B2 => 
                           n29222, ZN => n13105);
   U4235 : NAND2_X2 port map( A1 => n3867, A2 => n3864, ZN => n3863);
   U4239 : NAND2_X2 port map( A1 => n22300, A2 => n35431, ZN => n9941);
   U4254 : OAI21_X2 port map( A1 => n9723, A2 => n9722, B => n1608, ZN => 
                           n13073);
   U4278 : XOR2_X1 port map( A1 => n17756, A2 => n29974, Z => n3478);
   U4280 : AOI21_X2 port map( A1 => n30364, A2 => n8757, B => n462, ZN => n7150
                           );
   U4289 : XOR2_X1 port map( A1 => n14986, A2 => n27533, Z => n18060);
   U4294 : INV_X1 port map( I => n1740, ZN => n29163);
   U4306 : INV_X2 port map( I => n26729, ZN => n8814);
   U4320 : NOR2_X1 port map( A1 => n37160, A2 => n25630, ZN => n17855);
   U4328 : INV_X2 port map( I => n474, ZN => n12365);
   U4334 : NAND2_X2 port map( A1 => n2341, A2 => n17101, ZN => n15136);
   U4343 : NAND3_X2 port map( A1 => n4660, A2 => n15966, A3 => n5552, ZN => 
                           n4875);
   U4351 : INV_X4 port map( I => n19594, ZN => n1316);
   U4363 : XOR2_X1 port map( A1 => n485, A2 => n6802, Z => n6801);
   U4364 : XOR2_X1 port map( A1 => n4796, A2 => n11688, Z => n485);
   U4371 : INV_X2 port map( I => n8454, ZN => n12081);
   U4376 : NAND3_X2 port map( A1 => n22095, A2 => n22097, A3 => n22096, ZN => 
                           n22648);
   U4385 : INV_X4 port map( I => n22337, ZN => n22100);
   U4389 : INV_X2 port map( I => n22092, ZN => n22356);
   U4397 : XOR2_X1 port map( A1 => n31127, A2 => n29131, Z => n489);
   U4404 : OR2_X1 port map( A1 => n2257, A2 => n22019, Z => n2709);
   U4412 : NOR2_X2 port map( A1 => n19609, A2 => n19641, ZN => n21433);
   U4413 : XOR2_X1 port map( A1 => n2997, A2 => n27493, Z => n8425);
   U4441 : INV_X4 port map( I => n18144, ZN => n1200);
   U4445 : INV_X4 port map( I => n20476, ZN => n1354);
   U4456 : NAND2_X2 port map( A1 => n8971, A2 => n10044, ZN => n18059);
   U4457 : AOI21_X2 port map( A1 => n18059, A2 => n21371, B => n9253, ZN => 
                           n9251);
   U4477 : NAND2_X2 port map( A1 => n16642, A2 => n16643, ZN => n19847);
   U4482 : XOR2_X1 port map( A1 => n10653, A2 => n10622, Z => n6212);
   U4487 : XOR2_X1 port map( A1 => n18597, A2 => n509, Z => n784);
   U4492 : XOR2_X1 port map( A1 => n26482, A2 => n9398, Z => n3459);
   U4494 : INV_X1 port map( I => n26483, ZN => n2711);
   U4511 : XOR2_X1 port map( A1 => n514, A2 => n22057, Z => n9420);
   U4519 : NAND2_X2 port map( A1 => n25830, A2 => n1512, ZN => n25919);
   U4521 : OAI21_X1 port map( A1 => n11718, A2 => n902, B => n515, ZN => n11719
                           );
   U4525 : AND2_X1 port map( A1 => n10171, A2 => n2722, Z => n12213);
   U4528 : XOR2_X1 port map( A1 => n11355, A2 => n33936, Z => n11354);
   U4540 : OR3_X1 port map( A1 => n15354, A2 => n114, A3 => n1816, Z => n1766);
   U4553 : INV_X2 port map( I => n3526, ZN => n20405);
   U4558 : INV_X4 port map( I => n4553, ZN => n25978);
   U4570 : XOR2_X1 port map( A1 => n28999, A2 => n28998, Z => n18452);
   U4574 : XOR2_X1 port map( A1 => n525, A2 => n30479, Z => n1455);
   U4575 : XOR2_X1 port map( A1 => n16218, A2 => n11996, Z => n525);
   U4583 : INV_X2 port map( I => n11643, ZN => n19293);
   U4592 : NAND2_X2 port map( A1 => n34404, A2 => n9524, ZN => n9523);
   U4609 : INV_X2 port map( I => n855, ZN => n17515);
   U4618 : AOI22_X2 port map( A1 => n9705, A2 => n18112, B1 => n9886, B2 => 
                           n39650, ZN => n7759);
   U4623 : INV_X2 port map( I => n19978, ZN => n25623);
   U4638 : AOI21_X2 port map( A1 => n538, A2 => n21764, B => n15148, ZN => 
                           n15614);
   U4640 : AOI21_X2 port map( A1 => n14899, A2 => n33580, B => n14898, ZN => 
                           n14897);
   U4644 : XOR2_X1 port map( A1 => n540, A2 => n23684, Z => n16893);
   U4653 : XOR2_X1 port map( A1 => n10200, A2 => n1867, Z => n12410);
   U4660 : NAND2_X2 port map( A1 => n4597, A2 => n11434, ZN => n5044);
   U4677 : XOR2_X1 port map( A1 => n7944, A2 => n7148, Z => n19112);
   U4678 : NAND2_X2 port map( A1 => n7144, A2 => n7145, ZN => n7148);
   U4684 : AOI22_X2 port map( A1 => n919, A2 => n21833, B1 => n21834, B2 => 
                           n19620, ZN => n15951);
   U4686 : NOR2_X1 port map( A1 => n19349, A2 => n7905, ZN => n551);
   U4695 : AOI21_X2 port map( A1 => n18104, A2 => n38215, B => n29956, ZN => 
                           n19093);
   U4713 : INV_X2 port map( I => n39823, ZN => n11707);
   U4717 : NOR2_X2 port map( A1 => n13964, A2 => n13963, ZN => n13962);
   U4729 : XOR2_X1 port map( A1 => n562, A2 => n18301, Z => n16905);
   U4746 : OAI21_X2 port map( A1 => n24147, A2 => n5360, B => n5359, ZN => 
                           n24794);
   U4780 : INV_X2 port map( I => n21792, ZN => n21660);
   U4786 : INV_X2 port map( I => n21432, ZN => n21822);
   U4810 : XOR2_X1 port map( A1 => n588, A2 => n29983, Z => Ciphertext(137));
   U4811 : OAI22_X1 port map( A1 => n29982, A2 => n29981, B1 => n18200, B2 => 
                           n5678, ZN => n588);
   U4812 : AND2_X1 port map( A1 => n17867, A2 => n7883, Z => n2058);
   U4828 : AOI21_X2 port map( A1 => n13409, A2 => n10536, B => n19969, ZN => 
                           n28656);
   U4835 : NAND2_X2 port map( A1 => n5479, A2 => n5477, ZN => n12685);
   U4838 : NAND2_X2 port map( A1 => n13669, A2 => n13671, ZN => n13442);
   U4850 : INV_X2 port map( I => n38210, ZN => n25472);
   U4859 : NOR2_X1 port map( A1 => n35604, A2 => n15245, ZN => n15243);
   U4870 : INV_X2 port map( I => n9626, ZN => n22652);
   U4880 : NOR2_X2 port map( A1 => n9050, A2 => n23032, ZN => n22956);
   U4882 : XOR2_X1 port map( A1 => n17277, A2 => n18434, Z => n7327);
   U4883 : NAND2_X2 port map( A1 => n28272, A2 => n13609, ZN => n12644);
   U4884 : INV_X2 port map( I => n12644, ZN => n20663);
   U4888 : XOR2_X1 port map( A1 => n25124, A2 => n25125, Z => n606);
   U4890 : XOR2_X1 port map( A1 => n608, A2 => n16861, Z => n27538);
   U4916 : XOR2_X1 port map( A1 => n6635, A2 => n2979, Z => n2215);
   U4930 : INV_X2 port map( I => n615, ZN => n10896);
   U4931 : XOR2_X1 port map( A1 => n10899, A2 => n10897, Z => n615);
   U4934 : AOI21_X1 port map( A1 => n29480, A2 => n29466, B => n616, ZN => 
                           n29467);
   U4938 : AOI21_X1 port map( A1 => n619, A2 => n29753, B => n30555, ZN => 
                           n29725);
   U4939 : NAND2_X1 port map( A1 => n38143, A2 => n29740, ZN => n619);
   U4941 : NAND2_X2 port map( A1 => n27386, A2 => n7680, ZN => n27492);
   U4942 : NAND2_X2 port map( A1 => n21057, A2 => n21060, ZN => n21961);
   U4943 : XOR2_X1 port map( A1 => n23882, A2 => n23724, Z => n5412);
   U4947 : NOR2_X1 port map( A1 => n6202, A2 => n1183, ZN => n6201);
   U4965 : NOR2_X1 port map( A1 => n4613, A2 => n20391, ZN => n15719);
   U4973 : BUF_X4 port map( I => n4381, Z => n2625);
   U4978 : AOI21_X2 port map( A1 => n14118, A2 => n28129, B => n14117, ZN => 
                           n13690);
   U4980 : NAND2_X2 port map( A1 => n4978, A2 => n4977, ZN => n28207);
   U4983 : INV_X4 port map( I => n38204, ZN => n11700);
   U4985 : XOR2_X1 port map( A1 => n3203, A2 => n629, Z => n628);
   U4987 : INV_X4 port map( I => n13285, ZN => n1351);
   U4995 : XOR2_X1 port map( A1 => n18305, A2 => n13639, Z => n632);
   U4999 : XOR2_X1 port map( A1 => n2943, A2 => n8940, Z => n29148);
   U5001 : XOR2_X1 port map( A1 => n14977, A2 => n5873, Z => n635);
   U5003 : XOR2_X1 port map( A1 => n636, A2 => n18976, Z => n18269);
   U5005 : INV_X1 port map( I => n36735, ZN => n8970);
   U5011 : NOR3_X1 port map( A1 => n21693, A2 => n21410, A3 => n36735, ZN => 
                           n9040);
   U5012 : NAND2_X1 port map( A1 => n21814, A2 => n21352, ZN => n21431);
   U5013 : AOI21_X1 port map( A1 => n10822, A2 => n36735, B => n21693, ZN => 
                           n10821);
   U5017 : INV_X1 port map( I => n8026, ZN => n22590);
   U5044 : INV_X1 port map( I => n19775, ZN => n26330);
   U5049 : INV_X1 port map( I => n19929, ZN => n1727);
   U5056 : INV_X1 port map( I => n11562, ZN => n923);
   U5062 : NOR3_X1 port map( A1 => n36344, A2 => n19728, A3 => n38591, ZN => 
                           n27123);
   U5065 : INV_X1 port map( I => n19903, ZN => n1704);
   U5066 : NAND2_X1 port map( A1 => n27421, A2 => n30768, ZN => n27509);
   U5067 : INV_X1 port map( I => n19845, ZN => n19020);
   U5079 : INV_X1 port map( I => n29875, ZN => n28868);
   U5086 : INV_X1 port map( I => n19875, ZN => n29109);
   U5088 : INV_X1 port map( I => n29432, ZN => n15181);
   U5090 : INV_X1 port map( I => n29003, ZN => n1365);
   U5091 : INV_X1 port map( I => n19817, ZN => n29730);
   U5092 : INV_X1 port map( I => n19905, ZN => n15273);
   U5094 : INV_X1 port map( I => n19904, ZN => n15700);
   U5095 : INV_X1 port map( I => n19755, ZN => n1738);
   U5096 : AND2_X1 port map( A1 => n22188, A2 => n39607, Z => n637);
   U5097 : XNOR2_X1 port map( A1 => n23680, A2 => n30006, ZN => n638);
   U5098 : XNOR2_X1 port map( A1 => n22613, A2 => n15762, ZN => n639);
   U5105 : XNOR2_X1 port map( A1 => n29680, A2 => n1010, ZN => n646);
   U5108 : XNOR2_X1 port map( A1 => n4302, A2 => n27739, ZN => n650);
   U5111 : XNOR2_X1 port map( A1 => n35610, A2 => n21280, ZN => n654);
   U5112 : XNOR2_X1 port map( A1 => n18300, A2 => n17428, ZN => n655);
   U5113 : XNOR2_X1 port map( A1 => n17605, A2 => n37110, ZN => n656);
   U5114 : XNOR2_X1 port map( A1 => n25271, A2 => n19937, ZN => n657);
   U5115 : XNOR2_X1 port map( A1 => n22510, A2 => n20206, ZN => n658);
   U5118 : XNOR2_X1 port map( A1 => n24065, A2 => n29671, ZN => n661);
   U5119 : XNOR2_X1 port map( A1 => n16492, A2 => n28831, ZN => n662);
   U5120 : XNOR2_X1 port map( A1 => n30612, A2 => n31771, ZN => n663);
   U5121 : XNOR2_X1 port map( A1 => n25175, A2 => n19950, ZN => n664);
   U5122 : XNOR2_X1 port map( A1 => n35262, A2 => n29229, ZN => n665);
   U5124 : XNOR2_X1 port map( A1 => n23874, A2 => n23591, ZN => n666);
   U5126 : XNOR2_X1 port map( A1 => n36867, A2 => n22763, ZN => n669);
   U5129 : XNOR2_X1 port map( A1 => n24050, A2 => n19758, ZN => n672);
   U5130 : XNOR2_X1 port map( A1 => n27595, A2 => n19676, ZN => n673);
   U5131 : XNOR2_X1 port map( A1 => n34902, A2 => n15046, ZN => n674);
   U5132 : XNOR2_X1 port map( A1 => n23884, A2 => n29964, ZN => n675);
   U5134 : XNOR2_X1 port map( A1 => n27799, A2 => n1161, ZN => n677);
   U5135 : XNOR2_X1 port map( A1 => n23894, A2 => n1367, ZN => n678);
   U5137 : XNOR2_X1 port map( A1 => n29041, A2 => n19913, ZN => n680);
   U5138 : XNOR2_X1 port map( A1 => n29095, A2 => n1377, ZN => n681);
   U5139 : XNOR2_X1 port map( A1 => n27617, A2 => n30114, ZN => n682);
   U5142 : XOR2_X1 port map( A1 => Plaintext(10), A2 => Key(10), Z => n686);
   U5144 : INV_X2 port map( I => n22219, ZN => n1688);
   U5145 : XOR2_X1 port map( A1 => Plaintext(22), A2 => Key(22), Z => n688);
   U5148 : XNOR2_X1 port map( A1 => Plaintext(30), A2 => Key(30), ZN => n690);
   U5151 : XOR2_X1 port map( A1 => Plaintext(114), A2 => Key(114), Z => n694);
   U5152 : INV_X1 port map( I => n21805, ZN => n21693);
   U5153 : XNOR2_X1 port map( A1 => n22651, A2 => n22430, ZN => n696);
   U5154 : XNOR2_X1 port map( A1 => n22463, A2 => n16648, ZN => n697);
   U5155 : XNOR2_X1 port map( A1 => n4493, A2 => n19648, ZN => n698);
   U5156 : XNOR2_X1 port map( A1 => n22474, A2 => n32993, ZN => n699);
   U5157 : XNOR2_X1 port map( A1 => n32135, A2 => n19885, ZN => n700);
   U5158 : XNOR2_X1 port map( A1 => n10268, A2 => n10267, ZN => n701);
   U5160 : XNOR2_X1 port map( A1 => n20392, A2 => n29363, ZN => n704);
   U5161 : XNOR2_X1 port map( A1 => n22731, A2 => n19254, ZN => n705);
   U5162 : XNOR2_X1 port map( A1 => n22775, A2 => n29689, ZN => n706);
   U5163 : AND2_X1 port map( A1 => n21461, A2 => n21870, Z => n707);
   U5164 : XOR2_X1 port map( A1 => n17285, A2 => n17283, Z => n708);
   U5166 : XNOR2_X1 port map( A1 => n5185, A2 => n29320, ZN => n710);
   U5167 : XNOR2_X1 port map( A1 => n14322, A2 => n9496, ZN => n711);
   U5170 : XNOR2_X1 port map( A1 => n33672, A2 => n30253, ZN => n713);
   U5171 : XNOR2_X1 port map( A1 => n19932, A2 => n37957, ZN => n714);
   U5176 : XNOR2_X1 port map( A1 => n2145, A2 => n23658, ZN => n718);
   U5177 : XNOR2_X1 port map( A1 => n14385, A2 => n19876, ZN => n719);
   U5178 : XNOR2_X1 port map( A1 => n36218, A2 => n29411, ZN => n720);
   U5179 : XNOR2_X1 port map( A1 => n25301, A2 => n16618, ZN => n721);
   U5181 : XNOR2_X1 port map( A1 => n24932, A2 => n25160, ZN => n723);
   U5182 : XNOR2_X1 port map( A1 => n25216, A2 => n25123, ZN => n724);
   U5185 : XNOR2_X1 port map( A1 => n9701, A2 => n25296, ZN => n727);
   U5187 : XNOR2_X1 port map( A1 => n25030, A2 => n28934, ZN => n729);
   U5189 : XNOR2_X1 port map( A1 => n25241, A2 => n29649, ZN => n731);
   U5194 : XNOR2_X1 port map( A1 => n10012, A2 => n1733, ZN => n736);
   U5195 : XNOR2_X1 port map( A1 => n26262, A2 => n19761, ZN => n737);
   U5196 : XNOR2_X1 port map( A1 => n26455, A2 => n19677, ZN => n738);
   U5197 : XNOR2_X1 port map( A1 => n26340, A2 => n26357, ZN => n739);
   U5199 : XNOR2_X1 port map( A1 => n24933, A2 => n25177, ZN => n741);
   U5200 : XNOR2_X1 port map( A1 => n23970, A2 => n23697, ZN => n742);
   U5201 : XNOR2_X1 port map( A1 => n9246, A2 => n965, ZN => n743);
   U5203 : XNOR2_X1 port map( A1 => n5084, A2 => n29223, ZN => n745);
   U5205 : XNOR2_X1 port map( A1 => n26255, A2 => n1050, ZN => n747);
   U5206 : XNOR2_X1 port map( A1 => n6989, A2 => n29514, ZN => n748);
   U5207 : XNOR2_X1 port map( A1 => n6989, A2 => n29831, ZN => n749);
   U5208 : XNOR2_X1 port map( A1 => n26587, A2 => n19805, ZN => n750);
   U5211 : INV_X1 port map( I => n19226, ZN => n26895);
   U5215 : XNOR2_X1 port map( A1 => n27664, A2 => n19936, ZN => n756);
   U5219 : XNOR2_X1 port map( A1 => n35188, A2 => n30090, ZN => n760);
   U5220 : XNOR2_X1 port map( A1 => n31620, A2 => n35140, ZN => n761);
   U5221 : XNOR2_X1 port map( A1 => n27528, A2 => n19355, ZN => n763);
   U5222 : XNOR2_X1 port map( A1 => n28966, A2 => n30150, ZN => n764);
   U5223 : XNOR2_X1 port map( A1 => n28940, A2 => n1369, ZN => n765);
   U5226 : XNOR2_X1 port map( A1 => n13852, A2 => n19786, ZN => n769);
   U5227 : XNOR2_X1 port map( A1 => n10343, A2 => n29067, ZN => n770);
   U5229 : XNOR2_X1 port map( A1 => n31535, A2 => n19887, ZN => n772);
   U5230 : XNOR2_X1 port map( A1 => n35832, A2 => n1733, ZN => n774);
   U5233 : XNOR2_X1 port map( A1 => n6311, A2 => n22469, ZN => n778);
   U5238 : XOR2_X1 port map( A1 => n6610, A2 => n6608, Z => n782);
   U5253 : XNOR2_X1 port map( A1 => n23623, A2 => n29974, ZN => n790);
   U5257 : XNOR2_X1 port map( A1 => n23927, A2 => n20594, ZN => n794);
   U5267 : XOR2_X1 port map( A1 => n15730, A2 => n15728, Z => n801);
   U5269 : BUF_X2 port map( I => n24285, Z => n13970);
   U5271 : INV_X2 port map( I => n24307, ZN => n14371);
   U5282 : NAND2_X2 port map( A1 => n24300, A2 => n39815, ZN => n14206);
   U5283 : AND2_X1 port map( A1 => n24191, A2 => n18466, Z => n808);
   U5291 : XNOR2_X1 port map( A1 => n25241, A2 => n19677, ZN => n810);
   U5295 : XOR2_X1 port map( A1 => n39765, A2 => n30122, Z => n814);
   U5301 : NAND2_X2 port map( A1 => n12914, A2 => n4840, ZN => n6759);
   U5305 : XNOR2_X1 port map( A1 => n824, A2 => n741, ZN => n823);
   U5307 : XOR2_X1 port map( A1 => n4551, A2 => n4550, Z => n825);
   U5313 : XOR2_X1 port map( A1 => n3187, A2 => n3188, Z => n830);
   U5320 : AND2_X2 port map( A1 => n25714, A2 => n25713, Z => n834);
   U5326 : XOR2_X1 port map( A1 => n19384, A2 => n29282, Z => n837);
   U5334 : XNOR2_X1 port map( A1 => n26359, A2 => n30068, ZN => n838);
   U5335 : XNOR2_X1 port map( A1 => n25595, A2 => n25594, ZN => n839);
   U5342 : XNOR2_X1 port map( A1 => n26191, A2 => n26192, ZN => n845);
   U5345 : XNOR2_X1 port map( A1 => n26488, A2 => n8950, ZN => n848);
   U5354 : XNOR2_X1 port map( A1 => n14770, A2 => n14771, ZN => n856);
   U5359 : XNOR2_X1 port map( A1 => n9300, A2 => n9297, ZN => n859);
   U5364 : AND2_X1 port map( A1 => n26934, A2 => n17993, Z => n863);
   U5371 : XOR2_X1 port map( A1 => n26410, A2 => n3858, Z => n866);
   U5373 : INV_X1 port map( I => n867, ZN => n9690);
   U5385 : XNOR2_X1 port map( A1 => n35189, A2 => n27823, ZN => n869);
   U5386 : XNOR2_X1 port map( A1 => n27491, A2 => n900, ZN => n870);
   U5389 : XNOR2_X1 port map( A1 => n27513, A2 => n27514, ZN => n873);
   U5396 : XNOR2_X1 port map( A1 => n20140, A2 => n19421, ZN => n877);
   U5399 : INV_X1 port map( I => n20531, ZN => n28222);
   U5408 : XNOR2_X1 port map( A1 => n9139, A2 => n7764, ZN => n886);
   U5421 : BUF_X2 port map( I => n28883, Z => n29486);
   U5422 : BUF_X2 port map( I => n30243, Z => n6443);
   U5425 : XNOR2_X1 port map( A1 => n28574, A2 => n28493, ZN => n893);
   U5430 : AOI21_X2 port map( A1 => n16144, A2 => n7612, B => n14764, ZN => 
                           n3923);
   U5434 : OAI21_X2 port map( A1 => n9319, A2 => n9318, B => n9317, ZN => 
                           n22219);
   U5443 : NAND2_X1 port map( A1 => n5402, A2 => n6285, ZN => n28017);
   U5446 : OAI21_X2 port map( A1 => n4375, A2 => n28215, B => n3928, ZN => 
                           n28326);
   U5456 : AOI21_X2 port map( A1 => n1319, A2 => n1654, B => n5437, ZN => 
                           n22851);
   U5460 : NAND2_X1 port map( A1 => n918, A2 => n21478, ZN => n14527);
   U5461 : NAND2_X1 port map( A1 => n20266, A2 => n21478, ZN => n2278);
   U5462 : NAND2_X1 port map( A1 => n21478, A2 => n37200, ZN => n1814);
   U5469 : OAI21_X2 port map( A1 => n22927, A2 => n8141, B => n37087, ZN => 
                           n23611);
   U5505 : INV_X2 port map( I => n16382, ZN => n26780);
   U5507 : NOR2_X1 port map( A1 => n23057, A2 => n3310, ZN => n8142);
   U5508 : NAND2_X1 port map( A1 => n18450, A2 => n11576, ZN => n21450);
   U5509 : OAI21_X2 port map( A1 => n2237, A2 => n2236, B => n2233, ZN => n2082
                           );
   U5519 : BUF_X4 port map( I => n22813, Z => n23078);
   U5537 : AOI22_X2 port map( A1 => n3268, A2 => n22301, B1 => n22039, B2 => 
                           n22299, ZN => n3267);
   U5549 : OAI22_X2 port map( A1 => n7911, A2 => n9546, B1 => n3181, B2 => 
                           n22147, ZN => n1965);
   U5557 : NOR2_X1 port map( A1 => n7240, A2 => n1921, ZN => n8359);
   U5565 : OAI21_X1 port map( A1 => n9231, A2 => n30038, B => n30009, ZN => 
                           n5369);
   U5577 : NOR3_X1 port map( A1 => n12081, A2 => n30187, A3 => n30240, ZN => 
                           n6864);
   U5600 : BUF_X4 port map( I => n27908, Z => n28755);
   U5609 : INV_X4 port map( I => n876, ZN => n18392);
   U5612 : NAND3_X1 port map( A1 => n28054, A2 => n34008, A3 => n1072, ZN => 
                           n13697);
   U5618 : INV_X1 port map( I => n33958, ZN => n18451);
   U5640 : NAND3_X1 port map( A1 => n26976, A2 => n12065, A3 => n10902, ZN => 
                           n26977);
   U5653 : INV_X1 port map( I => n924, ZN => n13801);
   U5665 : INV_X1 port map( I => n26165, ZN => n1096);
   U5669 : NAND3_X1 port map( A1 => n37683, A2 => n25992, A3 => n1012, ZN => 
                           n8161);
   U5670 : INV_X2 port map( I => n33440, ZN => n1101);
   U5672 : INV_X2 port map( I => n7901, ZN => n14375);
   U5684 : INV_X4 port map( I => n11060, ZN => n17353);
   U5699 : NOR2_X1 port map( A1 => n24500, A2 => n933, ZN => n12207);
   U5725 : INV_X2 port map( I => n10659, ZN => n19682);
   U5749 : OAI21_X2 port map( A1 => n22959, A2 => n22960, B => n7639, ZN => 
                           n5357);
   U5755 : NOR2_X1 port map( A1 => n7960, A2 => n8151, ZN => n23057);
   U5766 : INV_X2 port map( I => n18433, ZN => n23053);
   U5779 : NOR3_X1 port map( A1 => n22038, A2 => n8899, A3 => n21802, ZN => 
                           n5698);
   U5804 : NAND2_X2 port map( A1 => n16014, A2 => n16015, ZN => n22122);
   U5817 : BUF_X2 port map( I => n33506, Z => n19470);
   U5839 : NOR3_X1 port map( A1 => n971, A2 => n16510, A3 => n21285, ZN => 
                           n9048);
   U5841 : NAND3_X1 port map( A1 => n3986, A2 => n4095, A3 => n1058, ZN => 
                           n11217);
   U5852 : INV_X1 port map( I => n9930, ZN => n12765);
   U5858 : NAND2_X2 port map( A1 => n28350, A2 => n28351, ZN => n28496);
   U5874 : NOR2_X1 port map( A1 => n1473, A2 => n35500, ZN => n4254);
   U5906 : INV_X1 port map( I => n17097, ZN => n26686);
   U5910 : INV_X2 port map( I => n18390, ZN => n26688);
   U5913 : INV_X2 port map( I => n14121, ZN => n924);
   U5939 : INV_X1 port map( I => n252, ZN => n14460);
   U5950 : OAI22_X1 port map( A1 => n24603, A2 => n1270, B1 => n32391, B2 => 
                           n5282, ZN => n20807);
   U5961 : NAND2_X2 port map( A1 => n10777, A2 => n10784, ZN => n20039);
   U5962 : INV_X4 port map( I => n13779, ZN => n933);
   U5963 : AND2_X1 port map( A1 => n1597, A2 => n1586, Z => n10069);
   U5966 : NOR2_X1 port map( A1 => n7364, A2 => n5986, ZN => n24335);
   U5981 : INV_X1 port map( I => n23582, ZN => n14855);
   U5988 : NAND2_X1 port map( A1 => n7584, A2 => n37815, ZN => n7071);
   U6007 : NAND3_X1 port map( A1 => n11091, A2 => n39075, A3 => n5497, ZN => 
                           n5496);
   U6009 : NAND2_X1 port map( A1 => n22325, A2 => n12365, ZN => n17781);
   U6011 : NAND3_X1 port map( A1 => n37113, A2 => n18253, A3 => n17976, ZN => 
                           n1864);
   U6012 : INV_X1 port map( I => n9485, ZN => n9483);
   U6018 : NOR2_X1 port map( A1 => n17440, A2 => n22047, ZN => n22111);
   U6026 : INV_X1 port map( I => n19017, ZN => n22496);
   U6031 : NAND3_X1 port map( A1 => n6420, A2 => n1690, A3 => n21762, ZN => 
                           n6419);
   U6034 : NOR2_X1 port map( A1 => n18784, A2 => n21881, ZN => n9669);
   U6039 : OAI21_X1 port map( A1 => n21551, A2 => n21762, B => n21308, ZN => 
                           n6672);
   U6040 : INV_X1 port map( I => n21765, ZN => n1690);
   U6049 : INV_X2 port map( I => n16496, ZN => n21668);
   U6050 : INV_X1 port map( I => n21641, ZN => n21908);
   U6051 : CLKBUF_X2 port map( I => Key(18), Z => n19677);
   U6052 : CLKBUF_X2 port map( I => Key(28), Z => n19732);
   U6056 : CLKBUF_X2 port map( I => Key(172), Z => n29689);
   U6060 : AOI22_X1 port map( A1 => n29340, A2 => n29339, B1 => n12848, B2 => 
                           n20481, ZN => n12847);
   U6071 : INV_X4 port map( I => n12726, ZN => n939);
   U6095 : INV_X1 port map( I => n30243, ZN => n30192);
   U6130 : AOI21_X1 port map( A1 => n984, A2 => n1205, B => n1072, ZN => n11147
                           );
   U6133 : INV_X2 port map( I => n28237, ZN => n982);
   U6140 : INV_X1 port map( I => n11694, ZN => n27848);
   U6146 : NAND2_X1 port map( A1 => n27337, A2 => n1225, ZN => n11431);
   U6150 : AOI21_X1 port map( A1 => n991, A2 => n32046, B => n4782, ZN => 
                           n16847);
   U6163 : INV_X1 port map( I => n35750, ZN => n27286);
   U6164 : INV_X1 port map( I => n27446, ZN => n27447);
   U6203 : NAND3_X1 port map( A1 => n26101, A2 => n1021, A3 => n35207, ZN => 
                           n26105);
   U6238 : NOR2_X1 port map( A1 => n39599, A2 => n1024, ZN => n25436);
   U6247 : INV_X1 port map( I => n25694, ZN => n25630);
   U6260 : NAND2_X1 port map( A1 => n24648, A2 => n15850, ZN => n15848);
   U6263 : NAND3_X1 port map( A1 => n16210, A2 => n24660, A3 => n24783, ZN => 
                           n12133);
   U6287 : NAND2_X1 port map( A1 => n1586, A2 => n18302, ZN => n13310);
   U6289 : NAND2_X1 port map( A1 => n32297, A2 => n8175, ZN => n24340);
   U6298 : INV_X1 port map( I => n36552, ZN => n14699);
   U6301 : NOR2_X1 port map( A1 => n7273, A2 => n17709, ZN => n23797);
   U6303 : NOR3_X1 port map( A1 => n14392, A2 => n37045, A3 => n24300, ZN => 
                           n3227);
   U6305 : BUF_X4 port map( I => n23934, Z => n1129);
   U6308 : INV_X1 port map( I => n8116, ZN => n20312);
   U6325 : OAI22_X1 port map( A1 => n23597, A2 => n23314, B1 => n23055, B2 => 
                           n23373, ZN => n23073);
   U6351 : OAI21_X1 port map( A1 => n23115, A2 => n9699, B => n1146, ZN => 
                           n12508);
   U6357 : NAND3_X1 port map( A1 => n11658, A2 => n23098, A3 => n21094, ZN => 
                           n12473);
   U6358 : NOR2_X1 port map( A1 => n33697, A2 => n35576, ZN => n22850);
   U6361 : NAND2_X1 port map( A1 => n23083, A2 => n23190, ZN => n2163);
   U6390 : INV_X1 port map( I => n22181, ZN => n2842);
   U6408 : OAI21_X1 port map( A1 => n21906, A2 => n9886, B => n21908, ZN => 
                           n5305);
   U6416 : NAND3_X1 port map( A1 => n21699, A2 => n1353, A3 => n19709, ZN => 
                           n9424);
   U6423 : NOR2_X1 port map( A1 => n21550, A2 => n21506, ZN => n21765);
   U6429 : INV_X1 port map( I => n695, ZN => n21555);
   U6432 : INV_X1 port map( I => n19516, ZN => n1367);
   U6438 : INV_X1 port map( I => n19822, ZN => n21539);
   U6447 : INV_X1 port map( I => n16333, ZN => n21888);
   U6449 : INV_X1 port map( I => n29657, ZN => n1724);
   U6452 : CLKBUF_X2 port map( I => Key(133), Z => n19816);
   U6458 : CLKBUF_X2 port map( I => Key(37), Z => n19905);
   U6478 : NOR2_X1 port map( A1 => n35187, A2 => n30107, ZN => n19033);
   U6479 : NOR2_X1 port map( A1 => n4378, A2 => n30079, ZN => n6687);
   U6483 : NOR2_X1 port map( A1 => n29721, A2 => n29719, ZN => n5779);
   U6531 : NAND3_X1 port map( A1 => n9143, A2 => n30052, A3 => n1057, ZN => 
                           n9142);
   U6532 : NAND2_X1 port map( A1 => n18816, A2 => n5471, ZN => n2860);
   U6535 : NOR2_X1 port map( A1 => n29862, A2 => n38215, ZN => n13132);
   U6539 : NOR2_X1 port map( A1 => n32906, A2 => n31279, ZN => n12880);
   U6543 : NOR3_X1 port map( A1 => n30154, A2 => n5414, A3 => n892, ZN => n5415
                           );
   U6548 : INV_X1 port map( I => n30049, ZN => n8731);
   U6551 : NAND2_X1 port map( A1 => n30153, A2 => n30192, ZN => n30244);
   U6569 : OR2_X1 port map( A1 => n14559, A2 => n29174, Z => n4387);
   U6576 : INV_X1 port map( I => n28983, ZN => n1413);
   U6586 : OAI21_X1 port map( A1 => n28720, A2 => n33646, B => n4980, ZN => 
                           n16474);
   U6597 : INV_X1 port map( I => n28454, ZN => n12990);
   U6601 : NAND2_X1 port map( A1 => n35182, A2 => n1433, ZN => n17801);
   U6607 : NAND2_X1 port map( A1 => n30304, A2 => n28728, ZN => n28061);
   U6612 : OAI21_X1 port map( A1 => n15792, A2 => n1197, B => n10369, ZN => 
                           n28658);
   U6669 : NAND2_X1 port map( A1 => n27997, A2 => n11461, ZN => n8523);
   U6670 : INV_X1 port map( I => n27997, ZN => n27876);
   U6675 : INV_X1 port map( I => n14456, ZN => n1447);
   U6693 : INV_X2 port map( I => n15410, ZN => n18689);
   U6694 : BUF_X4 port map( I => n18474, Z => n988);
   U6698 : INV_X2 port map( I => n15219, ZN => n16613);
   U6706 : AND3_X1 port map( A1 => n27409, A2 => n7706, A3 => n34689, Z => 
                           n27315);
   U6709 : NOR2_X1 port map( A1 => n18374, A2 => n18743, ZN => n15918);
   U6713 : NAND2_X1 port map( A1 => n27410, A2 => n32131, ZN => n4568);
   U6717 : INV_X1 port map( I => n19529, ZN => n20057);
   U6743 : NAND2_X1 port map( A1 => n8000, A2 => n26269, ZN => n4582);
   U6746 : INV_X1 port map( I => n27043, ZN => n17227);
   U6747 : NAND3_X1 port map( A1 => n26794, A2 => n26793, A3 => n36873, ZN => 
                           n12170);
   U6751 : NAND2_X1 port map( A1 => n26708, A2 => n5960, ZN => n14097);
   U6759 : AND2_X1 port map( A1 => n26815, A2 => n1490, Z => n18956);
   U6780 : OAI21_X1 port map( A1 => n13393, A2 => n26763, B => n26895, ZN => 
                           n12713);
   U6790 : INV_X2 port map( I => n17535, ZN => n1003);
   U6793 : BUF_X2 port map( I => n26803, Z => n1091);
   U6794 : INV_X1 port map( I => n11335, ZN => n26936);
   U6798 : INV_X1 port map( I => n14752, ZN => n16834);
   U6804 : INV_X2 port map( I => n26689, ZN => n17252);
   U6810 : INV_X2 port map( I => n26478, ZN => n1009);
   U6812 : AND2_X1 port map( A1 => n6179, A2 => n25875, Z => n6178);
   U6827 : NAND2_X1 port map( A1 => n15020, A2 => n37582, ZN => n10476);
   U6840 : NOR2_X1 port map( A1 => n7110, A2 => n1101, ZN => n15020);
   U6858 : INV_X1 port map( I => n25900, ZN => n26122);
   U6881 : OAI21_X1 port map( A1 => n25385, A2 => n10158, B => n7284, ZN => 
                           n25353);
   U6886 : NAND2_X1 port map( A1 => n25687, A2 => n14518, ZN => n20122);
   U6888 : NOR3_X1 port map( A1 => n25574, A2 => n18031, A3 => n25614, ZN => 
                           n12097);
   U6895 : NAND3_X1 port map( A1 => n7986, A2 => n8070, A3 => n4947, ZN => 
                           n8770);
   U6904 : NAND3_X1 port map( A1 => n25036, A2 => n19785, A3 => n17894, ZN => 
                           n8863);
   U6916 : INV_X1 port map( I => n25379, ZN => n11951);
   U6921 : INV_X2 port map( I => n25543, ZN => n1539);
   U6955 : NAND2_X1 port map( A1 => n7693, A2 => n5388, ZN => n5387);
   U6960 : NOR3_X1 port map( A1 => n10667, A2 => n934, A3 => n17658, ZN => 
                           n17663);
   U6976 : NOR2_X1 port map( A1 => n24782, A2 => n1121, ZN => n4775);
   U6981 : NOR3_X1 port map( A1 => n39513, A2 => n16502, A3 => n5768, ZN => 
                           n1996);
   U6997 : NAND2_X1 port map( A1 => n23797, A2 => n1586, ZN => n5740);
   U7011 : INV_X2 port map( I => n30447, ZN => n1595);
   U7026 : AND2_X1 port map( A1 => n24223, A2 => n24088, Z => n24089);
   U7031 : INV_X1 port map( I => n24327, ZN => n24229);
   U7034 : INV_X1 port map( I => n205, ZN => n1280);
   U7038 : INV_X1 port map( I => n12519, ZN => n17081);
   U7042 : INV_X4 port map( I => n24241, ZN => n1033);
   U7057 : NOR2_X1 port map( A1 => n5044, A2 => n33747, ZN => n23575);
   U7071 : OAI21_X1 port map( A1 => n13830, A2 => n23506, B => n13833, ZN => 
                           n13829);
   U7075 : NAND3_X1 port map( A1 => n35808, A2 => n9823, A3 => n5083, ZN => 
                           n4290);
   U7085 : NAND2_X1 port map( A1 => n960, A2 => n14477, ZN => n23748);
   U7090 : OAI21_X1 port map( A1 => n21247, A2 => n11970, B => n1862, ZN => 
                           n1861);
   U7098 : NOR2_X1 port map( A1 => n33840, A2 => n14477, ZN => n8239);
   U7107 : NAND2_X1 port map( A1 => n34506, A2 => n23472, ZN => n23746);
   U7120 : NAND3_X1 port map( A1 => n14234, A2 => n22934, A3 => n9699, ZN => 
                           n8101);
   U7133 : NAND3_X1 port map( A1 => n15151, A2 => n23099, A3 => n20570, ZN => 
                           n12472);
   U7139 : NOR3_X1 port map( A1 => n1647, A2 => n38524, A3 => n19865, ZN => 
                           n20362);
   U7145 : OAI21_X1 port map( A1 => n16419, A2 => n1646, B => n19469, ZN => 
                           n13093);
   U7147 : NAND3_X1 port map( A1 => n11913, A2 => n22937, A3 => n1141, ZN => 
                           n11912);
   U7148 : NAND2_X1 port map( A1 => n15330, A2 => n23098, ZN => n22905);
   U7149 : OAI21_X1 port map( A1 => n5581, A2 => n17226, B => n1313, ZN => 
                           n13640);
   U7166 : NAND2_X1 port map( A1 => n22993, A2 => n22866, ZN => n14749);
   U7173 : INV_X1 port map( I => n12315, ZN => n1646);
   U7174 : INV_X1 port map( I => n22857, ZN => n22890);
   U7183 : OR2_X2 port map( A1 => n2386, A2 => n2384, Z => n2383);
   U7191 : NOR2_X1 port map( A1 => n39075, A2 => n1149, ZN => n13570);
   U7192 : NAND2_X1 port map( A1 => n21002, A2 => n21001, ZN => n21000);
   U7193 : NAND3_X1 port map( A1 => n11345, A2 => n1812, A3 => n1866, ZN => 
                           n1865);
   U7195 : NAND2_X1 port map( A1 => n3840, A2 => n17530, ZN => n21958);
   U7200 : NOR2_X1 port map( A1 => n7916, A2 => n22239, ZN => n8118);
   U7207 : NAND3_X1 port map( A1 => n31940, A2 => n11327, A3 => n1672, ZN => 
                           n22218);
   U7214 : INV_X1 port map( I => n22243, ZN => n22241);
   U7218 : NAND3_X1 port map( A1 => n32107, A2 => n4239, A3 => n2910, ZN => 
                           n8623);
   U7228 : INV_X1 port map( I => n22019, ZN => n22084);
   U7231 : INV_X1 port map( I => n18303, ZN => n17086);
   U7233 : BUF_X2 port map( I => n22041, Z => n2839);
   U7237 : BUF_X4 port map( I => n17440, Z => n1048);
   U7239 : INV_X1 port map( I => n22113, ZN => n13191);
   U7243 : OAI21_X1 port map( A1 => n21901, A2 => n21902, B => n35921, ZN => 
                           n5822);
   U7255 : NAND2_X1 port map( A1 => n18576, A2 => n20266, ZN => n2157);
   U7257 : AND2_X1 port map( A1 => n21401, A2 => n668, Z => n9705);
   U7259 : NAND2_X1 port map( A1 => n21817, A2 => n32820, ZN => n21479);
   U7268 : INV_X1 port map( I => n21606, ZN => n2645);
   U7277 : INV_X1 port map( I => n21550, ZN => n21763);
   U7279 : INV_X1 port map( I => n21352, ZN => n4094);
   U7291 : INV_X1 port map( I => n13679, ZN => n21521);
   U7292 : NOR2_X1 port map( A1 => n20778, A2 => n19496, ZN => n21561);
   U7294 : INV_X1 port map( I => n30104, ZN => n1163);
   U7295 : CLKBUF_X2 port map( I => n21330, Z => n21697);
   U7297 : INV_X1 port map( I => n30150, ZN => n1161);
   U7298 : BUF_X2 port map( I => n21938, Z => n8700);
   U7302 : INV_X1 port map( I => n29970, ZN => n1162);
   U7303 : INV_X1 port map( I => n19805, ZN => n1167);
   U7307 : INV_X1 port map( I => n30126, ZN => n1165);
   U7308 : INV_X1 port map( I => n29831, ZN => n1169);
   U7309 : CLKBUF_X2 port map( I => Key(183), Z => n30126);
   U7312 : CLKBUF_X2 port map( I => Key(75), Z => n30179);
   U7320 : CLKBUF_X2 port map( I => Key(27), Z => n29371);
   U7324 : NAND3_X1 port map( A1 => n37632, A2 => n939, A3 => n13142, ZN => 
                           n12452);
   U7331 : NAND2_X1 port map( A1 => n29874, A2 => n17286, ZN => n10293);
   U7332 : NAND2_X1 port map( A1 => n29881, A2 => n17286, ZN => n10292);
   U7334 : OR2_X1 port map( A1 => n35180, A2 => n16084, Z => n16083);
   U7340 : NAND2_X1 port map( A1 => n37632, A2 => n939, ZN => n11973);
   U7341 : AOI21_X1 port map( A1 => n18039, A2 => n15509, B => n939, ZN => 
                           n12033);
   U7342 : NAND2_X1 port map( A1 => n31160, A2 => n8955, ZN => n5813);
   U7349 : NAND2_X1 port map( A1 => n31569, A2 => n29929, ZN => n29912);
   U7351 : INV_X1 port map( I => n31569, ZN => n8561);
   U7354 : INV_X1 port map( I => n29722, ZN => n5951);
   U7357 : NOR2_X1 port map( A1 => n30086, A2 => n30096, ZN => n2484);
   U7376 : AND2_X1 port map( A1 => n2858, A2 => n5579, Z => n2507);
   U7377 : NOR2_X1 port map( A1 => n4377, A2 => n30076, ZN => n30056);
   U7378 : AOI22_X1 port map( A1 => n29708, A2 => n29721, B1 => n29720, B2 => 
                           n14337, ZN => n16577);
   U7383 : INV_X1 port map( I => n4449, ZN => n4447);
   U7384 : NOR2_X1 port map( A1 => n3861, A2 => n5579, ZN => n2073);
   U7387 : INV_X1 port map( I => n13786, ZN => n11701);
   U7392 : NOR2_X1 port map( A1 => n12081, A2 => n19544, ZN => n6863);
   U7405 : NOR2_X1 port map( A1 => n12940, A2 => n33928, ZN => n15584);
   U7406 : NOR2_X1 port map( A1 => n1177, A2 => n1399, ZN => n2321);
   U7411 : NAND3_X1 port map( A1 => n11415, A2 => n30046, A3 => n30162, ZN => 
                           n3819);
   U7416 : OAI21_X1 port map( A1 => n9572, A2 => n13132, B => n18104, ZN => 
                           n9569);
   U7421 : NOR2_X1 port map( A1 => n31511, A2 => n37061, ZN => n28744);
   U7430 : AOI21_X1 port map( A1 => n2160, A2 => n8529, B => n16224, ZN => 
                           n18445);
   U7433 : INV_X1 port map( I => n30232, ZN => n15062);
   U7436 : NAND2_X1 port map( A1 => n19137, A2 => n29892, ZN => n6803);
   U7450 : NOR2_X1 port map( A1 => n19050, A2 => n30220, ZN => n4807);
   U7455 : NOR2_X1 port map( A1 => n21167, A2 => n39828, ZN => n15301);
   U7456 : AND2_X1 port map( A1 => n18816, A2 => n3631, Z => n4445);
   U7457 : NAND2_X1 port map( A1 => n29998, A2 => n30043, ZN => n4858);
   U7464 : AND3_X1 port map( A1 => n19765, A2 => n10590, A3 => n30229, Z => 
                           n9996);
   U7465 : NAND2_X1 port map( A1 => n17597, A2 => n19783, ZN => n29317);
   U7473 : NOR2_X1 port map( A1 => n30238, A2 => n31788, ZN => n11886);
   U7496 : INV_X1 port map( I => n4341, ZN => n29048);
   U7506 : NOR2_X1 port map( A1 => n28360, A2 => n14677, ZN => n16475);
   U7520 : OAI21_X1 port map( A1 => n35172, A2 => n28484, B => n32543, ZN => 
                           n6694);
   U7524 : INV_X2 port map( I => n5115, ZN => n1065);
   U7533 : OAI22_X1 port map( A1 => n28765, A2 => n35203, B1 => n28812, B2 => 
                           n5465, ZN => n12545);
   U7537 : NOR2_X1 port map( A1 => n1431, A2 => n28553, ZN => n8759);
   U7548 : NAND3_X1 port map( A1 => n15447, A2 => n39355, A3 => n19827, ZN => 
                           n6071);
   U7551 : NAND2_X1 port map( A1 => n976, A2 => n35203, ZN => n8914);
   U7559 : NAND2_X1 port map( A1 => n9329, A2 => n17771, ZN => n10676);
   U7563 : NAND3_X1 port map( A1 => n15112, A2 => n9141, A3 => n5093, ZN => 
                           n16183);
   U7564 : INV_X1 port map( I => n1882, ZN => n18369);
   U7571 : NOR2_X1 port map( A1 => n5383, A2 => n39435, ZN => n12611);
   U7576 : NOR2_X1 port map( A1 => n2790, A2 => n28723, ZN => n2785);
   U7580 : NOR2_X1 port map( A1 => n28323, A2 => n30304, ZN => n17596);
   U7600 : INV_X1 port map( I => n28569, ZN => n28614);
   U7608 : NAND2_X1 port map( A1 => n10825, A2 => n27980, ZN => n10824);
   U7618 : NAND2_X1 port map( A1 => n8787, A2 => n20445, ZN => n28612);
   U7637 : OAI21_X1 port map( A1 => n28064, A2 => n16513, B => n981, ZN => 
                           n6980);
   U7638 : AOI21_X1 port map( A1 => n27624, A2 => n37056, B => n16576, ZN => 
                           n7365);
   U7641 : AOI21_X1 port map( A1 => n16576, A2 => n8960, B => n35694, ZN => 
                           n9170);
   U7653 : NAND3_X1 port map( A1 => n10836, A2 => n983, A3 => n28050, ZN => 
                           n10443);
   U7660 : NAND2_X1 port map( A1 => n27900, A2 => n16461, ZN => n8525);
   U7672 : AND2_X1 port map( A1 => n14397, A2 => n1200, Z => n4456);
   U7673 : NAND2_X1 port map( A1 => n2716, A2 => n5266, ZN => n5905);
   U7679 : NOR2_X1 port map( A1 => n37, A2 => n1448, ZN => n11838);
   U7726 : INV_X1 port map( I => n27964, ZN => n28137);
   U7736 : BUF_X2 port map( I => n16339, Z => n11461);
   U7747 : INV_X1 port map( I => n17378, ZN => n27997);
   U7749 : INV_X1 port map( I => n39442, ZN => n7755);
   U7753 : INV_X1 port map( I => n27556, ZN => n14325);
   U7755 : INV_X1 port map( I => n27574, ZN => n1215);
   U7765 : NAND2_X1 port map( A1 => n30871, A2 => n35115, ZN => n18050);
   U7768 : AOI21_X1 port map( A1 => n26941, A2 => n12156, B => n18489, ZN => 
                           n26942);
   U7787 : AND2_X1 port map( A1 => n4434, A2 => n34689, Z => n11735);
   U7789 : OR2_X1 port map( A1 => n39065, A2 => n1470, Z => n26967);
   U7791 : OAI21_X1 port map( A1 => n33593, A2 => n36496, B => n16782, ZN => 
                           n4231);
   U7794 : NAND2_X1 port map( A1 => n992, A2 => n1227, ZN => n2259);
   U7822 : AND2_X1 port map( A1 => n34562, A2 => n19203, Z => n4610);
   U7831 : NOR3_X1 port map( A1 => n20402, A2 => n17795, A3 => n27123, ZN => 
                           n6415);
   U7837 : NOR2_X1 port map( A1 => n33503, A2 => n7975, ZN => n6975);
   U7838 : INV_X2 port map( I => n7611, ZN => n12156);
   U7840 : OAI21_X1 port map( A1 => n26767, A2 => n9690, B => n33396, ZN => 
                           n8331);
   U7843 : OR2_X1 port map( A1 => n11467, A2 => n14412, Z => n3809);
   U7849 : NOR2_X1 port map( A1 => n26639, A2 => n17515, ZN => n26767);
   U7854 : NOR2_X1 port map( A1 => n26859, A2 => n32256, ZN => n14469);
   U7864 : OAI21_X1 port map( A1 => n19206, A2 => n19207, B => n38797, ZN => 
                           n9891);
   U7865 : OR2_X1 port map( A1 => n13854, A2 => n26988, Z => n13334);
   U7883 : NOR2_X1 port map( A1 => n19448, A2 => n8556, ZN => n11130);
   U7885 : NAND2_X1 port map( A1 => n3350, A2 => n7527, ZN => n3349);
   U7889 : NAND2_X1 port map( A1 => n26962, A2 => n17601, ZN => n17600);
   U7893 : NAND3_X1 port map( A1 => n13605, A2 => n5405, A3 => n35912, ZN => 
                           n26642);
   U7900 : AND2_X1 port map( A1 => n26922, A2 => n26895, Z => n26304);
   U7923 : AND2_X1 port map( A1 => n26961, A2 => n20936, Z => n3224);
   U7929 : OAI21_X1 port map( A1 => n14355, A2 => n7752, B => n3351, ZN => 
                           n3350);
   U7955 : INV_X1 port map( I => n26666, ZN => n26179);
   U7959 : NAND2_X1 port map( A1 => n11105, A2 => n26598, ZN => n3098);
   U7974 : AND2_X1 port map( A1 => n26000, A2 => n13971, Z => n16239);
   U7981 : NAND2_X1 port map( A1 => n16200, A2 => n1017, ZN => n10138);
   U7987 : NOR2_X1 port map( A1 => n2835, A2 => n2833, ZN => n2832);
   U7995 : AND2_X1 port map( A1 => n25847, A2 => n1514, Z => n11770);
   U8005 : OAI21_X1 port map( A1 => n25867, A2 => n37306, B => n26022, ZN => 
                           n21198);
   U8011 : OAI21_X1 port map( A1 => n4190, A2 => n26125, B => n929, ZN => n6883
                           );
   U8023 : NAND3_X1 port map( A1 => n31192, A2 => n2888, A3 => n4772, ZN => 
                           n12448);
   U8025 : NAND2_X1 port map( A1 => n18289, A2 => n26075, ZN => n26076);
   U8048 : AND2_X1 port map( A1 => n1521, A2 => n2534, Z => n11386);
   U8056 : NAND2_X1 port map( A1 => n26029, A2 => n18320, ZN => n25922);
   U8063 : NAND2_X1 port map( A1 => n31133, A2 => n31626, ZN => n8255);
   U8064 : OAI21_X1 port map( A1 => n8883, A2 => n18142, B => n17791, ZN => 
                           n7732);
   U8073 : INV_X2 port map( I => n18320, ZN => n1102);
   U8074 : BUF_X2 port map( I => n7136, Z => n7110);
   U8089 : OR2_X1 port map( A1 => n13467, A2 => n954, Z => n13466);
   U8091 : NAND3_X1 port map( A1 => n5860, A2 => n32105, A3 => n25452, ZN => 
                           n5858);
   U8097 : NAND2_X1 port map( A1 => n4455, A2 => n13129, ZN => n4452);
   U8101 : NOR2_X1 port map( A1 => n728, A2 => n2799, ZN => n5455);
   U8113 : NAND2_X1 port map( A1 => n1539, A2 => n25482, ZN => n2250);
   U8115 : NAND3_X1 port map( A1 => n1253, A2 => n16677, A3 => n24896, ZN => 
                           n17303);
   U8119 : AND2_X1 port map( A1 => n17029, A2 => n36708, Z => n9429);
   U8121 : NOR2_X1 port map( A1 => n5227, A2 => n12500, ZN => n5010);
   U8135 : OAI22_X1 port map( A1 => n14081, A2 => n14082, B1 => n25642, B2 => 
                           n25674, ZN => n14056);
   U8143 : NAND3_X1 port map( A1 => n1545, A2 => n6747, A3 => n25361, ZN => 
                           n9145);
   U8155 : OAI21_X1 port map( A1 => n16933, A2 => n25482, B => n25548, ZN => 
                           n10786);
   U8179 : INV_X1 port map( I => n20924, ZN => n25533);
   U8180 : OR2_X1 port map( A1 => n15052, A2 => n15051, Z => n25548);
   U8186 : INV_X1 port map( I => n25722, ZN => n25721);
   U8190 : BUF_X4 port map( I => n3785, Z => n25361);
   U8196 : INV_X2 port map( I => n825, ZN => n1257);
   U8198 : INV_X1 port map( I => n11497, ZN => n7876);
   U8201 : INV_X1 port map( I => n25176, ZN => n1554);
   U8203 : NAND3_X1 port map( A1 => n25203, A2 => n7968, A3 => n7969, ZN => 
                           n3653);
   U8208 : OR2_X1 port map( A1 => n20800, A2 => n4973, Z => n16747);
   U8215 : NAND2_X1 port map( A1 => n7065, A2 => n24608, ZN => n4908);
   U8244 : NOR2_X1 port map( A1 => n7693, A2 => n10116, ZN => n20689);
   U8249 : AND2_X1 port map( A1 => n24887, A2 => n15467, Z => n16745);
   U8263 : NOR2_X1 port map( A1 => n7286, A2 => n19420, ZN => n8954);
   U8274 : INV_X1 port map( I => n24565, ZN => n1573);
   U8277 : INV_X2 port map( I => n24673, ZN => n16547);
   U8284 : NOR2_X1 port map( A1 => n1586, A2 => n37227, ZN => n19027);
   U8290 : AOI21_X1 port map( A1 => n4666, A2 => n24153, B => n16377, ZN => 
                           n24154);
   U8291 : OAI21_X1 port map( A1 => n19466, A2 => n24303, B => n21310, ZN => 
                           n11170);
   U8293 : NOR3_X1 port map( A1 => n15240, A2 => n12975, A3 => n1608, ZN => 
                           n20653);
   U8294 : INV_X1 port map( I => n3133, ZN => n8175);
   U8300 : NOR2_X1 port map( A1 => n12366, A2 => n7086, ZN => n7085);
   U8317 : OR2_X1 port map( A1 => n6933, A2 => n33450, Z => n12974);
   U8322 : NAND2_X1 port map( A1 => n33712, A2 => n24245, ZN => n24582);
   U8323 : NOR2_X1 port map( A1 => n24274, A2 => n35954, ZN => n5358);
   U8327 : OAI21_X1 port map( A1 => n12975, A2 => n24087, B => n1608, ZN => 
                           n7406);
   U8331 : INV_X1 port map( I => n38224, ZN => n19653);
   U8341 : INV_X2 port map( I => n39816, ZN => n1596);
   U8357 : CLKBUF_X2 port map( I => n39814, Z => n7440);
   U8371 : AOI22_X1 port map( A1 => n21251, A2 => n21130, B1 => n1633, B2 => 
                           n21250, ZN => n12175);
   U8375 : NAND2_X1 port map( A1 => n3715, A2 => n31644, ZN => n2919);
   U8380 : NOR3_X1 port map( A1 => n10480, A2 => n9395, A3 => n33496, ZN => 
                           n1918);
   U8385 : NOR2_X1 port map( A1 => n1290, A2 => n9862, ZN => n12851);
   U8388 : OAI21_X1 port map( A1 => n20841, A2 => n1308, B => n33349, ZN => 
                           n17442);
   U8421 : NOR2_X1 port map( A1 => n36810, A2 => n33703, ZN => n23243);
   U8431 : NAND2_X1 port map( A1 => n19559, A2 => n13733, ZN => n1862);
   U8439 : INV_X4 port map( I => n2600, ZN => n23567);
   U8443 : INV_X1 port map( I => n23516, ZN => n1623);
   U8466 : OAI22_X1 port map( A1 => n20637, A2 => n23209, B1 => n5464, B2 => 
                           n23135, ZN => n23136);
   U8469 : NAND2_X1 port map( A1 => n35442, A2 => n8812, ZN => n19181);
   U8470 : NOR2_X1 port map( A1 => n1319, A2 => n1654, ZN => n6500);
   U8473 : OAI21_X1 port map( A1 => n1645, A2 => n23124, B => n22875, ZN => 
                           n13450);
   U8486 : NOR2_X1 port map( A1 => n22890, A2 => n22682, ZN => n15242);
   U8489 : NAND2_X1 port map( A1 => n38601, A2 => n23212, ZN => n3041);
   U8494 : OR2_X1 port map( A1 => n18229, A2 => n19697, Z => n13337);
   U8512 : OR2_X1 port map( A1 => n39810, A2 => n2047, Z => n2049);
   U8517 : OAI21_X1 port map( A1 => n19440, A2 => n19134, B => n23124, ZN => 
                           n14187);
   U8542 : INV_X1 port map( I => n34757, ZN => n23172);
   U8545 : INV_X2 port map( I => n13572, ZN => n1145);
   U8548 : INV_X1 port map( I => n23122, ZN => n11295);
   U8552 : BUF_X2 port map( I => n12315, Z => n5657);
   U8563 : AND2_X2 port map( A1 => n5205, A2 => n5204, Z => n5203);
   U8564 : NAND2_X1 port map( A1 => n37089, A2 => n34808, ZN => n4851);
   U8568 : NAND2_X1 port map( A1 => n22340, A2 => n20238, ZN => n10630);
   U8569 : NOR2_X1 port map( A1 => n30800, A2 => n11329, ZN => n7896);
   U8570 : NAND2_X1 port map( A1 => n22143, A2 => n34808, ZN => n8753);
   U8574 : NAND2_X1 port map( A1 => n19261, A2 => n1329, ZN => n5877);
   U8580 : AND3_X1 port map( A1 => n31940, A2 => n11171, A3 => n22361, Z => 
                           n4800);
   U8584 : NAND2_X1 port map( A1 => n32889, A2 => n5929, ZN => n21969);
   U8585 : NOR2_X1 port map( A1 => n11329, A2 => n5302, ZN => n9484);
   U8598 : OR2_X1 port map( A1 => n32889, A2 => n5929, Z => n11511);
   U8599 : NOR2_X1 port map( A1 => n21503, A2 => n30306, ZN => n19453);
   U8605 : NAND2_X1 port map( A1 => n474, A2 => n14349, ZN => n2211);
   U8610 : NOR2_X1 port map( A1 => n6576, A2 => n36397, ZN => n5617);
   U8612 : NOR2_X1 port map( A1 => n32107, A2 => n14423, ZN => n8622);
   U8614 : NAND2_X1 port map( A1 => n17685, A2 => n12077, ZN => n12930);
   U8615 : NAND3_X1 port map( A1 => n18360, A2 => n1344, A3 => n22086, ZN => 
                           n9341);
   U8620 : NOR2_X1 port map( A1 => n2839, A2 => n1338, ZN => n14028);
   U8621 : NAND2_X1 port map( A1 => n19958, A2 => n6297, ZN => n14233);
   U8627 : NOR2_X1 port map( A1 => n1338, A2 => n18303, ZN => n7434);
   U8629 : AOI21_X1 port map( A1 => n6347, A2 => n22019, B => n36006, ZN => 
                           n5462);
   U8632 : INV_X2 port map( I => n4179, ZN => n12814);
   U8635 : NOR2_X1 port map( A1 => n6347, A2 => n2696, ZN => n21664);
   U8636 : BUF_X2 port map( I => n22497, Z => n7131);
   U8638 : NAND4_X1 port map( A1 => n5304, A2 => n5303, A3 => n5305, A4 => 
                           n7608, ZN => n5302);
   U8641 : NAND2_X1 port map( A1 => n7357, A2 => n22364, ZN => n12169);
   U8649 : INV_X2 port map( I => n22354, ZN => n1152);
   U8650 : NAND3_X1 port map( A1 => n2278, A2 => n21817, A3 => n2092, ZN => 
                           n2276);
   U8656 : OAI22_X1 port map( A1 => n13701, A2 => n21898, B1 => n21838, B2 => 
                           n10120, ZN => n10085);
   U8659 : AOI22_X1 port map( A1 => n543, A2 => n6418, B1 => n33771, B2 => 
                           n21765, ZN => n6417);
   U8667 : AOI22_X1 port map( A1 => n15031, A2 => n275, B1 => n21440, B2 => 
                           n18152, ZN => n5823);
   U8668 : OR2_X1 port map( A1 => n2759, A2 => n18219, Z => n9746);
   U8669 : NAND3_X1 port map( A1 => n20898, A2 => n21899, A3 => n21897, ZN => 
                           n3438);
   U8670 : NAND2_X1 port map( A1 => n38011, A2 => n5531, ZN => n5023);
   U8676 : NOR2_X1 port map( A1 => n18774, A2 => n14373, ZN => n19554);
   U8685 : NOR2_X1 port map( A1 => n9642, A2 => n20328, ZN => n15706);
   U8688 : NOR2_X1 port map( A1 => n33771, A2 => n21761, ZN => n6418);
   U8692 : NOR2_X1 port map( A1 => n1346, A2 => n5751, ZN => n9286);
   U8693 : NOR2_X1 port map( A1 => n15839, A2 => n3784, ZN => n15523);
   U8696 : NAND2_X1 port map( A1 => n7703, A2 => n7654, ZN => n10822);
   U8700 : INV_X1 port map( I => n21475, ZN => n6350);
   U8701 : NAND2_X1 port map( A1 => n33154, A2 => n21912, ZN => n13437);
   U8704 : NOR2_X1 port map( A1 => n8799, A2 => n21898, ZN => n15369);
   U8706 : NAND2_X1 port map( A1 => n8293, A2 => n21339, ZN => n7367);
   U8707 : AND2_X1 port map( A1 => n21666, A2 => n690, Z => n10464);
   U8709 : INV_X1 port map( I => n21905, ZN => n21462);
   U8710 : INV_X1 port map( I => n21894, ZN => n21581);
   U8720 : INV_X1 port map( I => n21898, ZN => n1694);
   U8724 : NAND2_X1 port map( A1 => n7304, A2 => n526, ZN => n16035);
   U8725 : INV_X2 port map( I => n18450, ZN => n21897);
   U8726 : INV_X1 port map( I => n13997, ZN => n18496);
   U8727 : NOR2_X1 port map( A1 => n19395, A2 => n21875, ZN => n11916);
   U8728 : AOI21_X1 port map( A1 => n21546, A2 => n21696, B => n21330, ZN => 
                           n11917);
   U8732 : INV_X1 port map( I => n29649, ZN => n1708);
   U8733 : INV_X1 port map( I => n19804, ZN => n1371);
   U8734 : INV_X1 port map( I => n29666, ZN => n1361);
   U8735 : INV_X1 port map( I => n15370, ZN => n12044);
   U8737 : INV_X1 port map( I => n19683, ZN => n1356);
   U8739 : INV_X1 port map( I => n19720, ZN => n1370);
   U8740 : INV_X1 port map( I => n19622, ZN => n1358);
   U8741 : INV_X1 port map( I => n29506, ZN => n1357);
   U8744 : INV_X1 port map( I => n30010, ZN => n1374);
   U8746 : BUF_X2 port map( I => n19871, Z => n20328);
   U8750 : INV_X1 port map( I => n18270, ZN => n23591);
   U8752 : INV_X1 port map( I => n19800, ZN => n1366);
   U8753 : INV_X1 port map( I => n29978, ZN => n1368);
   U8756 : CLKBUF_X2 port map( I => Key(62), Z => n19800);
   U8759 : CLKBUF_X2 port map( I => Key(153), Z => n19786);
   U8762 : CLKBUF_X2 port map( I => Key(157), Z => n19720);
   U8763 : CLKBUF_X2 port map( I => Key(24), Z => n19925);
   U8764 : CLKBUF_X2 port map( I => Key(17), Z => n30101);
   U8765 : CLKBUF_X2 port map( I => Key(118), Z => n19683);
   U8767 : CLKBUF_X2 port map( I => Key(15), Z => n30016);
   U8768 : CLKBUF_X2 port map( I => Key(10), Z => n19622);
   U8772 : CLKBUF_X2 port map( I => Key(94), Z => n19516);
   U8773 : CLKBUF_X2 port map( I => Key(168), Z => n19902);
   U8781 : CLKBUF_X2 port map( I => Key(173), Z => n19940);
   U8789 : CLKBUF_X2 port map( I => Key(78), Z => n19629);
   U8790 : CLKBUF_X2 port map( I => Key(113), Z => n29538);
   U8794 : NAND3_X1 port map( A1 => n29369, A2 => n11067, A3 => n15768, ZN => 
                           n4669);
   U8795 : OAI21_X1 port map( A1 => n1380, A2 => n6147, B => n7600, ZN => 
                           n16472);
   U8802 : NOR2_X1 port map( A1 => n17369, A2 => n16598, ZN => n16597);
   U8804 : NOR2_X1 port map( A1 => n2489, A2 => n6147, ZN => n2488);
   U8806 : INV_X1 port map( I => n1385, ZN => n11448);
   U8808 : AOI21_X1 port map( A1 => n969, A2 => n38200, B => n6341, ZN => n6340
                           );
   U8811 : INV_X1 port map( I => n29219, ZN => n1378);
   U8812 : OAI21_X1 port map( A1 => n29812, A2 => n29811, B => n38141, ZN => 
                           n6441);
   U8815 : AOI21_X1 port map( A1 => n11898, A2 => n29859, B => n36764, ZN => 
                           n2506);
   U8816 : OAI21_X1 port map( A1 => n15601, A2 => n8955, B => n968, ZN => 
                           n11972);
   U8818 : AOI21_X1 port map( A1 => n8561, A2 => n19097, B => n18081, ZN => 
                           n8560);
   U8819 : AOI21_X1 port map( A1 => n29851, A2 => n11898, B => n29855, ZN => 
                           n5580);
   U8826 : BUF_X2 port map( I => n33966, Z => n10003);
   U8828 : NAND2_X1 port map( A1 => n29318, A2 => n38156, ZN => n9627);
   U8829 : AOI21_X1 port map( A1 => n6147, A2 => n30096, B => n13559, ZN => 
                           n6149);
   U8830 : NAND2_X1 port map( A1 => n13442, A2 => n29574, ZN => n14075);
   U8832 : NOR2_X1 port map( A1 => n2944, A2 => n5579, ZN => n29846);
   U8834 : OAI21_X1 port map( A1 => n29756, A2 => n29754, B => n29739, ZN => 
                           n8063);
   U8838 : INV_X2 port map( I => n29980, ZN => n1170);
   U8849 : OAI21_X1 port map( A1 => n30192, A2 => n30153, B => n30152, ZN => 
                           n5300);
   U8857 : NAND2_X1 port map( A1 => n28996, A2 => n1057, ZN => n7167);
   U8859 : NOR3_X1 port map( A1 => n31629, A2 => n6019, A3 => n34179, ZN => 
                           n6372);
   U8860 : AOI21_X1 port map( A1 => n6851, A2 => n8918, B => n32946, ZN => 
                           n12992);
   U8864 : NAND2_X1 port map( A1 => n7208, A2 => n4169, ZN => n21052);
   U8873 : NOR2_X1 port map( A1 => n29777, A2 => n17726, ZN => n15424);
   U8876 : NOR2_X1 port map( A1 => n7789, A2 => n29059, ZN => n7989);
   U8878 : NAND2_X1 port map( A1 => n29595, A2 => n1404, ZN => n6254);
   U8881 : NOR2_X1 port map( A1 => n16907, A2 => n7790, ZN => n7479);
   U8882 : NOR2_X1 port map( A1 => n29904, A2 => n6204, ZN => n6203);
   U8883 : NOR2_X1 port map( A1 => n1402, A2 => n29776, ZN => n7448);
   U8886 : NOR2_X1 port map( A1 => n21074, A2 => n30041, ZN => n9817);
   U8888 : NOR2_X1 port map( A1 => n30041, A2 => n21074, ZN => n20125);
   U8890 : NOR2_X1 port map( A1 => n5736, A2 => n3986, ZN => n3154);
   U8893 : BUF_X2 port map( I => n14438, Z => n2121);
   U8897 : NOR2_X1 port map( A1 => n29992, A2 => n775, ZN => n3169);
   U8898 : NOR2_X1 port map( A1 => n1060, A2 => n29699, ZN => n9000);
   U8899 : NOR2_X1 port map( A1 => n14891, A2 => n18667, ZN => n11635);
   U8910 : INV_X1 port map( I => n29450, ZN => n29418);
   U8917 : INV_X1 port map( I => n29907, ZN => n29955);
   U8919 : INV_X2 port map( I => n29493, ZN => n1179);
   U8920 : INV_X1 port map( I => n16009, ZN => n19994);
   U8928 : NAND3_X1 port map( A1 => n28632, A2 => n28634, A3 => n14209, ZN => 
                           n28636);
   U8937 : NAND2_X1 port map( A1 => n10303, A2 => n32014, ZN => n10302);
   U8945 : NAND3_X1 port map( A1 => n28453, A2 => n13379, A3 => n9668, ZN => 
                           n13378);
   U8948 : NOR2_X1 port map( A1 => n28759, A2 => n3014, ZN => n28408);
   U8955 : NAND2_X1 port map( A1 => n17800, A2 => n11164, ZN => n14239);
   U8964 : AOI21_X1 port map( A1 => n8093, A2 => n3845, B => n28473, ZN => 
                           n8159);
   U8965 : NOR2_X1 port map( A1 => n28514, A2 => n28716, ZN => n5243);
   U8968 : INV_X2 port map( I => n9878, ZN => n11488);
   U8971 : NAND2_X1 port map( A1 => n5343, A2 => n28735, ZN => n5342);
   U8974 : NOR2_X1 port map( A1 => n2639, A2 => n8476, ZN => n13061);
   U8986 : NAND2_X1 port map( A1 => n28570, A2 => n39020, ZN => n19322);
   U9004 : INV_X1 port map( I => n28715, ZN => n28509);
   U9005 : NAND2_X1 port map( A1 => n3899, A2 => n979, ZN => n4119);
   U9013 : INV_X2 port map( I => n9597, ZN => n13508);
   U9022 : NOR2_X1 port map( A1 => n39786, A2 => n32080, ZN => n11743);
   U9031 : OAI21_X1 port map( A1 => n28048, A2 => n28258, B => n11025, ZN => 
                           n11024);
   U9049 : NOR2_X1 port map( A1 => n27915, A2 => n1451, ZN => n19748);
   U9053 : NOR2_X1 port map( A1 => n11461, A2 => n28001, ZN => n8801);
   U9054 : OR2_X1 port map( A1 => n1439, A2 => n1441, Z => n18777);
   U9063 : NAND2_X1 port map( A1 => n28206, A2 => n156, ZN => n4977);
   U9072 : NOR2_X1 port map( A1 => n32783, A2 => n15357, ZN => n10236);
   U9077 : NOR2_X1 port map( A1 => n28258, A2 => n34410, ZN => n27883);
   U9083 : NOR2_X1 port map( A1 => n28236, A2 => n2262, ZN => n4153);
   U9086 : NAND3_X1 port map( A1 => n27894, A2 => n17410, A3 => n28273, ZN => 
                           n20639);
   U9090 : NAND2_X1 port map( A1 => n36517, A2 => n13366, ZN => n11407);
   U9094 : NOR3_X1 port map( A1 => n13927, A2 => n11461, A3 => n28200, ZN => 
                           n13906);
   U9102 : AND2_X1 port map( A1 => n15357, A2 => n1447, Z => n14615);
   U9103 : NAND2_X1 port map( A1 => n28236, A2 => n28237, ZN => n12623);
   U9104 : INV_X1 port map( I => n38202, ZN => n3511);
   U9116 : NOR2_X1 port map( A1 => n17410, A2 => n14399, ZN => n12477);
   U9117 : NAND2_X1 port map( A1 => n12257, A2 => n28230, ZN => n27063);
   U9137 : INV_X2 port map( I => n18383, ZN => n1212);
   U9142 : INV_X2 port map( I => n15287, ZN => n1214);
   U9151 : NAND2_X1 port map( A1 => n9037, A2 => n27395, ZN => n3851);
   U9156 : NOR2_X1 port map( A1 => n38488, A2 => n6191, ZN => n7499);
   U9159 : NAND3_X1 port map( A1 => n13213, A2 => n7975, A3 => n7676, ZN => 
                           n21232);
   U9160 : NAND2_X1 port map( A1 => n27084, A2 => n5675, ZN => n16360);
   U9163 : NOR2_X1 port map( A1 => n9488, A2 => n1481, ZN => n9487);
   U9176 : NOR2_X1 port map( A1 => n1473, A2 => n17132, ZN => n17422);
   U9184 : AND2_X1 port map( A1 => n26074, A2 => n1470, Z => n11485);
   U9185 : OAI21_X1 port map( A1 => n10581, A2 => n9633, B => n38193, ZN => 
                           n10577);
   U9199 : NAND2_X1 port map( A1 => n39628, A2 => n15616, ZN => n7921);
   U9208 : NAND2_X1 port map( A1 => n27285, A2 => n33254, ZN => n10284);
   U9211 : NAND2_X1 port map( A1 => n1480, A2 => n33503, ZN => n27119);
   U9213 : OR2_X1 port map( A1 => n19455, A2 => n27197, Z => n6507);
   U9221 : NAND2_X1 port map( A1 => n5089, A2 => n27284, ZN => n27285);
   U9224 : NOR2_X1 port map( A1 => n27357, A2 => n15360, ZN => n5559);
   U9231 : NAND2_X1 port map( A1 => n7975, A2 => n9144, ZN => n6972);
   U9235 : NOR2_X1 port map( A1 => n27127, A2 => n27126, ZN => n27128);
   U9247 : NAND2_X1 port map( A1 => n12373, A2 => n9690, ZN => n4325);
   U9252 : NOR2_X1 port map( A1 => n15594, A2 => n26804, ZN => n10891);
   U9256 : OAI21_X1 port map( A1 => n32168, A2 => n26970, B => n2226, ZN => 
                           n26250);
   U9263 : NOR2_X1 port map( A1 => n2079, A2 => n36801, ZN => n2078);
   U9269 : NAND2_X1 port map( A1 => n18870, A2 => n15485, ZN => n26750);
   U9275 : NOR3_X1 port map( A1 => n20120, A2 => n26802, A3 => n8479, ZN => 
                           n2801);
   U9278 : NAND3_X1 port map( A1 => n33333, A2 => n6606, A3 => n26932, ZN => 
                           n14457);
   U9295 : NOR2_X1 port map( A1 => n19762, A2 => n36882, ZN => n18901);
   U9296 : AND2_X1 port map( A1 => n26719, A2 => n10111, Z => n26471);
   U9298 : OR2_X1 port map( A1 => n20936, A2 => n33858, Z => n12505);
   U9304 : NAND2_X1 port map( A1 => n34160, A2 => n26968, ZN => n2079);
   U9306 : NAND2_X1 port map( A1 => n17515, A2 => n6454, ZN => n16402);
   U9312 : NOR2_X1 port map( A1 => n26862, A2 => n17712, ZN => n9731);
   U9313 : AOI21_X1 port map( A1 => n26783, A2 => n8814, B => n8817, ZN => 
                           n26784);
   U9314 : INV_X2 port map( I => n26768, ZN => n10355);
   U9332 : NOR2_X1 port map( A1 => n26734, A2 => n4138, ZN => n10202);
   U9337 : NAND2_X1 port map( A1 => n14382, A2 => n13004, ZN => n7778);
   U9338 : NAND3_X1 port map( A1 => n13777, A2 => n875, A3 => n26937, ZN => 
                           n18024);
   U9342 : INV_X1 port map( I => n3449, ZN => n26773);
   U9347 : NOR2_X1 port map( A1 => n34005, A2 => n26901, ZN => n5174);
   U9352 : INV_X1 port map( I => n9117, ZN => n26910);
   U9354 : INV_X2 port map( I => n11188, ZN => n26961);
   U9355 : INV_X2 port map( I => n20974, ZN => n26935);
   U9356 : BUF_X2 port map( I => n26713, Z => n19425);
   U9368 : AOI22_X1 port map( A1 => n25846, A2 => n25928, B1 => n25847, B2 => 
                           n26116, ZN => n12489);
   U9372 : NAND3_X1 port map( A1 => n11552, A2 => n18406, A3 => n318, ZN => 
                           n25896);
   U9376 : NOR2_X1 port map( A1 => n25928, A2 => n4154, ZN => n7544);
   U9377 : OAI21_X1 port map( A1 => n25971, A2 => n951, B => n14215, ZN => 
                           n3916);
   U9381 : OAI21_X1 port map( A1 => n31192, A2 => n7961, B => n26088, ZN => 
                           n20490);
   U9386 : OAI21_X1 port map( A1 => n25868, A2 => n31375, B => n5885, ZN => 
                           n5884);
   U9392 : OR2_X1 port map( A1 => n25822, A2 => n1511, Z => n14660);
   U9399 : OAI21_X1 port map( A1 => n26125, A2 => n4190, B => n4515, ZN => 
                           n26011);
   U9403 : NOR2_X1 port map( A1 => n14703, A2 => n6222, ZN => n12449);
   U9406 : NAND3_X1 port map( A1 => n31375, A2 => n26020, A3 => n25867, ZN => 
                           n5885);
   U9423 : NAND3_X1 port map( A1 => n38247, A2 => n18801, A3 => n25820, ZN => 
                           n25706);
   U9427 : NAND2_X1 port map( A1 => n36546, A2 => n2888, ZN => n14703);
   U9429 : NOR2_X1 port map( A1 => n25829, A2 => n17624, ZN => n6062);
   U9431 : NOR2_X1 port map( A1 => n26055, A2 => n38198, ZN => n25744);
   U9433 : NAND2_X1 port map( A1 => n26185, A2 => n38185, ZN => n17952);
   U9438 : INV_X1 port map( I => n25936, ZN => n26130);
   U9441 : NOR2_X1 port map( A1 => n19121, A2 => n35138, ZN => n19120);
   U9445 : INV_X1 port map( I => n4382, ZN => n4385);
   U9466 : NAND2_X1 port map( A1 => n25349, A2 => n25073, ZN => n25108);
   U9471 : OAI21_X1 port map( A1 => n15543, A2 => n15541, B => n15542, ZN => 
                           n15184);
   U9480 : OR2_X1 port map( A1 => n35157, A2 => n15541, Z => n25593);
   U9481 : AOI21_X1 port map( A1 => n4726, A2 => n25575, B => n25574, ZN => 
                           n16466);
   U9484 : NAND2_X1 port map( A1 => n19095, A2 => n19171, ZN => n20358);
   U9485 : NOR3_X1 port map( A1 => n12896, A2 => n6747, A3 => n25361, ZN => 
                           n6748);
   U9486 : AOI22_X1 port map( A1 => n8879, A2 => n31780, B1 => n953, B2 => 
                           n1548, ZN => n12062);
   U9490 : OAI22_X1 port map( A1 => n1117, A2 => n25380, B1 => n19863, B2 => 
                           n1109, ZN => n7173);
   U9492 : INV_X1 port map( I => n33950, ZN => n18894);
   U9493 : NAND2_X1 port map( A1 => n25571, A2 => n19235, ZN => n19234);
   U9494 : NAND2_X1 port map( A1 => n25480, A2 => n10786, ZN => n10785);
   U9496 : NAND3_X1 port map( A1 => n18298, A2 => n25649, A3 => n32291, ZN => 
                           n25650);
   U9513 : NAND2_X1 port map( A1 => n13218, A2 => n19235, ZN => n20876);
   U9519 : NAND2_X1 port map( A1 => n25481, A2 => n25543, ZN => n12625);
   U9521 : NAND2_X1 port map( A1 => n1535, A2 => n10938, ZN => n6762);
   U9522 : NOR2_X1 port map( A1 => n6696, A2 => n7583, ZN => n6763);
   U9524 : NAND2_X1 port map( A1 => n25601, A2 => n33947, ZN => n3058);
   U9526 : NAND2_X1 port map( A1 => n34576, A2 => n17594, ZN => n2721);
   U9533 : NOR2_X1 port map( A1 => n220, A2 => n2366, ZN => n3005);
   U9542 : NOR2_X1 port map( A1 => n37050, A2 => n1552, ZN => n8738);
   U9543 : OAI21_X1 port map( A1 => n19581, A2 => n12825, B => n20052, ZN => 
                           n10082);
   U9552 : NOR2_X1 port map( A1 => n5541, A2 => n31509, ZN => n5483);
   U9558 : NOR2_X1 port map( A1 => n14436, A2 => n835, ZN => n6573);
   U9576 : INV_X1 port map( I => n25552, ZN => n12828);
   U9582 : INV_X1 port map( I => n21031, ZN => n17183);
   U9586 : NAND2_X1 port map( A1 => n1560, A2 => n11601, ZN => n7263);
   U9589 : INV_X1 port map( I => n25218, ZN => n24873);
   U9590 : INV_X2 port map( I => n33132, ZN => n1258);
   U9598 : INV_X1 port map( I => n19670, ZN => n6598);
   U9602 : NOR2_X1 port map( A1 => n16745, A2 => n17270, ZN => n20000);
   U9606 : INV_X2 port map( I => n19691, ZN => n1261);
   U9610 : INV_X2 port map( I => n25140, ZN => n1262);
   U9616 : NOR2_X1 port map( A1 => n13583, A2 => n24806, ZN => n13582);
   U9620 : NAND2_X1 port map( A1 => n1567, A2 => n7831, ZN => n24491);
   U9622 : NAND2_X1 port map( A1 => n7248, A2 => n38073, ZN => n7245);
   U9631 : NAND2_X1 port map( A1 => n6273, A2 => n24529, ZN => n1784);
   U9633 : NAND2_X1 port map( A1 => n1583, A2 => n7177, ZN => n7176);
   U9635 : NAND2_X1 port map( A1 => n19484, A2 => n24680, ZN => n6335);
   U9642 : AOI21_X1 port map( A1 => n24692, A2 => n30764, B => n24717, ZN => 
                           n6539);
   U9643 : AOI21_X1 port map( A1 => n35250, A2 => n37395, B => n14211, ZN => 
                           n20505);
   U9647 : NAND2_X1 port map( A1 => n24785, A2 => n32045, ZN => n13817);
   U9658 : INV_X1 port map( I => n24613, ZN => n1567);
   U9659 : NOR2_X1 port map( A1 => n1583, A2 => n16238, ZN => n8803);
   U9663 : AOI21_X1 port map( A1 => n19431, A2 => n34458, B => n37341, ZN => 
                           n13553);
   U9664 : OAI21_X1 port map( A1 => n20155, A2 => n24712, B => n19279, ZN => 
                           n20154);
   U9670 : NOR2_X1 port map( A1 => n38749, A2 => n24515, ZN => n24776);
   U9673 : NOR2_X1 port map( A1 => n1030, A2 => n3697, ZN => n4176);
   U9677 : NAND2_X1 port map( A1 => n24707, A2 => n34526, ZN => n6274);
   U9678 : INV_X1 port map( I => n24866, ZN => n19339);
   U9683 : INV_X2 port map( I => n20728, ZN => n14999);
   U9684 : NAND2_X1 port map( A1 => n24148, A2 => n24274, ZN => n5360);
   U9687 : NAND2_X1 port map( A1 => n8846, A2 => n1598, ZN => n8845);
   U9712 : AOI21_X1 port map( A1 => n6998, A2 => n13692, B => n1595, ZN => 
                           n6997);
   U9719 : OAI21_X1 port map( A1 => n24272, A2 => n1604, B => n24273, ZN => 
                           n10713);
   U9721 : AOI21_X1 port map( A1 => n38224, A2 => n8690, B => n12692, ZN => 
                           n9362);
   U9731 : NAND2_X1 port map( A1 => n24231, A2 => n1127, ZN => n18256);
   U9737 : NOR2_X1 port map( A1 => n13808, A2 => n1598, ZN => n9634);
   U9751 : OAI21_X1 port map( A1 => n24406, A2 => n37934, B => n24410, ZN => 
                           n18615);
   U9762 : OAI22_X1 port map( A1 => n16884, A2 => n1596, B1 => n250, B2 => 
                           n24442, ZN => n10783);
   U9763 : NAND2_X1 port map( A1 => n39467, A2 => n19880, ZN => n9584);
   U9765 : NAND2_X1 port map( A1 => n19402, A2 => n6515, ZN => n9822);
   U9776 : NAND2_X1 port map( A1 => n4243, A2 => n36500, ZN => n3453);
   U9784 : NOR2_X1 port map( A1 => n18304, A2 => n7210, ZN => n24123);
   U9795 : NOR2_X1 port map( A1 => n24146, A2 => n232, ZN => n12692);
   U9797 : OR2_X1 port map( A1 => n13144, A2 => n30280, Z => n23855);
   U9799 : INV_X1 port map( I => n24445, ZN => n24448);
   U9807 : INV_X2 port map( I => n15865, ZN => n24469);
   U9813 : NAND2_X1 port map( A1 => n24294, A2 => n33939, ZN => n24297);
   U9826 : BUF_X2 port map( I => n24431, Z => n12975);
   U9832 : INV_X1 port map( I => n23794, ZN => n23670);
   U9839 : NAND2_X1 port map( A1 => n23751, A2 => n11452, ZN => n23987);
   U9846 : NOR2_X1 port map( A1 => n12638, A2 => n23399, ZN => n11723);
   U9857 : NAND2_X1 port map( A1 => n2961, A2 => n23588, ZN => n2960);
   U9865 : NOR2_X1 port map( A1 => n1918, A2 => n23622, ZN => n1917);
   U9866 : NOR2_X1 port map( A1 => n23251, A2 => n23592, ZN => n17888);
   U9868 : NOR2_X1 port map( A1 => n4207, A2 => n14235, ZN => n10840);
   U9880 : NAND2_X1 port map( A1 => n52, A2 => n33496, ZN => n15842);
   U9881 : NAND2_X1 port map( A1 => n23243, A2 => n38981, ZN => n12641);
   U9885 : INV_X1 port map( I => n11669, ZN => n4637);
   U9887 : NOR2_X1 port map( A1 => n32424, A2 => n1635, ZN => n6993);
   U9889 : OAI21_X1 port map( A1 => n32377, A2 => n23578, B => n1138, ZN => 
                           n10612);
   U9899 : INV_X1 port map( I => n23637, ZN => n23641);
   U9915 : NOR2_X1 port map( A1 => n16443, A2 => n35506, ZN => n9621);
   U9916 : NAND3_X1 port map( A1 => n37622, A2 => n38042, A3 => n23515, ZN => 
                           n11842);
   U9922 : NAND2_X1 port map( A1 => n4207, A2 => n14235, ZN => n10711);
   U9924 : NOR2_X1 port map( A1 => n23458, A2 => n23238, ZN => n4707);
   U9929 : NAND3_X1 port map( A1 => n6303, A2 => n6176, A3 => n23484, ZN => 
                           n23362);
   U9935 : NOR2_X1 port map( A1 => n20835, A2 => n16013, ZN => n13602);
   U9937 : INV_X1 port map( I => n38724, ZN => n19665);
   U9945 : OAI21_X1 port map( A1 => n36829, A2 => n30574, B => n37014, ZN => 
                           n9796);
   U9949 : INV_X1 port map( I => n23517, ZN => n6373);
   U9953 : NAND2_X1 port map( A1 => n7335, A2 => n23624, ZN => n3498);
   U9966 : NAND2_X1 port map( A1 => n6827, A2 => n6826, ZN => n11245);
   U9967 : OAI22_X1 port map( A1 => n2049, A2 => n1989, B1 => n20439, B2 => 
                           n23146, ZN => n23147);
   U9970 : INV_X1 port map( I => n3713, ZN => n3717);
   U9972 : NAND2_X1 port map( A1 => n6916, A2 => n20373, ZN => n4959);
   U9978 : AOI21_X1 port map( A1 => n6581, A2 => n4472, B => n15388, ZN => 
                           n6826);
   U9979 : NOR2_X1 port map( A1 => n19469, A2 => n8462, ZN => n8461);
   U9991 : NAND3_X1 port map( A1 => n17131, A2 => n22368, A3 => n1143, ZN => 
                           n6916);
   U10002 : AOI21_X1 port map( A1 => n11307, A2 => n23111, B => n12392, ZN => 
                           n13262);
   U10004 : OR3_X1 port map( A1 => n8809, A2 => n32677, A3 => n31300, Z => 
                           n22805);
   U10005 : AND2_X1 port map( A1 => n38524, A2 => n1647, Z => n2927);
   U10011 : AND3_X1 port map( A1 => n37791, A2 => n22368, A3 => n2047, Z => 
                           n5942);
   U10013 : NOR2_X1 port map( A1 => n1650, A2 => n6499, ZN => n6498);
   U10014 : NAND2_X1 port map( A1 => n1645, A2 => n14187, ZN => n14186);
   U10022 : NAND2_X1 port map( A1 => n23214, A2 => n4472, ZN => n3040);
   U10025 : NAND2_X1 port map( A1 => n22682, A2 => n22921, ZN => n13515);
   U10033 : NAND2_X1 port map( A1 => n272, A2 => n1655, ZN => n21062);
   U10034 : NOR2_X1 port map( A1 => n17080, A2 => n22920, ZN => n22922);
   U10038 : NAND2_X1 port map( A1 => n22890, A2 => n17080, ZN => n22924);
   U10046 : NOR2_X1 port map( A1 => n5657, A2 => n19645, ZN => n8458);
   U10050 : AND3_X1 port map( A1 => n33934, A2 => n19586, A3 => n33745, Z => 
                           n23187);
   U10051 : AND2_X1 port map( A1 => n18750, A2 => n3273, Z => n3543);
   U10058 : INV_X1 port map( I => n12925, ZN => n22901);
   U10060 : NOR2_X1 port map( A1 => n9472, A2 => n10074, ZN => n22860);
   U10062 : INV_X1 port map( I => n23088, ZN => n23090);
   U10066 : NAND2_X1 port map( A1 => n12392, A2 => n23108, ZN => n13339);
   U10068 : NOR2_X1 port map( A1 => n23111, A2 => n23110, ZN => n23112);
   U10069 : NOR2_X1 port map( A1 => n8197, A2 => n12630, ZN => n22908);
   U10076 : NOR2_X1 port map( A1 => n22709, A2 => n550, ZN => n5214);
   U10077 : NOR2_X1 port map( A1 => n18708, A2 => n1654, ZN => n4162);
   U10079 : NOR2_X1 port map( A1 => n3906, A2 => n23142, ZN => n2116);
   U10083 : NAND2_X1 port map( A1 => n1648, A2 => n16104, ZN => n20175);
   U10090 : CLKBUF_X2 port map( I => n22897, Z => n10074);
   U10107 : INV_X1 port map( I => n22862, ZN => n18708);
   U10114 : INV_X1 port map( I => n22610, ZN => n2838);
   U10115 : OAI21_X1 port map( A1 => n13565, A2 => n13566, B => n22348, ZN => 
                           n3024);
   U10117 : INV_X1 port map( I => n22622, ZN => n1657);
   U10118 : INV_X1 port map( I => n22657, ZN => n1660);
   U10129 : NAND2_X1 port map( A1 => n19515, A2 => n12023, ZN => n8343);
   U10131 : NAND2_X1 port map( A1 => n22055, A2 => n8089, ZN => n13765);
   U10137 : OAI21_X1 port map( A1 => n22143, A2 => n8754, B => n8753, ZN => 
                           n8752);
   U10153 : NAND2_X1 port map( A1 => n5053, A2 => n22286, ZN => n3954);
   U10154 : NOR2_X1 port map( A1 => n11542, A2 => n22388, ZN => n5204);
   U10156 : OAI21_X1 port map( A1 => n21958, A2 => n17531, B => n16989, ZN => 
                           n2386);
   U10160 : NAND2_X1 port map( A1 => n1672, A2 => n5617, ZN => n5616);
   U10161 : NAND2_X1 port map( A1 => n35822, A2 => n12793, ZN => n12812);
   U10165 : OAI22_X1 port map( A1 => n31092, A2 => n22324, B1 => n1812, B2 => 
                           n22323, ZN => n21830);
   U10171 : NAND2_X1 port map( A1 => n21090, A2 => n22326, ZN => n8342);
   U10179 : NAND2_X1 port map( A1 => n22181, A2 => n2840, ZN => n9843);
   U10181 : AOI21_X1 port map( A1 => n4239, A2 => n19873, B => n14423, ZN => 
                           n5207);
   U10183 : AND2_X1 port map( A1 => n11149, A2 => n19773, Z => n12023);
   U10188 : NAND2_X1 port map( A1 => n7955, A2 => n12230, ZN => n7818);
   U10193 : NOR2_X1 port map( A1 => n37217, A2 => n22132, ZN => n14311);
   U10194 : NAND2_X1 port map( A1 => n6128, A2 => n22295, ZN => n5497);
   U10198 : AND2_X1 port map( A1 => n22265, A2 => n19515, Z => n13900);
   U10210 : NAND2_X1 port map( A1 => n9387, A2 => n1688, ZN => n11013);
   U10211 : NAND2_X1 port map( A1 => n1686, A2 => n36371, ZN => n14020);
   U10212 : NAND2_X1 port map( A1 => n8520, A2 => n8518, ZN => n5053);
   U10218 : AOI21_X1 port map( A1 => n33168, A2 => n9422, B => n20376, ZN => 
                           n21363);
   U10219 : AND2_X1 port map( A1 => n1680, A2 => n6128, Z => n13627);
   U10222 : AND2_X1 port map( A1 => n22143, A2 => n37089, Z => n8687);
   U10238 : AOI21_X1 port map( A1 => n33860, A2 => n22177, B => n6451, ZN => 
                           n5878);
   U10241 : AND2_X1 port map( A1 => n35526, A2 => n22264, Z => n19211);
   U10256 : NAND2_X1 port map( A1 => n22226, A2 => n22225, ZN => n20123);
   U10261 : AND2_X1 port map( A1 => n19373, A2 => n9165, Z => n22249);
   U10264 : OAI21_X1 port map( A1 => n33168, A2 => n5821, B => n31649, ZN => 
                           n21364);
   U10272 : NAND2_X1 port map( A1 => n3325, A2 => n21583, ZN => n3323);
   U10278 : NAND2_X1 port map( A1 => n3676, A2 => n32817, ZN => n3680);
   U10280 : NOR2_X1 port map( A1 => n33168, A2 => n19017, ZN => n20374);
   U10289 : OAI22_X1 port map( A1 => n3692, A2 => n938, B1 => n1155, B2 => 
                           n5132, ZN => n3691);
   U10296 : AOI21_X1 port map( A1 => n8438, A2 => n21838, B => n1159, ZN => 
                           n8442);
   U10297 : NOR2_X1 port map( A1 => n10875, A2 => n37678, ZN => n10125);
   U10302 : INV_X2 port map( I => n8040, ZN => n1342);
   U10303 : NOR3_X1 port map( A1 => n38546, A2 => n21712, A3 => n17266, ZN => 
                           n17265);
   U10305 : AOI21_X1 port map( A1 => n21551, A2 => n19871, B => n21550, ZN => 
                           n11238);
   U10306 : AND2_X1 port map( A1 => n21654, A2 => n6732, Z => n12546);
   U10312 : AOI22_X1 port map( A1 => n8598, A2 => n19543, B1 => n17792, B2 => 
                           n8600, ZN => n15382);
   U10318 : AOI22_X1 port map( A1 => n8466, A2 => n19323, B1 => n8468, B2 => 
                           n670, ZN => n5417);
   U10319 : OAI21_X1 port map( A1 => n21911, A2 => n21910, B => n21909, ZN => 
                           n7608);
   U10322 : AOI21_X1 port map( A1 => n21665, A2 => n919, B => n21833, ZN => 
                           n9319);
   U10324 : NAND2_X1 port map( A1 => n21723, A2 => n1689, ZN => n4924);
   U10328 : AOI22_X1 port map( A1 => n1156, A2 => n21691, B1 => n21690, B2 => 
                           n21339, ZN => n7998);
   U10330 : NAND2_X1 port map( A1 => n13996, A2 => n13998, ZN => n12513);
   U10334 : NOR2_X1 port map( A1 => n21410, A2 => n21804, ZN => n21371);
   U10339 : INV_X1 port map( I => n21885, ZN => n2045);
   U10340 : OAI21_X1 port map( A1 => n18542, A2 => n17792, B => n21561, ZN => 
                           n21562);
   U10342 : INV_X1 port map( I => n20328, ZN => n21764);
   U10344 : AND2_X1 port map( A1 => n1159, A2 => n21897, Z => n11008);
   U10346 : AOI21_X1 port map( A1 => n17848, A2 => n21450, B => n17242, ZN => 
                           n17544);
   U10347 : NAND2_X1 port map( A1 => n21784, A2 => n37111, ZN => n18339);
   U10349 : NOR2_X1 port map( A1 => n19620, A2 => n8936, ZN => n8434);
   U10351 : OAI22_X1 port map( A1 => n293, A2 => n670, B1 => n18412, B2 => 
                           n34867, ZN => n13098);
   U10352 : OAI21_X1 port map( A1 => n7935, A2 => n21923, B => n4116, ZN => 
                           n5187);
   U10354 : AND2_X1 port map( A1 => n21565, A2 => n17534, Z => n3912);
   U10357 : NAND2_X1 port map( A1 => n1816, A2 => n15839, ZN => n13859);
   U10358 : NAND2_X1 port map( A1 => n1816, A2 => n15338, ZN => n13861);
   U10360 : NOR3_X1 port map( A1 => n917, A2 => n21928, A3 => n19372, ZN => 
                           n7640);
   U10362 : NAND2_X1 port map( A1 => n33771, A2 => n21762, ZN => n17886);
   U10364 : NAND2_X1 port map( A1 => n21640, A2 => n21923, ZN => n4925);
   U10367 : OAI21_X1 port map( A1 => n275, A2 => n21440, B => n16035, ZN => 
                           n21442);
   U10368 : NOR2_X1 port map( A1 => n21887, A2 => n19850, ZN => n5980);
   U10369 : NOR2_X1 port map( A1 => n21450, A2 => n1694, ZN => n16901);
   U10373 : AND2_X1 port map( A1 => n1694, A2 => n452, Z => n12439);
   U10375 : NAND2_X1 port map( A1 => n21899, A2 => n10120, ZN => n11007);
   U10379 : INV_X1 port map( I => n37200, ZN => n2277);
   U10390 : INV_X1 port map( I => n1697, ZN => n8951);
   U10392 : INV_X1 port map( I => n21688, ZN => n1693);
   U10395 : NAND2_X1 port map( A1 => n21893, A2 => n3294, ZN => n3295);
   U10396 : NOR2_X1 port map( A1 => n37200, A2 => n20266, ZN => n2187);
   U10397 : NAND2_X1 port map( A1 => n21730, A2 => n10211, ZN => n21554);
   U10400 : BUF_X2 port map( I => n21577, Z => n19238);
   U10401 : NOR2_X1 port map( A1 => n2533, A2 => n2532, ZN => n2531);
   U10403 : BUF_X2 port map( I => n21750, Z => n21889);
   U10404 : INV_X1 port map( I => n19733, ZN => n1734);
   U10405 : INV_X1 port map( I => n19874, ZN => n1695);
   U10408 : INV_X1 port map( I => n19616, ZN => n1710);
   U10410 : INV_X1 port map( I => n29785, ZN => n1711);
   U10415 : INV_X1 port map( I => n28831, ZN => n1723);
   U10421 : INV_X1 port map( I => n19527, ZN => n1707);
   U10422 : INV_X1 port map( I => n19722, ZN => n1714);
   U10424 : INV_X1 port map( I => n21428, ZN => n21682);
   U10425 : CLKBUF_X2 port map( I => n10212, Z => n9863);
   U10430 : INV_X1 port map( I => n19770, ZN => n1700);
   U10432 : INV_X1 port map( I => n29509, ZN => n1699);
   U10433 : INV_X1 port map( I => n29647, ZN => n1725);
   U10436 : INV_X1 port map( I => n29357, ZN => n1717);
   U10438 : CLKBUF_X2 port map( I => Key(174), Z => n29785);
   U10440 : CLKBUF_X2 port map( I => Key(188), Z => n29221);
   U10443 : CLKBUF_X2 port map( I => Key(38), Z => n29808);
   U10444 : CLKBUF_X2 port map( I => Key(90), Z => n29711);
   U10446 : CLKBUF_X2 port map( I => Key(104), Z => n30253);
   U10449 : CLKBUF_X2 port map( I => Key(26), Z => n29334);
   U10453 : CLKBUF_X2 port map( I => Key(191), Z => n29357);
   U10455 : CLKBUF_X2 port map( I => Key(182), Z => n30114);
   U10459 : CLKBUF_X2 port map( I => Key(144), Z => n19616);
   U10460 : CLKBUF_X2 port map( I => Key(116), Z => n29657);
   U10461 : CLKBUF_X2 port map( I => Key(158), Z => n19831);
   U10463 : CLKBUF_X2 port map( I => Key(125), Z => n30063);
   U10466 : CLKBUF_X2 port map( I => Key(135), Z => n29285);
   U10469 : CLKBUF_X2 port map( I => Key(55), Z => n19929);
   U10470 : CLKBUF_X2 port map( I => Key(48), Z => n30207);
   U10471 : CLKBUF_X2 port map( I => Key(149), Z => n29875);
   U10472 : CLKBUF_X2 port map( I => Key(179), Z => n30006);
   U10474 : CLKBUF_X2 port map( I => Key(117), Z => n29680);
   U10477 : CLKBUF_X2 port map( I => Key(23), Z => n19770);
   U10478 : CLKBUF_X2 port map( I => Key(68), Z => n29920);
   U10479 : CLKBUF_X2 port map( I => Key(185), Z => n30203);
   U10481 : CLKBUF_X2 port map( I => Key(119), Z => n28831);
   U10484 : CLKBUF_X2 port map( I => Key(136), Z => n19733);
   U10485 : CLKBUF_X2 port map( I => Key(122), Z => n28910);
   U10486 : CLKBUF_X2 port map( I => Key(56), Z => n29141);
   U10487 : CLKBUF_X2 port map( I => Key(2), Z => n29474);
   U10488 : CLKBUF_X2 port map( I => Key(77), Z => n19875);
   U10490 : CLKBUF_X2 port map( I => Key(29), Z => n29463);
   U10492 : CLKBUF_X2 port map( I => Key(105), Z => n29206);
   U10493 : NOR2_X1 port map( A1 => n5369, A2 => n30010, ZN => n5194);
   U10497 : NAND2_X1 port map( A1 => n12942, A2 => n29369, ZN => n29362);
   U10510 : NAND2_X1 port map( A1 => n6440, A2 => n29802, ZN => n6438);
   U10513 : AOI21_X1 port map( A1 => n14073, A2 => n29572, B => n14072, ZN => 
                           n29573);
   U10515 : AOI21_X1 port map( A1 => n12033, A2 => n5813, B => n5811, ZN => 
                           n15600);
   U10516 : AOI21_X1 port map( A1 => n29543, A2 => n29560, B => n21177, ZN => 
                           n29019);
   U10519 : OR2_X1 port map( A1 => n9591, A2 => n29932, Z => n16187);
   U10522 : NAND2_X1 port map( A1 => n9837, A2 => n19380, ZN => n29552);
   U10526 : NAND2_X1 port map( A1 => n7015, A2 => n5970, ZN => n6440);
   U10532 : AOI21_X1 port map( A1 => n3287, A2 => n29318, B => n3285, ZN => 
                           n3284);
   U10540 : AOI21_X1 port map( A1 => n29372, A2 => n29373, B => n29355, ZN => 
                           n15957);
   U10542 : NAND2_X1 port map( A1 => n18041, A2 => n31538, ZN => n3118);
   U10543 : NOR2_X1 port map( A1 => n6342, A2 => n29468, ZN => n6341);
   U10544 : OAI21_X1 port map( A1 => n19097, A2 => n29922, B => n8560, ZN => 
                           n18085);
   U10546 : AOI21_X1 port map( A1 => n29932, A2 => n29922, B => n1174, ZN => 
                           n29919);
   U10550 : OAI22_X1 port map( A1 => n30099, A2 => n30098, B1 => n30097, B2 => 
                           n6149, ZN => n6148);
   U10554 : OAI21_X1 port map( A1 => n14007, A2 => n4910, B => n29807, ZN => 
                           n29809);
   U10561 : NAND2_X1 port map( A1 => n6843, A2 => n16233, ZN => n11394);
   U10562 : NAND2_X1 port map( A1 => n29207, A2 => n920, ZN => n13143);
   U10565 : OAI22_X1 port map( A1 => n5580, A2 => n29860, B1 => n1171, B2 => 
                           n8727, ZN => n5065);
   U10567 : NAND2_X1 port map( A1 => n29923, A2 => n39709, ZN => n21283);
   U10571 : NOR2_X1 port map( A1 => n14009, A2 => n14008, ZN => n4910);
   U10574 : NAND2_X1 port map( A1 => n29540, A2 => n29541, ZN => n7435);
   U10575 : NAND2_X1 port map( A1 => n29846, A2 => n29851, ZN => n5108);
   U10579 : NOR2_X1 port map( A1 => n21146, A2 => n29739, ZN => n8064);
   U10580 : NAND2_X1 port map( A1 => n29275, A2 => n3378, ZN => n6842);
   U10581 : NAND2_X1 port map( A1 => n29795, A2 => n32050, ZN => n5467);
   U10582 : AOI21_X1 port map( A1 => n19090, A2 => n16233, B => n29277, ZN => 
                           n16232);
   U10589 : NAND2_X1 port map( A1 => n14414, A2 => n15841, ZN => n12340);
   U10590 : OAI21_X1 port map( A1 => n29437, A2 => n29441, B => n29433, ZN => 
                           n12339);
   U10591 : NAND2_X1 port map( A1 => n13363, A2 => n30257, ZN => n30247);
   U10592 : NOR3_X1 port map( A1 => n29677, A2 => n20672, A3 => n1173, ZN => 
                           n9610);
   U10597 : NAND2_X1 port map( A1 => n29670, A2 => n5067, ZN => n2110);
   U10598 : NAND2_X1 port map( A1 => n29979, A2 => n29980, ZN => n5018);
   U10600 : NOR2_X1 port map( A1 => n969, A2 => n29477, ZN => n9103);
   U10603 : INV_X1 port map( I => n15259, ZN => n11940);
   U10605 : NAND2_X1 port map( A1 => n12301, A2 => n30183, ZN => n10513);
   U10606 : AOI21_X1 port map( A1 => n2113, A2 => n29675, B => n2112, ZN => 
                           n2111);
   U10609 : INV_X2 port map( I => n7303, ZN => n13433);
   U10611 : AOI21_X1 port map( A1 => n19663, A2 => n1172, B => n11700, ZN => 
                           n13991);
   U10612 : NAND2_X1 port map( A1 => n8955, A2 => n13142, ZN => n13014);
   U10615 : NOR2_X1 port map( A1 => n2944, A2 => n2858, ZN => n2205);
   U10616 : AND2_X1 port map( A1 => n6720, A2 => n16803, Z => n11182);
   U10619 : INV_X1 port map( I => n3614, ZN => n3611);
   U10621 : AND2_X1 port map( A1 => n29806, A2 => n38141, Z => n14007);
   U10622 : NAND2_X1 port map( A1 => n29858, A2 => n3725, ZN => n2945);
   U10626 : OAI21_X1 port map( A1 => n29439, A2 => n15841, B => n18502, ZN => 
                           n15131);
   U10630 : NAND2_X1 port map( A1 => n17192, A2 => n17469, ZN => n9264);
   U10631 : OR2_X1 port map( A1 => n8287, A2 => n20274, Z => n10289);
   U10632 : INV_X1 port map( I => n8063, ZN => n8062);
   U10633 : INV_X1 port map( I => n36096, ZN => n29791);
   U10635 : INV_X1 port map( I => n30033, ZN => n18780);
   U10636 : AND4_X1 port map( A1 => n29273, A2 => n29272, A3 => n29270, A4 => 
                           n29271, Z => n29274);
   U10641 : OR2_X1 port map( A1 => n29407, A2 => n9790, Z => n20131);
   U10642 : NAND2_X1 port map( A1 => n16683, A2 => n9839, ZN => n7376);
   U10643 : AOI21_X1 port map( A1 => n31539, A2 => n29683, B => n18042, ZN => 
                           n29674);
   U10648 : AND4_X1 port map( A1 => n30174, A2 => n10101, A3 => n30173, A4 => 
                           n30172, Z => n30175);
   U10654 : OR2_X1 port map( A1 => n17262, A2 => n29574, Z => n29572);
   U10667 : CLKBUF_X2 port map( I => n29687, Z => n5067);
   U10670 : INV_X1 port map( I => n29687, ZN => n29676);
   U10684 : NAND2_X1 port map( A1 => n9573, A2 => n29957, ZN => n9570);
   U10690 : NAND2_X1 port map( A1 => n20436, A2 => n20435, ZN => n20434);
   U10698 : OAI22_X1 port map( A1 => n29499, A2 => n36275, B1 => n29498, B2 => 
                           n29497, ZN => n29503);
   U10700 : NAND2_X1 port map( A1 => n5300, A2 => n33784, ZN => n5299);
   U10706 : INV_X1 port map( I => n9885, ZN => n9884);
   U10707 : INV_X1 port map( I => n4220, ZN => n9818);
   U10712 : OAI21_X1 port map( A1 => n16116, A2 => n1179, B => n4655, ZN => 
                           n29496);
   U10722 : NAND2_X1 port map( A1 => n37544, A2 => n15584, ZN => n15583);
   U10728 : NAND2_X1 port map( A1 => n18658, A2 => n19994, ZN => n6257);
   U10731 : INV_X1 port map( I => n14281, ZN => n12657);
   U10733 : AOI21_X1 port map( A1 => n39830, A2 => n21023, B => n344, ZN => 
                           n20435);
   U10736 : NOR2_X1 port map( A1 => n15267, A2 => n7194, ZN => n7191);
   U10741 : NOR2_X1 port map( A1 => n30152, A2 => n33784, ZN => n10976);
   U10743 : NAND2_X1 port map( A1 => n29702, A2 => n9000, ZN => n8999);
   U10746 : OAI21_X1 port map( A1 => n7790, A2 => n30240, B => n31603, ZN => 
                           n8338);
   U10748 : INV_X1 port map( I => n13069, ZN => n11218);
   U10752 : NOR2_X1 port map( A1 => n2001, A2 => n19878, ZN => n9572);
   U10755 : OAI21_X1 port map( A1 => n2001, A2 => n29960, B => n29955, ZN => 
                           n9573);
   U10762 : INV_X1 port map( I => n7166, ZN => n7163);
   U10765 : NAND2_X1 port map( A1 => n34086, A2 => n7167, ZN => n7164);
   U10769 : NAND2_X1 port map( A1 => n13657, A2 => n12992, ZN => n12991);
   U10770 : NAND2_X1 port map( A1 => n13942, A2 => n16116, ZN => n7614);
   U10774 : NAND2_X1 port map( A1 => n8477, A2 => n29997, ZN => n8419);
   U10775 : NAND2_X1 port map( A1 => n7448, A2 => n29779, ZN => n21038);
   U10780 : NOR2_X1 port map( A1 => n30153, A2 => n1059, ZN => n8716);
   U10784 : NOR2_X1 port map( A1 => n21168, A2 => n21167, ZN => n21166);
   U10788 : OR2_X1 port map( A1 => n6851, A2 => n8918, Z => n10452);
   U10792 : NOR2_X1 port map( A1 => n8529, A2 => n30049, ZN => n29864);
   U10794 : OR2_X1 port map( A1 => n29643, A2 => n19734, Z => n29485);
   U10796 : NAND2_X1 port map( A1 => n14151, A2 => n29494, ZN => n28902);
   U10800 : OAI21_X1 port map( A1 => n34006, A2 => n20979, B => n19962, ZN => 
                           n28885);
   U10806 : NAND2_X1 port map( A1 => n1059, A2 => n30192, ZN => n8031);
   U10807 : OAI21_X1 port map( A1 => n29006, A2 => n1058, B => n29992, ZN => 
                           n13069);
   U10809 : NOR2_X1 port map( A1 => n3700, A2 => n5471, ZN => n3246);
   U10813 : AND2_X1 port map( A1 => n19508, A2 => n3700, Z => n29703);
   U10816 : CLKBUF_X2 port map( I => n37083, Z => n10101);
   U10826 : NAND2_X1 port map( A1 => n9872, A2 => n10590, ZN => n7193);
   U10829 : AND2_X1 port map( A1 => n29701, A2 => n5977, Z => n14511);
   U10833 : NOR2_X1 port map( A1 => n16490, A2 => n29940, ZN => n7363);
   U10834 : INV_X1 port map( I => n11677, ZN => n9836);
   U10836 : NOR2_X1 port map( A1 => n10702, A2 => n7789, ZN => n8892);
   U10845 : INV_X1 port map( I => n9649, ZN => n2001);
   U10846 : OR2_X1 port map( A1 => n29450, A2 => n28899, Z => n29380);
   U10847 : INV_X1 port map( I => n29904, ZN => n29902);
   U10849 : AND2_X1 port map( A1 => n10569, A2 => n6938, Z => n28788);
   U10852 : AND2_X1 port map( A1 => n16224, A2 => n16060, Z => n15521);
   U10853 : NOR3_X1 port map( A1 => n14449, A2 => n29310, A3 => n1406, ZN => 
                           n29078);
   U10863 : INV_X1 port map( I => n15293, ZN => n18461);
   U10865 : INV_X1 port map( I => n35551, ZN => n11826);
   U10866 : NOR2_X1 port map( A1 => n15293, A2 => n20018, ZN => n12056);
   U10867 : INV_X2 port map( I => n34175, ZN => n29635);
   U10868 : INV_X1 port map( I => n14438, ZN => n7295);
   U10870 : NAND2_X1 port map( A1 => n20931, A2 => n3986, ZN => n3951);
   U10872 : INV_X1 port map( I => n30058, ZN => n3671);
   U10873 : INV_X1 port map( I => n20508, ZN => n13349);
   U10874 : AND2_X1 port map( A1 => n30042, A2 => n30041, Z => n29150);
   U10875 : AND2_X1 port map( A1 => n2216, A2 => n29957, Z => n11830);
   U10876 : OR2_X1 port map( A1 => n39828, A2 => n20102, Z => n29173);
   U10877 : NOR2_X1 port map( A1 => n28882, A2 => n21023, ZN => n17681);
   U10878 : NOR2_X1 port map( A1 => n971, A2 => n39745, ZN => n9049);
   U10882 : OR2_X1 port map( A1 => n30047, A2 => n16217, Z => n14664);
   U10883 : INV_X1 port map( I => n29347, ZN => n14178);
   U10884 : AND2_X1 port map( A1 => n15651, A2 => n5414, Z => n18962);
   U10886 : CLKBUF_X2 port map( I => n29907, Z => n19878);
   U10887 : INV_X4 port map( I => n29185, ZN => n1400);
   U10894 : NOR2_X1 port map( A1 => n21187, A2 => n29862, ZN => n2216);
   U10897 : INV_X2 port map( I => n19599, ZN => n29760);
   U10902 : CLKBUF_X2 port map( I => n14405, Z => n12353);
   U10915 : INV_X1 port map( I => n29049, ZN => n12574);
   U10917 : INV_X1 port map( I => n29153, ZN => n5041);
   U10918 : INV_X1 port map( I => n29114, ZN => n9436);
   U10921 : NAND2_X1 port map( A1 => n15006, A2 => n15005, ZN => n3551);
   U10922 : INV_X1 port map( I => n29026, ZN => n2914);
   U10924 : INV_X1 port map( I => n38147, ZN => n6854);
   U10925 : INV_X1 port map( I => n29162, ZN => n2995);
   U10927 : NAND2_X1 port map( A1 => n7384, A2 => n28747, ZN => n28751);
   U10928 : NAND2_X1 port map( A1 => n19957, A2 => n7296, ZN => n13484);
   U10936 : INV_X1 port map( I => n15271, ZN => n11347);
   U10944 : INV_X1 port map( I => n28852, ZN => n28707);
   U10946 : INV_X1 port map( I => n28529, ZN => n28343);
   U10955 : NAND2_X1 port map( A1 => n28522, A2 => n28747, ZN => n12608);
   U10961 : NAND2_X1 port map( A1 => n18473, A2 => n18470, ZN => n28953);
   U10968 : AOI21_X1 port map( A1 => n20314, A2 => n28331, B => n29474, ZN => 
                           n15007);
   U10972 : NAND2_X1 port map( A1 => n28480, A2 => n32575, ZN => n4665);
   U10976 : AND2_X1 port map( A1 => n6405, A2 => n3927, Z => n8323);
   U10980 : INV_X1 port map( I => n1815, ZN => n4371);
   U11003 : OR2_X1 port map( A1 => n28095, A2 => n19827, Z => n14049);
   U11006 : INV_X1 port map( I => n28747, ZN => n4025);
   U11026 : NAND2_X1 port map( A1 => n20952, A2 => n28748, ZN => n20951);
   U11032 : AND2_X1 port map( A1 => n6287, A2 => n37204, Z => n12882);
   U11033 : NOR2_X1 port map( A1 => n28289, A2 => n1187, ZN => n13963);
   U11035 : INV_X1 port map( I => n28455, ZN => n12883);
   U11041 : OR3_X1 port map( A1 => n28720, A2 => n28722, A3 => n38145, Z => 
                           n13593);
   U11044 : INV_X1 port map( I => n28431, ZN => n16307);
   U11057 : AND2_X1 port map( A1 => n28612, A2 => n7454, Z => n2060);
   U11060 : AND2_X1 port map( A1 => n6892, A2 => n12237, Z => n12238);
   U11065 : AND2_X1 port map( A1 => n9878, A2 => n32146, Z => n28528);
   U11067 : NOR2_X1 port map( A1 => n10544, A2 => n10543, ZN => n13563);
   U11069 : INV_X1 port map( I => n28576, ZN => n2703);
   U11077 : NOR2_X1 port map( A1 => n39355, A2 => n28464, ZN => n28302);
   U11081 : INV_X1 port map( I => n28535, ZN => n7869);
   U11082 : INV_X1 port map( I => n15752, ZN => n5399);
   U11092 : NOR2_X1 port map( A1 => n1190, A2 => n30894, ZN => n17542);
   U11095 : NAND2_X1 port map( A1 => n13508, A2 => n28408, ZN => n20878);
   U11099 : AND2_X1 port map( A1 => n28551, A2 => n28659, Z => n14652);
   U11100 : AND2_X1 port map( A1 => n10907, A2 => n18871, Z => n10857);
   U11102 : NAND2_X1 port map( A1 => n3903, A2 => n28569, ZN => n28571);
   U11105 : OR2_X1 port map( A1 => n28606, A2 => n8349, Z => n12045);
   U11106 : NOR2_X1 port map( A1 => n28391, A2 => n28486, ZN => n12343);
   U11107 : NAND2_X1 port map( A1 => n28313, A2 => n19844, ZN => n28209);
   U11110 : AND2_X1 port map( A1 => n28532, A2 => n36796, Z => n13894);
   U11113 : AND2_X1 port map( A1 => n28759, A2 => n2022, Z => n13237);
   U11114 : NOR2_X1 port map( A1 => n7251, A2 => n31554, ZN => n5343);
   U11118 : INV_X1 port map( I => n28515, ZN => n9638);
   U11120 : INV_X1 port map( I => n1193, ZN => n5152);
   U11124 : AND2_X1 port map( A1 => n28433, A2 => n28434, Z => n8322);
   U11126 : AND2_X1 port map( A1 => n28681, A2 => n15473, Z => n14677);
   U11128 : INV_X1 port map( I => n13601, ZN => n6017);
   U11129 : OAI21_X1 port map( A1 => n38998, A2 => n36623, B => n5028, ZN => 
                           n3191);
   U11130 : NOR2_X1 port map( A1 => n28606, A2 => n2639, ZN => n10757);
   U11134 : NOR2_X1 port map( A1 => n20199, A2 => n20198, ZN => n20197);
   U11136 : NAND2_X1 port map( A1 => n13133, A2 => n496, ZN => n8714);
   U11140 : OR2_X1 port map( A1 => n8349, A2 => n36827, Z => n14339);
   U11141 : AND2_X1 port map( A1 => n18369, A2 => n28717, Z => n4428);
   U11144 : AND2_X1 port map( A1 => n28772, A2 => n17771, Z => n28773);
   U11147 : NOR2_X1 port map( A1 => n31597, A2 => n14760, ZN => n28635);
   U11151 : INV_X1 port map( I => n28444, ZN => n14003);
   U11153 : INV_X1 port map( I => n1192, ZN => n11128);
   U11156 : NAND3_X1 port map( A1 => n28424, A2 => n17818, A3 => n28423, ZN => 
                           n9405);
   U11165 : OAI21_X1 port map( A1 => n1206, A2 => n3231, B => n3230, ZN => 
                           n4028);
   U11178 : NOR2_X1 port map( A1 => n18020, A2 => n17447, ZN => n17057);
   U11195 : NAND2_X1 port map( A1 => n11743, A2 => n37623, ZN => n11742);
   U11200 : AND4_X1 port map( A1 => n28347, A2 => n28346, A3 => n28345, A4 => 
                           n28344, Z => n28348);
   U11204 : AND3_X1 port map( A1 => n20019, A2 => n20020, A3 => n28104, Z => 
                           n14596);
   U11205 : INV_X1 port map( I => n11717, ZN => n12061);
   U11208 : INV_X1 port map( I => n10167, ZN => n3534);
   U11216 : NAND2_X1 port map( A1 => n1198, A2 => n27892, ZN => n13755);
   U11223 : NAND2_X1 port map( A1 => n28053, A2 => n18392, ZN => n13847);
   U11235 : NAND2_X1 port map( A1 => n8290, A2 => n1073, ZN => n8289);
   U11243 : NAND2_X1 port map( A1 => n1445, A2 => n981, ZN => n17856);
   U11245 : INV_X1 port map( I => n8819, ZN => n28243);
   U11252 : NAND2_X1 port map( A1 => n28022, A2 => n27951, ZN => n11705);
   U11257 : NAND2_X1 port map( A1 => n27948, A2 => n28022, ZN => n19039);
   U11259 : NAND2_X1 port map( A1 => n11024, A2 => n28260, ZN => n10150);
   U11260 : OAI21_X1 port map( A1 => n7719, A2 => n984, B => n7718, ZN => 
                           n28058);
   U11262 : OAI21_X1 port map( A1 => n4767, A2 => n14389, B => n4766, ZN => 
                           n28185);
   U11268 : NAND2_X1 port map( A1 => n18530, A2 => n19743, ZN => n18529);
   U11272 : NOR2_X1 port map( A1 => n27963, A2 => n14404, ZN => n21318);
   U11276 : NAND2_X1 port map( A1 => n28259, A2 => n28258, ZN => n9990);
   U11277 : NOR2_X1 port map( A1 => n16115, A2 => n580, ZN => n6693);
   U11278 : NAND2_X1 port map( A1 => n5939, A2 => n28045, ZN => n4889);
   U11293 : INV_X1 port map( I => n13984, ZN => n10536);
   U11296 : AND2_X1 port map( A1 => n1202, A2 => n16115, Z => n6245);
   U11299 : OAI21_X1 port map( A1 => n8801, A2 => n18061, B => n27998, ZN => 
                           n4788);
   U11307 : INV_X1 port map( I => n6777, ZN => n3198);
   U11311 : INV_X1 port map( I => n28223, ZN => n28227);
   U11312 : INV_X1 port map( I => n15695, ZN => n15693);
   U11313 : NAND2_X1 port map( A1 => n8291, A2 => n17032, ZN => n8290);
   U11314 : AOI21_X1 port map( A1 => n33980, A2 => n13457, B => n36844, ZN => 
                           n3067);
   U11316 : OAI21_X1 port map( A1 => n16461, A2 => n878, B => n4507, ZN => 
                           n4506);
   U11319 : NOR2_X1 port map( A1 => n33957, A2 => n28283, ZN => n13993);
   U11330 : INV_X1 port map( I => n28235, ZN => n3832);
   U11335 : INV_X1 port map( I => n28285, ZN => n6374);
   U11341 : OR2_X1 port map( A1 => n1211, A2 => n28089, Z => n6118);
   U11351 : NAND2_X1 port map( A1 => n2302, A2 => n17314, ZN => n27888);
   U11353 : OR2_X1 port map( A1 => n1209, A2 => n882, Z => n27911);
   U11354 : INV_X1 port map( I => n11408, ZN => n8351);
   U11359 : AND3_X1 port map( A1 => n33656, A2 => n37783, A3 => n288, Z => 
                           n6115);
   U11361 : OAI21_X1 port map( A1 => n27772, A2 => n36877, B => n30846, ZN => 
                           n10825);
   U11363 : NOR2_X1 port map( A1 => n5940, A2 => n6990, ZN => n5939);
   U11369 : OR2_X1 port map( A1 => n18841, A2 => n16065, Z => n4825);
   U11371 : NAND2_X1 port map( A1 => n28257, A2 => n3989, ZN => n3164);
   U11375 : NAND2_X1 port map( A1 => n12623, A2 => n28238, ZN => n2983);
   U11386 : AND2_X1 port map( A1 => n759, A2 => n28205, Z => n14791);
   U11391 : INV_X1 port map( I => n27901, ZN => n4507);
   U11394 : INV_X1 port map( I => n28282, ZN => n12807);
   U11396 : INV_X1 port map( I => n10009, ZN => n14829);
   U11400 : INV_X2 port map( I => n12298, ZN => n27910);
   U11405 : OR2_X1 port map( A1 => n27995, A2 => n16461, Z => n4502);
   U11406 : OR2_X1 port map( A1 => n5266, A2 => n20053, Z => n20993);
   U11409 : AND2_X1 port map( A1 => n19667, A2 => n28137, Z => n16987);
   U11411 : NOR2_X1 port map( A1 => n36854, A2 => n11283, ZN => n2613);
   U11412 : INV_X1 port map( I => n12663, ZN => n19525);
   U11413 : BUF_X2 port map( I => n19855, Z => n6643);
   U11414 : NAND2_X1 port map( A1 => n39488, A2 => n28237, ZN => n2982);
   U11417 : NOR2_X1 port map( A1 => n16115, A2 => n39571, ZN => n15048);
   U11418 : INV_X2 port map( I => n17177, ZN => n1445);
   U11419 : INV_X1 port map( I => n28127, ZN => n28124);
   U11424 : INV_X2 port map( I => n9791, ZN => n15925);
   U11425 : CLKBUF_X2 port map( I => n28132, Z => n19946);
   U11428 : BUF_X2 port map( I => n28127, Z => n11891);
   U11429 : INV_X4 port map( I => n28236, ZN => n1453);
   U11430 : INV_X1 port map( I => n27675, ZN => n6471);
   U11432 : INV_X1 port map( I => n14977, ZN => n3499);
   U11433 : INV_X1 port map( I => n27732, ZN => n27733);
   U11441 : OAI21_X1 port map( A1 => n13291, A2 => n13290, B => n27523, ZN => 
                           n12240);
   U11451 : INV_X1 port map( I => n13293, ZN => n13290);
   U11453 : NAND2_X2 port map( A1 => n12415, A2 => n26967, ZN => n12556);
   U11455 : NAND2_X1 port map( A1 => n27466, A2 => n19877, ZN => n17686);
   U11459 : AND2_X1 port map( A1 => n27346, A2 => n27345, Z => n6689);
   U11463 : NOR2_X1 port map( A1 => n10576, A2 => n10575, ZN => n10573);
   U11471 : OAI21_X1 port map( A1 => n17524, A2 => n21110, B => n17523, ZN => 
                           n4419);
   U11476 : INV_X1 port map( I => n26942, ZN => n10575);
   U11477 : INV_X1 port map( I => n13245, ZN => n27597);
   U11481 : INV_X1 port map( I => n27178, ZN => n27860);
   U11482 : INV_X1 port map( I => n10580, ZN => n10576);
   U11487 : INV_X1 port map( I => n27549, ZN => n27863);
   U11489 : NAND2_X1 port map( A1 => n27199, A2 => n35919, ZN => n9202);
   U11493 : AND3_X1 port map( A1 => n27563, A2 => n27562, A3 => n27561, Z => 
                           n18927);
   U11497 : INV_X1 port map( I => n27501, ZN => n7910);
   U11499 : INV_X1 port map( I => n27632, ZN => n12970);
   U11501 : INV_X1 port map( I => n27509, ZN => n15245);
   U11502 : INV_X2 port map( I => n27541, ZN => n1466);
   U11505 : INV_X2 port map( I => n27755, ZN => n1467);
   U11508 : NAND2_X1 port map( A1 => n30981, A2 => n27368, ZN => n13462);
   U11514 : NAND2_X1 port map( A1 => n27351, A2 => n11682, ZN => n8168);
   U11516 : INV_X1 port map( I => n10177, ZN => n10176);
   U11517 : NAND2_X1 port map( A1 => n27559, A2 => n8252, ZN => n27563);
   U11531 : NAND3_X1 port map( A1 => n20143, A2 => n20145, A3 => n27288, ZN => 
                           n12446);
   U11534 : NAND2_X1 port map( A1 => n8931, A2 => n36159, ZN => n7312);
   U11536 : NAND2_X1 port map( A1 => n27351, A2 => n8988, ZN => n27051);
   U11540 : AND3_X1 port map( A1 => n27428, A2 => n4964, A3 => n10461, Z => 
                           n9452);
   U11557 : NAND2_X1 port map( A1 => n27366, A2 => n9310, ZN => n5774);
   U11563 : OR3_X1 port map( A1 => n39711, A2 => n35904, A3 => n1084, Z => 
                           n14116);
   U11566 : NOR2_X1 port map( A1 => n5101, A2 => n6534, ZN => n7894);
   U11578 : NOR2_X1 port map( A1 => n2259, A2 => n5559, ZN => n2258);
   U11579 : OAI21_X1 port map( A1 => n38305, A2 => n27197, B => n19455, ZN => 
                           n16127);
   U11580 : NAND3_X1 port map( A1 => n27412, A2 => n36200, A3 => n997, ZN => 
                           n20203);
   U11588 : OR2_X1 port map( A1 => n18562, A2 => n12018, Z => n12017);
   U11597 : NAND2_X1 port map( A1 => n27430, A2 => n10051, ZN => n10755);
   U11616 : NAND2_X1 port map( A1 => n9512, A2 => n27009, ZN => n10574);
   U11621 : NAND2_X1 port map( A1 => n27220, A2 => n39546, ZN => n6192);
   U11627 : OR2_X1 port map( A1 => n27289, A2 => n1223, Z => n14682);
   U11628 : NAND2_X1 port map( A1 => n27020, A2 => n11140, ZN => n16919);
   U11633 : NAND2_X1 port map( A1 => n1080, A2 => n17662, ZN => n17465);
   U11636 : NOR2_X1 port map( A1 => n27248, A2 => n6972, ZN => n11853);
   U11637 : NAND2_X1 port map( A1 => n991, A2 => n3531, ZN => n8932);
   U11643 : NAND2_X1 port map( A1 => n26428, A2 => n35299, ZN => n9680);
   U11652 : NAND2_X1 port map( A1 => n994, A2 => n35258, ZN => n1798);
   U11654 : AND2_X1 port map( A1 => n27484, A2 => n1218, Z => n11042);
   U11658 : NAND2_X1 port map( A1 => n18549, A2 => n34562, ZN => n12018);
   U11664 : NAND2_X1 port map( A1 => n11039, A2 => n39296, ZN => n7227);
   U11665 : AND2_X1 port map( A1 => n27387, A2 => n6908, Z => n20870);
   U11669 : NAND2_X1 port map( A1 => n18669, A2 => n14881, ZN => n18668);
   U11674 : AND2_X1 port map( A1 => n27385, A2 => n34562, Z => n5219);
   U11682 : AND2_X1 port map( A1 => n39671, A2 => n20740, Z => n14482);
   U11693 : NAND2_X1 port map( A1 => n27298, A2 => n8137, ZN => n4038);
   U11696 : INV_X1 port map( I => n5630, ZN => n2006);
   U11700 : INV_X1 port map( I => n27128, ZN => n6416);
   U11702 : NOR2_X1 port map( A1 => n31672, A2 => n27269, ZN => n3466);
   U11706 : NAND2_X1 port map( A1 => n27383, A2 => n27064, ZN => n12022);
   U11720 : NOR2_X1 port map( A1 => n12685, A2 => n27417, ZN => n7175);
   U11722 : INV_X1 port map( I => n20871, ZN => n2846);
   U11723 : AOI21_X1 port map( A1 => n31672, A2 => n27267, B => n27372, ZN => 
                           n15748);
   U11739 : NAND2_X1 port map( A1 => n26612, A2 => n14496, ZN => n17467);
   U11740 : NAND2_X1 port map( A1 => n26037, A2 => n10890, ZN => n12510);
   U11742 : NAND2_X1 port map( A1 => n20797, A2 => n10187, ZN => n7912);
   U11743 : INV_X2 port map( I => n9144, ZN => n26870);
   U11762 : NAND2_X1 port map( A1 => n38120, A2 => n26515, ZN => n4489);
   U11780 : NAND2_X1 port map( A1 => n20462, A2 => n21202, ZN => n10203);
   U11784 : INV_X1 port map( I => n8311, ZN => n26684);
   U11792 : NAND2_X1 port map( A1 => n26731, A2 => n17712, ZN => n9075);
   U11817 : NAND2_X1 port map( A1 => n26697, A2 => n26269, ZN => n4937);
   U11824 : OR2_X1 port map( A1 => n7742, A2 => n4218, Z => n20912);
   U11825 : NOR2_X1 port map( A1 => n14825, A2 => n17047, ZN => n13159);
   U11833 : NOR2_X1 port map( A1 => n3368, A2 => n1229, ZN => n20549);
   U11836 : OR2_X1 port map( A1 => n16773, A2 => n3388, Z => n26138);
   U11838 : NAND2_X1 port map( A1 => n4486, A2 => n11334, ZN => n4485);
   U11840 : NAND2_X1 port map( A1 => n26926, A2 => n26470, ZN => n6503);
   U11843 : NAND2_X1 port map( A1 => n26283, A2 => n19353, ZN => n13252);
   U11846 : NAND2_X1 port map( A1 => n14382, A2 => n860, ZN => n8746);
   U11848 : NOR2_X1 port map( A1 => n26299, A2 => n26763, ZN => n7320);
   U11856 : NAND2_X1 port map( A1 => n17655, A2 => n13110, ZN => n17823);
   U11857 : NAND2_X1 port map( A1 => n17466, A2 => n36392, ZN => n11388);
   U11859 : NOR2_X1 port map( A1 => n15124, A2 => n13181, ZN => n4173);
   U11864 : NAND2_X1 port map( A1 => n19206, A2 => n19425, ZN => n26717);
   U11866 : INV_X2 port map( I => n19762, ZN => n26826);
   U11868 : OAI21_X1 port map( A1 => n26842, A2 => n34004, B => n9650, ZN => 
                           n21181);
   U11871 : OR2_X1 port map( A1 => n26671, A2 => n26672, Z => n14583);
   U11879 : NAND2_X1 port map( A1 => n26734, A2 => n9188, ZN => n9763);
   U11880 : NAND2_X1 port map( A1 => n10913, A2 => n26978, ZN => n5438);
   U11883 : INV_X1 port map( I => n18792, ZN => n4887);
   U11886 : AND2_X1 port map( A1 => n26686, A2 => n26979, Z => n17098);
   U11894 : NOR2_X1 port map( A1 => n26819, A2 => n37104, ZN => n13948);
   U11898 : NOR2_X1 port map( A1 => n13110, A2 => n26993, ZN => n4656);
   U11899 : NOR2_X1 port map( A1 => n38491, A2 => n19332, ZN => n18706);
   U11914 : OR2_X1 port map( A1 => n33726, A2 => n3328, Z => n26813);
   U11915 : NAND2_X1 port map( A1 => n5869, A2 => n26932, ZN => n16633);
   U11923 : AND2_X1 port map( A1 => n13758, A2 => n3134, Z => n3135);
   U11924 : NOR2_X1 port map( A1 => n3574, A2 => n1008, ZN => n3573);
   U11925 : OAI22_X1 port map( A1 => n26979, A2 => n26978, B1 => n17097, B2 => 
                           n17252, ZN => n26981);
   U11929 : OR3_X1 port map( A1 => n26901, A2 => n10231, A3 => n19821, Z => 
                           n26902);
   U11931 : NOR2_X1 port map( A1 => n26930, A2 => n19222, ZN => n7523);
   U11932 : INV_X1 port map( I => n14347, ZN => n16970);
   U11935 : INV_X1 port map( I => n26926, ZN => n26928);
   U11938 : NOR2_X1 port map( A1 => n1232, A2 => n19371, ZN => n8989);
   U11939 : NOR2_X1 port map( A1 => n2966, A2 => n19338, ZN => n2965);
   U11940 : INV_X1 port map( I => n13777, ZN => n4486);
   U11941 : INV_X1 port map( I => n33561, ZN => n19045);
   U11944 : OR2_X1 port map( A1 => n26724, A2 => n14355, Z => n26725);
   U11956 : AND2_X1 port map( A1 => n6190, A2 => n10440, Z => n8010);
   U11960 : NOR2_X1 port map( A1 => n26708, A2 => n17034, ZN => n4946);
   U11974 : INV_X1 port map( I => n13131, ZN => n26346);
   U11975 : INV_X1 port map( I => n26309, ZN => n13928);
   U11977 : INV_X1 port map( I => n34009, ZN => n19882);
   U11979 : INV_X1 port map( I => n26348, ZN => n7474);
   U11986 : INV_X1 port map( I => n26154, ZN => n7571);
   U11987 : INV_X1 port map( I => n26201, ZN => n3802);
   U11991 : INV_X1 port map( I => n9001, ZN => n6413);
   U11993 : INV_X1 port map( I => n26434, ZN => n3639);
   U12000 : INV_X1 port map( I => n3219, ZN => n3218);
   U12002 : INV_X1 port map( I => n17757, ZN => n26291);
   U12007 : NAND2_X1 port map( A1 => n14546, A2 => n26333, ZN => n12859);
   U12010 : INV_X1 port map( I => n7481, ZN => n2178);
   U12013 : INV_X1 port map( I => n5241, ZN => n5691);
   U12017 : INV_X1 port map( I => n36522, ZN => n26550);
   U12019 : INV_X1 port map( I => n26514, ZN => n12915);
   U12033 : OR2_X1 port map( A1 => n10724, A2 => n25989, Z => n20336);
   U12039 : NAND2_X1 port map( A1 => n4293, A2 => n37502, ZN => n4292);
   U12041 : NOR2_X1 port map( A1 => n33440, A2 => n26001, ZN => n9375);
   U12048 : OAI21_X1 port map( A1 => n424, A2 => n927, B => n5162, ZN => n5161)
                           ;
   U12052 : NAND2_X1 port map( A1 => n18958, A2 => n7544, ZN => n12490);
   U12060 : NAND2_X1 port map( A1 => n8710, A2 => n26027, ZN => n8709);
   U12061 : NOR2_X1 port map( A1 => n26214, A2 => n5908, ZN => n17125);
   U12062 : NAND2_X1 port map( A1 => n25958, A2 => n25959, ZN => n2125);
   U12070 : INV_X1 port map( I => n14157, ZN => n26238);
   U12071 : AND2_X1 port map( A1 => n26187, A2 => n14375, Z => n16878);
   U12073 : INV_X1 port map( I => n26190, ZN => n3333);
   U12077 : NAND2_X1 port map( A1 => n17035, A2 => n25970, ZN => n9811);
   U12078 : AND2_X1 port map( A1 => n25770, A2 => n25941, Z => n14685);
   U12084 : NAND2_X1 port map( A1 => n8898, A2 => n26045, ZN => n20965);
   U12091 : NAND2_X1 port map( A1 => n6883, A2 => n11904, ZN => n1850);
   U12092 : NAND2_X1 port map( A1 => n1239, A2 => n25744, ZN => n7415);
   U12094 : OAI21_X1 port map( A1 => n4163, A2 => n3517, B => n5356, ZN => 
                           n3516);
   U12097 : NAND2_X1 port map( A1 => n37306, A2 => n5886, ZN => n5883);
   U12101 : AND3_X1 port map( A1 => n19259, A2 => n2830, A3 => n1021, Z => 
                           n4794);
   U12105 : AND2_X1 port map( A1 => n26010, A2 => n26012, Z => n3555);
   U12107 : INV_X1 port map( I => n26131, ZN => n14146);
   U12108 : AND2_X1 port map( A1 => n14133, A2 => n14131, Z => n25938);
   U12111 : OAI22_X1 port map( A1 => n7369, A2 => n31205, B1 => n1014, B2 => 
                           n26024, ZN => n6400);
   U12113 : INV_X1 port map( I => n6180, ZN => n25875);
   U12118 : NAND2_X1 port map( A1 => n18037, A2 => n25961, ZN => n13164);
   U12124 : NAND2_X1 port map( A1 => n17439, A2 => n840, ZN => n5683);
   U12127 : OAI21_X1 port map( A1 => n25982, A2 => n25981, B => n39375, ZN => 
                           n25983);
   U12133 : OAI21_X1 port map( A1 => n4190, A2 => n5098, B => n10834, ZN => 
                           n11904);
   U12135 : AOI21_X1 port map( A1 => n26111, A2 => n14228, B => n951, ZN => 
                           n6589);
   U12139 : AOI21_X1 port map( A1 => n926, A2 => n26018, B => n1020, ZN => 
                           n11763);
   U12142 : NAND2_X1 port map( A1 => n950, A2 => n4699, ZN => n12522);
   U12146 : NAND2_X1 port map( A1 => n11762, A2 => n34898, ZN => n13586);
   U12147 : AND3_X1 port map( A1 => n32690, A2 => n34961, A3 => n38835, Z => 
                           n4884);
   U12153 : NAND2_X1 port map( A1 => n25915, A2 => n25978, ZN => n16977);
   U12156 : NOR2_X1 port map( A1 => n25852, A2 => n13391, ZN => n13067);
   U12160 : NAND2_X1 port map( A1 => n25927, A2 => n5356, ZN => n18958);
   U12165 : NAND2_X1 port map( A1 => n7370, A2 => n26024, ZN => n7369);
   U12167 : INV_X1 port map( I => n17008, ZN => n20530);
   U12170 : AOI21_X1 port map( A1 => n26109, A2 => n14228, B => n1019, ZN => 
                           n17035);
   U12171 : NAND2_X1 port map( A1 => n33293, A2 => n36922, ZN => n4832);
   U12176 : OR2_X1 port map( A1 => n25852, A2 => n31523, Z => n2946);
   U12181 : INV_X1 port map( I => n26110, ZN => n11945);
   U12183 : AND3_X1 port map( A1 => n1240, A2 => n26330, A3 => n931, Z => 
                           n14407);
   U12191 : CLKBUF_X2 port map( I => n26328, Z => n19574);
   U12198 : NAND2_X1 port map( A1 => n26130, A2 => n9916, ZN => n7370);
   U12203 : INV_X1 port map( I => n26113, ZN => n8393);
   U12207 : AND2_X1 port map( A1 => n18162, A2 => n17180, Z => n25783);
   U12208 : INV_X1 port map( I => n26024, ZN => n20769);
   U12215 : NAND2_X1 port map( A1 => n15575, A2 => n17624, ZN => n10234);
   U12216 : NOR3_X1 port map( A1 => n26108, A2 => n1017, A3 => n38760, ZN => 
                           n10137);
   U12218 : NOR2_X1 port map( A1 => n31205, A2 => n25813, ZN => n7699);
   U12220 : NOR2_X1 port map( A1 => n4385, A2 => n2625, ZN => n8376);
   U12224 : NAND2_X1 port map( A1 => n5753, A2 => n33440, ZN => n7134);
   U12235 : INV_X1 port map( I => n36546, ZN => n6221);
   U12246 : AND2_X1 port map( A1 => n25836, A2 => n33997, Z => n14694);
   U12250 : NAND2_X1 port map( A1 => n25567, A2 => n19438, ZN => n16569);
   U12257 : NOR2_X1 port map( A1 => n4048, A2 => n8906, ZN => n8905);
   U12269 : NAND2_X1 port map( A1 => n13195, A2 => n19367, ZN => n13194);
   U12274 : INV_X1 port map( I => n17305, ZN => n4433);
   U12275 : NOR2_X1 port map( A1 => n7853, A2 => n5519, ZN => n5711);
   U12286 : NAND2_X1 port map( A1 => n20876, A2 => n19237, ZN => n20875);
   U12296 : NAND2_X1 port map( A1 => n6762, A2 => n6763, ZN => n1932);
   U12298 : INV_X1 port map( I => n38825, ZN => n25904);
   U12300 : CLKBUF_X2 port map( I => n26124, Z => n9682);
   U12307 : INV_X1 port map( I => n25479, ZN => n8978);
   U12308 : AND3_X1 port map( A1 => n25719, A2 => n18519, A3 => n18831, Z => 
                           n8689);
   U12310 : NOR2_X1 port map( A1 => n7235, A2 => n25721, ZN => n7234);
   U12313 : AND2_X1 port map( A1 => n39289, A2 => n953, Z => n8878);
   U12318 : OAI21_X1 port map( A1 => n25437, A2 => n39389, B => n39599, ZN => 
                           n25438);
   U12323 : OAI21_X1 port map( A1 => n25427, A2 => n19302, B => n34150, ZN => 
                           n25714);
   U12337 : OAI21_X1 port map( A1 => n12478, A2 => n33950, B => n20648, ZN => 
                           n11333);
   U12340 : OAI21_X1 port map( A1 => n25698, A2 => n17774, B => n11641, ZN => 
                           n16229);
   U12343 : AND2_X1 port map( A1 => n17303, A2 => n25389, Z => n4988);
   U12344 : NAND2_X1 port map( A1 => n1022, A2 => n36019, ZN => n18694);
   U12345 : NAND2_X1 port map( A1 => n38178, A2 => n8033, ZN => n8032);
   U12349 : AND2_X1 port map( A1 => n25719, A2 => n25557, Z => n17282);
   U12350 : NAND2_X1 port map( A1 => n14056, A2 => n34464, ZN => n14192);
   U12352 : NAND2_X1 port map( A1 => n17450, A2 => n18831, ZN => n13195);
   U12356 : NOR2_X1 port map( A1 => n24894, A2 => n25449, ZN => n8122);
   U12365 : NOR2_X1 port map( A1 => n32101, A2 => n7802, ZN => n18988);
   U12368 : AND2_X1 port map( A1 => n38359, A2 => n3736, Z => n3735);
   U12371 : NAND2_X1 port map( A1 => n14947, A2 => n11874, ZN => n5901);
   U12373 : NAND2_X1 port map( A1 => n25577, A2 => n25660, ZN => n11806);
   U12374 : OR2_X1 port map( A1 => n1109, A2 => n25660, Z => n13826);
   U12376 : NAND2_X1 port map( A1 => n25012, A2 => n25337, ZN => n6939);
   U12378 : NOR2_X1 port map( A1 => n32419, A2 => n4048, ZN => n4047);
   U12380 : NAND2_X1 port map( A1 => n33826, A2 => n25425, ZN => n4791);
   U12386 : NAND2_X1 port map( A1 => n4755, A2 => n5798, ZN => n4754);
   U12389 : OAI21_X1 port map( A1 => n25448, A2 => n38782, B => n17304, ZN => 
                           n4989);
   U12390 : NAND2_X1 port map( A1 => n18734, A2 => n1256, ZN => n7878);
   U12397 : INV_X1 port map( I => n25548, ZN => n12417);
   U12398 : OR2_X1 port map( A1 => n18909, A2 => n21254, Z => n4976);
   U12409 : AND3_X1 port map( A1 => n25689, A2 => n19548, A3 => n31557, Z => 
                           n25506);
   U12410 : NAND3_X1 port map( A1 => n25681, A2 => n25680, A3 => n25679, ZN => 
                           n13589);
   U12413 : INV_X1 port map( I => n9441, ZN => n9241);
   U12414 : AND3_X1 port map( A1 => n25540, A2 => n5042, A3 => n25513, Z => 
                           n14613);
   U12425 : AND2_X1 port map( A1 => n12500, A2 => n7866, Z => n12768);
   U12432 : AND2_X1 port map( A1 => n541, A2 => n319, Z => n14666);
   U12433 : OR2_X1 port map( A1 => n20052, A2 => n25477, Z => n11924);
   U12434 : OR2_X1 port map( A1 => n33130, A2 => n14460, Z => n14490);
   U12444 : AND2_X1 port map( A1 => n25355, A2 => n24896, Z => n4674);
   U12445 : NOR2_X1 port map( A1 => n14472, A2 => n24963, ZN => n10973);
   U12446 : OAI21_X1 port map( A1 => n14475, A2 => n15180, B => n25401, ZN => 
                           n20859);
   U12449 : NAND2_X1 port map( A1 => n17281, A2 => n18519, ZN => n7238);
   U12452 : OR2_X1 port map( A1 => n19701, A2 => n16933, Z => n25333);
   U12455 : NAND2_X1 port map( A1 => n17183, A2 => n14602, ZN => n11063);
   U12458 : INV_X1 port map( I => n19636, ZN => n25385);
   U12460 : OR2_X1 port map( A1 => n25670, A2 => n18164, Z => n11647);
   U12461 : NAND2_X1 port map( A1 => n25408, A2 => n25606, ZN => n4647);
   U12465 : INV_X1 port map( I => n25725, ZN => n25633);
   U12472 : AND2_X1 port map( A1 => n25412, A2 => n25307, Z => n16911);
   U12476 : AND2_X1 port map( A1 => n8304, A2 => n37926, Z => n14475);
   U12486 : NAND3_X1 port map( A1 => n8764, A2 => n5501, A3 => n7990, ZN => 
                           n5500);
   U12492 : INV_X1 port map( I => n25022, ZN => n8764);
   U12496 : OAI21_X1 port map( A1 => n9183, A2 => n9182, B => n7967, ZN => 
                           n9181);
   U12500 : INV_X1 port map( I => n9177, ZN => n5501);
   U12505 : INV_X1 port map( I => n39541, ZN => n9564);
   U12506 : INV_X1 port map( I => n16819, ZN => n16420);
   U12508 : INV_X1 port map( I => n6759, ZN => n8447);
   U12509 : INV_X1 port map( I => n7968, ZN => n7966);
   U12511 : INV_X1 port map( I => n17904, ZN => n9182);
   U12518 : INV_X1 port map( I => n25127, ZN => n17445);
   U12519 : INV_X1 port map( I => n18211, ZN => n6896);
   U12521 : INV_X2 port map( I => n18395, ZN => n1553);
   U12523 : INV_X1 port map( I => n16581, ZN => n9438);
   U12526 : NAND2_X1 port map( A1 => n1118, A2 => n2747, ZN => n16820);
   U12527 : INV_X1 port map( I => n16751, ZN => n8608);
   U12531 : NOR2_X1 port map( A1 => n10988, A2 => n10648, ZN => n2847);
   U12533 : INV_X1 port map( I => n15945, ZN => n8607);
   U12534 : INV_X1 port map( I => n4063, ZN => n4062);
   U12546 : INV_X1 port map( I => n9528, ZN => n17100);
   U12548 : NAND2_X1 port map( A1 => n13582, A2 => n13581, ZN => n14534);
   U12549 : INV_X1 port map( I => n24813, ZN => n9183);
   U12564 : NAND2_X1 port map( A1 => n36955, A2 => n3750, ZN => n3749);
   U12567 : NAND2_X1 port map( A1 => n1907, A2 => n19279, ZN => n1906);
   U12569 : NOR2_X1 port map( A1 => n15527, A2 => n5933, ZN => n15526);
   U12570 : OAI21_X1 port map( A1 => n10114, A2 => n9849, B => n24735, ZN => 
                           n4688);
   U12571 : INV_X1 port map( I => n7969, ZN => n7972);
   U12572 : INV_X1 port map( I => n24540, ZN => n16750);
   U12587 : NAND2_X1 port map( A1 => n24755, A2 => n19339, ZN => n17962);
   U12592 : NAND2_X1 port map( A1 => n7242, A2 => n24691, ZN => n7241);
   U12594 : NAND2_X1 port map( A1 => n24733, A2 => n16815, ZN => n3630);
   U12598 : NAND2_X1 port map( A1 => n13553, A2 => n13554, ZN => n12363);
   U12604 : NAND2_X1 port map( A1 => n8428, A2 => n8426, ZN => n11610);
   U12609 : NOR2_X1 port map( A1 => n2634, A2 => n1029, ZN => n20926);
   U12612 : NOR2_X1 port map( A1 => n6038, A2 => n36186, ZN => n6037);
   U12613 : NAND2_X1 port map( A1 => n14167, A2 => n24820, ZN => n4349);
   U12615 : INV_X1 port map( I => n24704, ZN => n2697);
   U12616 : INV_X1 port map( I => n24494, ZN => n13214);
   U12623 : NOR2_X1 port map( A1 => n31722, A2 => n18508, ZN => n13628);
   U12632 : NAND2_X1 port map( A1 => n35250, A2 => n14211, ZN => n24842);
   U12639 : INV_X1 port map( I => n24581, ZN => n16871);
   U12651 : NAND2_X1 port map( A1 => n4008, A2 => n24764, ZN => n10353);
   U12652 : INV_X1 port map( I => n24602, ZN => n3374);
   U12672 : INV_X1 port map( I => n24591, ZN => n6838);
   U12674 : NAND2_X1 port map( A1 => n5934, A2 => n16547, ZN => n5933);
   U12677 : INV_X1 port map( I => n5934, ZN => n2537);
   U12681 : INV_X1 port map( I => n32831, ZN => n13518);
   U12686 : NAND2_X1 port map( A1 => n24788, A2 => n24787, ZN => n7065);
   U12697 : NAND2_X1 port map( A1 => n17618, A2 => n14276, ZN => n14275);
   U12705 : INV_X1 port map( I => n24847, ZN => n11714);
   U12707 : NAND2_X1 port map( A1 => n24614, A2 => n24812, ZN => n12160);
   U12708 : NOR2_X1 port map( A1 => n39523, A2 => n38317, ZN => n2698);
   U12712 : NAND2_X1 port map( A1 => n24818, A2 => n17618, ZN => n4350);
   U12714 : NOR2_X1 port map( A1 => n1029, A2 => n19422, ZN => n20013);
   U12715 : INV_X1 port map( I => n24779, ZN => n7515);
   U12722 : NAND3_X1 port map( A1 => n8842, A2 => n8843, A3 => n8839, ZN => 
                           n18508);
   U12733 : NOR2_X1 port map( A1 => n8841, A2 => n8840, ZN => n8839);
   U12734 : OR2_X1 port map( A1 => n19422, A2 => n17101, Z => n18771);
   U12736 : NOR2_X1 port map( A1 => n24811, A2 => n24810, ZN => n3626);
   U12738 : NAND2_X1 port map( A1 => n16238, A2 => n35981, ZN => n9149);
   U12740 : NAND2_X1 port map( A1 => n24874, A2 => n31519, ZN => n5607);
   U12744 : INV_X2 port map( I => n24878, ZN => n1570);
   U12756 : NAND2_X1 port map( A1 => n20654, A2 => n24222, ZN => n5712);
   U12760 : INV_X1 port map( I => n15365, ZN => n8841);
   U12761 : INV_X1 port map( I => n7813, ZN => n7812);
   U12771 : AOI21_X1 port map( A1 => n2400, A2 => n16106, B => n24330, ZN => 
                           n15497);
   U12779 : NOR2_X1 port map( A1 => n11316, A2 => n23797, ZN => n7624);
   U12795 : NAND2_X1 port map( A1 => n24441, A2 => n24440, ZN => n10784);
   U12799 : NAND3_X1 port map( A1 => n16313, A2 => n24086, A3 => n13513, ZN => 
                           n16312);
   U12809 : NAND2_X1 port map( A1 => n24297, A2 => n8847, ZN => n8846);
   U12813 : NAND2_X1 port map( A1 => n1031, A2 => n19895, ZN => n2977);
   U12818 : NAND2_X1 port map( A1 => n12665, A2 => n38431, ZN => n20172);
   U12824 : OAI21_X1 port map( A1 => n39818, A2 => n7210, B => n24121, ZN => 
                           n24125);
   U12827 : OAI21_X1 port map( A1 => n35712, A2 => n19653, B => n4687, ZN => 
                           n5140);
   U12830 : INV_X1 port map( I => n21114, ZN => n8842);
   U12839 : NAND2_X1 port map( A1 => n7773, A2 => n7772, ZN => n24096);
   U12848 : NAND2_X1 port map( A1 => n24355, A2 => n1128, ZN => n8361);
   U12850 : NAND2_X1 port map( A1 => n24141, A2 => n24359, ZN => n13227);
   U12855 : NAND2_X1 port map( A1 => n11134, A2 => n1285, ZN => n6954);
   U12872 : NAND2_X1 port map( A1 => n11261, A2 => n1035, ZN => n11260);
   U12880 : INV_X1 port map( I => n10421, ZN => n24627);
   U12882 : NAND2_X1 port map( A1 => n8501, A2 => n8500, ZN => n8499);
   U12890 : NAND2_X1 port map( A1 => n3142, A2 => n37047, ZN => n24377);
   U12898 : NAND2_X1 port map( A1 => n12248, A2 => n20839, ZN => n13808);
   U12900 : AND2_X1 port map( A1 => n24303, A2 => n1126, Z => n24304);
   U12902 : INV_X1 port map( I => n23855, ZN => n6175);
   U12904 : NAND2_X1 port map( A1 => n24400, A2 => n1284, ZN => n23817);
   U12905 : OR2_X1 port map( A1 => n24275, A2 => n24180, Z => n14654);
   U12907 : NAND2_X1 port map( A1 => n12759, A2 => n1276, ZN => n13692);
   U12909 : NOR2_X1 port map( A1 => n20312, A2 => n15320, ZN => n2268);
   U12912 : NAND2_X1 port map( A1 => n24198, A2 => n32891, ZN => n24199);
   U12914 : AND2_X1 port map( A1 => n18466, A2 => n24373, Z => n24374);
   U12915 : NOR2_X1 port map( A1 => n3453, A2 => n30454, ZN => n14898);
   U12919 : NOR2_X1 port map( A1 => n24223, A2 => n24432, ZN => n5714);
   U12921 : NOR2_X1 port map( A1 => n24360, A2 => n39814, ZN => n15256);
   U12924 : NAND2_X1 port map( A1 => n24426, A2 => n38972, ZN => n18532);
   U12927 : NOR2_X1 port map( A1 => n1276, A2 => n5985, ZN => n12277);
   U12929 : OR2_X1 port map( A1 => n24238, A2 => n20313, Z => n13636);
   U12931 : NOR2_X1 port map( A1 => n23855, A2 => n12771, ZN => n10691);
   U12934 : AND2_X1 port map( A1 => n37229, A2 => n21125, Z => n21124);
   U12935 : NAND2_X1 port map( A1 => n19990, A2 => n24461, ZN => n24460);
   U12939 : AOI21_X1 port map( A1 => n1274, A2 => n19653, B => n13970, ZN => 
                           n9360);
   U12946 : AND2_X1 port map( A1 => n14255, A2 => n24119, Z => n7950);
   U12950 : NAND3_X1 port map( A1 => n14718, A2 => n14717, A3 => n24309, ZN => 
                           n13548);
   U12952 : OR2_X1 port map( A1 => n24152, A2 => n14491, Z => n5432);
   U12953 : NAND2_X1 port map( A1 => n14699, A2 => n20537, ZN => n12120);
   U12955 : AND2_X1 port map( A1 => n24446, A2 => n24445, Z => n24447);
   U12958 : AND2_X1 port map( A1 => n24296, A2 => n8825, Z => n9084);
   U12961 : AND2_X1 port map( A1 => n23819, A2 => n24116, Z => n8500);
   U12967 : AND2_X1 port map( A1 => n24309, A2 => n24446, Z => n18141);
   U12969 : NAND2_X1 port map( A1 => n24232, A2 => n545, ZN => n4361);
   U12976 : INV_X2 port map( I => n39467, ZN => n1587);
   U12978 : NAND2_X1 port map( A1 => n24446, A2 => n24445, ZN => n14717);
   U12980 : INV_X1 port map( I => n5985, ZN => n18295);
   U12984 : OR2_X1 port map( A1 => n24267, A2 => n24445, Z => n13513);
   U12985 : INV_X1 port map( I => n24207, ZN => n24218);
   U12989 : NOR3_X1 port map( A1 => n94, A2 => n3869, A3 => n370, ZN => n15205)
                           ;
   U12997 : NAND2_X1 port map( A1 => n1282, A2 => n1288, ZN => n13040);
   U12999 : INV_X2 port map( I => n13444, ZN => n19007);
   U13001 : NAND2_X1 port map( A1 => n24372, A2 => n24225, ZN => n16644);
   U13002 : NOR2_X1 port map( A1 => n5985, A2 => n19915, ZN => n20068);
   U13003 : NAND2_X1 port map( A1 => n36380, A2 => n1131, ZN => n16141);
   U13007 : OR2_X1 port map( A1 => n800, A2 => n33937, Z => n14686);
   U13008 : NOR2_X1 port map( A1 => n17871, A2 => n14491, ZN => n7880);
   U13012 : NOR2_X1 port map( A1 => n37230, A2 => n20404, ZN => n7835);
   U13023 : INV_X2 port map( I => n11795, ZN => n18697);
   U13026 : INV_X1 port map( I => n24245, ZN => n9519);
   U13039 : OR2_X1 port map( A1 => n24445, A2 => n24266, Z => n14718);
   U13040 : NOR2_X1 port map( A1 => n39815, A2 => n24110, ZN => n10800);
   U13044 : INV_X1 port map( I => n14471, ZN => n11004);
   U13051 : INV_X2 port map( I => n13540, ZN => n1609);
   U13055 : INV_X1 port map( I => n23920, ZN => n5441);
   U13057 : INV_X1 port map( I => n23802, ZN => n7673);
   U13058 : NAND2_X1 port map( A1 => n12820, A2 => n12819, ZN => n15971);
   U13061 : INV_X1 port map( I => n12798, ZN => n5005);
   U13066 : INV_X1 port map( I => n24062, ZN => n20715);
   U13077 : INV_X1 port map( I => n12821, ZN => n12820);
   U13080 : INV_X1 port map( I => n33322, ZN => n23805);
   U13081 : INV_X1 port map( I => n38175, ZN => n23919);
   U13083 : NOR2_X1 port map( A1 => n22806, A2 => n10174, ZN => n10614);
   U13084 : INV_X1 port map( I => n23710, ZN => n23769);
   U13085 : INV_X1 port map( I => n5841, ZN => n11116);
   U13090 : INV_X1 port map( I => n15800, ZN => n5914);
   U13097 : INV_X1 port map( I => n24047, ZN => n6626);
   U13098 : NOR2_X1 port map( A1 => n10205, A2 => n10204, ZN => n10110);
   U13100 : INV_X1 port map( I => n24053, ZN => n12842);
   U13105 : INV_X1 port map( I => n23685, ZN => n23851);
   U13116 : NAND2_X1 port map( A1 => n9795, A2 => n9794, ZN => n18889);
   U13119 : INV_X1 port map( I => n10207, ZN => n10204);
   U13120 : INV_X1 port map( I => n10208, ZN => n10205);
   U13129 : INV_X2 port map( I => n14219, ZN => n1618);
   U13132 : NAND2_X1 port map( A1 => n17888, A2 => n23315, ZN => n16370);
   U13140 : NAND2_X1 port map( A1 => n11723, A2 => n23400, ZN => n18918);
   U13141 : INV_X1 port map( I => n17423, ZN => n8986);
   U13152 : INV_X1 port map( I => n6561, ZN => n21046);
   U13166 : INV_X1 port map( I => n23217, ZN => n2599);
   U13173 : NAND2_X1 port map( A1 => n6637, A2 => n6993, ZN => n6992);
   U13177 : NOR2_X1 port map( A1 => n23512, A2 => n23513, ZN => n7333);
   U13185 : AOI21_X1 port map( A1 => n23247, A2 => n14011, B => n7008, ZN => 
                           n20118);
   U13192 : NAND2_X1 port map( A1 => n23471, A2 => n23636, ZN => n20504);
   U13201 : NOR2_X1 port map( A1 => n21051, A2 => n8965, ZN => n8964);
   U13205 : NAND2_X1 port map( A1 => n37209, A2 => n37757, ZN => n22824);
   U13208 : NAND2_X1 port map( A1 => n21156, A2 => n23641, ZN => n3274);
   U13209 : NAND2_X1 port map( A1 => n23575, A2 => n20955, ZN => n3743);
   U13210 : INV_X1 port map( I => n9796, ZN => n9795);
   U13214 : NAND3_X1 port map( A1 => n8432, A2 => n11186, A3 => n15176, ZN => 
                           n11185);
   U13219 : NAND2_X1 port map( A1 => n6217, A2 => n6216, ZN => n14623);
   U13221 : INV_X1 port map( I => n20100, ZN => n3383);
   U13231 : INV_X1 port map( I => n17875, ZN => n7146);
   U13232 : OR2_X1 port map( A1 => n23194, A2 => n33349, Z => n20629);
   U13241 : NAND2_X1 port map( A1 => n36829, A2 => n1039, ZN => n9794);
   U13242 : NAND2_X1 port map( A1 => n1295, A2 => n34506, ZN => n17768);
   U13243 : NAND2_X1 port map( A1 => n38248, A2 => n14477, ZN => n19068);
   U13251 : INV_X1 port map( I => n11186, ZN => n11187);
   U13253 : OAI21_X1 port map( A1 => n17511, A2 => n1139, B => n20343, ZN => 
                           n12011);
   U13263 : NAND2_X1 port map( A1 => n38244, A2 => n1306, ZN => n2961);
   U13269 : NAND2_X1 port map( A1 => n23747, A2 => n39805, ZN => n23752);
   U13274 : AOI21_X1 port map( A1 => n39300, A2 => n10216, B => n32366, ZN => 
                           n4534);
   U13276 : AOI21_X1 port map( A1 => n22987, A2 => n22986, B => n18762, ZN => 
                           n16033);
   U13283 : NOR2_X1 port map( A1 => n31908, A2 => n13414, ZN => n23555);
   U13289 : INV_X1 port map( I => n23543, ZN => n2921);
   U13292 : INV_X1 port map( I => n8249, ZN => n2812);
   U13294 : NAND2_X1 port map( A1 => n3716, A2 => n4618, ZN => n2928);
   U13301 : AND2_X1 port map( A1 => n32377, A2 => n13150, Z => n13560);
   U13303 : NAND2_X1 port map( A1 => n9321, A2 => n14477, ZN => n2683);
   U13305 : INV_X1 port map( I => n23576, ZN => n6301);
   U13312 : OR2_X1 port map( A1 => n35331, A2 => n14235, Z => n10122);
   U13313 : AND2_X1 port map( A1 => n52, A2 => n37431, Z => n19379);
   U13314 : NAND2_X1 port map( A1 => n34012, A2 => n8249, ZN => n1894);
   U13320 : AND2_X1 port map( A1 => n33894, A2 => n7335, Z => n16575);
   U13325 : AND2_X1 port map( A1 => n23580, A2 => n10174, Z => n23257);
   U13327 : AND2_X1 port map( A1 => n34959, A2 => n18866, Z => n9192);
   U13336 : NAND2_X1 port map( A1 => n13095, A2 => n11588, ZN => n13094);
   U13337 : NAND2_X1 port map( A1 => n3717, A2 => n23566, ZN => n3716);
   U13339 : NAND2_X1 port map( A1 => n9340, A2 => n23158, ZN => n6346);
   U13355 : NAND2_X1 port map( A1 => n22369, A2 => n3289, ZN => n6917);
   U13360 : NAND2_X1 port map( A1 => n22858, A2 => n13515, ZN => n16301);
   U13365 : AND2_X1 port map( A1 => n5657, A2 => n38282, Z => n8459);
   U13366 : NAND2_X1 port map( A1 => n16053, A2 => n22894, ZN => n22896);
   U13375 : NOR2_X1 port map( A1 => n15947, A2 => n23120, ZN => n13095);
   U13381 : NAND2_X1 port map( A1 => n9472, A2 => n36453, ZN => n15345);
   U13383 : NAND2_X1 port map( A1 => n11197, A2 => n14725, ZN => n18856);
   U13390 : AND2_X1 port map( A1 => n23042, A2 => n1144, Z => n9322);
   U13392 : NOR2_X1 port map( A1 => n22791, A2 => n23172, ZN => n20076);
   U13397 : AND3_X1 port map( A1 => n11584, A2 => n11582, A3 => n34184, Z => 
                           n11583);
   U13398 : AOI21_X1 port map( A1 => n20175, A2 => n20174, B => n20173, ZN => 
                           n22885);
   U13400 : NOR2_X1 port map( A1 => n23046, A2 => n11582, ZN => n4963);
   U13402 : NOR2_X1 port map( A1 => n19082, A2 => n1143, ZN => n5806);
   U13403 : NAND2_X1 port map( A1 => n16957, A2 => n16956, ZN => n12253);
   U13408 : INV_X1 port map( I => n23044, ZN => n2726);
   U13413 : OR2_X1 port map( A1 => n23005, A2 => n19823, Z => n5895);
   U13416 : NAND2_X1 port map( A1 => n22909, A2 => n22908, ZN => n21229);
   U13419 : NAND2_X1 port map( A1 => n22792, A2 => n22804, ZN => n8806);
   U13433 : NOR2_X1 port map( A1 => n15741, A2 => n32032, ZN => n15740);
   U13437 : NOR2_X1 port map( A1 => n22947, A2 => n23175, ZN => n15742);
   U13438 : INV_X1 port map( I => n23072, ZN => n16617);
   U13440 : INV_X1 port map( I => n22947, ZN => n22960);
   U13441 : INV_X1 port map( I => n22924, ZN => n5747);
   U13472 : INV_X1 port map( I => n13373, ZN => n18462);
   U13487 : OR2_X2 port map( A1 => n34073, A2 => n16692, Z => n7130);
   U13498 : NAND2_X1 port map( A1 => n22916, A2 => n19870, ZN => n8143);
   U13505 : AOI21_X1 port map( A1 => n33082, A2 => n11658, B => n34184, ZN => 
                           n16957);
   U13507 : AND2_X1 port map( A1 => n38282, A2 => n23198, Z => n10552);
   U13512 : NAND2_X1 port map( A1 => n22850, A2 => n37335, ZN => n14658);
   U13513 : AND2_X1 port map( A1 => n5515, A2 => n14442, Z => n5786);
   U13516 : NOR2_X1 port map( A1 => n640, A2 => n39527, ZN => n6902);
   U13517 : INV_X1 port map( I => n11704, ZN => n9660);
   U13527 : INV_X1 port map( I => n23030, ZN => n5621);
   U13528 : NAND2_X1 port map( A1 => n11295, A2 => n23124, ZN => n22769);
   U13532 : INV_X1 port map( I => n19319, ZN => n23068);
   U13538 : AND2_X1 port map( A1 => n22915, A2 => n23163, Z => n22916);
   U13540 : NOR2_X1 port map( A1 => n36724, A2 => n19535, ZN => n19246);
   U13543 : CLKBUF_X2 port map( I => n10071, Z => n9725);
   U13544 : INV_X1 port map( I => n12032, ZN => n22807);
   U13550 : NAND2_X1 port map( A1 => n10634, A2 => n19859, ZN => n7013);
   U13556 : AND2_X1 port map( A1 => n39155, A2 => n18415, Z => n6385);
   U13557 : CLKBUF_X2 port map( I => n22857, Z => n7537);
   U13570 : INV_X2 port map( I => n9176, ZN => n18415);
   U13582 : NAND2_X1 port map( A1 => n9334, A2 => n4413, ZN => n10729);
   U13583 : INV_X1 port map( I => n9334, ZN => n22587);
   U13584 : NAND2_X1 port map( A1 => n10556, A2 => n10555, ZN => n11255);
   U13587 : INV_X1 port map( I => n15413, ZN => n12194);
   U13589 : INV_X1 port map( I => n22654, ZN => n13354);
   U13590 : INV_X1 port map( I => n3969, ZN => n2236);
   U13592 : INV_X1 port map( I => n22531, ZN => n22291);
   U13596 : INV_X1 port map( I => n22500, ZN => n3623);
   U13599 : INV_X1 port map( I => n14309, ZN => n7593);
   U13603 : NAND2_X1 port map( A1 => n38099, A2 => n9483, ZN => n8549);
   U13610 : INV_X2 port map( I => n22348, ZN => n1658);
   U13615 : INV_X1 port map( I => n22488, ZN => n10862);
   U13616 : CLKBUF_X2 port map( I => n19328, Z => n4819);
   U13619 : INV_X1 port map( I => n9116, ZN => n9115);
   U13620 : INV_X1 port map( I => n8552, ZN => n22666);
   U13621 : INV_X1 port map( I => n22485, ZN => n2986);
   U13622 : INV_X2 port map( I => n16667, ZN => n1661);
   U13624 : INV_X1 port map( I => n19221, ZN => n22675);
   U13626 : AOI21_X1 port map( A1 => n12567, A2 => n22162, B => n19890, ZN => 
                           n6773);
   U13627 : INV_X1 port map( I => n12324, ZN => n6121);
   U13628 : NOR2_X1 port map( A1 => n12325, A2 => n19801, ZN => n6120);
   U13629 : OAI21_X1 port map( A1 => n12324, A2 => n12325, B => n19801, ZN => 
                           n6125);
   U13630 : INV_X1 port map( I => n31504, ZN => n14322);
   U13631 : NAND3_X1 port map( A1 => n12661, A2 => n29334, A3 => n12660, ZN => 
                           n10555);
   U13635 : NAND2_X1 port map( A1 => n22381, A2 => n22380, ZN => n22637);
   U13636 : INV_X2 port map( I => n36886, ZN => n1663);
   U13642 : INV_X1 port map( I => n22298, ZN => n6015);
   U13645 : NAND2_X1 port map( A1 => n19976, A2 => n17096, ZN => n3236);
   U13647 : OAI21_X1 port map( A1 => n8749, A2 => n37089, B => n4851, ZN => 
                           n7058);
   U13648 : NAND2_X1 port map( A1 => n18950, A2 => n18953, ZN => n17041);
   U13649 : NAND2_X1 port map( A1 => n13570, A2 => n11091, ZN => n4662);
   U13654 : INV_X1 port map( I => n3967, ZN => n2237);
   U13657 : NAND2_X1 port map( A1 => n22242, A2 => n8749, ZN => n2590);
   U13661 : NAND2_X1 port map( A1 => n13279, A2 => n17147, ZN => n7490);
   U13665 : OAI21_X1 port map( A1 => n39075, A2 => n1149, B => n10092, ZN => 
                           n19284);
   U13675 : AND2_X1 port map( A1 => n21801, A2 => n33886, Z => n19292);
   U13677 : NAND2_X1 port map( A1 => n22123, A2 => n11149, ZN => n12345);
   U13692 : NAND2_X1 port map( A1 => n22134, A2 => n1327, ZN => n11047);
   U13693 : NAND2_X1 port map( A1 => n7818, A2 => n7817, ZN => n7816);
   U13696 : NAND2_X1 port map( A1 => n22271, A2 => n12814, ZN => n5149);
   U13700 : AND2_X1 port map( A1 => n22325, A2 => n31092, Z => n14535);
   U13705 : NOR2_X1 port map( A1 => n21363, A2 => n31649, ZN => n6557);
   U13711 : NOR2_X1 port map( A1 => n22089, A2 => n18656, ZN => n13279);
   U13714 : OAI21_X1 port map( A1 => n37089, A2 => n34808, B => n13055, ZN => 
                           n22403);
   U13718 : OAI22_X1 port map( A1 => n6722, A2 => n10261, B1 => n5819, B2 => 
                           n22189, ZN => n6721);
   U13719 : NAND2_X1 port map( A1 => n1149, A2 => n6129, ZN => n4661);
   U13720 : INV_X1 port map( I => n10631, ZN => n7771);
   U13729 : NOR2_X1 port map( A1 => n22349, A2 => n916, ZN => n5577);
   U13730 : OAI21_X1 port map( A1 => n14423, A2 => n1332, B => n19873, ZN => 
                           n5576);
   U13733 : NOR3_X1 port map( A1 => n3003, A2 => n3001, A3 => n17359, ZN => 
                           n3002);
   U13738 : INV_X1 port map( I => n5302, ZN => n20759);
   U13742 : INV_X1 port map( I => n4283, ZN => n18675);
   U13743 : NOR2_X1 port map( A1 => n22147, A2 => n22239, ZN => n13633);
   U13746 : NOR2_X1 port map( A1 => n22267, A2 => n33782, ZN => n21262);
   U13747 : NAND2_X1 port map( A1 => n10434, A2 => n32889, ZN => n10433);
   U13748 : NAND2_X1 port map( A1 => n19486, A2 => n22282, ZN => n13980);
   U13749 : OR2_X1 port map( A1 => n22360, A2 => n31939, Z => n14683);
   U13750 : AOI21_X1 port map( A1 => n22289, A2 => n22041, B => n2840, ZN => 
                           n13420);
   U13751 : NOR2_X1 port map( A1 => n22367, A2 => n22365, ZN => n13296);
   U13753 : NAND2_X1 port map( A1 => n1331, A2 => n36237, ZN => n4629);
   U13755 : NAND2_X1 port map( A1 => n22151, A2 => n33678, ZN => n17973);
   U13764 : INV_X1 port map( I => n16511, ZN => n16772);
   U13766 : NOR2_X1 port map( A1 => n20869, A2 => n2910, ZN => n11542);
   U13769 : NAND2_X1 port map( A1 => n17639, A2 => n22184, ZN => n17638);
   U13770 : NOR2_X1 port map( A1 => n10681, A2 => n34488, ZN => n4110);
   U13771 : INV_X1 port map( I => n22111, ZN => n4932);
   U13772 : NAND2_X1 port map( A1 => n36151, A2 => n15493, ZN => n7294);
   U13776 : NAND2_X1 port map( A1 => n9224, A2 => n9223, ZN => n9222);
   U13784 : OR2_X1 port map( A1 => n22030, A2 => n5075, Z => n9126);
   U13785 : OR2_X1 port map( A1 => n34813, A2 => n19873, Z => n5206);
   U13788 : AND4_X1 port map( A1 => n10650, A2 => n685, A3 => n10649, A4 => 
                           n10652, Z => n10651);
   U13794 : NOR2_X1 port map( A1 => n17307, A2 => n19773, ZN => n21261);
   U13796 : NOR3_X1 port map( A1 => n22263, A2 => n22262, A3 => n22264, ZN => 
                           n4336);
   U13797 : AND2_X1 port map( A1 => n21961, A2 => n22130, Z => n12255);
   U13799 : AND2_X1 port map( A1 => n21961, A2 => n12892, Z => n6722);
   U13807 : INV_X2 port map( I => n21973, ZN => n22184);
   U13813 : OR2_X1 port map( A1 => n22086, A2 => n36006, Z => n13837);
   U13817 : CLKBUF_X2 port map( I => n22215, Z => n9938);
   U13818 : INV_X1 port map( I => n18656, ZN => n9129);
   U13823 : INV_X1 port map( I => n37089, ZN => n8439);
   U13824 : NAND2_X1 port map( A1 => n1342, A2 => n20679, ZN => n3678);
   U13826 : NAND2_X1 port map( A1 => n21891, A2 => n18758, ZN => n10417);
   U13834 : NAND2_X1 port map( A1 => n5451, A2 => n5391, ZN => n5448);
   U13835 : NOR2_X1 port map( A1 => n12513, A2 => n21733, ZN => n12512);
   U13842 : AOI21_X1 port map( A1 => n21708, A2 => n19271, B => n21886, ZN => 
                           n21709);
   U13843 : INV_X1 port map( I => n21695, ZN => n10325);
   U13845 : NAND2_X1 port map( A1 => n21710, A2 => n20535, ZN => n10323);
   U13849 : NOR2_X1 port map( A1 => n2458, A2 => n29411, ZN => n17940);
   U13852 : NAND2_X1 port map( A1 => n20037, A2 => n21910, ZN => n13240);
   U13854 : INV_X1 port map( I => n9102, ZN => n7183);
   U13856 : NAND2_X1 port map( A1 => n7414, A2 => n9863, ZN => n4241);
   U13857 : NAND2_X1 port map( A1 => n13098, A2 => n21557, ZN => n6799);
   U13867 : OAI21_X1 port map( A1 => n12737, A2 => n4116, B => n5187, ZN => 
                           n12358);
   U13869 : OR2_X1 port map( A1 => n21843, A2 => n15031, Z => n14572);
   U13872 : AOI21_X1 port map( A1 => n19822, A2 => n14493, B => n19708, ZN => 
                           n19707);
   U13873 : INV_X1 port map( I => n21867, ZN => n10657);
   U13875 : NAND2_X1 port map( A1 => n21550, A2 => n20328, ZN => n6420);
   U13877 : AND2_X1 port map( A1 => n16951, A2 => n21789, Z => n21796);
   U13888 : NAND2_X1 port map( A1 => n21443, A2 => n15031, ZN => n2479);
   U13889 : NAND2_X1 port map( A1 => n21442, A2 => n33285, ZN => n2478);
   U13892 : NAND2_X1 port map( A1 => n2045, A2 => n11274, ZN => n21708);
   U13893 : NAND2_X1 port map( A1 => n2990, A2 => n18205, ZN => n17965);
   U13896 : NAND2_X1 port map( A1 => n17886, A2 => n21653, ZN => n7601);
   U13897 : AOI21_X1 port map( A1 => n21373, A2 => n21372, B => n35973, ZN => 
                           n21374);
   U13898 : NAND2_X1 port map( A1 => n8969, A2 => n21410, ZN => n21127);
   U13899 : NAND2_X1 port map( A1 => n14909, A2 => n21833, ZN => n14908);
   U13901 : AND2_X1 port map( A1 => n21901, A2 => n21900, Z => n14526);
   U13904 : OR2_X1 port map( A1 => n33771, A2 => n11851, Z => n11850);
   U13907 : INV_X2 port map( I => n19091, ZN => n18710);
   U13909 : AND2_X1 port map( A1 => n13959, A2 => n13997, Z => n13685);
   U13911 : NOR2_X1 port map( A1 => n21569, A2 => n3326, ZN => n3325);
   U13912 : NAND2_X1 port map( A1 => n15381, A2 => n6504, ZN => n15380);
   U13913 : AND2_X1 port map( A1 => n21750, A2 => n2532, Z => n16163);
   U13914 : NAND2_X1 port map( A1 => n17233, A2 => n32370, ZN => n13348);
   U13915 : NAND2_X1 port map( A1 => n19169, A2 => n18496, ZN => n10263);
   U13917 : NAND2_X1 port map( A1 => n21545, A2 => n19650, ZN => n13522);
   U13921 : AOI21_X1 port map( A1 => n21923, A2 => n21640, B => n12738, ZN => 
                           n12737);
   U13926 : INV_X1 port map( I => n10875, ZN => n9253);
   U13929 : NAND2_X1 port map( A1 => n19768, A2 => n4094, ZN => n21372);
   U13933 : INV_X1 port map( I => n11851, ZN => n11239);
   U13935 : NOR2_X1 port map( A1 => n21718, A2 => n1352, ZN => n5503);
   U13939 : INV_X1 port map( I => n1814, ZN => n1813);
   U13940 : INV_X1 port map( I => n21450, ZN => n16873);
   U13941 : NOR2_X1 port map( A1 => n21749, A2 => n21748, ZN => n18274);
   U13942 : INV_X1 port map( I => n17848, ZN => n12109);
   U13944 : OR3_X1 port map( A1 => n4759, A2 => n21029, A3 => n19850, Z => 
                           n21891);
   U13945 : NAND2_X1 port map( A1 => n20587, A2 => n21509, ZN => n17820);
   U13946 : NAND2_X1 port map( A1 => n13997, A2 => n10211, ZN => n13158);
   U13951 : AND2_X1 port map( A1 => n10212, A2 => n695, Z => n21397);
   U13952 : CLKBUF_X2 port map( I => n21688, Z => n21853);
   U13956 : NOR2_X1 port map( A1 => n21465, A2 => n34922, ZN => n20752);
   U13960 : NOR2_X1 port map( A1 => n19699, A2 => n21894, ZN => n3326);
   U13962 : AND2_X1 port map( A1 => n21699, A2 => n18266, Z => n19037);
   U13966 : INV_X2 port map( I => n8799, ZN => n7278);
   U13972 : AND2_X1 port map( A1 => n19542, A2 => n21748, Z => n14542);
   U13976 : CLKBUF_X2 port map( I => n21506, Z => n9642);
   U13980 : CLKBUF_X2 port map( I => n21846, Z => n19392);
   U13986 : INV_X1 port map( I => n29689, ZN => n29690);
   U13987 : INV_X1 port map( I => n30179, ZN => n3711);
   U13993 : INV_X1 port map( I => n29661, ZN => n16641);
   U13994 : INV_X1 port map( I => n29849, ZN => n18691);
   U13995 : INV_X1 port map( I => n30006, ZN => n30007);
   U13998 : CLKBUF_X2 port map( I => n21849, Z => n18219);
   U14001 : INV_X1 port map( I => n30114, ZN => n30115);
   U14003 : INV_X1 port map( I => n19950, ZN => n6462);
   U14004 : INV_X1 port map( I => n19801, ZN => n6429);
   U14005 : INV_X1 port map( I => n29857, ZN => n20420);
   U14009 : INV_X1 port map( I => n19758, ZN => n17316);
   U14010 : INV_X1 port map( I => n29808, ZN => n22285);
   U14011 : INV_X1 port map( I => n29320, ZN => n29321);
   U14013 : CLKBUF_X2 port map( I => n21776, Z => n19350);
   U14014 : INV_X1 port map( I => n29238, ZN => n29239);
   U14015 : INV_X1 port map( I => n19732, ZN => n21048);
   U14017 : INV_X2 port map( I => n8653, ZN => n8799);
   U14019 : INV_X1 port map( I => n19761, ZN => n15599);
   U14020 : INV_X1 port map( I => n19583, ZN => n15888);
   U14023 : INV_X1 port map( I => n15009, ZN => n21782);
   U14024 : CLKBUF_X2 port map( I => Key(134), Z => n19913);
   U14025 : INV_X1 port map( I => Key(178), ZN => n11200);
   U14030 : CLKBUF_X2 port map( I => Key(87), Z => n28934);
   U14035 : CLKBUF_X2 port map( I => Key(131), Z => n30248);
   U14037 : CLKBUF_X2 port map( I => Key(83), Z => n29432);
   U14038 : CLKBUF_X2 port map( I => Key(152), Z => n19883);
   U14039 : CLKBUF_X2 port map( I => Key(53), Z => n29319);
   U14042 : INV_X1 port map( I => n29295, ZN => n1706);
   U14045 : CLKBUF_X2 port map( I => Key(111), Z => n19814);
   U14046 : CLKBUF_X2 port map( I => Key(89), Z => n29671);
   U14048 : CLKBUF_X2 port map( I => Key(71), Z => n10027);
   U14050 : CLKBUF_X2 port map( I => Key(32), Z => n28968);
   U14051 : CLKBUF_X2 port map( I => Key(57), Z => n29476);
   U14056 : CLKBUF_X2 port map( I => Key(101), Z => n29298);
   U14057 : CLKBUF_X2 port map( I => Key(186), Z => n19936);
   U14058 : INV_X1 port map( I => n19825, ZN => n1726);
   U14059 : CLKBUF_X2 port map( I => Key(35), Z => n29707);
   U14060 : CLKBUF_X2 port map( I => Key(161), Z => n29229);
   U14064 : CLKBUF_X2 port map( I => Key(128), Z => n19649);
   U14066 : CLKBUF_X2 port map( I => Key(171), Z => n29661);
   U14067 : INV_X1 port map( I => n30063, ZN => n1737);
   U14069 : CLKBUF_X2 port map( I => Key(59), Z => n29562);
   U14070 : CLKBUF_X2 port map( I => Key(178), Z => n19749);
   U14071 : XOR2_X1 port map( A1 => n1740, A2 => n4041, Z => n1769);
   U14082 : NOR3_X1 port map( A1 => n14791, A2 => n9514, A3 => n1753, ZN => 
                           n1752);
   U14086 : XOR2_X1 port map( A1 => n36895, A2 => n23609, Z => n23771);
   U14087 : XOR2_X1 port map( A1 => n17478, A2 => n36895, Z => n10885);
   U14088 : NOR2_X1 port map( A1 => n20873, A2 => n906, ZN => n18851);
   U14089 : XOR2_X1 port map( A1 => n1758, A2 => n22385, Z => n17628);
   U14092 : NAND2_X1 port map( A1 => n1759, A2 => n15038, ZN => n19327);
   U14095 : NAND2_X2 port map( A1 => n3380, A2 => n1760, ZN => n26553);
   U14099 : XOR2_X1 port map( A1 => n10026, A2 => n16134, Z => n18966);
   U14105 : XOR2_X1 port map( A1 => n22416, A2 => n22417, Z => n1765);
   U14107 : NAND2_X2 port map( A1 => n3226, A2 => n1284, ZN => n23818);
   U14113 : NAND2_X1 port map( A1 => n1771, A2 => n13113, ZN => n13047);
   U14114 : NAND2_X1 port map( A1 => n1771, A2 => n13112, ZN => n13048);
   U14115 : XOR2_X1 port map( A1 => n29029, A2 => n9952, Z => n2217);
   U14120 : XOR2_X1 port map( A1 => n1775, A2 => n28783, Z => n28945);
   U14122 : XOR2_X1 port map( A1 => n1775, A2 => n19816, Z => n8774);
   U14123 : XOR2_X1 port map( A1 => n1775, A2 => n29831, Z => n29834);
   U14125 : NAND3_X1 port map( A1 => n35287, A2 => n4434, A3 => n38079, ZN => 
                           n27317);
   U14130 : NAND2_X1 port map( A1 => n27298, A2 => n1788, ZN => n5082);
   U14136 : XOR2_X1 port map( A1 => n13395, A2 => n19733, Z => n1790);
   U14137 : XOR2_X1 port map( A1 => n23712, A2 => n18006, Z => n24062);
   U14138 : NOR2_X2 port map( A1 => n16033, A2 => n16032, ZN => n18006);
   U14145 : XOR2_X1 port map( A1 => n29073, A2 => n1793, Z => n1792);
   U14146 : XOR2_X1 port map( A1 => n20452, A2 => n29509, Z => n1793);
   U14150 : XOR2_X1 port map( A1 => n13289, A2 => n19875, Z => n18182);
   U14151 : AOI21_X2 port map( A1 => n34036, A2 => n35258, B => n1796, ZN => 
                           n13293);
   U14152 : OAI21_X1 port map( A1 => n29862, A2 => n29960, B => n29955, ZN => 
                           n15140);
   U14154 : NOR2_X2 port map( A1 => n24863, A2 => n13966, ZN => n24862);
   U14155 : NAND2_X2 port map( A1 => n4178, A2 => n4177, ZN => n24863);
   U14158 : INV_X1 port map( I => n29844, ZN => n5972);
   U14159 : NAND2_X1 port map( A1 => n1063, A2 => n20284, ZN => n29844);
   U14163 : XOR2_X1 port map( A1 => n16898, A2 => n1808, Z => n1807);
   U14164 : XOR2_X1 port map( A1 => n17908, A2 => n22568, Z => n1809);
   U14168 : NAND2_X1 port map( A1 => n11344, A2 => n1812, ZN => n21989);
   U14170 : INV_X2 port map( I => n1816, ZN => n21886);
   U14177 : INV_X2 port map( I => n10962, ZN => n13042);
   U14178 : INV_X1 port map( I => n23080, ZN => n23104);
   U14179 : XOR2_X1 port map( A1 => n10963, A2 => n7708, Z => n10962);
   U14185 : NOR2_X1 port map( A1 => n425, A2 => n1827, ZN => n20850);
   U14187 : NAND2_X1 port map( A1 => n25738, A2 => n34485, ZN => n5236);
   U14188 : XOR2_X1 port map( A1 => n35215, A2 => n16296, Z => n16338);
   U14191 : MUX2_X1 port map( I0 => n1836, I1 => n1835, S => n34520, Z => n1834
                           );
   U14192 : NAND2_X1 port map( A1 => n30358, A2 => n27390, ZN => n1836);
   U14198 : OAI22_X2 port map( A1 => n8316, A2 => n38369, B1 => n8315, B2 => 
                           n1844, ZN => n24985);
   U14206 : XOR2_X1 port map( A1 => n23833, A2 => n23801, Z => n21268);
   U14207 : XOR2_X1 port map( A1 => n23695, A2 => n23707, Z => n23833);
   U14220 : XOR2_X1 port map( A1 => n22758, A2 => n1868, Z => n1867);
   U14228 : XOR2_X1 port map( A1 => n1878, A2 => n19627, Z => n4853);
   U14229 : XNOR2_X1 port map( A1 => n10965, A2 => n26554, ZN => n19627);
   U14231 : XOR2_X1 port map( A1 => n1880, A2 => n1879, Z => n1878);
   U14237 : XOR2_X1 port map( A1 => n16864, A2 => n19843, Z => n1884);
   U14239 : XOR2_X1 port map( A1 => n24857, A2 => n25132, Z => n1885);
   U14241 : XOR2_X1 port map( A1 => n25016, A2 => n25266, Z => n19797);
   U14245 : MUX2_X1 port map( I0 => n30134, I1 => n37117, S => n35234, Z => 
                           n3898);
   U14256 : XOR2_X1 port map( A1 => n1897, A2 => n10617, Z => n1896);
   U14259 : XOR2_X1 port map( A1 => n39637, A2 => n29357, Z => n1902);
   U14260 : INV_X2 port map( I => n5966, ZN => n2716);
   U14268 : XOR2_X1 port map( A1 => n1913, A2 => n1912, Z => n1911);
   U14269 : XOR2_X1 port map( A1 => n5652, A2 => n39082, Z => n1912);
   U14271 : XOR2_X1 port map( A1 => n28948, A2 => n38195, Z => n1913);
   U14276 : NAND2_X2 port map( A1 => n15321, A2 => n15323, ZN => n29147);
   U14288 : NAND2_X1 port map( A1 => n5570, A2 => n2121, ZN => n2856);
   U14292 : NAND3_X1 port map( A1 => n25480, A2 => n36083, A3 => n1539, ZN => 
                           n25332);
   U14301 : XOR2_X1 port map( A1 => n1930, A2 => n25015, Z => n2623);
   U14307 : NAND2_X1 port map( A1 => n10015, A2 => n26215, ZN => n1934);
   U14311 : OAI21_X2 port map( A1 => n10336, A2 => n10337, B => n9493, ZN => 
                           n19606);
   U14322 : XOR2_X1 port map( A1 => n1945, A2 => n1947, Z => n17564);
   U14323 : XOR2_X1 port map( A1 => n22723, A2 => n1946, Z => n1945);
   U14324 : XOR2_X1 port map( A1 => n22444, A2 => n30803, Z => n1946);
   U14334 : NAND3_X1 port map( A1 => n26101, A2 => n11148, A3 => n35207, ZN => 
                           n1954);
   U14340 : INV_X2 port map( I => n1961, ZN => n20673);
   U14346 : OR2_X1 port map( A1 => n22145, A2 => n19180, Z => n1966);
   U14350 : NAND2_X2 port map( A1 => n1003, A2 => n865, ZN => n26743);
   U14351 : XOR2_X1 port map( A1 => n7543, A2 => n857, Z => n9618);
   U14362 : XOR2_X1 port map( A1 => n38180, A2 => n1366, Z => n1980);
   U14364 : XOR2_X1 port map( A1 => n26165, A2 => n26180, Z => n26229);
   U14372 : INV_X2 port map( I => n13994, ZN => n2047);
   U14376 : AND2_X1 port map( A1 => n25528, A2 => n36083, Z => n1991);
   U14380 : OAI21_X2 port map( A1 => n2698, A2 => n19836, B => n1995, ZN => 
                           n19725);
   U14388 : XOR2_X1 port map( A1 => n2004, A2 => n2003, Z => n2002);
   U14389 : XOR2_X1 port map( A1 => n29247, A2 => n19681, Z => n2003);
   U14393 : XOR2_X1 port map( A1 => n36596, A2 => n35559, Z => n10201);
   U14396 : NAND2_X1 port map( A1 => n21925, A2 => n2008, ZN => n3437);
   U14399 : OAI21_X2 port map( A1 => n2017, A2 => n2016, B => n2013, ZN => 
                           n29672);
   U14404 : INV_X1 port map( I => n24404, ZN => n13443);
   U14409 : NAND2_X2 port map( A1 => n20200, A2 => n20201, ZN => n9597);
   U14414 : XOR2_X1 port map( A1 => n25183, A2 => n24936, Z => n2025);
   U14419 : NOR2_X1 port map( A1 => n2423, A2 => n2029, ZN => n17371);
   U14420 : NOR2_X1 port map( A1 => n30302, A2 => n2029, ZN => n25847);
   U14421 : NOR2_X1 port map( A1 => n5356, A2 => n2029, ZN => n4154);
   U14427 : XOR2_X1 port map( A1 => n2032, A2 => n28871, Z => n2031);
   U14429 : XOR2_X1 port map( A1 => n29289, A2 => n28790, Z => n28871);
   U14433 : NOR2_X2 port map( A1 => n16968, A2 => n3093, ZN => n3092);
   U14438 : XOR2_X1 port map( A1 => n35241, A2 => n11755, Z => n2041);
   U14449 : XOR2_X1 port map( A1 => n15202, A2 => n2044, Z => n23739);
   U14452 : NAND2_X1 port map( A1 => n7210, A2 => n24383, ZN => n6570);
   U14460 : XOR2_X1 port map( A1 => n14260, A2 => n29647, Z => n20513);
   U14461 : NOR2_X2 port map( A1 => n21110, A2 => n21109, ZN => n14260);
   U14469 : XOR2_X1 port map( A1 => n37312, A2 => n1559, Z => n2064);
   U14471 : XOR2_X1 port map( A1 => n9939, A2 => n657, Z => n2065);
   U14477 : XOR2_X1 port map( A1 => n31062, A2 => n35238, Z => n2067);
   U14482 : AOI21_X2 port map( A1 => n25924, A2 => n25961, B => n25805, ZN => 
                           n26554);
   U14484 : XOR2_X1 port map( A1 => n2070, A2 => n1367, Z => Ciphertext(119));
   U14486 : XOR2_X1 port map( A1 => n34564, A2 => n19730, Z => n16555);
   U14489 : NAND2_X1 port map( A1 => n1573, A2 => n24812, ZN => n2075);
   U14490 : NAND2_X1 port map( A1 => n24615, A2 => n18983, ZN => n2076);
   U14492 : OAI21_X2 port map( A1 => n31214, A2 => n2233, B => n2082, ZN => 
                           n2234);
   U14493 : AOI21_X2 port map( A1 => n3972, A2 => n22204, B => n3971, ZN => 
                           n2233);
   U14497 : INV_X2 port map( I => n3021, ZN => n18576);
   U14498 : NAND2_X1 port map( A1 => n21820, A2 => n18722, ZN => n2092);
   U14499 : INV_X2 port map( I => n2094, ZN => n18815);
   U14502 : XOR2_X1 port map( A1 => n28835, A2 => n2097, Z => n2096);
   U14503 : XOR2_X1 port map( A1 => n14039, A2 => n19947, Z => n2097);
   U14506 : XOR2_X1 port map( A1 => n542, A2 => n9035, Z => n28834);
   U14513 : AOI21_X2 port map( A1 => n24780, A2 => n24783, B => n17936, ZN => 
                           n25298);
   U14517 : INV_X2 port map( I => n21277, ZN => n26959);
   U14518 : XOR2_X1 port map( A1 => n27690, A2 => n2281, Z => n27756);
   U14523 : XOR2_X1 port map( A1 => n2106, A2 => n2105, Z => n2104);
   U14524 : XOR2_X1 port map( A1 => n23728, A2 => n29522, Z => n2105);
   U14528 : NOR3_X1 port map( A1 => n29683, A2 => n31538, A3 => n38206, ZN => 
                           n2112);
   U14540 : XOR2_X1 port map( A1 => n2122, A2 => n28841, Z => n14438);
   U14551 : XOR2_X1 port map( A1 => n32298, A2 => n29221, Z => n2135);
   U14552 : XOR2_X1 port map( A1 => n33470, A2 => n27862, Z => n2136);
   U14553 : NAND2_X2 port map( A1 => n27375, A2 => n27376, ZN => n27862);
   U14557 : XOR2_X1 port map( A1 => n38144, A2 => n27178, Z => n2138);
   U14568 : NAND2_X1 port map( A1 => n2147, A2 => n28745, ZN => n4024);
   U14584 : XOR2_X1 port map( A1 => n29840, A2 => n4268, Z => n2162);
   U14585 : XOR2_X1 port map( A1 => n29070, A2 => n28948, Z => n29840);
   U14592 : OAI21_X2 port map( A1 => n25430, A2 => n30633, B => n2167, ZN => 
                           n17180);
   U14597 : XOR2_X1 port map( A1 => n24043, A2 => n24042, Z => n2170);
   U14606 : XOR2_X1 port map( A1 => n2177, A2 => n39579, Z => n2176);
   U14607 : XOR2_X1 port map( A1 => n18051, A2 => n2178, Z => n2177);
   U14617 : XOR2_X1 port map( A1 => n25263, A2 => n19359, Z => n2185);
   U14620 : NOR2_X1 port map( A1 => n2187, A2 => n18576, ZN => n2189);
   U14623 : NAND2_X1 port map( A1 => n16237, A2 => n8537, ZN => n16243);
   U14627 : OAI21_X1 port map( A1 => n31875, A2 => n16237, B => n8538, ZN => 
                           n8534);
   U14631 : XOR2_X1 port map( A1 => n36758, A2 => n18180, Z => n2195);
   U14636 : XOR2_X1 port map( A1 => n2199, A2 => n14609, Z => n2198);
   U14637 : XOR2_X1 port map( A1 => n1659, A2 => n4139, Z => n2199);
   U14641 : AOI21_X2 port map( A1 => n22849, A2 => n12925, B => n6018, ZN => 
                           n23200);
   U14643 : NOR2_X1 port map( A1 => n22849, A2 => n36369, ZN => n2202);
   U14644 : XOR2_X1 port map( A1 => n2203, A2 => n19874, Z => Ciphertext(118));
   U14645 : NAND2_X1 port map( A1 => n21018, A2 => n524, ZN => n21017);
   U14647 : XOR2_X1 port map( A1 => n4135, A2 => n2209, Z => n4137);
   U14652 : XOR2_X1 port map( A1 => n2215, A2 => n2214, Z => n20687);
   U14653 : XOR2_X1 port map( A1 => n2978, A2 => n11151, Z => n2214);
   U14659 : XOR2_X1 port map( A1 => n2221, A2 => n32973, Z => n2220);
   U14663 : XOR2_X1 port map( A1 => n24031, A2 => n24032, Z => n2222);
   U14664 : NOR2_X2 port map( A1 => n10109, A2 => n2223, ZN => n24031);
   U14670 : AOI21_X1 port map( A1 => n3697, A2 => n1030, B => n20728, ZN => 
                           n2231);
   U14671 : XOR2_X1 port map( A1 => n8083, A2 => n34553, Z => n2235);
   U14672 : NAND2_X2 port map( A1 => n2707, A2 => n2705, ZN => n8083);
   U14674 : XOR2_X1 port map( A1 => n2234, A2 => n2235, Z => n3999);
   U14675 : INV_X2 port map( I => n8083, ZN => n7287);
   U14682 : NAND2_X2 port map( A1 => n35059, A2 => n26039, ZN => n26214);
   U14689 : XOR2_X1 port map( A1 => n828, A2 => n2263, Z => n15050);
   U14691 : XOR2_X1 port map( A1 => n449, A2 => n29602, Z => n2263);
   U14692 : INV_X2 port map( I => n2264, ZN => n28163);
   U14694 : MUX2_X1 port map( I0 => n4945, I1 => n16363, S => n28163, Z => 
                           n28164);
   U14698 : NAND2_X2 port map( A1 => n2270, A2 => n28308, ZN => n29122);
   U14703 : NAND3_X1 port map( A1 => n23521, A2 => n30835, A3 => n2273, ZN => 
                           n23406);
   U14706 : AOI22_X1 port map( A1 => n21821, A2 => n38246, B1 => n22240, B2 => 
                           n22239, ZN => n19012);
   U14707 : NOR2_X1 port map( A1 => n1349, A2 => n2277, ZN => n2279);
   U14708 : AND2_X1 port map( A1 => n918, A2 => n19388, Z => n2280);
   U14714 : XOR2_X1 port map( A1 => n29066, A2 => n2285, Z => n2284);
   U14715 : XOR2_X1 port map( A1 => n1413, A2 => n19571, Z => n2285);
   U14731 : XOR2_X1 port map( A1 => n2301, A2 => Plaintext(65), Z => n3021);
   U14732 : INV_X1 port map( I => Key(65), ZN => n2301);
   U14736 : INV_X2 port map( I => n2309, ZN => n19966);
   U14742 : XOR2_X1 port map( A1 => n35062, A2 => n23846, Z => n7127);
   U14743 : XOR2_X1 port map( A1 => n24061, A2 => n35062, Z => n23711);
   U14745 : XOR2_X1 port map( A1 => n35062, A2 => n36895, Z => n16004);
   U14754 : AOI21_X1 port map( A1 => n26039, A2 => n31340, B => n20813, ZN => 
                           n2326);
   U14757 : NAND2_X2 port map( A1 => n2328, A2 => n2327, ZN => n28850);
   U14758 : OR2_X1 port map( A1 => n18875, A2 => n31663, Z => n2330);
   U14759 : MUX2_X1 port map( I0 => n28735, I1 => n32682, S => n31554, Z => 
                           n2331);
   U14760 : AOI21_X2 port map( A1 => n28058, A2 => n28057, B => n28056, ZN => 
                           n28735);
   U14766 : INV_X1 port map( I => n11390, ZN => n2335);
   U14773 : NOR2_X1 port map( A1 => n35187, A2 => n10118, ZN => n16275);
   U14776 : OR2_X1 port map( A1 => n10734, A2 => n16792, Z => n15701);
   U14777 : XOR2_X1 port map( A1 => n12200, A2 => n15987, Z => n10734);
   U14784 : XOR2_X1 port map( A1 => n3475, A2 => n37974, Z => n2354);
   U14794 : NAND2_X1 port map( A1 => n38364, A2 => n38013, ZN => n14444);
   U14797 : NOR2_X1 port map( A1 => n10938, A2 => n2366, ZN => n10444);
   U14799 : XOR2_X1 port map( A1 => n23807, A2 => n2367, Z => n3376);
   U14800 : XOR2_X1 port map( A1 => n23910, A2 => n1369, Z => n2367);
   U14803 : OAI21_X2 port map( A1 => n2369, A2 => n17454, B => n2368, ZN => 
                           n5841);
   U14810 : XOR2_X1 port map( A1 => n12430, A2 => n39359, Z => n2371);
   U14819 : NOR2_X2 port map( A1 => n19918, A2 => n7974, ZN => n27027);
   U14820 : NAND2_X2 port map( A1 => n27249, A2 => n7974, ZN => n27250);
   U14821 : NAND2_X1 port map( A1 => n29441, A2 => n29437, ZN => n29423);
   U14822 : XOR2_X1 port map( A1 => n2382, A2 => n2379, Z => n20032);
   U14823 : XOR2_X1 port map( A1 => n35266, A2 => n1698, Z => n2379);
   U14826 : XOR2_X1 port map( A1 => n27850, A2 => n27672, Z => n2382);
   U14830 : XOR2_X1 port map( A1 => n17398, A2 => n2389, Z => n2387);
   U14831 : XOR2_X1 port map( A1 => n19194, A2 => n9271, Z => n2388);
   U14832 : XOR2_X1 port map( A1 => n2390, A2 => n12972, Z => n19194);
   U14833 : XOR2_X1 port map( A1 => n16138, A2 => n19845, Z => n2389);
   U14836 : INV_X2 port map( I => n2391, ZN => n28033);
   U14855 : XOR2_X1 port map( A1 => n23677, A2 => n23891, Z => n2402);
   U14858 : NOR2_X2 port map( A1 => n21557, A2 => n21917, ZN => n21622);
   U14864 : INV_X2 port map( I => n10665, ZN => n25365);
   U14870 : INV_X1 port map( I => n2424, ZN => n26068);
   U14872 : NAND2_X1 port map( A1 => n38914, A2 => n26070, ZN => n25371);
   U14886 : XOR2_X1 port map( A1 => n38219, A2 => n29838, Z => n14772);
   U14888 : XOR2_X1 port map( A1 => n13496, A2 => n38218, Z => n26374);
   U14893 : XOR2_X1 port map( A1 => n24970, A2 => n2446, Z => n2445);
   U14894 : XNOR2_X1 port map( A1 => n20707, A2 => n25163, ZN => n24970);
   U14897 : NAND2_X1 port map( A1 => n9103, A2 => n13433, ZN => n2450);
   U14900 : INV_X2 port map( I => n25636, ZN => n25637);
   U14911 : NOR2_X1 port map( A1 => n2467, A2 => n28128, ZN => n14117);
   U14915 : XOR2_X1 port map( A1 => n20335, A2 => n22790, Z => n22654);
   U14918 : NOR2_X2 port map( A1 => n22024, A2 => n22023, ZN => n22491);
   U14920 : XOR2_X1 port map( A1 => n2476, A2 => n2475, Z => n2474);
   U14921 : XOR2_X1 port map( A1 => n23776, A2 => n1711, Z => n2475);
   U14929 : NAND2_X2 port map( A1 => n2479, A2 => n2478, ZN => n8431);
   U14930 : NAND2_X2 port map( A1 => n2482, A2 => n2481, ZN => n4424);
   U14931 : OAI21_X1 port map( A1 => n16873, A2 => n12109, B => n5733, ZN => 
                           n2482);
   U14933 : XOR2_X1 port map( A1 => n2485, A2 => n1713, Z => Ciphertext(152));
   U14935 : XOR2_X1 port map( A1 => n35404, A2 => n32765, Z => n9695);
   U14937 : XOR2_X1 port map( A1 => n25214, A2 => n32765, Z => n3427);
   U14938 : XOR2_X1 port map( A1 => n32765, A2 => n17395, Z => n10617);
   U14955 : XOR2_X1 port map( A1 => n23865, A2 => n7129, Z => n2510);
   U14956 : XOR2_X1 port map( A1 => n23712, A2 => n3601, Z => n23865);
   U14959 : XOR2_X1 port map( A1 => n20509, A2 => n2656, Z => n7129);
   U14961 : NOR2_X2 port map( A1 => n6911, A2 => n6910, ZN => n2656);
   U14970 : XOR2_X1 port map( A1 => n31537, A2 => n14069, Z => n2515);
   U14972 : XOR2_X1 port map( A1 => n2526, A2 => n2525, Z => n2524);
   U14973 : XOR2_X1 port map( A1 => n24049, A2 => n1370, Z => n2525);
   U14977 : XOR2_X1 port map( A1 => n3609, A2 => n17462, Z => n2529);
   U14980 : XOR2_X1 port map( A1 => n38581, A2 => n31543, Z => n24892);
   U14982 : XOR2_X1 port map( A1 => n35707, A2 => n31543, Z => n13918);
   U14986 : XNOR2_X1 port map( A1 => Plaintext(106), A2 => Key(106), ZN => 
                           n2533);
   U14988 : NAND2_X1 port map( A1 => n11033, A2 => n2534, ZN => n2679);
   U14997 : NAND2_X2 port map( A1 => n16820, A2 => n2537, ZN => n16819);
   U14999 : XOR2_X1 port map( A1 => Plaintext(128), A2 => Key(128), Z => n11702
                           );
   U15001 : XOR2_X1 port map( A1 => n35208, A2 => n37110, Z => n2543);
   U15003 : XOR2_X1 port map( A1 => n871, A2 => n2544, Z => n14174);
   U15004 : XOR2_X1 port map( A1 => n27749, A2 => n19815, Z => n2544);
   U15009 : NAND3_X1 port map( A1 => n30699, A2 => n37983, A3 => n32882, ZN => 
                           n24748);
   U15020 : NAND2_X2 port map( A1 => n939, A2 => n3462, ZN => n11939);
   U15021 : INV_X2 port map( I => n2572, ZN => n20309);
   U15023 : NAND2_X2 port map( A1 => n2667, A2 => n2666, ZN => n6287);
   U15039 : XOR2_X1 port map( A1 => n26491, A2 => n26493, Z => n2592);
   U15043 : XOR2_X1 port map( A1 => n2596, A2 => n18179, Z => n19142);
   U15048 : OAI21_X1 port map( A1 => n2599, A2 => n2601, B => n2598, ZN => 
                           n23219);
   U15055 : XOR2_X1 port map( A1 => n13090, A2 => n5090, Z => n20406);
   U15058 : NAND2_X1 port map( A1 => n24581, A2 => n24904, ZN => n2610);
   U15065 : INV_X2 port map( I => n13207, ZN => n17105);
   U15067 : NAND2_X1 port map( A1 => n17351, A2 => n2616, ZN => n24800);
   U15072 : XOR2_X1 port map( A1 => n25148, A2 => n724, Z => n2622);
   U15075 : XOR2_X1 port map( A1 => n282, A2 => n2627, Z => n6351);
   U15076 : XOR2_X1 port map( A1 => n2627, A2 => n27540, Z => n12495);
   U15077 : XOR2_X1 port map( A1 => n2627, A2 => n19952, Z => n12855);
   U15079 : XOR2_X1 port map( A1 => n2627, A2 => n27802, Z => n27630);
   U15081 : INV_X1 port map( I => n33703, ZN => n23263);
   U15089 : NOR2_X2 port map( A1 => n6636, A2 => n2340, ZN => n10988);
   U15090 : NAND2_X1 port map( A1 => n2634, A2 => n9825, ZN => n24662);
   U15093 : OR2_X1 port map( A1 => n18573, A2 => n1029, Z => n2635);
   U15095 : XOR2_X1 port map( A1 => n28836, A2 => n770, Z => n2637);
   U15100 : XOR2_X1 port map( A1 => n2646, A2 => n2648, Z => n11224);
   U15101 : XOR2_X1 port map( A1 => n26241, A2 => n2647, Z => n2646);
   U15102 : XOR2_X1 port map( A1 => n26439, A2 => n36958, Z => n2647);
   U15103 : XOR2_X1 port map( A1 => n15010, A2 => n2649, Z => n2648);
   U15104 : XOR2_X1 port map( A1 => n9989, A2 => n3413, Z => n2649);
   U15105 : OAI21_X2 port map( A1 => n18273, A2 => n34148, B => n7862, ZN => 
                           n15010);
   U15106 : XOR2_X1 port map( A1 => n2650, A2 => n711, Z => n22897);
   U15108 : XOR2_X1 port map( A1 => n9497, A2 => n2838, Z => n2651);
   U15110 : XOR2_X1 port map( A1 => n2653, A2 => n25290, Z => n25291);
   U15113 : NAND2_X1 port map( A1 => n21982, A2 => n2654, ZN => n3137);
   U15117 : XOR2_X1 port map( A1 => n2656, A2 => n29838, Z => n10402);
   U15118 : XOR2_X1 port map( A1 => n2656, A2 => n19683, Z => n17006);
   U15128 : NOR2_X1 port map( A1 => n7355, A2 => n32434, ZN => n2671);
   U15130 : OAI21_X2 port map( A1 => n2677, A2 => n2674, B => n2675, ZN => 
                           n16502);
   U15131 : AND2_X1 port map( A1 => n24162, A2 => n1603, Z => n2677);
   U15136 : NAND2_X2 port map( A1 => n26447, A2 => n14682, ZN => n27556);
   U15151 : NAND3_X1 port map( A1 => n1337, A2 => n36006, A3 => n32434, ZN => 
                           n22021);
   U15152 : OAI21_X1 port map( A1 => n22019, A2 => n2816, B => n32434, ZN => 
                           n2705);
   U15159 : XOR2_X1 port map( A1 => n2714, A2 => n2713, Z => n2712);
   U15160 : XOR2_X1 port map( A1 => n26531, A2 => n19592, Z => n2713);
   U15165 : NOR2_X1 port map( A1 => n27305, A2 => n34853, ZN => n12427);
   U15171 : XOR2_X1 port map( A1 => n3126, A2 => n2728, Z => n2727);
   U15173 : XOR2_X1 port map( A1 => n37059, A2 => n18430, Z => n2728);
   U15180 : AOI21_X2 port map( A1 => n9580, A2 => n9581, B => n9579, ZN => 
                           n24674);
   U15181 : XOR2_X1 port map( A1 => n22552, A2 => n22743, Z => n18943);
   U15184 : XOR2_X1 port map( A1 => n23894, A2 => n3601, Z => n23663);
   U15191 : XOR2_X1 port map( A1 => n9979, A2 => n23695, Z => n2738);
   U15196 : XOR2_X1 port map( A1 => n15165, A2 => n3110, Z => n11603);
   U15203 : INV_X2 port map( I => n2742, ZN => n8245);
   U15205 : XOR2_X1 port map( A1 => n22438, A2 => n5247, Z => n2743);
   U15212 : XOR2_X1 port map( A1 => n20212, A2 => n14569, Z => n2753);
   U15218 : NOR2_X1 port map( A1 => n4105, A2 => n36840, ZN => n9489);
   U15220 : NAND2_X1 port map( A1 => n9756, A2 => n36840, ZN => n27113);
   U15224 : XOR2_X1 port map( A1 => n27565, A2 => n674, Z => n2757);
   U15225 : XOR2_X1 port map( A1 => n27829, A2 => n27766, Z => n27565);
   U15233 : NOR2_X1 port map( A1 => n34808, A2 => n2765, ZN => n22242);
   U15248 : INV_X2 port map( I => n2778, ZN => n7705);
   U15253 : XOR2_X1 port map( A1 => n2781, A2 => n2780, Z => n22813);
   U15254 : XOR2_X1 port map( A1 => n9206, A2 => n9207, Z => n2780);
   U15258 : NOR2_X2 port map( A1 => n10052, A2 => n17254, ZN => n28722);
   U15269 : XOR2_X1 port map( A1 => n10582, A2 => n25245, Z => n2800);
   U15270 : XOR2_X1 port map( A1 => n27831, A2 => n15736, Z => n2815);
   U15273 : NAND2_X1 port map( A1 => n25484, A2 => n2803, ZN => n25375);
   U15274 : NAND2_X1 port map( A1 => n32904, A2 => n2803, ZN => n25462);
   U15277 : XOR2_X1 port map( A1 => n2806, A2 => n2808, Z => n2805);
   U15279 : XOR2_X1 port map( A1 => n24038, A2 => n23886, Z => n2808);
   U15282 : OAI21_X2 port map( A1 => n2814, A2 => n34245, B => n2813, ZN => 
                           n23894);
   U15283 : INV_X2 port map( I => n2819, ZN => n26863);
   U15290 : XOR2_X1 port map( A1 => n39798, A2 => n39482, Z => n2825);
   U15294 : INV_X2 port map( I => n9133, ZN => n24366);
   U15312 : XOR2_X1 port map( A1 => n26275, A2 => n17428, Z => n2864);
   U15314 : INV_X1 port map( I => n2867, ZN => n5900);
   U15316 : XOR2_X1 port map( A1 => n29964, A2 => n2867, Z => n9270);
   U15317 : XOR2_X1 port map( A1 => n2867, A2 => n27776, Z => n16551);
   U15318 : NAND2_X2 port map( A1 => n3468, A2 => n3467, ZN => n2867);
   U15319 : INV_X2 port map( I => n19888, ZN => n28224);
   U15325 : NAND3_X2 port map( A1 => n2873, A2 => n2874, A3 => n2872, ZN => 
                           n3538);
   U15331 : INV_X2 port map( I => n2881, ZN => n4472);
   U15333 : XOR2_X1 port map( A1 => n3999, A2 => n4000, Z => n2881);
   U15335 : INV_X2 port map( I => n2895, ZN => n24536);
   U15340 : XOR2_X1 port map( A1 => n467, A2 => n29131, Z => n29047);
   U15351 : INV_X2 port map( I => n16704, ZN => n30238);
   U15361 : NAND2_X2 port map( A1 => n2920, A2 => n2919, ZN => n23774);
   U15362 : OAI21_X2 port map( A1 => n19281, A2 => n13262, B => n23086, ZN => 
                           n17017);
   U15369 : XOR2_X1 port map( A1 => n27466, A2 => n29238, Z => n8397);
   U15373 : NAND2_X2 port map( A1 => n14351, A2 => n14352, ZN => n4618);
   U15374 : XOR2_X1 port map( A1 => n25263, A2 => n31568, Z => n13711);
   U15375 : XOR2_X1 port map( A1 => n25182, A2 => n31568, Z => n20805);
   U15377 : XOR2_X1 port map( A1 => n13076, A2 => n2931, Z => n15451);
   U15379 : XOR2_X1 port map( A1 => n23996, A2 => n38880, Z => n9271);
   U15384 : XOR2_X1 port map( A1 => n22648, A2 => n19950, Z => n2935);
   U15388 : NOR2_X2 port map( A1 => n20226, A2 => n20225, ZN => n9878);
   U15390 : AOI21_X1 port map( A1 => n15360, A2 => n32020, B => n27357, ZN => 
                           n21169);
   U15391 : MUX2_X1 port map( I0 => n27066, I1 => n27067, S => n1000, Z => 
                           n27068);
   U15399 : XOR2_X1 port map( A1 => n2943, A2 => n5652, Z => n16587);
   U15400 : XOR2_X1 port map( A1 => n2943, A2 => n28886, Z => n28794);
   U15405 : AOI21_X1 port map( A1 => n2947, A2 => n495, B => n27406, ZN => 
                           n2949);
   U15406 : XNOR2_X1 port map( A1 => n23419, A2 => n23965, ZN => n24026);
   U15410 : AND2_X1 port map( A1 => n13468, A2 => n6894, Z => n2957);
   U15422 : XOR2_X1 port map( A1 => n29142, A2 => n19035, Z => n2978);
   U15424 : XOR2_X1 port map( A1 => n38222, A2 => n31548, Z => n2979);
   U15426 : XOR2_X1 port map( A1 => n3649, A2 => n8447, Z => n3651);
   U15428 : NAND2_X2 port map( A1 => n18571, A2 => n20410, ZN => n3014);
   U15430 : XOR2_X1 port map( A1 => n22699, A2 => n39136, Z => n18834);
   U15432 : XOR2_X1 port map( A1 => n2988, A2 => n2985, Z => n20874);
   U15433 : XOR2_X1 port map( A1 => n2986, A2 => n3953, Z => n2985);
   U15434 : NAND2_X2 port map( A1 => n2987, A2 => n3954, ZN => n3953);
   U15435 : AND2_X1 port map( A1 => n22198, A2 => n22199, Z => n2987);
   U15439 : NAND2_X2 port map( A1 => n5006, A2 => n2991, ZN => n7497);
   U15444 : XOR2_X1 port map( A1 => n28889, A2 => n5862, Z => n29162);
   U15445 : XOR2_X1 port map( A1 => n29164, A2 => n29163, Z => n2996);
   U15450 : XOR2_X1 port map( A1 => n12114, A2 => n12111, Z => n7742);
   U15451 : NAND2_X2 port map( A1 => n15801, A2 => n15804, ZN => n3003);
   U15465 : NOR2_X1 port map( A1 => n22022, A2 => n39010, ZN => n22023);
   U15466 : XOR2_X1 port map( A1 => n22661, A2 => n18888, Z => n3022);
   U15469 : XOR2_X1 port map( A1 => n15311, A2 => n11908, Z => n3023);
   U15474 : OAI21_X2 port map( A1 => n3464, A2 => n29059, B => n3463, ZN => 
                           n3462);
   U15476 : INV_X2 port map( I => n3027, ZN => n22895);
   U15477 : NAND2_X1 port map( A1 => n16104, A2 => n20174, ZN => n22884);
   U15479 : XNOR2_X1 port map( A1 => n35220, A2 => n38201, ZN => n14563);
   U15489 : XOR2_X1 port map( A1 => n3036, A2 => n3037, Z => n3035);
   U15490 : XOR2_X1 port map( A1 => n38844, A2 => n1704, Z => n3036);
   U15491 : XOR2_X1 port map( A1 => n26594, A2 => n10221, Z => n3037);
   U15497 : NAND2_X1 port map( A1 => n3045, A2 => n39828, ZN => n3599);
   U15506 : XOR2_X1 port map( A1 => n3060, A2 => n38189, Z => n29169);
   U15507 : XOR2_X1 port map( A1 => n3082, A2 => n29300, Z => n3060);
   U15514 : OAI21_X2 port map( A1 => n3072, A2 => n1000, B => n3071, ZN => 
                           n27663);
   U15516 : AOI21_X1 port map( A1 => n34952, A2 => n3313, B => n32557, ZN => 
                           n3072);
   U15525 : XOR2_X1 port map( A1 => n10638, A2 => n10635, Z => n12480);
   U15532 : OAI21_X2 port map( A1 => n17531, A2 => n22182, B => n3085, ZN => 
                           n16487);
   U15537 : XOR2_X1 port map( A1 => n27785, A2 => n29785, Z => n3090);
   U15542 : NOR2_X1 port map( A1 => n18257, A2 => n3096, ZN => n20963);
   U15551 : XOR2_X1 port map( A1 => n26194, A2 => n26360, Z => n4022);
   U15554 : XOR2_X1 port map( A1 => n12282, A2 => n3105, Z => n7708);
   U15555 : XOR2_X1 port map( A1 => n22476, A2 => n19866, Z => n3105);
   U15557 : OAI22_X2 port map( A1 => n8549, A2 => n3107, B1 => n8552, B2 => 
                           n3106, ZN => n12282);
   U15564 : AOI21_X1 port map( A1 => n37093, A2 => n31944, B => n38173, ZN => 
                           n20809);
   U15565 : NOR2_X1 port map( A1 => n1642, A2 => n37093, ZN => n15519);
   U15566 : NOR2_X1 port map( A1 => n1633, A2 => n37093, ZN => n21251);
   U15572 : AOI22_X1 port map( A1 => n28708, A2 => n16108, B1 => n18369, B2 => 
                           n28716, ZN => n3128);
   U15573 : OAI21_X2 port map( A1 => n27458, A2 => n36609, B => n3129, ZN => 
                           n28943);
   U15575 : INV_X2 port map( I => n5410, ZN => n20313);
   U15576 : INV_X2 port map( I => n3134, ZN => n26837);
   U15581 : INV_X2 port map( I => n16102, ZN => n18261);
   U15587 : XOR2_X1 port map( A1 => n791, A2 => n3141, Z => n24427);
   U15592 : XOR2_X1 port map( A1 => n38584, A2 => n33515, Z => n3150);
   U15594 : XOR2_X1 port map( A1 => n26595, A2 => n18004, Z => n3152);
   U15599 : AND2_X1 port map( A1 => n5736, A2 => n29182, Z => n3155);
   U15600 : OR2_X1 port map( A1 => n775, A2 => n4095, Z => n3156);
   U15615 : NAND2_X2 port map( A1 => n25441, A2 => n25440, ZN => n18051);
   U15621 : NAND3_X2 port map( A1 => n28173, A2 => n18192, A3 => n3164, ZN => 
                           n28673);
   U15626 : XOR2_X1 port map( A1 => n16523, A2 => n19991, Z => n3166);
   U15629 : XOR2_X1 port map( A1 => n22729, A2 => n29671, Z => n3172);
   U15639 : XOR2_X1 port map( A1 => n27664, A2 => n27663, Z => n27835);
   U15642 : OAI22_X1 port map( A1 => n21826, A2 => n34407, B1 => n21827, B2 => 
                           n3181, ZN => n21828);
   U15644 : INV_X2 port map( I => n21187, ZN => n18104);
   U15647 : XOR2_X1 port map( A1 => n14639, A2 => n25035, Z => n3186);
   U15649 : XOR2_X1 port map( A1 => n15531, A2 => n20069, Z => n3188);
   U15661 : XOR2_X1 port map( A1 => n6560, A2 => n35196, Z => n5915);
   U15662 : XOR2_X1 port map( A1 => n6560, A2 => n23902, Z => n14230);
   U15664 : MUX2_X1 port map( I0 => n1069, I1 => n989, S => n28023, Z => n3199)
                           ;
   U15666 : OAI21_X1 port map( A1 => n1042, A2 => n33817, B => n3200, ZN => 
                           n17202);
   U15671 : XOR2_X1 port map( A1 => n13035, A2 => n27839, Z => n3206);
   U15675 : XOR2_X1 port map( A1 => n27581, A2 => n27580, Z => n27837);
   U15677 : XOR2_X1 port map( A1 => n39093, A2 => n35200, Z => n18106);
   U15678 : XOR2_X1 port map( A1 => n39093, A2 => n12838, Z => n10920);
   U15680 : NAND3_X2 port map( A1 => n24964, A2 => n3214, A3 => n16785, ZN => 
                           n25274);
   U15681 : OAI22_X1 port map( A1 => n3215, A2 => n2277, B1 => n21479, B2 => 
                           n18576, ZN => n21481);
   U15682 : AOI21_X1 port map( A1 => n1349, A2 => n3215, B => n21820, ZN => 
                           n21480);
   U15683 : NAND3_X1 port map( A1 => n6844, A2 => n6845, A3 => n1377, ZN => 
                           n3217);
   U15685 : XOR2_X1 port map( A1 => n35654, A2 => n29983, Z => n17363);
   U15688 : XOR2_X1 port map( A1 => n35867, A2 => n29269, Z => n3223);
   U15692 : XOR2_X1 port map( A1 => n3229, A2 => n4235, Z => n25636);
   U15694 : NAND2_X2 port map( A1 => n8096, A2 => n25358, ZN => n9743);
   U15696 : NOR2_X2 port map( A1 => n5592, A2 => n23313, ZN => n6561);
   U15699 : NAND2_X1 port map( A1 => n13539, A2 => n3235, ZN => n28146);
   U15702 : OAI21_X2 port map( A1 => n1663, A2 => n4139, B => n3237, ZN => 
                           n22663);
   U15707 : XOR2_X1 port map( A1 => n22663, A2 => n8136, Z => n3240);
   U15708 : XOR2_X1 port map( A1 => n3242, A2 => n10718, Z => n3241);
   U15709 : XOR2_X1 port map( A1 => n33690, A2 => n31620, Z => n3242);
   U15710 : AOI21_X2 port map( A1 => n12375, A2 => n16041, B => n12374, ZN => 
                           n10621);
   U15715 : NOR2_X2 port map( A1 => n23468, A2 => n3256, ZN => n23635);
   U15723 : XOR2_X1 port map( A1 => n3262, A2 => n27819, Z => n3261);
   U15724 : NOR2_X2 port map( A1 => n27489, A2 => n27488, ZN => n27819);
   U15725 : XOR2_X1 port map( A1 => n19642, A2 => n1160, Z => n3262);
   U15727 : NAND3_X1 port map( A1 => n29236, A2 => n3263, A3 => n8728, ZN => 
                           n29234);
   U15729 : OAI22_X1 port map( A1 => n14198, A2 => n3263, B1 => n14199, B2 => 
                           n29231, ZN => n14197);
   U15730 : NAND2_X1 port map( A1 => n29230, A2 => n3263, ZN => n15026);
   U15735 : OAI22_X2 port map( A1 => n3271, A2 => n21810, B1 => n3270, B2 => 
                           n19470, ZN => n21214);
   U15739 : XOR2_X1 port map( A1 => n28852, A2 => n3280, Z => n29023);
   U15741 : XOR2_X1 port map( A1 => n3280, A2 => n1374, Z => n29250);
   U15742 : XOR2_X1 port map( A1 => n3280, A2 => n13639, Z => n5648);
   U15747 : INV_X2 port map( I => n14060, ZN => n19914);
   U15751 : XOR2_X1 port map( A1 => n3284, A2 => n14969, Z => Ciphertext(24));
   U15754 : NAND2_X1 port map( A1 => n3288, A2 => n29333, ZN => n3287);
   U15757 : XOR2_X1 port map( A1 => n26393, A2 => n11057, Z => n3290);
   U15758 : XOR2_X1 port map( A1 => n26421, A2 => n26436, Z => n11057);
   U15774 : XOR2_X1 port map( A1 => n7287, A2 => n38920, Z => n3301);
   U15775 : XOR2_X1 port map( A1 => n12437, A2 => n22775, Z => n3303);
   U15776 : XOR2_X1 port map( A1 => n3305, A2 => n16131, Z => n3304);
   U15777 : XOR2_X1 port map( A1 => n15513, A2 => n4139, Z => n3305);
   U15783 : AOI22_X1 port map( A1 => n3312, A2 => n13754, B1 => n27282, B2 => 
                           n3313, ZN => n17697);
   U15784 : NOR2_X1 port map( A1 => n1227, A2 => n3313, ZN => n3312);
   U15786 : NAND2_X2 port map( A1 => n16147, A2 => n9008, ZN => n20333);
   U15789 : XOR2_X1 port map( A1 => n5820, A2 => n23964, Z => n3316);
   U15797 : XOR2_X1 port map( A1 => n26311, A2 => n26232, Z => n3331);
   U15798 : OAI21_X1 port map( A1 => n21574, A2 => n3337, B => n21571, ZN => 
                           n20581);
   U15800 : INV_X1 port map( I => n29023, ZN => n3342);
   U15801 : INV_X2 port map( I => n14834, ZN => n13153);
   U15808 : XOR2_X1 port map( A1 => n11739, A2 => n19879, Z => n3346);
   U15810 : INV_X1 port map( I => n8705, ZN => n3352);
   U15822 : OAI21_X2 port map( A1 => n23318, A2 => n23589, B => n3364, ZN => 
                           n23883);
   U15829 : OAI21_X1 port map( A1 => n34177, A2 => n30141, B => n18588, ZN => 
                           n3373);
   U15831 : XOR2_X1 port map( A1 => n23835, A2 => n16781, Z => n3375);
   U15834 : NAND2_X1 port map( A1 => n6843, A2 => n29278, ZN => n6841);
   U15842 : NOR3_X1 port map( A1 => n34813, A2 => n19873, A3 => n22349, ZN => 
                           n22388);
   U15846 : XOR2_X1 port map( A1 => n57, A2 => n1163, Z => n3387);
   U15847 : NAND2_X1 port map( A1 => n26666, A2 => n3388, ZN => n9646);
   U15848 : NAND2_X1 port map( A1 => n11523, A2 => n3388, ZN => n11522);
   U15849 : XOR2_X1 port map( A1 => n3604, A2 => n8874, Z => n8741);
   U15873 : AOI21_X2 port map( A1 => n3412, A2 => n36662, B => n3409, ZN => 
                           n13733);
   U15875 : MUX2_X1 port map( I0 => n19698, I1 => n4846, S => n13042, Z => 
                           n3412);
   U15878 : AOI21_X2 port map( A1 => n25955, A2 => n365, B => n9589, ZN => 
                           n4828);
   U15880 : XOR2_X1 port map( A1 => n32190, A2 => n18279, Z => n13025);
   U15881 : XOR2_X1 port map( A1 => n23832, A2 => n32190, Z => n13102);
   U15886 : XOR2_X1 port map( A1 => n29098, A2 => n3127, Z => n29100);
   U15892 : XOR2_X1 port map( A1 => Plaintext(187), A2 => Key(187), Z => n3443)
                           ;
   U15896 : XOR2_X1 port map( A1 => n8885, A2 => n26247, Z => n3422);
   U15897 : INV_X2 port map( I => n14122, ZN => n17709);
   U15902 : XOR2_X1 port map( A1 => n3424, A2 => n7329, Z => n15051);
   U15911 : NAND2_X2 port map( A1 => n6214, A2 => n14654, ZN => n17658);
   U15916 : INV_X2 port map( I => n3445, ZN => n5988);
   U15917 : XNOR2_X1 port map( A1 => n3446, A2 => n3603, ZN => n3445);
   U15919 : XOR2_X1 port map( A1 => n27749, A2 => n9981, Z => n3447);
   U15922 : NAND2_X2 port map( A1 => n12269, A2 => n12268, ZN => n3448);
   U15924 : INV_X1 port map( I => Plaintext(191), ZN => n3450);
   U15925 : XOR2_X1 port map( A1 => n3450, A2 => Key(191), Z => n3507);
   U15926 : NAND2_X1 port map( A1 => n3452, A2 => n17464, ZN => n23003);
   U15933 : XOR2_X1 port map( A1 => n3458, A2 => n3457, Z => n3456);
   U15934 : XOR2_X1 port map( A1 => n34768, A2 => n3413, Z => n3457);
   U15935 : XOR2_X1 port map( A1 => n1009, A2 => n26480, Z => n3458);
   U15940 : XOR2_X1 port map( A1 => n3473, A2 => n3472, Z => n3471);
   U15941 : XOR2_X1 port map( A1 => n27796, A2 => n37112, Z => n3472);
   U15942 : XOR2_X1 port map( A1 => n27633, A2 => n8059, Z => n3473);
   U15953 : MUX2_X1 port map( I0 => n19322, I1 => n28571, S => n31513, Z => 
                           n28573);
   U15954 : AOI21_X1 port map( A1 => n37938, A2 => n18854, B => n35290, ZN => 
                           n18952);
   U15958 : INV_X2 port map( I => n3486, ZN => n17993);
   U15961 : NAND2_X1 port map( A1 => n3760, A2 => n30464, ZN => n5401);
   U15964 : XOR2_X1 port map( A1 => n17399, A2 => n3488, Z => n3489);
   U15965 : XOR2_X1 port map( A1 => n29047, A2 => n29046, Z => n3490);
   U15970 : XOR2_X1 port map( A1 => n25240, A2 => n19947, Z => n3493);
   U15979 : NAND2_X2 port map( A1 => n23433, A2 => n23431, ZN => n23624);
   U15981 : NAND2_X2 port map( A1 => n23434, A2 => n23432, ZN => n7335);
   U15982 : INV_X2 port map( I => n3507, ZN => n4116);
   U15986 : NAND2_X1 port map( A1 => n24909, A2 => n3510, ZN => n24729);
   U15992 : NAND3_X2 port map( A1 => n26579, A2 => n26580, A3 => n26581, ZN => 
                           n5831);
   U15995 : AND2_X1 port map( A1 => n26116, A2 => n30302, Z => n3517);
   U15996 : XOR2_X1 port map( A1 => n3521, A2 => n19897, Z => n6781);
   U15998 : XOR2_X1 port map( A1 => n3521, A2 => n19902, Z => n23995);
   U15999 : XOR2_X1 port map( A1 => n3521, A2 => n19887, Z => n15862);
   U16003 : XOR2_X1 port map( A1 => n3523, A2 => n25003, Z => n3522);
   U16004 : XOR2_X1 port map( A1 => n33038, A2 => n31891, Z => n3523);
   U16005 : XNOR2_X1 port map( A1 => n38581, A2 => n25115, ZN => n25003);
   U16006 : XOR2_X1 port map( A1 => n24970, A2 => n4015, Z => n3525);
   U16009 : OAI21_X2 port map( A1 => n33861, A2 => n30196, B => n37083, ZN => 
                           n3527);
   U16011 : INV_X4 port map( I => n20405, ZN => n30196);
   U16015 : NOR2_X1 port map( A1 => n34014, A2 => n3273, ZN => n3546);
   U16016 : INV_X1 port map( I => n13688, ZN => n3547);
   U16017 : XOR2_X1 port map( A1 => n6635, A2 => n3549, Z => n3548);
   U16018 : XOR2_X1 port map( A1 => n29165, A2 => n35249, Z => n3549);
   U16020 : XOR2_X1 port map( A1 => n3552, A2 => n3551, Z => n3550);
   U16023 : XOR2_X1 port map( A1 => n26363, A2 => n3554, Z => n3553);
   U16024 : XOR2_X1 port map( A1 => n18012, A2 => n39082, Z => n3554);
   U16025 : XOR2_X1 port map( A1 => n26587, A2 => n26387, Z => n26363);
   U16026 : NAND2_X2 port map( A1 => n3555, A2 => n26011, ZN => n26387);
   U16027 : NOR2_X2 port map( A1 => n7517, A2 => n26017, ZN => n26587);
   U16041 : XOR2_X1 port map( A1 => Plaintext(99), A2 => Key(99), Z => n3839);
   U16042 : XOR2_X1 port map( A1 => Key(101), A2 => Plaintext(101), Z => n7696)
                           ;
   U16043 : INV_X2 port map( I => n10629, ZN => n21870);
   U16059 : NOR2_X1 port map( A1 => n6390, A2 => n3575, ZN => n6179);
   U16065 : OAI21_X2 port map( A1 => n24209, A2 => n326, B => n23816, ZN => 
                           n8646);
   U16069 : AOI21_X1 port map( A1 => n17618, A2 => n8646, B => n7529, ZN => 
                           n23824);
   U16072 : XOR2_X1 port map( A1 => n25269, A2 => n449, Z => n3576);
   U16073 : XOR2_X1 port map( A1 => n6778, A2 => n3578, Z => n3577);
   U16074 : XOR2_X1 port map( A1 => n25115, A2 => n24944, Z => n3578);
   U16077 : XOR2_X1 port map( A1 => n3585, A2 => n3584, Z => n8765);
   U16078 : XOR2_X1 port map( A1 => n4301, A2 => n698, Z => n3584);
   U16087 : NAND2_X1 port map( A1 => n23529, A2 => n31685, ZN => n6611);
   U16089 : NOR2_X1 port map( A1 => n18883, A2 => n28578, ZN => n14516);
   U16096 : XOR2_X1 port map( A1 => n3601, A2 => n19534, Z => n23984);
   U16097 : XOR2_X1 port map( A1 => n39014, A2 => n19674, Z => n23809);
   U16098 : XOR2_X1 port map( A1 => n39014, A2 => n19903, Z => n23842);
   U16104 : XOR2_X1 port map( A1 => n3604, A2 => n27750, Z => n3603);
   U16107 : NAND2_X1 port map( A1 => n35427, A2 => n11820, ZN => n18488);
   U16110 : NOR2_X1 port map( A1 => n3606, A2 => n13393, ZN => n17024);
   U16111 : NAND2_X1 port map( A1 => n26897, A2 => n3606, ZN => n9203);
   U16114 : XOR2_X1 port map( A1 => n3609, A2 => n19816, Z => n13023);
   U16115 : XOR2_X1 port map( A1 => n3609, A2 => n19843, Z => n23759);
   U16116 : XOR2_X1 port map( A1 => n16858, A2 => n34844, Z => n24015);
   U16117 : XOR2_X1 port map( A1 => n2585, A2 => n29017, Z => n22690);
   U16120 : XOR2_X1 port map( A1 => n23931, A2 => n23609, Z => n3616);
   U16126 : XOR2_X1 port map( A1 => n3621, A2 => n13845, Z => n8694);
   U16128 : XOR2_X1 port map( A1 => n22634, A2 => n3623, Z => n3622);
   U16134 : OAI21_X2 port map( A1 => n3627, A2 => n3626, B => n33821, ZN => 
                           n17904);
   U16135 : XOR2_X1 port map( A1 => n17907, A2 => n17909, Z => n3952);
   U16136 : INV_X2 port map( I => n20482, ZN => n22795);
   U16139 : XOR2_X1 port map( A1 => n28836, A2 => n665, Z => n3632);
   U16141 : INV_X2 port map( I => n11784, ZN => n8527);
   U16143 : XOR2_X1 port map( A1 => n3639, A2 => n13154, Z => n3638);
   U16145 : XOR2_X1 port map( A1 => n26437, A2 => n1506, Z => n3641);
   U16147 : NAND2_X1 port map( A1 => n8393, A2 => n3642, ZN => n8392);
   U16152 : XNOR2_X1 port map( A1 => n19156, A2 => n25030, ZN => n25201);
   U16158 : XOR2_X1 port map( A1 => n3657, A2 => n3651, Z => n3650);
   U16159 : XOR2_X1 port map( A1 => n3656, A2 => n25043, Z => n3652);
   U16160 : XOR2_X1 port map( A1 => n39541, A2 => n19874, Z => n3656);
   U16162 : XOR2_X1 port map( A1 => n26403, A2 => n18432, Z => n15717);
   U16172 : NAND2_X1 port map( A1 => n28654, A2 => n3664, ZN => n28443);
   U16174 : XOR2_X1 port map( A1 => n39798, A2 => n29165, Z => n3666);
   U16184 : XOR2_X1 port map( A1 => n38816, A2 => n29514, Z => n16606);
   U16186 : INV_X2 port map( I => n3675, ZN => n4947);
   U16187 : XOR2_X1 port map( A1 => n1664, A2 => n22604, Z => n4270);
   U16188 : NAND2_X2 port map( A1 => n3679, A2 => n3677, ZN => n10488);
   U16189 : XOR2_X1 port map( A1 => n7848, A2 => n28610, Z => n28959);
   U16197 : OAI21_X1 port map( A1 => n13900, A2 => n11684, B => n3687, ZN => 
                           n11683);
   U16200 : NOR2_X1 port map( A1 => n15996, A2 => n3694, ZN => n20882);
   U16203 : XNOR2_X1 port map( A1 => n22635, A2 => n22619, ZN => n3695);
   U16204 : XOR2_X1 port map( A1 => n19819, A2 => n13564, Z => n22619);
   U16206 : XOR2_X1 port map( A1 => n22760, A2 => n8890, Z => n3696);
   U16211 : NAND2_X1 port map( A1 => n4449, A2 => n3700, ZN => n4448);
   U16213 : XOR2_X1 port map( A1 => n10382, A2 => n14648, Z => n3701);
   U16222 : NOR2_X2 port map( A1 => n18364, A2 => n28518, ZN => n29042);
   U16225 : XOR2_X1 port map( A1 => n9776, A2 => n3711, Z => n3710);
   U16228 : XOR2_X1 port map( A1 => n13155, A2 => n38979, Z => n3712);
   U16232 : INV_X1 port map( I => n30076, ZN => n30081);
   U16233 : NOR2_X1 port map( A1 => n20078, A2 => n30076, ZN => n30060);
   U16235 : NOR2_X2 port map( A1 => n23567, A2 => n23566, ZN => n3715);
   U16238 : NOR2_X1 port map( A1 => n29856, A2 => n3725, ZN => n14160);
   U16241 : XOR2_X1 port map( A1 => n27497, A2 => n3727, Z => n3726);
   U16242 : XOR2_X1 port map( A1 => n27672, A2 => n28831, Z => n3727);
   U16244 : XOR2_X1 port map( A1 => n34829, A2 => n27556, Z => n27673);
   U16248 : XOR2_X1 port map( A1 => n26487, A2 => n39129, Z => n3731);
   U16256 : NOR2_X1 port map( A1 => n19863, A2 => n25498, ZN => n3736);
   U16259 : XOR2_X1 port map( A1 => n25163, A2 => n25096, Z => n24987);
   U16260 : XOR2_X1 port map( A1 => n25163, A2 => n1369, Z => n14687);
   U16263 : XOR2_X1 port map( A1 => n23938, A2 => n9518, Z => n23387);
   U16267 : XOR2_X1 port map( A1 => n12101, A2 => n12282, Z => n3747);
   U16269 : XOR2_X1 port map( A1 => n17651, A2 => n22782, Z => n3748);
   U16270 : OAI21_X2 port map( A1 => n3751, A2 => n24731, B => n3749, ZN => 
                           n15186);
   U16279 : XOR2_X1 port map( A1 => n26522, A2 => n3769, Z => n4412);
   U16280 : XOR2_X1 port map( A1 => n291, A2 => n1723, Z => n3769);
   U16285 : INV_X2 port map( I => n3770, ZN => n16363);
   U16286 : INV_X2 port map( I => n3771, ZN => n4945);
   U16293 : INV_X2 port map( I => n31775, ZN => n3917);
   U16297 : XOR2_X1 port map( A1 => n35320, A2 => n14307, Z => n3776);
   U16298 : XOR2_X1 port map( A1 => n8585, A2 => n30324, Z => n3777);
   U16299 : XOR2_X1 port map( A1 => n38495, A2 => n35251, Z => n3778);
   U16301 : NAND2_X1 port map( A1 => n2302, A2 => n3779, ZN => n12486);
   U16302 : XOR2_X1 port map( A1 => n3780, A2 => n3782, Z => n19436);
   U16304 : NAND2_X2 port map( A1 => n25795, A2 => n25794, ZN => n26396);
   U16306 : NAND2_X2 port map( A1 => n14145, A2 => n25938, ZN => n12649);
   U16307 : XOR2_X1 port map( A1 => n26497, A2 => n30471, Z => n3782);
   U16315 : XOR2_X1 port map( A1 => n33310, A2 => n19925, Z => n3787);
   U16319 : XOR2_X1 port map( A1 => n33584, A2 => n1215, Z => n3790);
   U16320 : XOR2_X1 port map( A1 => n27845, A2 => n31551, Z => n3791);
   U16325 : NOR2_X1 port map( A1 => n28622, A2 => n9917, ZN => n3799);
   U16326 : XOR2_X1 port map( A1 => n3800, A2 => n3801, Z => n12770);
   U16328 : XOR2_X1 port map( A1 => n22689, A2 => n22410, Z => n3801);
   U16330 : NAND2_X2 port map( A1 => n17155, A2 => n17154, ZN => n22775);
   U16331 : INV_X2 port map( I => n26265, ZN => n10440);
   U16337 : XOR2_X1 port map( A1 => n5086, A2 => n3804, Z => n6331);
   U16349 : INV_X1 port map( I => n10029, ZN => n3826);
   U16352 : XOR2_X1 port map( A1 => n15581, A2 => n14969, Z => n11882);
   U16353 : OAI21_X1 port map( A1 => n22299, A2 => n22073, B => n22038, ZN => 
                           n3833);
   U16354 : NAND2_X2 port map( A1 => n33886, A2 => n4388, ZN => n22304);
   U16359 : NAND2_X1 port map( A1 => n39098, A2 => n24764, ZN => n6038);
   U16362 : AOI21_X1 port map( A1 => n36186, A2 => n39098, B => n5896, ZN => 
                           n8579);
   U16364 : OAI21_X1 port map( A1 => n1269, A2 => n39098, B => n4008, ZN => 
                           n7242);
   U16371 : INV_X2 port map( I => n3852, ZN => n8805);
   U16373 : NOR2_X2 port map( A1 => n9016, A2 => n10712, ZN => n11923);
   U16377 : XOR2_X1 port map( A1 => n39698, A2 => n38160, Z => n3855);
   U16380 : OR2_X1 port map( A1 => n3951, A2 => n29182, Z => n3857);
   U16381 : XOR2_X1 port map( A1 => n26408, A2 => n26409, Z => n3858);
   U16383 : NOR2_X1 port map( A1 => n3860, A2 => n31570, ZN => n18083);
   U16384 : NAND2_X1 port map( A1 => n3860, A2 => n39709, ZN => n29913);
   U16387 : OAI21_X1 port map( A1 => n12439, A2 => n7278, B => n3868, ZN => 
                           n3867);
   U16391 : XOR2_X1 port map( A1 => n3929, A2 => n7783, Z => n3872);
   U16396 : AND2_X1 port map( A1 => n19005, A2 => n23381, Z => n3884);
   U16406 : XOR2_X1 port map( A1 => n31620, A2 => n38154, Z => n3891);
   U16409 : XOR2_X1 port map( A1 => n3895, A2 => n3894, Z => n3893);
   U16410 : XOR2_X1 port map( A1 => n9325, A2 => n9324, Z => n3894);
   U16411 : XOR2_X1 port map( A1 => n15186, A2 => n37357, Z => n3895);
   U16413 : NAND2_X2 port map( A1 => n28014, A2 => n28013, ZN => n28570);
   U16418 : XOR2_X1 port map( A1 => n23780, A2 => n3917, Z => n6628);
   U16432 : NAND2_X1 port map( A1 => n9711, A2 => n39489, ZN => n3930);
   U16433 : MUX2_X1 port map( I0 => n6361, I1 => n22069, S => n22327, Z => 
                           n20090);
   U16446 : AOI21_X2 port map( A1 => n14971, A2 => n17190, B => n28754, ZN => 
                           n28852);
   U16447 : XOR2_X1 port map( A1 => n28943, A2 => n19845, Z => n3941);
   U16449 : NOR2_X2 port map( A1 => n34016, A2 => n6241, ZN => n10961);
   U16454 : XNOR2_X1 port map( A1 => n25179, A2 => n20707, ZN => n14644);
   U16457 : XOR2_X1 port map( A1 => n20212, A2 => n11057, Z => n3956);
   U16461 : XOR2_X1 port map( A1 => n2711, A2 => n4258, Z => n4257);
   U16462 : XOR2_X1 port map( A1 => n10653, A2 => n21121, Z => n18893);
   U16464 : XOR2_X1 port map( A1 => n27535, A2 => n10653, Z => n9732);
   U16470 : INV_X2 port map( I => n3973, ZN => n19615);
   U16473 : XOR2_X1 port map( A1 => n11399, A2 => n14293, Z => n3975);
   U16479 : XOR2_X1 port map( A1 => n4273, A2 => n816, Z => n16203);
   U16485 : INV_X2 port map( I => n28174, ZN => n28258);
   U16494 : XOR2_X1 port map( A1 => n8785, A2 => n22505, Z => n4000);
   U16495 : NOR2_X2 port map( A1 => n7041, A2 => n7042, ZN => n4117);
   U16498 : XOR2_X1 port map( A1 => n654, A2 => n27628, Z => n4009);
   U16500 : OR2_X1 port map( A1 => n9334, A2 => n4413, Z => n4010);
   U16502 : NAND3_X2 port map( A1 => n11921, A2 => n22217, A3 => n22218, ZN => 
                           n22615);
   U16506 : XOR2_X1 port map( A1 => n25301, A2 => n29432, Z => n4015);
   U16507 : INV_X2 port map( I => n4016, ZN => n22920);
   U16508 : XOR2_X1 port map( A1 => n14106, A2 => n7593, Z => n15331);
   U16514 : XOR2_X1 port map( A1 => n33308, A2 => n2150, Z => n4021);
   U16518 : XOR2_X1 port map( A1 => n5848, A2 => n39652, Z => n4039);
   U16520 : XOR2_X1 port map( A1 => n29303, A2 => n29934, Z => n4041);
   U16528 : INV_X2 port map( I => n17084, ZN => n24360);
   U16538 : XOR2_X1 port map( A1 => n25330, A2 => n18898, Z => n4061);
   U16542 : XOR2_X1 port map( A1 => n4066, A2 => n4065, Z => n4064);
   U16543 : XOR2_X1 port map( A1 => n27525, A2 => n30207, Z => n4065);
   U16544 : XOR2_X1 port map( A1 => n33584, A2 => n27663, Z => n4066);
   U16554 : XOR2_X1 port map( A1 => n792, A2 => n23940, Z => n4070);
   U16559 : OAI21_X2 port map( A1 => n4429, A2 => n4428, B => n4076, ZN => 
                           n18362);
   U16562 : XOR2_X1 port map( A1 => n39637, A2 => n1357, Z => n4079);
   U16563 : XOR2_X1 port map( A1 => n26571, A2 => n8585, Z => n4080);
   U16569 : XOR2_X1 port map( A1 => n22625, A2 => n22650, Z => n4085);
   U16573 : NOR2_X2 port map( A1 => n10025, A2 => n20042, ZN => n19221);
   U16580 : XOR2_X1 port map( A1 => n32349, A2 => n4092, Z => n4091);
   U16582 : XOR2_X1 port map( A1 => n5026, A2 => n24923, Z => n4090);
   U16585 : XOR2_X1 port map( A1 => n7352, A2 => n15186, Z => n4092);
   U16586 : NOR2_X2 port map( A1 => n23148, A2 => n23147, ZN => n23560);
   U16588 : AOI22_X1 port map( A1 => n19262, A2 => n4093, B1 => n21812, B2 => 
                           n4094, ZN => n18825);
   U16589 : NOR2_X1 port map( A1 => n19768, A2 => n4094, ZN => n4093);
   U16591 : OR2_X1 port map( A1 => n22871, A2 => n19293, Z => n4100);
   U16594 : NOR2_X1 port map( A1 => n38193, A2 => n27253, ZN => n4104);
   U16598 : NAND2_X2 port map( A1 => n4111, A2 => n4109, ZN => n19152);
   U16600 : INV_X1 port map( I => n4108, ZN => n4114);
   U16603 : XOR2_X1 port map( A1 => n20586, A2 => n5185, Z => n23565);
   U16608 : NOR2_X2 port map( A1 => n21374, A2 => n21375, ZN => n22131);
   U16611 : XOR2_X1 port map( A1 => n8875, A2 => n38174, Z => n27750);
   U16619 : XOR2_X1 port map( A1 => n25202, A2 => n24918, Z => n4129);
   U16622 : XOR2_X1 port map( A1 => n5293, A2 => n718, Z => n4131);
   U16626 : XOR2_X1 port map( A1 => n35972, A2 => n19862, Z => n4136);
   U16627 : INV_X2 port map( I => n4137, ZN => n10414);
   U16628 : XOR2_X1 port map( A1 => n4139, A2 => n1356, Z => n4436);
   U16629 : XOR2_X1 port map( A1 => n4441, A2 => n4139, Z => n19956);
   U16630 : XOR2_X1 port map( A1 => n28969, A2 => n29840, Z => n4140);
   U16632 : XOR2_X1 port map( A1 => n11997, A2 => n4142, Z => n11996);
   U16633 : INV_X1 port map( I => n27828, ZN => n4142);
   U16654 : NOR2_X1 port map( A1 => n954, A2 => n728, ZN => n5453);
   U16659 : NAND2_X2 port map( A1 => n17142, A2 => n35500, ZN => n27328);
   U16662 : MUX2_X1 port map( I0 => n24378, I1 => n24377, S => n8041, Z => 
                           n4177);
   U16671 : NOR2_X1 port map( A1 => n17217, A2 => n38377, ZN => n4194);
   U16677 : XOR2_X1 port map( A1 => n4201, A2 => n9027, Z => n9026);
   U16678 : XOR2_X1 port map( A1 => n4201, A2 => n11392, Z => n6906);
   U16683 : XOR2_X1 port map( A1 => n334, A2 => n10027, Z => n4204);
   U16685 : XOR2_X1 port map( A1 => n4205, A2 => n26477, Z => n20536);
   U16689 : NOR2_X1 port map( A1 => n35915, A2 => n31931, ZN => n5723);
   U16693 : NAND3_X1 port map( A1 => n1231, A2 => n33858, A3 => n4211, ZN => 
                           n26964);
   U16696 : NAND2_X1 port map( A1 => n25584, A2 => n25449, ZN => n4214);
   U16700 : XOR2_X1 port map( A1 => n38221, A2 => n4222, Z => n4221);
   U16701 : XOR2_X1 port map( A1 => n7710, A2 => n29325, Z => n4222);
   U16709 : NAND2_X2 port map( A1 => n13073, A2 => n13072, ZN => n13966);
   U16711 : XOR2_X1 port map( A1 => Plaintext(11), A2 => Key(11), Z => n5131);
   U16714 : OAI21_X1 port map( A1 => n18453, A2 => n4232, B => n10544, ZN => 
                           n18398);
   U16715 : NAND3_X1 port map( A1 => n10544, A2 => n18453, A3 => n4232, ZN => 
                           n17045);
   U16720 : XOR2_X1 port map( A1 => n4237, A2 => n25276, Z => n4235);
   U16721 : XOR2_X1 port map( A1 => n18600, A2 => n25275, Z => n4237);
   U16731 : XOR2_X1 port map( A1 => n4256, A2 => n4257, Z => n20995);
   U16733 : XOR2_X1 port map( A1 => n19450, A2 => n19583, Z => n4258);
   U16741 : XOR2_X1 port map( A1 => n16096, A2 => n23591, Z => n4268);
   U16744 : XOR2_X1 port map( A1 => n20668, A2 => n4270, Z => n4269);
   U16745 : XOR2_X1 port map( A1 => n10525, A2 => n22525, Z => n4271);
   U16746 : NAND2_X2 port map( A1 => n22856, A2 => n17080, ZN => n22923);
   U16756 : XOR2_X1 port map( A1 => n22615, A2 => n29920, Z => n4277);
   U16757 : XOR2_X1 port map( A1 => n10558, A2 => n4493, Z => n4278);
   U16765 : XOR2_X1 port map( A1 => n14023, A2 => n9272, Z => n4282);
   U16768 : NAND2_X1 port map( A1 => n14927, A2 => n4283, ZN => n14926);
   U16769 : NAND2_X2 port map( A1 => n22315, A2 => n9616, ZN => n4283);
   U16771 : NOR2_X1 port map( A1 => n35911, A2 => n1414, ZN => n17115);
   U16772 : MUX2_X1 port map( I0 => n28113, I1 => n28112, S => n1414, Z => 
                           n28122);
   U16773 : NAND2_X1 port map( A1 => n32796, A2 => n9677, ZN => n22840);
   U16775 : NAND2_X1 port map( A1 => n31601, A2 => n30096, ZN => n18134);
   U16777 : NOR2_X1 port map( A1 => n9543, A2 => n4294, ZN => n13408);
   U16778 : NAND2_X1 port map( A1 => n33431, A2 => n10334, ZN => n4294);
   U16779 : INV_X2 port map( I => n4300, ZN => n11496);
   U16797 : XOR2_X1 port map( A1 => n29824, A2 => n29785, Z => n4313);
   U16798 : XOR2_X1 port map( A1 => n4314, A2 => n15157, Z => n29129);
   U16806 : OR2_X1 port map( A1 => n16999, A2 => n37067, Z => n4321);
   U16814 : XOR2_X1 port map( A1 => n4327, A2 => n12174, Z => n4326);
   U16815 : NAND2_X2 port map( A1 => n5946, A2 => n4328, ZN => n4644);
   U16816 : OAI21_X1 port map( A1 => n15230, A2 => n22833, B => n11914, ZN => 
                           n4329);
   U16817 : XOR2_X1 port map( A1 => n21098, A2 => n18322, Z => n4330);
   U16819 : XOR2_X1 port map( A1 => n4332, A2 => n4334, Z => n5050);
   U16820 : XOR2_X1 port map( A1 => n24610, A2 => n4333, Z => n4332);
   U16821 : XOR2_X1 port map( A1 => n6066, A2 => n965, Z => n4333);
   U16823 : XOR2_X1 port map( A1 => n25254, A2 => n4335, Z => n4334);
   U16824 : XOR2_X1 port map( A1 => n38665, A2 => n32195, Z => n4335);
   U16826 : NAND2_X1 port map( A1 => n4340, A2 => n1648, ZN => n20971);
   U16830 : INV_X2 port map( I => n4342, ZN => n22335);
   U16831 : XOR2_X1 port map( A1 => n32239, A2 => n19774, Z => n23782);
   U16836 : XOR2_X1 port map( A1 => n22624, A2 => n34239, Z => n4346);
   U16839 : XOR2_X1 port map( A1 => n5566, A2 => n5565, Z => n5402);
   U16840 : INV_X2 port map( I => n4352, ZN => n25601);
   U16842 : NAND2_X2 port map( A1 => n19495, A2 => n25601, ZN => n17613);
   U16845 : NAND3_X1 port map( A1 => n27199, A2 => n13471, A3 => n4353, ZN => 
                           n26915);
   U16848 : XOR2_X1 port map( A1 => n29060, A2 => n4357, Z => n4355);
   U16850 : INV_X2 port map( I => n4356, ZN => n14559);
   U16851 : XOR2_X1 port map( A1 => n15960, A2 => n30682, Z => n4357);
   U16860 : NAND2_X2 port map( A1 => n8169, A2 => n8168, ZN => n9013);
   U16862 : OAI21_X1 port map( A1 => n30181, A2 => n12198, B => n4368, ZN => 
                           n30182);
   U16867 : INV_X2 port map( I => n4386, ZN => n30161);
   U16875 : NOR2_X1 port map( A1 => n28458, A2 => n39423, ZN => n28098);
   U16877 : XOR2_X1 port map( A1 => n4399, A2 => n4398, Z => n4397);
   U16878 : XOR2_X1 port map( A1 => n19561, A2 => n17428, Z => n4398);
   U16879 : XOR2_X1 port map( A1 => n282, A2 => n27504, Z => n4399);
   U16885 : INV_X2 port map( I => n4409, ZN => n13605);
   U16891 : MUX2_X1 port map( I0 => n4417, I1 => n788, S => n1298, Z => n4416);
   U16895 : NAND2_X2 port map( A1 => n15982, A2 => n15985, ZN => n27754);
   U16898 : AOI21_X1 port map( A1 => n6938, A2 => n1399, B => n19050, ZN => 
                           n4423);
   U16899 : INV_X1 port map( I => n4424, ZN => n15663);
   U16901 : NAND2_X1 port map( A1 => n22063, A2 => n4424, ZN => n16499);
   U16913 : XNOR2_X1 port map( A1 => n26514, A2 => n26245, ZN => n26287);
   U16925 : NAND2_X1 port map( A1 => n13982, A2 => n4439, ZN => n23513);
   U16926 : XOR2_X1 port map( A1 => n4440, A2 => n4443, Z => n4442);
   U16927 : XOR2_X1 port map( A1 => n37699, A2 => n1707, Z => n4443);
   U16931 : MUX2_X1 port map( I0 => n28181, I1 => n36573, S => n14397, Z => 
                           n27742);
   U16932 : MUX2_X1 port map( I0 => n1200, I1 => n1074, S => n14397, Z => 
                           n27904);
   U16933 : NOR2_X1 port map( A1 => n4458, A2 => n2752, ZN => n9014);
   U16937 : XOR2_X1 port map( A1 => n38212, A2 => n1362, Z => n15785);
   U16939 : INV_X1 port map( I => n4469, ZN => n25645);
   U16944 : INV_X1 port map( I => n9155, ZN => n8339);
   U16945 : INV_X2 port map( I => n12900, ZN => n14561);
   U16948 : XOR2_X1 port map( A1 => n4477, A2 => n1464, Z => n4476);
   U16949 : XOR2_X1 port map( A1 => n7106, A2 => n19825, Z => n4477);
   U16959 : OAI21_X1 port map( A1 => n30041, A2 => n30042, B => n4498, ZN => 
                           n8477);
   U16961 : XOR2_X1 port map( A1 => n4499, A2 => n4501, Z => n25722);
   U16962 : XOR2_X1 port map( A1 => n25206, A2 => n4500, Z => n4499);
   U16963 : XOR2_X1 port map( A1 => n449, A2 => n30063, Z => n4500);
   U16964 : XOR2_X1 port map( A1 => n25301, A2 => n24984, Z => n25206);
   U16975 : AOI21_X1 port map( A1 => n9559, A2 => n1391, B => n4518, ZN => 
                           n18137);
   U16976 : OAI21_X1 port map( A1 => n29318, A2 => n29333, B => n4519, ZN => 
                           n4518);
   U16988 : XOR2_X1 port map( A1 => n36516, A2 => n12972, Z => n23922);
   U16989 : NAND2_X1 port map( A1 => n8416, A2 => n23414, ZN => n4536);
   U16991 : XOR2_X1 port map( A1 => n360, A2 => n9246, Z => n4540);
   U16994 : XOR2_X1 port map( A1 => n25046, A2 => n4549, Z => n4551);
   U16995 : XOR2_X1 port map( A1 => n16897, A2 => n31771, Z => n4549);
   U16997 : XOR2_X1 port map( A1 => n19967, A2 => n4552, Z => n4550);
   U16999 : XOR2_X1 port map( A1 => n1555, A2 => n3110, Z => n4552);
   U17002 : NAND2_X2 port map( A1 => n19258, A2 => n19257, ZN => n4553);
   U17008 : XOR2_X1 port map( A1 => n38850, A2 => n19534, Z => n4558);
   U17010 : XOR2_X1 port map( A1 => n22637, A2 => n31214, Z => n4559);
   U17014 : XOR2_X1 port map( A1 => n39310, A2 => n30104, Z => n4561);
   U17018 : NAND2_X2 port map( A1 => n5186, A2 => n16393, ZN => n5185);
   U17020 : XOR2_X1 port map( A1 => n4572, A2 => n10230, Z => n9235);
   U17023 : NAND3_X2 port map( A1 => n26104, A2 => n10234, A3 => n26105, ZN => 
                           n26436);
   U17030 : XNOR2_X1 port map( A1 => n778, A2 => n6308, ZN => n4574);
   U17037 : XOR2_X1 port map( A1 => n4591, A2 => n739, Z => n4587);
   U17038 : XOR2_X1 port map( A1 => n11667, A2 => n19516, Z => n4589);
   U17042 : XOR2_X1 port map( A1 => n4592, A2 => n23783, Z => n15160);
   U17052 : XOR2_X1 port map( A1 => n12838, A2 => n8585, Z => n6526);
   U17077 : AOI21_X2 port map( A1 => n4611, A2 => n20971, B => n14544, ZN => 
                           n23307);
   U17084 : NOR2_X2 port map( A1 => n15915, A2 => n27111, ZN => n27478);
   U17095 : INV_X1 port map( I => n19366, ZN => n28147);
   U17099 : OR2_X1 port map( A1 => n29687, A2 => n29678, Z => n29673);
   U17101 : NAND2_X1 port map( A1 => n5357, A2 => n23251, ZN => n19358);
   U17102 : CLKBUF_X2 port map( I => Key(177), Z => n29887);
   U17106 : INV_X2 port map( I => n11782, ZN => n20522);
   U17111 : OAI21_X1 port map( A1 => n15246, A2 => n27506, B => n15243, ZN => 
                           n16861);
   U17114 : INV_X1 port map( I => n20546, ZN => n7468);
   U17119 : NAND2_X1 port map( A1 => n7303, A2 => n38200, ZN => n4621);
   U17124 : NAND2_X2 port map( A1 => n11141, A2 => n11143, ZN => n12015);
   U17128 : OAI21_X2 port map( A1 => n22224, A2 => n22166, B => n13008, ZN => 
                           n22485);
   U17129 : AND2_X1 port map( A1 => n16261, A2 => n1208, Z => n9850);
   U17130 : XOR2_X1 port map( A1 => n29122, A2 => n29072, Z => n28917);
   U17133 : NAND2_X1 port map( A1 => n19060, A2 => n11067, ZN => n4631);
   U17134 : OR2_X1 port map( A1 => n27150, A2 => n27149, Z => n27151);
   U17139 : INV_X2 port map( I => n4632, ZN => n29643);
   U17140 : XOR2_X1 port map( A1 => n27944, A2 => n4834, Z => n4632);
   U17141 : INV_X1 port map( I => n22647, ZN => n7056);
   U17142 : INV_X2 port map( I => n4633, ZN => n20638);
   U17143 : XOR2_X1 port map( A1 => n24935, A2 => n11698, Z => n12181);
   U17149 : XNOR2_X1 port map( A1 => n18765, A2 => n18764, ZN => n5517);
   U17150 : OAI22_X1 port map( A1 => n24720, A2 => n24719, B1 => n30764, B2 => 
                           n24723, ZN => n24726);
   U17151 : XOR2_X1 port map( A1 => n30179, A2 => n16017, Z => n7548);
   U17162 : NAND3_X1 port map( A1 => n20314, A2 => n28331, A3 => n29474, ZN => 
                           n15005);
   U17163 : NAND2_X2 port map( A1 => n10798, A2 => n10799, ZN => n10667);
   U17166 : XOR2_X1 port map( A1 => n5794, A2 => n23378, Z => n5793);
   U17171 : XOR2_X1 port map( A1 => n17552, A2 => n17553, Z => n9748);
   U17174 : XOR2_X1 port map( A1 => n27460, A2 => n1461, Z => n4646);
   U17179 : INV_X1 port map( I => n19088, ZN => n6862);
   U17183 : XOR2_X1 port map( A1 => n5649, A2 => n5651, Z => n28186);
   U17184 : XOR2_X1 port map( A1 => n29085, A2 => n17832, Z => n6855);
   U17185 : OAI21_X2 port map( A1 => n6866, A2 => n17821, B => n6865, ZN => 
                           n16233);
   U17197 : XOR2_X1 port map( A1 => n5889, A2 => n19186, Z => n4658);
   U17199 : AND2_X1 port map( A1 => n18077, A2 => n10004, Z => n17332);
   U17217 : NOR2_X2 port map( A1 => n4670, A2 => n10751, ZN => n24492);
   U17221 : NOR2_X1 port map( A1 => n26847, A2 => n26945, ZN => n15669);
   U17228 : XOR2_X1 port map( A1 => n9776, A2 => n26588, Z => n4673);
   U17238 : NAND2_X1 port map( A1 => n29946, A2 => n105, ZN => n10146);
   U17239 : XNOR2_X1 port map( A1 => n17937, A2 => n30114, ZN => n14053);
   U17246 : XOR2_X1 port map( A1 => n13235, A2 => n5861, Z => n17461);
   U17262 : XNOR2_X1 port map( A1 => n24525, A2 => n24524, ZN => n7957);
   U17268 : OAI21_X1 port map( A1 => n38173, A2 => n15519, B => n23450, ZN => 
                           n22913);
   U17269 : XOR2_X1 port map( A1 => n23954, A2 => n23953, Z => n11575);
   U17277 : NOR2_X2 port map( A1 => n4704, A2 => n22885, ZN => n23296);
   U17278 : XOR2_X1 port map( A1 => n39739, A2 => n29857, Z => n10040);
   U17282 : NAND2_X1 port map( A1 => n22910, A2 => n10828, ZN => n12697);
   U17292 : OR2_X1 port map( A1 => n15320, A2 => n14471, Z => n10937);
   U17293 : AOI21_X2 port map( A1 => n1249, A2 => n20924, B => n4715, ZN => 
                           n25491);
   U17302 : OR2_X1 port map( A1 => n15267, A2 => n9872, Z => n20994);
   U17316 : OAI21_X1 port map( A1 => n19686, A2 => n37757, B => n9856, ZN => 
                           n22823);
   U17319 : XOR2_X1 port map( A1 => n9626, A2 => n29229, Z => n4720);
   U17325 : INV_X1 port map( I => n5762, ZN => n21324);
   U17327 : OR2_X1 port map( A1 => n18815, A2 => n7295, Z => n29187);
   U17334 : OR2_X1 port map( A1 => n26634, A2 => n26905, Z => n26579);
   U17336 : XOR2_X1 port map( A1 => n8703, A2 => n10364, Z => n5583);
   U17337 : AOI21_X1 port map( A1 => n29527, A2 => n29526, B => n4730, ZN => 
                           n29529);
   U17340 : OR2_X1 port map( A1 => n9177, A2 => n25022, Z => n4736);
   U17343 : XOR2_X1 port map( A1 => n19973, A2 => n26314, Z => n9577);
   U17346 : XOR2_X1 port map( A1 => n4738, A2 => n13680, Z => n17918);
   U17350 : XOR2_X1 port map( A1 => n36750, A2 => n19681, Z => n15765);
   U17356 : INV_X2 port map( I => n21074, ZN => n30042);
   U17358 : XOR2_X1 port map( A1 => n4739, A2 => n1730, Z => Ciphertext(123));
   U17371 : NOR2_X1 port map( A1 => n27904, A2 => n18832, ZN => n13976);
   U17377 : NAND3_X1 port map( A1 => n16630, A2 => n16628, A3 => n20499, ZN => 
                           n7589);
   U17380 : XOR2_X1 port map( A1 => n25072, A2 => n6410, Z => n25270);
   U17384 : NAND2_X1 port map( A1 => n13097, A2 => n26956, ZN => n13096);
   U17402 : OR2_X1 port map( A1 => n18168, A2 => n24768, Z => n9418);
   U17404 : XOR2_X1 port map( A1 => n4752, A2 => n27803, Z => n15995);
   U17421 : NAND2_X1 port map( A1 => n2910, A2 => n32107, ZN => n7817);
   U17422 : NAND2_X2 port map( A1 => n8578, A2 => n7971, ZN => n25203);
   U17433 : XOR2_X1 port map( A1 => n17138, A2 => n17139, Z => n28179);
   U17440 : INV_X1 port map( I => n13018, ZN => n20648);
   U17441 : AND2_X1 port map( A1 => n25692, A2 => n12500, Z => n5011);
   U17450 : NAND3_X2 port map( A1 => n22972, A2 => n22970, A3 => n22971, ZN => 
                           n17478);
   U17468 : XOR2_X1 port map( A1 => n4780, A2 => n33515, Z => Ciphertext(179));
   U17470 : XOR2_X1 port map( A1 => n9137, A2 => n779, Z => n4899);
   U17476 : INV_X2 port map( I => n17064, ZN => n20010);
   U17480 : OR2_X1 port map( A1 => n16671, A2 => n24737, Z => n14681);
   U17481 : INV_X2 port map( I => n4786, ZN => n14417);
   U17483 : XOR2_X1 port map( A1 => n13177, A2 => n16310, Z => n13176);
   U17489 : NAND2_X2 port map( A1 => n4897, A2 => n13905, ZN => n15224);
   U17493 : XOR2_X1 port map( A1 => n22454, A2 => n35590, Z => n21134);
   U17494 : NAND2_X2 port map( A1 => n8135, A2 => n16070, ZN => n8585);
   U17499 : AND2_X1 port map( A1 => n30162, A2 => n1400, Z => n17842);
   U17511 : XOR2_X1 port map( A1 => n6642, A2 => n9887, Z => n6641);
   U17512 : NAND2_X2 port map( A1 => n9053, A2 => n11605, ZN => n14425);
   U17513 : NOR2_X1 port map( A1 => n14618, A2 => n6643, ZN => n13620);
   U17517 : AND2_X1 port map( A1 => n3977, A2 => n3092, Z => n11088);
   U17530 : INV_X1 port map( I => n29174, ZN => n30046);
   U17532 : INV_X1 port map( I => n22346, ZN => n13565);
   U17537 : NAND3_X1 port map( A1 => n5110, A2 => n18708, A3 => n10074, ZN => 
                           n16202);
   U17538 : OR2_X1 port map( A1 => n25825, A2 => n18162, Z => n25784);
   U17542 : XOR2_X1 port map( A1 => n11779, A2 => n697, Z => n11778);
   U17551 : NAND3_X2 port map( A1 => n10056, A2 => n24598, A3 => n24599, ZN => 
                           n24991);
   U17566 : XNOR2_X1 port map( A1 => n1065, A2 => n29067, ZN => n9054);
   U17569 : XNOR2_X1 port map( A1 => n27942, A2 => n27943, ZN => n4834);
   U17579 : AND2_X1 port map( A1 => n25539, A2 => n30317, Z => n12908);
   U17584 : NAND2_X1 port map( A1 => n1120, A2 => n24764, ZN => n9417);
   U17590 : INV_X2 port map( I => n4850, ZN => n17424);
   U17597 : NAND3_X1 port map( A1 => n28717, A2 => n28716, A3 => n16108, ZN => 
                           n16505);
   U17598 : OR2_X1 port map( A1 => n5044, A2 => n23542, Z => n6235);
   U17606 : NAND3_X1 port map( A1 => n13586, A2 => n26077, A3 => n9883, ZN => 
                           n13585);
   U17615 : XOR2_X1 port map( A1 => n35376, A2 => n23846, Z => n10888);
   U17616 : NAND2_X2 port map( A1 => n23279, A2 => n15562, ZN => n23846);
   U17618 : AND2_X1 port map( A1 => n906, A2 => n4862, Z => n10018);
   U17627 : INV_X2 port map( I => n4866, ZN => n17412);
   U17628 : XOR2_X1 port map( A1 => n4869, A2 => n11960, Z => n13827);
   U17636 : XOR2_X1 port map( A1 => n4876, A2 => n16641, Z => Ciphertext(82));
   U17637 : NOR3_X1 port map( A1 => n20443, A2 => n21032, A3 => n20444, ZN => 
                           n4876);
   U17649 : XOR2_X1 port map( A1 => n18843, A2 => n22694, Z => n4883);
   U17658 : XOR2_X1 port map( A1 => n17403, A2 => n17402, Z => n14367);
   U17668 : AND2_X1 port map( A1 => n21310, A2 => n19864, Z => n14617);
   U17673 : NOR2_X1 port map( A1 => n5669, A2 => n16704, ZN => n4893);
   U17674 : OAI21_X1 port map( A1 => n13123, A2 => n13771, B => n10190, ZN => 
                           n10189);
   U17677 : AND2_X1 port map( A1 => n19750, A2 => n10836, Z => n10518);
   U17681 : XOR2_X1 port map( A1 => n4894, A2 => n12330, Z => n5080);
   U17682 : OAI21_X1 port map( A1 => n4713, A2 => n12952, B => n4895, ZN => 
                           n16006);
   U17690 : NAND2_X1 port map( A1 => n17202, A2 => n935, ZN => n17201);
   U17691 : OR2_X1 port map( A1 => n28203, A2 => n28001, Z => n4897);
   U17693 : INV_X2 port map( I => n4899, ZN => n20408);
   U17695 : XOR2_X1 port map( A1 => n29027, A2 => n681, Z => n4900);
   U17702 : NAND2_X2 port map( A1 => n4901, A2 => n18108, ZN => n26109);
   U17704 : OR2_X1 port map( A1 => n21989, A2 => n12365, Z => n15652);
   U17706 : XOR2_X1 port map( A1 => n11319, A2 => n16460, Z => n11318);
   U17707 : XNOR2_X1 port map( A1 => n3528, A2 => n17727, ZN => n8785);
   U17711 : XOR2_X1 port map( A1 => n17554, A2 => n9748, Z => n20194);
   U17716 : NAND2_X2 port map( A1 => n28467, A2 => n16840, ZN => n29247);
   U17728 : NAND2_X1 port map( A1 => n6488, A2 => n6489, ZN => n6487);
   U17730 : OR2_X1 port map( A1 => n22783, A2 => n38725, Z => n15375);
   U17731 : OR2_X1 port map( A1 => n20407, A2 => n20408, Z => n13373);
   U17735 : XOR2_X1 port map( A1 => n29837, A2 => n28840, Z => n6536);
   U17742 : NAND2_X1 port map( A1 => n18670, A2 => n29341, ZN => n4919);
   U17745 : AND2_X1 port map( A1 => n12964, A2 => n36006, Z => n5461);
   U17751 : NOR2_X2 port map( A1 => n12537, A2 => n32535, ZN => n11438);
   U17755 : XOR2_X1 port map( A1 => n14955, A2 => n21279, Z => n4929);
   U17772 : XOR2_X1 port map( A1 => n13012, A2 => n13013, Z => n13286);
   U17776 : NAND2_X2 port map( A1 => n4936, A2 => n20302, ZN => n13038);
   U17777 : XOR2_X1 port map( A1 => n26181, A2 => n26182, Z => n17922);
   U17779 : XNOR2_X1 port map( A1 => n22670, A2 => n2383, ZN => n12806);
   U17790 : NOR2_X2 port map( A1 => n11443, A2 => n27010, ZN => n19642);
   U17795 : OR2_X1 port map( A1 => n25327, A2 => n5080, Z => n25535);
   U17798 : NAND3_X2 port map( A1 => n10577, A2 => n10578, A3 => n27106, ZN => 
                           n20976);
   U17800 : NAND2_X1 port map( A1 => n30845, A2 => n7529, ZN => n14276);
   U17802 : INV_X2 port map( I => n21846, ZN => n21672);
   U17807 : OAI21_X1 port map( A1 => n14551, A2 => n18755, B => n21751, ZN => 
                           n10419);
   U17812 : XOR2_X1 port map( A1 => n22699, A2 => n13768, Z => n10382);
   U17813 : NAND2_X2 port map( A1 => n8649, A2 => n22106, ZN => n22699);
   U17816 : AOI21_X1 port map( A1 => n29806, A2 => n29811, B => n39018, ZN => 
                           n5144);
   U17817 : XOR2_X1 port map( A1 => n25029, A2 => n24588, Z => n6109);
   U17823 : XOR2_X1 port map( A1 => n5291, A2 => n4958, Z => n19995);
   U17824 : INV_X1 port map( I => n27538, ZN => n4958);
   U17825 : NOR2_X1 port map( A1 => n11300, A2 => n22856, ZN => n11299);
   U17826 : NOR2_X2 port map( A1 => n24717, A2 => n6944, ZN => n24591);
   U17827 : NOR2_X2 port map( A1 => n6917, A2 => n4959, ZN => n18425);
   U17831 : NAND2_X2 port map( A1 => n13075, A2 => n7884, ZN => n23832);
   U17834 : NAND2_X1 port map( A1 => n11202, A2 => n22008, ZN => n5618);
   U17841 : XOR2_X1 port map( A1 => n21087, A2 => n5742, Z => n4967);
   U17842 : NAND2_X1 port map( A1 => n35506, A2 => n1308, ZN => n4968);
   U17843 : INV_X1 port map( I => n10419, ZN => n10418);
   U17846 : INV_X1 port map( I => n27690, ZN => n15547);
   U17849 : INV_X1 port map( I => n13420, ZN => n13419);
   U17853 : XOR2_X1 port map( A1 => n35303, A2 => n27672, Z => n6026);
   U17856 : NAND2_X2 port map( A1 => n11822, A2 => n4972, ZN => n12028);
   U17860 : XNOR2_X1 port map( A1 => n17567, A2 => n29818, ZN => n5636);
   U17862 : XOR2_X1 port map( A1 => n27692, A2 => n756, Z => n6927);
   U17871 : NOR2_X1 port map( A1 => n6322, A2 => n6321, ZN => n6320);
   U17881 : NAND2_X1 port map( A1 => n9725, A2 => n7537, ZN => n11300);
   U17883 : XOR2_X1 port map( A1 => n26375, A2 => n16046, Z => n26377);
   U17885 : XOR2_X1 port map( A1 => n25180, A2 => n4987, Z => n15517);
   U17886 : XOR2_X1 port map( A1 => n24926, A2 => n19904, Z => n4987);
   U17887 : AND2_X1 port map( A1 => n16250, A2 => n35003, Z => n13885);
   U17890 : XOR2_X1 port map( A1 => n5443, A2 => n23919, Z => n5442);
   U17892 : AOI22_X1 port map( A1 => n13143, A2 => n11981, B1 => n13141, B2 => 
                           n19303, ZN => n13140);
   U17897 : XOR2_X1 port map( A1 => n29096, A2 => n29253, Z => n28767);
   U17901 : XOR2_X1 port map( A1 => n13729, A2 => n16245, Z => n20384);
   U17905 : NAND2_X1 port map( A1 => n19994, A2 => n17644, ZN => n17684);
   U17909 : XOR2_X1 port map( A1 => n29074, A2 => n5648, Z => n4999);
   U17916 : XOR2_X1 port map( A1 => n34009, A2 => n15717, Z => n5003);
   U17923 : NOR2_X2 port map( A1 => n6999, A2 => n6997, ZN => n24829);
   U17928 : AOI21_X2 port map( A1 => n23605, A2 => n23604, B => n23603, ZN => 
                           n23654);
   U17929 : NAND2_X1 port map( A1 => n24232, A2 => n5985, ZN => n6998);
   U17938 : INV_X2 port map( I => n5012, ZN => n11795);
   U17944 : NOR2_X1 port map( A1 => n30059, A2 => n36166, ZN => n21168);
   U17946 : OR2_X1 port map( A1 => n6623, A2 => n29980, Z => n5019);
   U17956 : XOR2_X1 port map( A1 => n29304, A2 => n29305, Z => n14872);
   U17957 : XOR2_X1 port map( A1 => n29113, A2 => n29254, Z => n29305);
   U17963 : NAND2_X2 port map( A1 => n6110, A2 => n27122, ZN => n27786);
   U17966 : XOR2_X1 port map( A1 => n5033, A2 => n24915, Z => n19572);
   U17968 : NAND2_X1 port map( A1 => n32450, A2 => n7467, ZN => n7466);
   U17969 : OAI22_X1 port map( A1 => n9954, A2 => n14390, B1 => n34073, B2 => 
                           n23071, ZN => n16693);
   U17973 : XOR2_X1 port map( A1 => n18094, A2 => n5037, Z => n5525);
   U17974 : XOR2_X1 port map( A1 => n27628, A2 => n27627, Z => n5037);
   U17977 : INV_X1 port map( I => n23686, ZN => n6227);
   U17980 : AND2_X1 port map( A1 => n25851, A2 => n11858, Z => n6399);
   U17984 : XOR2_X1 port map( A1 => n21235, A2 => n5048, Z => n21234);
   U17985 : XOR2_X1 port map( A1 => n18526, A2 => n31515, Z => n5048);
   U17996 : XOR2_X1 port map( A1 => n17195, A2 => n1050, Z => n12598);
   U18003 : OR2_X1 port map( A1 => n8245, A2 => n12631, Z => n7626);
   U18005 : NAND2_X2 port map( A1 => n5054, A2 => n18589, ZN => n20307);
   U18009 : XOR2_X1 port map( A1 => n28946, A2 => n28945, Z => n5587);
   U18013 : XOR2_X1 port map( A1 => n3953, A2 => n17189, Z => n5055);
   U18015 : NAND2_X1 port map( A1 => n9616, A2 => n22155, ZN => n15435);
   U18019 : XOR2_X1 port map( A1 => n8401, A2 => n15197, Z => n5651);
   U18020 : NAND2_X2 port map( A1 => n5623, A2 => n5622, ZN => n8401);
   U18021 : XOR2_X1 port map( A1 => n25253, A2 => n19022, Z => n5058);
   U18028 : AOI21_X2 port map( A1 => n11869, A2 => n19055, B => n11868, ZN => 
                           n11867);
   U18031 : XOR2_X1 port map( A1 => n5065, A2 => n14820, Z => Ciphertext(115));
   U18033 : XOR2_X1 port map( A1 => n15758, A2 => n25178, Z => n17108);
   U18034 : XOR2_X1 port map( A1 => n23965, A2 => n5071, Z => n23966);
   U18035 : XOR2_X1 port map( A1 => n5073, A2 => n19950, Z => Ciphertext(106));
   U18041 : NOR2_X1 port map( A1 => n29719, A2 => n5921, ZN => n16629);
   U18049 : NAND2_X2 port map( A1 => n8961, A2 => n12974, ZN => n13779);
   U18051 : OR2_X1 port map( A1 => n17496, A2 => n16841, Z => n17495);
   U18061 : NAND2_X1 port map( A1 => n5773, A2 => n5772, ZN => n5771);
   U18065 : XOR2_X1 port map( A1 => n5088, A2 => n19845, Z => Ciphertext(19));
   U18070 : XOR2_X1 port map( A1 => n29086, A2 => n13497, Z => n5090);
   U18071 : NAND2_X1 port map( A1 => n8231, A2 => n39083, ZN => n8229);
   U18072 : XOR2_X1 port map( A1 => n7031, A2 => n5091, Z => n28961);
   U18073 : XOR2_X1 port map( A1 => n29026, A2 => n28849, Z => n5091);
   U18077 : XOR2_X1 port map( A1 => n5094, A2 => n23910, Z => n5293);
   U18086 : XOR2_X1 port map( A1 => n16218, A2 => n677, Z => n5096);
   U18091 : OR2_X1 port map( A1 => n31564, A2 => n17790, Z => n23958);
   U18097 : NAND3_X2 port map( A1 => n6521, A2 => n6520, A3 => n9988, ZN => 
                           n6527);
   U18107 : XOR2_X1 port map( A1 => n25164, A2 => n10431, Z => n5114);
   U18112 : XOR2_X1 port map( A1 => n5119, A2 => n5120, Z => n5118);
   U18113 : XOR2_X1 port map( A1 => n26531, A2 => n26305, Z => n5120);
   U18118 : NAND2_X1 port map( A1 => n5126, A2 => n26128, ZN => n25892);
   U18119 : NAND2_X1 port map( A1 => n26126, A2 => n5126, ZN => n5687);
   U18128 : XOR2_X1 port map( A1 => n16781, A2 => n5142, Z => n14258);
   U18129 : XOR2_X1 port map( A1 => n14219, A2 => n23658, Z => n5142);
   U18130 : XOR2_X1 port map( A1 => n5143, A2 => n20781, Z => Ciphertext(108));
   U18132 : XOR2_X1 port map( A1 => n5153, A2 => n28889, Z => n29036);
   U18133 : NOR2_X2 port map( A1 => n5151, A2 => n5150, ZN => n28889);
   U18140 : OAI21_X1 port map( A1 => n27385, A2 => n27064, B => n34562, ZN => 
                           n5167);
   U18141 : XOR2_X1 port map( A1 => n5171, A2 => n13564, Z => n6310);
   U18142 : XOR2_X1 port map( A1 => n5171, A2 => n22598, Z => n13844);
   U18143 : XOR2_X1 port map( A1 => n5171, A2 => n4624, Z => n22686);
   U18152 : XOR2_X1 port map( A1 => n5185, A2 => n14820, Z => n14819);
   U18154 : NAND2_X1 port map( A1 => n5192, A2 => n5188, ZN => Ciphertext(139))
                           ;
   U18155 : NAND2_X1 port map( A1 => n5189, A2 => n5369, ZN => n5188);
   U18156 : NOR2_X1 port map( A1 => n5191, A2 => n5190, ZN => n5189);
   U18157 : NAND2_X1 port map( A1 => n5270, A2 => n30010, ZN => n5190);
   U18158 : NOR2_X1 port map( A1 => n30032, A2 => n39407, ZN => n5191);
   U18159 : NOR3_X1 port map( A1 => n5195, A2 => n5194, A3 => n5193, ZN => 
                           n5192);
   U18160 : NOR2_X1 port map( A1 => n5270, A2 => n30010, ZN => n5193);
   U18161 : NOR3_X1 port map( A1 => n30032, A2 => n39407, A3 => n30010, ZN => 
                           n5195);
   U18164 : INV_X2 port map( I => n11727, ZN => n25727);
   U18166 : OAI22_X2 port map( A1 => n25491, A2 => n14947, B1 => n25142, B2 => 
                           n30470, ZN => n9833);
   U18171 : INV_X2 port map( I => n18707, ZN => n22709);
   U18173 : XOR2_X1 port map( A1 => n28500, A2 => n1160, Z => n28793);
   U18176 : XOR2_X1 port map( A1 => n13853, A2 => n26162, Z => n5226);
   U18177 : XOR2_X1 port map( A1 => n25063, A2 => n5271, Z => n5228);
   U18178 : XNOR2_X1 port map( A1 => n25266, A2 => n25290, ZN => n5271);
   U18180 : XOR2_X1 port map( A1 => n25159, A2 => n813, Z => n5229);
   U18186 : XOR2_X1 port map( A1 => n20353, A2 => n29432, Z => n5235);
   U18188 : XOR2_X1 port map( A1 => n7148, A2 => n30065, Z => n5238);
   U18190 : XOR2_X1 port map( A1 => n5241, A2 => n26325, Z => n8189);
   U18193 : XOR2_X1 port map( A1 => n5242, A2 => n4413, Z => n11967);
   U18194 : XOR2_X1 port map( A1 => n5242, A2 => n29282, Z => n22057);
   U18199 : XOR2_X1 port map( A1 => n19094, A2 => n21048, Z => n5247);
   U18201 : AND2_X1 port map( A1 => n25618, A2 => n19264, Z => n5249);
   U18203 : INV_X1 port map( I => n31767, ZN => n5251);
   U18215 : NAND2_X2 port map( A1 => n9231, A2 => n15643, ZN => n5270);
   U18226 : XOR2_X1 port map( A1 => n19781, A2 => n5285, Z => n19692);
   U18227 : XOR2_X1 port map( A1 => n5286, A2 => n22487, Z => n5285);
   U18228 : XOR2_X1 port map( A1 => n22644, A2 => n5284, Z => n5286);
   U18232 : XOR2_X1 port map( A1 => n6559, A2 => n5290, Z => n18622);
   U18235 : XOR2_X1 port map( A1 => n32464, A2 => n18004, Z => n8780);
   U18238 : NAND3_X1 port map( A1 => n36989, A2 => n6445, A3 => n8137, ZN => 
                           n5295);
   U18242 : INV_X2 port map( I => n19224, ZN => n30153);
   U18254 : XOR2_X1 port map( A1 => n10424, A2 => n9309, Z => n5316);
   U18257 : XOR2_X1 port map( A1 => n5320, A2 => n17859, Z => n5318);
   U18265 : XNOR2_X1 port map( A1 => n5338, A2 => n5339, ZN => n5337);
   U18269 : XOR2_X1 port map( A1 => n5340, A2 => n14530, Z => n5339);
   U18283 : INV_X1 port map( I => n12916, ZN => n5367);
   U18285 : XOR2_X1 port map( A1 => n14333, A2 => Key(71), Z => n21518);
   U18286 : MUX2_X1 port map( I0 => n21039, I1 => n36404, S => n25975, Z => 
                           n16201);
   U18288 : NOR2_X1 port map( A1 => n14838, A2 => n3487, ZN => n10089);
   U18289 : XOR2_X1 port map( A1 => n16524, A2 => n23814, Z => n23676);
   U18291 : XOR2_X1 port map( A1 => n5323, A2 => n29514, Z => n5370);
   U18294 : XOR2_X1 port map( A1 => n27566, A2 => n27767, Z => n27721);
   U18296 : OR2_X1 port map( A1 => n27220, A2 => n37077, Z => n5377);
   U18297 : NOR2_X1 port map( A1 => n3273, A2 => n5380, ZN => n15885);
   U18298 : NAND2_X1 port map( A1 => n5929, A2 => n8882, ZN => n10434);
   U18301 : NAND2_X2 port map( A1 => n23994, A2 => n23993, ZN => n24814);
   U18306 : XOR2_X1 port map( A1 => n5625, A2 => n11755, Z => n5394);
   U18308 : XOR2_X1 port map( A1 => n27716, A2 => n7801, Z => n5395);
   U18316 : XOR2_X1 port map( A1 => n8163, A2 => n1361, Z => n5407);
   U18321 : INV_X2 port map( I => n11543, ZN => n30154);
   U18325 : NAND3_X1 port map( A1 => n30177, A2 => n35899, A3 => n30184, ZN => 
                           n5422);
   U18326 : INV_X1 port map( I => Plaintext(9), ZN => n5423);
   U18327 : XOR2_X1 port map( A1 => n5423, A2 => Key(9), Z => n13397);
   U18331 : AOI21_X1 port map( A1 => n30069, A2 => n30071, B => n30078, ZN => 
                           n20948);
   U18332 : XOR2_X1 port map( A1 => n35215, A2 => n17850, Z => n23920);
   U18333 : XOR2_X1 port map( A1 => n39038, A2 => n19833, Z => n5443);
   U18334 : XOR2_X1 port map( A1 => n20540, A2 => n1096, Z => n26373);
   U18336 : XOR2_X1 port map( A1 => n5447, A2 => n5445, Z => n5444);
   U18337 : XOR2_X1 port map( A1 => n5446, A2 => n26244, Z => n5445);
   U18338 : XOR2_X1 port map( A1 => n26252, A2 => n19866, Z => n5446);
   U18341 : OAI21_X1 port map( A1 => n29338, A2 => n16889, B => n31532, ZN => 
                           n12848);
   U18350 : NOR2_X1 port map( A1 => n28812, A2 => n5465, ZN => n18471);
   U18351 : NAND2_X1 port map( A1 => n28811, A2 => n5465, ZN => n18473);
   U18354 : XOR2_X1 port map( A1 => n39600, A2 => n25074, Z => n5472);
   U18356 : XOR2_X1 port map( A1 => n6352, A2 => n12438, Z => n5473);
   U18365 : XOR2_X1 port map( A1 => n27745, A2 => n29661, Z => n5486);
   U18366 : OAI21_X2 port map( A1 => n21140, A2 => n38305, B => n21139, ZN => 
                           n27745);
   U18367 : INV_X4 port map( I => n23634, ZN => n23468);
   U18368 : OAI21_X2 port map( A1 => n23635, A2 => n5491, B => n5488, ZN => 
                           n24050);
   U18371 : NAND2_X1 port map( A1 => n5798, A2 => n1530, ZN => n15882);
   U18375 : XOR2_X1 port map( A1 => n5510, A2 => n5511, Z => n24104);
   U18379 : XOR2_X1 port map( A1 => n13977, A2 => n23674, Z => n5511);
   U18386 : INV_X1 port map( I => n5709, ZN => n18810);
   U18392 : XOR2_X1 port map( A1 => n35270, A2 => n5524, Z => n5522);
   U18394 : NAND2_X1 port map( A1 => n28286, A2 => n11375, ZN => n6375);
   U18395 : XOR2_X1 port map( A1 => n9030, A2 => n26396, Z => n25853);
   U18396 : XOR2_X1 port map( A1 => n9030, A2 => n19885, Z => n14102);
   U18397 : INV_X1 port map( I => n5527, ZN => n20147);
   U18401 : NOR2_X1 port map( A1 => n5530, A2 => n29284, ZN => n29276);
   U18402 : NOR2_X1 port map( A1 => n37157, A2 => n5530, ZN => n9445);
   U18403 : OAI21_X1 port map( A1 => n18611, A2 => n18610, B => n36676, ZN => 
                           n29280);
   U18406 : XOR2_X1 port map( A1 => n7464, A2 => n8475, Z => n12400);
   U18409 : XOR2_X1 port map( A1 => n5540, A2 => n5538, Z => n13572);
   U18410 : XOR2_X1 port map( A1 => n17413, A2 => n5539, Z => n5538);
   U18411 : XOR2_X1 port map( A1 => n13564, A2 => n29514, Z => n5539);
   U18424 : NAND2_X1 port map( A1 => n36763, A2 => n936, ZN => n23141);
   U18432 : AOI21_X2 port map( A1 => n20504, A2 => n20503, B => n15564, ZN => 
                           n23710);
   U18433 : XOR2_X1 port map( A1 => n5561, A2 => n5562, Z => n5986);
   U18434 : XOR2_X1 port map( A1 => n23756, A2 => n7017, Z => n5561);
   U18435 : XOR2_X1 port map( A1 => n5563, A2 => n23653, Z => n5562);
   U18436 : XOR2_X1 port map( A1 => n8045, A2 => n5564, Z => n5563);
   U18438 : XOR2_X1 port map( A1 => n27713, A2 => n761, Z => n5565);
   U18446 : XOR2_X1 port map( A1 => n22567, A2 => n2383, Z => n17528);
   U18450 : XOR2_X1 port map( A1 => n12464, A2 => n5583, Z => n8943);
   U18452 : XOR2_X1 port map( A1 => n5639, A2 => n18609, Z => n5584);
   U18453 : XOR2_X1 port map( A1 => n10079, A2 => n29050, Z => n5586);
   U18459 : NOR2_X1 port map( A1 => n20924, A2 => n16114, ZN => n5596);
   U18461 : NAND2_X1 port map( A1 => n19587, A2 => n686, ZN => n5598);
   U18462 : XOR2_X1 port map( A1 => n743, A2 => n17680, Z => n5600);
   U18488 : AOI21_X2 port map( A1 => n15651, A2 => n30239, B => n5632, ZN => 
                           n30262);
   U18492 : XOR2_X1 port map( A1 => n5637, A2 => n5636, Z => n5635);
   U18495 : NAND2_X1 port map( A1 => n10836, A2 => n11890, ZN => n27915);
   U18499 : NAND2_X2 port map( A1 => n5930, A2 => n5931, ZN => n5929);
   U18505 : XOR2_X1 port map( A1 => n31550, A2 => n6854, Z => n6853);
   U18506 : XOR2_X1 port map( A1 => n29024, A2 => n5647, Z => n5646);
   U18507 : XOR2_X1 port map( A1 => n29122, A2 => n19897, Z => n5647);
   U18513 : XOR2_X1 port map( A1 => n27781, A2 => n27637, Z => n5650);
   U18516 : XOR2_X1 port map( A1 => n5652, A2 => n29071, Z => n10258);
   U18517 : XOR2_X1 port map( A1 => n5652, A2 => n1165, Z => n17832);
   U18518 : XOR2_X1 port map( A1 => n27823, A2 => n35229, Z => n5655);
   U18519 : INV_X2 port map( I => n5656, ZN => n19469);
   U18526 : XOR2_X1 port map( A1 => n9719, A2 => n1167, Z => n11189);
   U18528 : INV_X1 port map( I => n11166, ZN => n5670);
   U18529 : NAND2_X1 port map( A1 => n28159, A2 => n6548, ZN => n11166);
   U18532 : NAND2_X1 port map( A1 => n1104, A2 => n26055, ZN => n5674);
   U18536 : AOI21_X1 port map( A1 => n29977, A2 => n5678, B => n13705, ZN => 
                           n5677);
   U18537 : OAI21_X1 port map( A1 => n26126, A2 => n15677, B => n5687, ZN => 
                           n5686);
   U18541 : XOR2_X1 port map( A1 => n5692, A2 => n5691, Z => n5690);
   U18544 : XOR2_X1 port map( A1 => n12865, A2 => n18487, Z => n5694);
   U18546 : XOR2_X1 port map( A1 => n1460, A2 => n27676, Z => n5697);
   U18547 : XOR2_X1 port map( A1 => n10370, A2 => n18981, Z => n18980);
   U18549 : XOR2_X1 port map( A1 => n23924, A2 => n5699, Z => n17874);
   U18554 : MUX2_X1 port map( I0 => n27866, I1 => n27928, S => n28193, Z => 
                           n5707);
   U18558 : INV_X2 port map( I => n5717, ZN => n18342);
   U18561 : XOR2_X1 port map( A1 => n6951, A2 => n6952, Z => n5719);
   U18564 : XOR2_X1 port map( A1 => n9567, A2 => n16093, Z => n5722);
   U18568 : XOR2_X1 port map( A1 => n5726, A2 => n5725, Z => n5724);
   U18569 : XOR2_X1 port map( A1 => n29819, A2 => n29818, Z => n5725);
   U18570 : AOI21_X2 port map( A1 => n20951, A2 => n28750, B => n13656, ZN => 
                           n29818);
   U18571 : XOR2_X1 port map( A1 => n38160, A2 => n15617, Z => n5726);
   U18575 : XOR2_X1 port map( A1 => n25247, A2 => n30126, Z => n5730);
   U18577 : XOR2_X1 port map( A1 => n25245, A2 => n11905, Z => n5731);
   U18579 : INV_X1 port map( I => n31528, ZN => n24071);
   U18580 : XOR2_X1 port map( A1 => n15916, A2 => n31528, Z => n7017);
   U18582 : XOR2_X1 port map( A1 => n31528, A2 => n19646, Z => n20045);
   U18584 : XOR2_X1 port map( A1 => n5737, A2 => n12412, Z => n14121);
   U18590 : XOR2_X1 port map( A1 => n29045, A2 => n1163, Z => n14195);
   U18591 : XOR2_X1 port map( A1 => n5741, A2 => n28707, Z => n7665);
   U18592 : XOR2_X1 port map( A1 => n35266, A2 => n29298, Z => n5742);
   U18596 : XOR2_X1 port map( A1 => n15368, A2 => n1214, Z => n5744);
   U18597 : AOI21_X2 port map( A1 => n5748, A2 => n5837, B => n5747, ZN => 
                           n23610);
   U18599 : XOR2_X1 port map( A1 => n5750, A2 => n29506, Z => n18487);
   U18604 : XOR2_X1 port map( A1 => n37044, A2 => n661, Z => n5760);
   U18605 : XOR2_X1 port map( A1 => n24031, A2 => n11267, Z => n5761);
   U18607 : OAI22_X1 port map( A1 => n29869, A2 => n5762, B1 => n20793, B2 => 
                           n4879, ZN => n5971);
   U18609 : XOR2_X1 port map( A1 => n5766, A2 => n5763, Z => n18210);
   U18610 : XOR2_X1 port map( A1 => n5765, A2 => n5764, Z => n5763);
   U18611 : XOR2_X1 port map( A1 => n26402, A2 => n37109, Z => n5764);
   U18614 : XOR2_X1 port map( A1 => n12429, A2 => n26242, Z => n5766);
   U18616 : OAI21_X1 port map( A1 => n1581, A2 => n5768, B => n36395, ZN => 
                           n19836);
   U18618 : OR2_X1 port map( A1 => n27270, A2 => n5772, Z => n5775);
   U18620 : XOR2_X1 port map( A1 => n5778, A2 => n29718, Z => Ciphertext(93));
   U18621 : XOR2_X1 port map( A1 => n28958, A2 => n28959, Z => n5781);
   U18627 : XOR2_X1 port map( A1 => n25257, A2 => n24960, Z => n5789);
   U18628 : AOI21_X2 port map( A1 => n11769, A2 => n11768, B => n17663, ZN => 
                           n6066);
   U18629 : XOR2_X1 port map( A1 => n18427, A2 => n5793, Z => n24202);
   U18630 : INV_X1 port map( I => n23945, ZN => n5794);
   U18631 : XOR2_X1 port map( A1 => n23929, A2 => n24040, Z => n23945);
   U18636 : XOR2_X1 port map( A1 => n17623, A2 => n24962, Z => n5801);
   U18638 : XOR2_X1 port map( A1 => n15288, A2 => n25865, Z => n5803);
   U18640 : XOR2_X1 port map( A1 => n26492, A2 => n26210, Z => n5804);
   U18643 : NAND2_X2 port map( A1 => n5807, A2 => n5805, ZN => n18866);
   U18644 : XOR2_X1 port map( A1 => n5814, A2 => n6112, Z => n5815);
   U18645 : XOR2_X1 port map( A1 => n15186, A2 => n25079, Z => n5814);
   U18653 : AND2_X1 port map( A1 => n22282, A2 => n5819, Z => n6485);
   U18656 : XOR2_X1 port map( A1 => n23873, A2 => n29711, Z => n5820);
   U18657 : OAI21_X2 port map( A1 => n5823, A2 => n526, B => n5822, ZN => n8071
                           );
   U18663 : XOR2_X1 port map( A1 => n5830, A2 => n1554, Z => n5829);
   U18664 : XOR2_X1 port map( A1 => n6759, A2 => n29661, Z => n5830);
   U18672 : NAND2_X2 port map( A1 => n8358, A2 => n8361, ZN => n24764);
   U18674 : XOR2_X1 port map( A1 => n5841, A2 => n15203, Z => n5842);
   U18675 : XOR2_X1 port map( A1 => n23714, A2 => n23883, Z => n24068);
   U18678 : XOR2_X1 port map( A1 => n15531, A2 => n5844, Z => n5843);
   U18679 : XOR2_X1 port map( A1 => n25216, A2 => n19516, Z => n5844);
   U18680 : AOI22_X2 port map( A1 => n21028, A2 => n24749, B1 => n20944, B2 => 
                           n18858, ZN => n25216);
   U18682 : NAND2_X2 port map( A1 => n24965, A2 => n16819, ZN => n24942);
   U18691 : XOR2_X1 port map( A1 => n9719, A2 => n7056, Z => n22516);
   U18692 : XOR2_X1 port map( A1 => n37660, A2 => n1361, Z => n5861);
   U18693 : XOR2_X1 port map( A1 => n5862, A2 => n29034, Z => n28888);
   U18694 : XOR2_X1 port map( A1 => n28982, A2 => n5862, Z => n12561);
   U18697 : AOI21_X2 port map( A1 => n14339, A2 => n11680, B => n7647, ZN => 
                           n5862);
   U18701 : XOR2_X1 port map( A1 => n23686, A2 => n29562, Z => n5866);
   U18704 : XOR2_X1 port map( A1 => n10253, A2 => n10252, Z => n5867);
   U18708 : NAND2_X1 port map( A1 => n5871, A2 => n31679, ZN => n24539);
   U18710 : XOR2_X1 port map( A1 => n27736, A2 => n19874, Z => n5873);
   U18716 : NOR3_X1 port map( A1 => n4674, A2 => n17091, A3 => n36792, ZN => 
                           n25450);
   U18725 : NAND3_X1 port map( A1 => n24709, A2 => n5897, A3 => n34526, ZN => 
                           n7595);
   U18726 : OAI21_X1 port map( A1 => n24708, A2 => n24529, B => n5897, ZN => 
                           n6083);
   U18736 : INV_X2 port map( I => n18186, ZN => n27866);
   U18741 : XOR2_X1 port map( A1 => n360, A2 => n5914, Z => n5913);
   U18744 : XOR2_X1 port map( A1 => n10424, A2 => n723, Z => n5917);
   U18745 : XOR2_X1 port map( A1 => n6896, A2 => n25271, Z => n10424);
   U18747 : XOR2_X1 port map( A1 => n23868, A2 => n5919, Z => n5918);
   U18748 : XOR2_X1 port map( A1 => n23774, A2 => n23686, Z => n5919);
   U18749 : NAND2_X2 port map( A1 => n10208, A2 => n10207, ZN => n19656);
   U18750 : XOR2_X1 port map( A1 => n23740, A2 => n23687, Z => n5920);
   U18756 : NAND2_X1 port map( A1 => n21377, A2 => n21565, ZN => n5931);
   U18760 : XOR2_X1 port map( A1 => n23848, A2 => n16258, Z => n5936);
   U18761 : XOR2_X1 port map( A1 => n24031, A2 => n16257, Z => n5937);
   U18762 : AND2_X1 port map( A1 => n34279, A2 => n31433, Z => n5941);
   U18764 : AOI21_X1 port map( A1 => n17731, A2 => n29719, B => n5921, ZN => 
                           n5949);
   U18768 : OAI21_X1 port map( A1 => n7835, A2 => n1288, B => n5953, ZN => 
                           n24485);
   U18770 : XOR2_X1 port map( A1 => n5956, A2 => n13681, Z => n8812);
   U18771 : XOR2_X1 port map( A1 => n17569, A2 => n22321, Z => n5956);
   U18778 : XOR2_X1 port map( A1 => n10635, A2 => n34848, Z => n5959);
   U18786 : NAND2_X2 port map( A1 => n5969, A2 => n5968, ZN => n20460);
   U18788 : INV_X2 port map( I => n5975, ZN => n19823);
   U18792 : XOR2_X1 port map( A1 => n12863, A2 => n12861, Z => n5974);
   U18801 : NAND3_X2 port map( A1 => n17393, A2 => n17391, A3 => n14457, ZN => 
                           n7611);
   U18802 : INV_X2 port map( I => n5986, ZN => n19915);
   U18807 : XOR2_X1 port map( A1 => n5993, A2 => n5992, Z => n5991);
   U18810 : OAI22_X1 port map( A1 => n33864, A2 => n30299, B1 => n23381, B2 => 
                           n31594, ZN => n5999);
   U18812 : NOR2_X1 port map( A1 => n29220, A2 => n35264, ZN => n13123);
   U18814 : AOI21_X1 port map( A1 => n31772, A2 => n18240, B => n6002, ZN => 
                           n13108);
   U18815 : NOR2_X1 port map( A1 => n10685, A2 => n6002, ZN => n10050);
   U18817 : NAND2_X1 port map( A1 => n13761, A2 => n6002, ZN => n6001);
   U18819 : XOR2_X1 port map( A1 => n26358, A2 => n6008, Z => n6007);
   U18820 : XOR2_X1 port map( A1 => n26596, A2 => n19751, Z => n6008);
   U18821 : NOR3_X1 port map( A1 => n5314, A2 => n10882, A3 => n953, ZN => 
                           n11944);
   U18827 : XOR2_X1 port map( A1 => n5284, A2 => n22743, Z => n7277);
   U18828 : OAI21_X2 port map( A1 => n22305, A2 => n6015, B => n22304, ZN => 
                           n22743);
   U18830 : INV_X2 port map( I => n8694, ZN => n12925);
   U18831 : OR2_X2 port map( A1 => n20649, A2 => n6449, Z => n16468);
   U18832 : NAND2_X1 port map( A1 => n30053, A2 => n6019, ZN => n29180);
   U18834 : XOR2_X1 port map( A1 => n12053, A2 => n6029, Z => n7462);
   U18835 : XOR2_X1 port map( A1 => n7854, A2 => n6030, Z => n6029);
   U18836 : XOR2_X1 port map( A1 => n35240, A2 => n33811, Z => n6030);
   U18842 : XOR2_X1 port map( A1 => n6035, A2 => n22563, Z => n6034);
   U18843 : XOR2_X1 port map( A1 => n22485, A2 => n33661, Z => n6035);
   U18845 : NOR2_X1 port map( A1 => n19089, A2 => n6036, ZN => n13910);
   U18847 : OAI21_X1 port map( A1 => n22156, A2 => n6036, B => n16935, ZN => 
                           n13912);
   U18850 : INV_X4 port map( I => n19604, ZN => n6036);
   U18851 : OAI21_X2 port map( A1 => n15955, A2 => n24094, B => n9909, ZN => 
                           n24878);
   U18856 : INV_X1 port map( I => n4441, ZN => n9074);
   U18857 : XOR2_X1 port map( A1 => n4441, A2 => n4123, Z => n6047);
   U18868 : NAND2_X1 port map( A1 => n23583, A2 => n1626, ZN => n6053);
   U18871 : XOR2_X1 port map( A1 => n6412, A2 => n26206, Z => n6057);
   U18874 : XOR2_X1 port map( A1 => n6066, A2 => n25184, Z => n25042);
   U18886 : INV_X2 port map( I => n7140, ZN => n20931);
   U18887 : XOR2_X1 port map( A1 => n6092, A2 => n6090, Z => n17660);
   U18890 : XOR2_X1 port map( A1 => n19608, A2 => n29554, Z => n6091);
   U18892 : OAI21_X2 port map( A1 => n28531, A2 => n6095, B => n6094, ZN => 
                           n29082);
   U18896 : XOR2_X1 port map( A1 => n12251, A2 => n6108, Z => n6107);
   U18897 : XOR2_X1 port map( A1 => n13917, A2 => n39765, Z => n6108);
   U18899 : XNOR2_X1 port map( A1 => n27786, A2 => n27632, ZN => n16066);
   U18904 : XOR2_X1 port map( A1 => n33921, A2 => n19749, Z => n6112);
   U18905 : NAND2_X1 port map( A1 => n6121, A2 => n6120, ZN => n6126);
   U18909 : NAND2_X1 port map( A1 => n6126, A2 => n6125, ZN => n6124);
   U18911 : NAND3_X1 port map( A1 => n5061, A2 => n6128, A3 => n22248, ZN => 
                           n21739);
   U18914 : XOR2_X1 port map( A1 => n9085, A2 => n6131, Z => n6133);
   U18921 : NOR2_X1 port map( A1 => n35990, A2 => n27267, ZN => n27055);
   U18923 : AOI21_X1 port map( A1 => n27129, A2 => n27128, B => n36177, ZN => 
                           n9727);
   U18924 : NOR2_X1 port map( A1 => n19662, A2 => n35990, ZN => n27130);
   U18925 : XOR2_X1 port map( A1 => n6148, A2 => n19903, Z => Ciphertext(155));
   U18929 : XOR2_X1 port map( A1 => n13961, A2 => n17117, Z => n17060);
   U18933 : NAND2_X2 port map( A1 => n18748, A2 => n19177, ZN => n6159);
   U18934 : XOR2_X1 port map( A1 => Key(131), A2 => Plaintext(131), Z => n6161)
                           ;
   U18935 : INV_X2 port map( I => n6161, ZN => n21308);
   U18938 : NAND2_X1 port map( A1 => n19941, A2 => n25449, ZN => n6172);
   U18940 : XOR2_X1 port map( A1 => n11165, A2 => n11266, Z => n13144);
   U18941 : XOR2_X1 port map( A1 => n6177, A2 => n29298, Z => n20232);
   U18948 : NOR2_X1 port map( A1 => n11126, A2 => n39268, ZN => n6189);
   U18950 : NOR2_X1 port map( A1 => n19951, A2 => n6190, ZN => n10442);
   U18957 : NAND2_X1 port map( A1 => n6198, A2 => n21667, ZN => n6197);
   U18959 : AOI21_X1 port map( A1 => n13574, A2 => n1407, B => n14158, ZN => 
                           n6207);
   U18962 : XOR2_X1 port map( A1 => n6677, A2 => n6212, Z => n6211);
   U18964 : NAND2_X1 port map( A1 => n23528, A2 => n6218, ZN => n23221);
   U18965 : INV_X1 port map( I => n6218, ZN => n6216);
   U18966 : NAND2_X1 port map( A1 => n18086, A2 => n6218, ZN => n20978);
   U18967 : NOR2_X2 port map( A1 => n15588, A2 => n15589, ZN => n6218);
   U18968 : XOR2_X1 port map( A1 => n6224, A2 => n6225, Z => n6223);
   U18970 : XOR2_X1 port map( A1 => n12243, A2 => n19860, Z => n6225);
   U18974 : XOR2_X1 port map( A1 => n6233, A2 => n6231, Z => n25322);
   U18976 : XOR2_X1 port map( A1 => n31579, A2 => n1167, Z => n6232);
   U18983 : NAND2_X1 port map( A1 => n6241, A2 => n261, ZN => n14124);
   U18984 : NAND2_X2 port map( A1 => n17534, A2 => n6241, ZN => n9102);
   U18988 : NOR2_X1 port map( A1 => n39140, A2 => n38198, ZN => n6783);
   U18990 : XOR2_X1 port map( A1 => n6527, A2 => n23776, Z => n23804);
   U18992 : XOR2_X1 port map( A1 => n39231, A2 => n6429, Z => n6428);
   U18993 : XOR2_X1 port map( A1 => n38207, A2 => n1938, Z => n8896);
   U18999 : INV_X2 port map( I => n11084, ZN => n16828);
   U19006 : XOR2_X1 port map( A1 => n22656, A2 => n17428, Z => n12125);
   U19007 : XOR2_X1 port map( A1 => n22656, A2 => n13564, Z => n11289);
   U19017 : INV_X2 port map( I => n21214, ZN => n22146);
   U19023 : XOR2_X1 port map( A1 => n19960, A2 => n6281, Z => n19959);
   U19024 : XOR2_X1 port map( A1 => n23709, A2 => n8929, Z => n6281);
   U19025 : XOR2_X1 port map( A1 => n8447, A2 => n24927, Z => n6283);
   U19027 : OAI22_X2 port map( A1 => n6286, A2 => n39812, B1 => n23553, B2 => 
                           n18747, ZN => n14219);
   U19028 : OAI21_X1 port map( A1 => n6287, A2 => n1420, B => n38155, ZN => 
                           n15964);
   U19031 : XOR2_X1 port map( A1 => n7944, A2 => n29649, Z => n6289);
   U19032 : XOR2_X1 port map( A1 => n26400, A2 => n1509, Z => n26555);
   U19033 : XOR2_X1 port map( A1 => n35239, A2 => n26359, Z => n26400);
   U19035 : XOR2_X1 port map( A1 => n6294, A2 => n20136, Z => n20135);
   U19036 : INV_X1 port map( I => n17493, ZN => n6294);
   U19042 : NAND2_X1 port map( A1 => n26060, A2 => n6302, ZN => n7677);
   U19044 : MUX2_X1 port map( I0 => n18176, I1 => n26063, S => n25943, Z => 
                           n26065);
   U19047 : XOR2_X1 port map( A1 => n6305, A2 => n6306, Z => n6304);
   U19048 : XOR2_X1 port map( A1 => n5021, A2 => n1727, Z => n6305);
   U19050 : XOR2_X1 port map( A1 => n25272, A2 => n19797, Z => n6307);
   U19051 : XOR2_X1 port map( A1 => n6310, A2 => n6309, Z => n6308);
   U19052 : XOR2_X1 port map( A1 => n22620, A2 => n22488, Z => n6309);
   U19056 : INV_X2 port map( I => n18574, ZN => n26893);
   U19063 : XOR2_X1 port map( A1 => n28909, A2 => n6319, Z => n6318);
   U19064 : XOR2_X1 port map( A1 => n10343, A2 => n29849, Z => n6319);
   U19067 : XOR2_X1 port map( A1 => n6320, A2 => n33811, Z => Ciphertext(53));
   U19068 : NAND2_X1 port map( A1 => n9913, A2 => n38200, ZN => n6323);
   U19070 : XOR2_X1 port map( A1 => n6325, A2 => n20047, Z => n6324);
   U19074 : XOR2_X1 port map( A1 => n6329, A2 => n14979, Z => n6328);
   U19076 : INV_X2 port map( I => n6331, ZN => n7834);
   U19082 : NOR2_X1 port map( A1 => n32091, A2 => n6756, ZN => n6706);
   U19085 : NOR2_X1 port map( A1 => n9105, A2 => n9913, ZN => n6339);
   U19087 : NAND2_X2 port map( A1 => n29472, A2 => n29469, ZN => n29477);
   U19088 : NAND2_X1 port map( A1 => n38629, A2 => n34695, ZN => n28112);
   U19092 : XOR2_X1 port map( A1 => n6351, A2 => n16606, Z => n16605);
   U19093 : OAI21_X1 port map( A1 => n39495, A2 => n10211, B => n33148, ZN => 
                           n19169);
   U19094 : XOR2_X1 port map( A1 => n6352, A2 => n24325, Z => n15989);
   U19095 : NOR2_X1 port map( A1 => n6355, A2 => n34969, ZN => n8538);
   U19096 : NAND2_X1 port map( A1 => n6355, A2 => n34969, ZN => n8642);
   U19105 : XOR2_X1 port map( A1 => n23885, A2 => n39161, Z => n6360);
   U19115 : XOR2_X1 port map( A1 => n22542, A2 => n19952, Z => n6368);
   U19116 : XNOR2_X1 port map( A1 => n22488, A2 => n19254, ZN => n22372);
   U19118 : XOR2_X1 port map( A1 => n13564, A2 => n7659, Z => n18153);
   U19127 : AOI21_X2 port map( A1 => n26749, A2 => n11682, B => n6383, ZN => 
                           n13569);
   U19130 : XOR2_X1 port map( A1 => n28850, A2 => n6384, Z => n29031);
   U19131 : XOR2_X1 port map( A1 => n31599, A2 => n19808, Z => n6387);
   U19132 : XOR2_X1 port map( A1 => n6389, A2 => n6467, Z => n20801);
   U19135 : XOR2_X1 port map( A1 => n6395, A2 => n6392, Z => n7281);
   U19136 : XOR2_X1 port map( A1 => n6394, A2 => n6393, Z => n6392);
   U19137 : XOR2_X1 port map( A1 => n27710, A2 => n1707, Z => n6393);
   U19138 : XOR2_X1 port map( A1 => n5625, A2 => n21093, Z => n6394);
   U19142 : NAND3_X2 port map( A1 => n17312, A2 => n6397, A3 => n6396, ZN => 
                           n26519);
   U19143 : OAI21_X2 port map( A1 => n6399, A2 => n17311, B => n6398, ZN => 
                           n26259);
   U19148 : NAND3_X1 port map( A1 => n30078, A2 => n20078, A3 => n3815, ZN => 
                           n30074);
   U19155 : XOR2_X1 port map( A1 => n6413, A2 => n26476, Z => n6412);
   U19164 : AOI21_X2 port map( A1 => n15457, A2 => n19892, B => n33318, ZN => 
                           n10712);
   U19167 : XOR2_X1 port map( A1 => n21108, A2 => n6428, Z => n6427);
   U19169 : XOR2_X1 port map( A1 => n34091, A2 => n29138, Z => n6430);
   U19170 : XOR2_X1 port map( A1 => n6431, A2 => n6432, Z => n6991);
   U19171 : XOR2_X1 port map( A1 => n34829, A2 => n30006, Z => n6431);
   U19172 : XOR2_X1 port map( A1 => n15368, A2 => n13289, Z => n6432);
   U19173 : XOR2_X1 port map( A1 => n6433, A2 => n19761, Z => n29248);
   U19174 : XOR2_X1 port map( A1 => n6433, A2 => n19839, Z => n28785);
   U19176 : XOR2_X1 port map( A1 => n18886, A2 => n769, Z => n6436);
   U19179 : INV_X2 port map( I => n13258, ZN => n7062);
   U19185 : INV_X1 port map( I => Key(134), ZN => n6447);
   U19193 : XOR2_X1 port map( A1 => n26335, A2 => n9554, Z => n6455);
   U19195 : XOR2_X1 port map( A1 => n6458, A2 => n6457, Z => n6456);
   U19199 : XOR2_X1 port map( A1 => n25274, A2 => n6461, Z => n6460);
   U19201 : XOR2_X1 port map( A1 => n23707, A2 => n6462, Z => n6881);
   U19207 : INV_X2 port map( I => n20801, ZN => n24244);
   U19208 : XOR2_X1 port map( A1 => n6468, A2 => n23906, Z => n6467);
   U19212 : XOR2_X1 port map( A1 => n27626, A2 => n6471, Z => n6470);
   U19215 : AOI21_X1 port map( A1 => n6481, A2 => n6480, B => n6479, ZN => 
                           n16249);
   U19216 : NOR3_X1 port map( A1 => n31534, A2 => n29237, A3 => n14933, ZN => 
                           n6479);
   U19217 : OAI21_X1 port map( A1 => n29237, A2 => n1387, B => n1388, ZN => 
                           n6480);
   U19218 : NAND3_X1 port map( A1 => n29228, A2 => n8728, A3 => n38945, ZN => 
                           n6481);
   U19219 : INV_X2 port map( I => n6484, ZN => n19543);
   U19220 : XNOR2_X1 port map( A1 => Plaintext(74), A2 => Key(74), ZN => n6484)
                           ;
   U19221 : NAND2_X2 port map( A1 => n9328, A2 => n9327, ZN => n28768);
   U19223 : NAND2_X1 port map( A1 => n30067, A2 => n31120, ZN => n6486);
   U19226 : NAND2_X2 port map( A1 => n23818, A2 => n13881, ZN => n23796);
   U19229 : INV_X2 port map( I => n6493, ZN => n14562);
   U19232 : NAND2_X2 port map( A1 => n15343, A2 => n6497, ZN => n18762);
   U19235 : INV_X1 port map( I => n19455, ZN => n27276);
   U19236 : NAND2_X1 port map( A1 => n20027, A2 => n37480, ZN => n6509);
   U19239 : XOR2_X1 port map( A1 => n22597, A2 => n6512, Z => n6511);
   U19240 : XOR2_X1 port map( A1 => n12243, A2 => n19905, Z => n6512);
   U19241 : XOR2_X1 port map( A1 => n22658, A2 => n18634, Z => n6513);
   U19242 : XOR2_X1 port map( A1 => n11541, A2 => n5203, Z => n22658);
   U19246 : XOR2_X1 port map( A1 => n12839, A2 => n18296, Z => n6525);
   U19248 : XOR2_X1 port map( A1 => n6530, A2 => n6528, Z => n19576);
   U19250 : XOR2_X1 port map( A1 => n23794, A2 => n1699, Z => n6531);
   U19252 : XOR2_X1 port map( A1 => n6536, A2 => n28820, Z => n6535);
   U19256 : NAND2_X2 port map( A1 => n24717, A2 => n6944, ZN => n24724);
   U19257 : NOR2_X2 port map( A1 => n6543, A2 => n19580, ZN => n25862);
   U19259 : XOR2_X1 port map( A1 => n10705, A2 => n22448, Z => n6544);
   U19260 : XOR2_X1 port map( A1 => n57, A2 => n22784, Z => n22448);
   U19267 : XOR2_X1 port map( A1 => n27413, A2 => n11365, Z => n6549);
   U19274 : XOR2_X1 port map( A1 => n6562, A2 => n6563, Z => n18602);
   U19275 : XOR2_X1 port map( A1 => n31581, A2 => n23785, Z => n6562);
   U19276 : XOR2_X1 port map( A1 => n23316, A2 => n6564, Z => n6563);
   U19285 : XOR2_X1 port map( A1 => n6817, A2 => n6580, Z => n6581);
   U19286 : XOR2_X1 port map( A1 => n6633, A2 => n6632, Z => n6580);
   U19287 : XOR2_X1 port map( A1 => n6630, A2 => n17513, Z => n6817);
   U19292 : OAI21_X2 port map( A1 => n14665, A2 => n15702, B => n14012, ZN => 
                           n10635);
   U19294 : NAND2_X2 port map( A1 => n6587, A2 => n6586, ZN => n28807);
   U19295 : NAND2_X1 port map( A1 => n28288, A2 => n11375, ZN => n6586);
   U19296 : NAND2_X1 port map( A1 => n6590, A2 => n13712, ZN => n25970);
   U19304 : XOR2_X1 port map( A1 => n13919, A2 => n13918, Z => n6595);
   U19310 : OAI21_X1 port map( A1 => n6600, A2 => n11861, B => n16510, ZN => 
                           n6599);
   U19316 : XOR2_X1 port map( A1 => n22442, A2 => n6609, Z => n6608);
   U19317 : XOR2_X1 port map( A1 => n11201, A2 => n1661, Z => n6609);
   U19321 : XOR2_X1 port map( A1 => n22484, A2 => n22459, Z => n22441);
   U19326 : INV_X1 port map( I => n26088, ZN => n20545);
   U19328 : AOI21_X1 port map( A1 => n29979, A2 => n29980, B => n6623, ZN => 
                           n18200);
   U19331 : NAND2_X1 port map( A1 => n6623, A2 => n29979, ZN => n6622);
   U19332 : NAND2_X2 port map( A1 => n17983, A2 => n29961, ZN => n6623);
   U19333 : XOR2_X1 port map( A1 => n6624, A2 => n6627, Z => n7364);
   U19334 : XOR2_X1 port map( A1 => n24013, A2 => n6625, Z => n6624);
   U19335 : XOR2_X1 port map( A1 => n24079, A2 => n6626, Z => n6625);
   U19337 : XOR2_X1 port map( A1 => n6628, A2 => n19623, Z => n6627);
   U19338 : OR2_X1 port map( A1 => n6629, A2 => n8082, Z => n6697);
   U19343 : XOR2_X1 port map( A1 => n17189, A2 => n22508, Z => n6632);
   U19345 : NAND2_X1 port map( A1 => n6772, A2 => n6771, ZN => n6634);
   U19347 : NOR2_X2 port map( A1 => n10648, A2 => n10988, ZN => n10987);
   U19349 : XOR2_X1 port map( A1 => n6644, A2 => n16886, Z => n19855);
   U19355 : OAI21_X1 port map( A1 => n10096, A2 => n29870, B => n20793, ZN => 
                           n20895);
   U19360 : MUX2_X1 port map( I0 => n841, I1 => n6656, S => n25669, Z => n19971
                           );
   U19365 : NOR3_X1 port map( A1 => n38529, A2 => n28695, A3 => n28696, ZN => 
                           n10680);
   U19367 : NAND2_X2 port map( A1 => n10304, A2 => n10302, ZN => n29054);
   U19373 : OR2_X1 port map( A1 => n1486, A2 => n34001, Z => n6668);
   U19382 : XOR2_X1 port map( A1 => n12101, A2 => n6676, Z => n9595);
   U19383 : XOR2_X1 port map( A1 => n22703, A2 => n19676, Z => n6676);
   U19385 : XOR2_X1 port map( A1 => n2281, A2 => n27736, Z => n6677);
   U19395 : INV_X2 port map( I => n4378, ZN => n30071);
   U19397 : XOR2_X1 port map( A1 => n10653, A2 => n1738, Z => n6688);
   U19401 : XOR2_X1 port map( A1 => n12763, A2 => n10059, Z => n16217);
   U19402 : INV_X2 port map( I => n8532, ZN => n16639);
   U19404 : INV_X1 port map( I => n8082, ZN => n6698);
   U19409 : XOR2_X1 port map( A1 => n22634, A2 => n5203, Z => n6711);
   U19411 : NAND2_X2 port map( A1 => n1275, A2 => n39699, ZN => n6715);
   U19412 : XOR2_X1 port map( A1 => n8402, A2 => n11755, Z => n6717);
   U19417 : XOR2_X1 port map( A1 => n38161, A2 => n29394, Z => n28372);
   U19418 : XOR2_X1 port map( A1 => n30856, A2 => n38161, Z => n29138);
   U19424 : XOR2_X1 port map( A1 => n26370, A2 => n26323, Z => n12228);
   U19429 : AOI21_X2 port map( A1 => n27297, A2 => n35473, B => n27296, ZN => 
                           n27525);
   U19431 : XOR2_X1 port map( A1 => n25153, A2 => n20803, Z => n6728);
   U19433 : XOR2_X1 port map( A1 => n25152, A2 => n20805, Z => n6729);
   U19437 : OAI21_X1 port map( A1 => n21654, A2 => n33771, B => n6732, ZN => 
                           n11849);
   U19447 : XOR2_X1 port map( A1 => n26510, A2 => n36579, Z => n26172);
   U19449 : XOR2_X1 port map( A1 => n26233, A2 => n25930, Z => n6739);
   U19450 : XOR2_X1 port map( A1 => n26157, A2 => n26389, Z => n26233);
   U19452 : XOR2_X1 port map( A1 => n16254, A2 => n22693, Z => n6741);
   U19460 : XOR2_X1 port map( A1 => n16066, A2 => n6752, Z => n6751);
   U19461 : XOR2_X1 port map( A1 => n27729, A2 => n37101, Z => n6752);
   U19462 : XOR2_X1 port map( A1 => n27515, A2 => n10766, Z => n6753);
   U19463 : XOR2_X1 port map( A1 => n5284, A2 => n19904, Z => n18843);
   U19464 : XOR2_X1 port map( A1 => n6014, A2 => n29649, Z => n18941);
   U19465 : XOR2_X1 port map( A1 => n5284, A2 => n19677, Z => n22427);
   U19466 : NAND3_X1 port map( A1 => n36376, A2 => n36920, A3 => n38884, ZN => 
                           n8109);
   U19468 : XOR2_X1 port map( A1 => n6757, A2 => n19877, Z => n25865);
   U19470 : XOR2_X1 port map( A1 => n38584, A2 => n6757, Z => n13814);
   U19472 : XOR2_X1 port map( A1 => n38195, A2 => n19874, Z => n28306);
   U19474 : XOR2_X1 port map( A1 => n19725, A2 => n61, Z => n25075);
   U19479 : XOR2_X1 port map( A1 => n6765, A2 => n34815, Z => n6764);
   U19480 : XOR2_X1 port map( A1 => n1613, A2 => n23900, Z => n6765);
   U19490 : NAND3_X1 port map( A1 => n12567, A2 => n22162, A3 => n19890, ZN => 
                           n6771);
   U19491 : INV_X1 port map( I => n6773, ZN => n6772);
   U19493 : INV_X2 port map( I => n29943, ZN => n16353);
   U19495 : NOR2_X1 port map( A1 => n6776, A2 => n9727, ZN => n6775);
   U19501 : XOR2_X1 port map( A1 => n35379, A2 => n19875, Z => n6778);
   U19502 : XOR2_X1 port map( A1 => n6782, A2 => n6781, Z => n6780);
   U19503 : XOR2_X1 port map( A1 => n6527, A2 => n23829, Z => n6782);
   U19507 : XOR2_X1 port map( A1 => n22689, A2 => n2234, Z => n7346);
   U19509 : INV_X2 port map( I => n6801, ZN => n12162);
   U19510 : XOR2_X1 port map( A1 => n24946, A2 => n11689, Z => n6802);
   U19516 : XOR2_X1 port map( A1 => n7352, A2 => n25123, Z => n25011);
   U19518 : NOR2_X1 port map( A1 => n23502, A2 => n32366, ZN => n23048);
   U19521 : OAI21_X2 port map( A1 => n19104, A2 => n21622, B => n18900, ZN => 
                           n22364);
   U19527 : XOR2_X1 port map( A1 => Plaintext(21), A2 => Key(21), Z => n8267);
   U19531 : XOR2_X1 port map( A1 => n12442, A2 => n15158, Z => n6825);
   U19538 : XOR2_X1 port map( A1 => n6835, A2 => n6834, Z => n6836);
   U19540 : INV_X2 port map( I => n6836, ZN => n30055);
   U19542 : INV_X1 port map( I => n9310, ZN => n27271);
   U19545 : XOR2_X1 port map( A1 => n12730, A2 => n31562, Z => n11908);
   U19546 : XOR2_X1 port map( A1 => n31562, A2 => n1718, Z => n16753);
   U19547 : XOR2_X1 port map( A1 => n31562, A2 => n19761, Z => n13846);
   U19552 : NAND2_X1 port map( A1 => n6851, A2 => n20018, ZN => n12994);
   U19554 : OAI21_X1 port map( A1 => n18461, A2 => n13153, B => n6851, ZN => 
                           n16121);
   U19556 : XOR2_X1 port map( A1 => n29031, A2 => n6853, Z => n6852);
   U19568 : INV_X1 port map( I => n34001, ZN => n27196);
   U19570 : NAND2_X1 port map( A1 => n27368, A2 => n5772, ZN => n6874);
   U19571 : XOR2_X1 port map( A1 => n6879, A2 => n6878, Z => n6877);
   U19572 : XOR2_X1 port map( A1 => n26234, A2 => n1362, Z => n6878);
   U19573 : XOR2_X1 port map( A1 => n208, A2 => n6881, Z => n6880);
   U19577 : NAND2_X1 port map( A1 => n31533, A2 => n16803, ZN => n10294);
   U19578 : NAND2_X1 port map( A1 => n31533, A2 => n967, ZN => n17885);
   U19580 : XOR2_X1 port map( A1 => n6886, A2 => n12076, Z => n8069);
   U19581 : XOR2_X1 port map( A1 => n25126, A2 => n6887, Z => n6886);
   U19582 : XOR2_X1 port map( A1 => n25080, A2 => n19733, Z => n6887);
   U19583 : XOR2_X1 port map( A1 => n25259, A2 => n25216, Z => n25126);
   U19585 : NAND2_X2 port map( A1 => n10826, A2 => n10824, ZN => n6892);
   U19588 : XOR2_X1 port map( A1 => n35112, A2 => n22615, Z => n22479);
   U19591 : XOR2_X1 port map( A1 => n10424, A2 => n6895, Z => n9808);
   U19592 : XOR2_X1 port map( A1 => n35053, A2 => n1697, Z => n6895);
   U19598 : XOR2_X1 port map( A1 => n7416, A2 => n11391, Z => n6905);
   U19602 : NAND2_X1 port map( A1 => n6908, A2 => n27389, ZN => n26428);
   U19611 : XOR2_X1 port map( A1 => n6923, A2 => n25262, Z => n6922);
   U19613 : XOR2_X1 port map( A1 => n15779, A2 => n13711, Z => n6924);
   U19619 : XOR2_X1 port map( A1 => n6930, A2 => n30006, Z => n29068);
   U19620 : XOR2_X1 port map( A1 => n6930, A2 => n29671, Z => n29028);
   U19622 : XOR2_X1 port map( A1 => n38703, A2 => n29538, Z => n20136);
   U19625 : NAND3_X2 port map( A1 => n10476, A2 => n10475, A3 => n25378, ZN => 
                           n7133);
   U19627 : XOR2_X1 port map( A1 => n19384, A2 => n26244, Z => n9490);
   U19631 : XOR2_X1 port map( A1 => n6942, A2 => n6941, Z => n6940);
   U19632 : XOR2_X1 port map( A1 => n23658, A2 => n29357, Z => n6941);
   U19633 : XOR2_X1 port map( A1 => n33322, A2 => n24002, Z => n6942);
   U19636 : OAI21_X1 port map( A1 => n24590, A2 => n5056, B => n6944, ZN => 
                           n16077);
   U19640 : NOR2_X2 port map( A1 => n8496, A2 => n9165, ZN => n21995);
   U19641 : NOR2_X1 port map( A1 => n36303, A2 => n39489, ZN => n6948);
   U19642 : INV_X1 port map( I => n17478, ZN => n10560);
   U19643 : XOR2_X1 port map( A1 => n23888, A2 => n18006, Z => n6951);
   U19644 : XOR2_X1 port map( A1 => n23988, A2 => n23609, Z => n6952);
   U19645 : XNOR2_X1 port map( A1 => n17478, A2 => n23762, ZN => n23745);
   U19648 : AOI21_X2 port map( A1 => n6956, A2 => n23828, B => n6955, ZN => 
                           n24696);
   U19649 : NAND2_X1 port map( A1 => n39196, A2 => n24805, ZN => n6957);
   U19666 : OAI22_X1 port map( A1 => n6981, A2 => n22157, B1 => n22225, B2 => 
                           n6982, ZN => n22087);
   U19667 : NAND2_X1 port map( A1 => n6982, A2 => n7357, ZN => n6981);
   U19669 : NAND2_X1 port map( A1 => n8275, A2 => n22364, ZN => n6982);
   U19670 : NAND2_X2 port map( A1 => n21625, A2 => n15468, ZN => n8275);
   U19674 : XOR2_X1 port map( A1 => n6987, A2 => n6986, Z => n6985);
   U19675 : XOR2_X1 port map( A1 => n23903, A2 => n29476, Z => n6986);
   U19677 : NAND3_X2 port map( A1 => n6994, A2 => n11842, A3 => n6992, ZN => 
                           n23755);
   U19680 : XOR2_X1 port map( A1 => n24982, A2 => n29223, Z => n6996);
   U19685 : NAND3_X1 port map( A1 => n1595, A2 => n1127, A3 => n15385, ZN => 
                           n7000);
   U19690 : OAI21_X2 port map( A1 => n7007, A2 => n7006, B => n7005, ZN => 
                           n9144);
   U19694 : NAND2_X2 port map( A1 => n21213, A2 => n7009, ZN => n23331);
   U19703 : AOI21_X1 port map( A1 => n24804, A2 => n24829, B => n15664, ZN => 
                           n10521);
   U19705 : INV_X2 port map( I => n14367, ZN => n23042);
   U19707 : NAND2_X2 port map( A1 => n28565, A2 => n28564, ZN => n28983);
   U19711 : XOR2_X1 port map( A1 => n19571, A2 => n29303, Z => n7032);
   U19716 : XOR2_X1 port map( A1 => n7039, A2 => n7038, Z => n7037);
   U19720 : XOR2_X1 port map( A1 => n37023, A2 => n22167, Z => n7040);
   U19726 : NAND2_X1 port map( A1 => n7046, A2 => n33713, ZN => n18951);
   U19727 : INV_X1 port map( I => n21795, ZN => n7047);
   U19731 : XOR2_X1 port map( A1 => n27672, A2 => n29229, Z => n7060);
   U19738 : NAND3_X1 port map( A1 => n10906, A2 => n28686, A3 => n36663, ZN => 
                           n28587);
   U19741 : OAI21_X1 port map( A1 => n24789, A2 => n31161, B => n20039, ZN => 
                           n7066);
   U19747 : XOR2_X1 port map( A1 => n19606, A2 => n29411, Z => n7069);
   U19748 : XOR2_X1 port map( A1 => n29824, A2 => n19722, Z => n7070);
   U19755 : XOR2_X1 port map( A1 => n10794, A2 => n1370, Z => n7089);
   U19770 : NAND2_X1 port map( A1 => n9875, A2 => n27197, ZN => n12031);
   U19775 : XOR2_X1 port map( A1 => n12838, A2 => n29849, Z => n7101);
   U19780 : AOI21_X1 port map( A1 => n20376, A2 => n19017, B => n1154, ZN => 
                           n7104);
   U19785 : XOR2_X1 port map( A1 => n23970, A2 => n39482, Z => n7113);
   U19790 : XOR2_X1 port map( A1 => n1658, A2 => n19127, Z => n7119);
   U19792 : INV_X2 port map( I => n18732, ZN => n28205);
   U19793 : XOR2_X1 port map( A1 => n7120, A2 => n7123, Z => n22864);
   U19796 : XOR2_X1 port map( A1 => n7510, A2 => n17153, Z => n7123);
   U19797 : INV_X2 port map( I => n7124, ZN => n7304);
   U19798 : XNOR2_X1 port map( A1 => Plaintext(20), A2 => Key(20), ZN => n7124)
                           ;
   U19799 : XOR2_X1 port map( A1 => n24925, A2 => n15912, Z => n18584);
   U19800 : XOR2_X1 port map( A1 => n15912, A2 => n30065, Z => n25035);
   U19803 : XOR2_X1 port map( A1 => n7127, A2 => n7126, Z => n7125);
   U19804 : XOR2_X1 port map( A1 => n24040, A2 => n1362, Z => n7126);
   U19809 : XOR2_X1 port map( A1 => n26244, A2 => n1096, Z => n10317);
   U19811 : NOR2_X1 port map( A1 => n15121, A2 => n7134, ZN => n15021);
   U19814 : NAND2_X2 port map( A1 => n22211, A2 => n22210, ZN => n22665);
   U19817 : NAND2_X1 port map( A1 => n7146, A2 => n23229, ZN => n7145);
   U19820 : XOR2_X1 port map( A1 => n25254, A2 => n25001, Z => n7152);
   U19821 : XOR2_X1 port map( A1 => n20333, A2 => n38148, Z => n25001);
   U19822 : XOR2_X1 port map( A1 => n25002, A2 => n10905, Z => n7153);
   U19824 : XOR2_X1 port map( A1 => n25118, A2 => n24982, Z => n25002);
   U19833 : XOR2_X1 port map( A1 => n57, A2 => n7162, Z => n7161);
   U19834 : AOI21_X2 port map( A1 => n34086, A2 => n7167, B => n7166, ZN => 
                           n17469);
   U19839 : XOR2_X1 port map( A1 => n15216, A2 => n18905, Z => n7180);
   U19844 : XOR2_X1 port map( A1 => n39631, A2 => n1413, Z => n7182);
   U19853 : NOR2_X1 port map( A1 => n13088, A2 => n7195, ZN => n13951);
   U19860 : XOR2_X1 port map( A1 => n1662, A2 => n17195, Z => n7200);
   U19862 : XOR2_X1 port map( A1 => n19071, A2 => n7202, Z => n9894);
   U19863 : XOR2_X1 port map( A1 => n19656, A2 => n29229, Z => n7202);
   U19864 : XOR2_X1 port map( A1 => n7203, A2 => n7206, Z => n17764);
   U19865 : XOR2_X1 port map( A1 => n25313, A2 => n7204, Z => n7203);
   U19866 : XOR2_X1 port map( A1 => n39295, A2 => n24926, Z => n7204);
   U19867 : XOR2_X1 port map( A1 => n35237, A2 => n20828, Z => n7206);
   U19869 : NAND2_X1 port map( A1 => n29952, A2 => n7208, ZN => n29953);
   U19873 : XOR2_X1 port map( A1 => n3082, A2 => n15617, Z => n8285);
   U19874 : XOR2_X1 port map( A1 => n35320, A2 => n3082, Z => n20137);
   U19875 : AND2_X1 port map( A1 => n19017, A2 => n1154, Z => n22149);
   U19878 : OAI21_X2 port map( A1 => n7232, A2 => n7230, B => n26998, ZN => 
                           n27503);
   U19879 : NAND2_X2 port map( A1 => n37393, A2 => n33263, ZN => n25940);
   U19882 : INV_X2 port map( I => n25719, ZN => n19237);
   U19883 : XNOR2_X1 port map( A1 => n27854, A2 => n38158, ZN => n27628);
   U19884 : XOR2_X1 port map( A1 => n10782, A2 => n7257, Z => n7256);
   U19886 : XOR2_X1 port map( A1 => n27674, A2 => n1467, Z => n7257);
   U19888 : NAND2_X1 port map( A1 => n37160, A2 => n32722, ZN => n14840);
   U19890 : NAND2_X1 port map( A1 => n1147, A2 => n7266, ZN => n23191);
   U19892 : NAND3_X1 port map( A1 => n7267, A2 => n24799, A3 => n17350, ZN => 
                           n16570);
   U19893 : AOI21_X1 port map( A1 => n7267, A2 => n19679, B => n33409, ZN => 
                           n8575);
   U19896 : NAND2_X2 port map( A1 => n17980, A2 => n17982, ZN => n29980);
   U19898 : XOR2_X1 port map( A1 => n16667, A2 => n17310, Z => n7275);
   U19899 : XOR2_X1 port map( A1 => n37023, A2 => n7277, Z => n7276);
   U19901 : INV_X2 port map( I => n12951, ZN => n19857);
   U19903 : NAND2_X1 port map( A1 => n21383, A2 => n21384, ZN => n19911);
   U19912 : NAND2_X1 port map( A1 => n23639, A2 => n35232, ZN => n23470);
   U19914 : AND2_X1 port map( A1 => n17648, A2 => n23617, Z => n12426);
   U19923 : NAND2_X1 port map( A1 => n27278, A2 => n7291, ZN => n7300);
   U19928 : INV_X1 port map( I => n10413, ZN => n7737);
   U19932 : XNOR2_X1 port map( A1 => n39063, A2 => n19851, ZN => n17921);
   U19937 : XOR2_X1 port map( A1 => n7316, A2 => n7667, Z => n28841);
   U19938 : XOR2_X1 port map( A1 => n29145, A2 => n14956, Z => n7316);
   U19947 : OAI21_X1 port map( A1 => n20538, A2 => n20342, B => n7318, ZN => 
                           n10409);
   U19950 : NAND2_X2 port map( A1 => n18641, A2 => n18640, ZN => n27830);
   U19952 : NOR2_X1 port map( A1 => n9276, A2 => n17087, ZN => n9849);
   U19955 : AND2_X1 port map( A1 => n18406, A2 => n9413, Z => n11835);
   U19957 : XOR2_X1 port map( A1 => n17455, A2 => n19919, Z => n17396);
   U19958 : XOR2_X1 port map( A1 => n23912, A2 => n29857, Z => n10312);
   U19966 : XOR2_X1 port map( A1 => n11318, A2 => n24988, Z => n7329);
   U19967 : NOR2_X2 port map( A1 => n13922, A2 => n20356, ZN => n9626);
   U19969 : NAND2_X1 port map( A1 => n34004, A2 => n35269, ZN => n9650);
   U19975 : XOR2_X1 port map( A1 => n18267, A2 => n26368, Z => n26832);
   U19976 : NAND2_X1 port map( A1 => n8000, A2 => n17934, ZN => n12844);
   U19983 : AND2_X1 port map( A1 => n24335, A2 => n545, Z => n14581);
   U19987 : XOR2_X1 port map( A1 => n22755, A2 => n704, Z => n7341);
   U19988 : OAI21_X2 port map( A1 => n27661, A2 => n27557, B => n10801, ZN => 
                           n27648);
   U19991 : NOR2_X2 port map( A1 => n26853, A2 => n7349, ZN => n27320);
   U19992 : NOR3_X1 port map( A1 => n26944, A2 => n19425, A3 => n15670, ZN => 
                           n7349);
   U19999 : XOR2_X1 port map( A1 => n27606, A2 => n18817, Z => n7353);
   U20000 : XOR2_X1 port map( A1 => n22712, A2 => n22617, Z => n13840);
   U20001 : INV_X1 port map( I => n14991, ZN => n14990);
   U20006 : XOR2_X1 port map( A1 => n24060, A2 => n7360, Z => n7359);
   U20019 : NAND3_X1 port map( A1 => n8568, A2 => n15173, A3 => n36708, ZN => 
                           n7362);
   U20022 : INV_X2 port map( I => n25782, ZN => n26108);
   U20030 : XOR2_X1 port map( A1 => n334, A2 => n30169, Z => n7698);
   U20037 : OR2_X1 port map( A1 => n29794, A2 => n18257, Z => n29787);
   U20045 : XOR2_X1 port map( A1 => n25000, A2 => n810, Z => n7380);
   U20047 : XOR2_X1 port map( A1 => n28985, A2 => n765, Z => n7382);
   U20052 : MUX2_X1 port map( I0 => n27363, I1 => n34001, S => n21101, Z => 
                           n27056);
   U20056 : INV_X1 port map( I => n13004, ZN => n7393);
   U20058 : NOR2_X1 port map( A1 => n18377, A2 => n22991, ZN => n8011);
   U20060 : OAI21_X1 port map( A1 => n9460, A2 => n9459, B => n10220, ZN => 
                           n10219);
   U20072 : OR2_X1 port map( A1 => n10634, A2 => n18072, Z => n21120);
   U20074 : XNOR2_X1 port map( A1 => n26246, A2 => n35212, ZN => n26166);
   U20079 : AND2_X1 port map( A1 => n20734, A2 => n31452, Z => n8927);
   U20082 : INV_X1 port map( I => n20243, ZN => n15058);
   U20100 : XOR2_X1 port map( A1 => n27825, A2 => n27540, Z => n27667);
   U20104 : XOR2_X1 port map( A1 => n8199, A2 => n11475, Z => n10970);
   U20106 : XOR2_X1 port map( A1 => n8401, A2 => n27577, Z => n8403);
   U20109 : AOI21_X1 port map( A1 => n7303, A2 => n38200, B => n969, ZN => 
                           n29466);
   U20113 : AND2_X1 port map( A1 => n29662, A2 => n19297, Z => n29654);
   U20115 : XOR2_X1 port map( A1 => n23680, A2 => n7917, Z => n10279);
   U20118 : NOR2_X1 port map( A1 => n26133, A2 => n13678, ZN => n13677);
   U20119 : NAND2_X1 port map( A1 => n20807, A2 => n20696, ZN => n11963);
   U20122 : XOR2_X1 port map( A1 => n22435, A2 => n12598, Z => n7498);
   U20123 : NOR2_X2 port map( A1 => n7443, A2 => n9148, ZN => n17184);
   U20124 : XOR2_X1 port map( A1 => n1667, A2 => n22766, Z => n22606);
   U20125 : OAI21_X2 port map( A1 => n17409, A2 => n17408, B => n17407, ZN => 
                           n22766);
   U20127 : XOR2_X1 port map( A1 => n29070, A2 => n1409, Z => n20675);
   U20128 : INV_X1 port map( I => n25897, ZN => n16444);
   U20129 : OR2_X1 port map( A1 => n29218, A2 => n29219, Z => n13104);
   U20138 : XOR2_X1 port map( A1 => n7451, A2 => n15432, Z => Ciphertext(72));
   U20139 : AOI22_X1 port map( A1 => n20126, A2 => n29618, B1 => n29601, B2 => 
                           n29616, ZN => n7451);
   U20146 : OR3_X1 port map( A1 => n34906, A2 => n24733, A3 => n24839, Z => 
                           n11367);
   U20149 : AND2_X1 port map( A1 => n22900, A2 => n2350, Z => n14483);
   U20152 : XOR2_X1 port map( A1 => n26497, A2 => n26496, Z => n26502);
   U20154 : INV_X2 port map( I => n7459, ZN => n8818);
   U20157 : INV_X2 port map( I => n7462, ZN => n14459);
   U20163 : OAI21_X1 port map( A1 => n17262, A2 => n29567, B => n1053, ZN => 
                           n13926);
   U20165 : OR2_X1 port map( A1 => n27233, A2 => n12306, Z => n7472);
   U20172 : NAND2_X1 port map( A1 => n17939, A2 => n16534, ZN => n16533);
   U20173 : AOI21_X1 port map( A1 => n14582, A2 => n30323, B => n16533, ZN => 
                           n16532);
   U20174 : INV_X1 port map( I => n16179, ZN => n24294);
   U20175 : NAND2_X1 port map( A1 => n25937, A2 => n1105, ZN => n14133);
   U20176 : XOR2_X1 port map( A1 => n13035, A2 => n18800, Z => n8564);
   U20177 : XOR2_X1 port map( A1 => n26396, A2 => n12649, Z => n19051);
   U20178 : NAND3_X2 port map( A1 => n25478, A2 => n11063, A3 => n25460, ZN => 
                           n11064);
   U20180 : AOI22_X1 port map( A1 => n17318, A2 => n1389, B1 => n17317, B2 => 
                           n29437, ZN => n7572);
   U20184 : XOR2_X1 port map( A1 => n27728, A2 => n17721, Z => n8975);
   U20190 : INV_X2 port map( I => n7492, ZN => n25540);
   U20191 : INV_X1 port map( I => n1283, ZN => n13185);
   U20193 : AND2_X1 port map( A1 => n36162, A2 => n3985, Z => n25373);
   U20199 : AOI21_X1 port map( A1 => n7502, A2 => n29633, B => n29700, ZN => 
                           n29198);
   U20206 : AND3_X1 port map( A1 => n13770, A2 => n26811, A3 => n26810, Z => 
                           n7628);
   U20208 : XNOR2_X1 port map( A1 => n31823, A2 => n18273, ZN => n10546);
   U20210 : XOR2_X1 port map( A1 => n32298, A2 => n27830, Z => n27657);
   U20213 : XOR2_X1 port map( A1 => n7507, A2 => n29964, Z => Ciphertext(132));
   U20214 : OAI22_X1 port map( A1 => n29963, A2 => n29977, B1 => n29962, B2 => 
                           n1170, ZN => n7507);
   U20224 : NOR2_X2 port map( A1 => n31569, A2 => n29927, ZN => n29923);
   U20234 : NAND2_X1 port map( A1 => n32865, A2 => n11700, ZN => n19164);
   U20237 : AND2_X1 port map( A1 => n30158, A2 => n20541, Z => n14539);
   U20238 : OAI22_X2 port map( A1 => n21553, A2 => n21908, B1 => n7526, B2 => 
                           n21645, ZN => n19604);
   U20246 : OR2_X1 port map( A1 => n22324, A2 => n22322, Z => n11345);
   U20252 : NOR2_X1 port map( A1 => n12168, A2 => n11330, ZN => n7539);
   U20254 : XOR2_X1 port map( A1 => n10668, A2 => n16591, Z => n7543);
   U20256 : XOR2_X1 port map( A1 => n29159, A2 => n7546, Z => n28805);
   U20257 : XOR2_X1 port map( A1 => n973, A2 => n29828, Z => n7546);
   U20258 : XOR2_X1 port map( A1 => n10156, A2 => n7547, Z => n10155);
   U20259 : XOR2_X1 port map( A1 => n28914, A2 => n7548, Z => n7547);
   U20260 : NAND2_X2 port map( A1 => n9382, A2 => n9381, ZN => n9385);
   U20261 : NAND3_X1 port map( A1 => n26635, A2 => n26634, A3 => n4748, ZN => 
                           n26638);
   U20263 : INV_X4 port map( I => n10632, ZN => n22342);
   U20270 : OR2_X1 port map( A1 => n26976, A2 => n36262, Z => n10853);
   U20271 : NAND2_X1 port map( A1 => n9737, A2 => n13997, ZN => n11124);
   U20272 : XOR2_X1 port map( A1 => n26537, A2 => n26538, Z => n8020);
   U20280 : NAND2_X1 port map( A1 => n12526, A2 => n12525, ZN => n12524);
   U20287 : XOR2_X1 port map( A1 => n25072, A2 => n7569, Z => n7762);
   U20288 : XOR2_X1 port map( A1 => n25179, A2 => n35707, Z => n7569);
   U20289 : XOR2_X1 port map( A1 => n7570, A2 => n846, Z => n7959);
   U20290 : XOR2_X1 port map( A1 => n11374, A2 => n7571, Z => n7570);
   U20291 : XOR2_X1 port map( A1 => n7572, A2 => n17316, Z => Ciphertext(44));
   U20293 : XOR2_X1 port map( A1 => n26276, A2 => n11902, Z => n7573);
   U20302 : OAI21_X1 port map( A1 => n19570, A2 => n19569, B => n27286, ZN => 
                           n11487);
   U20309 : XNOR2_X1 port map( A1 => n29026, A2 => n14689, ZN => n11405);
   U20310 : NAND3_X1 port map( A1 => n5921, A2 => n29721, A3 => n20498, ZN => 
                           n29713);
   U20314 : XOR2_X1 port map( A1 => n7589, A2 => n19953, Z => Ciphertext(94));
   U20327 : XNOR2_X1 port map( A1 => n27825, A2 => n35229, ZN => n11031);
   U20329 : XOR2_X1 port map( A1 => n20811, A2 => n28829, Z => n16380);
   U20330 : XOR2_X1 port map( A1 => n28991, A2 => n29247, Z => n28829);
   U20344 : AND2_X1 port map( A1 => n23550, A2 => n35191, Z => n18617);
   U20350 : INV_X1 port map( I => n28523, ZN => n12609);
   U20352 : XOR2_X1 port map( A1 => n13247, A2 => n23995, Z => n13246);
   U20354 : XOR2_X1 port map( A1 => n23889, A2 => n32230, Z => n23724);
   U20356 : XOR2_X1 port map( A1 => n20101, A2 => n839, Z => n14440);
   U20358 : OR2_X1 port map( A1 => n13415, A2 => n34666, Z => n18264);
   U20363 : XOR2_X1 port map( A1 => n9120, A2 => n738, Z => n7623);
   U20373 : AOI21_X1 port map( A1 => n16722, A2 => n30109, B => n1052, ZN => 
                           n16721);
   U20377 : XOR2_X1 port map( A1 => n19112, A2 => n23672, Z => n7981);
   U20379 : XOR2_X1 port map( A1 => n25161, A2 => n17457, Z => n11161);
   U20385 : OAI22_X1 port map( A1 => n11939, A2 => n15509, B1 => n8955, B2 => 
                           n15535, ZN => n7637);
   U20389 : XOR2_X1 port map( A1 => n18133, A2 => n28982, Z => n28913);
   U20392 : OR2_X1 port map( A1 => n1630, A2 => n23325, Z => n19666);
   U20399 : XOR2_X1 port map( A1 => n8563, A2 => n8564, Z => n16327);
   U20401 : NAND3_X1 port map( A1 => n1172, A2 => n13786, A3 => n38204, ZN => 
                           n18231);
   U20407 : XOR2_X1 port map( A1 => n7661, A2 => n26455, Z => n26309);
   U20412 : XOR2_X1 port map( A1 => n7663, A2 => n9270, Z => n18923);
   U20413 : XOR2_X1 port map( A1 => n18924, A2 => n27672, Z => n7663);
   U20417 : XOR2_X1 port map( A1 => n28710, A2 => n7665, Z => n7664);
   U20418 : INV_X2 port map( I => n7666, ZN => n10422);
   U20422 : NOR3_X1 port map( A1 => n3989, A2 => n19467, A3 => n28255, ZN => 
                           n9880);
   U20433 : NAND2_X1 port map( A1 => n25769, A2 => n25943, ZN => n7678);
   U20434 : XOR2_X1 port map( A1 => n7681, A2 => n1362, Z => Ciphertext(191));
   U20438 : XNOR2_X1 port map( A1 => n13243, A2 => n13242, ZN => n7720);
   U20444 : XOR2_X1 port map( A1 => n27539, A2 => n12495, Z => n12494);
   U20453 : XOR2_X1 port map( A1 => n9980, A2 => n12283, Z => n22862);
   U20459 : XOR2_X1 port map( A1 => n7698, A2 => n8585, Z => n8586);
   U20473 : XOR2_X1 port map( A1 => n25204, A2 => n1735, Z => n24962);
   U20474 : AOI21_X2 port map( A1 => n13893, A2 => n13894, B => n8733, ZN => 
                           n7710);
   U20484 : AND3_X1 port map( A1 => n27048, A2 => n27047, A3 => n27046, Z => 
                           n7716);
   U20493 : XNOR2_X1 port map( A1 => n29253, A2 => n19730, ZN => n10087);
   U20494 : NAND2_X1 port map( A1 => n14132, A2 => n25813, ZN => n7724);
   U20496 : OR3_X1 port map( A1 => n1276, A2 => n1127, A3 => n24232, Z => 
                           n18759);
   U20497 : NOR2_X1 port map( A1 => n16924, A2 => n9178, ZN => n20462);
   U20498 : OR2_X1 port map( A1 => n11805, A2 => n35919, Z => n26913);
   U20507 : NAND3_X2 port map( A1 => n16312, A2 => n24268, A3 => n16311, ZN => 
                           n24912);
   U20509 : XOR2_X1 port map( A1 => n31627, A2 => n26287, Z => n10967);
   U20512 : XOR2_X1 port map( A1 => n31339, A2 => n35596, Z => n22321);
   U20524 : XNOR2_X1 port map( A1 => n38152, A2 => n19592, ZN => n7801);
   U20538 : XOR2_X1 port map( A1 => n14219, A2 => n16055, Z => n23715);
   U20549 : XOR2_X1 port map( A1 => n35505, A2 => n7287, Z => n9093);
   U20554 : XOR2_X1 port map( A1 => n7763, A2 => n18371, Z => n8002);
   U20557 : XOR2_X1 port map( A1 => n27813, A2 => n673, Z => n7764);
   U20561 : OR2_X2 port map( A1 => n29198, A2 => n7765, Z => n29732);
   U20562 : OAI21_X1 port map( A1 => n29197, A2 => n29702, B => n34180, ZN => 
                           n7765);
   U20563 : XOR2_X1 port map( A1 => n12265, A2 => n12266, Z => n12759);
   U20565 : OAI21_X1 port map( A1 => n29611, A2 => n29618, B => n9045, ZN => 
                           n9044);
   U20568 : XOR2_X1 port map( A1 => n7779, A2 => n7780, Z => n26768);
   U20569 : XOR2_X1 port map( A1 => n26442, A2 => n15750, Z => n7779);
   U20573 : XOR2_X1 port map( A1 => n18849, A2 => n1368, Z => n7783);
   U20576 : XOR2_X1 port map( A1 => n26324, A2 => n1237, Z => n7785);
   U20577 : XOR2_X1 port map( A1 => n20425, A2 => n7787, Z => n7786);
   U20578 : XNOR2_X1 port map( A1 => n26223, A2 => n26598, ZN => n20425);
   U20579 : NOR2_X1 port map( A1 => n5077, A2 => n22215, ZN => n11202);
   U20580 : NAND2_X1 port map( A1 => n9938, A2 => n5077, ZN => n22009);
   U20581 : NAND2_X1 port map( A1 => n15488, A2 => n5077, ZN => n15487);
   U20586 : AOI21_X1 port map( A1 => n30214, A2 => n14387, B => n30217, ZN => 
                           n7795);
   U20587 : NAND2_X1 port map( A1 => n7892, A2 => n30210, ZN => n7796);
   U20600 : XOR2_X1 port map( A1 => n23700, A2 => n7832, Z => n13369);
   U20601 : XOR2_X1 port map( A1 => n7833, A2 => n23973, Z => n7832);
   U20606 : NOR2_X2 port map( A1 => n15072, A2 => n14526, ZN => n7843);
   U20608 : XOR2_X1 port map( A1 => n23980, A2 => n21046, Z => n21045);
   U20609 : XOR2_X1 port map( A1 => n7848, A2 => n29021, Z => n28333);
   U20610 : NAND3_X1 port map( A1 => n1438, A2 => n39235, A3 => n9514, ZN => 
                           n14790);
   U20622 : NAND2_X2 port map( A1 => n7868, A2 => n7867, ZN => n20352);
   U20623 : XOR2_X1 port map( A1 => n7870, A2 => n10794, Z => n19308);
   U20624 : XOR2_X1 port map( A1 => n9108, A2 => n19929, Z => n7870);
   U20625 : INV_X2 port map( I => n12686, ZN => n19420);
   U20629 : OR2_X1 port map( A1 => n19731, A2 => n21132, Z => n22947);
   U20630 : XOR2_X1 port map( A1 => n21133, A2 => n22415, Z => n19731);
   U20635 : XOR2_X1 port map( A1 => n8473, A2 => n8939, Z => n12357);
   U20644 : INV_X1 port map( I => n7914, ZN => n14713);
   U20646 : NAND2_X1 port map( A1 => n7914, A2 => n28625, ZN => n21004);
   U20648 : XOR2_X1 port map( A1 => n11938, A2 => n23696, Z => n7920);
   U20651 : XOR2_X1 port map( A1 => n1618, A2 => n1357, Z => n7919);
   U20656 : XOR2_X1 port map( A1 => n8729, A2 => n35262, Z => n28987);
   U20658 : XOR2_X1 port map( A1 => n29820, A2 => n1050, Z => n7929);
   U20659 : XOR2_X1 port map( A1 => n7931, A2 => n7932, Z => n13635);
   U20662 : XOR2_X1 port map( A1 => n18595, A2 => n22411, Z => n22447);
   U20664 : NAND3_X1 port map( A1 => n34179, A2 => n9918, A3 => n31629, ZN => 
                           n7933);
   U20665 : NOR2_X2 port map( A1 => n7591, A2 => n20053, ZN => n8498);
   U20672 : AOI22_X2 port map( A1 => n20037, A2 => n21645, B1 => n21462, B2 => 
                           n21910, ZN => n21553);
   U20673 : NOR2_X2 port map( A1 => n20037, A2 => n39650, ZN => n21719);
   U20677 : XOR2_X1 port map( A1 => n7980, A2 => n7979, Z => n26704);
   U20680 : NAND2_X2 port map( A1 => n7969, A2 => n7968, ZN => n25278);
   U20683 : XOR2_X1 port map( A1 => n25853, A2 => n747, Z => n7979);
   U20690 : OAI22_X2 port map( A1 => n21439, A2 => n21853, B1 => n21438, B2 => 
                           n21687, ZN => n8040);
   U20693 : OAI22_X2 port map( A1 => n33978, A2 => n9312, B1 => n9320, B2 => 
                           n18801, ZN => n26180);
   U20696 : NAND3_X1 port map( A1 => n36183, A2 => n1225, A3 => n27337, ZN => 
                           n18268);
   U20706 : NOR2_X2 port map( A1 => n8012, A2 => n8011, ZN => n23607);
   U20710 : XOR2_X1 port map( A1 => n16270, A2 => n14053, Z => n8015);
   U20715 : NAND4_X1 port map( A1 => n8213, A2 => n8211, A3 => n18381, A4 => 
                           n18382, ZN => n8023);
   U20718 : NOR2_X2 port map( A1 => n21855, A2 => n21856, ZN => n22243);
   U20720 : NAND2_X1 port map( A1 => n6443, A2 => n30153, ZN => n8030);
   U20722 : XOR2_X1 port map( A1 => n22629, A2 => n29602, Z => n8037);
   U20723 : XOR2_X1 port map( A1 => n12267, A2 => n39548, Z => n8038);
   U20725 : NOR2_X1 port map( A1 => n30022, A2 => n8039, ZN => n30009);
   U20731 : INV_X1 port map( I => n11956, ZN => n28548);
   U20732 : INV_X1 port map( I => n28735, ZN => n16206);
   U20739 : XOR2_X1 port map( A1 => n19910, A2 => n8059, Z => n19183);
   U20741 : XOR2_X1 port map( A1 => n8060, A2 => n1169, Z => Ciphertext(98));
   U20743 : XOR2_X1 port map( A1 => n8067, A2 => n8066, Z => n8065);
   U20744 : XOR2_X1 port map( A1 => n36750, A2 => n29051, Z => n8066);
   U20745 : XOR2_X1 port map( A1 => n22620, A2 => n12243, Z => n8067);
   U20747 : OAI21_X2 port map( A1 => n17358, A2 => n20798, B => n17356, ZN => 
                           n22371);
   U20749 : XOR2_X1 port map( A1 => n8075, A2 => n26600, Z => n8074);
   U20751 : NOR2_X1 port map( A1 => n14837, A2 => n33899, ZN => n8076);
   U20753 : NOR2_X1 port map( A1 => n20632, A2 => n8078, ZN => n10806);
   U20756 : XNOR2_X1 port map( A1 => n17276, A2 => n17273, ZN => n8078);
   U20758 : NOR2_X1 port map( A1 => n28486, A2 => n8082, ZN => n28031);
   U20759 : NAND2_X1 port map( A1 => n1066, A2 => n8082, ZN => n28392);
   U20760 : NOR2_X1 port map( A1 => n28483, A2 => n8082, ZN => n19610);
   U20761 : NOR2_X1 port map( A1 => n16559, A2 => n8082, ZN => n8658);
   U20762 : NAND2_X1 port map( A1 => n12343, A2 => n8082, ZN => n12342);
   U20763 : NAND2_X1 port map( A1 => n36573, A2 => n18144, ZN => n8085);
   U20768 : XOR2_X1 port map( A1 => n27712, A2 => n16759, Z => n8100);
   U20771 : AND2_X1 port map( A1 => n24681, A2 => n8109, Z => n8108);
   U20775 : NOR2_X1 port map( A1 => n124, A2 => n20313, ZN => n11757);
   U20777 : XOR2_X1 port map( A1 => n6522, A2 => n21003, Z => n8119);
   U20778 : NOR2_X1 port map( A1 => n24895, A2 => n25583, ZN => n8123);
   U20782 : OAI21_X2 port map( A1 => n8127, A2 => n24877, B => n8125, ZN => 
                           n21028);
   U20783 : INV_X2 port map( I => n8128, ZN => n16080);
   U20789 : XOR2_X1 port map( A1 => n26476, A2 => n8585, Z => n8132);
   U20790 : XOR2_X1 port map( A1 => n38951, A2 => n19717, Z => n8136);
   U20795 : NAND2_X2 port map( A1 => n13748, A2 => n13747, ZN => n8139);
   U20798 : INV_X2 port map( I => n8151, ZN => n22915);
   U20804 : XOR2_X1 port map( A1 => n8163, A2 => n19624, Z => n25260);
   U20805 : XOR2_X1 port map( A1 => n8163, A2 => n29238, Z => n24952);
   U20811 : XOR2_X1 port map( A1 => n8171, A2 => n17060, Z => n23152);
   U20812 : XOR2_X1 port map( A1 => n8172, A2 => n13295, Z => n8171);
   U20813 : XOR2_X1 port map( A1 => n8176, A2 => n8180, Z => n26746);
   U20815 : XOR2_X1 port map( A1 => n12839, A2 => n35984, Z => n8177);
   U20817 : XOR2_X1 port map( A1 => n8502, A2 => n9018, Z => n8180);
   U20823 : INV_X2 port map( I => n8186, ZN => n14383);
   U20824 : XNOR2_X1 port map( A1 => n8187, A2 => n8188, ZN => n8186);
   U20826 : XOR2_X1 port map( A1 => n8189, A2 => n26429, Z => n8188);
   U20829 : NAND2_X1 port map( A1 => n8201, A2 => n8193, ZN => n8200);
   U20831 : OAI21_X2 port map( A1 => n8338, A2 => n8892, B => n8202, ZN => 
                           n13786);
   U20833 : NAND2_X2 port map( A1 => n9251, A2 => n21127, ZN => n8882);
   U20834 : INV_X2 port map( I => n8205, ZN => n14478);
   U20835 : NOR2_X2 port map( A1 => n8205, A2 => n16081, ZN => n10815);
   U20836 : NAND2_X1 port map( A1 => n7424, A2 => n14949, ZN => n27035);
   U20839 : NOR2_X2 port map( A1 => n27036, A2 => n19034, ZN => n27570);
   U20840 : XOR2_X1 port map( A1 => n31214, A2 => n19877, Z => n18969);
   U20848 : XOR2_X1 port map( A1 => n32448, A2 => n21280, Z => n14476);
   U20849 : XOR2_X1 port map( A1 => n32448, A2 => n33320, Z => n28857);
   U20851 : MUX2_X1 port map( I0 => n8236, I1 => n26077, S => n11807, Z => 
                           n8235);
   U20854 : XOR2_X1 port map( A1 => n8244, A2 => n8242, Z => n11497);
   U20855 : XOR2_X1 port map( A1 => n25081, A2 => n8243, Z => n8242);
   U20856 : XOR2_X1 port map( A1 => n16627, A2 => n1358, Z => n8243);
   U20857 : XOR2_X1 port map( A1 => n25032, A2 => n25314, Z => n8244);
   U20859 : XOR2_X1 port map( A1 => n8247, A2 => n8246, Z => n12634);
   U20860 : XOR2_X1 port map( A1 => n26560, A2 => n30473, Z => n8246);
   U20861 : XOR2_X1 port map( A1 => n26594, A2 => n26305, Z => n26560);
   U20864 : NAND2_X1 port map( A1 => n27560, A2 => n8253, ZN => n27561);
   U20867 : NOR2_X1 port map( A1 => n27456, A2 => n27455, ZN => n8257);
   U20869 : NAND2_X2 port map( A1 => n26638, A2 => n26637, ZN => n27240);
   U20878 : XOR2_X1 port map( A1 => n25080, A2 => n1260, Z => n8276);
   U20883 : XOR2_X1 port map( A1 => n27464, A2 => n27503, Z => n27650);
   U20884 : XOR2_X1 port map( A1 => n27848, A2 => n35189, Z => n8280);
   U20888 : XOR2_X1 port map( A1 => n38190, A2 => n30324, Z => n8283);
   U20892 : NAND2_X1 port map( A1 => n8287, A2 => n20274, ZN => n20510);
   U20895 : INV_X2 port map( I => n12001, ZN => n9751);
   U20901 : XOR2_X1 port map( A1 => n8299, A2 => n15160, Z => n8298);
   U20903 : XOR2_X1 port map( A1 => n25303, A2 => n25252, Z => n17804);
   U20906 : XOR2_X1 port map( A1 => n8303, A2 => n29978, Z => n12003);
   U20907 : XOR2_X1 port map( A1 => n16096, A2 => n8303, Z => n17643);
   U20908 : XOR2_X1 port map( A1 => n8303, A2 => n30016, Z => n28607);
   U20909 : NOR2_X1 port map( A1 => n8304, A2 => n16080, ZN => n14515);
   U20910 : OAI21_X1 port map( A1 => n34150, A2 => n8305, B => n15180, ZN => 
                           n25712);
   U20922 : XOR2_X1 port map( A1 => n8335, A2 => n8334, Z => n8333);
   U20923 : XOR2_X1 port map( A1 => n27778, A2 => n1704, Z => n8334);
   U20928 : XOR2_X1 port map( A1 => n26495, A2 => n29229, Z => n8340);
   U20935 : NOR2_X1 port map( A1 => n10940, A2 => n15873, ZN => n24410);
   U20937 : NAND2_X1 port map( A1 => n21929, A2 => n917, ZN => n21060);
   U20938 : NAND2_X2 port map( A1 => n20525, A2 => n20522, ZN => n30245);
   U20950 : AOI21_X1 port map( A1 => n5675, A2 => n32191, B => n33662, ZN => 
                           n8384);
   U20952 : AOI21_X1 port map( A1 => n23049, A2 => n8491, B => n8386, ZN => 
                           n23051);
   U20957 : XOR2_X1 port map( A1 => n18633, A2 => n8397, Z => n8396);
   U20964 : XOR2_X1 port map( A1 => n26448, A2 => n7602, Z => n8409);
   U20965 : XOR2_X1 port map( A1 => n26449, A2 => n9152, Z => n8410);
   U20967 : NAND2_X1 port map( A1 => n8412, A2 => n27211, ZN => n27096);
   U20970 : OAI21_X1 port map( A1 => n27438, A2 => n4771, B => n8412, ZN => 
                           n12916);
   U20975 : XOR2_X1 port map( A1 => n31293, A2 => n26519, Z => n26176);
   U20978 : XOR2_X1 port map( A1 => n8425, A2 => n27494, Z => n8424);
   U20985 : NAND2_X1 port map( A1 => n18148, A2 => n8430, ZN => n11609);
   U20987 : NAND3_X1 port map( A1 => n32817, A2 => n20679, A3 => n3676, ZN => 
                           n14904);
   U20988 : AOI21_X1 port map( A1 => n1341, A2 => n32817, B => n3676, ZN => 
                           n9223);
   U20990 : NAND2_X1 port map( A1 => n8799, A2 => n31381, ZN => n8438);
   U20994 : NAND3_X1 port map( A1 => n7278, A2 => n17242, A3 => n21898, ZN => 
                           n8441);
   U20995 : INV_X2 port map( I => n8443, ZN => n30057);
   U21002 : NAND2_X1 port map( A1 => n8463, A2 => n24294, ZN => n24208);
   U21004 : AOI21_X2 port map( A1 => n20680, A2 => n20682, B => n15490, ZN => 
                           n20679);
   U21008 : OAI21_X1 port map( A1 => n293, A2 => n8468, B => n19323, ZN => 
                           n21734);
   U21009 : NOR2_X1 port map( A1 => n18926, A2 => n8468, ZN => n8466);
   U21012 : XOR2_X1 port map( A1 => n8474, A2 => n8470, Z => n8469);
   U21013 : XOR2_X1 port map( A1 => n29147, A2 => n19498, Z => n8470);
   U21014 : XOR2_X1 port map( A1 => n8472, A2 => n29148, Z => n8471);
   U21015 : NAND2_X2 port map( A1 => n27914, A2 => n27913, ZN => n8476);
   U21019 : NOR2_X2 port map( A1 => n1245, A2 => n834, ZN => n18884);
   U21021 : XOR2_X1 port map( A1 => n25295, A2 => n8483, Z => n8482);
   U21022 : XOR2_X1 port map( A1 => n19359, A2 => n29509, Z => n8483);
   U21023 : XOR2_X1 port map( A1 => n2145, A2 => n23805, Z => n8632);
   U21026 : XOR2_X1 port map( A1 => n22574, A2 => n22576, Z => n13550);
   U21031 : NAND2_X1 port map( A1 => n19604, A2 => n396, ZN => n16936);
   U21032 : NOR2_X1 port map( A1 => n22313, A2 => n396, ZN => n15294);
   U21033 : NAND2_X1 port map( A1 => n13912, A2 => n396, ZN => n13911);
   U21036 : NOR2_X1 port map( A1 => n21929, A2 => n8495, ZN => n21059);
   U21037 : OAI22_X2 port map( A1 => n14813, A2 => n21928, B1 => n14811, B2 => 
                           n8495, ZN => n22337);
   U21038 : INV_X1 port map( I => n21927, ZN => n8495);
   U21044 : XOR2_X1 port map( A1 => n8671, A2 => n13215, Z => n8505);
   U21050 : XOR2_X1 port map( A1 => n8512, A2 => n8511, Z => n13904);
   U21051 : XOR2_X1 port map( A1 => n23918, A2 => n12553, Z => n8511);
   U21054 : XOR2_X1 port map( A1 => n13483, A2 => n8515, Z => n8514);
   U21055 : XOR2_X1 port map( A1 => n18785, A2 => n19835, Z => n8515);
   U21058 : XNOR2_X1 port map( A1 => Plaintext(12), A2 => Key(12), ZN => n8517)
                           ;
   U21062 : XOR2_X1 port map( A1 => n12690, A2 => n8528, Z => n11870);
   U21063 : XOR2_X1 port map( A1 => n19355, A2 => n1702, Z => n8528);
   U21066 : XOR2_X1 port map( A1 => n29823, A2 => n8531, Z => n8530);
   U21067 : XOR2_X1 port map( A1 => n31524, A2 => n30964, Z => n29823);
   U21070 : XOR2_X1 port map( A1 => n29824, A2 => n8532, Z => n8531);
   U21071 : XOR2_X1 port map( A1 => n29822, A2 => n29827, Z => n8533);
   U21072 : XOR2_X1 port map( A1 => n8852, A2 => n28943, Z => n29822);
   U21073 : NAND2_X1 port map( A1 => n8517, A2 => n21898, ZN => n20898);
   U21074 : INV_X2 port map( I => n14217, ZN => n14426);
   U21075 : XOR2_X1 port map( A1 => n27619, A2 => n27618, Z => n8540);
   U21077 : XOR2_X1 port map( A1 => n30761, A2 => n32218, Z => n16843);
   U21078 : XOR2_X1 port map( A1 => n25149, A2 => n30761, Z => n24953);
   U21080 : XOR2_X1 port map( A1 => n30761, A2 => n25014, Z => n24631);
   U21081 : NOR2_X1 port map( A1 => n29951, A2 => n29997, ZN => n19197);
   U21087 : XOR2_X1 port map( A1 => n10579, A2 => n27467, Z => n8553);
   U21091 : XOR2_X1 port map( A1 => n1503, A2 => n16735, Z => n8559);
   U21092 : INV_X1 port map( I => Plaintext(116), ZN => n8562);
   U21093 : XOR2_X1 port map( A1 => n8562, A2 => Key(116), Z => n9308);
   U21095 : XOR2_X1 port map( A1 => n8566, A2 => n18482, Z => n8565);
   U21096 : XOR2_X1 port map( A1 => n10526, A2 => n23931, Z => n18482);
   U21097 : XOR2_X1 port map( A1 => n24043, A2 => n23763, Z => n8567);
   U21098 : OR2_X1 port map( A1 => n21969, A2 => n34015, Z => n8570);
   U21104 : AOI21_X1 port map( A1 => n16187, A2 => n8584, B => n8582, ZN => 
                           n19138);
   U21105 : AOI21_X1 port map( A1 => n31570, A2 => n9591, B => n1174, ZN => 
                           n8584);
   U21110 : NAND3_X1 port map( A1 => n8731, A2 => n33256, A3 => n16224, ZN => 
                           n8590);
   U21111 : NAND2_X1 port map( A1 => n30049, A2 => n29936, ZN => n8593);
   U21120 : XOR2_X1 port map( A1 => n26432, A2 => n26517, Z => n8625);
   U21122 : XOR2_X1 port map( A1 => n26431, A2 => n14148, Z => n8626);
   U21127 : XOR2_X1 port map( A1 => n8632, A2 => n23806, Z => n8631);
   U21128 : INV_X2 port map( I => n8824, ZN => n13453);
   U21132 : XNOR2_X1 port map( A1 => Plaintext(15), A2 => Key(15), ZN => n8653)
                           ;
   U21136 : NAND2_X1 port map( A1 => n29901, A2 => n13607, ZN => n8666);
   U21146 : OR2_X1 port map( A1 => n23078, A2 => n20873, Z => n8674);
   U21149 : OAI21_X2 port map( A1 => n21143, A2 => n23076, B => n23078, ZN => 
                           n14804);
   U21150 : XOR2_X1 port map( A1 => n8678, A2 => n15808, Z => n14403);
   U21154 : NAND2_X1 port map( A1 => n22243, A2 => n37089, ZN => n8754);
   U21155 : NOR2_X1 port map( A1 => n37089, A2 => n21864, ZN => n8688);
   U21162 : XOR2_X1 port map( A1 => Plaintext(164), A2 => Key(164), Z => n21938
                           );
   U21163 : NOR3_X1 port map( A1 => n22349, A2 => n14423, A3 => n7955, ZN => 
                           n8701);
   U21165 : INV_X2 port map( I => n10733, ZN => n13584);
   U21174 : NAND3_X1 port map( A1 => n1477, A2 => n27412, A3 => n34969, ZN => 
                           n27159);
   U21180 : XOR2_X1 port map( A1 => n13374, A2 => n38962, Z => n8723);
   U21186 : NAND2_X1 port map( A1 => n14933, A2 => n8728, ZN => n14199);
   U21187 : AOI21_X1 port map( A1 => n16837, A2 => n16839, B => n8728, ZN => 
                           n16838);
   U21191 : XOR2_X1 port map( A1 => n29829, A2 => n29832, Z => n8732);
   U21192 : INV_X2 port map( I => n8736, ZN => n21436);
   U21193 : XNOR2_X1 port map( A1 => Plaintext(33), A2 => Key(33), ZN => n8736)
                           ;
   U21195 : NAND2_X1 port map( A1 => n955, A2 => n8738, ZN => n8737);
   U21205 : XOR2_X1 port map( A1 => n27502, A2 => n8748, Z => n8747);
   U21206 : XOR2_X1 port map( A1 => n29292, A2 => n29291, Z => n8755);
   U21211 : XOR2_X1 port map( A1 => n38154, A2 => n1938, Z => n11153);
   U21213 : NAND2_X1 port map( A1 => n8762, A2 => n29704, ZN => n20436);
   U21214 : NAND2_X1 port map( A1 => n28843, A2 => n29635, ZN => n20474);
   U21216 : XOR2_X1 port map( A1 => n28838, A2 => n8774, Z => n8773);
   U21217 : XOR2_X1 port map( A1 => n28920, A2 => n8776, Z => n8775);
   U21219 : XOR2_X1 port map( A1 => n28977, A2 => n10079, Z => n8776);
   U21224 : XOR2_X1 port map( A1 => n27662, A2 => n19953, Z => n8782);
   U21226 : OAI21_X1 port map( A1 => n22165, A2 => n8792, B => n22221, ZN => 
                           n18804);
   U21227 : XOR2_X1 port map( A1 => n37899, A2 => n35215, Z => n23975);
   U21229 : XOR2_X1 port map( A1 => n27665, A2 => n8794, Z => n8793);
   U21230 : XOR2_X1 port map( A1 => n13569, A2 => n1699, Z => n8794);
   U21232 : XOR2_X1 port map( A1 => n25215, A2 => n19800, Z => n8796);
   U21236 : NAND2_X1 port map( A1 => n8799, A2 => n21898, ZN => n17847);
   U21237 : XNOR2_X1 port map( A1 => n27540, A2 => n9013, ZN => n14986);
   U21238 : NOR2_X2 port map( A1 => n11463, A2 => n11462, ZN => n27540);
   U21242 : INV_X2 port map( I => n8812, ZN => n22368);
   U21249 : INV_X2 port map( I => n12634, ZN => n12755);
   U21251 : XOR2_X1 port map( A1 => n23802, A2 => n23803, Z => n8826);
   U21261 : NAND3_X1 port map( A1 => n15121, A2 => n9380, A3 => n34577, ZN => 
                           n25378);
   U21276 : NAND2_X1 port map( A1 => n8882, A2 => n22131, ZN => n21968);
   U21277 : AOI21_X1 port map( A1 => n36457, A2 => n31573, B => n35780, ZN => 
                           n14323);
   U21278 : XOR2_X1 port map( A1 => n38041, A2 => n29051, Z => n8885);
   U21281 : XOR2_X1 port map( A1 => n29260, A2 => n31591, Z => n8887);
   U21283 : INV_X2 port map( I => n8889, ZN => n10436);
   U21284 : XOR2_X1 port map( A1 => n4819, A2 => n1713, Z => n8890);
   U21285 : INV_X1 port map( I => Plaintext(97), ZN => n8891);
   U21286 : XOR2_X1 port map( A1 => n8891, A2 => Key(97), Z => n9552);
   U21296 : XOR2_X1 port map( A1 => n8902, A2 => n8901, Z => n8900);
   U21297 : XOR2_X1 port map( A1 => n35239, A2 => n1370, Z => n8901);
   U21300 : NAND2_X1 port map( A1 => n32419, A2 => n833, ZN => n8906);
   U21306 : INV_X2 port map( I => n14170, ZN => n14415);
   U21314 : AND2_X1 port map( A1 => n5282, A2 => n1270, Z => n24516);
   U21316 : XOR2_X1 port map( A1 => n23590, A2 => n29223, Z => n8929);
   U21319 : XOR2_X1 port map( A1 => n8939, A2 => n29206, Z => n28887);
   U21320 : AND2_X1 port map( A1 => n9745, A2 => n28508, Z => n8934);
   U21322 : NOR2_X1 port map( A1 => n1158, A2 => n8936, ZN => n20681);
   U21323 : XNOR2_X1 port map( A1 => Plaintext(31), A2 => Key(31), ZN => n8936)
                           ;
   U21324 : XOR2_X1 port map( A1 => n19991, A2 => n8938, Z => n8937);
   U21327 : XOR2_X1 port map( A1 => n23831, A2 => n19729, Z => n8938);
   U21330 : XOR2_X1 port map( A1 => n8940, A2 => n1167, Z => n13497);
   U21332 : AOI21_X1 port map( A1 => n22221, A2 => n22219, B => n9387, ZN => 
                           n8949);
   U21335 : XOR2_X1 port map( A1 => n26489, A2 => n8951, Z => n8950);
   U21336 : XOR2_X1 port map( A1 => n10621, A2 => n19835, Z => n8952);
   U21339 : XOR2_X1 port map( A1 => n37129, A2 => n28868, Z => n8957);
   U21341 : INV_X2 port map( I => n16907, ZN => n29059);
   U21344 : XOR2_X1 port map( A1 => Plaintext(79), A2 => Key(79), Z => n17209);
   U21345 : NOR2_X1 port map( A1 => n8970, A2 => n7536, ZN => n8969);
   U21348 : XOR2_X1 port map( A1 => n33083, A2 => n1010, Z => n26468);
   U21352 : XOR2_X1 port map( A1 => n27729, A2 => n17884, Z => n8974);
   U21357 : XOR2_X1 port map( A1 => n38208, A2 => n19801, Z => n8982);
   U21359 : INV_X2 port map( I => n8983, ZN => n25696);
   U21360 : XOR2_X1 port map( A1 => n15361, A2 => n17255, Z => n8983);
   U21362 : XOR2_X1 port map( A1 => n24071, A2 => n8985, Z => n12912);
   U21363 : XOR2_X1 port map( A1 => n15916, A2 => n8986, Z => n8985);
   U21364 : NAND3_X1 port map( A1 => n34379, A2 => n7916, A3 => n38246, ZN => 
                           n22032);
   U21368 : XOR2_X1 port map( A1 => n23852, A2 => n23853, Z => n9003);
   U21373 : XOR2_X1 port map( A1 => n25280, A2 => n1371, Z => n9005);
   U21376 : XOR2_X1 port map( A1 => n9010, A2 => n9009, Z => n19840);
   U21377 : XOR2_X1 port map( A1 => n22650, A2 => n22649, Z => n9009);
   U21378 : XOR2_X1 port map( A1 => n10384, A2 => n14194, Z => n9010);
   U21381 : XOR2_X1 port map( A1 => n26396, A2 => n26460, Z => n9018);
   U21383 : AOI22_X2 port map( A1 => n15554, A2 => n9021, B1 => n18744, B2 => 
                           n15553, ZN => n25160);
   U21384 : NAND2_X2 port map( A1 => n16999, A2 => n37067, ZN => n9021);
   U21385 : XOR2_X1 port map( A1 => n9023, A2 => n9022, Z => n14709);
   U21391 : NOR2_X2 port map( A1 => n16230, A2 => n16229, ZN => n18142);
   U21393 : XOR2_X1 port map( A1 => n9013, A2 => n1733, Z => n9027);
   U21394 : XOR2_X1 port map( A1 => n15653, A2 => n22441, Z => n9028);
   U21397 : XOR2_X1 port map( A1 => n9030, A2 => n35251, Z => n26293);
   U21398 : OR2_X1 port map( A1 => n24607, A2 => n29285, Z => n9032);
   U21399 : XOR2_X1 port map( A1 => n24610, A2 => n9033, Z => n13938);
   U21402 : AOI21_X1 port map( A1 => n29613, A2 => n29612, B => n9044, ZN => 
                           n29615);
   U21403 : OAI21_X2 port map( A1 => n9049, A2 => n21289, B => n9047, ZN => 
                           n29859);
   U21404 : XOR2_X1 port map( A1 => n9054, A2 => n11347, Z => n11349);
   U21406 : NOR2_X1 port map( A1 => n9062, A2 => n15411, ZN => n9058);
   U21407 : AOI21_X1 port map( A1 => n9061, A2 => n9060, B => n11226, ZN => 
                           n9059);
   U21414 : INV_X2 port map( I => n16160, ZN => n26619);
   U21417 : XOR2_X1 port map( A1 => n17519, A2 => n17516, Z => n16179);
   U21421 : XOR2_X1 port map( A1 => n9246, A2 => n15916, Z => n9247);
   U21422 : XOR2_X1 port map( A1 => n9093, A2 => n9092, Z => n9091);
   U21423 : XOR2_X1 port map( A1 => n22483, A2 => n29238, Z => n9092);
   U21424 : XOR2_X1 port map( A1 => n13596, A2 => n9095, Z => n9094);
   U21425 : XOR2_X1 port map( A1 => n25243, A2 => n19592, Z => n9095);
   U21431 : XOR2_X1 port map( A1 => n9114, A2 => n1713, Z => n10485);
   U21432 : XOR2_X1 port map( A1 => n9114, A2 => n17428, Z => n19824);
   U21433 : XOR2_X1 port map( A1 => n25093, A2 => n9113, Z => n25095);
   U21434 : XOR2_X1 port map( A1 => n9114, A2 => n25192, Z => n17555);
   U21435 : XOR2_X1 port map( A1 => n26454, A2 => n26453, Z => n9119);
   U21436 : XOR2_X1 port map( A1 => n26259, A2 => n26402, Z => n26453);
   U21438 : XOR2_X1 port map( A1 => n26456, A2 => n32528, Z => n9120);
   U21446 : XOR2_X1 port map( A1 => n17140, A2 => n655, Z => n9123);
   U21449 : NAND2_X1 port map( A1 => n1331, A2 => n18656, ZN => n14590);
   U21450 : NOR2_X1 port map( A1 => n22229, A2 => n9129, ZN => n22088);
   U21454 : AOI21_X2 port map( A1 => n1024, A2 => n25637, B => n14410, ZN => 
                           n12866);
   U21459 : XOR2_X1 port map( A1 => n27657, A2 => n27463, Z => n9139);
   U21462 : AOI21_X1 port map( A1 => n24795, A2 => n9149, B => n24646, ZN => 
                           n9148);
   U21464 : NOR2_X1 port map( A1 => n3944, A2 => n14448, ZN => n28468);
   U21468 : XOR2_X1 port map( A1 => n26532, A2 => n19407, Z => n9152);
   U21469 : XOR2_X1 port map( A1 => n39163, A2 => n19738, Z => n9153);
   U21470 : AND2_X1 port map( A1 => n26927, A2 => n735, Z => n9156);
   U21472 : XOR2_X1 port map( A1 => n9160, A2 => n16161, Z => n9159);
   U21477 : NAND2_X2 port map( A1 => n18769, A2 => n18767, ZN => n27730);
   U21484 : XOR2_X1 port map( A1 => n7475, A2 => n28821, Z => n9244);
   U21486 : INV_X1 port map( I => Plaintext(39), ZN => n9180);
   U21487 : XOR2_X1 port map( A1 => n9180, A2 => Key(39), Z => n20361);
   U21488 : NOR2_X1 port map( A1 => n15663, A2 => n1342, ZN => n21451);
   U21489 : AOI21_X1 port map( A1 => n1341, A2 => n1342, B => n32817, ZN => 
                           n13411);
   U21495 : INV_X2 port map( I => n14440, ZN => n9188);
   U21499 : XOR2_X1 port map( A1 => n33587, A2 => n30203, Z => n9195);
   U21502 : XOR2_X1 port map( A1 => n22637, A2 => n32218, Z => n9206);
   U21503 : XOR2_X1 port map( A1 => n12015, A2 => n16226, Z => n9207);
   U21508 : AOI21_X2 port map( A1 => n23909, A2 => n9909, B => n23908, ZN => 
                           n9218);
   U21512 : XOR2_X1 port map( A1 => n23920, A2 => n9220, Z => n9219);
   U21513 : XOR2_X1 port map( A1 => n23890, A2 => n1162, Z => n9220);
   U21515 : NAND2_X1 port map( A1 => n18567, A2 => n14833, ZN => n9224);
   U21517 : XOR2_X1 port map( A1 => n38165, A2 => n17428, Z => n9230);
   U21519 : INV_X2 port map( I => n9235, ZN => n19821);
   U21524 : XOR2_X1 port map( A1 => n9247, A2 => n9244, Z => n9243);
   U21534 : XOR2_X1 port map( A1 => n33197, A2 => n29657, Z => n9272);
   U21535 : XOR2_X1 port map( A1 => n22429, A2 => n22762, Z => n19342);
   U21536 : XOR2_X1 port map( A1 => n21149, A2 => n9275, Z => n9274);
   U21537 : XOR2_X1 port map( A1 => n27549, A2 => n1724, Z => n9275);
   U21538 : NAND2_X1 port map( A1 => n10589, A2 => n34786, ZN => n9278);
   U21546 : AND2_X1 port map( A1 => n31669, A2 => n25696, Z => n9292);
   U21547 : AOI21_X1 port map( A1 => n11734, A2 => n36666, B => n1103, ZN => 
                           n9294);
   U21548 : XOR2_X1 port map( A1 => n29021, A2 => n12707, Z => n11077);
   U21549 : XOR2_X1 port map( A1 => n12707, A2 => n31515, Z => n28406);
   U21550 : XOR2_X1 port map( A1 => n9299, A2 => n9298, Z => n9297);
   U21551 : XOR2_X1 port map( A1 => n26519, A2 => n1714, Z => n9298);
   U21552 : XOR2_X1 port map( A1 => n26516, A2 => n26518, Z => n9299);
   U21559 : INV_X2 port map( I => n9308, ZN => n14493);
   U21560 : XOR2_X1 port map( A1 => n25193, A2 => n29805, Z => n9309);
   U21562 : AOI21_X1 port map( A1 => n1511, A2 => n31133, B => n37378, ZN => 
                           n9312);
   U21565 : NAND2_X2 port map( A1 => n10580, A2 => n26942, ZN => n9315);
   U21567 : NOR2_X2 port map( A1 => n12122, A2 => n12121, ZN => n9920);
   U21570 : NAND2_X1 port map( A1 => n9326, A2 => n4602, ZN => n25891);
   U21574 : OAI21_X2 port map( A1 => n25644, A2 => n25361, B => n9337, ZN => 
                           n11589);
   U21575 : INV_X2 port map( I => n10686, ZN => n25644);
   U21576 : INV_X2 port map( I => n9338, ZN => n25699);
   U21577 : INV_X1 port map( I => n9698, ZN => n9340);
   U21582 : NAND3_X1 port map( A1 => n33987, A2 => n24709, A3 => n6273, ZN => 
                           n9357);
   U21586 : NAND2_X1 port map( A1 => n32891, A2 => n9371, ZN => n23799);
   U21587 : AOI21_X1 port map( A1 => n39605, A2 => n31452, B => n9371, ZN => 
                           n9821);
   U21588 : INV_X2 port map( I => n24280, ZN => n9371);
   U21590 : INV_X2 port map( I => n9373, ZN => n14389);
   U21591 : INV_X2 port map( I => n9374, ZN => n18144);
   U21594 : XOR2_X1 port map( A1 => n38149, A2 => n26567, Z => n20139);
   U21599 : XOR2_X1 port map( A1 => n9390, A2 => n24929, Z => n19742);
   U21600 : NAND2_X1 port map( A1 => n5669, A2 => n21299, ZN => n16171);
   U21601 : NAND3_X1 port map( A1 => n5414, A2 => n30238, A3 => n5669, ZN => 
                           n12232);
   U21603 : XOR2_X1 port map( A1 => n26481, A2 => n29221, Z => n9398);
   U21609 : XOR2_X1 port map( A1 => n26386, A2 => n26474, Z => n9408);
   U21612 : XOR2_X1 port map( A1 => n9411, A2 => n9410, Z => n9409);
   U21613 : XOR2_X1 port map( A1 => n26390, A2 => n29978, Z => n9410);
   U21614 : XOR2_X1 port map( A1 => n9776, A2 => n37024, Z => n9411);
   U21615 : XOR2_X1 port map( A1 => n25201, A2 => n11899, Z => n9550);
   U21617 : NOR2_X2 port map( A1 => n19740, A2 => n9413, ZN => n25996);
   U21618 : MUX2_X1 port map( I0 => n24763, I1 => n9417, S => n24691, Z => 
                           n9416);
   U21623 : XOR2_X1 port map( A1 => n18857, A2 => n9431, Z => n9430);
   U21624 : XOR2_X1 port map( A1 => n23885, A2 => n34672, Z => n9431);
   U21630 : XOR2_X1 port map( A1 => n22755, A2 => n19145, Z => n9448);
   U21631 : NAND3_X1 port map( A1 => n32050, A2 => n29794, A3 => n15867, ZN => 
                           n9457);
   U21635 : NOR2_X1 port map( A1 => n16663, A2 => n26932, ZN => n17394);
   U21636 : NOR2_X1 port map( A1 => n26933, A2 => n26932, ZN => n17392);
   U21637 : XOR2_X1 port map( A1 => n14902, A2 => n15171, Z => n9469);
   U21638 : XOR2_X1 port map( A1 => n22669, A2 => n22556, Z => n9468);
   U21643 : XOR2_X1 port map( A1 => n22503, A2 => n7432, Z => n9496);
   U21644 : XOR2_X1 port map( A1 => n22744, A2 => n35211, Z => n22616);
   U21648 : OAI21_X1 port map( A1 => n1654, A2 => n18708, B => n9507, ZN => 
                           n9506);
   U21649 : INV_X2 port map( I => n9509, ZN => n22802);
   U21652 : NAND2_X2 port map( A1 => n9513, A2 => n27121, ZN => n27776);
   U21655 : INV_X2 port map( I => n14306, ZN => n9520);
   U21657 : INV_X1 port map( I => n9529, ZN => n12624);
   U21668 : NAND2_X1 port map( A1 => n9546, A2 => n7916, ZN => n21816);
   U21669 : NAND3_X1 port map( A1 => n16888, A2 => n13632, A3 => n9546, ZN => 
                           n21815);
   U21671 : XOR2_X1 port map( A1 => n23922, A2 => n23901, Z => n9549);
   U21672 : XOR2_X1 port map( A1 => n9550, A2 => n17878, Z => n20614);
   U21673 : INV_X2 port map( I => n9552, ZN => n21869);
   U21675 : XOR2_X1 port map( A1 => n3413, A2 => n15046, Z => n9554);
   U21682 : NOR2_X2 port map( A1 => n12371, A2 => n12372, ZN => n16889);
   U21685 : OAI21_X1 port map( A1 => n9321, A2 => n14477, B => n33840, ZN => 
                           n17875);
   U21686 : XOR2_X1 port map( A1 => n9565, A2 => n9564, Z => n9563);
   U21687 : XOR2_X1 port map( A1 => n12233, A2 => n39559, Z => n9565);
   U21691 : OAI22_X2 port map( A1 => n20180, A2 => n14827, B1 => n24729, B2 => 
                           n1273, ZN => n24922);
   U21695 : NAND2_X1 port map( A1 => n28380, A2 => n7555, ZN => n28099);
   U21699 : XOR2_X1 port map( A1 => n19973, A2 => n26282, Z => n12735);
   U21703 : OR2_X1 port map( A1 => n12471, A2 => n39811, Z => n15151);
   U21705 : NOR2_X1 port map( A1 => n26813, A2 => n11138, ZN => n15352);
   U21706 : NAND3_X1 port map( A1 => n17308, A2 => n33782, A3 => n21458, ZN => 
                           n11672);
   U21713 : NAND2_X1 port map( A1 => n30156, A2 => n16786, ZN => n10210);
   U21715 : AND2_X1 port map( A1 => n26724, A2 => n14318, Z => n18225);
   U21716 : NOR2_X1 port map( A1 => n33230, A2 => n24759, ZN => n13903);
   U21719 : OR2_X1 port map( A1 => n33368, A2 => n14428, Z => n13723);
   U21724 : AND2_X1 port map( A1 => n19609, A2 => n455, Z => n21343);
   U21726 : INV_X2 port map( I => n9604, ZN => n13285);
   U21727 : XOR2_X1 port map( A1 => Plaintext(143), A2 => Key(143), Z => n9604)
                           ;
   U21730 : NAND2_X1 port map( A1 => n39140, A2 => n38198, ZN => n9605);
   U21732 : AOI21_X1 port map( A1 => n12978, A2 => n29218, B => n1378, ZN => 
                           n9607);
   U21733 : INV_X4 port map( I => n11304, ZN => n12077);
   U21734 : XNOR2_X1 port map( A1 => n28970, A2 => n20137, ZN => n9853);
   U21735 : NAND2_X1 port map( A1 => n22684, A2 => n37589, ZN => n9608);
   U21736 : NAND2_X2 port map( A1 => n21061, A2 => n21064, ZN => n23639);
   U21741 : NAND2_X1 port map( A1 => n14497, A2 => n28468, ZN => n28471);
   U21743 : XOR2_X1 port map( A1 => n25268, A2 => n814, Z => n9624);
   U21750 : OAI21_X1 port map( A1 => n32697, A2 => n9633, B => n9632, ZN => 
                           n27116);
   U21752 : NOR2_X2 port map( A1 => n27045, A2 => n27044, ZN => n27253);
   U21753 : OR2_X1 port map( A1 => n13300, A2 => n24683, Z => n14657);
   U21754 : INV_X1 port map( I => n29531, ZN => n29516);
   U21756 : XOR2_X1 port map( A1 => n18612, A2 => n35561, Z => n9643);
   U21758 : AND2_X1 port map( A1 => n19085, A2 => n38142, Z => n18611);
   U21763 : NAND2_X1 port map( A1 => n9917, A2 => n28622, ZN => n20952);
   U21774 : AND2_X1 port map( A1 => n28576, A2 => n35199, Z => n28177);
   U21783 : XOR2_X1 port map( A1 => n25196, A2 => n19670, Z => n24958);
   U21789 : NOR2_X1 port map( A1 => n15256, A2 => n24359, ZN => n10439);
   U21790 : AND3_X1 port map( A1 => n16154, A2 => n28141, A3 => n281, Z => 
                           n15975);
   U21791 : XOR2_X1 port map( A1 => n22713, A2 => n22195, Z => n22203);
   U21800 : XOR2_X1 port map( A1 => n39636, A2 => n23841, Z => n16697);
   U21803 : NAND2_X2 port map( A1 => n10349, A2 => n11705, ZN => n28313);
   U21809 : XOR2_X1 port map( A1 => n11810, A2 => n11809, Z => n9687);
   U21810 : XOR2_X1 port map( A1 => n26597, A2 => n19627, Z => n19772);
   U21831 : INV_X1 port map( I => n6523, ZN => n10904);
   U21837 : XOR2_X1 port map( A1 => n12157, A2 => n28100, Z => n9712);
   U21839 : NOR2_X2 port map( A1 => n10174, A2 => n23582, ZN => n23508);
   U21845 : XOR2_X1 port map( A1 => n10113, A2 => n20279, Z => n20891);
   U21846 : NAND2_X1 port map( A1 => n16854, A2 => n16855, ZN => n12385);
   U21848 : XOR2_X1 port map( A1 => n20454, A2 => n29887, Z => n19766);
   U21849 : NAND2_X2 port map( A1 => n948, A2 => n26660, ZN => n27141);
   U21852 : AND2_X1 port map( A1 => n12032, A2 => n7575, Z => n13157);
   U21857 : XOR2_X1 port map( A1 => n9732, A2 => n27536, Z => n12104);
   U21862 : INV_X2 port map( I => n9737, ZN => n13998);
   U21863 : XOR2_X1 port map( A1 => Plaintext(179), A2 => Key(179), Z => n9737)
                           ;
   U21865 : OR2_X1 port map( A1 => n32105, A2 => n25349, Z => n12923);
   U21873 : INV_X1 port map( I => n10012, ZN => n24678);
   U21875 : INV_X1 port map( I => n10847, ZN => n10846);
   U21887 : XOR2_X1 port map( A1 => n36039, A2 => n721, Z => n12000);
   U21903 : XOR2_X1 port map( A1 => n9766, A2 => n25226, Z => n13575);
   U21904 : XOR2_X1 port map( A1 => n25323, A2 => n25006, Z => n9766);
   U21909 : NOR2_X1 port map( A1 => n15420, A2 => n14869, ZN => n15419);
   U21910 : INV_X1 port map( I => n13219, ZN => n10754);
   U21917 : INV_X2 port map( I => n9780, ZN => n16836);
   U21923 : NOR2_X1 port map( A1 => n21071, A2 => n21069, ZN => n29539);
   U21932 : INV_X2 port map( I => n19313, ZN => n20476);
   U21934 : NAND2_X1 port map( A1 => n15003, A2 => n26092, ZN => n25883);
   U21938 : INV_X2 port map( I => n9813, ZN => n10334);
   U21939 : XOR2_X1 port map( A1 => n22233, A2 => n22232, Z => n9813);
   U21941 : XOR2_X1 port map( A1 => n17987, A2 => n12806, Z => n12805);
   U21942 : XOR2_X1 port map( A1 => n13155, A2 => n29337, Z => n13154);
   U21951 : XOR2_X1 port map( A1 => Plaintext(4), A2 => Key(4), Z => n12225);
   U21954 : OAI22_X1 port map( A1 => n7876, A2 => n7284, B1 => n19637, B2 => 
                           n1256, ZN => n25352);
   U21957 : XOR2_X1 port map( A1 => n9829, A2 => n10027, Z => Ciphertext(150));
   U21958 : OAI22_X1 port map( A1 => n30084, A2 => n30093, B1 => n30086, B2 => 
                           n30083, ZN => n9829);
   U21962 : AND2_X1 port map( A1 => n1548, A2 => n10882, Z => n14625);
   U21964 : NOR2_X2 port map( A1 => n16078, A2 => n16076, ZN => n24925);
   U21969 : XOR2_X1 port map( A1 => n18447, A2 => n18449, Z => n9845);
   U21973 : NOR2_X1 port map( A1 => n13646, A2 => n29359, ZN => n9857);
   U21975 : OAI21_X2 port map( A1 => n22634, A2 => n12243, B => n12242, ZN => 
                           n18751);
   U21977 : AND3_X1 port map( A1 => n914, A2 => n14558, A3 => n20313, Z => 
                           n11758);
   U21979 : XOR2_X1 port map( A1 => n9852, A2 => n14867, Z => n14866);
   U21980 : XOR2_X1 port map( A1 => n37024, A2 => n36171, Z => n9852);
   U21984 : XNOR2_X1 port map( A1 => n22717, A2 => n37094, ZN => n14109);
   U21988 : INV_X2 port map( I => n15621, ZN => n29452);
   U21989 : XOR2_X1 port map( A1 => n20135, A2 => n9853, Z => n15621);
   U21990 : XOR2_X1 port map( A1 => n12300, A2 => n26400, Z => n20098);
   U21992 : XOR2_X1 port map( A1 => n15011, A2 => n25100, Z => n14859);
   U21996 : XOR2_X1 port map( A1 => n9857, A2 => n29360, Z => Ciphertext(31));
   U22001 : OAI22_X1 port map( A1 => n9865, A2 => n14417, B1 => n29596, B2 => 
                           n31667, ZN => n28585);
   U22004 : NOR2_X2 port map( A1 => n13000, A2 => n9869, ZN => n12726);
   U22008 : NOR2_X2 port map( A1 => n21401, A2 => n21645, ZN => n9886);
   U22012 : NAND2_X2 port map( A1 => n3293, A2 => n21895, ZN => n21582);
   U22018 : XOR2_X1 port map( A1 => n14986, A2 => n754, Z => n27827);
   U22020 : XOR2_X1 port map( A1 => n29002, A2 => n20324, Z => n20323);
   U22024 : XOR2_X1 port map( A1 => n35227, A2 => n16613, Z => n9887);
   U22026 : XOR2_X1 port map( A1 => n26259, A2 => n29711, Z => n16427);
   U22027 : NAND2_X2 port map( A1 => n9891, A2 => n10535, ZN => n27407);
   U22028 : INV_X2 port map( I => n9895, ZN => n14636);
   U22029 : XOR2_X1 port map( A1 => n16425, A2 => n16423, Z => n9895);
   U22031 : XOR2_X1 port map( A1 => Plaintext(73), A2 => Key(73), Z => n20778);
   U22037 : XNOR2_X1 port map( A1 => n22450, A2 => n22451, ZN => n13667);
   U22039 : XOR2_X1 port map( A1 => n10225, A2 => n1356, Z => n11902);
   U22041 : NAND2_X1 port map( A1 => n13107, A2 => n10803, ZN => n9907);
   U22044 : NOR2_X1 port map( A1 => n19310, A2 => n29262, ZN => n19475);
   U22045 : XOR2_X1 port map( A1 => n11437, A2 => n22522, Z => n9911);
   U22048 : AND2_X1 port map( A1 => n18451, A2 => n14451, Z => n14484);
   U22049 : AND2_X1 port map( A1 => n27150, A2 => n20740, Z => n26966);
   U22059 : XOR2_X1 port map( A1 => n25245, A2 => n25187, Z => n10928);
   U22065 : XOR2_X1 port map( A1 => n35532, A2 => n37094, Z => n9937);
   U22067 : NAND2_X1 port map( A1 => n20997, A2 => n31586, ZN => n9988);
   U22068 : AND2_X1 port map( A1 => n13370, A2 => n32377, Z => n23583);
   U22069 : XNOR2_X1 port map( A1 => Key(18), A2 => Plaintext(18), ZN => n9942)
                           ;
   U22071 : NAND2_X1 port map( A1 => n17965, A2 => n13257, ZN => n15803);
   U22072 : XOR2_X1 port map( A1 => n1412, A2 => n38150, Z => n18493);
   U22074 : OAI22_X1 port map( A1 => n21507, A2 => n21509, B1 => n21484, B2 => 
                           n21593, ZN => n21485);
   U22080 : XOR2_X1 port map( A1 => n736, A2 => n11989, Z => n9948);
   U22088 : XOR2_X1 port map( A1 => n15581, A2 => n15181, Z => n9952);
   U22089 : XOR2_X1 port map( A1 => n9953, A2 => n29887, Z => Ciphertext(124));
   U22093 : NOR2_X1 port map( A1 => n34049, A2 => n21626, ZN => n21627);
   U22095 : NAND3_X1 port map( A1 => n29621, A2 => n29622, A3 => n29627, ZN => 
                           n9957);
   U22100 : NOR2_X2 port map( A1 => n10041, A2 => n11544, ZN => n9959);
   U22102 : XOR2_X1 port map( A1 => n9960, A2 => n20824, Z => n11856);
   U22108 : XOR2_X1 port map( A1 => n9967, A2 => n29109, Z => Ciphertext(0));
   U22109 : OAI21_X1 port map( A1 => n10681, A2 => n1681, B => n6361, ZN => 
                           n10979);
   U22110 : XOR2_X1 port map( A1 => n14638, A2 => n29245, Z => n14136);
   U22113 : XOR2_X1 port map( A1 => Plaintext(14), A2 => Key(14), Z => n10925);
   U22115 : INV_X2 port map( I => n9973, ZN => n14422);
   U22116 : XOR2_X1 port map( A1 => n19443, A2 => n750, Z => n18973);
   U22121 : XOR2_X1 port map( A1 => n37044, A2 => n14651, Z => n9976);
   U22124 : XOR2_X1 port map( A1 => n1555, A2 => n15625, Z => n9977);
   U22125 : XOR2_X1 port map( A1 => n12282, A2 => n22501, Z => n9980);
   U22133 : XOR2_X1 port map( A1 => n9986, A2 => n823, Z => n11046);
   U22136 : NAND2_X1 port map( A1 => n9991, A2 => n9990, ZN => n28264);
   U22137 : INV_X1 port map( I => n9992, ZN => n9991);
   U22138 : AOI21_X1 port map( A1 => n28048, A2 => n28255, B => n28258, ZN => 
                           n9992);
   U22140 : BUF_X2 port map( I => n29493, Z => n9993);
   U22141 : XOR2_X1 port map( A1 => n33322, A2 => n7917, Z => n23848);
   U22143 : XNOR2_X1 port map( A1 => n35245, A2 => n25274, ZN => n10644);
   U22145 : XOR2_X1 port map( A1 => n1259, A2 => n10791, Z => n24914);
   U22149 : NAND3_X2 port map( A1 => n14903, A2 => n5795, A3 => n14904, ZN => 
                           n16798);
   U22154 : XOR2_X1 port map( A1 => n19002, A2 => n10001, Z => n19001);
   U22155 : XOR2_X1 port map( A1 => n18751, A2 => n658, Z => n10001);
   U22158 : XNOR2_X1 port map( A1 => n26343, A2 => n19099, ZN => n10230);
   U22167 : AND2_X1 port map( A1 => n19941, A2 => n36794, Z => n17304);
   U22170 : XOR2_X1 port map( A1 => n10583, A2 => n10585, Z => n10584);
   U22171 : XOR2_X1 port map( A1 => n23688, A2 => n23849, Z => n10014);
   U22172 : NAND2_X1 port map( A1 => n16567, A2 => n13851, ZN => n13600);
   U22174 : XOR2_X1 port map( A1 => n11620, A2 => n11621, Z => n19423);
   U22175 : XOR2_X1 port map( A1 => n22506, A2 => n11230, Z => n15218);
   U22183 : XOR2_X1 port map( A1 => n22622, A2 => n33990, Z => n15610);
   U22186 : AOI22_X1 port map( A1 => n10031, A2 => n30139, B1 => n19098, B2 => 
                           n30138, ZN => n30140);
   U22188 : OR2_X1 port map( A1 => n13786, A2 => n11700, Z => n11022);
   U22189 : XOR2_X1 port map( A1 => n13229, A2 => n1469, Z => n10036);
   U22193 : XOR2_X1 port map( A1 => n14388, A2 => n21097, Z => n21096);
   U22196 : XOR2_X1 port map( A1 => n28662, A2 => n10040, Z => n13234);
   U22197 : XNOR2_X1 port map( A1 => n15270, A2 => n29067, ZN => n11127);
   U22202 : NOR2_X1 port map( A1 => n27152, A2 => n19750, ZN => n10393);
   U22204 : XOR2_X1 port map( A1 => n29128, A2 => n29107, Z => n11946);
   U22217 : INV_X1 port map( I => n27252, ZN => n18717);
   U22220 : AND2_X1 port map( A1 => n34561, A2 => n12612, Z => n16779);
   U22221 : OAI21_X1 port map( A1 => n34007, A2 => n32146, B => n10058, ZN => 
                           n28342);
   U22223 : NAND2_X1 port map( A1 => n28068, A2 => n28067, ZN => n13512);
   U22224 : XOR2_X1 port map( A1 => n29836, A2 => n29839, Z => n10059);
   U22226 : AOI21_X1 port map( A1 => n28634, A2 => n28635, B => n28633, ZN => 
                           n10061);
   U22231 : XOR2_X1 port map( A1 => n25257, A2 => n642, Z => n10070);
   U22233 : XOR2_X1 port map( A1 => n12356, A2 => n12354, Z => n14405);
   U22239 : NAND3_X2 port map( A1 => n18125, A2 => n21004, A3 => n28627, ZN => 
                           n10080);
   U22241 : XOR2_X1 port map( A1 => n29037, A2 => n10087, Z => n11747);
   U22242 : NAND2_X1 port map( A1 => n27138, A2 => n18074, ZN => n18073);
   U22245 : XOR2_X1 port map( A1 => n19289, A2 => n33866, Z => n14569);
   U22246 : XOR2_X1 port map( A1 => n29140, A2 => n19078, Z => n10391);
   U22248 : NAND3_X1 port map( A1 => n1202, A2 => n15704, A3 => n11676, ZN => 
                           n15446);
   U22253 : NAND2_X1 port map( A1 => n20965, A2 => n37306, ZN => n26052);
   U22265 : NOR2_X1 port map( A1 => n24814, A2 => n21231, ZN => n10114);
   U22267 : XOR2_X1 port map( A1 => Plaintext(17), A2 => Key(17), Z => n11576);
   U22269 : XOR2_X1 port map( A1 => n33178, A2 => n1165, Z => n10131);
   U22270 : XOR2_X1 port map( A1 => n10136, A2 => n10134, Z => n10679);
   U22276 : XOR2_X1 port map( A1 => n11724, A2 => n11725, Z => n14471);
   U22278 : INV_X2 port map( I => n10155, ZN => n19424);
   U22285 : AOI21_X1 port map( A1 => n21322, A2 => n28119, B => n28139, ZN => 
                           n10167);
   U22289 : XOR2_X1 port map( A1 => n27496, A2 => n12351, Z => n10169);
   U22291 : INV_X2 port map( I => n12950, ZN => n24274);
   U22292 : XOR2_X1 port map( A1 => n10182, A2 => n10181, Z => n12950);
   U22294 : XOR2_X1 port map( A1 => n21227, A2 => n18683, Z => n10182);
   U22298 : XOR2_X1 port map( A1 => n10189, A2 => n29223, Z => Ciphertext(10));
   U22302 : XOR2_X1 port map( A1 => n10197, A2 => n10196, Z => n10195);
   U22303 : XOR2_X1 port map( A1 => n35953, A2 => n19833, Z => n10196);
   U22304 : XOR2_X1 port map( A1 => n37312, A2 => n25226, Z => n10197);
   U22305 : XOR2_X1 port map( A1 => n10201, A2 => n16458, Z => n10200);
   U22307 : XOR2_X1 port map( A1 => Plaintext(177), A2 => Key(177), Z => n10212
                           );
   U22308 : NOR2_X1 port map( A1 => n21730, A2 => n9863, ZN => n21731);
   U22310 : XOR2_X1 port map( A1 => n7287, A2 => n19516, Z => n10214);
   U22314 : XOR2_X1 port map( A1 => n27539, A2 => n27826, Z => n10226);
   U22327 : XOR2_X1 port map( A1 => n10240, A2 => n27761, Z => n10673);
   U22328 : XOR2_X1 port map( A1 => n27664, A2 => n19616, Z => n10240);
   U22331 : AOI21_X1 port map( A1 => n17411, A2 => n22252, B => n10242, ZN => 
                           n17408);
   U22332 : XOR2_X1 port map( A1 => n10243, A2 => n10245, Z => n26666);
   U22333 : XOR2_X1 port map( A1 => n21034, A2 => n10244, Z => n10243);
   U22335 : XOR2_X1 port map( A1 => n19760, A2 => n33194, Z => n10244);
   U22336 : XOR2_X1 port map( A1 => n10246, A2 => n26085, Z => n10245);
   U22337 : XOR2_X1 port map( A1 => n12934, A2 => n26518, Z => n10246);
   U22338 : INV_X2 port map( I => n10247, ZN => n20077);
   U22339 : NAND2_X1 port map( A1 => n38725, A2 => n20077, ZN => n19054);
   U22340 : XOR2_X1 port map( A1 => n17706, A2 => n10250, Z => n10248);
   U22341 : XOR2_X1 port map( A1 => n25149, A2 => n19670, Z => n10250);
   U22342 : INV_X2 port map( I => n10251, ZN => n24271);
   U22343 : XOR2_X1 port map( A1 => n24064, A2 => n23073, Z => n10252);
   U22349 : XOR2_X1 port map( A1 => n10258, A2 => n12357, Z => n12356);
   U22355 : XOR2_X1 port map( A1 => n22749, A2 => n29647, Z => n10267);
   U22356 : XOR2_X1 port map( A1 => n18595, A2 => n22580, Z => n10268);
   U22358 : XOR2_X1 port map( A1 => n24033, A2 => n10276, Z => n10275);
   U22359 : XOR2_X1 port map( A1 => n19656, A2 => n30248, Z => n10276);
   U22361 : XOR2_X1 port map( A1 => n24022, A2 => n10279, Z => n10278);
   U22362 : XOR2_X1 port map( A1 => n23933, A2 => n15202, Z => n24022);
   U22363 : NAND2_X1 port map( A1 => n1084, A2 => n35750, ZN => n17900);
   U22364 : INV_X2 port map( I => n10282, ZN => n12953);
   U22369 : XOR2_X1 port map( A1 => n17937, A2 => n23968, Z => n12799);
   U22370 : NAND2_X2 port map( A1 => n15073, A2 => n23228, ZN => n23968);
   U22375 : XOR2_X1 port map( A1 => n32931, A2 => n35318, Z => n13750);
   U22387 : XOR2_X1 port map( A1 => n10319, A2 => n10318, Z => n10315);
   U22389 : XOR2_X1 port map( A1 => n26584, A2 => n29474, Z => n10318);
   U22392 : INV_X1 port map( I => n22209, ZN => n22207);
   U22394 : OAI21_X2 port map( A1 => n10325, A2 => n21759, B => n10324, ZN => 
                           n22354);
   U22395 : NAND2_X2 port map( A1 => n19650, A2 => n21697, ZN => n21759);
   U22397 : XOR2_X1 port map( A1 => n35222, A2 => n1730, Z => n10328);
   U22398 : XOR2_X1 port map( A1 => n10333, A2 => n10330, Z => n20595);
   U22399 : XOR2_X1 port map( A1 => n10332, A2 => n10331, Z => n10330);
   U22400 : XOR2_X1 port map( A1 => n25182, A2 => n34848, Z => n10331);
   U22401 : XOR2_X1 port map( A1 => n6727, A2 => n25181, Z => n10332);
   U22405 : XOR2_X1 port map( A1 => n30856, A2 => n10343, Z => n28854);
   U22407 : INV_X2 port map( I => n20883, ZN => n21270);
   U22412 : XOR2_X1 port map( A1 => n39548, A2 => n30063, Z => n10364);
   U22415 : XOR2_X1 port map( A1 => n10371, A2 => n16029, Z => n10636);
   U22421 : XOR2_X1 port map( A1 => n10387, A2 => n10386, Z => n23992);
   U22422 : XOR2_X1 port map( A1 => n15777, A2 => n10389, Z => n10386);
   U22423 : XOR2_X1 port map( A1 => n23981, A2 => n10388, Z => n10387);
   U22424 : XOR2_X1 port map( A1 => n36143, A2 => n35181, Z => n10388);
   U22425 : XOR2_X1 port map( A1 => n23982, A2 => n19498, Z => n10389);
   U22427 : AOI21_X2 port map( A1 => n10394, A2 => n27063, B => n27062, ZN => 
                           n28537);
   U22432 : XOR2_X1 port map( A1 => n10400, A2 => n11464, Z => n10534);
   U22434 : XOR2_X1 port map( A1 => n10402, A2 => n24005, Z => n10401);
   U22436 : XOR2_X1 port map( A1 => n25161, A2 => n14687, Z => n10406);
   U22438 : NAND2_X1 port map( A1 => n30171, A2 => n30177, ZN => n10410);
   U22439 : XOR2_X1 port map( A1 => n10412, A2 => n18927, Z => n27784);
   U22444 : XOR2_X1 port map( A1 => n37094, A2 => n22621, Z => n15608);
   U22446 : XOR2_X1 port map( A1 => n18857, A2 => n663, Z => n10426);
   U22450 : OAI21_X1 port map( A1 => n29220, A2 => n29222, B => n9914, ZN => 
                           n10428);
   U22451 : XOR2_X1 port map( A1 => n10430, A2 => n20560, Z => n10658);
   U22452 : XOR2_X1 port map( A1 => n12534, A2 => n19933, Z => n10431);
   U22458 : XOR2_X1 port map( A1 => n12251, A2 => n19131, Z => n10447);
   U22462 : NAND3_X1 port map( A1 => n21599, A2 => n16305, A3 => n21870, ZN => 
                           n10649);
   U22467 : INV_X2 port map( I => n10455, ZN => n23198);
   U22469 : OAI21_X1 port map( A1 => n10051, A2 => n10461, B => n20133, ZN => 
                           n16966);
   U22470 : NOR2_X1 port map( A1 => n10461, A2 => n27428, ZN => n26941);
   U22475 : XOR2_X1 port map( A1 => n10884, A2 => n10885, Z => n10478);
   U22477 : XOR2_X1 port map( A1 => n17284, A2 => n708, Z => n10482);
   U22480 : XOR2_X1 port map( A1 => n20304, A2 => n25291, Z => n10486);
   U22482 : XOR2_X1 port map( A1 => n26258, A2 => n38502, Z => n26385);
   U22483 : XOR2_X1 port map( A1 => n14386, A2 => n10493, Z => n11661);
   U22484 : XOR2_X1 port map( A1 => n11098, A2 => n29337, Z => n10493);
   U22487 : XOR2_X1 port map( A1 => n16743, A2 => n27785, Z => n27494);
   U22489 : XOR2_X1 port map( A1 => n22541, A2 => n669, Z => n10502);
   U22494 : INV_X1 port map( I => n24829, ZN => n18654);
   U22495 : XOR2_X1 port map( A1 => n17935, A2 => n845, Z => n10523);
   U22498 : INV_X2 port map( I => n10534, ZN => n13444);
   U22500 : XOR2_X1 port map( A1 => n32931, A2 => n19950, Z => n10538);
   U22506 : XOR2_X1 port map( A1 => n10541, A2 => n15071, Z => n29495);
   U22507 : OAI21_X1 port map( A1 => n37804, A2 => n36827, B => n10542, ZN => 
                           n14362);
   U22508 : NOR2_X1 port map( A1 => n28690, A2 => n36827, ZN => n28691);
   U22510 : XOR2_X1 port map( A1 => n23898, A2 => n23779, Z => n10548);
   U22512 : XOR2_X1 port map( A1 => n23781, A2 => n12107, Z => n10549);
   U22518 : XOR2_X1 port map( A1 => n13083, A2 => n10561, Z => n13082);
   U22519 : XOR2_X1 port map( A1 => n10562, A2 => n27638, Z => n10561);
   U22520 : XOR2_X1 port map( A1 => n34345, A2 => n29875, Z => n20047);
   U22521 : XOR2_X1 port map( A1 => n37466, A2 => n1717, Z => n15214);
   U22522 : XOR2_X1 port map( A1 => n2383, A2 => n34345, Z => n22432);
   U22531 : XOR2_X1 port map( A1 => n10586, A2 => n664, Z => n10585);
   U22532 : XOR2_X1 port map( A1 => n1554, A2 => n24927, Z => n10586);
   U22537 : XOR2_X1 port map( A1 => n33216, A2 => n26334, Z => n10593);
   U22539 : XOR2_X1 port map( A1 => n29093, A2 => n29146, Z => n29065);
   U22540 : NAND2_X2 port map( A1 => n10596, A2 => n20430, ZN => n29146);
   U22543 : INV_X2 port map( I => n14061, ZN => n14408);
   U22544 : XOR2_X1 port map( A1 => n10599, A2 => n10597, Z => n14061);
   U22545 : XOR2_X1 port map( A1 => n26204, A2 => n10598, Z => n10597);
   U22547 : XOR2_X1 port map( A1 => n26150, A2 => n16998, Z => n10599);
   U22552 : XOR2_X1 port map( A1 => n10616, A2 => n25027, Z => n10615);
   U22554 : INV_X1 port map( I => n25959, ZN => n25334);
   U22556 : XOR2_X1 port map( A1 => n10620, A2 => n10619, Z => n24307);
   U22557 : XOR2_X1 port map( A1 => n24045, A2 => n24048, Z => n10619);
   U22558 : XOR2_X1 port map( A1 => n33690, A2 => n27736, Z => n10706);
   U22561 : NAND2_X2 port map( A1 => n21884, A2 => n13856, ZN => n22042);
   U22566 : XNOR2_X1 port map( A1 => Plaintext(96), A2 => Key(96), ZN => n10629
                           );
   U22580 : XNOR2_X1 port map( A1 => Plaintext(100), A2 => Key(100), ZN => 
                           n10656);
   U22582 : MUX2_X1 port map( I0 => n11034, I1 => n2678, S => n910, Z => n11036
                           );
   U22583 : XOR2_X1 port map( A1 => n19956, A2 => n10663, Z => n10662);
   U22584 : XOR2_X1 port map( A1 => n30322, A2 => n19717, Z => n10663);
   U22585 : NOR2_X1 port map( A1 => n15282, A2 => n10667, ZN => n12409);
   U22589 : XOR2_X1 port map( A1 => n17937, A2 => n1366, Z => n10684);
   U22593 : XOR2_X1 port map( A1 => n13245, A2 => n27534, Z => n10707);
   U22594 : XOR2_X1 port map( A1 => n35268, A2 => n19910, Z => n11401);
   U22595 : XOR2_X1 port map( A1 => n1614, A2 => n35181, Z => n22957);
   U22596 : XOR2_X1 port map( A1 => n10717, A2 => n10714, Z => n21031);
   U22597 : XOR2_X1 port map( A1 => n10715, A2 => n10716, Z => n10714);
   U22598 : XOR2_X1 port map( A1 => n35268, A2 => n20748, Z => n10715);
   U22599 : XOR2_X1 port map( A1 => n7250, A2 => n19096, Z => n10716);
   U22600 : INV_X1 port map( I => n33178, ZN => n10718);
   U22601 : XOR2_X1 port map( A1 => n36596, A2 => n19674, Z => n22518);
   U22606 : OAI21_X1 port map( A1 => n31564, A2 => n38839, B => n20864, ZN => 
                           n23962);
   U22609 : XOR2_X1 port map( A1 => n10737, A2 => n14101, Z => n14170);
   U22611 : AOI21_X1 port map( A1 => n22045, A2 => n38448, B => n10743, ZN => 
                           n10742);
   U22614 : XOR2_X1 port map( A1 => n14023, A2 => n18992, Z => n10748);
   U22618 : XOR2_X1 port map( A1 => n8402, A2 => n1051, Z => n10766);
   U22626 : OR2_X1 port map( A1 => n24872, A2 => n31161, Z => n10773);
   U22629 : NAND2_X1 port map( A1 => n21256, A2 => n9178, ZN => n21255);
   U22632 : XOR2_X1 port map( A1 => n39320, A2 => n25086, Z => n15126);
   U22636 : XOR2_X1 port map( A1 => n38950, A2 => n10791, Z => n25000);
   U22637 : XOR2_X1 port map( A1 => n10791, A2 => n19808, Z => n19986);
   U22638 : XOR2_X1 port map( A1 => n10797, A2 => n16783, Z => n11503);
   U22641 : OAI21_X1 port map( A1 => n13107, A2 => n10803, B => n29224, ZN => 
                           n29226);
   U22646 : INV_X2 port map( I => n10810, ZN => n12235);
   U22647 : INV_X2 port map( I => n16931, ZN => n18164);
   U22649 : INV_X2 port map( I => n10816, ZN => n14158);
   U22650 : XOR2_X1 port map( A1 => n27757, A2 => n12769, Z => n10819);
   U22652 : XOR2_X1 port map( A1 => n26441, A2 => n29857, Z => n10823);
   U22653 : XOR2_X1 port map( A1 => n26438, A2 => n6131, Z => n26523);
   U22654 : XOR2_X1 port map( A1 => n28928, A2 => n10830, Z => n10829);
   U22655 : XOR2_X1 port map( A1 => n28927, A2 => n10794, Z => n10830);
   U22656 : AOI21_X1 port map( A1 => n10831, A2 => n17750, B => n17748, ZN => 
                           n17747);
   U22657 : NOR2_X1 port map( A1 => n39454, A2 => n32979, ZN => n25749);
   U22658 : INV_X2 port map( I => n10835, ZN => n11150);
   U22662 : XOR2_X1 port map( A1 => n26450, A2 => n17858, Z => n10855);
   U22663 : XOR2_X1 port map( A1 => n22688, A2 => n10859, Z => n10858);
   U22664 : XOR2_X1 port map( A1 => n5203, A2 => n19843, Z => n10859);
   U22668 : XOR2_X1 port map( A1 => n27606, A2 => n10864, Z => n10863);
   U22669 : XOR2_X1 port map( A1 => n27776, A2 => n29849, Z => n10864);
   U22673 : XOR2_X1 port map( A1 => n3649, A2 => n35169, Z => n25044);
   U22674 : XOR2_X1 port map( A1 => n32195, A2 => n3649, Z => n17879);
   U22675 : XOR2_X1 port map( A1 => n10872, A2 => n10874, Z => n13248);
   U22679 : XOR2_X1 port map( A1 => n9344, A2 => n23996, Z => n10874);
   U22686 : XOR2_X1 port map( A1 => n21093, A2 => n1367, Z => n27808);
   U22687 : XOR2_X1 port map( A1 => n27858, A2 => n21093, Z => n15068);
   U22688 : XOR2_X1 port map( A1 => n21093, A2 => n27781, Z => n27615);
   U22689 : XOR2_X1 port map( A1 => n39636, A2 => n1375, Z => n10884);
   U22691 : XOR2_X1 port map( A1 => n20509, A2 => n33452, Z => n10887);
   U22696 : XOR2_X1 port map( A1 => n10898, A2 => n764, Z => n10897);
   U22697 : XOR2_X1 port map( A1 => n33961, A2 => n35249, Z => n10898);
   U22699 : XOR2_X1 port map( A1 => n25247, A2 => n29554, Z => n10905);
   U22706 : INV_X2 port map( I => n10925, ZN => n18450);
   U22711 : INV_X1 port map( I => Plaintext(59), ZN => n10929);
   U22713 : NOR2_X1 port map( A1 => n1416, A2 => n2022, ZN => n18701);
   U22714 : AOI22_X1 port map( A1 => n33100, A2 => n9597, B1 => n18571, B2 => 
                           n20197, ZN => n28409);
   U22728 : XOR2_X1 port map( A1 => n17999, A2 => n656, Z => n10955);
   U22730 : XOR2_X1 port map( A1 => n23774, A2 => n23680, Z => n10957);
   U22735 : XOR2_X1 port map( A1 => n10967, A2 => n10966, Z => n18933);
   U22736 : XOR2_X1 port map( A1 => n26222, A2 => n18934, Z => n10966);
   U22737 : XOR2_X1 port map( A1 => n10965, A2 => n26359, Z => n26222);
   U22740 : OR2_X1 port map( A1 => n19159, A2 => n10979, Z => n19158);
   U22743 : XOR2_X1 port map( A1 => n13374, A2 => n11755, Z => n10983);
   U22744 : XOR2_X1 port map( A1 => n27807, A2 => n27808, Z => n10984);
   U22746 : XOR2_X1 port map( A1 => n10987, A2 => n29474, Z => n24929);
   U22747 : XOR2_X1 port map( A1 => n10987, A2 => n16460, Z => n17836);
   U22750 : XOR2_X1 port map( A1 => n18180, A2 => n30114, Z => n13064);
   U22760 : XOR2_X1 port map( A1 => n15617, A2 => n29300, Z => n11016);
   U22765 : NOR2_X1 port map( A1 => n25533, A2 => n9594, ZN => n11018);
   U22768 : NOR2_X1 port map( A1 => n11020, A2 => n15135, ZN => n27589);
   U22773 : XOR2_X1 port map( A1 => n27697, A2 => n27503, Z => n27826);
   U22775 : NOR2_X1 port map( A1 => n30758, A2 => n17095, ZN => n11043);
   U22776 : INV_X2 port map( I => n11046, ZN => n19696);
   U22781 : NAND2_X2 port map( A1 => n21242, A2 => n21241, ZN => n17986);
   U22787 : AOI21_X1 port map( A1 => n15958, A2 => n12943, B => n11067, ZN => 
                           n15956);
   U22789 : XOR2_X1 port map( A1 => n12393, A2 => n29857, Z => n14505);
   U22792 : XOR2_X1 port map( A1 => Plaintext(153), A2 => Key(153), Z => n15009
                           );
   U22794 : XOR2_X1 port map( A1 => n29090, A2 => n11075, Z => n11074);
   U22795 : XOR2_X1 port map( A1 => n296, A2 => n29808, Z => n11075);
   U22796 : XOR2_X1 port map( A1 => n29022, A2 => n11077, Z => n11076);
   U22798 : INV_X1 port map( I => n24152, ZN => n21148);
   U22799 : XOR2_X1 port map( A1 => n11372, A2 => n24011, Z => n23915);
   U22800 : XOR2_X1 port map( A1 => n11372, A2 => n19947, Z => n17725);
   U22804 : XNOR2_X1 port map( A1 => n16742, A2 => n16740, ZN => n11084);
   U22806 : OAI21_X2 port map( A1 => n27902, A2 => n21020, B => n16994, ZN => 
                           n28689);
   U22807 : XOR2_X1 port map( A1 => n11098, A2 => n29411, Z => n23316);
   U22808 : XOR2_X1 port map( A1 => n23695, A2 => n11098, Z => n15974);
   U22810 : XOR2_X1 port map( A1 => n11102, A2 => n25075, Z => n11103);
   U22814 : XOR2_X1 port map( A1 => n11115, A2 => n23977, Z => n11114);
   U22819 : NOR2_X1 port map( A1 => n11120, A2 => n16619, ZN => n18971);
   U22821 : NAND2_X1 port map( A1 => n25998, A2 => n39165, ZN => n25842);
   U22831 : NAND2_X1 port map( A1 => n20328, A2 => n11146, ZN => n17219);
   U22832 : XOR2_X1 port map( A1 => n16254, A2 => n649, Z => n22412);
   U22834 : NAND3_X2 port map( A1 => n16028, A2 => n21998, A3 => n18401, ZN => 
                           n22644);
   U22836 : OAI22_X2 port map( A1 => n12546, A2 => n11239, B1 => n11238, B2 => 
                           n543, ZN => n11149);
   U22837 : NOR2_X1 port map( A1 => n11149, A2 => n19515, ZN => n13899);
   U22838 : XOR2_X1 port map( A1 => n28966, A2 => n28968, Z => n11151);
   U22840 : XOR2_X1 port map( A1 => n679, A2 => n11153, Z => n11152);
   U22841 : XOR2_X1 port map( A1 => n10129, A2 => n11155, Z => n11154);
   U22845 : XOR2_X1 port map( A1 => n11267, A2 => n722, Z => n11165);
   U22852 : OAI21_X2 port map( A1 => n14189, A2 => n14188, B => n14186, ZN => 
                           n17511);
   U22858 : XOR2_X1 port map( A1 => n11200, A2 => Plaintext(178), Z => n13996);
   U22860 : XOR2_X1 port map( A1 => n11201, A2 => n3953, Z => n22694);
   U22866 : XOR2_X1 port map( A1 => n27865, A2 => n11211, Z => n11210);
   U22867 : XOR2_X1 port map( A1 => n20454, A2 => n27738, Z => n11211);
   U22871 : INV_X1 port map( I => n11214, ZN => n18746);
   U22872 : NAND2_X2 port map( A1 => n11218, A2 => n11217, ZN => n17192);
   U22877 : XOR2_X1 port map( A1 => n11233, A2 => n22291, Z => n22506);
   U22879 : XOR2_X1 port map( A1 => n11236, A2 => n27479, Z => n11235);
   U22882 : NAND2_X1 port map( A1 => n15299, A2 => n7577, ZN => n23249);
   U22883 : XOR2_X1 port map( A1 => n11255, A2 => n11254, Z => n11253);
   U22885 : OAI21_X2 port map( A1 => n26940, A2 => n26939, B => n26938, ZN => 
                           n27184);
   U22886 : OAI21_X1 port map( A1 => n13971, A2 => n7317, B => n11257, ZN => 
                           n25955);
   U22887 : XOR2_X1 port map( A1 => n518, A2 => n1051, Z => n20592);
   U22888 : XOR2_X1 port map( A1 => n1558, A2 => n13531, Z => n13530);
   U22889 : NOR2_X1 port map( A1 => n15049, A2 => n1275, ZN => n11261);
   U22891 : NAND2_X1 port map( A1 => n14492, A2 => n11274, ZN => n16165);
   U22892 : XOR2_X1 port map( A1 => Plaintext(95), A2 => Key(95), Z => n15354);
   U22898 : XOR2_X1 port map( A1 => n22688, A2 => n11289, Z => n11288);
   U22899 : XOR2_X1 port map( A1 => n22544, A2 => n22409, Z => n11290);
   U22901 : INV_X1 port map( I => Plaintext(160), ZN => n11291);
   U22902 : XOR2_X1 port map( A1 => n11291, A2 => Key(160), Z => n12036);
   U22905 : XOR2_X1 port map( A1 => n22524, A2 => n22523, Z => n22857);
   U22907 : AOI21_X2 port map( A1 => n21636, A2 => n11303, B => n11302, ZN => 
                           n11304);
   U22909 : XOR2_X1 port map( A1 => n11311, A2 => n11310, Z => n11309);
   U22910 : XOR2_X1 port map( A1 => n22621, A2 => n19953, Z => n11310);
   U22912 : XOR2_X1 port map( A1 => n11314, A2 => n11313, Z => n11312);
   U22913 : XOR2_X1 port map( A1 => n9116, A2 => n19221, Z => n11313);
   U22915 : XOR2_X1 port map( A1 => n14304, A2 => n1745, Z => n21201);
   U22916 : INV_X2 port map( I => n15051, ZN => n25543);
   U22918 : XOR2_X1 port map( A1 => n11321, A2 => n25218, Z => n25219);
   U22924 : OAI22_X2 port map( A1 => n24689, A2 => n24690, B1 => n10019, B2 => 
                           n13002, ZN => n25237);
   U22926 : NAND2_X1 port map( A1 => n1314, A2 => n33745, ZN => n15081);
   U22929 : XOR2_X1 port map( A1 => n24994, A2 => n25127, Z => n25171);
   U22933 : XOR2_X1 port map( A1 => n15270, A2 => n5755, Z => n11346);
   U22936 : XOR2_X1 port map( A1 => n22606, A2 => n11356, Z => n11355);
   U22937 : XOR2_X1 port map( A1 => n22699, A2 => n11308, Z => n11356);
   U22941 : XOR2_X1 port map( A1 => n33027, A2 => n26554, Z => n26307);
   U22942 : XOR2_X1 port map( A1 => n33027, A2 => n19464, Z => n20539);
   U22943 : XOR2_X1 port map( A1 => n38937, A2 => n1374, Z => n11365);
   U22950 : XOR2_X1 port map( A1 => n11377, A2 => n11376, Z => n23122);
   U22951 : XOR2_X1 port map( A1 => n16278, A2 => n22646, Z => n11376);
   U22952 : XOR2_X1 port map( A1 => n22643, A2 => n22644, Z => n16278);
   U22958 : XOR2_X1 port map( A1 => n20294, A2 => n22636, Z => n11382);
   U22960 : XOR2_X1 port map( A1 => n11384, A2 => n28814, Z => n11783);
   U22961 : INV_X1 port map( I => n37295, ZN => n28769);
   U22964 : XOR2_X1 port map( A1 => n27773, A2 => n31295, Z => n11391);
   U22965 : XOR2_X1 port map( A1 => n27774, A2 => n36384, Z => n11392);
   U22969 : NAND2_X1 port map( A1 => n19090, A2 => n19085, ZN => n11397);
   U22974 : XOR2_X1 port map( A1 => n14843, A2 => n11405, Z => n11406);
   U22975 : NAND2_X1 port map( A1 => n11406, A2 => n12049, ZN => n15293);
   U22978 : XOR2_X1 port map( A1 => n11419, A2 => n11417, Z => n11416);
   U22979 : XOR2_X1 port map( A1 => n30964, A2 => n11418, Z => n11417);
   U22980 : INV_X1 port map( I => n28851, ZN => n11418);
   U22981 : XOR2_X1 port map( A1 => n13639, A2 => n15745, Z => n11419);
   U22987 : XOR2_X1 port map( A1 => n11425, A2 => n29974, Z => n17760);
   U22988 : XOR2_X1 port map( A1 => n4622, A2 => n11425, Z => n12587);
   U22989 : XOR2_X1 port map( A1 => n35065, A2 => n23880, Z => n23737);
   U22990 : XOR2_X1 port map( A1 => n22416, A2 => n1657, Z => n12205);
   U22995 : NAND2_X2 port map( A1 => n30128, A2 => n20274, ZN => n30127);
   U23001 : XOR2_X1 port map( A1 => n27539, A2 => n27029, Z => n11458);
   U23002 : INV_X2 port map( I => n11459, ZN => n12257);
   U23005 : INV_X1 port map( I => n23926, ZN => n11464);
   U23006 : NAND2_X1 port map( A1 => n26829, A2 => n11467, ZN => n21182);
   U23007 : NAND3_X2 port map( A1 => n11473, A2 => n23180, A3 => n11472, ZN => 
                           n23631);
   U23010 : XOR2_X1 port map( A1 => n25194, A2 => n1706, Z => n11475);
   U23011 : NAND2_X2 port map( A1 => n18393, A2 => n18394, ZN => n25194);
   U23012 : NAND2_X1 port map( A1 => n11476, A2 => n22722, ZN => n22730);
   U23013 : NAND2_X1 port map( A1 => n37954, A2 => n24328, ZN => n11477);
   U23018 : INV_X2 port map( I => n11482, ZN => n17240);
   U23020 : NOR2_X1 port map( A1 => n24206, A2 => n37264, ZN => n11494);
   U23025 : INV_X2 port map( I => n18502, ZN => n11506);
   U23030 : XOR2_X1 port map( A1 => n11519, A2 => n11520, Z => n13018);
   U23032 : XOR2_X1 port map( A1 => n25162, A2 => n24945, Z => n11520);
   U23034 : NOR2_X1 port map( A1 => n26666, A2 => n924, ZN => n11523);
   U23041 : NAND3_X1 port map( A1 => n31523, A2 => n39729, A3 => n33237, ZN => 
                           n26094);
   U23042 : NAND2_X1 port map( A1 => n17008, A2 => n11533, ZN => n20833);
   U23052 : XOR2_X1 port map( A1 => n1258, A2 => n11554, Z => n11553);
   U23053 : NAND2_X1 port map( A1 => n11556, A2 => n11555, ZN => n11554);
   U23054 : OAI21_X1 port map( A1 => n24495, A2 => n24496, B => n19128, ZN => 
                           n11555);
   U23055 : NAND2_X1 port map( A1 => n11558, A2 => n11557, ZN => n11556);
   U23056 : NOR2_X1 port map( A1 => n24496, A2 => n19128, ZN => n11557);
   U23057 : INV_X1 port map( I => n24495, ZN => n11558);
   U23058 : XOR2_X1 port map( A1 => n38213, A2 => n13054, Z => n11559);
   U23061 : INV_X1 port map( I => n20840, ZN => n23175);
   U23063 : XOR2_X1 port map( A1 => n19072, A2 => n11572, Z => n11571);
   U23064 : XOR2_X1 port map( A1 => n25242, A2 => n25241, Z => n11572);
   U23067 : XOR2_X1 port map( A1 => n13439, A2 => n17423, Z => n23953);
   U23068 : XOR2_X1 port map( A1 => n27607, A2 => n27707, Z => n27608);
   U23070 : NAND2_X1 port map( A1 => n5892, A2 => n35994, ZN => n23036);
   U23071 : INV_X2 port map( I => n11586, ZN => n14379);
   U23073 : AND2_X1 port map( A1 => n29237, A2 => n12141, Z => n14529);
   U23076 : XOR2_X1 port map( A1 => n14425, A2 => n11603, Z => n11602);
   U23079 : XOR2_X1 port map( A1 => n11612, A2 => n11611, Z => n12103);
   U23080 : XOR2_X1 port map( A1 => n2281, A2 => n27534, Z => n11611);
   U23082 : XOR2_X1 port map( A1 => n19608, A2 => n39559, Z => n11615);
   U23084 : XOR2_X1 port map( A1 => n12824, A2 => n26350, Z => n11621);
   U23086 : INV_X2 port map( I => n11622, ZN => n14436);
   U23090 : INV_X2 port map( I => n11627, ZN => n15163);
   U23091 : INV_X4 port map( I => n13609, ZN => n11628);
   U23092 : INV_X2 port map( I => n13787, ZN => n13609);
   U23097 : NAND2_X1 port map( A1 => n20092, A2 => n27438, ZN => n11637);
   U23099 : XOR2_X1 port map( A1 => n10213, A2 => n11644, Z => n22662);
   U23100 : XOR2_X1 port map( A1 => n11644, A2 => n1375, Z => n14609);
   U23101 : XOR2_X1 port map( A1 => n15448, A2 => n11644, Z => n20350);
   U23105 : INV_X2 port map( I => n11663, ZN => n15320);
   U23108 : NAND2_X1 port map( A1 => n5657, A2 => n22889, ZN => n23509);
   U23114 : XOR2_X1 port map( A1 => n30068, A2 => n24932, Z => n11688);
   U23115 : XOR2_X1 port map( A1 => n25133, A2 => n37296, Z => n11689);
   U23120 : XOR2_X1 port map( A1 => n11694, A2 => n29269, Z => n27477);
   U23121 : XOR2_X1 port map( A1 => n27669, A2 => n282, Z => n18548);
   U23123 : XOR2_X1 port map( A1 => n3703, A2 => n3665, Z => n28662);
   U23124 : XOR2_X1 port map( A1 => n11698, A2 => n30170, Z => n17134);
   U23125 : XOR2_X1 port map( A1 => n12534, A2 => n11698, Z => n25295);
   U23126 : XOR2_X1 port map( A1 => n24978, A2 => n11698, Z => n19073);
   U23127 : INV_X2 port map( I => n11699, ZN => n20517);
   U23129 : NOR2_X1 port map( A1 => n22901, A2 => n11704, ZN => n22468);
   U23133 : AND2_X1 port map( A1 => n15540, A2 => n31418, Z => n11718);
   U23136 : XOR2_X1 port map( A1 => n23663, A2 => n15094, Z => n11725);
   U23137 : OAI21_X1 port map( A1 => n26954, A2 => n26957, B => n11726, ZN => 
                           n13097);
   U23142 : NAND3_X1 port map( A1 => n30621, A2 => n425, A3 => n11734, ZN => 
                           n25404);
   U23143 : INV_X1 port map( I => n26521, ZN => n26347);
   U23147 : OAI21_X2 port map( A1 => n14503, A2 => n17125, B => n26218, ZN => 
                           n26407);
   U23149 : XOR2_X1 port map( A1 => n29036, A2 => n29035, Z => n11746);
   U23150 : XOR2_X1 port map( A1 => n11750, A2 => n11748, Z => n16593);
   U23151 : XOR2_X1 port map( A1 => n5463, A2 => n11749, Z => n11748);
   U23152 : XOR2_X1 port map( A1 => n22531, A2 => n11974, Z => n11749);
   U23154 : XOR2_X1 port map( A1 => n37951, A2 => n31591, Z => n16695);
   U23156 : XOR2_X1 port map( A1 => n11756, A2 => n25278, Z => n25279);
   U23157 : XOR2_X1 port map( A1 => n39541, A2 => n11756, Z => n11905);
   U23161 : NAND2_X2 port map( A1 => n25573, A2 => n25572, ZN => n26116);
   U23164 : XOR2_X1 port map( A1 => n22533, A2 => n22462, Z => n11779);
   U23166 : NOR2_X2 port map( A1 => n21103, A2 => n21104, ZN => n22582);
   U23167 : OAI21_X2 port map( A1 => n22010, A2 => n21105, B => n14683, ZN => 
                           n18778);
   U23168 : INV_X2 port map( I => n11780, ZN => n12931);
   U23170 : OR2_X1 port map( A1 => n11783, A2 => n20522, Z => n29010);
   U23172 : XOR2_X1 port map( A1 => n11790, A2 => n11788, Z => n21187);
   U23173 : XOR2_X1 port map( A1 => n28979, A2 => n11789, Z => n11788);
   U23174 : XOR2_X1 port map( A1 => n36905, A2 => n19932, Z => n11789);
   U23175 : XOR2_X1 port map( A1 => n28984, A2 => n19600, Z => n11790);
   U23177 : XOR2_X1 port map( A1 => n22717, A2 => n22514, Z => n11791);
   U23180 : XOR2_X1 port map( A1 => n22515, A2 => n1371, Z => n11793);
   U23185 : NOR2_X1 port map( A1 => n18029, A2 => n25614, ZN => n12096);
   U23186 : INV_X4 port map( I => n39827, ZN => n29185);
   U23188 : AND2_X1 port map( A1 => n7693, A2 => n19868, Z => n20690);
   U23192 : NAND3_X1 port map( A1 => n22212, A2 => n22213, A3 => n22361, ZN => 
                           n11921);
   U23195 : XOR2_X1 port map( A1 => n963, A2 => n29983, Z => n16061);
   U23196 : XOR2_X1 port map( A1 => n963, A2 => n19730, Z => n22720);
   U23198 : XOR2_X1 port map( A1 => n24023, A2 => n29875, Z => n23806);
   U23202 : XOR2_X1 port map( A1 => n22595, A2 => n37042, Z => n11809);
   U23206 : XOR2_X1 port map( A1 => n31181, A2 => n29785, Z => n12180);
   U23207 : XOR2_X1 port map( A1 => n31181, A2 => n30010, Z => n19074);
   U23208 : XOR2_X1 port map( A1 => n35972, A2 => n19845, Z => n24950);
   U23211 : XOR2_X1 port map( A1 => n507, A2 => n14969, Z => n24588);
   U23216 : XOR2_X1 port map( A1 => n6559, A2 => n13617, Z => n19984);
   U23217 : XOR2_X1 port map( A1 => n16639, A2 => n32836, Z => n14487);
   U23219 : NAND2_X2 port map( A1 => n13913, A2 => n14658, ZN => n23515);
   U23224 : AOI21_X2 port map( A1 => n21653, A2 => n11850, B => n11849, ZN => 
                           n19737);
   U23230 : INV_X2 port map( I => n13499, ZN => n28141);
   U23232 : XOR2_X1 port map( A1 => n27474, A2 => n15068, Z => n11871);
   U23238 : XOR2_X1 port map( A1 => n1410, A2 => n15780, Z => n11883);
   U23242 : OAI21_X1 port map( A1 => n11890, A2 => n28123, B => n11891, ZN => 
                           n11895);
   U23245 : INV_X1 port map( I => Plaintext(169), ZN => n11901);
   U23251 : NAND2_X1 port map( A1 => n13512, A2 => n36877, ZN => n14766);
   U23254 : XOR2_X1 port map( A1 => n16566, A2 => n11926, Z => n11925);
   U23255 : XOR2_X1 port map( A1 => n35202, A2 => n19874, Z => n11926);
   U23258 : XOR2_X1 port map( A1 => n18051, A2 => n35200, Z => n14285);
   U23262 : XOR2_X1 port map( A1 => n11962, A2 => n11961, Z => n11960);
   U23263 : XOR2_X1 port map( A1 => n33038, A2 => n19770, Z => n11961);
   U23264 : XOR2_X1 port map( A1 => n25071, A2 => n10273, Z => n11962);
   U23265 : NAND2_X2 port map( A1 => n20697, A2 => n11963, ZN => n25071);
   U23266 : XOR2_X1 port map( A1 => n14258, A2 => n11965, Z => n12612);
   U23267 : XOR2_X1 port map( A1 => n11966, A2 => n23795, Z => n11965);
   U23268 : XOR2_X1 port map( A1 => n36842, A2 => n29394, Z => n11966);
   U23271 : INV_X2 port map( I => n11975, ZN => n13770);
   U23273 : XOR2_X1 port map( A1 => n27788, A2 => n11977, Z => n11976);
   U23274 : XOR2_X1 port map( A1 => n17884, A2 => n21226, Z => n11977);
   U23281 : XOR2_X1 port map( A1 => n22677, A2 => n22715, Z => n11984);
   U23282 : XOR2_X1 port map( A1 => n20980, A2 => n22675, Z => n11985);
   U23283 : NAND2_X1 port map( A1 => n11987, A2 => n11986, ZN => n14140);
   U23284 : NAND3_X1 port map( A1 => n36701, A2 => n36011, A3 => n1695, ZN => 
                           n11986);
   U23287 : XOR2_X1 port map( A1 => n38641, A2 => n25090, Z => n11989);
   U23291 : XOR2_X1 port map( A1 => n27564, A2 => n27640, Z => n11994);
   U23292 : XOR2_X1 port map( A1 => n26221, A2 => n26143, Z => n11998);
   U23293 : XOR2_X1 port map( A1 => n26454, A2 => n26413, Z => n11999);
   U23294 : XOR2_X1 port map( A1 => n12000, A2 => n18869, Z => n12001);
   U23295 : NAND2_X1 port map( A1 => n2771, A2 => n37984, ZN => n22826);
   U23302 : NAND2_X2 port map( A1 => n12025, A2 => n12024, ZN => n19773);
   U23306 : XOR2_X1 port map( A1 => n13430, A2 => n639, Z => n23196);
   U23307 : AOI22_X2 port map( A1 => n25819, A2 => n25940, B1 => n25817, B2 => 
                           n25818, ZN => n20600);
   U23310 : INV_X2 port map( I => n12036, ZN => n21770);
   U23313 : XOR2_X1 port map( A1 => n18924, A2 => n35178, Z => n15222);
   U23318 : NAND2_X2 port map( A1 => n8127, A2 => n24668, ZN => n18858);
   U23321 : XOR2_X1 port map( A1 => n26160, A2 => n31605, Z => n12053);
   U23330 : XOR2_X1 port map( A1 => n25170, A2 => n24958, Z => n12076);
   U23331 : INV_X1 port map( I => n21213, ZN => n23638);
   U23333 : NAND2_X2 port map( A1 => n1424, A2 => n496, ZN => n28544);
   U23336 : INV_X1 port map( I => n24162, ZN => n24173);
   U23337 : XOR2_X1 port map( A1 => n12086, A2 => n12085, Z => n12084);
   U23338 : XOR2_X1 port map( A1 => n33323, A2 => n19845, Z => n12085);
   U23339 : XOR2_X1 port map( A1 => n22668, A2 => n7432, Z => n12086);
   U23344 : XOR2_X1 port map( A1 => n23778, A2 => n19910, Z => n12107);
   U23345 : XOR2_X1 port map( A1 => Plaintext(82), A2 => Key(82), Z => n12670);
   U23346 : NAND2_X1 port map( A1 => n9916, A2 => n25813, ZN => n13678);
   U23349 : XOR2_X1 port map( A1 => n12113, A2 => n12112, Z => n12111);
   U23350 : XOR2_X1 port map( A1 => n26455, A2 => n31771, Z => n12112);
   U23351 : NAND3_X2 port map( A1 => n26095, A2 => n26096, A3 => n26094, ZN => 
                           n26455);
   U23352 : XOR2_X1 port map( A1 => n26403, A2 => n26541, Z => n12113);
   U23353 : NAND2_X2 port map( A1 => n12490, A2 => n12489, ZN => n26541);
   U23356 : NOR2_X1 port map( A1 => n26185, A2 => n38185, ZN => n12115);
   U23359 : OAI21_X1 port map( A1 => n15456, A2 => n18152, B => n21840, ZN => 
                           n12118);
   U23360 : NAND2_X1 port map( A1 => n23111, A2 => n20783, ZN => n12123);
   U23362 : XOR2_X1 port map( A1 => n10329, A2 => n731, Z => n12132);
   U23363 : NAND2_X1 port map( A1 => n9913, A2 => n7303, ZN => n12547);
   U23364 : OAI22_X1 port map( A1 => n29462, A2 => n7303, B1 => n29464, B2 => 
                           n969, ZN => n13431);
   U23369 : XOR2_X1 port map( A1 => n7148, A2 => n19722, Z => n12139);
   U23370 : NAND3_X1 port map( A1 => n1388, A2 => n35185, A3 => n29236, ZN => 
                           n29233);
   U23371 : NOR2_X1 port map( A1 => n1388, A2 => n35185, ZN => n15028);
   U23373 : NAND3_X2 port map( A1 => n25950, A2 => n25949, A3 => n12151, ZN => 
                           n26438);
   U23375 : OAI22_X2 port map( A1 => n20996, A2 => n133, B1 => n22047, B2 => 
                           n21973, ZN => n22188);
   U23382 : XOR2_X1 port map( A1 => n557, A2 => n19890, Z => n12165);
   U23385 : XOR2_X1 port map( A1 => n35065, A2 => n1165, Z => n23674);
   U23390 : XOR2_X1 port map( A1 => n23745, A2 => n12184, Z => n12183);
   U23391 : XOR2_X1 port map( A1 => n23789, A2 => n35235, Z => n12184);
   U23392 : XOR2_X1 port map( A1 => n12185, A2 => n20093, Z => n28250);
   U23393 : XOR2_X1 port map( A1 => n379, A2 => n37242, Z => n12185);
   U23400 : XOR2_X1 port map( A1 => n22750, A2 => n12197, Z => n12196);
   U23401 : XOR2_X1 port map( A1 => n35824, A2 => n29506, Z => n12197);
   U23402 : NAND2_X1 port map( A1 => n30106, A2 => n18829, ZN => n12204);
   U23405 : INV_X2 port map( I => n18188, ZN => n19435);
   U23406 : INV_X2 port map( I => n15774, ZN => n19667);
   U23412 : INV_X2 port map( I => n12225, ZN => n18412);
   U23413 : XOR2_X1 port map( A1 => n22695, A2 => n36362, Z => n20048);
   U23415 : XOR2_X1 port map( A1 => n30865, A2 => n12233, Z => n24525);
   U23417 : XOR2_X1 port map( A1 => Plaintext(176), A2 => Key(176), Z => n12535
                           );
   U23418 : XOR2_X1 port map( A1 => n15286, A2 => n27843, Z => n12432);
   U23420 : XOR2_X1 port map( A1 => n12243, A2 => n19876, Z => n22545);
   U23422 : XOR2_X1 port map( A1 => n19516, A2 => n39536, Z => n28493);
   U23429 : XOR2_X1 port map( A1 => n24043, A2 => n23892, Z => n12265);
   U23430 : XOR2_X1 port map( A1 => n21316, A2 => n23656, Z => n12266);
   U23431 : INV_X2 port map( I => n12759, ZN => n24232);
   U23432 : XOR2_X1 port map( A1 => n12267, A2 => n30122, Z => n21225);
   U23433 : XOR2_X1 port map( A1 => n21227, A2 => n12973, Z => n18582);
   U23434 : NOR2_X1 port map( A1 => n16224, A2 => n29935, ZN => n12273);
   U23441 : NOR2_X1 port map( A1 => n23226, A2 => n12289, ZN => n16394);
   U23442 : NAND2_X1 port map( A1 => n23226, A2 => n12289, ZN => n15075);
   U23444 : NOR2_X1 port map( A1 => n31331, A2 => n12289, ZN => n23278);
   U23452 : XOR2_X1 port map( A1 => n17884, A2 => n29442, Z => n15726);
   U23453 : XOR2_X1 port map( A1 => n12970, A2 => n17884, Z => n12969);
   U23454 : INV_X2 port map( I => n12302, ZN => n20739);
   U23457 : NOR2_X1 port map( A1 => n12306, A2 => n27233, ZN => n27234);
   U23460 : XOR2_X1 port map( A1 => n25089, A2 => n25088, Z => n12310);
   U23464 : XOR2_X1 port map( A1 => n12316, A2 => n1377, Z => Ciphertext(47));
   U23465 : AOI21_X1 port map( A1 => n15841, A2 => n12318, B => n11506, ZN => 
                           n12317);
   U23466 : NAND2_X1 port map( A1 => n29439, A2 => n29438, ZN => n12318);
   U23472 : INV_X2 port map( I => n12334, ZN => n14399);
   U23475 : XOR2_X1 port map( A1 => n6522, A2 => n12337, Z => n12834);
   U23476 : XOR2_X1 port map( A1 => n9576, A2 => n33184, Z => n12337);
   U23480 : INV_X1 port map( I => n17777, ZN => n20632);
   U23482 : XOR2_X1 port map( A1 => n35218, A2 => n4709, Z => n12351);
   U23483 : INV_X2 port map( I => n14405, ZN => n15651);
   U23484 : XOR2_X1 port map( A1 => n28969, A2 => n12355, Z => n12354);
   U23485 : XOR2_X1 port map( A1 => n28850, A2 => n19950, Z => n12355);
   U23489 : NAND2_X1 port map( A1 => n24403, A2 => n20517, ZN => n12367);
   U23492 : INV_X2 port map( I => n17198, ZN => n19147);
   U23496 : XOR2_X1 port map( A1 => n27792, A2 => n27511, Z => n27569);
   U23502 : INV_X2 port map( I => n12403, ZN => n21898);
   U23503 : XNOR2_X1 port map( A1 => Plaintext(13), A2 => Key(13), ZN => n12403
                           );
   U23504 : NOR2_X1 port map( A1 => n13142, A2 => n3462, ZN => n13141);
   U23506 : INV_X2 port map( I => n12414, ZN => n29241);
   U23507 : XOR2_X1 port map( A1 => n12556, A2 => n1169, Z => n27000);
   U23509 : XOR2_X1 port map( A1 => n29260, A2 => n19804, Z => n13287);
   U23511 : XOR2_X1 port map( A1 => n25263, A2 => n19897, Z => n12438);
   U23515 : XOR2_X1 port map( A1 => n35188, A2 => n29522, Z => n27618);
   U23518 : NAND3_X1 port map( A1 => n14433, A2 => n20901, A3 => n12450, ZN => 
                           n14850);
   U23520 : XOR2_X1 port map( A1 => n12454, A2 => n28549, Z => n12453);
   U23521 : XOR2_X1 port map( A1 => n35262, A2 => n38160, Z => n12454);
   U23526 : XOR2_X1 port map( A1 => n12470, A2 => n12468, Z => n14076);
   U23527 : XOR2_X1 port map( A1 => n28589, A2 => n12469, Z => n12468);
   U23528 : XOR2_X1 port map( A1 => n19513, A2 => n28889, Z => n28589);
   U23530 : XOR2_X1 port map( A1 => n29092, A2 => n19751, Z => n12469);
   U23531 : XOR2_X1 port map( A1 => n14388, A2 => n29114, Z => n12470);
   U23532 : XOR2_X1 port map( A1 => n28865, A2 => n31396, Z => n29114);
   U23533 : NAND2_X2 port map( A1 => n19482, A2 => n28488, ZN => n29115);
   U23542 : XOR2_X1 port map( A1 => n12493, A2 => n12492, Z => n12491);
   U23543 : XOR2_X1 port map( A1 => n27631, A2 => n19681, Z => n12492);
   U23544 : XOR2_X1 port map( A1 => n27541, A2 => n20976, Z => n12493);
   U23545 : NOR2_X1 port map( A1 => n28271, A2 => n11628, ZN => n12498);
   U23546 : NAND3_X1 port map( A1 => n19290, A2 => n28271, A3 => n28272, ZN => 
                           n12499);
   U23551 : NOR2_X1 port map( A1 => n24603, A2 => n36058, ZN => n18055);
   U23552 : XOR2_X1 port map( A1 => n27302, A2 => n12507, Z => n18847);
   U23553 : XOR2_X1 port map( A1 => n23695, A2 => n14289, Z => n23786);
   U23557 : XOR2_X1 port map( A1 => n12516, A2 => n14309, Z => n12515);
   U23558 : INV_X2 port map( I => n18933, ZN => n19332);
   U23563 : NAND2_X1 port map( A1 => n25957, A2 => n18406, ZN => n12525);
   U23564 : INV_X2 port map( I => n12535, ZN => n13997);
   U23565 : XOR2_X1 port map( A1 => n29252, A2 => n29253, Z => n14171);
   U23568 : XOR2_X1 port map( A1 => n37101, A2 => n19894, Z => n27193);
   U23570 : XOR2_X1 port map( A1 => n18160, A2 => n29528, Z => n12553);
   U23574 : NOR2_X1 port map( A1 => n32580, A2 => n5519, ZN => n12558);
   U23579 : XOR2_X1 port map( A1 => n12562, A2 => n12561, Z => n12560);
   U23580 : XOR2_X1 port map( A1 => n28866, A2 => n16685, Z => n12563);
   U23584 : XOR2_X1 port map( A1 => n29292, A2 => n12576, Z => n12575);
   U23585 : XOR2_X1 port map( A1 => n16356, A2 => n19741, Z => n29049);
   U23586 : XOR2_X1 port map( A1 => n4341, A2 => n29832, Z => n12576);
   U23588 : XOR2_X1 port map( A1 => n26286, A2 => n12587, Z => n12586);
   U23589 : XOR2_X1 port map( A1 => n11298, A2 => n18180, Z => n12588);
   U23593 : XOR2_X1 port map( A1 => n12593, A2 => n25034, Z => n12592);
   U23594 : XOR2_X1 port map( A1 => n37943, A2 => n25160, Z => n12593);
   U23596 : XOR2_X1 port map( A1 => n14214, A2 => n25033, Z => n12594);
   U23597 : NAND2_X1 port map( A1 => n37105, A2 => n24912, ZN => n13610);
   U23598 : NAND2_X1 port map( A1 => n36634, A2 => n32825, ZN => n12654);
   U23601 : XOR2_X1 port map( A1 => n18568, A2 => n22511, Z => n22435);
   U23605 : XOR2_X1 port map( A1 => n12622, A2 => n16381, Z => n16382);
   U23606 : INV_X2 port map( I => n17313, ZN => n28236);
   U23607 : INV_X2 port map( I => n20945, ZN => n29815);
   U23608 : NAND2_X1 port map( A1 => n21397, A2 => n19483, ZN => n13682);
   U23609 : NAND2_X1 port map( A1 => n19327, A2 => n12644, ZN => n28011);
   U23611 : XOR2_X1 port map( A1 => n26197, A2 => n12655, Z => n20501);
   U23612 : XOR2_X1 port map( A1 => n29562, A2 => n12839, Z => n12655);
   U23613 : XOR2_X1 port map( A1 => n5848, A2 => n29875, Z => n26314);
   U23614 : XOR2_X1 port map( A1 => n14307, A2 => n29298, Z => n29299);
   U23615 : XOR2_X1 port map( A1 => n33452, A2 => n19894, Z => n12664);
   U23617 : XOR2_X1 port map( A1 => n6131, A2 => n19649, Z => n26228);
   U23618 : XOR2_X1 port map( A1 => n6131, A2 => n36544, Z => n12728);
   U23622 : XOR2_X1 port map( A1 => n33041, A2 => n30085, Z => n28928);
   U23625 : XOR2_X1 port map( A1 => n16376, A2 => n26594, Z => n12683);
   U23626 : XOR2_X1 port map( A1 => Plaintext(159), A2 => Key(159), Z => n12722
                           );
   U23629 : OR2_X1 port map( A1 => n20852, A2 => n20851, Z => n12689);
   U23630 : XOR2_X1 port map( A1 => n12570, A2 => n16697, Z => n16696);
   U23631 : NOR2_X1 port map( A1 => n13849, A2 => n34010, ZN => n12703);
   U23633 : AOI21_X2 port map( A1 => n34459, A2 => n975, B => n12715, ZN => 
                           n28799);
   U23634 : XOR2_X1 port map( A1 => n18601, A2 => n1718, Z => n29324);
   U23635 : INV_X2 port map( I => n12722, ZN => n12754);
   U23636 : OAI21_X1 port map( A1 => n19601, A2 => n27882, B => n19467, ZN => 
                           n12723);
   U23639 : XOR2_X1 port map( A1 => n12728, A2 => n12727, Z => n13183);
   U23640 : XOR2_X1 port map( A1 => n5031, A2 => n1730, Z => n12727);
   U23642 : XOR2_X1 port map( A1 => n12730, A2 => n1697, Z => n12862);
   U23643 : XOR2_X1 port map( A1 => n12730, A2 => n22762, Z => n16690);
   U23644 : INV_X2 port map( I => n12732, ZN => n29591);
   U23645 : XOR2_X1 port map( A1 => n12903, A2 => n26281, Z => n12736);
   U23646 : XOR2_X1 port map( A1 => n12741, A2 => n1738, Z => n28826);
   U23657 : XOR2_X1 port map( A1 => n22757, A2 => n16061, Z => n12762);
   U23660 : NAND2_X1 port map( A1 => n15332, A2 => n3120, ZN => n15333);
   U23661 : OAI21_X1 port map( A1 => n33344, A2 => n24847, B => n3120, ZN => 
                           n24540);
   U23663 : XOR2_X1 port map( A1 => n27758, A2 => n30179, Z => n12769);
   U23664 : INV_X2 port map( I => n12770, ZN => n21132);
   U23672 : XOR2_X1 port map( A1 => n39025, A2 => n29649, Z => n12796);
   U23673 : OAI21_X2 port map( A1 => n39467, A2 => n19880, B => n24395, ZN => 
                           n12804);
   U23677 : AOI21_X2 port map( A1 => n25834, A2 => n39291, B => n25833, ZN => 
                           n26253);
   U23679 : MUX2_X1 port map( I0 => n19581, I1 => n31580, S => n12828, Z => 
                           n12826);
   U23682 : XOR2_X1 port map( A1 => n25003, A2 => n25004, Z => n12833);
   U23683 : XOR2_X1 port map( A1 => n12835, A2 => n12834, Z => n12836);
   U23684 : XOR2_X1 port map( A1 => n7055, A2 => n32174, Z => n22697);
   U23687 : XOR2_X1 port map( A1 => n12847, A2 => n1734, Z => Ciphertext(29));
   U23688 : NAND2_X1 port map( A1 => n20566, A2 => n29241, ZN => n29287);
   U23689 : XOR2_X1 port map( A1 => n20976, A2 => n900, Z => n12854);
   U23691 : XOR2_X1 port map( A1 => n14230, A2 => n666, Z => n12858);
   U23693 : XOR2_X1 port map( A1 => n18446, A2 => n12862, Z => n12861);
   U23695 : XOR2_X1 port map( A1 => n25285, A2 => n16843, Z => n12871);
   U23701 : NAND3_X1 port map( A1 => n12885, A2 => n28352, A3 => n28351, ZN => 
                           n28353);
   U23702 : NAND2_X1 port map( A1 => n28535, A2 => n28495, ZN => n12888);
   U23705 : XOR2_X1 port map( A1 => n20412, A2 => n12897, Z => n12899);
   U23706 : XOR2_X1 port map( A1 => n17195, A2 => n22580, Z => n12897);
   U23707 : XOR2_X1 port map( A1 => n12898, A2 => n12899, Z => n12900);
   U23711 : XOR2_X1 port map( A1 => n22511, A2 => n18296, Z => n12901);
   U23712 : XOR2_X1 port map( A1 => n12902, A2 => Plaintext(23), Z => n21441);
   U23713 : INV_X1 port map( I => Key(23), ZN => n12902);
   U23717 : XOR2_X1 port map( A1 => n39172, A2 => n12915, Z => n17946);
   U23718 : XOR2_X1 port map( A1 => n2782, A2 => n12939, Z => n12918);
   U23719 : XOR2_X1 port map( A1 => n14756, A2 => n17817, Z => n12919);
   U23720 : XOR2_X1 port map( A1 => n12922, A2 => n790, Z => n12920);
   U23722 : XOR2_X1 port map( A1 => n23912, A2 => n23667, Z => n12922);
   U23724 : XOR2_X1 port map( A1 => n24944, A2 => n24984, Z => n25029);
   U23725 : NAND2_X1 port map( A1 => n12926, A2 => n370, ZN => n24481);
   U23733 : NOR2_X1 port map( A1 => n9839, A2 => n29367, ZN => n19059);
   U23736 : NOR2_X1 port map( A1 => n35023, A2 => n28695, ZN => n17320);
   U23738 : NAND2_X1 port map( A1 => n12950, A2 => n12951, ZN => n24273);
   U23742 : OAI21_X2 port map( A1 => n17724, A2 => n16660, B => n16659, ZN => 
                           n17685);
   U23746 : XOR2_X1 port map( A1 => n23812, A2 => n23220, Z => n12976);
   U23750 : NAND2_X1 port map( A1 => n38953, A2 => n16250, ZN => n12984);
   U23751 : XOR2_X1 port map( A1 => n29045, A2 => n29730, Z => n12985);
   U23752 : XOR2_X1 port map( A1 => n29289, A2 => n12989, Z => n29290);
   U23754 : XOR2_X1 port map( A1 => n24932, A2 => n25006, Z => n25234);
   U23755 : OAI22_X2 port map( A1 => n24726, A2 => n24725, B1 => n24724, B2 => 
                           n9656, ZN => n25006);
   U23756 : NAND2_X2 port map( A1 => n24415, A2 => n24414, ZN => n24932);
   U23759 : NAND2_X1 port map( A1 => n30171, A2 => n17997, ZN => n13006);
   U23760 : XOR2_X1 port map( A1 => n22485, A2 => n19925, Z => n13255);
   U23761 : NOR2_X1 port map( A1 => n13300, A2 => n24515, ZN => n24292);
   U23764 : XNOR2_X1 port map( A1 => n25303, A2 => n18991, ZN => n25329);
   U23765 : XOR2_X1 port map( A1 => n25330, A2 => n25331, Z => n13013);
   U23766 : NAND2_X1 port map( A1 => n21892, A2 => n12670, ZN => n19376);
   U23767 : XOR2_X1 port map( A1 => n13024, A2 => n13022, Z => n14122);
   U23768 : XOR2_X1 port map( A1 => n23741, A2 => n13023, Z => n13022);
   U23769 : XOR2_X1 port map( A1 => n23972, A2 => n13025, Z => n13024);
   U23774 : INV_X1 port map( I => n20342, ZN => n30181);
   U23777 : NOR2_X1 port map( A1 => n35506, A2 => n13038, ZN => n19924);
   U23782 : XOR2_X1 port map( A1 => n13054, A2 => n30094, Z => n16161);
   U23784 : XOR2_X1 port map( A1 => n39063, A2 => n26365, Z => n26398);
   U23793 : INV_X2 port map( I => n13082, ZN => n17410);
   U23794 : XOR2_X1 port map( A1 => n27636, A2 => n27639, Z => n13083);
   U23806 : XOR2_X1 port map( A1 => n23831, A2 => n1726, Z => n13101);
   U23807 : AND2_X1 port map( A1 => n25826, A2 => n25825, Z => n13103);
   U23813 : INV_X2 port map( I => n13124, ZN => n15290);
   U23815 : INV_X2 port map( I => n13127, ZN => n14962);
   U23816 : NAND3_X1 port map( A1 => n25630, A2 => n13129, A3 => n911, ZN => 
                           n25369);
   U23820 : INV_X1 port map( I => n13132, ZN => n29906);
   U23821 : XOR2_X1 port map( A1 => n37943, A2 => n14374, Z => n25231);
   U23822 : XOR2_X1 port map( A1 => n35953, A2 => n14374, Z => n25091);
   U23824 : XOR2_X1 port map( A1 => n25193, A2 => n14374, Z => n17553);
   U23826 : XOR2_X1 port map( A1 => n18543, A2 => n18546, Z => n13138);
   U23827 : XOR2_X1 port map( A1 => n5021, A2 => n19720, Z => n16093);
   U23828 : XOR2_X1 port map( A1 => n29024, A2 => n13139, Z => n14835);
   U23829 : XOR2_X1 port map( A1 => n19887, A2 => n29824, Z => n13139);
   U23830 : XOR2_X1 port map( A1 => n13140, A2 => n16498, Z => Ciphertext(1));
   U23835 : NAND2_X1 port map( A1 => n13153, A2 => n37060, ZN => n13657);
   U23836 : NAND2_X1 port map( A1 => n13158, A2 => n13998, ZN => n13557);
   U23837 : NAND2_X1 port map( A1 => n13170, A2 => n31542, ZN => n14222);
   U23839 : XOR2_X1 port map( A1 => n22661, A2 => n22660, Z => n13172);
   U23841 : XOR2_X1 port map( A1 => n13716, A2 => n13183, Z => n26968);
   U23842 : XOR2_X1 port map( A1 => n13188, A2 => n15835, Z => n13187);
   U23843 : XOR2_X1 port map( A1 => n29040, A2 => n30964, Z => n13188);
   U23846 : XOR2_X1 port map( A1 => n24417, A2 => n25133, Z => n13190);
   U23848 : XOR2_X1 port map( A1 => n22710, A2 => n36513, Z => n13199);
   U23852 : NAND2_X1 port map( A1 => n29763, A2 => n13208, ZN => n28963);
   U23853 : AND2_X1 port map( A1 => n13207, A2 => n28961, Z => n13208);
   U23855 : NOR2_X1 port map( A1 => n7676, A2 => n7973, ZN => n13212);
   U23857 : XOR2_X1 port map( A1 => n18279, A2 => n30068, Z => n13215);
   U23862 : NOR2_X1 port map( A1 => n22368, A2 => n13995, ZN => n13226);
   U23864 : XOR2_X1 port map( A1 => n26274, A2 => n39172, Z => n13232);
   U23866 : XOR2_X1 port map( A1 => n29024, A2 => n29823, Z => n21079);
   U23869 : XOR2_X1 port map( A1 => n26389, A2 => n19755, Z => n13242);
   U23870 : XOR2_X1 port map( A1 => n26437, A2 => n26567, Z => n13243);
   U23871 : XOR2_X1 port map( A1 => n31599, A2 => n7944, Z => n13247);
   U23872 : OR2_X1 port map( A1 => n29673, A2 => n18042, Z => n18795);
   U23873 : INV_X2 port map( I => n19948, ZN => n29764);
   U23875 : XOR2_X1 port map( A1 => n13255, A2 => n7432, Z => n13254);
   U23878 : NAND2_X2 port map( A1 => n19268, A2 => n21967, ZN => n22621);
   U23881 : XOR2_X1 port map( A1 => Plaintext(77), A2 => Key(77), Z => n17833);
   U23882 : NAND2_X2 port map( A1 => n29403, A2 => n29400, ZN => n29410);
   U23884 : XOR2_X1 port map( A1 => n33509, A2 => n29522, Z => n17243);
   U23887 : INV_X1 port map( I => n13278, ZN => n20708);
   U23888 : XOR2_X1 port map( A1 => n13283, A2 => n27658, Z => n27659);
   U23892 : INV_X2 port map( I => n13286, ZN => n13545);
   U23895 : INV_X1 port map( I => n13292, ZN => n13291);
   U23896 : XOR2_X1 port map( A1 => n22595, A2 => n28934, Z => n13295);
   U23897 : OR2_X1 port map( A1 => n29493, A2 => n15621, Z => n13302);
   U23898 : NOR2_X1 port map( A1 => n13959, A2 => n13997, ZN => n13556);
   U23903 : AOI21_X2 port map( A1 => n24278, A2 => n13310, B => n24277, ZN => 
                           n24515);
   U23904 : XOR2_X1 port map( A1 => n13315, A2 => n13312, Z => n13317);
   U23906 : XOR2_X1 port map( A1 => n9035, A2 => n19800, Z => n13313);
   U23908 : INV_X2 port map( I => n13317, ZN => n29493);
   U23909 : NOR3_X1 port map( A1 => n21397, A2 => n13318, A3 => n13997, ZN => 
                           n13684);
   U23910 : NOR2_X1 port map( A1 => n695, A2 => n18959, ZN => n13318);
   U23913 : XOR2_X1 port map( A1 => n25247, A2 => n20479, Z => n13326);
   U23917 : XOR2_X1 port map( A1 => n8894, A2 => n27735, Z => n27547);
   U23918 : XOR2_X1 port map( A1 => n13329, A2 => n19929, Z => Ciphertext(38));
   U23921 : INV_X2 port map( I => n13332, ZN => n28283);
   U23922 : XOR2_X1 port map( A1 => n31579, A2 => n19786, Z => n15405);
   U23924 : MUX2_X1 port map( I0 => n19737, I1 => n18656, S => n22228, Z => 
                           n22027);
   U23932 : XOR2_X1 port map( A1 => n22651, A2 => n22652, Z => n13356);
   U23934 : XOR2_X1 port map( A1 => n29123, A2 => n14244, Z => n13358);
   U23937 : XNOR2_X1 port map( A1 => Plaintext(54), A2 => Key(54), ZN => n13359
                           );
   U23939 : INV_X2 port map( I => n22837, ZN => n23101);
   U23940 : XOR2_X1 port map( A1 => n13362, A2 => n13361, Z => n22837);
   U23941 : XOR2_X1 port map( A1 => n17988, A2 => n14894, Z => n13361);
   U23942 : XOR2_X1 port map( A1 => n22774, A2 => n22662, Z => n13362);
   U23943 : XOR2_X1 port map( A1 => n23971, A2 => n13368, Z => n13367);
   U23944 : XOR2_X1 port map( A1 => n24049, A2 => n19937, Z => n13368);
   U23945 : XOR2_X1 port map( A1 => n26573, A2 => n29334, Z => n26575);
   U23946 : AND2_X1 port map( A1 => n28466, A2 => n13372, Z => n16840);
   U23953 : XOR2_X1 port map( A1 => n13544, A2 => n26294, Z => n13543);
   U23954 : INV_X2 port map( I => n13397, ZN => n21912);
   U23957 : XOR2_X1 port map( A1 => n16651, A2 => n33990, Z => n16650);
   U23959 : OAI21_X1 port map( A1 => n19007, A2 => n13412, B => n1032, ZN => 
                           n17301);
   U23960 : INV_X2 port map( I => n13413, ZN => n18909);
   U23961 : NAND2_X1 port map( A1 => n13415, A2 => n1121, ZN => n24413);
   U23964 : MUX2_X1 port map( I0 => n16853, I1 => n35224, S => n14193, Z => 
                           n13424);
   U23965 : INV_X1 port map( I => n26177, ZN => n26703);
   U23966 : INV_X2 port map( I => n13425, ZN => n19951);
   U23968 : INV_X2 port map( I => n13429, ZN => n17693);
   U23969 : XOR2_X1 port map( A1 => n14303, A2 => n22611, Z => n13430);
   U23970 : AOI21_X1 port map( A1 => n20964, A2 => n34534, B => n13433, ZN => 
                           n13432);
   U23971 : INV_X1 port map( I => n17594, ZN => n25575);
   U23972 : XOR2_X1 port map( A1 => n13439, A2 => n23880, Z => n23660);
   U23975 : XOR2_X1 port map( A1 => n27864, A2 => n29476, Z => n13448);
   U23976 : AND2_X1 port map( A1 => n1645, A2 => n19351, Z => n13451);
   U23977 : INV_X2 port map( I => n14332, ZN => n25539);
   U23978 : XOR2_X1 port map( A1 => Plaintext(69), A2 => Key(69), Z => n13473);
   U23979 : XOR2_X1 port map( A1 => n13477, A2 => n13475, Z => n21291);
   U23980 : XOR2_X1 port map( A1 => n13476, A2 => n22565, Z => n13475);
   U23981 : XOR2_X1 port map( A1 => n19254, A2 => n22732, Z => n13476);
   U23983 : XOR2_X1 port map( A1 => n13479, A2 => n11541, Z => n13478);
   U23984 : XOR2_X1 port map( A1 => n17605, A2 => n19720, Z => n13479);
   U23991 : XOR2_X1 port map( A1 => n31504, A2 => n29320, Z => n22200);
   U23997 : INV_X2 port map( I => n13503, ZN => n24445);
   U24000 : XOR2_X1 port map( A1 => n27782, A2 => n13510, Z => n13969);
   U24001 : XOR2_X1 port map( A1 => n27781, A2 => n19749, Z => n13510);
   U24003 : NAND2_X2 port map( A1 => n13523, A2 => n13525, ZN => n17757);
   U24008 : NAND3_X1 port map( A1 => n1340, A2 => n4200, A3 => n13519, ZN => 
                           n21334);
   U24013 : NOR2_X1 port map( A1 => n8304, A2 => n1551, ZN => n19302);
   U24014 : XOR2_X1 port map( A1 => n29104, A2 => n29306, Z => n28869);
   U24022 : AND2_X1 port map( A1 => n25717, A2 => n25716, Z => n13538);
   U24023 : MUX2_X1 port map( I0 => n28141, I1 => n20184, S => n281, Z => 
                           n13539);
   U24025 : XOR2_X1 port map( A1 => n23996, A2 => n38813, Z => n23684);
   U24031 : XOR2_X1 port map( A1 => n28574, A2 => n13552, Z => n13551);
   U24032 : XOR2_X1 port map( A1 => n29837, A2 => n19613, Z => n13552);
   U24036 : OAI21_X1 port map( A1 => n16472, A2 => n13559, B => n13558, ZN => 
                           n16469);
   U24037 : AOI22_X1 port map( A1 => n16471, A2 => n30093, B1 => n16470, B2 => 
                           n13559, ZN => n13558);
   U24039 : INV_X2 port map( I => n13561, ZN => n23020);
   U24042 : XOR2_X1 port map( A1 => n22659, A2 => n15909, Z => n20865);
   U24043 : INV_X1 port map( I => n22347, ZN => n13566);
   U24044 : XOR2_X1 port map( A1 => n13569, A2 => n19817, Z => n27513);
   U24053 : XOR2_X1 port map( A1 => n15216, A2 => n28912, Z => n17905);
   U24057 : XOR2_X1 port map( A1 => n13592, A2 => n22559, Z => n13591);
   U24058 : XOR2_X1 port map( A1 => n22773, A2 => n29661, Z => n13592);
   U24063 : INV_X2 port map( I => n13595, ZN => n28036);
   U24065 : XOR2_X1 port map( A1 => n23830, A2 => n18828, Z => n17581);
   U24076 : NAND2_X1 port map( A1 => n16065, A2 => n19855, ZN => n13623);
   U24080 : XOR2_X1 port map( A1 => n13634, A2 => n29399, Z => n24936);
   U24085 : XOR2_X1 port map( A1 => n23688, A2 => n23465, Z => n13649);
   U24087 : XOR2_X1 port map( A1 => n21332, A2 => Key(102), Z => n19387);
   U24089 : XOR2_X1 port map( A1 => n35824, A2 => n2383, Z => n22520);
   U24093 : XOR2_X1 port map( A1 => n13658, A2 => n19492, Z => n18135);
   U24095 : XOR2_X1 port map( A1 => n17565, A2 => n13667, Z => n13668);
   U24096 : INV_X2 port map( I => n13668, ZN => n14442);
   U24097 : NOR2_X1 port map( A1 => n19704, A2 => n33368, ZN => n13672);
   U24098 : XOR2_X1 port map( A1 => n17757, A2 => n12649, Z => n13674);
   U24100 : XOR2_X1 port map( A1 => Plaintext(72), A2 => Key(72), Z => n13679);
   U24101 : XOR2_X1 port map( A1 => n705, A2 => n5203, Z => n13680);
   U24102 : XOR2_X1 port map( A1 => n22700, A2 => n14022, Z => n13681);
   U24103 : NAND2_X2 port map( A1 => n13683, A2 => n13682, ZN => n22315);
   U24104 : XOR2_X1 port map( A1 => n25137, A2 => n13689, Z => n25138);
   U24105 : XOR2_X1 port map( A1 => n1258, A2 => n16864, Z => n13689);
   U24112 : NAND2_X1 port map( A1 => n26856, A2 => n11334, ZN => n13698);
   U24115 : NAND2_X1 port map( A1 => n1641, A2 => n35689, ZN => n23617);
   U24116 : XOR2_X1 port map( A1 => n386, A2 => n1718, Z => n16709);
   U24118 : XOR2_X1 port map( A1 => n35505, A2 => n16226, Z => n22664);
   U24121 : NOR2_X1 port map( A1 => n24309, A2 => n807, ZN => n13710);
   U24126 : XOR2_X1 port map( A1 => n26364, A2 => n26482, Z => n13716);
   U24128 : INV_X2 port map( I => n13725, ZN => n15153);
   U24129 : XOR2_X1 port map( A1 => n23756, A2 => n16244, Z => n13729);
   U24131 : INV_X2 port map( I => n16993, ZN => n21484);
   U24132 : XOR2_X1 port map( A1 => Plaintext(86), A2 => Key(86), Z => n16993);
   U24134 : INV_X2 port map( I => n13745, ZN => n23107);
   U24135 : XOR2_X1 port map( A1 => n13750, A2 => n27521, Z => n13749);
   U24136 : NAND2_X1 port map( A1 => n13786, A2 => n30262, ZN => n13990);
   U24137 : NOR2_X1 port map( A1 => n13753, A2 => n35114, ZN => n27331);
   U24139 : NOR2_X1 port map( A1 => n11039, A2 => n13753, ZN => n27332);
   U24141 : INV_X2 port map( I => n13759, ZN => n26839);
   U24148 : NAND2_X2 port map( A1 => n13789, A2 => n13788, ZN => n19515);
   U24151 : XOR2_X1 port map( A1 => n29245, A2 => n29244, Z => n13797);
   U24153 : NOR2_X1 port map( A1 => n26137, A2 => n13801, ZN => n15684);
   U24154 : XOR2_X1 port map( A1 => n13802, A2 => n19879, Z => n27087);
   U24155 : XOR2_X1 port map( A1 => n27679, A2 => n13802, Z => n27042);
   U24156 : INV_X2 port map( I => n13827, ZN => n19863);
   U24162 : AND2_X1 port map( A1 => n13834, A2 => n13833, Z => n13832);
   U24165 : XOR2_X1 port map( A1 => n22608, A2 => n13846, Z => n13845);
   U24167 : INV_X2 port map( I => n13862, ZN => n14404);
   U24175 : XOR2_X1 port map( A1 => n900, A2 => n19761, Z => n13878);
   U24176 : OAI21_X1 port map( A1 => n16778, A2 => n33843, B => n13879, ZN => 
                           n14931);
   U24179 : OR2_X1 port map( A1 => n37157, A2 => n19085, Z => n13886);
   U24182 : NOR2_X1 port map( A1 => n11413, A2 => n8944, ZN => n13892);
   U24185 : MUX2_X1 port map( I0 => n27876, I1 => n28200, S => n18061, Z => 
                           n13907);
   U24189 : XOR2_X1 port map( A1 => n20352, A2 => n9626, Z => n22533);
   U24197 : XOR2_X1 port map( A1 => n34178, A2 => n29300, Z => n13933);
   U24199 : XOR2_X1 port map( A1 => n21108, A2 => n29110, Z => n13934);
   U24200 : XOR2_X1 port map( A1 => n14639, A2 => n16417, Z => n13937);
   U24201 : XOR2_X1 port map( A1 => n25277, A2 => n33661, Z => n13939);
   U24203 : OAI21_X1 port map( A1 => n14409, A2 => n33925, B => n13945, ZN => 
                           n23206);
   U24209 : XOR2_X1 port map( A1 => n39765, A2 => n17646, Z => n13967);
   U24212 : NOR2_X1 port map( A1 => n28231, A2 => n18451, ZN => n13983);
   U24216 : INV_X2 port map( I => n14000, ZN => n19762);
   U24218 : NAND3_X1 port map( A1 => n14006, A2 => n22817, A3 => n6646, ZN => 
                           n22819);
   U24219 : OAI21_X1 port map( A1 => n29810, A2 => n966, B => n15189, ZN => 
                           n14008);
   U24221 : INV_X2 port map( I => n14016, ZN => n19395);
   U24222 : XNOR2_X1 port map( A1 => Plaintext(108), A2 => Key(108), ZN => 
                           n14016);
   U24225 : XOR2_X1 port map( A1 => n22515, A2 => n30120, Z => n14022);
   U24228 : XOR2_X1 port map( A1 => n20723, A2 => n18539, Z => n14031);
   U24230 : XOR2_X1 port map( A1 => n12839, A2 => n26476, Z => n14143);
   U24231 : NOR3_X1 port map( A1 => n2839, A2 => n14027, A3 => n36428, ZN => 
                           n14034);
   U24232 : NOR2_X1 port map( A1 => n17664, A2 => n2839, ZN => n14035);
   U24233 : XOR2_X1 port map( A1 => n25264, A2 => n719, Z => n14043);
   U24234 : XOR2_X1 port map( A1 => n17837, A2 => n24966, Z => n14046);
   U24237 : NAND2_X1 port map( A1 => n34074, A2 => n37377, ZN => n14050);
   U24241 : XOR2_X1 port map( A1 => n7942, A2 => n14063, Z => n14062);
   U24242 : XOR2_X1 port map( A1 => n22741, A2 => n31863, Z => n14063);
   U24244 : XOR2_X1 port map( A1 => n26590, A2 => n29689, Z => n14069);
   U24250 : XOR2_X1 port map( A1 => n14128, A2 => n31547, Z => n14099);
   U24252 : XOR2_X1 port map( A1 => n23676, A2 => n14105, Z => n14104);
   U24253 : XOR2_X1 port map( A1 => n23890, A2 => n19681, Z => n14105);
   U24256 : INV_X1 port map( I => n22603, ZN => n19118);
   U24258 : XOR2_X1 port map( A1 => n35824, A2 => n28831, Z => n14112);
   U24259 : XOR2_X1 port map( A1 => n22787, A2 => n22447, Z => n14113);
   U24270 : XOR2_X1 port map( A1 => n27567, A2 => n27568, Z => n14147);
   U24271 : XOR2_X1 port map( A1 => n33252, A2 => n30065, Z => n14148);
   U24273 : AOI21_X2 port map( A1 => n29496, A2 => n14151, B => n14150, ZN => 
                           n20208);
   U24275 : OR2_X1 port map( A1 => n37227, A2 => n17693, Z => n14154);
   U24279 : XOR2_X1 port map( A1 => n5208, A2 => n31543, Z => n24542);
   U24281 : XOR2_X1 port map( A1 => Plaintext(88), A2 => Key(88), Z => n21882);
   U24284 : XOR2_X1 port map( A1 => n22668, A2 => n22563, Z => n21994);
   U24286 : NAND2_X2 port map( A1 => n23800, A2 => n14169, ZN => n24821);
   U24287 : XOR2_X1 port map( A1 => n31566, A2 => n19851, Z => n14173);
   U24288 : INV_X1 port map( I => n28290, ZN => n28155);
   U24291 : XOR2_X1 port map( A1 => n9116, A2 => n33990, Z => n22698);
   U24296 : XOR2_X1 port map( A1 => n22647, A2 => n22772, Z => n14194);
   U24297 : NAND2_X2 port map( A1 => n20487, A2 => n27572, ZN => n15745);
   U24298 : AOI21_X1 port map( A1 => n17973, A2 => n17972, B => n14196, ZN => 
                           n20670);
   U24302 : XOR2_X1 port map( A1 => n37499, A2 => n38212, Z => n18579);
   U24303 : NAND2_X1 port map( A1 => n25971, A2 => n35151, ZN => n14215);
   U24305 : XOR2_X1 port map( A1 => n36218, A2 => n19755, Z => n24524);
   U24306 : XOR2_X1 port map( A1 => n36218, A2 => n24982, Z => n24861);
   U24307 : NAND2_X2 port map( A1 => n15038, A2 => n14426, ZN => n14232);
   U24310 : XOR2_X1 port map( A1 => n31522, A2 => n20658, Z => n14244);
   U24312 : XNOR2_X1 port map( A1 => Plaintext(49), A2 => Key(49), ZN => n14245
                           );
   U24316 : OAI21_X2 port map( A1 => n14252, A2 => n14251, B => n14248, ZN => 
                           n22594);
   U24321 : XNOR2_X1 port map( A1 => n24065, A2 => n23905, ZN => n16781);
   U24326 : NOR2_X1 port map( A1 => n19193, A2 => n17238, ZN => n14282);
   U24328 : XOR2_X1 port map( A1 => Key(127), A2 => Plaintext(127), Z => n19871
                           );
   U24329 : INV_X2 port map( I => n14287, ZN => n19594);
   U24331 : XOR2_X1 port map( A1 => n33252, A2 => n19904, Z => n14293);
   U24332 : XOR2_X1 port map( A1 => n22771, A2 => n14295, Z => n14294);
   U24333 : XOR2_X1 port map( A1 => n22528, A2 => n11308, Z => n14295);
   U24336 : XOR2_X1 port map( A1 => n26457, A2 => n837, Z => n14302);
   U24337 : XOR2_X1 port map( A1 => n14304, A2 => n14309, Z => n14303);
   U24339 : XOR2_X1 port map( A1 => n14307, A2 => n15203, Z => n16583);
   U24343 : XOR2_X1 port map( A1 => n33038, A2 => n29849, Z => n19131);
   U24350 : XOR2_X1 port map( A1 => n1458, A2 => n27556, Z => n27573);
   U24351 : XOR2_X1 port map( A1 => n27461, A2 => n14325, Z => n27462);
   U24354 : INV_X1 port map( I => Plaintext(71), ZN => n14333);
   U24357 : MUX2_X1 port map( I0 => n28006, I1 => n28007, S => n941, Z => 
                           n28010);
   U24358 : OAI22_X2 port map( A1 => n22878, A2 => n14343, B1 => n22877, B2 => 
                           n23121, ZN => n23461);
   U24365 : XOR2_X1 port map( A1 => n39637, A2 => n29647, Z => n26344);
   U24369 : XOR2_X1 port map( A1 => n18300, A2 => n23675, Z => n23741);
   U24370 : OAI21_X2 port map( A1 => n14363, A2 => n19292, B => n21803, ZN => 
                           n22773);
   U24371 : XOR2_X1 port map( A1 => n6435, A2 => n32174, Z => n14364);
   U24373 : NOR2_X1 port map( A1 => n25048, A2 => n24912, ZN => n15633);
   U24375 : AOI21_X1 port map( A1 => n23311, A2 => n39626, B => n19869, ZN => 
                           n23015);
   U24386 : NOR2_X1 port map( A1 => n28675, A2 => n28676, ZN => n15631);
   U24390 : NOR2_X1 port map( A1 => n14450, A2 => n1354, ZN => n17724);
   U24393 : NAND2_X1 port map( A1 => n19594, A2 => n20590, ZN => n19361);
   U24394 : INV_X1 port map( I => n27862, ZN => n20310);
   U24395 : NAND2_X1 port map( A1 => n17942, A2 => n17551, ZN => n16534);
   U24397 : NOR2_X1 port map( A1 => n11307, A2 => n20782, ZN => n23113);
   U24406 : NAND2_X1 port map( A1 => n16159, A2 => n10477, ZN => n16158);
   U24408 : NOR2_X1 port map( A1 => n24854, A2 => n24853, ZN => n18537);
   U24414 : NAND2_X1 port map( A1 => n36954, A2 => n20010, ZN => n19996);
   U24415 : NAND2_X1 port map( A1 => n5020, A2 => n28282, ZN => n28068);
   U24418 : NAND3_X1 port map( A1 => n31604, A2 => n21672, A3 => n21667, ZN => 
                           n14912);
   U24419 : NAND2_X1 port map( A1 => n18266, A2 => n694, ZN => n16763);
   U24423 : OAI21_X1 port map( A1 => n21551, A2 => n11851, B => n1690, ZN => 
                           n20330);
   U24430 : NAND2_X1 port map( A1 => n1678, A2 => n9685, ZN => n16455);
   U24433 : INV_X1 port map( I => n20518, ZN => n23063);
   U24436 : NAND2_X1 port map( A1 => n22928, A2 => n22990, ZN => n18377);
   U24444 : NOR2_X1 port map( A1 => n17076, A2 => n24461, ZN => n20002);
   U24447 : NAND3_X1 port map( A1 => n1634, A2 => n23552, A3 => n14845, ZN => 
                           n18915);
   U24448 : NAND2_X1 port map( A1 => n6849, A2 => n24469, ZN => n19053);
   U24451 : INV_X1 port map( I => n20394, ZN => n24156);
   U24459 : NAND2_X1 port map( A1 => n16999, A2 => n39317, ZN => n19643);
   U24460 : INV_X1 port map( I => n37943, ZN => n16350);
   U24462 : INV_X1 port map( I => n20627, ZN => n25390);
   U24463 : INV_X1 port map( I => n25724, ZN => n16317);
   U24464 : NAND2_X1 port map( A1 => n15180, A2 => n37926, ZN => n25399);
   U24469 : INV_X1 port map( I => n26163, ZN => n19464);
   U24474 : NAND2_X1 port map( A1 => n27321, A2 => n14881, ZN => n18251);
   U24477 : INV_X1 port map( I => n16169, ZN => n17051);
   U24478 : INV_X1 port map( I => n27606, ZN => n27609);
   U24479 : NAND2_X1 port map( A1 => n17686, A2 => n17699, ZN => n15162);
   U24480 : NAND3_X1 port map( A1 => n27449, A2 => n33893, A3 => n16043, ZN => 
                           n15277);
   U24481 : INV_X1 port map( I => n27507, ZN => n15246);
   U24482 : INV_X1 port map( I => n17349, ZN => n20721);
   U24484 : NAND2_X1 port map( A1 => n27989, A2 => n38996, ZN => n18687);
   U24489 : NAND2_X1 port map( A1 => n20053, A2 => n7591, ZN => n19324);
   U24490 : NAND2_X1 port map( A1 => n38874, A2 => n18948, ZN => n19325);
   U24493 : NAND2_X1 port map( A1 => n27984, A2 => n37204, ZN => n19957);
   U24494 : NAND2_X1 port map( A1 => n16777, A2 => n17542, ZN => n17541);
   U24495 : INV_X1 port map( I => n7667, ZN => n28931);
   U24498 : NAND2_X1 port map( A1 => n21550, A2 => n21506, ZN => n15149);
   U24500 : INV_X1 port map( I => n21753, ZN => n21698);
   U24502 : NOR3_X1 port map( A1 => n20535, A2 => n3562, A3 => n21870, ZN => 
                           n15155);
   U24506 : NOR2_X1 port map( A1 => n21862, A2 => n21823, ZN => n15097);
   U24507 : OR2_X1 port map( A1 => n19016, A2 => n21858, Z => n15099);
   U24508 : INV_X1 port map( I => n21841, ZN => n21903);
   U24517 : OAI21_X1 port map( A1 => n37200, A2 => n1349, B => n1990, ZN => 
                           n19320);
   U24520 : NAND2_X1 port map( A1 => n39680, A2 => n21488, ZN => n19377);
   U24521 : NAND2_X1 port map( A1 => n39680, A2 => n21568, ZN => n14919);
   U24522 : NOR2_X1 port map( A1 => n20799, A2 => n1333, ZN => n18728);
   U24523 : NAND2_X1 port map( A1 => n9942, A2 => n18152, ZN => n21843);
   U24524 : NAND2_X1 port map( A1 => n21890, A2 => n15910, ZN => n18758);
   U24525 : NOR2_X1 port map( A1 => n21784, A2 => n20241, ZN => n21505);
   U24527 : NOR2_X1 port map( A1 => n19850, A2 => n16333, ZN => n21694);
   U24529 : NOR2_X1 port map( A1 => n34282, A2 => n17989, ZN => n20280);
   U24530 : NAND2_X1 port map( A1 => n21593, A2 => n21484, ZN => n21590);
   U24534 : OAI21_X1 port map( A1 => n32525, A2 => n18028, B => n1354, ZN => 
                           n21935);
   U24535 : AOI21_X1 port map( A1 => n20003, A2 => n20476, B => n16537, ZN => 
                           n16536);
   U24539 : OAI21_X1 port map( A1 => n18412, A2 => n21917, B => n19105, ZN => 
                           n19104);
   U24541 : NAND2_X1 port map( A1 => n21917, A2 => n34867, ZN => n19105);
   U24544 : NOR2_X1 port map( A1 => n9543, A2 => n23042, ZN => n14851);
   U24553 : NOR2_X1 port map( A1 => n22865, A2 => n12331, ZN => n15239);
   U24554 : NOR2_X1 port map( A1 => n18071, A2 => n18072, ZN => n18506);
   U24555 : NAND2_X1 port map( A1 => n33933, A2 => n23076, ZN => n15039);
   U24558 : INV_X1 port map( I => n22934, ZN => n22083);
   U24559 : NAND2_X1 port map( A1 => n18850, A2 => n23308, ZN => n23309);
   U24568 : INV_X1 port map( I => n23420, ZN => n17224);
   U24572 : NAND2_X1 port map( A1 => n22992, A2 => n22993, ZN => n20024);
   U24573 : NAND2_X1 port map( A1 => n16292, A2 => n16291, ZN => n16150);
   U24574 : OAI21_X1 port map( A1 => n23346, A2 => n1634, B => n23550, ZN => 
                           n18618);
   U24575 : INV_X1 port map( I => n24077, ZN => n15477);
   U24578 : NAND2_X1 port map( A1 => n24311, A2 => n19584, ZN => n16918);
   U24579 : NAND3_X1 port map( A1 => n9078, A2 => n20972, A3 => n4542, ZN => 
                           n15534);
   U24582 : NAND2_X1 port map( A1 => n32069, A2 => n39074, ZN => n24153);
   U24583 : NAND2_X1 port map( A1 => n24795, A2 => n16238, ZN => n17453);
   U24585 : NOR2_X1 port map( A1 => n24419, A2 => n30494, ZN => n24090);
   U24592 : NAND2_X1 port map( A1 => n24660, A2 => n18110, ZN => n18263);
   U24593 : INV_X1 port map( I => n24784, ZN => n24785);
   U24596 : OAI21_X1 port map( A1 => n596, A2 => n26061, B => n9530, ZN => 
                           n25740);
   U24601 : NOR2_X1 port map( A1 => n26185, A2 => n25934, ZN => n26187);
   U24603 : INV_X1 port map( I => n26338, ZN => n26418);
   U24606 : NAND2_X1 port map( A1 => n9859, A2 => n25849, ZN => n14839);
   U24609 : NOR2_X1 port map( A1 => n25754, A2 => n25699, ZN => n21233);
   U24610 : NOR2_X1 port map( A1 => n24896, A2 => n25390, ZN => n17091);
   U24611 : INV_X1 port map( I => n25418, ZN => n25600);
   U24614 : NOR2_X1 port map( A1 => n36249, A2 => n19637, ZN => n16810);
   U24620 : NAND2_X1 port map( A1 => n26923, A2 => n13393, ZN => n17025);
   U24626 : INV_X1 port map( I => n18146, ZN => n18145);
   U24630 : NAND2_X1 port map( A1 => n26803, A2 => n26802, ZN => n20797);
   U24631 : NAND2_X1 port map( A1 => n20669, A2 => n26961, ZN => n17601);
   U24636 : OAI21_X1 port map( A1 => n26937, A2 => n875, B => n17993, ZN => 
                           n26856);
   U24638 : NOR2_X1 port map( A1 => n26734, A2 => n9188, ZN => n16924);
   U24639 : NAND2_X1 port map( A1 => n13758, A2 => n13757, ZN => n14861);
   U24641 : NAND2_X1 port map( A1 => n27347, A2 => n993, ZN => n18651);
   U24642 : INV_X1 port map( I => n18652, ZN => n27138);
   U24658 : NOR3_X1 port map( A1 => n26672, A2 => n17158, A3 => n36480, ZN => 
                           n14989);
   U24659 : NOR2_X1 port map( A1 => n1207, A2 => n34166, ZN => n20305);
   U24661 : NAND2_X1 port map( A1 => n3158, A2 => n13457, ZN => n21224);
   U24664 : NAND2_X1 port map( A1 => n27875, A2 => n17378, ZN => n27901);
   U24671 : NOR3_X1 port map( A1 => n17253, A2 => n1212, A3 => n15357, ZN => 
                           n17254);
   U24675 : NAND3_X1 port map( A1 => n17410, A2 => n988, A3 => n13081, ZN => 
                           n28075);
   U24677 : INV_X1 port map( I => n29223, ZN => n15395);
   U24680 : NAND2_X1 port map( A1 => n16343, A2 => n28598, ZN => n16272);
   U24682 : INV_X1 port map( I => n29034, ZN => n18523);
   U24683 : NAND2_X1 port map( A1 => n28577, A2 => n28674, ZN => n28307);
   U24684 : NAND2_X1 port map( A1 => n17644, A2 => n39830, ZN => n20288);
   U24686 : INV_X1 port map( I => n29768, ZN => n29692);
   U24687 : NOR2_X1 port map( A1 => n19424, A2 => n29900, ZN => n17779);
   U24688 : INV_X1 port map( I => n30233, ZN => n14891);
   U24691 : NAND2_X1 port map( A1 => n14428, A2 => n21269, ZN => n28880);
   U24693 : NOR2_X1 port map( A1 => n31444, A2 => n29774, ZN => n18221);
   U24695 : NOR2_X1 port map( A1 => n21285, A2 => n32571, ZN => n17632);
   U24696 : INV_X2 port map( I => n20080, ZN => n30043);
   U24698 : INV_X1 port map( I => n19050, ZN => n20251);
   U24699 : NAND2_X1 port map( A1 => n29438, A2 => n29439, ZN => n16960);
   U24701 : AOI21_X1 port map( A1 => n29543, A2 => n21072, B => n29559, ZN => 
                           n21071);
   U24702 : NAND2_X1 port map( A1 => n19272, A2 => n29548, ZN => n21072);
   U24703 : AOI21_X1 port map( A1 => n29546, A2 => n29548, B => n29558, ZN => 
                           n29542);
   U24704 : INV_X1 port map( I => n29558, ZN => n29550);
   U24706 : NAND2_X1 port map( A1 => n29567, A2 => n29574, ZN => n15308);
   U24707 : NAND2_X1 port map( A1 => n29797, A2 => n18257, ZN => n21012);
   U24710 : NAND2_X1 port map( A1 => n15466, A2 => n20277, ZN => n21058);
   U24712 : OAI21_X1 port map( A1 => n21666, A2 => n21833, B => n21436, ZN => 
                           n21361);
   U24716 : NOR2_X1 port map( A1 => n22019, A2 => n36006, ZN => n19958);
   U24717 : OAI22_X1 port map( A1 => n21431, A2 => n21682, B1 => n21681, B2 => 
                           n21683, ZN => n21356);
   U24718 : NAND2_X1 port map( A1 => n35973, A2 => n21681, ZN => n21354);
   U24721 : NAND3_X1 port map( A1 => n33771, A2 => n21762, A3 => n11851, ZN => 
                           n15613);
   U24723 : NAND2_X1 port map( A1 => n21964, A2 => n10261, ZN => n20043);
   U24727 : NAND2_X1 port map( A1 => n19850, A2 => n17102, ZN => n16231);
   U24730 : NAND2_X1 port map( A1 => n9970, A2 => n22234, ZN => n18064);
   U24731 : NOR2_X1 port map( A1 => n9970, A2 => n1329, ZN => n16228);
   U24735 : NAND2_X1 port map( A1 => n21863, A2 => n19609, ZN => n14995);
   U24739 : NOR2_X1 port map( A1 => n22236, A2 => n22235, ZN => n18129);
   U24743 : INV_X1 port map( I => n15268, ZN => n18272);
   U24748 : NAND2_X1 port map( A1 => n13855, A2 => n21885, ZN => n15816);
   U24750 : AOI21_X1 port map( A1 => n19416, A2 => n18266, B => n1353, ZN => 
                           n16762);
   U24753 : NOR2_X1 port map( A1 => n21656, A2 => n17938, ZN => n17433);
   U24757 : INV_X1 port map( I => n16347, ZN => n16345);
   U24758 : NOR2_X1 port map( A1 => n39594, A2 => n21478, ZN => n14945);
   U24761 : NOR2_X1 port map( A1 => n17869, A2 => n1676, ZN => n17334);
   U24763 : AOI21_X1 port map( A1 => n18657, A2 => n21924, B => n21923, ZN => 
                           n20844);
   U24765 : NOR2_X1 port map( A1 => n20681, A2 => n21837, ZN => n20680);
   U24767 : OAI21_X1 port map( A1 => n1372, A2 => n19709, B => n21703, ZN => 
                           n21704);
   U24768 : OAI21_X1 port map( A1 => n16302, A2 => n21887, B => n21889, ZN => 
                           n15929);
   U24770 : NOR2_X1 port map( A1 => n18542, A2 => n19543, ZN => n18561);
   U24772 : AOI21_X1 port map( A1 => n21591, A2 => n21590, B => n19434, ZN => 
                           n21598);
   U24773 : NAND2_X1 port map( A1 => n33086, A2 => n22262, ZN => n16625);
   U24774 : NAND2_X1 port map( A1 => n18926, A2 => n21920, ZN => n21736);
   U24776 : NOR2_X1 port map( A1 => n18205, A2 => n21528, ZN => n17967);
   U24777 : NAND2_X1 port map( A1 => n32525, A2 => n15560, ZN => n21657);
   U24779 : NOR2_X1 port map( A1 => n1354, A2 => n18028, ZN => n15560);
   U24780 : AND2_X1 port map( A1 => n22915, A2 => n23164, Z => n14628);
   U24781 : NOR2_X1 port map( A1 => n36095, A2 => n19293, ZN => n16604);
   U24782 : NAND2_X1 port map( A1 => n39418, A2 => n23171, ZN => n19177);
   U24784 : INV_X1 port map( I => n12392, ZN => n21292);
   U24793 : NAND2_X1 port map( A1 => n1310, A2 => n23637, ZN => n23471);
   U24794 : AOI21_X1 port map( A1 => n38604, A2 => n9699, B => n19229, ZN => 
                           n19228);
   U24796 : NOR2_X1 port map( A1 => n36839, A2 => n23213, ZN => n16198);
   U24798 : NAND2_X1 port map( A1 => n22918, A2 => n18679, ZN => n14738);
   U24801 : NAND2_X1 port map( A1 => n31234, A2 => n39070, ZN => n23194);
   U24805 : NAND2_X1 port map( A1 => n1300, A2 => n18236, ZN => n18235);
   U24807 : NOR2_X1 port map( A1 => n23548, A2 => n9321, ZN => n17674);
   U24814 : OAI21_X1 port map( A1 => n23184, A2 => n19538, B => n1314, ZN => 
                           n22965);
   U24815 : NAND2_X1 port map( A1 => n21094, A2 => n23098, ZN => n16956);
   U24816 : NOR2_X1 port map( A1 => n23060, A2 => n14560, ZN => n23062);
   U24817 : NAND2_X1 port map( A1 => n17127, A2 => n39810, ZN => n19083);
   U24818 : NOR2_X1 port map( A1 => n19823, A2 => n3452, ZN => n16615);
   U24819 : INV_X1 port map( I => n22870, ZN => n22998);
   U24820 : NAND3_X1 port map( A1 => n32815, A2 => n19293, A3 => n22996, ZN => 
                           n20214);
   U24821 : NOR2_X1 port map( A1 => n1648, A2 => n16104, ZN => n22894);
   U24822 : INV_X1 port map( I => n24065, ZN => n19102);
   U24823 : NOR2_X1 port map( A1 => n38282, A2 => n12029, ZN => n16419);
   U24825 : NAND2_X1 port map( A1 => n23087, A2 => n531, ZN => n23093);
   U24830 : AOI21_X1 port map( A1 => n31049, A2 => n19469, B => n1044, ZN => 
                           n15588);
   U24831 : NOR3_X1 port map( A1 => n20408, A2 => n23211, A3 => n20407, ZN => 
                           n21119);
   U24832 : INV_X1 port map( I => n20788, ZN => n23614);
   U24840 : NAND2_X1 port map( A1 => n15320, A2 => n11004, ZN => n24238);
   U24844 : INV_X1 port map( I => n24223, ZN => n20655);
   U24845 : NAND3_X1 port map( A1 => n14265, A2 => n24761, A3 => n33230, ZN => 
                           n20787);
   U24849 : NAND2_X1 port map( A1 => n24327, A2 => n1589, ZN => n16106);
   U24850 : NAND2_X1 port map( A1 => n19745, A2 => n24267, ZN => n16313);
   U24854 : NAND2_X1 port map( A1 => n24348, A2 => n24347, ZN => n24349);
   U24857 : OAI21_X1 port map( A1 => n20058, A2 => n37227, B => n24143, ZN => 
                           n24145);
   U24860 : NAND3_X1 port map( A1 => n24157, A2 => n24465, A3 => n17546, ZN => 
                           n24159);
   U24862 : NAND2_X1 port map( A1 => n23962, A2 => n6849, ZN => n21241);
   U24863 : NAND2_X1 port map( A1 => n24510, A2 => n24608, ZN => n15208);
   U24866 : NAND2_X1 port map( A1 => n24258, A2 => n38972, ZN => n19069);
   U24867 : NOR2_X1 port map( A1 => n34547, A2 => n20839, ZN => n18937);
   U24873 : AOI21_X1 port map( A1 => n24118, A2 => n24373, B => n24191, ZN => 
                           n18456);
   U24875 : NAND2_X1 port map( A1 => n17246, A2 => n955, ZN => n17451);
   U24879 : NAND2_X1 port map( A1 => n25106, A2 => n24896, ZN => n24895);
   U24884 : NOR2_X1 port map( A1 => n911, A2 => n19767, ZN => n20216);
   U24886 : OAI21_X1 port map( A1 => n17645, A2 => n9682, B => n26125, ZN => 
                           n14983);
   U24888 : NAND3_X1 port map( A1 => n25741, A2 => n25742, A3 => n596, ZN => 
                           n16137);
   U24899 : INV_X1 port map( I => n18031, ZN => n19514);
   U24902 : NOR2_X1 port map( A1 => n25431, A2 => n25649, ZN => n17182);
   U24908 : NAND2_X1 port map( A1 => n1102, A2 => n25965, ZN => n18038);
   U24909 : NOR2_X1 port map( A1 => n33644, A2 => n37502, ZN => n20235);
   U24914 : NAND2_X1 port map( A1 => n834, A2 => n17212, ZN => n15178);
   U24915 : NOR2_X1 port map( A1 => n25721, A2 => n18519, ZN => n25723);
   U24916 : NOR2_X1 port map( A1 => n2752, A2 => n35580, ZN => n26037);
   U24917 : NOR2_X1 port map( A1 => n20699, A2 => n32986, ZN => n20103);
   U24921 : NAND2_X1 port map( A1 => n26934, A2 => n17993, ZN => n19939);
   U24924 : NAND3_X1 port map( A1 => n12290, A2 => n26688, A3 => n26979, ZN => 
                           n26659);
   U24927 : NAND3_X1 port map( A1 => n12162, A2 => n25721, A3 => n33826, ZN => 
                           n25572);
   U24928 : OAI22_X1 port map( A1 => n26101, A2 => n35207, B1 => n25779, B2 => 
                           n25780, ZN => n20738);
   U24929 : NOR2_X1 port map( A1 => n25866, A2 => n2830, ZN => n25774);
   U24930 : NAND2_X1 port map( A1 => n1021, A2 => n35207, ZN => n16181);
   U24933 : NAND2_X1 port map( A1 => n34279, A2 => n39417, ZN => n17662);
   U24934 : NOR2_X1 port map( A1 => n17575, A2 => n33279, ZN => n17574);
   U24937 : NAND2_X1 port map( A1 => n32191, A2 => n38211, ZN => n20244);
   U24938 : NAND2_X1 port map( A1 => n26776, A2 => n38120, ZN => n21021);
   U24939 : NAND2_X1 port map( A1 => n19222, A2 => n26905, ZN => n15897);
   U24940 : INV_X1 port map( I => n27436, ZN => n16173);
   U24945 : NOR2_X1 port map( A1 => n33050, A2 => n27364, ZN => n18232);
   U24946 : NOR2_X1 port map( A1 => n1484, A2 => n34001, ZN => n19619);
   U24959 : NAND2_X1 port map( A1 => n31254, A2 => n26734, ZN => n21202);
   U24960 : INV_X1 port map( I => n7974, ZN => n27248);
   U24966 : NAND2_X1 port map( A1 => n4411, A2 => n17392, ZN => n17391);
   U24968 : OAI21_X1 port map( A1 => n14862, A2 => n20211, B => n14861, ZN => 
                           n20546);
   U24969 : INV_X1 port map( I => n26982, ZN => n26983);
   U24971 : NOR2_X1 port map( A1 => n26996, A2 => n13111, ZN => n17824);
   U24974 : INV_X1 port map( I => n19855, ZN => n28221);
   U24975 : AOI21_X1 port map( A1 => n26671, A2 => n33726, B => n11138, ZN => 
                           n14991);
   U24978 : INV_X1 port map( I => n20200, ZN => n20198);
   U24979 : NAND2_X1 port map( A1 => n20201, A2 => n20410, ZN => n20199);
   U24983 : NAND2_X1 port map( A1 => n28324, A2 => n33331, ZN => n27867);
   U24985 : NAND2_X1 port map( A1 => n17322, A2 => n28698, ZN => n19591);
   U24987 : NAND2_X1 port map( A1 => n3899, A2 => n37018, ZN => n19321);
   U24991 : NAND3_X1 port map( A1 => n28532, A2 => n38159, A3 => n11413, ZN => 
                           n28508);
   U24999 : NAND3_X1 port map( A1 => n28652, A2 => n28653, A3 => n28386, ZN => 
                           n28387);
   U25000 : NAND2_X1 port map( A1 => n18341, A2 => n19039, ZN => n28327);
   U25001 : NOR2_X1 port map( A1 => n28283, A2 => n28282, ZN => n20398);
   U25002 : AOI21_X1 port map( A1 => n1426, A2 => n3014, B => n1415, ZN => 
                           n19795);
   U25003 : AND2_X1 port map( A1 => n18036, A2 => n28656, Z => n14621);
   U25005 : NAND2_X1 port map( A1 => n28310, A2 => n28723, ZN => n14816);
   U25006 : NOR2_X1 port map( A1 => n28724, A2 => n28722, ZN => n28310);
   U25011 : NOR2_X1 port map( A1 => n1397, A2 => n10702, ZN => n16988);
   U25013 : NAND2_X1 port map( A1 => n20830, A2 => n29455, ZN => n29457);
   U25015 : NAND2_X1 port map( A1 => n29764, A2 => n29696, ZN => n29636);
   U25018 : NOR2_X1 port map( A1 => n29698, A2 => n1060, ZN => n16392);
   U25019 : OAI21_X1 port map( A1 => n29761, A2 => n31516, B => n19567, ZN => 
                           n29697);
   U25020 : AOI21_X1 port map( A1 => n31516, A2 => n19568, B => n19599, ZN => 
                           n19567);
   U25021 : INV_X1 port map( I => n29940, ZN => n29989);
   U25025 : OAI21_X1 port map( A1 => n1387, A2 => n1388, B => n29236, ZN => 
                           n15482);
   U25026 : NOR2_X1 port map( A1 => n907, A2 => n19088, ZN => n17821);
   U25027 : NAND2_X1 port map( A1 => n29351, A2 => n12876, ZN => n29309);
   U25028 : AOI21_X1 port map( A1 => n1055, A2 => n29314, B => n29313, ZN => 
                           n19130);
   U25029 : NAND2_X1 port map( A1 => n29315, A2 => n357, ZN => n19129);
   U25030 : NOR2_X1 port map( A1 => n16123, A2 => n29317, ZN => n14787);
   U25031 : NAND2_X1 port map( A1 => n12943, A2 => n29367, ZN => n29373);
   U25034 : NAND2_X1 port map( A1 => n38200, A2 => n29478, ZN => n29462);
   U25038 : NAND2_X1 port map( A1 => n28619, A2 => n505, ZN => n18726);
   U25040 : NAND2_X1 port map( A1 => n1390, A2 => n29664, ZN => n16596);
   U25041 : NAND2_X1 port map( A1 => n29641, A2 => n29660, ZN => n21033);
   U25045 : NAND2_X1 port map( A1 => n17684, A2 => n33358, ZN => n17683);
   U25046 : AOI22_X1 port map( A1 => n17681, A2 => n4849, B1 => n39830, B2 => 
                           n21023, ZN => n16996);
   U25048 : OAI21_X1 port map( A1 => n29761, A2 => n29760, B => n16962, ZN => 
                           n29767);
   U25049 : NOR2_X1 port map( A1 => n29763, A2 => n17105, ZN => n16962);
   U25051 : NAND2_X1 port map( A1 => n1063, A2 => n29870, ZN => n19393);
   U25052 : NAND2_X1 port map( A1 => n19093, A2 => n18104, ZN => n15138);
   U25053 : INV_X1 port map( I => n28980, ZN => n15141);
   U25056 : NAND2_X1 port map( A1 => n29949, A2 => n35809, ZN => n29951);
   U25057 : NAND2_X1 port map( A1 => n21166, A2 => n30058, ZN => n17982);
   U25058 : NOR2_X1 port map( A1 => n11861, A2 => n29996, ZN => n17633);
   U25060 : NAND2_X1 port map( A1 => n16180, A2 => n35187, ZN => n16722);
   U25063 : INV_X1 port map( I => n32415, ZN => n29183);
   U25064 : NOR2_X1 port map( A1 => n30177, A2 => n20342, ZN => n14998);
   U25066 : NOR2_X1 port map( A1 => n37659, A2 => n33280, ZN => n18755);
   U25070 : OAI21_X1 port map( A1 => n16016, A2 => n2532, B => n21889, ZN => 
                           n16014);
   U25075 : INV_X1 port map( I => n1048, ZN => n17639);
   U25079 : NOR2_X1 port map( A1 => n36237, A2 => n20799, ZN => n20798);
   U25080 : NAND2_X1 port map( A1 => n17940, A2 => n15175, ZN => n17939);
   U25081 : NAND2_X1 port map( A1 => n9970, A2 => n20943, ZN => n22061);
   U25082 : NAND2_X1 port map( A1 => n16262, A2 => n21288, ZN => n16453);
   U25084 : NOR2_X1 port map( A1 => n1152, A2 => n16265, ZN => n16452);
   U25085 : INV_X1 port map( I => n2233, ZN => n22445);
   U25086 : INV_X1 port map( I => n22495, ZN => n18189);
   U25087 : NAND3_X1 port map( A1 => n22209, A2 => n30315, A3 => n22208, ZN => 
                           n22210);
   U25090 : NAND2_X1 port map( A1 => n22345, A2 => n22341, ZN => n21967);
   U25098 : INV_X1 port map( I => n16348, ZN => n16346);
   U25099 : INV_X1 port map( I => n22645, ZN => n20718);
   U25100 : NAND2_X1 port map( A1 => n22190, A2 => n9987, ZN => n22191);
   U25101 : OAI21_X1 port map( A1 => n19486, A2 => n22189, B => n9987, ZN => 
                           n22193);
   U25102 : INV_X1 port map( I => n22743, ZN => n17513);
   U25103 : NAND2_X1 port map( A1 => n17341, A2 => n30323, ZN => n17339);
   U25105 : NAND3_X1 port map( A1 => n30315, A2 => n22204, A3 => n21288, ZN => 
                           n22096);
   U25110 : INV_X1 port map( I => n22043, ZN => n17668);
   U25111 : INV_X1 port map( I => n22044, ZN => n17669);
   U25112 : NAND2_X1 port map( A1 => n22944, A2 => n23166, ZN => n16955);
   U25127 : NAND3_X1 port map( A1 => n4147, A2 => n17887, A3 => n23493, ZN => 
                           n22970);
   U25128 : INV_X1 port map( I => n32226, ZN => n20503);
   U25130 : AOI21_X1 port map( A1 => n15579, A2 => n23461, B => n23238, ZN => 
                           n20322);
   U25132 : AOI21_X1 port map( A1 => n22988, A2 => n1135, B => n36829, ZN => 
                           n16032);
   U25135 : NOR2_X1 port map( A1 => n19481, A2 => n19686, ZN => n21118);
   U25137 : NAND2_X1 port map( A1 => n20817, A2 => n39001, ZN => n18389);
   U25141 : NAND2_X1 port map( A1 => n23547, A2 => n1295, ZN => n17677);
   U25143 : AND2_X1 port map( A1 => n1038, A2 => n23515, Z => n14665);
   U25148 : NAND2_X1 port map( A1 => n23264, A2 => n38724, ZN => n16058);
   U25151 : OAI21_X1 port map( A1 => n16443, A2 => n34307, B => n35068, ZN => 
                           n23557);
   U25155 : AOI22_X1 port map( A1 => n20661, A2 => n20343, B1 => n17511, B2 => 
                           n23477, ZN => n23466);
   U25156 : INV_X1 port map( I => n23969, ZN => n23698);
   U25159 : NAND2_X1 port map( A1 => n23630, A2 => n39070, ZN => n19922);
   U25161 : NOR2_X1 port map( A1 => n23351, A2 => n17090, ZN => n14720);
   U25162 : NAND2_X1 port map( A1 => n20100, A2 => n31331, ZN => n23118);
   U25163 : INV_X1 port map( I => n23762, ZN => n18172);
   U25165 : OAI21_X1 port map( A1 => n23039, A2 => n20620, B => n15797, ZN => 
                           n15800);
   U25166 : NOR2_X1 port map( A1 => n15949, A2 => n15798, ZN => n15797);
   U25167 : NOR2_X1 port map( A1 => n17995, A2 => n20620, ZN => n15798);
   U25169 : OAI21_X1 port map( A1 => n20002, A2 => n15210, B => n39067, ZN => 
                           n18552);
   U25170 : NOR2_X1 port map( A1 => n19466, A2 => n21310, ZN => n18551);
   U25171 : INV_X1 port map( I => n24669, ZN => n24670);
   U25172 : NOR2_X1 port map( A1 => n24668, A2 => n3076, ZN => n24671);
   U25174 : AND2_X1 port map( A1 => n20787, A2 => n24762, Z => n14548);
   U25181 : INV_X1 port map( I => n24965, ZN => n16421);
   U25185 : AND2_X1 port map( A1 => n37229, A2 => n24433, Z => n14538);
   U25186 : NAND2_X1 port map( A1 => n20027, A2 => n24271, ZN => n19690);
   U25187 : AOI21_X1 port map( A1 => n24738, A2 => n24737, B => n37389, ZN => 
                           n16670);
   U25191 : NAND2_X1 port map( A1 => n24117, A2 => n16547, ZN => n16785);
   U25193 : INV_X1 port map( I => n16900, ZN => n15158);
   U25194 : NAND3_X1 port map( A1 => n9892, A2 => n1240, A3 => n931, ZN => 
                           n26326);
   U25195 : AOI22_X1 port map( A1 => n1515, A2 => n26330, B1 => n14407, B2 => 
                           n9892, ZN => n15194);
   U25197 : INV_X1 port map( I => n17891, ZN => n24606);
   U25200 : INV_X1 port map( I => n16542, ZN => n16540);
   U25201 : INV_X1 port map( I => n17613, ZN => n25347);
   U25216 : OAI21_X1 port map( A1 => n31557, A2 => n25689, B => n25690, ZN => 
                           n18146);
   U25218 : NAND2_X1 port map( A1 => n25803, A2 => n25965, ZN => n25585);
   U25220 : NOR2_X1 port map( A1 => n4699, A2 => n26098, ZN => n25785);
   U25221 : NAND2_X1 port map( A1 => n1528, A2 => n11848, ZN => n25817);
   U25222 : INV_X1 port map( I => n17372, ZN => n17261);
   U25223 : NAND2_X1 port map( A1 => n951, A2 => n26109, ZN => n14810);
   U25224 : INV_X1 port map( I => n35209, ZN => n18371);
   U25225 : NOR2_X1 port map( A1 => n25812, A2 => n26131, ZN => n21305);
   U25226 : NAND2_X1 port map( A1 => n1097, A2 => n4604, ZN => n18282);
   U25232 : INV_X1 port map( I => n26006, ZN => n20051);
   U25241 : INV_X1 port map( I => n25841, ZN => n16424);
   U25243 : NOR2_X1 port map( A1 => n27054, A2 => n27341, ZN => n20915);
   U25244 : NOR2_X1 port map( A1 => n25803, A2 => n25965, ZN => n18037);
   U25245 : NAND2_X1 port map( A1 => n19980, A2 => n12162, ZN => n25559);
   U25246 : NOR2_X1 port map( A1 => n25558, A2 => n25557, ZN => n19980);
   U25250 : OAI21_X1 port map( A1 => n27230, A2 => n27415, B => n27109, ZN => 
                           n15915);
   U25252 : NAND2_X1 port map( A1 => n39065, A2 => n27069, ZN => n20145);
   U25261 : NAND2_X1 port map( A1 => n20738, A2 => n32193, ZN => n15869);
   U25265 : NAND2_X1 port map( A1 => n8696, A2 => n27586, ZN => n27041);
   U25266 : INV_X1 port map( I => n19352, ZN => n27175);
   U25270 : OAI21_X1 port map( A1 => n15433, A2 => n15434, B => n15432, ZN => 
                           n15430);
   U25273 : INV_X1 port map( I => n27076, ZN => n18170);
   U25274 : INV_X1 port map( I => n27441, ZN => n27444);
   U25275 : OAI21_X1 port map( A1 => n27306, A2 => n27583, B => n27585, ZN => 
                           n27307);
   U25278 : NAND2_X1 port map( A1 => n38571, A2 => n7291, ZN => n27146);
   U25279 : NAND2_X1 port map( A1 => n27145, A2 => n7291, ZN => n17058);
   U25283 : NAND3_X1 port map( A1 => n27429, A2 => n27428, A3 => n12156, ZN => 
                           n27431);
   U25284 : OR2_X1 port map( A1 => n27167, A2 => n27166, Z => n14586);
   U25291 : INV_X1 port map( I => n16848, ZN => n19669);
   U25295 : INV_X1 port map( I => n28650, ZN => n18961);
   U25296 : NAND2_X1 port map( A1 => n32543, A2 => n28484, ZN => n28483);
   U25297 : NAND3_X1 port map( A1 => n28756, A2 => n28755, A3 => n16691, ZN => 
                           n28757);
   U25298 : NAND2_X1 port map( A1 => n28666, A2 => n28665, ZN => n21212);
   U25303 : NAND2_X1 port map( A1 => n37956, A2 => n14968, ZN => n14967);
   U25305 : INV_X1 port map( I => n29142, ZN => n21056);
   U25309 : INV_X1 port map( I => n15015, ZN => n28670);
   U25312 : NAND2_X1 port map( A1 => n28061, A2 => n28060, ZN => n28062);
   U25315 : NOR2_X1 port map( A1 => n18472, A2 => n18471, ZN => n18470);
   U25316 : NOR2_X1 port map( A1 => n28758, A2 => n978, ZN => n19055);
   U25322 : NAND2_X1 port map( A1 => n28323, A2 => n30304, ZN => n19754);
   U25325 : INV_X1 port map( I => n28943, ZN => n16640);
   U25328 : OAI21_X1 port map( A1 => n20931, A2 => n8805, B => n37013, ZN => 
                           n29006);
   U25332 : NAND2_X1 port map( A1 => n28715, A2 => n19844, ZN => n28210);
   U25335 : NOR2_X1 port map( A1 => n29777, A2 => n29781, ZN => n21037);
   U25337 : INV_X1 port map( I => n35272, ZN => n29390);
   U25340 : NAND2_X1 port map( A1 => n29525, A2 => n29535, ZN => n16084);
   U25341 : NAND2_X1 port map( A1 => n29546, A2 => n29558, ZN => n19380);
   U25342 : NAND2_X1 port map( A1 => n29721, A2 => n29720, ZN => n17731);
   U25343 : NAND2_X1 port map( A1 => n30022, A2 => n9231, ZN => n18782);
   U25345 : NOR2_X1 port map( A1 => n30109, A2 => n35186, ZN => n19032);
   U25348 : OAI21_X1 port map( A1 => n18611, A2 => n29274, B => n19090, ZN => 
                           n17955);
   U25353 : NOR2_X1 port map( A1 => n29409, A2 => n17849, ZN => n29405);
   U25354 : AOI21_X1 port map( A1 => n29423, A2 => n29440, B => n1383, ZN => 
                           n19618);
   U25355 : NAND2_X1 port map( A1 => n1389, A2 => n29438, ZN => n15127);
   U25356 : NOR2_X1 port map( A1 => n29440, A2 => n17293, ZN => n15128);
   U25357 : NAND2_X1 port map( A1 => n29540, A2 => n29550, ZN => n28906);
   U25359 : OAI21_X1 port map( A1 => n29570, A2 => n29571, B => n1393, ZN => 
                           n20701);
   U25360 : NAND3_X1 port map( A1 => n29570, A2 => n31899, A3 => n29571, ZN => 
                           n15310);
   U25362 : NOR2_X1 port map( A1 => n30295, A2 => n19318, ZN => n29656);
   U25363 : NOR3_X1 port map( A1 => n6181, A2 => n19297, A3 => n39689, ZN => 
                           n21032);
   U25364 : NOR2_X1 port map( A1 => n21033, A2 => n19318, ZN => n20444);
   U25366 : INV_X1 port map( I => n18042, ZN => n29686);
   U25368 : NAND3_X1 port map( A1 => n20498, A2 => n5921, A3 => n29722, ZN => 
                           n20499);
   U25369 : AOI21_X1 port map( A1 => n21013, A2 => n29788, B => n21010, ZN => 
                           n21009);
   U25371 : NAND2_X1 port map( A1 => n18085, A2 => n18082, ZN => n29915);
   U25373 : INV_X1 port map( I => n30078, ZN => n19550);
   U25374 : AOI21_X1 port map( A1 => n16723, A2 => n30111, B => n16721, ZN => 
                           n16720);
   U25377 : AOI21_X1 port map( A1 => n10289, A2 => n31527, B => n17192, ZN => 
                           n21006);
   U25378 : AOI21_X1 port map( A1 => n13384, A2 => n10813, B => n17193, ZN => 
                           n21005);
   U25379 : NAND2_X1 port map( A1 => n20538, A2 => n14998, ZN => n14997);
   U25380 : NAND2_X1 port map( A1 => n30176, A2 => n17997, ZN => n17168);
   U25386 : OR2_X1 port map( A1 => n16052, A2 => n21606, Z => n14420);
   U25389 : OR2_X1 port map( A1 => n25387, A2 => n25386, Z => n14431);
   U25390 : NAND2_X1 port map( A1 => n1177, A2 => n10569, ZN => n14435);
   U25399 : NOR2_X1 port map( A1 => n21885, A2 => n15839, ZN => n14492);
   U25400 : XOR2_X1 port map( A1 => n22781, A2 => n22780, Z => n14494);
   U25404 : XNOR2_X1 port map( A1 => n24861, A2 => n24860, ZN => n14507);
   U25407 : OR2_X1 port map( A1 => n1076, A2 => n28150, Z => n14513);
   U25408 : OR2_X1 port map( A1 => n25690, A2 => n25689, Z => n14518);
   U25410 : OR2_X1 port map( A1 => n29675, A2 => n29683, Z => n14522);
   U25412 : XNOR2_X1 port map( A1 => n10027, A2 => n22749, ZN => n14530);
   U25414 : XNOR2_X1 port map( A1 => n9576, A2 => n19875, ZN => n14533);
   U25416 : INV_X1 port map( I => n19819, ZN => n22565);
   U25418 : INV_X1 port map( I => n37229, ZN => n24434);
   U25419 : AND2_X1 port map( A1 => n35357, A2 => n28812, Z => n14543);
   U25421 : AND2_X1 port map( A1 => n15194, A2 => n26332, Z => n14546);
   U25422 : INV_X1 port map( I => n22674, ZN => n23135);
   U25424 : NOR2_X1 port map( A1 => n8700, A2 => n19350, ZN => n14549);
   U25425 : AND2_X1 port map( A1 => n19850, A2 => n21887, Z => n14551);
   U25428 : XNOR2_X1 port map( A1 => n38184, A2 => n35267, ZN => n14565);
   U25430 : INV_X1 port map( I => n29696, ZN => n19568);
   U25431 : XNOR2_X1 port map( A1 => n14264, A2 => n20706, ZN => n14566);
   U25433 : XNOR2_X1 port map( A1 => n33194, A2 => n30207, ZN => n14568);
   U25434 : XNOR2_X1 port map( A1 => n23357, A2 => n1621, ZN => n14571);
   U25436 : AND2_X1 port map( A1 => n18884, A2 => n11848, Z => n14579);
   U25437 : BUF_X2 port map( I => n21655, Z => n17938);
   U25438 : AND2_X1 port map( A1 => n17943, A2 => n29411, Z => n14582);
   U25442 : INV_X1 port map( I => n22204, ZN => n22351);
   U25443 : OR2_X1 port map( A1 => n24687, A2 => n14857, Z => n14593);
   U25444 : AND2_X1 port map( A1 => n23107, A2 => n22005, Z => n14594);
   U25445 : NAND2_X1 port map( A1 => n22101, A2 => n20234, ZN => n14597);
   U25449 : XNOR2_X1 port map( A1 => n16017, A2 => n19775, ZN => n14603);
   U25458 : AND2_X1 port map( A1 => n27163, A2 => n20981, Z => n14626);
   U25459 : AND2_X1 port map( A1 => n20919, A2 => n28053, Z => n14632);
   U25463 : INV_X1 port map( I => n314, ZN => n21073);
   U25467 : XNOR2_X1 port map( A1 => n25094, A2 => n25095, ZN => n14646);
   U25469 : XNOR2_X1 port map( A1 => n19221, A2 => n20479, ZN => n14648);
   U25470 : XNOR2_X1 port map( A1 => n24002, A2 => n1723, ZN => n14651);
   U25473 : XNOR2_X1 port map( A1 => n39063, A2 => n19913, ZN => n14670);
   U25476 : XNOR2_X1 port map( A1 => n22790, A2 => n29707, ZN => n14673);
   U25478 : INV_X1 port map( I => n21880, ZN => n21509);
   U25479 : XNOR2_X1 port map( A1 => n26394, A2 => n28934, ZN => n14675);
   U25482 : INV_X1 port map( I => n25502, ZN => n15647);
   U25484 : INV_X1 port map( I => n22773, ZN => n16531);
   U25487 : XNOR2_X1 port map( A1 => n29252, A2 => n1734, ZN => n14689);
   U25488 : XNOR2_X1 port map( A1 => n20311, A2 => n20310, ZN => n14691);
   U25491 : XNOR2_X1 port map( A1 => n27746, A2 => n35702, ZN => n14693);
   U25492 : NOR2_X1 port map( A1 => n438, A2 => n759, ZN => n14696);
   U25499 : INV_X1 port map( I => n27129, ZN => n20402);
   U25501 : INV_X1 port map( I => n19879, ZN => n17078);
   U25502 : INV_X1 port map( I => n19760, ZN => n18981);
   U25503 : INV_X1 port map( I => n19937, ZN => n20206);
   U25504 : INV_X1 port map( I => n19876, ZN => n16320);
   U25505 : INV_X1 port map( I => n29554, ZN => n21121);
   U25506 : INV_X1 port map( I => n30090, ZN => n18109);
   U25507 : INV_X1 port map( I => n19866, ZN => n17603);
   U25509 : INV_X1 port map( I => n19808, ZN => n20658);
   U25510 : INV_X1 port map( I => n9981, ZN => n18432);
   U25511 : INV_X1 port map( I => n10027, ZN => n16618);
   U25512 : INV_X1 port map( I => n29411, ZN => n17551);
   U25513 : INV_X1 port map( I => n30169, ZN => n15203);
   U25517 : INV_X1 port map( I => n19936, ZN => n16562);
   U25518 : INV_X1 port map( I => n19613, ZN => n16332);
   U25520 : INV_X1 port map( I => n29221, ZN => n17257);
   U25521 : INV_X1 port map( I => n19860, ZN => n17463);
   U25522 : INV_X1 port map( I => n29269, ZN => n19128);
   U25524 : INV_X1 port map( I => n30068, ZN => n21294);
   U25525 : INV_X1 port map( I => n30248, ZN => n18296);
   U25526 : INV_X1 port map( I => n29602, ZN => n15432);
   U25527 : BUF_X2 port map( I => Key(65), Z => n29801);
   U25532 : XOR2_X1 port map( A1 => n19862, A2 => n29320, Z => n18015);
   U25536 : XOR2_X1 port map( A1 => n25246, A2 => n14716, Z => n14715);
   U25537 : XOR2_X1 port map( A1 => n19156, A2 => n25280, Z => n14716);
   U25538 : XOR2_X1 port map( A1 => n16318, A2 => n16321, Z => n24308);
   U25540 : NOR2_X1 port map( A1 => n8597, A2 => n21587, ZN => n21589);
   U25541 : AOI21_X2 port map( A1 => n15491, A2 => n14721, B => n14720, ZN => 
                           n23667);
   U25543 : NOR2_X1 port map( A1 => n22964, A2 => n14725, ZN => n15084);
   U25550 : XOR2_X1 port map( A1 => n27594, A2 => n15776, Z => n14756);
   U25551 : INV_X2 port map( I => n14758, ZN => n22682);
   U25552 : NOR2_X1 port map( A1 => n23533, A2 => n14759, ZN => n16395);
   U25553 : XOR2_X1 port map( A1 => n18273, A2 => n39183, Z => n19493);
   U25555 : NAND2_X1 port map( A1 => n25946, A2 => n39729, ZN => n14762);
   U25556 : XOR2_X1 port map( A1 => n15288, A2 => n14772, Z => n14771);
   U25561 : XOR2_X1 port map( A1 => n15165, A2 => n24999, Z => n25087);
   U25563 : XOR2_X1 port map( A1 => Plaintext(171), A2 => Key(171), Z => n15370
                           );
   U25564 : OR2_X1 port map( A1 => n20021, A2 => n14488, Z => n14798);
   U25569 : NAND2_X1 port map( A1 => n1126, A2 => n19864, ZN => n24069);
   U25575 : XOR2_X1 port map( A1 => n14808, A2 => n27834, Z => n27472);
   U25577 : XOR2_X1 port map( A1 => n14818, A2 => n14821, Z => n19806);
   U25578 : XOR2_X1 port map( A1 => n24058, A2 => n14819, Z => n14818);
   U25582 : XOR2_X1 port map( A1 => Plaintext(173), A2 => Key(173), Z => n15152
                           );
   U25585 : MUX2_X1 port map( I0 => n28647, I1 => n15296, S => n30805, Z => 
                           n15295);
   U25586 : XOR2_X1 port map( A1 => n29027, A2 => n14844, Z => n14843);
   U25587 : XOR2_X1 port map( A1 => n19513, A2 => n14956, Z => n14844);
   U25591 : XOR2_X1 port map( A1 => n25101, A2 => n14859, Z => n18121);
   U25592 : XOR2_X1 port map( A1 => n7728, A2 => n16492, Z => n25100);
   U25595 : XOR2_X1 port map( A1 => n26511, A2 => n26510, Z => n14867);
   U25600 : XOR2_X1 port map( A1 => n14425, A2 => n24919, Z => n24920);
   U25602 : NAND2_X1 port map( A1 => n23595, A2 => n23596, ZN => n23314);
   U25605 : XOR2_X1 port map( A1 => n35231, A2 => n1734, Z => n14887);
   U25606 : XOR2_X1 port map( A1 => n22465, A2 => n22600, Z => n14888);
   U25609 : NAND2_X1 port map( A1 => n39322, A2 => n14891, ZN => n29203);
   U25612 : XOR2_X1 port map( A1 => n2233, A2 => n19735, Z => n14894);
   U25615 : NOR2_X1 port map( A1 => n28559, A2 => n1197, ZN => n14900);
   U25618 : XOR2_X1 port map( A1 => n27855, A2 => n19885, Z => n14907);
   U25620 : NOR2_X1 port map( A1 => n1158, A2 => n21837, ZN => n14911);
   U25623 : XOR2_X1 port map( A1 => n18974, A2 => n18973, Z => n26668);
   U25630 : XOR2_X1 port map( A1 => n24018, A2 => n35196, Z => n23981);
   U25632 : NAND2_X2 port map( A1 => n25516, A2 => n19209, ZN => n25798);
   U25638 : XOR2_X1 port map( A1 => n28953, A2 => n14956, Z => n28813);
   U25640 : XOR2_X1 port map( A1 => n25071, A2 => n14970, Z => n17457);
   U25643 : XOR2_X1 port map( A1 => n26348, A2 => n1096, Z => n14978);
   U25644 : INV_X1 port map( I => n23992, ZN => n24311);
   U25645 : XOR2_X1 port map( A1 => n22703, A2 => n4413, Z => n14979);
   U25646 : NOR2_X2 port map( A1 => n21976, A2 => n17027, ZN => n19931);
   U25647 : INV_X2 port map( I => n19685, ZN => n23028);
   U25648 : XNOR2_X1 port map( A1 => n14981, A2 => n14982, ZN => n14980);
   U25650 : XOR2_X1 port map( A1 => n18127, A2 => n29097, Z => n14982);
   U25651 : OAI22_X1 port map( A1 => n3826, A2 => n17158, B1 => n11226, B2 => 
                           n38377, ZN => n26829);
   U25654 : OAI21_X1 port map( A1 => n15269, A2 => n14500, B => n33516, ZN => 
                           n28013);
   U25655 : NAND3_X2 port map( A1 => n17221, A2 => n27093, A3 => n27094, ZN => 
                           n17220);
   U25656 : INV_X1 port map( I => n15007, ZN => n15006);
   U25658 : XOR2_X1 port map( A1 => n15012, A2 => n21278, Z => n22674);
   U25660 : XOR2_X1 port map( A1 => n38850, A2 => n19592, Z => n15013);
   U25661 : OAI22_X1 port map( A1 => n28800, A2 => n28799, B1 => n19905, B2 => 
                           n15015, ZN => n28801);
   U25662 : NAND2_X1 port map( A1 => n15015, A2 => n19905, ZN => n28800);
   U25664 : OAI21_X1 port map( A1 => n21950, A2 => n32664, B => n15019, ZN => 
                           n21952);
   U25666 : XOR2_X1 port map( A1 => n27516, A2 => n35188, Z => n27169);
   U25669 : INV_X2 port map( I => n15036, ZN => n25660);
   U25672 : INV_X2 port map( I => n15052, ZN => n25481);
   U25674 : AOI21_X2 port map( A1 => n18340, A2 => n15053, B => n18338, ZN => 
                           n22058);
   U25677 : XOR2_X1 port map( A1 => n38158, A2 => n35266, Z => n15056);
   U25678 : NOR2_X2 port map( A1 => n32791, A2 => n28753, ZN => n28754);
   U25679 : XOR2_X1 port map( A1 => n17423, A2 => n18849, Z => n15972);
   U25680 : XOR2_X1 port map( A1 => n25163, A2 => n33184, Z => n18643);
   U25681 : XOR2_X1 port map( A1 => n38951, A2 => n15888, Z => n15753);
   U25682 : OAI21_X1 port map( A1 => n29497, A2 => n15063, B => n29498, ZN => 
                           n20720);
   U25683 : NOR2_X1 port map( A1 => n38051, A2 => n17424, ZN => n15063);
   U25685 : XOR2_X1 port map( A1 => n28603, A2 => n28607, Z => n15071);
   U25686 : NAND2_X1 port map( A1 => n19871, A2 => n20703, ZN => n21654);
   U25687 : OAI22_X1 port map( A1 => n21904, A2 => n21903, B1 => n21900, B2 => 
                           n21902, ZN => n15072);
   U25689 : NOR2_X1 port map( A1 => n36530, A2 => n15075, ZN => n15074);
   U25692 : MUX2_X1 port map( I0 => n27484, I1 => n1218, S => n3977, Z => 
                           n27485);
   U25696 : XOR2_X1 port map( A1 => n29297, A2 => n4816, Z => n15090);
   U25699 : XOR2_X1 port map( A1 => n37874, A2 => n29295, Z => n15093);
   U25700 : XOR2_X1 port map( A1 => n23931, A2 => n19732, Z => n15094);
   U25703 : AOI21_X1 port map( A1 => n28717, A2 => n28716, B => n5093, ZN => 
                           n27941);
   U25710 : XOR2_X1 port map( A1 => n15126, A2 => n18584, Z => n15516);
   U25712 : OAI21_X1 port map( A1 => n29435, A2 => n29437, B => n11506, ZN => 
                           n15132);
   U25714 : AOI21_X1 port map( A1 => n29960, A2 => n29957, B => n15140, ZN => 
                           n15139);
   U25719 : INV_X2 port map( I => n15152, ZN => n18293);
   U25720 : XOR2_X1 port map( A1 => n15156, A2 => n19629, Z => n28710);
   U25721 : XOR2_X1 port map( A1 => n15156, A2 => n20804, Z => n29155);
   U25723 : OR2_X1 port map( A1 => n22976, A2 => n15163, Z => n21245);
   U25725 : XOR2_X1 port map( A1 => n22749, A2 => n1700, Z => n15171);
   U25730 : XOR2_X1 port map( A1 => Plaintext(144), A2 => Key(144), Z => n15619
                           );
   U25733 : XOR2_X1 port map( A1 => n15186, A2 => n1377, Z => n15226);
   U25737 : INV_X2 port map( I => n27985, ZN => n28054);
   U25738 : INV_X2 port map( I => n15195, ZN => n21254);
   U25740 : XOR2_X1 port map( A1 => n27858, A2 => n19932, Z => n15197);
   U25744 : OAI21_X1 port map( A1 => n15209, A2 => n17262, B => n29574, ZN => 
                           n29575);
   U25748 : NOR2_X1 port map( A1 => n1126, A2 => n21310, ZN => n15210);
   U25749 : NOR2_X2 port map( A1 => n16467, A2 => n27921, ZN => n19844);
   U25750 : XOR2_X1 port map( A1 => n15213, A2 => n15212, Z => n18308);
   U25751 : XOR2_X1 port map( A1 => n22557, A2 => n22556, Z => n15212);
   U25752 : XOR2_X1 port map( A1 => n18778, A2 => n22629, Z => n22556);
   U25753 : XOR2_X1 port map( A1 => n22411, A2 => n36290, Z => n22557);
   U25754 : XOR2_X1 port map( A1 => n17987, A2 => n15214, Z => n15213);
   U25756 : XOR2_X1 port map( A1 => n28860, A2 => n28946, Z => n21271);
   U25757 : XOR2_X1 port map( A1 => n28827, A2 => n19741, Z => n28860);
   U25758 : XOR2_X1 port map( A1 => n15216, A2 => n28777, Z => n16554);
   U25759 : XOR2_X1 port map( A1 => n15220, A2 => n19986, Z => n15938);
   U25762 : XOR2_X1 port map( A1 => n21380, A2 => Key(130), Z => n21761);
   U25765 : XOR2_X1 port map( A1 => n17606, A2 => n25217, Z => n15227);
   U25767 : NAND2_X2 port map( A1 => n19999, A2 => n20000, ZN => n25127);
   U25770 : NAND2_X1 port map( A1 => n15233, A2 => n19362, ZN => n15232);
   U25774 : INV_X2 port map( I => n18308, ZN => n22929);
   U25776 : NAND2_X1 port map( A1 => n24193, A2 => n15240, ZN => n16882);
   U25781 : XOR2_X1 port map( A1 => n14454, A2 => n23280, Z => n15250);
   U25783 : NAND3_X1 port map( A1 => n24359, A2 => n24360, A3 => n38431, ZN => 
                           n15257);
   U25790 : XOR2_X1 port map( A1 => n27842, A2 => n31438, Z => n15286);
   U25791 : XOR2_X1 port map( A1 => Plaintext(172), A2 => Key(172), Z => n18968
                           );
   U25795 : XOR2_X1 port map( A1 => n28925, A2 => n3633, Z => n15303);
   U25797 : XOR2_X1 port map( A1 => n14638, A2 => n14476, Z => n15305);
   U25798 : NAND2_X1 port map( A1 => n29571, A2 => n29570, ZN => n29563);
   U25801 : XOR2_X1 port map( A1 => n15316, A2 => n15315, Z => n18544);
   U25802 : XOR2_X1 port map( A1 => n25093, A2 => n24931, Z => n15315);
   U25807 : MUX2_X1 port map( I0 => n15172, I1 => n9751, S => n15443, Z => 
                           n15444);
   U25811 : XOR2_X1 port map( A1 => n15340, A2 => n22621, Z => n15339);
   U25812 : XOR2_X1 port map( A1 => n22647, A2 => n19755, Z => n15340);
   U25815 : XOR2_X1 port map( A1 => n871, A2 => n15349, Z => n15348);
   U25816 : XOR2_X1 port map( A1 => n27730, A2 => n19763, Z => n15349);
   U25818 : OAI22_X1 port map( A1 => n18558, A2 => n15350, B1 => n9876, B2 => 
                           n22341, ZN => n19270);
   U25820 : NOR2_X1 port map( A1 => n36754, A2 => n11274, ZN => n21573);
   U25823 : XOR2_X1 port map( A1 => n10647, A2 => n14565, Z => n15361);
   U25825 : NOR2_X1 port map( A1 => n14783, A2 => n19372, ZN => n21629);
   U25826 : NAND2_X1 port map( A1 => n18968, A2 => n14783, ZN => n21726);
   U25830 : NOR2_X1 port map( A1 => n17792, A2 => n19397, ZN => n15381);
   U25831 : NAND2_X1 port map( A1 => n29687, A2 => n38206, ZN => n29667);
   U25832 : INV_X2 port map( I => n19741, ZN => n29829);
   U25834 : XOR2_X1 port map( A1 => n19308, A2 => n28860, Z => n15384);
   U25835 : INV_X2 port map( I => n15386, ZN => n17217);
   U25836 : INV_X1 port map( I => n8585, ZN => n26477);
   U25837 : XOR2_X1 port map( A1 => Plaintext(76), A2 => Key(76), Z => n18542);
   U25838 : INV_X2 port map( I => n25544, ZN => n16933);
   U25841 : XOR2_X1 port map( A1 => n28914, A2 => n15394, Z => n15393);
   U25842 : XOR2_X1 port map( A1 => n13852, A2 => n15395, Z => n15394);
   U25845 : XOR2_X1 port map( A1 => n27683, A2 => n1356, Z => n15398);
   U25851 : XOR2_X1 port map( A1 => n39116, A2 => n19929, Z => n18604);
   U25852 : XOR2_X1 port map( A1 => n36750, A2 => n19729, Z => n22278);
   U25853 : INV_X2 port map( I => n15412, ZN => n22935);
   U25862 : INV_X1 port map( I => n18880, ZN => n19171);
   U25867 : NAND2_X1 port map( A1 => n22277, A2 => n9616, ZN => n15436);
   U25869 : XOR2_X1 port map( A1 => n38896, A2 => n37024, Z => n15442);
   U25873 : XOR2_X1 port map( A1 => n15450, A2 => n15451, Z => n16062);
   U25878 : INV_X2 port map( I => n15463, ZN => n23163);
   U25880 : NOR2_X1 port map( A1 => n24602, A2 => n34011, ZN => n17270);
   U25885 : XOR2_X1 port map( A1 => n5841, A2 => n15679, Z => n20486);
   U25887 : XOR2_X1 port map( A1 => n15476, A2 => n24078, Z => n20270);
   U25888 : XOR2_X1 port map( A1 => n24079, A2 => n15477, Z => n15476);
   U25891 : XOR2_X1 port map( A1 => n35222, A2 => n1724, Z => n15481);
   U25892 : XOR2_X1 port map( A1 => n26548, A2 => n29003, Z => n25985);
   U25893 : XOR2_X1 port map( A1 => n26548, A2 => n19081, Z => n18808);
   U25894 : XOR2_X1 port map( A1 => n20956, A2 => n26548, Z => n15529);
   U25898 : XOR2_X1 port map( A1 => n9757, A2 => n19732, Z => n15500);
   U25899 : NOR2_X1 port map( A1 => n37200, A2 => n918, ZN => n21524);
   U25900 : INV_X2 port map( I => n20591, ZN => n20590);
   U25902 : XOR2_X1 port map( A1 => n23843, A2 => n15507, Z => n24106);
   U25903 : XOR2_X1 port map( A1 => n14454, A2 => n23839, Z => n15507);
   U25904 : XOR2_X1 port map( A1 => n26489, A2 => n1727, Z => n15508);
   U25906 : INV_X2 port map( I => n19928, ZN => n15515);
   U25908 : NAND2_X2 port map( A1 => n19701, A2 => n15515, ZN => n25528);
   U25910 : OAI21_X1 port map( A1 => n15357, A2 => n31832, B => n15518, ZN => 
                           n28008);
   U25911 : MUX2_X1 port map( I0 => n36850, I1 => n29864, S => n29938, Z => 
                           n29866);
   U25912 : INV_X1 port map( I => n18115, ZN => n25019);
   U25916 : XOR2_X1 port map( A1 => n22495, A2 => n16199, Z => n18416);
   U25918 : XOR2_X1 port map( A1 => n20452, A2 => n29025, Z => n28780);
   U25919 : XOR2_X1 port map( A1 => n38844, A2 => n19624, Z => n26059);
   U25920 : XOR2_X1 port map( A1 => n38844, A2 => n1361, Z => n18322);
   U25921 : XOR2_X1 port map( A1 => n11667, A2 => n38844, Z => n26557);
   U25922 : XOR2_X1 port map( A1 => n27688, A2 => n15546, Z => n15545);
   U25923 : XOR2_X1 port map( A1 => n15547, A2 => n27689, Z => n15546);
   U25927 : XOR2_X1 port map( A1 => n25236, A2 => n25235, Z => n19644);
   U25928 : XOR2_X1 port map( A1 => n25323, A2 => n25160, Z => n25232);
   U25932 : XOR2_X1 port map( A1 => n39739, A2 => n38181, Z => n15565);
   U25934 : NAND2_X1 port map( A1 => n39112, A2 => n28228, ZN => n15572);
   U25936 : XOR2_X1 port map( A1 => n33511, A2 => n21294, Z => n20811);
   U25937 : XOR2_X1 port map( A1 => n33511, A2 => n19738, Z => n28870);
   U25939 : XOR2_X1 port map( A1 => n22542, A2 => n19738, Z => n18888);
   U25940 : XOR2_X1 port map( A1 => n15591, A2 => n7602, Z => n26073);
   U25943 : INV_X2 port map( I => n15598, ZN => n20896);
   U25944 : XOR2_X1 port map( A1 => n15600, A2 => n15599, Z => Ciphertext(2));
   U25946 : XOR2_X1 port map( A1 => n22624, A2 => n30179, Z => n15607);
   U25949 : NOR2_X1 port map( A1 => n30184, A2 => n30178, ZN => n15615);
   U25950 : NOR2_X2 port map( A1 => n15684, A2 => n15685, ZN => n15616);
   U25956 : XOR2_X1 port map( A1 => n23779, A2 => n37842, Z => n23691);
   U25961 : NAND2_X1 port map( A1 => n9394, A2 => n15651, ZN => n29201);
   U25966 : XOR2_X1 port map( A1 => n22743, A2 => n15654, Z => n15653);
   U25967 : XOR2_X1 port map( A1 => n33323, A2 => n19760, Z => n15654);
   U25969 : XOR2_X1 port map( A1 => n26587, A2 => n33735, Z => n15656);
   U25971 : XOR2_X1 port map( A1 => n34469, A2 => n30094, Z => n15660);
   U25973 : NAND3_X1 port map( A1 => n24804, A2 => n15664, A3 => n14064, ZN => 
                           n15689);
   U25974 : MUX2_X1 port map( I0 => n34354, I1 => n15664, S => n36471, Z => 
                           n24573);
   U25976 : AOI21_X1 port map( A1 => n28323, A2 => n13601, B => n3845, ZN => 
                           n28060);
   U25977 : XOR2_X1 port map( A1 => n15674, A2 => n15672, Z => n20063);
   U25979 : XOR2_X1 port map( A1 => n26595, A2 => n26594, Z => n15673);
   U25982 : XOR2_X1 port map( A1 => n24030, A2 => n15679, Z => n23681);
   U25983 : XOR2_X1 port map( A1 => n35936, A2 => n15679, Z => n23562);
   U25984 : NAND2_X2 port map( A1 => n23557, A2 => n23558, ZN => n15679);
   U25986 : AOI21_X2 port map( A1 => n23363, A2 => n23364, B => n15681, ZN => 
                           n24040);
   U25989 : OAI22_X2 port map( A1 => n18025, A2 => n17923, B1 => n21607, B2 => 
                           n18026, ZN => n15697);
   U25991 : XOR2_X1 port map( A1 => Plaintext(147), A2 => Key(147), Z => n21933
                           );
   U25994 : AOI21_X2 port map( A1 => n28083, A2 => n986, B => n28082, ZN => 
                           n28638);
   U26001 : XOR2_X1 port map( A1 => n27794, A2 => n16618, Z => n15721);
   U26002 : XOR2_X1 port map( A1 => n35303, A2 => n27754, Z => n15722);
   U26004 : XOR2_X1 port map( A1 => n27498, A2 => n27850, Z => n27795);
   U26009 : XOR2_X1 port map( A1 => n23662, A2 => n15729, Z => n15728);
   U26010 : XOR2_X1 port map( A1 => n23888, A2 => n19624, Z => n15729);
   U26011 : XOR2_X1 port map( A1 => n12570, A2 => n24028, Z => n15730);
   U26012 : XOR2_X1 port map( A1 => n22588, A2 => n17078, Z => n22525);
   U26014 : INV_X2 port map( I => n15839, ZN => n21579);
   U26015 : NOR3_X1 port map( A1 => n31530, A2 => n35137, A3 => n9197, ZN => 
                           n15735);
   U26017 : NOR2_X1 port map( A1 => n23174, A2 => n14130, ZN => n15739);
   U26020 : XOR2_X1 port map( A1 => n18242, A2 => n15745, Z => n29251);
   U26022 : NAND3_X1 port map( A1 => n1139, A2 => n17511, A3 => n34558, ZN => 
                           n16098);
   U26023 : NOR2_X1 port map( A1 => n16094, A2 => n34558, ZN => n20661);
   U26024 : XOR2_X1 port map( A1 => n38816, A2 => n19561, Z => n27550);
   U26026 : XOR2_X1 port map( A1 => n10221, A2 => n29934, Z => n15750);
   U26028 : XOR2_X1 port map( A1 => n27707, A2 => n36894, Z => n27816);
   U26029 : XOR2_X1 port map( A1 => n27524, A2 => n27522, Z => n15757);
   U26030 : XOR2_X1 port map( A1 => n15758, A2 => n30435, Z => n19198);
   U26033 : XOR2_X1 port map( A1 => n22763, A2 => n35211, Z => n15762);
   U26036 : NOR2_X1 port map( A1 => n26135, A2 => n36798, ZN => n15767);
   U26037 : INV_X1 port map( I => n15768, ZN => n29355);
   U26040 : INV_X2 port map( I => n16339, ZN => n16461);
   U26041 : NAND2_X1 port map( A1 => n7975, A2 => n7974, ZN => n19276);
   U26042 : NAND2_X1 port map( A1 => n7973, A2 => n7975, ZN => n27028);
   U26043 : NOR2_X1 port map( A1 => n26870, A2 => n7975, ZN => n26871);
   U26044 : XOR2_X1 port map( A1 => n26435, A2 => n38279, Z => n18975);
   U26046 : NAND2_X1 port map( A1 => n15773, A2 => n29883, ZN => n29876);
   U26047 : XOR2_X1 port map( A1 => n27799, A2 => n15776, Z => n27800);
   U26048 : XOR2_X1 port map( A1 => n15776, A2 => n19851, Z => n18539);
   U26054 : XOR2_X1 port map( A1 => n29159, A2 => n21172, Z => n15782);
   U26059 : AOI21_X1 port map( A1 => n28654, A2 => n28617, B => n15792, ZN => 
                           n28562);
   U26062 : NAND2_X1 port map( A1 => n17967, A2 => n39627, ZN => n15804);
   U26063 : NAND2_X2 port map( A1 => n15806, A2 => n15805, ZN => n22160);
   U26064 : NAND2_X1 port map( A1 => n21663, A2 => n21662, ZN => n15806);
   U26065 : XOR2_X1 port map( A1 => n15810, A2 => n15809, Z => n15808);
   U26066 : XOR2_X1 port map( A1 => n29050, A2 => n19820, Z => n15809);
   U26068 : XOR2_X1 port map( A1 => n21142, A2 => n15819, Z => n15818);
   U26075 : XOR2_X1 port map( A1 => n9719, A2 => n33990, Z => n15824);
   U26079 : XOR2_X1 port map( A1 => n18242, A2 => n19677, Z => n15835);
   U26086 : XOR2_X1 port map( A1 => n29253, A2 => n29238, Z => n29161);
   U26088 : NAND2_X1 port map( A1 => n22354, A2 => n22353, ZN => n16266);
   U26090 : INV_X1 port map( I => n16658, ZN => n16656);
   U26091 : NOR3_X1 port map( A1 => n31542, A2 => n35203, A3 => n1187, ZN => 
                           n18472);
   U26092 : OAI21_X1 port map( A1 => n17942, A2 => n1670, B => n22676, ZN => 
                           n17340);
   U26097 : NAND2_X1 port map( A1 => n12537, A2 => n28340, ZN => n28341);
   U26098 : OAI21_X1 port map( A1 => n19657, A2 => n27866, B => n16476, ZN => 
                           n28195);
   U26101 : NOR2_X1 port map( A1 => n29704, A2 => n29635, ZN => n20433);
   U26108 : NAND2_X1 port map( A1 => n19404, A2 => n9993, ZN => n18494);
   U26111 : OAI21_X1 port map( A1 => n18408, A2 => n22274, B => n35771, ZN => 
                           n16351);
   U26114 : NAND2_X1 port map( A1 => n7265, A2 => n39160, ZN => n25368);
   U26115 : NAND2_X1 port map( A1 => n7644, A2 => n32024, ZN => n16726);
   U26123 : NOR2_X1 port map( A1 => n26089, A2 => n9743, ZN => n17439);
   U26125 : NAND2_X1 port map( A1 => n20348, A2 => n1351, ZN => n17483);
   U26129 : AOI21_X1 port map( A1 => n1679, A2 => n22316, B => n9824, ZN => 
                           n22320);
   U26130 : OAI21_X1 port map( A1 => n14422, A2 => n14400, B => n29446, ZN => 
                           n17089);
   U26140 : NOR2_X1 port map( A1 => n37089, A2 => n22243, ZN => n22244);
   U26141 : NOR2_X1 port map( A1 => n19084, A2 => n16128, ZN => n16130);
   U26151 : INV_X1 port map( I => n10747, ZN => n18479);
   U26153 : INV_X1 port map( I => n18806, ZN => n19508);
   U26156 : INV_X1 port map( I => n8473, ZN => n18623);
   U26163 : NAND2_X1 port map( A1 => n28193, A2 => n27866, ZN => n16476);
   U26166 : INV_X1 port map( I => Key(94), ZN => n15838);
   U26170 : XOR2_X1 port map( A1 => n38147, A2 => n34239, Z => n21157);
   U26171 : XOR2_X1 port map( A1 => n38147, A2 => n29554, Z => n28502);
   U26172 : NAND2_X1 port map( A1 => n15841, A2 => n29439, ZN => n15840);
   U26173 : OAI22_X1 port map( A1 => n18495, A2 => n15841, B1 => n29435, B2 => 
                           n29434, ZN => n19689);
   U26180 : XOR2_X1 port map( A1 => n25174, A2 => n15858, Z => n15857);
   U26181 : XOR2_X1 port map( A1 => n25155, A2 => n19952, Z => n15858);
   U26182 : XOR2_X1 port map( A1 => n15862, A2 => n15861, Z => n15859);
   U26183 : XOR2_X1 port map( A1 => n23671, A2 => n12972, Z => n15861);
   U26186 : INV_X1 port map( I => n15867, ZN => n21011);
   U26187 : NOR2_X1 port map( A1 => n15867, A2 => n29792, ZN => n29783);
   U26188 : MUX2_X1 port map( I0 => n15867, I1 => n18257, S => n29792, Z => 
                           n29790);
   U26189 : OAI21_X1 port map( A1 => n29782, A2 => n15867, B => n29789, ZN => 
                           n21013);
   U26193 : NAND2_X1 port map( A1 => n31412, A2 => n15868, ZN => n17972);
   U26194 : NAND2_X2 port map( A1 => n23859, A2 => n23858, ZN => n25269);
   U26200 : MUX2_X1 port map( I0 => n24490, I1 => n15878, S => n9212, Z => 
                           n15877);
   U26204 : NAND2_X1 port map( A1 => n16302, A2 => n33280, ZN => n15891);
   U26206 : XNOR2_X1 port map( A1 => n20550, A2 => n15893, ZN => n15892);
   U26207 : XOR2_X1 port map( A1 => n20777, A2 => n15894, Z => n15893);
   U26208 : XOR2_X1 port map( A1 => n3917, A2 => n36065, Z => n15894);
   U26210 : INV_X2 port map( I => n15903, ZN => n24296);
   U26211 : AOI22_X2 port map( A1 => n34547, A2 => n24296, B1 => n13453, B2 => 
                           n33939, ZN => n24209);
   U26214 : XOR2_X1 port map( A1 => n24038, A2 => n23893, Z => n24006);
   U26217 : INV_X2 port map( I => n15913, ZN => n26802);
   U26222 : XOR2_X1 port map( A1 => n15916, A2 => n19775, Z => n16244);
   U26223 : XOR2_X1 port map( A1 => n35245, A2 => n29334, Z => n20678);
   U26232 : NAND3_X1 port map( A1 => n37040, A2 => n27416, A3 => n33773, ZN => 
                           n18640);
   U26233 : XOR2_X1 port map( A1 => n1468, A2 => n27802, Z => n15932);
   U26240 : XOR2_X1 port map( A1 => n32354, A2 => n34017, Z => n17721);
   U26242 : XOR2_X1 port map( A1 => n20082, A2 => n26392, Z => n16440);
   U26249 : XOR2_X1 port map( A1 => n18482, A2 => n23847, Z => n15987);
   U26250 : XOR2_X1 port map( A1 => n15989, A2 => n16775, Z => n25392);
   U26257 : OAI21_X2 port map( A1 => n17683, A2 => n17682, B => n16996, ZN => 
                           n29719);
   U26259 : MUX2_X1 port map( I0 => n23036, I1 => n23037, S => n1145, Z => 
                           n16007);
   U26261 : XOR2_X1 port map( A1 => n29037, A2 => n28589, Z => n16010);
   U26266 : XOR2_X1 port map( A1 => n23967, A2 => n39073, Z => n23790);
   U26268 : XOR2_X1 port map( A1 => n16022, A2 => n5116, Z => n16021);
   U26269 : XOR2_X1 port map( A1 => n23623, A2 => n1724, Z => n16022);
   U26271 : XOR2_X1 port map( A1 => n30612, A2 => n18432, Z => n16029);
   U26272 : XOR2_X1 port map( A1 => n23892, A2 => n16030, Z => n23773);
   U26274 : XOR2_X1 port map( A1 => n18006, A2 => n23655, Z => n23892);
   U26275 : NAND2_X1 port map( A1 => n16034, A2 => n14596, ZN => n28113);
   U26281 : XOR2_X1 port map( A1 => n38753, A2 => n20206, Z => n16046);
   U26283 : XOR2_X1 port map( A1 => n16054, A2 => n15960, Z => n28579);
   U26289 : NAND2_X2 port map( A1 => n16075, A2 => n30002, ZN => n30022);
   U26292 : NAND2_X1 port map( A1 => n25641, A2 => n38963, ZN => n16095);
   U26293 : OR2_X1 port map( A1 => n19713, A2 => n24874, Z => n16097);
   U26295 : XOR2_X1 port map( A1 => n18362, A2 => n29363, Z => n18363);
   U26296 : NOR2_X1 port map( A1 => n27030, A2 => n2522, ZN => n27033);
   U26297 : XOR2_X1 port map( A1 => n27692, A2 => n772, Z => n16103);
   U26302 : XOR2_X1 port map( A1 => n22758, A2 => n22419, Z => n22420);
   U26303 : XOR2_X1 port map( A1 => n29093, A2 => n29092, Z => n18127);
   U26309 : XOR2_X1 port map( A1 => n33916, A2 => n16332, Z => n16131);
   U26310 : XOR2_X1 port map( A1 => n16135, A2 => n25023, Z => n16134);
   U26311 : XOR2_X1 port map( A1 => n31112, A2 => n25165, Z => n16135);
   U26317 : XOR2_X1 port map( A1 => n16151, A2 => n16150, Z => n16149);
   U26318 : XOR2_X1 port map( A1 => n38880, A2 => n1622, Z => n16151);
   U26322 : XOR2_X1 port map( A1 => n16864, A2 => n1718, Z => n24575);
   U26325 : XOR2_X1 port map( A1 => n39575, A2 => n19883, Z => n16175);
   U26328 : INV_X1 port map( I => n16182, ZN => n23361);
   U26329 : NOR2_X1 port map( A1 => n16182, A2 => n23482, ZN => n22513);
   U26330 : XOR2_X1 port map( A1 => n35266, A2 => n29357, Z => n27555);
   U26336 : XOR2_X1 port map( A1 => n39756, A2 => n25193, Z => n16192);
   U26337 : XOR2_X1 port map( A1 => n16193, A2 => n16694, Z => n19838);
   U26340 : OAI21_X2 port map( A1 => n22851, A2 => n22861, B => n16202, ZN => 
                           n23352);
   U26341 : NAND2_X1 port map( A1 => n24072, A2 => n21310, ZN => n24083);
   U26343 : NOR2_X1 port map( A1 => n16209, A2 => n4849, ZN => n28375);
   U26344 : NOR2_X1 port map( A1 => n19994, A2 => n16209, ZN => n17682);
   U26347 : AND2_X1 port map( A1 => n13393, A2 => n26763, Z => n16221);
   U26349 : XOR2_X1 port map( A1 => n28913, A2 => n16705, Z => n16225);
   U26350 : XOR2_X1 port map( A1 => n26602, A2 => n30010, Z => n20261);
   U26351 : XOR2_X1 port map( A1 => n26602, A2 => n29320, Z => n26143);
   U26352 : XOR2_X1 port map( A1 => n26602, A2 => n19020, Z => n19019);
   U26353 : XOR2_X1 port map( A1 => n17798, A2 => n26602, Z => n17797);
   U26354 : INV_X1 port map( I => n16233, ZN => n17975);
   U26355 : NAND2_X1 port map( A1 => n29276, A2 => n16233, ZN => n29281);
   U26356 : XOR2_X1 port map( A1 => n35190, A2 => n19908, Z => n16269);
   U26357 : XOR2_X1 port map( A1 => n35189, A2 => n1697, Z => n20263);
   U26360 : XOR2_X1 port map( A1 => n26157, A2 => n20213, Z => n26434);
   U26361 : XOR2_X1 port map( A1 => n16249, A2 => n17705, Z => Ciphertext(12));
   U26362 : XOR2_X1 port map( A1 => n23764, A2 => n30063, Z => n16257);
   U26363 : XOR2_X1 port map( A1 => n31247, A2 => n32973, Z => n16258);
   U26365 : OAI21_X1 port map( A1 => n35272, A2 => n16260, B => n9790, ZN => 
                           n29406);
   U26366 : OAI21_X1 port map( A1 => n20724, A2 => n16260, B => n35272, ZN => 
                           n29392);
   U26368 : XOR2_X1 port map( A1 => n27630, A2 => n16269, Z => n16268);
   U26369 : XOR2_X1 port map( A1 => Plaintext(105), A2 => Key(105), Z => n18757
                           );
   U26370 : INV_X2 port map( I => n16356, ZN => n29828);
   U26375 : NAND3_X1 port map( A1 => n21067, A2 => n21066, A3 => n19933, ZN => 
                           n16291);
   U26376 : INV_X1 port map( I => n16293, ZN => n16292);
   U26377 : AOI21_X1 port map( A1 => n21067, A2 => n21066, B => n19933, ZN => 
                           n16293);
   U26378 : INV_X1 port map( I => n23885, ZN => n23964);
   U26379 : INV_X2 port map( I => n18741, ZN => n18870);
   U26380 : XOR2_X1 port map( A1 => n25275, A2 => n29141, Z => n24921);
   U26382 : XOR2_X1 port map( A1 => n16342, A2 => n34945, Z => n23465);
   U26383 : NOR2_X1 port map( A1 => n28754, A2 => n16303, ZN => n17007);
   U26386 : NAND3_X1 port map( A1 => n39656, A2 => n19549, A3 => n16305, ZN => 
                           n22116);
   U26392 : NAND2_X1 port map( A1 => n1405, A2 => n16328, ZN => n16874);
   U26393 : AOI21_X1 port map( A1 => n1405, A2 => n30043, B => n16328, ZN => 
                           n29952);
   U26394 : XOR2_X1 port map( A1 => n29072, A2 => n28972, Z => n28319);
   U26398 : XOR2_X1 port map( A1 => Key(103), A2 => Plaintext(103), Z => n16333
                           );
   U26401 : XOR2_X1 port map( A1 => n23758, A2 => n16338, Z => n16337);
   U26403 : NAND2_X1 port map( A1 => n26090, A2 => n19889, ZN => n18003);
   U26406 : XOR2_X1 port map( A1 => n973, A2 => n16357, Z => n17452);
   U26407 : XOR2_X1 port map( A1 => n25326, A2 => n16350, Z => n20151);
   U26408 : XOR2_X1 port map( A1 => n25093, A2 => n24922, Z => n25326);
   U26409 : XOR2_X1 port map( A1 => n29082, A2 => n20329, Z => n16358);
   U26411 : XOR2_X1 port map( A1 => n27690, A2 => n27736, Z => n16362);
   U26414 : XOR2_X1 port map( A1 => n32863, A2 => n19629, Z => n22745);
   U26415 : XOR2_X1 port map( A1 => n22643, A2 => n32863, Z => n22387);
   U26420 : XOR2_X1 port map( A1 => n16379, A2 => n28945, Z => n16378);
   U26421 : XOR2_X1 port map( A1 => n28927, A2 => n29081, Z => n16379);
   U26422 : XOR2_X1 port map( A1 => n26395, A2 => n14675, Z => n16381);
   U26423 : NAND2_X2 port map( A1 => n16390, A2 => n16389, ZN => n29720);
   U26424 : NOR2_X1 port map( A1 => n29700, A2 => n29699, ZN => n16391);
   U26426 : XOR2_X1 port map( A1 => n33916, A2 => n29838, Z => n16679);
   U26429 : NAND2_X1 port map( A1 => n28153, A2 => n28151, ZN => n16412);
   U26430 : XOR2_X1 port map( A1 => n1262, A2 => n19722, Z => n16417);
   U26431 : INV_X1 port map( I => n25149, ZN => n16422);
   U26432 : XOR2_X1 port map( A1 => n16424, A2 => n17051, Z => n16423);
   U26433 : XOR2_X1 port map( A1 => n26487, A2 => n26407, Z => n25841);
   U26436 : XOR2_X1 port map( A1 => n17349, A2 => n19897, Z => n16439);
   U26439 : AOI21_X1 port map( A1 => n16455, A2 => n22205, B => n21288, ZN => 
                           n16454);
   U26442 : XOR2_X1 port map( A1 => n16460, A2 => n19676, Z => n25331);
   U26443 : XOR2_X1 port map( A1 => n16460, A2 => n25194, Z => n17258);
   U26445 : XOR2_X1 port map( A1 => n16469, A2 => n30094, Z => Ciphertext(154))
                           ;
   U26446 : NOR2_X1 port map( A1 => n30097, A2 => n30096, ZN => n16470);
   U26450 : OR2_X1 port map( A1 => n35903, A2 => n26031, Z => n16478);
   U26451 : INV_X1 port map( I => n25615, ZN => n25617);
   U26454 : XOR2_X1 port map( A1 => n16492, A2 => n25298, Z => n25300);
   U26456 : XNOR2_X1 port map( A1 => Plaintext(28), A2 => Key(28), ZN => n16496
                           );
   U26457 : XOR2_X1 port map( A1 => n26404, A2 => n16498, Z => n16497);
   U26458 : INV_X1 port map( I => n17716, ZN => n26028);
   U26464 : NOR2_X1 port map( A1 => n14453, A2 => n26945, ZN => n16522);
   U26465 : XOR2_X1 port map( A1 => n29104, A2 => n29661, Z => n16529);
   U26469 : INV_X1 port map( I => n32637, ZN => n24810);
   U26471 : XOR2_X1 port map( A1 => n1460, A2 => n35178, Z => n16549);
   U26472 : XOR2_X1 port map( A1 => n27850, A2 => n29671, Z => n16550);
   U26474 : XOR2_X1 port map( A1 => n26225, A2 => n16557, Z => n16556);
   U26475 : XOR2_X1 port map( A1 => n12838, A2 => n10904, Z => n16557);
   U26477 : XOR2_X1 port map( A1 => n22508, A2 => n22645, Z => n22486);
   U26481 : XOR2_X1 port map( A1 => n22713, A2 => n16561, Z => n16560);
   U26482 : XOR2_X1 port map( A1 => n1323, A2 => n16562, Z => n16561);
   U26483 : XOR2_X1 port map( A1 => n22712, A2 => n21201, Z => n16563);
   U26485 : XOR2_X1 port map( A1 => n16743, A2 => n19722, Z => n16565);
   U26486 : XOR2_X1 port map( A1 => n22503, A2 => n16667, Z => n22569);
   U26488 : NAND2_X1 port map( A1 => n24394, A2 => n16449, ZN => n17947);
   U26490 : XOR2_X1 port map( A1 => n16584, A2 => n16582, Z => n28436);
   U26491 : XOR2_X1 port map( A1 => n28545, A2 => n16583, Z => n16582);
   U26495 : XOR2_X1 port map( A1 => n26404, A2 => n19763, Z => n16591);
   U26500 : NOR2_X1 port map( A1 => n1390, A2 => n19297, ZN => n16598);
   U26509 : XOR2_X1 port map( A1 => n38208, A2 => n30101, Z => n24067);
   U26510 : NAND2_X1 port map( A1 => n29708, A2 => n16629, ZN => n16628);
   U26511 : NAND2_X1 port map( A1 => n35771, A2 => n16635, ZN => n16634);
   U26512 : XOR2_X1 port map( A1 => n16639, A2 => n16640, Z => n16976);
   U26514 : NAND2_X1 port map( A1 => n35761, A2 => n33580, ZN => n16645);
   U26515 : XOR2_X1 port map( A1 => n22511, A2 => n1369, Z => n16648);
   U26516 : INV_X2 port map( I => n38901, ZN => n26972);
   U26518 : XOR2_X1 port map( A1 => n22594, A2 => n19775, Z => n16651);
   U26520 : NOR2_X1 port map( A1 => n35151, A2 => n39015, ZN => n20884);
   U26522 : XOR2_X1 port map( A1 => n26525, A2 => n1503, Z => n16665);
   U26523 : AOI21_X1 port map( A1 => n21012, A2 => n16682, B => n21011, ZN => 
                           n21010);
   U26526 : XOR2_X1 port map( A1 => n29254, A2 => n19736, Z => n16685);
   U26527 : XOR2_X1 port map( A1 => n22760, A2 => n16688, Z => n16687);
   U26528 : XOR2_X1 port map( A1 => n22761, A2 => n30068, Z => n16688);
   U26529 : XOR2_X1 port map( A1 => n22759, A2 => n16690, Z => n16689);
   U26531 : XOR2_X1 port map( A1 => n16695, A2 => n28887, Z => n16694);
   U26532 : XOR2_X1 port map( A1 => n23787, A2 => n17150, Z => n16698);
   U26534 : XOR2_X1 port map( A1 => n29093, A2 => n19674, Z => n16705);
   U26537 : NAND2_X1 port map( A1 => n19837, A2 => n16265, ZN => n18163);
   U26538 : NAND3_X1 port map( A1 => n22351, A2 => n19837, A3 => n35060, ZN => 
                           n22012);
   U26541 : XOR2_X1 port map( A1 => n16720, A2 => n1703, Z => Ciphertext(156));
   U26542 : OAI21_X1 port map( A1 => n30100, A2 => n10118, B => n30112, ZN => 
                           n16723);
   U26547 : XOR2_X1 port map( A1 => n4828, A2 => n29363, Z => n16735);
   U26549 : XOR2_X1 port map( A1 => n29064, A2 => n16741, Z => n16740);
   U26550 : XOR2_X1 port map( A1 => n19571, A2 => n29666, Z => n16741);
   U26551 : XOR2_X1 port map( A1 => n29066, A2 => n29065, Z => n16742);
   U26552 : XOR2_X1 port map( A1 => n16743, A2 => n19933, Z => n27695);
   U26559 : XOR2_X1 port map( A1 => n27534, A2 => n19814, Z => n16759);
   U26562 : XOR2_X1 port map( A1 => n12221, A2 => n26460, Z => n17487);
   U26564 : XOR2_X1 port map( A1 => n23869, A2 => n23699, Z => n16766);
   U26568 : XOR2_X1 port map( A1 => n39575, A2 => n28968, Z => n23665);
   U26571 : XOR2_X1 port map( A1 => n16771, A2 => n20748, Z => n20560);
   U26572 : XOR2_X1 port map( A1 => n16771, A2 => n18700, Z => n29143);
   U26573 : XOR2_X1 port map( A1 => n16771, A2 => n36513, Z => n19445);
   U26574 : NOR2_X1 port map( A1 => n9066, A2 => n33939, ZN => n24149);
   U26575 : OAI21_X1 port map( A1 => n19914, A2 => n14458, B => n16773, ZN => 
                           n26137);
   U26576 : XOR2_X1 port map( A1 => n1505, A2 => n26476, Z => n16998);
   U26577 : XOR2_X1 port map( A1 => n38171, A2 => n19359, Z => n16776);
   U26578 : XOR2_X1 port map( A1 => n11974, A2 => n29718, Z => n16783);
   U26582 : XOR2_X1 port map( A1 => n32776, A2 => n19943, Z => n23683);
   U26584 : NAND3_X1 port map( A1 => n10618, A2 => n35777, A3 => n17771, ZN => 
                           n16791);
   U26585 : XNOR2_X1 port map( A1 => n16795, A2 => n16793, ZN => n16792);
   U26586 : XOR2_X1 port map( A1 => n16794, A2 => n16796, Z => n16793);
   U26587 : XOR2_X1 port map( A1 => n1618, A2 => n23910, Z => n16794);
   U26589 : XOR2_X1 port map( A1 => n23905, A2 => n29298, Z => n16796);
   U26590 : XOR2_X1 port map( A1 => n38208, A2 => n23686, Z => n16797);
   U26591 : NAND2_X1 port map( A1 => n22818, A2 => n1315, ZN => n20177);
   U26592 : XOR2_X1 port map( A1 => n16802, A2 => n16799, Z => n19685);
   U26593 : XOR2_X1 port map( A1 => n16801, A2 => n16800, Z => n16799);
   U26594 : XOR2_X1 port map( A1 => n22790, A2 => n29394, Z => n16800);
   U26595 : XOR2_X1 port map( A1 => n22789, A2 => n36290, Z => n16801);
   U26597 : NAND2_X2 port map( A1 => n17287, A2 => n17302, ZN => n16803);
   U26598 : XOR2_X1 port map( A1 => n900, A2 => n19839, Z => n16806);
   U26603 : NAND2_X2 port map( A1 => n25018, A2 => n18115, ZN => n24965);
   U26605 : NOR2_X1 port map( A1 => n38193, A2 => n39583, ZN => n18716);
   U26610 : NAND2_X1 port map( A1 => n496, A2 => n16853, ZN => n19391);
   U26611 : NAND2_X1 port map( A1 => n28733, A2 => n16853, ZN => n27553);
   U26612 : NAND2_X1 port map( A1 => n24782, A2 => n24779, ZN => n16855);
   U26619 : NOR2_X1 port map( A1 => n26186, A2 => n16878, ZN => n26188);
   U26624 : OR2_X1 port map( A1 => n34171, A2 => n2937, Z => n28297);
   U26625 : NAND2_X1 port map( A1 => n18671, A2 => n32790, ZN => n16985);
   U26629 : XOR2_X1 port map( A1 => n31320, A2 => n27704, Z => n16886);
   U26630 : NOR2_X1 port map( A1 => n1492, A2 => n19712, ZN => n26148);
   U26637 : NOR2_X1 port map( A1 => n25892, A2 => n15677, ZN => n16904);
   U26641 : NAND3_X1 port map( A1 => n24783, A2 => n1121, A3 => n38658, ZN => 
                           n24414);
   U26644 : XOR2_X1 port map( A1 => n18291, A2 => n22666, Z => n16912);
   U26647 : NAND2_X2 port map( A1 => n16929, A2 => n23427, ZN => n23955);
   U26649 : AOI21_X1 port map( A1 => n29431, A2 => n29435, B => n19618, ZN => 
                           n19617);
   U26655 : AND2_X1 port map( A1 => n19692, A2 => n22895, Z => n20344);
   U26659 : NAND3_X1 port map( A1 => n38210, A2 => n10004, A3 => n25609, ZN => 
                           n19257);
   U26660 : XOR2_X1 port map( A1 => n21408, A2 => Key(163), Z => n18739);
   U26662 : XOR2_X1 port map( A1 => n22663, A2 => n22662, Z => n21278);
   U26664 : OAI21_X1 port map( A1 => n29440, A2 => n29438, B => n16960, ZN => 
                           n17317);
   U26668 : NAND2_X2 port map( A1 => n25775, A2 => n25777, ZN => n18827);
   U26671 : XOR2_X1 port map( A1 => n28944, A2 => n16976, Z => n16975);
   U26676 : NAND2_X1 port map( A1 => n18908, A2 => n29682, ZN => n29688);
   U26677 : NOR2_X1 port map( A1 => n25468, A2 => n25606, ZN => n17480);
   U26678 : NAND2_X1 port map( A1 => n19796, A2 => n19795, ZN => n19794);
   U26679 : XOR2_X1 port map( A1 => n16992, A2 => n38265, Z => Ciphertext(129))
                           ;
   U26684 : OAI21_X1 port map( A1 => n12290, A2 => n26686, B => n852, ZN => 
                           n17099);
   U26686 : INV_X1 port map( I => n27875, ZN => n27998);
   U26687 : XOR2_X1 port map( A1 => n25211, A2 => n24886, Z => n25178);
   U26688 : INV_X1 port map( I => n23394, ZN => n22912);
   U26690 : XOR2_X1 port map( A1 => n25299, A2 => n25300, Z => n18869);
   U26691 : XNOR2_X1 port map( A1 => n26599, A2 => n19876, ZN => n17858);
   U26699 : NAND2_X1 port map( A1 => n29551, A2 => n29558, ZN => n28907);
   U26701 : NAND2_X2 port map( A1 => n25731, A2 => n25732, ZN => n17915);
   U26702 : XOR2_X1 port map( A1 => n17028, A2 => n14646, Z => n25613);
   U26703 : XOR2_X1 port map( A1 => n25091, A2 => n25092, Z => n17028);
   U26704 : XOR2_X1 port map( A1 => n17030, A2 => n29978, Z => Ciphertext(136))
                           ;
   U26705 : NOR2_X1 port map( A1 => n22904, A2 => n22813, ZN => n22903);
   U26709 : XOR2_X1 port map( A1 => n27856, A2 => n17033, Z => n27857);
   U26710 : XOR2_X1 port map( A1 => n27854, A2 => n27855, Z => n17033);
   U26719 : NOR2_X1 port map( A1 => n21604, A2 => n21783, ZN => n18340);
   U26725 : XOR2_X1 port map( A1 => n29553, A2 => n29554, Z => Ciphertext(64));
   U26726 : NAND3_X1 port map( A1 => n17152, A2 => n39305, A3 => n27263, ZN => 
                           n17151);
   U26729 : NAND2_X1 port map( A1 => n36191, A2 => n23450, ZN => n17470);
   U26731 : XOR2_X1 port map( A1 => n17063, A2 => n25736, Z => n26796);
   U26734 : XOR2_X1 port map( A1 => n29115, A2 => n29252, Z => n28574);
   U26738 : NAND2_X1 port map( A1 => n1268, A2 => n24900, ZN => n17377);
   U26739 : XOR2_X1 port map( A1 => n29165, A2 => n29614, Z => n28824);
   U26740 : OR2_X1 port map( A1 => n21958, A2 => n17086, Z => n21959);
   U26741 : NAND2_X1 port map( A1 => n19134, A2 => n19840, ZN => n21065);
   U26743 : OR2_X1 port map( A1 => n22340, A2 => n22341, Z => n21988);
   U26745 : XOR2_X1 port map( A1 => n25197, A2 => n25283, Z => n25060);
   U26751 : OAI21_X1 port map( A1 => n17382, A2 => n29662, B => n1390, ZN => 
                           n17381);
   U26752 : XOR2_X1 port map( A1 => n17113, A2 => n1702, Z => Ciphertext(71));
   U26761 : NAND2_X1 port map( A1 => n21997, A2 => n22265, ZN => n18401);
   U26762 : INV_X2 port map( I => n17119, ZN => n17127);
   U26765 : XOR2_X1 port map( A1 => n25039, A2 => n25041, Z => n17129);
   U26766 : XOR2_X1 port map( A1 => n7432, A2 => n30207, Z => n19201);
   U26767 : XOR2_X1 port map( A1 => n38330, A2 => n7432, Z => n20719);
   U26770 : NAND3_X1 port map( A1 => n25374, A2 => n25375, A3 => n35508, ZN => 
                           n25376);
   U26772 : XOR2_X1 port map( A1 => n26458, A2 => n38177, Z => n17136);
   U26774 : XOR2_X1 port map( A1 => n26572, A2 => n26277, Z => n17137);
   U26776 : XOR2_X1 port map( A1 => n10579, A2 => n20263, Z => n17139);
   U26777 : XOR2_X1 port map( A1 => n35707, A2 => n17705, Z => n17704);
   U26778 : INV_X1 port map( I => n27325, ZN => n27400);
   U26782 : NAND2_X1 port map( A1 => n1333, A2 => n22228, ZN => n17147);
   U26784 : XOR2_X1 port map( A1 => n23886, A2 => n19919, Z => n17150);
   U26785 : XOR2_X1 port map( A1 => n37094, A2 => n29371, Z => n17153);
   U26786 : XOR2_X1 port map( A1 => n22453, A2 => n11308, Z => n22550);
   U26787 : NAND2_X2 port map( A1 => n21658, A2 => n21657, ZN => n19655);
   U26791 : NAND2_X1 port map( A1 => n14418, A2 => n21779, ZN => n17160);
   U26793 : XOR2_X1 port map( A1 => n39129, A2 => n30104, Z => n25734);
   U26794 : XOR2_X1 port map( A1 => n39129, A2 => n19817, Z => n26323);
   U26795 : XOR2_X1 port map( A1 => n17171, A2 => n17172, Z => n20389);
   U26797 : XOR2_X1 port map( A1 => n26154, A2 => n26156, Z => n17172);
   U26801 : XOR2_X1 port map( A1 => n27731, A2 => n31551, Z => n18511);
   U26802 : XOR2_X1 port map( A1 => n19231, A2 => n14691, Z => n17177);
   U26803 : NOR2_X2 port map( A1 => n20369, A2 => n29631, ZN => n29662);
   U26805 : XOR2_X1 port map( A1 => n17189, A2 => n30010, Z => n22001);
   U26806 : XOR2_X1 port map( A1 => n17189, A2 => n29785, Z => n22568);
   U26809 : XOR2_X1 port map( A1 => Plaintext(126), A2 => Key(126), Z => n20703
                           );
   U26810 : INV_X2 port map( I => n31596, ZN => n20979);
   U26812 : INV_X2 port map( I => n17210, ZN => n20267);
   U26813 : OAI21_X1 port map( A1 => n17212, A2 => n1245, B => n17211, ZN => 
                           n17213);
   U26814 : NAND3_X1 port map( A1 => n28143, A2 => n28142, A3 => n17114, ZN => 
                           n28145);
   U26815 : INV_X2 port map( I => n19806, ZN => n24461);
   U26817 : NOR2_X1 port map( A1 => n29347, A2 => n29120, ZN => n20508);
   U26819 : NOR3_X1 port map( A1 => n17233, A2 => n1351, A3 => n19202, ZN => 
                           n17678);
   U26821 : XOR2_X1 port map( A1 => n7667, A2 => n35702, Z => n17245);
   U26823 : XOR2_X1 port map( A1 => n25097, A2 => n24924, Z => n18765);
   U26825 : NAND2_X1 port map( A1 => n17249, A2 => n6604, ZN => n21552);
   U26828 : NOR2_X1 port map( A1 => n18603, A2 => n34120, ZN => n17253);
   U26829 : XOR2_X1 port map( A1 => n17256, A2 => n17258, Z => n17255);
   U26830 : XOR2_X1 port map( A1 => n25250, A2 => n17257, Z => n17256);
   U26833 : NOR2_X1 port map( A1 => n30731, A2 => n19542, ZN => n17264);
   U26835 : XOR2_X1 port map( A1 => n35241, A2 => n27858, Z => n17272);
   U26836 : XOR2_X1 port map( A1 => n27362, A2 => n17274, Z => n17273);
   U26837 : XOR2_X1 port map( A1 => n27564, A2 => n17275, Z => n17274);
   U26838 : XOR2_X1 port map( A1 => n27724, A2 => n27516, Z => n27362);
   U26841 : NOR2_X1 port map( A1 => n20223, A2 => n26619, ZN => n17278);
   U26843 : NAND2_X1 port map( A1 => n19367, A2 => n17281, ZN => n25571);
   U26844 : XOR2_X1 port map( A1 => n22728, A2 => n36290, Z => n17283);
   U26845 : XOR2_X1 port map( A1 => n22729, A2 => n30006, Z => n17285);
   U26847 : XOR2_X1 port map( A1 => n17292, A2 => n24859, Z => n25106);
   U26848 : AOI21_X1 port map( A1 => n29435, A2 => n18502, B => n17293, ZN => 
                           n17318);
   U26850 : NOR2_X1 port map( A1 => n25454, A2 => n31375, ZN => n17297);
   U26855 : INV_X1 port map( I => n28696, ZN => n17322);
   U26857 : XOR2_X1 port map( A1 => n29303, A2 => n28889, Z => n17325);
   U26859 : XOR2_X1 port map( A1 => n31112, A2 => n30090, Z => n17328);
   U26863 : NAND2_X2 port map( A1 => n22312, A2 => n22311, ZN => n22453);
   U26865 : NAND2_X1 port map( A1 => n14590, A2 => n17357, ZN => n17356);
   U26866 : AOI21_X1 port map( A1 => n1675, A2 => n22228, B => n1333, ZN => 
                           n17357);
   U26867 : OR2_X1 port map( A1 => n22089, A2 => n17359, Z => n17358);
   U26869 : XOR2_X1 port map( A1 => n26484, A2 => n21100, Z => n17361);
   U26870 : XOR2_X1 port map( A1 => n17366, A2 => n34945, Z => Ciphertext(68));
   U26872 : OR2_X1 port map( A1 => n26114, A2 => n31624, Z => n17373);
   U26873 : AOI21_X1 port map( A1 => n29658, A2 => n17382, B => n17381, ZN => 
                           n20443);
   U26876 : XOR2_X1 port map( A1 => Plaintext(148), A2 => Key(148), Z => n18027
                           );
   U26877 : XOR2_X1 port map( A1 => n7402, A2 => n19905, Z => n20730);
   U26879 : OAI21_X1 port map( A1 => n28679, A2 => n33646, B => n28719, ZN => 
                           n19304);
   U26881 : XOR2_X1 port map( A1 => n17850, A2 => n1713, Z => n17404);
   U26882 : XOR2_X1 port map( A1 => n27471, A2 => n27472, Z => n17406);
   U26883 : XOR2_X1 port map( A1 => n27728, A2 => n14693, Z => n20693);
   U26885 : XOR2_X1 port map( A1 => n22776, A2 => n39787, Z => n17429);
   U26889 : NAND3_X1 port map( A1 => n32616, A2 => n31234, A3 => n34307, ZN => 
                           n23632);
   U26892 : NOR2_X1 port map( A1 => n20364, A2 => n5515, ZN => n20363);
   U26899 : NAND2_X1 port map( A1 => n20274, A2 => n17469, ZN => n29008);
   U26901 : NOR2_X1 port map( A1 => n24713, A2 => n24899, ZN => n17473);
   U26906 : XOR2_X1 port map( A1 => n17492, A2 => n17489, Z => n19949);
   U26907 : XOR2_X1 port map( A1 => n17491, A2 => n17490, Z => n17489);
   U26908 : XOR2_X1 port map( A1 => n23686, A2 => n29849, Z => n17490);
   U26909 : XOR2_X1 port map( A1 => n23952, A2 => n35942, Z => n17491);
   U26911 : XOR2_X1 port map( A1 => n28867, A2 => n20033, Z => n17494);
   U26914 : XOR2_X1 port map( A1 => n38370, A2 => n19905, Z => n23940);
   U26915 : XOR2_X1 port map( A1 => n39038, A2 => n29051, Z => n23960);
   U26916 : XOR2_X1 port map( A1 => n17518, A2 => n17517, Z => n17516);
   U26917 : XOR2_X1 port map( A1 => n17462, A2 => n19929, Z => n17517);
   U26918 : XOR2_X1 port map( A1 => n23961, A2 => n17520, Z => n17519);
   U26919 : XOR2_X1 port map( A1 => n24050, A2 => n23814, Z => n17520);
   U26920 : OAI21_X1 port map( A1 => n21110, A2 => n21109, B => n30169, ZN => 
                           n17523);
   U26921 : OR2_X1 port map( A1 => n21109, A2 => n30169, Z => n17524);
   U26922 : XOR2_X1 port map( A1 => n22750, A2 => n17528, Z => n20836);
   U26923 : XOR2_X1 port map( A1 => n21378, A2 => Key(67), Z => n19370);
   U26926 : NAND2_X2 port map( A1 => n21513, A2 => n21512, ZN => n22322);
   U26933 : XOR2_X1 port map( A1 => n10012, A2 => n19905, Z => n17552);
   U26934 : XOR2_X1 port map( A1 => n25234, A2 => n17555, Z => n17554);
   U26935 : INV_X1 port map( I => n35529, ZN => n20025);
   U26936 : XOR2_X1 port map( A1 => n35255, A2 => n29131, Z => n29133);
   U26940 : INV_X1 port map( I => n22448, ZN => n17566);
   U26941 : NAND2_X2 port map( A1 => n29193, A2 => n29192, ZN => n29740);
   U26943 : NAND2_X1 port map( A1 => n17989, A2 => n17499, ZN => n22050);
   U26944 : XOR2_X1 port map( A1 => n17580, A2 => n38880, Z => n17579);
   U26949 : XOR2_X1 port map( A1 => n39797, A2 => n30006, Z => n17595);
   U26950 : XOR2_X1 port map( A1 => n31163, A2 => n17603, Z => n20311);
   U26951 : INV_X2 port map( I => n17604, ZN => n25557);
   U26952 : XOR2_X1 port map( A1 => n35238, A2 => n39172, Z => n26167);
   U26959 : XOR2_X1 port map( A1 => n27466, A2 => n35241, Z => n17621);
   U26962 : NAND2_X2 port map( A1 => n28063, A2 => n28062, ZN => n29254);
   U26963 : XOR2_X1 port map( A1 => n28983, A2 => n19527, Z => n17627);
   U26965 : NAND2_X1 port map( A1 => n906, A2 => n20873, ZN => n17630);
   U26966 : NAND2_X1 port map( A1 => n17636, A2 => n1048, ZN => n17635);
   U26967 : XOR2_X1 port map( A1 => n28306, A2 => n17643, Z => n17642);
   U26971 : INV_X2 port map( I => n17660, ZN => n24287);
   U26973 : NOR2_X1 port map( A1 => n21780, A2 => n12144, ZN => n17679);
   U26978 : NAND3_X1 port map( A1 => n17687, A2 => n18986, A3 => n27465, ZN => 
                           n17699);
   U26981 : XOR2_X1 port map( A1 => Plaintext(129), A2 => Key(129), Z => n20300
                           );
   U26982 : XOR2_X1 port map( A1 => n24801, A2 => n17704, Z => n18556);
   U26983 : XOR2_X1 port map( A1 => n16627, A2 => n1557, Z => n17706);
   U26984 : XOR2_X1 port map( A1 => n24991, A2 => n19534, Z => n17707);
   U26985 : INV_X1 port map( I => Plaintext(146), ZN => n17717);
   U26986 : XOR2_X1 port map( A1 => n17717, A2 => Key(146), Z => n17799);
   U26988 : INV_X2 port map( I => n17726, ZN => n29781);
   U26990 : XOR2_X1 port map( A1 => n467, A2 => n17738, Z => n17737);
   U26991 : XOR2_X1 port map( A1 => n29040, A2 => n13639, Z => n17738);
   U26992 : AND2_X1 port map( A1 => n23550, A2 => n17094, Z => n17744);
   U26994 : XOR2_X1 port map( A1 => n17747, A2 => n29879, Z => Ciphertext(122))
                           ;
   U26996 : NAND2_X1 port map( A1 => n39019, A2 => n17286, ZN => n17750);
   U27001 : INV_X2 port map( I => n17764, ZN => n25558);
   U27002 : INV_X2 port map( I => n25558, ZN => n25719);
   U27003 : INV_X2 port map( I => n17767, ZN => n18841);
   U27007 : XOR2_X1 port map( A1 => n8833, A2 => n29801, Z => n21003);
   U27008 : XOR2_X1 port map( A1 => n17776, A2 => n19714, Z => n20526);
   U27015 : AOI21_X1 port map( A1 => n25799, A2 => n31263, B => n38168, ZN => 
                           n19048);
   U27019 : MUX2_X1 port map( I0 => n23221, I1 => n23222, S => n18236, Z => 
                           n23223);
   U27020 : XOR2_X1 port map( A1 => n27830, A2 => n27862, Z => n17817);
   U27022 : XOR2_X1 port map( A1 => n23707, A2 => n19755, Z => n19344);
   U27024 : INV_X2 port map( I => n17830, ZN => n23108);
   U27025 : OR2_X1 port map( A1 => n20493, A2 => n20492, Z => n17831);
   U27028 : XOR2_X1 port map( A1 => n17836, A2 => n17835, Z => n17839);
   U27029 : XOR2_X1 port map( A1 => n1261, A2 => n25104, Z => n17835);
   U27035 : XOR2_X1 port map( A1 => n17854, A2 => n17853, Z => n17852);
   U27036 : XOR2_X1 port map( A1 => n39682, A2 => n18700, Z => n17853);
   U27038 : XOR2_X1 port map( A1 => n29071, A2 => n20479, Z => n17859);
   U27039 : NOR2_X1 port map( A1 => n17864, A2 => n22240, ZN => n19180);
   U27040 : OAI21_X1 port map( A1 => n24449, A2 => n24453, B => n17867, ZN => 
                           n24246);
   U27045 : XOR2_X1 port map( A1 => n23922, A2 => n37521, Z => n17872);
   U27046 : OAI21_X1 port map( A1 => n18720, A2 => n29494, B => n29451, ZN => 
                           n28619);
   U27048 : XOR2_X1 port map( A1 => n38137, A2 => n19738, Z => n26339);
   U27051 : XOR2_X1 port map( A1 => n17910, A2 => n22764, Z => n17909);
   U27052 : INV_X2 port map( I => n19959, ZN => n17911);
   U27053 : NOR2_X1 port map( A1 => n24195, A2 => n17911, ZN => n20734);
   U27056 : XOR2_X1 port map( A1 => n17921, A2 => n26183, Z => n17920);
   U27058 : XOR2_X1 port map( A1 => n17937, A2 => n23898, Z => n23669);
   U27059 : XOR2_X1 port map( A1 => n17945, A2 => n17944, Z => n20573);
   U27060 : XOR2_X1 port map( A1 => n844, A2 => n838, Z => n17944);
   U27061 : XOR2_X1 port map( A1 => n26263, A2 => n17946, Z => n17945);
   U27062 : XNOR2_X1 port map( A1 => Plaintext(91), A2 => Key(91), ZN => n17964
                           );
   U27063 : XOR2_X1 port map( A1 => n17974, A2 => n19592, Z => Ciphertext(23));
   U27066 : NAND2_X1 port map( A1 => n29958, A2 => n29959, ZN => n17983);
   U27067 : XOR2_X1 port map( A1 => n1667, A2 => n39136, Z => n18912);
   U27070 : XOR2_X1 port map( A1 => n22509, A2 => n39787, Z => n17999);
   U27071 : AOI21_X1 port map( A1 => n993, A2 => n27137, B => n19477, ZN => 
                           n18074);
   U27072 : NOR2_X1 port map( A1 => n7304, A2 => n1348, ZN => n18005);
   U27073 : XOR2_X1 port map( A1 => n18006, A2 => n39636, Z => n18410);
   U27074 : XOR2_X1 port map( A1 => n18012, A2 => n30016, Z => n18367);
   U27075 : XOR2_X1 port map( A1 => n18012, A2 => n29285, Z => n26295);
   U27076 : XOR2_X1 port map( A1 => n25152, A2 => n18015, Z => n18014);
   U27081 : NAND3_X1 port map( A1 => n20672, A2 => n1173, A3 => n18042, ZN => 
                           n20862);
   U27082 : INV_X1 port map( I => n14387, ZN => n30215);
   U27085 : XOR2_X1 port map( A1 => n18931, A2 => n12707, Z => n18317);
   U27086 : NAND2_X1 port map( A1 => n28717, A2 => n32759, ZN => n28497);
   U27088 : OAI21_X1 port map( A1 => n26122, A2 => n31719, B => n25903, ZN => 
                           n25905);
   U27089 : XOR2_X1 port map( A1 => n27862, A2 => n29295, Z => n27680);
   U27090 : XOR2_X1 port map( A1 => n20602, A2 => n18078, Z => n20601);
   U27091 : XOR2_X1 port map( A1 => n18080, A2 => n18079, Z => n18078);
   U27092 : XOR2_X1 port map( A1 => n23707, A2 => n29661, Z => n18079);
   U27095 : OAI21_X1 port map( A1 => n18084, A2 => n18083, B => n39709, ZN => 
                           n18082);
   U27096 : AND2_X1 port map( A1 => n31570, A2 => n29927, Z => n18084);
   U27098 : NAND2_X1 port map( A1 => n18089, A2 => n18088, ZN => n28770);
   U27105 : AND2_X1 port map( A1 => n37674, A2 => n23155, Z => n23157);
   U27107 : XOR2_X1 port map( A1 => n24012, A2 => n18109, Z => n19623);
   U27113 : XOR2_X1 port map( A1 => n23955, A2 => n24012, Z => n23717);
   U27115 : XOR2_X1 port map( A1 => n1466, A2 => n1468, Z => n18122);
   U27117 : NOR3_X1 port map( A1 => n15338, A2 => n15839, A3 => n21571, ZN => 
                           n20580);
   U27125 : XOR2_X1 port map( A1 => n18137, A2 => n39482, Z => Ciphertext(27));
   U27134 : INV_X2 port map( I => n18156, ZN => n20404);
   U27136 : XOR2_X1 port map( A1 => Plaintext(5), A2 => Key(5), Z => n18157);
   U27139 : XOR2_X1 port map( A1 => Plaintext(63), A2 => Key(63), Z => n18722);
   U27140 : XNOR2_X1 port map( A1 => n23879, A2 => n24014, ZN => n18179);
   U27145 : XOR2_X1 port map( A1 => n23730, A2 => n18172, Z => n21316);
   U27147 : XOR2_X1 port map( A1 => n18404, A2 => n18403, Z => n18178);
   U27150 : INV_X2 port map( I => n18183, ZN => n26751);
   U27152 : XOR2_X1 port map( A1 => n18184, A2 => n29707, Z => Ciphertext(90));
   U27153 : OAI22_X1 port map( A1 => n29706, A2 => n29722, B1 => n29705, B2 => 
                           n29712, ZN => n18184);
   U27156 : NAND2_X1 port map( A1 => n18952, A2 => n18951, ZN => n18950);
   U27159 : NAND3_X2 port map( A1 => n22014, A2 => n22012, A3 => n22013, ZN => 
                           n22790);
   U27162 : NOR2_X1 port map( A1 => n19367, A2 => n25558, ZN => n19236);
   U27163 : XNOR2_X1 port map( A1 => n19983, A2 => n19984, ZN => n19714);
   U27164 : NAND2_X2 port map( A1 => n18208, A2 => n28903, ZN => n29548);
   U27165 : NAND3_X1 port map( A1 => n28902, A2 => n18720, A3 => n29491, ZN => 
                           n18208);
   U27170 : XOR2_X1 port map( A1 => n26403, A2 => n26407, Z => n25986);
   U27171 : AND2_X1 port map( A1 => n23484, A2 => n22493, Z => n20992);
   U27179 : OR2_X1 port map( A1 => n29682, A2 => n33128, Z => n18945);
   U27182 : XOR2_X1 port map( A1 => n18243, A2 => n1724, Z => Ciphertext(81));
   U27185 : XOR2_X1 port map( A1 => n22699, A2 => n22715, Z => n18255);
   U27189 : NOR2_X1 port map( A1 => n19347, A2 => n29717, ZN => n29706);
   U27190 : BUF_X2 port map( I => n21753, Z => n18266);
   U27191 : XOR2_X1 port map( A1 => n26366, A2 => n26398, Z => n18267);
   U27192 : NAND2_X1 port map( A1 => n21698, A2 => n19709, ZN => n19036);
   U27196 : OAI22_X1 port map( A1 => n27584, A2 => n27585, B1 => n31955, B2 => 
                           n27586, ZN => n27591);
   U27198 : XOR2_X1 port map( A1 => n5836, A2 => n22418, Z => n22421);
   U27201 : XNOR2_X1 port map( A1 => n24011, A2 => n29718, ZN => n20973);
   U27203 : XOR2_X1 port map( A1 => n29042, A2 => n38290, Z => n18319);
   U27205 : NAND2_X2 port map( A1 => n24438, A2 => n24437, ZN => n25290);
   U27207 : XOR2_X1 port map( A1 => n36886, A2 => n19152, Z => n22495);
   U27211 : NAND2_X1 port map( A1 => n29617, A2 => n29612, ZN => n18306);
   U27214 : OAI21_X1 port map( A1 => n30031, A2 => n30030, B => n18313, ZN => 
                           Ciphertext(142));
   U27219 : XOR2_X1 port map( A1 => n25166, A2 => n24697, Z => n18327);
   U27222 : XOR2_X1 port map( A1 => n26142, A2 => n17551, Z => n18335);
   U27226 : INV_X2 port map( I => n18345, ZN => n24465);
   U27228 : INV_X2 port map( I => n7705, ZN => n25647);
   U27231 : XOR2_X1 port map( A1 => n26508, A2 => n18367, Z => n18366);
   U27233 : NAND2_X1 port map( A1 => n13336, A2 => n12392, ZN => n18386);
   U27235 : NOR3_X1 port map( A1 => n39574, A2 => n28233, A3 => n18392, ZN => 
                           n27062);
   U27236 : NAND2_X1 port map( A1 => n24504, A2 => n6977, ZN => n18394);
   U27238 : NAND2_X2 port map( A1 => n25458, A2 => n25457, ZN => n26020);
   U27239 : XOR2_X1 port map( A1 => n23937, A2 => n23330, Z => n18403);
   U27240 : XOR2_X1 port map( A1 => n14638, A2 => n29299, Z => n18405);
   U27242 : XOR2_X1 port map( A1 => n23985, A2 => n18410, Z => n18427);
   U27243 : XOR2_X1 port map( A1 => n18422, A2 => n25044, Z => n18421);
   U27244 : XOR2_X1 port map( A1 => n13342, A2 => n24927, Z => n18422);
   U27245 : XOR2_X1 port map( A1 => n25043, A2 => n25042, Z => n18423);
   U27248 : INV_X2 port map( I => n24202, ZN => n18907);
   U27253 : XOR2_X1 port map( A1 => n27042, A2 => n760, Z => n18449);
   U27256 : XOR2_X1 port map( A1 => n39631, A2 => n28953, Z => n28954);
   U27259 : NAND2_X1 port map( A1 => n18484, A2 => n24229, ZN => n24230);
   U27260 : OAI21_X1 port map( A1 => n20133, A2 => n11820, B => n18488, ZN => 
                           n27185);
   U27263 : XOR2_X1 port map( A1 => n31941, A2 => n26541, Z => n26431);
   U27265 : XOR2_X1 port map( A1 => n18526, A2 => n28806, Z => n18491);
   U27267 : OAI21_X1 port map( A1 => n27951, A2 => n12303, B => n18497, ZN => 
                           n27868);
   U27272 : XOR2_X1 port map( A1 => n24930, A2 => n19742, Z => n25720);
   U27273 : XOR2_X1 port map( A1 => n9930, A2 => n18523, Z => n18522);
   U27274 : INV_X2 port map( I => n18542, ZN => n19397);
   U27277 : XOR2_X1 port map( A1 => n5021, A2 => n33569, Z => n18546);
   U27280 : NOR2_X1 port map( A1 => n19203, A2 => n18549, ZN => n26273);
   U27282 : XOR2_X1 port map( A1 => n18554, A2 => n20329, Z => Ciphertext(158))
                           ;
   U27285 : XOR2_X1 port map( A1 => n25317, A2 => n25028, Z => n18557);
   U27287 : XOR2_X1 port map( A1 => Plaintext(75), A2 => Key(75), Z => n19496);
   U27291 : XOR2_X1 port map( A1 => n12690, A2 => n18579, Z => n18578);
   U27295 : XNOR2_X1 port map( A1 => Plaintext(51), A2 => Key(51), ZN => n18585
                           );
   U27304 : XOR2_X1 port map( A1 => n26532, A2 => n19721, Z => n18609);
   U27305 : NOR2_X1 port map( A1 => n38142, A2 => n29284, ZN => n18610);
   U27308 : XOR2_X1 port map( A1 => n23778, A2 => n29920, Z => n18612);
   U27310 : XOR2_X1 port map( A1 => n14386, A2 => n23834, Z => n18620);
   U27313 : XOR2_X1 port map( A1 => n22500, A2 => n18635, Z => n18634);
   U27315 : XOR2_X1 port map( A1 => n25208, A2 => n18643, Z => n18642);
   U27316 : NOR2_X1 port map( A1 => n11411, A2 => n4116, ZN => n18645);
   U27318 : NAND2_X1 port map( A1 => n18659, A2 => n29581, ZN => n18658);
   U27319 : NAND2_X1 port map( A1 => n28843, A2 => n39830, ZN => n18659);
   U27320 : NAND2_X1 port map( A1 => n13508, A2 => n28758, ZN => n19796);
   U27323 : NAND2_X1 port map( A1 => n23006, A2 => n18679, ZN => n23007);
   U27324 : XOR2_X1 port map( A1 => n18692, A2 => n18690, Z => n19954);
   U27325 : XOR2_X1 port map( A1 => n22728, A2 => n18691, Z => n18690);
   U27326 : XOR2_X1 port map( A1 => n20335, A2 => n22580, Z => n18692);
   U27328 : XOR2_X1 port map( A1 => n20976, A2 => n19720, Z => n27161);
   U27330 : XOR2_X1 port map( A1 => Plaintext(62), A2 => Key(62), Z => n18723);
   U27331 : XOR2_X1 port map( A1 => n27556, A2 => n27853, Z => n18709);
   U27332 : INV_X1 port map( I => n26804, ZN => n18719);
   U27333 : INV_X2 port map( I => n18723, ZN => n20266);
   U27334 : NAND2_X2 port map( A1 => n18726, A2 => n18725, ZN => n29574);
   U27336 : XOR2_X1 port map( A1 => n18738, A2 => n18735, Z => n18741);
   U27337 : XOR2_X1 port map( A1 => n18737, A2 => n18736, Z => n18735);
   U27343 : NOR2_X1 port map( A1 => n22797, A2 => n18750, ZN => n20109);
   U27345 : XOR2_X1 port map( A1 => n20698, A2 => n29394, Z => n18764);
   U27347 : XOR2_X1 port map( A1 => Plaintext(48), A2 => Key(48), Z => n18774);
   U27348 : INV_X2 port map( I => n18774, ZN => n21684);
   U27350 : OAI21_X1 port map( A1 => n19434, A2 => n21882, B => n18784, ZN => 
                           n21884);
   U27356 : AND2_X1 port map( A1 => n29672, A2 => n29684, Z => n18793);
   U27358 : XOR2_X1 port map( A1 => n26254, A2 => n18797, Z => n18796);
   U27359 : XOR2_X1 port map( A1 => n26244, A2 => n26349, Z => n18797);
   U27360 : XOR2_X1 port map( A1 => n27802, A2 => n30085, Z => n18800);
   U27361 : NAND3_X1 port map( A1 => n39048, A2 => n31626, A3 => n17791, ZN => 
                           n25705);
   U27362 : NAND2_X1 port map( A1 => n27247, A2 => n7973, ZN => n20455);
   U27363 : XOR2_X1 port map( A1 => n18811, A2 => n14571, Z => n20196);
   U27364 : XOR2_X1 port map( A1 => n7549, A2 => n30063, Z => n18817);
   U27366 : XOR2_X1 port map( A1 => n23829, A2 => n29003, Z => n18828);
   U27367 : MUX2_X1 port map( I0 => n10118, I1 => n30117, S => n30109, Z => 
                           n30118);
   U27369 : XOR2_X1 port map( A1 => n22700, A2 => n18834, Z => n18833);
   U27376 : XOR2_X1 port map( A1 => n18846, A2 => n18847, Z => n28132);
   U27378 : XOR2_X1 port map( A1 => n844, A2 => n1237, Z => n18852);
   U27380 : XOR2_X1 port map( A1 => Plaintext(188), A2 => Key(188), Z => n21722
                           );
   U27388 : XOR2_X1 port map( A1 => n33194, A2 => n29399, Z => n18887);
   U27389 : MUX2_X1 port map( I0 => n23295, I1 => n23294, S => n35001, Z => 
                           n18890);
   U27390 : XOR2_X1 port map( A1 => n39348, A2 => n13639, Z => n28876);
   U27393 : NAND2_X1 port map( A1 => n18897, A2 => n29981, ZN => n29965);
   U27395 : AOI21_X1 port map( A1 => n31512, A2 => n29980, B => n18897, ZN => 
                           n19143);
   U27397 : XOR2_X1 port map( A1 => n17653, A2 => n29808, Z => n18898);
   U27401 : XOR2_X1 port map( A1 => n28982, A2 => n19583, Z => n18905);
   U27402 : XOR2_X1 port map( A1 => n18211, A2 => n19681, Z => n24711);
   U27403 : XOR2_X1 port map( A1 => n18914, A2 => n18911, Z => n23102);
   U27404 : XOR2_X1 port map( A1 => n18913, A2 => n18912, Z => n18911);
   U27405 : XOR2_X1 port map( A1 => n22443, A2 => n22453, Z => n18913);
   U27409 : XOR2_X1 port map( A1 => n23734, A2 => n23733, Z => n18921);
   U27413 : XOR2_X1 port map( A1 => n25009, A2 => n20592, Z => n18930);
   U27414 : XOR2_X1 port map( A1 => n26163, A2 => n29325, Z => n18934);
   U27415 : XOR2_X1 port map( A1 => n23813, A2 => n23915, Z => n18935);
   U27416 : XOR2_X1 port map( A1 => n20753, A2 => n18943, Z => n18942);
   U27420 : NAND2_X1 port map( A1 => n23532, A2 => n6217, ZN => n23222);
   U27424 : INV_X2 port map( I => n18968, ZN => n21928);
   U27427 : XOR2_X1 port map( A1 => n23598, A2 => n18977, Z => n18976);
   U27428 : XOR2_X1 port map( A1 => n37701, A2 => n30203, Z => n18977);
   U27429 : MUX2_X1 port map( I0 => n1299, I1 => n23516, S => n12396, Z => 
                           n23520);
   U27430 : NOR2_X1 port map( A1 => n18985, A2 => n37758, ZN => n18984);
   U27431 : NAND2_X1 port map( A1 => n31663, A2 => n28661, ZN => n18985);
   U27434 : XOR2_X1 port map( A1 => n15930, A2 => n18993, Z => n18992);
   U27436 : INV_X2 port map( I => n19001, ZN => n23149);
   U27437 : INV_X2 port map( I => n19008, ZN => n19599);
   U27438 : XOR2_X1 port map( A1 => n28858, A2 => n28859, Z => n19008);
   U27442 : XOR2_X1 port map( A1 => n21201, A2 => n22579, Z => n19015);
   U27446 : XOR2_X1 port map( A1 => n26370, A2 => n19019, Z => n19018);
   U27449 : XOR2_X1 port map( A1 => n25240, A2 => n29920, Z => n19022);
   U27450 : XOR2_X1 port map( A1 => n334, A2 => n19940, Z => n19025);
   U27452 : XOR2_X1 port map( A1 => n19031, A2 => n30120, Z => Ciphertext(160))
                           ;
   U27453 : NAND2_X1 port map( A1 => n19709, A2 => n18266, ZN => n21392);
   U27454 : NOR2_X1 port map( A1 => n19416, A2 => n18266, ZN => n21541);
   U27455 : NAND2_X1 port map( A1 => n26988, A2 => n19045, ZN => n26991);
   U27457 : XOR2_X1 port map( A1 => n34564, A2 => n19613, Z => n20069);
   U27459 : XOR2_X1 port map( A1 => n518, A2 => n37357, Z => n19155);
   U27464 : XOR2_X1 port map( A1 => n19067, A2 => n28898, Z => n19066);
   U27465 : XOR2_X1 port map( A1 => n29242, A2 => n1719, Z => n19078);
   U27467 : NAND2_X1 port map( A1 => n19084, A2 => n21770, ZN => n21771);
   U27469 : NOR2_X1 port map( A1 => n38142, A2 => n19085, ZN => n29267);
   U27470 : NAND3_X1 port map( A1 => n19091, A2 => n21465, A3 => n34922, ZN => 
                           n20750);
   U27472 : XOR2_X1 port map( A1 => n24061, A2 => n14668, Z => n24063);
   U27473 : XOR2_X1 port map( A1 => n24005, A2 => n14668, Z => n24007);
   U27474 : NAND2_X1 port map( A1 => n19097, A2 => n29929, ZN => n29918);
   U27476 : XOR2_X1 port map( A1 => n26224, A2 => n26207, Z => n19099);
   U27478 : XOR2_X1 port map( A1 => n24068, A2 => n19101, Z => n19100);
   U27479 : XOR2_X1 port map( A1 => n24064, A2 => n19102, Z => n19101);
   U27482 : MUX2_X1 port map( I0 => n24704, I1 => n24705, S => n38674, Z => 
                           n24706);
   U27486 : XOR2_X1 port map( A1 => n29254, A2 => n19721, Z => n19126);
   U27487 : NAND2_X2 port map( A1 => n19129, A2 => n19130, ZN => n29339);
   U27488 : NAND2_X1 port map( A1 => n21285, A2 => n105, ZN => n19312);
   U27490 : XOR2_X1 port map( A1 => n19138, A2 => n1735, Z => Ciphertext(126));
   U27491 : XOR2_X1 port map( A1 => n11974, A2 => n29295, Z => n19145);
   U27495 : XOR2_X1 port map( A1 => n25315, A2 => n19155, Z => n19154);
   U27496 : NOR2_X1 port map( A1 => n19157, A2 => n29410, ZN => n20132);
   U27497 : XOR2_X1 port map( A1 => n29818, A2 => n1737, Z => n19160);
   U27498 : AOI21_X1 port map( A1 => n19164, A2 => n30252, B => n31529, ZN => 
                           n19163);
   U27500 : INV_X2 port map( I => n19170, ZN => n28237);
   U27502 : XOR2_X1 port map( A1 => n19185, A2 => n19182, Z => n27964);
   U27503 : XOR2_X1 port map( A1 => n19184, A2 => n19183, Z => n19182);
   U27504 : XOR2_X1 port map( A1 => n34332, A2 => n27862, Z => n19184);
   U27505 : XOR2_X1 port map( A1 => n27565, A2 => n27500, Z => n19185);
   U27506 : XOR2_X1 port map( A1 => n11923, A2 => n16618, Z => n19186);
   U27507 : XOR2_X1 port map( A1 => n9701, A2 => n25196, Z => n19187);
   U27509 : INV_X2 port map( I => n19955, ZN => n25606);
   U27510 : XOR2_X1 port map( A1 => n22713, A2 => n19201, Z => n19200);
   U27514 : NAND2_X1 port map( A1 => n27272, A2 => n35228, ZN => n19300);
   U27515 : XOR2_X1 port map( A1 => n27532, A2 => n35229, Z => n19213);
   U27518 : NOR2_X1 port map( A1 => n12672, A2 => n25048, ZN => n25049);
   U27519 : XOR2_X1 port map( A1 => n19824, A2 => n4348, Z => n19220);
   U27521 : NAND2_X1 port map( A1 => n20276, A2 => n33786, ZN => n23414);
   U27522 : NAND2_X2 port map( A1 => n20059, A2 => n20062, ZN => n26594);
   U27529 : NOR2_X1 port map( A1 => n27279, A2 => n21144, ZN => n19456);
   U27530 : NOR2_X1 port map( A1 => n33538, A2 => n23516, ZN => n19249);
   U27531 : XOR2_X1 port map( A1 => n22693, A2 => n21994, Z => n22004);
   U27532 : XOR2_X1 port map( A1 => n38641, A2 => n38993, Z => n24858);
   U27533 : XOR2_X1 port map( A1 => n25097, A2 => n25096, Z => n25099);
   U27534 : INV_X1 port map( I => n34914, ZN => n29583);
   U27535 : INV_X2 port map( I => n19266, ZN => n20053);
   U27538 : XOR2_X1 port map( A1 => n28542, A2 => n19277, Z => n28883);
   U27539 : XOR2_X1 port map( A1 => n28540, A2 => n28541, Z => n19277);
   U27541 : XOR2_X1 port map( A1 => n29140, A2 => n29119, Z => n20447);
   U27542 : NOR2_X1 port map( A1 => n13410, A2 => n25611, ZN => n25412);
   U27544 : NOR2_X1 port map( A1 => n26564, A2 => n26905, ZN => n19285);
   U27547 : XOR2_X1 port map( A1 => n22624, A2 => n22773, Z => n22514);
   U27548 : NAND2_X1 port map( A1 => n37230, A2 => n24241, ZN => n24242);
   U27551 : NAND2_X1 port map( A1 => n15509, A2 => n920, ZN => n19303);
   U27552 : NOR2_X2 port map( A1 => n19305, A2 => n19304, ZN => n19741);
   U27555 : OR2_X1 port map( A1 => n29764, A2 => n19568, Z => n28862);
   U27556 : XOR2_X1 port map( A1 => n28983, A2 => n1375, Z => n19309);
   U27557 : XOR2_X1 port map( A1 => Key(149), A2 => Plaintext(149), Z => n19313
                           );
   U27559 : XOR2_X1 port map( A1 => n19316, A2 => n1697, Z => Ciphertext(140));
   U27560 : NOR2_X1 port map( A1 => n30013, A2 => n30012, ZN => n19316);
   U27563 : BUF_X2 port map( I => n21735, Z => n19323);
   U27565 : XOR2_X1 port map( A1 => n22676, A2 => n30126, Z => n20980);
   U27568 : NOR2_X1 port map( A1 => n21734, A2 => n21919, ZN => n19335);
   U27569 : BUF_X2 port map( I => n21875, Z => n19337);
   U27572 : OR2_X1 port map( A1 => n22135, A2 => n11044, Z => n22018);
   U27573 : NOR2_X1 port map( A1 => n29708, A2 => n29721, ZN => n19347);
   U27579 : XOR2_X1 port map( A1 => n22569, A2 => n22449, Z => n22413);
   U27582 : NAND2_X2 port map( A1 => n25344, A2 => n25343, ZN => n25941);
   U27586 : XOR2_X1 port map( A1 => n23693, A2 => n23692, Z => n24095);
   U27589 : BUF_X2 port map( I => n26921, Z => n19371);
   U27592 : OAI21_X1 port map( A1 => n11171, A2 => n1672, B => n19385, ZN => 
                           n22010);
   U27597 : INV_X1 port map( I => n29419, ZN => n19404);
   U27598 : NOR2_X1 port map( A1 => n29652, A2 => n17382, ZN => n19411);
   U27601 : OAI21_X2 port map( A1 => n25439, A2 => n19400, B => n25438, ZN => 
                           n26041);
   U27604 : XOR2_X1 port map( A1 => n20747, A2 => n27573, Z => n19421);
   U27607 : NAND2_X1 port map( A1 => n24842, A2 => n24733, ZN => n19595);
   U27609 : INV_X1 port map( I => n27197, ZN => n27279);
   U27611 : OAI21_X1 port map( A1 => n1240, A2 => n33237, B => n19439, ZN => 
                           n26095);
   U27613 : XOR2_X1 port map( A1 => n21186, A2 => n19445, Z => n19444);
   U27614 : XOR2_X1 port map( A1 => n19446, A2 => n20822, Z => n20821);
   U27620 : INV_X2 port map( I => n19459, ZN => n26695);
   U27625 : XOR2_X1 port map( A1 => n21381, A2 => Key(140), Z => n21608);
   U27630 : BUF_X2 port map( I => n21777, Z => n19479);
   U27631 : XOR2_X1 port map( A1 => n19744, A2 => n19493, Z => n19492);
   U27633 : XOR2_X1 port map( A1 => n18273, A2 => n29808, Z => n26285);
   U27641 : AOI22_X2 port map( A1 => n21543, A2 => n21542, B1 => n21541, B2 => 
                           n21540, ZN => n21973);
   U27643 : INV_X2 port map( I => n29721, ZN => n29712);
   U27645 : OAI21_X1 port map( A1 => n25647, A2 => n25429, B => n19532, ZN => 
                           n25430);
   U27646 : XOR2_X1 port map( A1 => n19533, A2 => n26230, Z => n19867);
   U27647 : NOR2_X1 port map( A1 => n7725, A2 => n9188, ZN => n21256);
   U27648 : OAI21_X1 port map( A1 => n17568, A2 => n36839, B => n14561, ZN => 
                           n22684);
   U27649 : OR2_X1 port map( A1 => n30212, A2 => n39083, Z => n30205);
   U27650 : NAND2_X1 port map( A1 => n21812, A2 => n21683, ZN => n19552);
   U27655 : AOI21_X1 port map( A1 => n20725, A2 => n27201, B => n35895, ZN => 
                           n27076);
   U27656 : XOR2_X1 port map( A1 => n16897, A2 => n25086, Z => n25088);
   U27657 : INV_X1 port map( I => n28546, ZN => n28322);
   U27658 : INV_X2 port map( I => n19576, ZN => n24433);
   U27664 : XOR2_X1 port map( A1 => n26518, A2 => n26402, Z => n20260);
   U27668 : OR2_X1 port map( A1 => n37183, A2 => n18545, Z => n20644);
   U27674 : XOR2_X1 port map( A1 => n19617, A2 => n15181, Z => Ciphertext(42));
   U27676 : XOR2_X1 port map( A1 => n26561, A2 => n26562, Z => n19632);
   U27677 : XOR2_X1 port map( A1 => n11721, A2 => n28815, Z => n19640);
   U27683 : XOR2_X1 port map( A1 => n19652, A2 => n20096, Z => n20095);
   U27684 : INV_X1 port map( I => n12410, ZN => n20570);
   U27688 : INV_X1 port map( I => n25555, ZN => n20237);
   U27689 : NOR2_X1 port map( A1 => n14453, A2 => n26614, ZN => n26851);
   U27695 : XOR2_X1 port map( A1 => Plaintext(118), A2 => Key(118), Z => n19822
                           );
   U27697 : AND2_X1 port map( A1 => n33073, A2 => n35116, Z => n21661);
   U27698 : INV_X1 port map( I => n24420, ZN => n24442);
   U27699 : INV_X2 port map( I => n21752, ZN => n19709);
   U27701 : OAI21_X1 port map( A1 => n452, A2 => n10120, B => n7278, ZN => 
                           n21626);
   U27702 : XOR2_X1 port map( A1 => Key(135), A2 => Plaintext(135), Z => n21790
                           );
   U27704 : NAND2_X1 port map( A1 => n28381, A2 => n28382, ZN => n28385);
   U27705 : XOR2_X1 port map( A1 => n27687, A2 => n19775, Z => n20096);
   U27709 : XOR2_X1 port map( A1 => n26481, A2 => n26438, Z => n19744);
   U27710 : NOR2_X2 port map( A1 => n19747, A2 => n20473, ZN => n29684);
   U27712 : INV_X2 port map( I => n19764, ZN => n27969);
   U27716 : XOR2_X1 port map( A1 => n19784, A2 => n29476, Z => Ciphertext(52));
   U27717 : NAND2_X1 port map( A1 => n20809, A2 => n20808, ZN => n23289);
   U27718 : XOR2_X1 port map( A1 => n23691, A2 => n19792, Z => n23693);
   U27719 : XOR2_X1 port map( A1 => n23690, A2 => n39073, Z => n19792);
   U27720 : XOR2_X1 port map( A1 => n26223, A2 => n19799, Z => n19798);
   U27722 : XOR2_X1 port map( A1 => n27829, A2 => n29808, Z => n20796);
   U27724 : XOR2_X1 port map( A1 => n25188, A2 => n25190, Z => n19809);
   U27727 : OAI21_X1 port map( A1 => n22110, A2 => n22111, B => n133, ZN => 
                           n19812);
   U27728 : XOR2_X1 port map( A1 => n27564, A2 => n27799, Z => n27769);
   U27729 : INV_X1 port map( I => n21875, ZN => n21696);
   U27733 : INV_X2 port map( I => n19838, ZN => n20830);
   U27736 : INV_X1 port map( I => n29837, ZN => n28819);
   U27737 : NOR2_X1 port map( A1 => n22184, A2 => n1048, ZN => n22186);
   U27740 : INV_X1 port map( I => n24683, ZN => n24774);
   U27743 : INV_X2 port map( I => n21630, ZN => n21775);
   U27746 : OAI21_X2 port map( A1 => n27742, A2 => n27743, B => n27741, ZN => 
                           n28753);
   U27747 : INV_X2 port map( I => n19867, ZN => n26974);
   U27749 : XOR2_X1 port map( A1 => n9246, A2 => n29680, Z => n19983);
   U27751 : XOR2_X1 port map( A1 => n21142, A2 => n19882, Z => n19881);
   U27755 : XOR2_X1 port map( A1 => n26210, A2 => n26209, Z => n19900);
   U27756 : NAND2_X1 port map( A1 => n20833, A2 => n25945, ZN => n25946);
   U27757 : XOR2_X1 port map( A1 => n18273, A2 => n30150, Z => n25947);
   U27762 : INV_X2 port map( I => n19920, ZN => n29642);
   U27765 : OAI21_X1 port map( A1 => n13767, A2 => n19924, B => n1308, ZN => 
                           n19923);
   U27766 : BUF_X2 port map( I => Key(54), Z => n19933);
   U27770 : OR2_X1 port map( A1 => n21933, A2 => n20476, Z => n19985);
   U27772 : XOR2_X1 port map( A1 => n22433, A2 => n19954, Z => n22973);
   U27777 : INV_X2 port map( I => n18576, ZN => n21820);
   U27778 : INV_X1 port map( I => n29624, ZN => n29608);
   U27779 : XOR2_X1 port map( A1 => n27806, A2 => n19988, Z => n19987);
   U27780 : XOR2_X1 port map( A1 => n27749, A2 => n29320, Z => n19988);
   U27784 : NAND2_X2 port map( A1 => n20008, A2 => n20007, ZN => n25814);
   U27785 : NOR3_X1 port map( A1 => n15350, A2 => n22341, A3 => n22342, ZN => 
                           n22343);
   U27786 : XOR2_X1 port map( A1 => n29167, A2 => n28868, Z => n20033);
   U27789 : XOR2_X1 port map( A1 => n23876, A2 => n20045, Z => n20044);
   U27792 : INV_X1 port map( I => n19676, ZN => n20489);
   U27793 : XOR2_X1 port map( A1 => n24047, A2 => n19676, Z => n23690);
   U27795 : INV_X2 port map( I => n20063, ZN => n26852);
   U27796 : XOR2_X1 port map( A1 => n26254, A2 => n14670, Z => n20065);
   U27799 : INV_X2 port map( I => n24224, ZN => n24432);
   U27800 : NAND2_X2 port map( A1 => n20090, A2 => n20089, ZN => n22503);
   U27801 : XOR2_X1 port map( A1 => n27800, A2 => n27797, Z => n20093);
   U27802 : XOR2_X1 port map( A1 => n20098, A2 => n20097, Z => n20858);
   U27803 : XOR2_X1 port map( A1 => n26401, A2 => n749, Z => n20097);
   U27804 : XOR2_X1 port map( A1 => n26593, A2 => n26261, Z => n20101);
   U27807 : XOR2_X1 port map( A1 => n26347, A2 => n14568, Z => n20107);
   U27809 : OAI21_X1 port map( A1 => n29491, A2 => n29418, B => n20113, ZN => 
                           n29419);
   U27810 : XOR2_X1 port map( A1 => n26073, A2 => n26059, Z => n20117);
   U27811 : INV_X1 port map( I => n35273, ZN => n29604);
   U27812 : XOR2_X1 port map( A1 => n20129, A2 => n17275, Z => Ciphertext(39));
   U27816 : XOR2_X1 port map( A1 => n27607, A2 => n35270, Z => n20167);
   U27817 : INV_X1 port map( I => n24728, ZN => n24727);
   U27819 : INV_X2 port map( I => n20194, ZN => n25695);
   U27820 : INV_X2 port map( I => n20196, ZN => n24381);
   U27821 : XOR2_X1 port map( A1 => Plaintext(110), A2 => Key(110), Z => n21330
                           );
   U27822 : XOR2_X1 port map( A1 => n24047, A2 => n20205, Z => n23871);
   U27823 : XOR2_X1 port map( A1 => n23968, A2 => n20205, Z => n23720);
   U27824 : INV_X1 port map( I => n26207, ZN => n26472);
   U27828 : MUX2_X1 port map( I0 => n22098, I1 => n22099, S => n32609, Z => 
                           n22105);
   U27834 : XOR2_X1 port map( A1 => n20261, A2 => n20262, Z => n20257);
   U27836 : XOR2_X1 port map( A1 => n26487, A2 => n26520, Z => n20262);
   U27840 : XOR2_X1 port map( A1 => n26263, A2 => n25511, Z => n20268);
   U27843 : INV_X2 port map( I => n33999, ZN => n21712);
   U27846 : XOR2_X1 port map( A1 => n26461, A2 => n26464, Z => n20279);
   U27847 : XOR2_X1 port map( A1 => n18133, A2 => n28776, Z => n28777);
   U27852 : INV_X2 port map( I => n20300, ZN => n21506);
   U27855 : NOR2_X1 port map( A1 => n30145, A2 => n18588, ZN => n30147);
   U27856 : AOI21_X1 port map( A1 => n30145, A2 => n18588, B => n34177, ZN => 
                           n30138);
   U27857 : NOR2_X2 port map( A1 => n26733, A2 => n26732, ZN => n27267);
   U27860 : XOR2_X1 port map( A1 => n20325, A2 => n20323, Z => n29941);
   U27861 : XOR2_X1 port map( A1 => n29072, A2 => n29003, Z => n20324);
   U27863 : NOR2_X1 port map( A1 => n11851, A2 => n21762, ZN => n20332);
   U27864 : XOR2_X1 port map( A1 => n20333, A2 => n25278, Z => n25120);
   U27865 : INV_X2 port map( I => n26931, ZN => n26564);
   U27869 : INV_X1 port map( I => n23861, ZN => n24020);
   U27870 : NAND2_X1 port map( A1 => n20544, A2 => n21779, ZN => n20348);
   U27871 : XOR2_X1 port map( A1 => n16639, A2 => n30065, Z => n28318);
   U27872 : XOR2_X1 port map( A1 => n18180, A2 => n29522, Z => n26241);
   U27873 : INV_X2 port map( I => n20361, ZN => n21808);
   U27876 : XOR2_X1 port map( A1 => n20365, A2 => n24973, Z => n25418);
   U27881 : XOR2_X1 port map( A1 => n20392, A2 => n30090, Z => n22501);
   U27883 : XOR2_X1 port map( A1 => n27490, A2 => n27819, Z => n20400);
   U27884 : XOR2_X1 port map( A1 => n39295, A2 => n19936, Z => n20409);
   U27892 : XOR2_X1 port map( A1 => n28895, A2 => n28894, Z => n29344);
   U27894 : XOR2_X1 port map( A1 => n38150, A2 => n31548, Z => n20446);
   U27895 : XOR2_X1 port map( A1 => n21284, A2 => n27550, Z => n20448);
   U27897 : XOR2_X1 port map( A1 => n20452, A2 => n18432, Z => n29132);
   U27898 : XOR2_X1 port map( A1 => n20452, A2 => n30170, Z => n28853);
   U27900 : XOR2_X1 port map( A1 => n20452, A2 => n19815, Z => n28973);
   U27902 : NAND2_X1 port map( A1 => n25336, A2 => n25337, ZN => n20463);
   U27906 : XOR2_X1 port map( A1 => Plaintext(24), A2 => Key(24), Z => n21849);
   U27909 : XOR2_X1 port map( A1 => n26349, A2 => n20489, Z => n26526);
   U27910 : NAND2_X1 port map( A1 => n37776, A2 => n28380, ZN => n20497);
   U27911 : XOR2_X1 port map( A1 => n21225, A2 => n22673, Z => n20502);
   U27916 : XOR2_X1 port map( A1 => Plaintext(121), A2 => Key(121), Z => n21740
                           );
   U27918 : OAI21_X1 port map( A1 => n28028, A2 => n33331, B => n33307, ZN => 
                           n28029);
   U27919 : INV_X2 port map( I => n20526, ZN => n24408);
   U27926 : XOR2_X1 port map( A1 => n22420, A2 => n22421, Z => n20555);
   U27927 : INV_X2 port map( I => n20555, ZN => n23089);
   U27929 : XOR2_X1 port map( A1 => Plaintext(136), A2 => Key(136), Z => n21791
                           );
   U27931 : XOR2_X1 port map( A1 => n20559, A2 => n19925, Z => Ciphertext(13));
   U27933 : XOR2_X1 port map( A1 => n25191, A2 => n662, Z => n20571);
   U27935 : NAND2_X1 port map( A1 => n547, A2 => n21571, ZN => n20593);
   U27936 : XOR2_X1 port map( A1 => Plaintext(70), A2 => Key(70), Z => n20694);
   U27938 : XNOR2_X1 port map( A1 => n21426, A2 => Key(1), ZN => n20596);
   U27939 : INV_X2 port map( I => n20601, ZN => n24241);
   U27947 : NAND2_X1 port map( A1 => n23075, A2 => n23076, ZN => n20625);
   U27949 : NAND2_X1 port map( A1 => n23210, A2 => n20408, ZN => n20741);
   U27950 : XOR2_X1 port map( A1 => n33470, A2 => n27829, Z => n20641);
   U27953 : XOR2_X1 port map( A1 => n20656, A2 => n26377, Z => n21277);
   U27955 : NAND2_X1 port map( A1 => n26607, A2 => n20666, ZN => n26608);
   U27956 : XOR2_X1 port map( A1 => n20675, A2 => n28579, Z => n20674);
   U27957 : INV_X2 port map( I => n20677, ZN => n29598);
   U27958 : XOR2_X1 port map( A1 => n28829, A2 => n28828, Z => n20684);
   U27959 : INV_X2 port map( I => n20685, ZN => n21924);
   U27961 : INV_X2 port map( I => n20694, ZN => n21810);
   U27963 : INV_X2 port map( I => n20702, ZN => n21023);
   U27964 : XOR2_X1 port map( A1 => n20707, A2 => n29671, Z => n25143);
   U27965 : XOR2_X1 port map( A1 => n17758, A2 => n18700, Z => n20713);
   U27966 : XOR2_X1 port map( A1 => n24063, A2 => n20717, Z => n20716);
   U27967 : XOR2_X1 port map( A1 => n24059, A2 => n19751, Z => n20717);
   U27969 : XOR2_X1 port map( A1 => n27724, A2 => n27766, Z => n20723);
   U27970 : INV_X2 port map( I => n20726, ZN => n29455);
   U27973 : BUF_X2 port map( I => n25351, Z => n25616);
   U27978 : OAI21_X2 port map( A1 => n5059, A2 => n27405, B => n27083, ZN => 
                           n27799);
   U27979 : XOR2_X1 port map( A1 => n19770, A2 => n27754, Z => n20747);
   U27983 : OR2_X1 port map( A1 => n26355, A2 => n26354, Z => n20764);
   U27984 : XOR2_X1 port map( A1 => n37044, A2 => n23950, Z => n20767);
   U27985 : MUX2_X1 port map( I0 => n26023, I1 => n20771, S => n1105, Z => 
                           n20770);
   U27986 : XOR2_X1 port map( A1 => Plaintext(81), A2 => Key(81), Z => n21488);
   U27988 : XOR2_X1 port map( A1 => n25178, A2 => n20780, Z => n20779);
   U27989 : XOR2_X1 port map( A1 => n25301, A2 => n20781, Z => n20780);
   U27990 : XOR2_X1 port map( A1 => n22490, A2 => n22633, Z => n20794);
   U27992 : XOR2_X1 port map( A1 => n38201, A2 => n20804, Z => n20803);
   U27993 : XNOR2_X1 port map( A1 => Plaintext(58), A2 => Key(58), ZN => n20810
                           );
   U27995 : INV_X2 port map( I => n20821, ZN => n30049);
   U27996 : XOR2_X1 port map( A1 => n29830, A2 => n29834, Z => n20822);
   U27997 : XOR2_X1 port map( A1 => n30733, A2 => n20483, Z => n20824);
   U27998 : NAND3_X1 port map( A1 => n21422, A2 => n275, A3 => n21843, ZN => 
                           n20825);
   U27999 : XOR2_X1 port map( A1 => n6727, A2 => n18981, Z => n20828);
   U28000 : XOR2_X1 port map( A1 => n20836, A2 => n22753, Z => n23129);
   U28001 : OAI21_X1 port map( A1 => n21635, A2 => n21942, B => n19546, ZN => 
                           n21638);
   U28005 : INV_X2 port map( I => n20866, ZN => n29777);
   U28006 : INV_X1 port map( I => n27389, ZN => n27291);
   U28008 : XOR2_X1 port map( A1 => Plaintext(84), A2 => Key(84), Z => n21880);
   U28009 : XOR2_X1 port map( A1 => n26436, A2 => n26435, Z => n20886);
   U28010 : XNOR2_X1 port map( A1 => Plaintext(156), A2 => Key(156), ZN => 
                           n20887);
   U28014 : XOR2_X1 port map( A1 => Plaintext(158), A2 => Key(158), Z => n21496
                           );
   U28015 : XOR2_X1 port map( A1 => n24561, A2 => n20893, Z => n20892);
   U28016 : XOR2_X1 port map( A1 => n7247, A2 => n25274, Z => n20893);
   U28017 : NAND2_X1 port map( A1 => n1404, A2 => n14417, ZN => n20901);
   U28018 : NOR2_X1 port map( A1 => n24419, A2 => n1596, ZN => n20903);
   U28026 : XOR2_X1 port map( A1 => n20939, A2 => n1719, Z => Ciphertext(105));
   U28027 : INV_X2 port map( I => n29797, ZN => n29788);
   U28032 : NAND2_X1 port map( A1 => n29797, A2 => n20963, ZN => n20962);
   U28034 : NOR2_X1 port map( A1 => n26800, A2 => n20120, ZN => n26801);
   U28037 : XOR2_X1 port map( A1 => n21009, A2 => n1723, Z => Ciphertext(102));
   U28038 : INV_X2 port map( I => n28132, ZN => n28229);
   U28039 : XOR2_X1 port map( A1 => Plaintext(45), A2 => Key(45), Z => n21674);
   U28042 : XOR2_X1 port map( A1 => n10560, A2 => n23838, Z => n23839);
   U28043 : XOR2_X1 port map( A1 => n27863, A2 => n29974, Z => n21044);
   U28045 : XOR2_X1 port map( A1 => n25133, A2 => n33208, Z => n25134);
   U28046 : OR2_X1 port map( A1 => n272, A2 => n22875, Z => n21063);
   U28047 : MUX2_X1 port map( I0 => n21065, I1 => n22769, S => n32228, Z => 
                           n21064);
   U28050 : XOR2_X1 port map( A1 => n29125, A2 => n17039, Z => n21076);
   U28052 : XOR2_X1 port map( A1 => n39032, A2 => n37882, Z => n21086);
   U28053 : XOR2_X1 port map( A1 => n36905, A2 => n19903, Z => n21095);
   U28054 : XOR2_X1 port map( A1 => n29145, A2 => n29146, Z => n21097);
   U28055 : INV_X1 port map( I => n9151, ZN => n21100);
   U28059 : XOR2_X1 port map( A1 => n21134, A2 => n22414, Z => n21133);
   U28060 : NOR2_X1 port map( A1 => n2799, A2 => n954, ZN => n21135);
   U28061 : NOR2_X1 port map( A1 => n29732, A2 => n29754, ZN => n21146);
   U28062 : NAND2_X1 port map( A1 => n29741, A2 => n29754, ZN => n21147);
   U28065 : XOR2_X1 port map( A1 => n21158, A2 => n32218, Z => Ciphertext(65));
   U28067 : XOR2_X1 port map( A1 => n21162, A2 => n21161, Z => n29586);
   U28068 : XOR2_X1 port map( A1 => n28767, A2 => n28762, Z => n21161);
   U28074 : XOR2_X1 port map( A1 => n29833, A2 => n19758, Z => n21172);
   U28076 : XOR2_X1 port map( A1 => n24417, A2 => n24932, Z => n21174);
   U28077 : XOR2_X1 port map( A1 => n27000, A2 => n27650, Z => n21176);
   U28080 : NAND3_X1 port map( A1 => n37102, A2 => n26695, A3 => n946, ZN => 
                           n21191);
   U28082 : XOR2_X1 port map( A1 => n359, A2 => n19649, Z => n21197);
   U28084 : XOR2_X1 port map( A1 => n9074, A2 => n22445, Z => n21206);
   U28086 : NOR2_X1 port map( A1 => n28569, A2 => n3900, ZN => n28665);
   U28087 : XOR2_X1 port map( A1 => n21215, A2 => n22025, Z => n21217);
   U28088 : XOR2_X1 port map( A1 => n21217, A2 => n14673, Z => n21216);
   U28089 : XOR2_X1 port map( A1 => n22462, A2 => n21219, Z => n21218);
   U28090 : XOR2_X1 port map( A1 => n22566, A2 => n22670, Z => n21219);
   U28091 : XOR2_X1 port map( A1 => Plaintext(56), A2 => Key(56), Z => n21805);
   U28093 : NAND2_X1 port map( A1 => n7693, A2 => n21231, ZN => n24621);
   U28094 : NAND2_X1 port map( A1 => n24852, A2 => n21231, ZN => n24854);
   U28096 : INV_X2 port map( I => n21234, ZN => n30000);
   U28098 : XOR2_X1 port map( A1 => n29282, A2 => n25303, Z => n21252);
   U28099 : INV_X1 port map( I => n22783, ZN => n22818);
   U28102 : XOR2_X1 port map( A1 => n25113, A2 => n21280, Z => n21279);
   U28103 : NAND2_X1 port map( A1 => n21698, A2 => n1353, ZN => n21701);
   U28105 : AOI21_X1 port map( A1 => n21393, A2 => n1353, B => n19709, ZN => 
                           n21394);
   U28114 : NOR2_X1 port map( A1 => n30134, A2 => n37117, ZN => n30146);
   U28115 : OR2_X1 port map( A1 => n29202, A2 => n6938, Z => n28789);
   U28120 : NAND3_X1 port map( A1 => n28191, A2 => n28189, A3 => n16325, ZN => 
                           n27874);
   U28128 : NAND2_X1 port map( A1 => n23344, A2 => n23430, ZN => n23345);
   U28129 : INV_X1 port map( I => n24104, ZN => n24174);
   U28130 : NAND2_X1 port map( A1 => n25726, A2 => n16168, ZN => n25732);
   U28131 : INV_X1 port map( I => n26172, ZN => n26173);
   U28132 : NOR2_X1 port map( A1 => n21272, A2 => n27165, ZN => n27166);
   U28133 : INV_X1 port map( I => n8875, ZN => n27493);
   U28137 : XOR2_X1 port map( A1 => Key(119), A2 => Plaintext(119), Z => n21754
                           );
   U28138 : XOR2_X1 port map( A1 => Key(115), A2 => Plaintext(115), Z => n21753
                           );
   U28139 : XOR2_X1 port map( A1 => Key(117), A2 => Plaintext(117), Z => n21752
                           );
   U28140 : XOR2_X1 port map( A1 => Key(87), A2 => Plaintext(87), Z => n21577);
   U28141 : INV_X1 port map( I => Plaintext(85), ZN => n21326);
   U28142 : XOR2_X1 port map( A1 => n21326, A2 => Key(85), Z => n21575);
   U28143 : NAND3_X1 port map( A1 => n21593, A2 => n21507, A3 => n21594, ZN => 
                           n21327);
   U28147 : XOR2_X1 port map( A1 => Key(111), A2 => Plaintext(111), Z => n21875
                           );
   U28148 : XOR2_X1 port map( A1 => Key(113), A2 => Plaintext(113), Z => n21871
                           );
   U28150 : INV_X1 port map( I => n21330, ZN => n21876);
   U28151 : INV_X1 port map( I => Plaintext(112), ZN => n21329);
   U28152 : XOR2_X1 port map( A1 => n21329, A2 => Key(112), Z => n21872);
   U28153 : OAI21_X1 port map( A1 => n21546, A2 => n19395, B => n21697, ZN => 
                           n21331);
   U28154 : XOR2_X1 port map( A1 => Key(107), A2 => Plaintext(107), Z => n21750
                           );
   U28155 : INV_X1 port map( I => Plaintext(102), ZN => n21332);
   U28158 : INV_X1 port map( I => Plaintext(40), ZN => n21340);
   U28159 : XOR2_X1 port map( A1 => n21340, A2 => Key(40), Z => n21688);
   U28160 : XOR2_X1 port map( A1 => Plaintext(47), A2 => Key(47), Z => n21432);
   U28161 : INV_X1 port map( I => Plaintext(42), ZN => n21341);
   U28162 : XOR2_X1 port map( A1 => n21341, A2 => Key(42), Z => n21857);
   U28163 : OAI21_X1 port map( A1 => n33053, A2 => n18174, B => n21860, ZN => 
                           n21345);
   U28164 : XOR2_X1 port map( A1 => Key(43), A2 => Plaintext(43), Z => n21823);
   U28167 : INV_X1 port map( I => Plaintext(25), ZN => n21346);
   U28169 : INV_X1 port map( I => Plaintext(27), ZN => n21347);
   U28170 : XOR2_X1 port map( A1 => n21347, A2 => Key(27), Z => n21848);
   U28174 : INV_X1 port map( I => Plaintext(26), ZN => n21350);
   U28175 : XOR2_X1 port map( A1 => n21350, A2 => Key(26), Z => n21846);
   U28176 : XOR2_X1 port map( A1 => Key(19), A2 => Plaintext(19), Z => n21841);
   U28177 : INV_X1 port map( I => Plaintext(50), ZN => n21351);
   U28178 : XOR2_X1 port map( A1 => n21351, A2 => Key(50), Z => n21352);
   U28179 : XOR2_X1 port map( A1 => Key(53), A2 => Plaintext(53), Z => n21814);
   U28180 : XOR2_X1 port map( A1 => Key(52), A2 => Plaintext(52), Z => n21428);
   U28183 : INV_X1 port map( I => Plaintext(35), ZN => n21357);
   U28184 : XOR2_X1 port map( A1 => n21357, A2 => Key(35), Z => n21358);
   U28185 : XOR2_X1 port map( A1 => Key(32), A2 => Plaintext(32), Z => n21835);
   U28186 : XOR2_X1 port map( A1 => Key(34), A2 => Plaintext(34), Z => n21628);
   U28188 : NOR2_X1 port map( A1 => n21665, A2 => n21837, ZN => n21360);
   U28189 : INV_X1 port map( I => Plaintext(60), ZN => n21366);
   U28190 : XOR2_X1 port map( A1 => n21366, A2 => Key(60), Z => n21818);
   U28191 : XOR2_X1 port map( A1 => Key(78), A2 => Plaintext(78), Z => n21368);
   U28192 : INV_X1 port map( I => n21368, ZN => n21568);
   U28193 : INV_X1 port map( I => Plaintext(83), ZN => n21367);
   U28194 : XOR2_X1 port map( A1 => n21367, A2 => Key(83), Z => n21567);
   U28197 : NAND2_X1 port map( A1 => n1350, A2 => n14373, ZN => n21373);
   U28198 : INV_X1 port map( I => Plaintext(68), ZN => n21376);
   U28200 : INV_X1 port map( I => Plaintext(67), ZN => n21378);
   U28201 : INV_X1 port map( I => Plaintext(130), ZN => n21380);
   U28202 : XOR2_X1 port map( A1 => Key(141), A2 => Plaintext(141), Z => n21655
                           );
   U28203 : INV_X1 port map( I => Plaintext(140), ZN => n21381);
   U28204 : INV_X1 port map( I => Plaintext(137), ZN => n21382);
   U28205 : XOR2_X1 port map( A1 => n21382, A2 => Key(137), Z => n21792);
   U28207 : OAI21_X1 port map( A1 => n7062, A2 => n21787, B => n18205, ZN => 
                           n21383);
   U28209 : INV_X1 port map( I => Plaintext(125), ZN => n21386);
   U28211 : XOR2_X1 port map( A1 => Key(122), A2 => Plaintext(122), Z => n21743
                           );
   U28212 : INV_X1 port map( I => Plaintext(124), ZN => n21389);
   U28213 : XOR2_X1 port map( A1 => n21389, A2 => Key(124), Z => n21742);
   U28214 : INV_X1 port map( I => Plaintext(123), ZN => n21390);
   U28215 : XOR2_X1 port map( A1 => n21390, A2 => Key(123), Z => n21741);
   U28216 : AOI21_X1 port map( A1 => n21542, A2 => n21392, B => n19822, ZN => 
                           n21395);
   U28218 : XOR2_X1 port map( A1 => Key(170), A2 => Plaintext(170), Z => n21927
                           );
   U28220 : INV_X1 port map( I => Plaintext(181), ZN => n21398);
   U28221 : XOR2_X1 port map( A1 => n21398, A2 => Key(181), Z => n21905);
   U28222 : INV_X1 port map( I => Plaintext(183), ZN => n21399);
   U28225 : XOR2_X1 port map( A1 => Key(182), A2 => Plaintext(182), Z => n21721
                           );
   U28228 : XOR2_X1 port map( A1 => Key(184), A2 => Plaintext(184), Z => n21641
                           );
   U28229 : NAND2_X1 port map( A1 => n21782, A2 => n35116, ZN => n21402);
   U28230 : INV_X1 port map( I => Plaintext(152), ZN => n21403);
   U28231 : XOR2_X1 port map( A1 => n21403, A2 => Key(152), Z => n21602);
   U28232 : XOR2_X1 port map( A1 => Key(154), A2 => Plaintext(154), Z => n21951
                           );
   U28233 : INV_X1 port map( I => n32664, ZN => n21405);
   U28236 : NAND2_X1 port map( A1 => n21782, A2 => n32664, ZN => n21406);
   U28237 : INV_X1 port map( I => Plaintext(162), ZN => n21407);
   U28238 : XOR2_X1 port map( A1 => n21407, A2 => Key(162), Z => n21630);
   U28239 : XOR2_X1 port map( A1 => Key(165), A2 => Plaintext(165), Z => n21777
                           );
   U28240 : INV_X1 port map( I => Plaintext(163), ZN => n21408);
   U28241 : INV_X1 port map( I => Plaintext(167), ZN => n21409);
   U28242 : XOR2_X1 port map( A1 => n21409, A2 => Key(167), Z => n21937);
   U28243 : XOR2_X1 port map( A1 => Key(166), A2 => Plaintext(166), Z => n21776
                           );
   U28246 : NAND2_X1 port map( A1 => n21862, A2 => n18143, ZN => n21417);
   U28250 : INV_X1 port map( I => Plaintext(1), ZN => n21426);
   U28251 : XOR2_X1 port map( A1 => Key(0), A2 => Plaintext(0), Z => n21735);
   U28254 : AOI21_X1 port map( A1 => n21808, A2 => n21692, B => n38241, ZN => 
                           n21438);
   U28257 : INV_X1 port map( I => n21460, ZN => n22118);
   U28258 : INV_X1 port map( I => n21459, ZN => n22117);
   U28259 : NOR2_X1 port map( A1 => n21756, A2 => n19337, ZN => n21454);
   U28260 : NOR2_X1 port map( A1 => n21546, A2 => n21756, ZN => n21457);
   U28261 : NOR2_X1 port map( A1 => n21697, A2 => n19650, ZN => n21456);
   U28262 : NOR2_X1 port map( A1 => n19647, A2 => n21401, ZN => n21464);
   U28263 : NOR2_X1 port map( A1 => n21644, A2 => n21462, ZN => n21463);
   U28264 : NOR2_X1 port map( A1 => n14837, A2 => n21923, ZN => n21468);
   U28265 : NOR2_X1 port map( A1 => n37612, A2 => n21724, ZN => n21467);
   U28269 : NAND2_X1 port map( A1 => n21485, A2 => n32544, ZN => n21486);
   U28270 : MUX2_X1 port map( I0 => n17209, I1 => n21893, S => n21892, Z => 
                           n21491);
   U28272 : NAND2_X1 port map( A1 => n21806, A2 => n21492, ZN => n21493);
   U28273 : INV_X2 port map( I => n21496, ZN => n21944);
   U28274 : INV_X1 port map( I => n21770, ZN => n21635);
   U28276 : NOR2_X1 port map( A1 => n21507, A2 => n19434, ZN => n21508);
   U28279 : NAND2_X1 port map( A1 => n21476, A2 => n19543, ZN => n21519);
   U28280 : NAND2_X1 port map( A1 => n1157, A2 => n39192, ZN => n21532);
   U28282 : MUX2_X1 port map( I0 => n21532, I1 => n21531, S => n18417, Z => 
                           n21534);
   U28283 : NAND2_X1 port map( A1 => n21539, A2 => n21699, ZN => n21540);
   U28285 : OAI22_X1 port map( A1 => n21872, A2 => n21756, B1 => n21546, B2 => 
                           n19337, ZN => n21548);
   U28286 : NAND2_X1 port map( A1 => n21696, A2 => n21695, ZN => n21547);
   U28287 : OAI21_X2 port map( A1 => n21549, A2 => n21548, B => n21547, ZN => 
                           n22047);
   U28288 : NAND2_X1 port map( A1 => n293, A2 => n21111, ZN => n21556);
   U28289 : NOR2_X1 port map( A1 => n21575, A2 => n21883, ZN => n21881);
   U28290 : OAI21_X2 port map( A1 => n21598, A2 => n21597, B => n21596, ZN => 
                           n22170);
   U28292 : NOR2_X1 port map( A1 => n21782, A2 => n35116, ZN => n21604);
   U28293 : NOR2_X1 port map( A1 => n4342, A2 => n15697, ZN => n21616);
   U28294 : INV_X1 port map( I => n21612, ZN => n21610);
   U28299 : AOI22_X1 port map( A1 => n21624, A2 => n21900, B1 => n21623, B2 => 
                           n21840, ZN => n21625);
   U28300 : OAI21_X1 port map( A1 => n21939, A2 => n19350, B => n21632, ZN => 
                           n21633);
   U28301 : NOR2_X1 port map( A1 => n16128, A2 => n21770, ZN => n21639);
   U28303 : NAND2_X1 port map( A1 => n21401, A2 => n39650, ZN => n21642);
   U28305 : NOR2_X1 port map( A1 => n21645, A2 => n21909, ZN => n21646);
   U28306 : OAI21_X1 port map( A1 => n21720, A2 => n21646, B => n21910, ZN => 
                           n21647);
   U28315 : NOR2_X1 port map( A1 => n21813, A2 => n21684, ZN => n21685);
   U28318 : NAND2_X1 port map( A1 => n21699, A2 => n19822, ZN => n21700);
   U28319 : MUX2_X1 port map( I0 => n21701, I1 => n21700, S => n21702, Z => 
                           n21705);
   U28320 : NAND2_X1 port map( A1 => n21886, A2 => n15338, ZN => n21706);
   U28321 : OAI21_X1 port map( A1 => n21748, A2 => n1157, B => n39192, ZN => 
                           n21711);
   U28322 : NAND2_X1 port map( A1 => n21711, A2 => n19542, ZN => n21717);
   U28323 : NOR2_X1 port map( A1 => n21748, A2 => n21712, ZN => n21714);
   U28325 : INV_X1 port map( I => n21732, ZN => n21733);
   U28326 : NAND2_X1 port map( A1 => n670, A2 => n21111, ZN => n21737);
   U28327 : OAI22_X1 port map( A1 => n21737, A2 => n18412, B1 => n21736, B2 => 
                           n19323, ZN => n21738);
   U28328 : NOR2_X1 port map( A1 => n1157, A2 => n19287, ZN => n21745);
   U28329 : MUX2_X1 port map( I0 => n694, I1 => n18266, S => n19416, Z => 
                           n21755);
   U28330 : NAND2_X1 port map( A1 => n21874, A2 => n21756, ZN => n21760);
   U28331 : NOR2_X1 port map( A1 => n1692, A2 => n19337, ZN => n21758);
   U28332 : NAND2_X1 port map( A1 => n21872, A2 => n21756, ZN => n21757);
   U28335 : NAND2_X1 port map( A1 => n20923, A2 => n32138, ZN => n21772);
   U28336 : MUX2_X1 port map( I0 => n21772, I1 => n21771, S => n21944, Z => 
                           n21773);
   U28339 : NAND2_X1 port map( A1 => n9759, A2 => n18205, ZN => n21793);
   U28340 : AOI21_X1 port map( A1 => n21794, A2 => n21793, B => n16945, ZN => 
                           n21795);
   U28341 : INV_X1 port map( I => n22034, ZN => n21799);
   U28342 : NOR2_X1 port map( A1 => n21799, A2 => n22246, ZN => n21800);
   U28343 : NAND2_X1 port map( A1 => n21980, A2 => n22300, ZN => n21801);
   U28344 : NAND2_X1 port map( A1 => n22039, A2 => n22038, ZN => n21803);
   U28346 : NAND2_X1 port map( A1 => n1345, A2 => n1693, ZN => n21809);
   U28347 : OAI21_X1 port map( A1 => n13632, A2 => n21816, B => n21815, ZN => 
                           n21829);
   U28348 : NAND2_X1 port map( A1 => n21821, A2 => n22146, ZN => n21827);
   U28350 : NAND2_X1 port map( A1 => n21830, A2 => n11344, ZN => n21831);
   U28354 : NOR2_X1 port map( A1 => n21857, A2 => n21861, ZN => n21859);
   U28355 : OAI21_X1 port map( A1 => n21862, A2 => n21861, B => n21860, ZN => 
                           n21863);
   U28356 : NAND2_X1 port map( A1 => n22241, A2 => n1047, ZN => n21865);
   U28357 : XOR2_X1 port map( A1 => n7055, A2 => n22528, Z => n21866);
   U28361 : AOI21_X1 port map( A1 => n21877, A2 => n19395, B => n21876, ZN => 
                           n21878);
   U28362 : NOR2_X1 port map( A1 => n2533, A2 => n21889, ZN => n21890);
   U28363 : NOR2_X1 port map( A1 => n19647, A2 => n21909, ZN => n21906);
   U28364 : NOR2_X1 port map( A1 => n21908, A2 => n21401, ZN => n21911);
   U28367 : NAND2_X1 port map( A1 => n32164, A2 => n20003, ZN => n21931);
   U28368 : NOR2_X1 port map( A1 => n14769, A2 => n20003, ZN => n21934);
   U28369 : OAI21_X1 port map( A1 => n6722, A2 => n22130, B => n22282, ZN => 
                           n21957);
   U28370 : INV_X1 port map( I => n21945, ZN => n21947);
   U28371 : NAND2_X2 port map( A1 => n21953, A2 => n21952, ZN => n22281);
   U28372 : NOR2_X1 port map( A1 => n22282, A2 => n19486, ZN => n21954);
   U28374 : INV_X1 port map( I => n21963, ZN => n21960);
   U28375 : NAND2_X1 port map( A1 => n22281, A2 => n22189, ZN => n21964);
   U28378 : NOR2_X1 port map( A1 => n22344, A2 => n22342, ZN => n21986);
   U28380 : NAND3_X1 port map( A1 => n19471, A2 => n21990, A3 => n32313, ZN => 
                           n21993);
   U28381 : NAND3_X1 port map( A1 => n22265, A2 => n33623, A3 => n22266, ZN => 
                           n21998);
   U28382 : NOR2_X1 port map( A1 => n32259, A2 => n22267, ZN => n21997);
   U28383 : INV_X1 port map( I => n22644, ZN => n21999);
   U28385 : XOR2_X1 port map( A1 => n22002, A2 => n22001, Z => n22003);
   U28389 : NAND3_X1 port map( A1 => n22204, A2 => n9685, A3 => n19837, ZN => 
                           n22013);
   U28391 : NAND2_X1 port map( A1 => n9736, A2 => n22100, ZN => n22060);
   U28392 : NOR2_X1 port map( A1 => n22268, A2 => n22266, ZN => n22072);
   U28393 : OAI21_X1 port map( A1 => n22140, A2 => n18854, B => n9265, ZN => 
                           n22078);
   U28394 : NOR2_X1 port map( A1 => n22246, A2 => n37938, ZN => n22077);
   U28395 : NAND2_X1 port map( A1 => n19471, A2 => n14139, ZN => n22081);
   U28396 : XOR2_X1 port map( A1 => n22583, A2 => n29562, Z => n22082);
   U28398 : NOR2_X1 port map( A1 => n22356, A2 => n22353, ZN => n22093);
   U28399 : NAND2_X1 port map( A1 => n22334, A2 => n22100, ZN => n22099);
   U28401 : NAND2_X1 port map( A1 => n22172, A2 => n19873, ZN => n22106);
   U28402 : NOR2_X1 port map( A1 => n22108, A2 => n22184, ZN => n22110);
   U28403 : NAND2_X1 port map( A1 => n1049, A2 => n1334, ZN => n22115);
   U28404 : NAND3_X1 port map( A1 => n22118, A2 => n22117, A3 => n22116, ZN => 
                           n22121);
   U28405 : INV_X1 port map( I => n22119, ZN => n22120);
   U28406 : OAI22_X1 port map( A1 => n22265, A2 => n22122, B1 => n22121, B2 => 
                           n22120, ZN => n22123);
   U28411 : NAND2_X1 port map( A1 => n22985, A2 => n35288, ZN => n22168);
   U28412 : NAND3_X1 port map( A1 => n22225, A2 => n35618, A3 => n22365, ZN => 
                           n22159);
   U28414 : NOR2_X1 port map( A1 => n22165, A2 => n196, ZN => n22166);
   U28415 : XOR2_X1 port map( A1 => n22485, A2 => n29399, Z => n22167);
   U28417 : XOR2_X1 port map( A1 => n22610, A2 => n31576, Z => n22195);
   U28418 : NOR2_X1 port map( A1 => n22282, A2 => n22281, ZN => n22192);
   U28419 : XOR2_X1 port map( A1 => n22459, A2 => n3953, Z => n22201);
   U28423 : NAND2_X1 port map( A1 => n22216, A2 => n9938, ZN => n22217);
   U28424 : XOR2_X1 port map( A1 => n22439, A2 => n28910, Z => n22231);
   U28425 : XOR2_X1 port map( A1 => n22452, A2 => n22231, Z => n22232);
   U28427 : XOR2_X1 port map( A1 => n22391, A2 => n22761, Z => n22279);
   U28430 : MUX2_X1 port map( I0 => n22309, I1 => n22308, S => n14024, Z => 
                           n22312);
   U28431 : NAND3_X1 port map( A1 => n1335, A2 => n22310, A3 => n31651, ZN => 
                           n22311);
   U28433 : XOR2_X1 port map( A1 => n22634, A2 => n29805, Z => n22370);
   U28434 : INV_X1 port map( I => n22376, ZN => n22374);
   U28435 : INV_X1 port map( I => n22375, ZN => n22373);
   U28436 : NAND3_X1 port map( A1 => n22374, A2 => n18270, A3 => n22373, ZN => 
                           n22378);
   U28437 : OAI21_X1 port map( A1 => n22376, A2 => n22375, B => n23591, ZN => 
                           n22377);
   U28438 : NAND2_X1 port map( A1 => n22378, A2 => n22377, ZN => n22379);
   U28439 : XOR2_X1 port map( A1 => n359, A2 => n30114, Z => n22383);
   U28440 : XOR2_X1 port map( A1 => n22729, A2 => n22749, Z => n22384);
   U28441 : XOR2_X1 port map( A1 => n22567, A2 => n22384, Z => n22385);
   U28442 : XOR2_X1 port map( A1 => n22715, A2 => n29206, Z => n22393);
   U28444 : XOR2_X1 port map( A1 => n34678, A2 => n19875, Z => n22394);
   U28447 : INV_X1 port map( I => n22398, ZN => n22404);
   U28448 : OAI22_X1 port map( A1 => n22404, A2 => n22403, B1 => n22402, B2 => 
                           n22401, ZN => n22405);
   U28449 : NAND3_X1 port map( A1 => n23103, A2 => n23104, A3 => n903, ZN => 
                           n22407);
   U28450 : XOR2_X1 port map( A1 => n11541, A2 => n19825, Z => n22409);
   U28453 : XOR2_X1 port map( A1 => n22700, A2 => n22550, Z => n22415);
   U28454 : XOR2_X1 port map( A1 => n9874, A2 => n28821, Z => n22414);
   U28455 : XOR2_X1 port map( A1 => n9116, A2 => n19874, Z => n22417);
   U28456 : XOR2_X1 port map( A1 => n16226, A2 => n19721, Z => n22418);
   U28458 : XOR2_X1 port map( A1 => n31863, A2 => n30950, Z => n22422);
   U28459 : XOR2_X1 port map( A1 => n22422, A2 => n22755, Z => n22425);
   U28462 : XOR2_X1 port map( A1 => n31576, A2 => n22563, Z => n22426);
   U28464 : XOR2_X1 port map( A1 => n22566, A2 => n21215, Z => n22431);
   U28465 : XOR2_X1 port map( A1 => n22432, A2 => n22431, Z => n22433);
   U28466 : XOR2_X1 port map( A1 => n34678, A2 => n29319, Z => n22436);
   U28467 : XOR2_X1 port map( A1 => n39804, A2 => n29003, Z => n22442);
   U28468 : XOR2_X1 port map( A1 => n36596, A2 => n19903, Z => n22446);
   U28469 : XOR2_X1 port map( A1 => n22643, A2 => n22763, Z => n22451);
   U28472 : XOR2_X1 port map( A1 => n22509, A2 => n19774, Z => n22469);
   U28473 : XOR2_X1 port map( A1 => n18568, A2 => n22580, Z => n22470);
   U28477 : XOR2_X1 port map( A1 => n31339, A2 => n9874, Z => n22474);
   U28478 : XOR2_X1 port map( A1 => n39682, A2 => n19947, Z => n22478);
   U28479 : XOR2_X1 port map( A1 => n9982, A2 => n19897, Z => n22487);
   U28481 : XOR2_X1 port map( A1 => n22575, A2 => n19624, Z => n22494);
   U28482 : MUX2_X1 port map( I0 => n22496, I1 => n36245, S => n20376, Z => 
                           n22498);
   U28483 : XOR2_X1 port map( A1 => n15439, A2 => n29442, Z => n22505);
   U28484 : XOR2_X1 port map( A1 => n34718, A2 => n22562, Z => n22519);
   U28485 : XOR2_X1 port map( A1 => n22583, A2 => n29801, Z => n22521);
   U28486 : XOR2_X1 port map( A1 => n22522, A2 => n22521, Z => n22523);
   U28487 : NAND2_X1 port map( A1 => n15770, A2 => n22890, ZN => n22526);
   U28490 : XOR2_X1 port map( A1 => n37428, A2 => n22582, Z => n22537);
   U28491 : XOR2_X1 port map( A1 => n17195, A2 => n29964, Z => n22536);
   U28492 : XOR2_X1 port map( A1 => n22536, A2 => n22537, Z => n22538);
   U28494 : XOR2_X1 port map( A1 => n20294, A2 => n22544, Z => n22548);
   U28495 : XOR2_X1 port map( A1 => n22546, A2 => n22545, Z => n22547);
   U28496 : XOR2_X1 port map( A1 => n22548, A2 => n22547, Z => n22853);
   U28498 : NAND2_X1 port map( A1 => n19288, A2 => n22928, ZN => n22558);
   U28499 : XOR2_X1 port map( A1 => n22647, A2 => n22621, Z => n22560);
   U28500 : XOR2_X1 port map( A1 => n22610, A2 => n19887, Z => n22564);
   U28503 : XOR2_X1 port map( A1 => n35920, A2 => n19622, Z => n22576);
   U28504 : XOR2_X1 port map( A1 => n22668, A2 => n14309, Z => n22579);
   U28505 : XOR2_X1 port map( A1 => n16798, A2 => n22582, Z => n22584);
   U28507 : XOR2_X1 port map( A1 => n22601, A2 => n2383, Z => n22602);
   U28508 : XOR2_X1 port map( A1 => n36867, A2 => n22610, Z => n22611);
   U28509 : XOR2_X1 port map( A1 => n39804, A2 => n19722, Z => n22613);
   U28510 : XOR2_X1 port map( A1 => n38330, A2 => n19933, Z => n22617);
   U28511 : XOR2_X1 port map( A1 => n19094, A2 => n19894, Z => n22618);
   U28512 : XOR2_X1 port map( A1 => n22629, A2 => n22749, Z => n22630);
   U28514 : XOR2_X1 port map( A1 => n22634, A2 => n19833, Z => n22636);
   U28515 : XOR2_X1 port map( A1 => n39682, A2 => n19913, Z => n22641);
   U28516 : XOR2_X1 port map( A1 => n22645, A2 => n19808, Z => n22646);
   U28517 : XOR2_X1 port map( A1 => n22648, A2 => n29554, Z => n22649);
   U28518 : XOR2_X1 port map( A1 => n17195, A2 => n29538, Z => n22653);
   U28519 : XOR2_X1 port map( A1 => n22659, A2 => n19820, Z => n22660);
   U28520 : XOR2_X1 port map( A1 => n22671, A2 => n22670, Z => n22673);
   U28524 : XOR2_X1 port map( A1 => n3475, A2 => n19910, Z => n22704);
   U28527 : NAND2_X1 port map( A1 => n23012, A2 => n33972, ZN => n22708);
   U28528 : XOR2_X1 port map( A1 => n22715, A2 => n30016, Z => n22716);
   U28529 : XOR2_X1 port map( A1 => n22717, A2 => n22716, Z => n22718);
   U28530 : XOR2_X1 port map( A1 => n22718, A2 => n22719, Z => n23140);
   U28532 : XOR2_X1 port map( A1 => n22778, A2 => n22761, Z => n22726);
   U28533 : XOR2_X1 port map( A1 => n22724, A2 => n19758, Z => n22725);
   U28534 : XOR2_X1 port map( A1 => n22726, A2 => n22725, Z => n22727);
   U28535 : XOR2_X1 port map( A1 => n35559, A2 => n19780, Z => n22734);
   U28537 : XOR2_X1 port map( A1 => n1657, A2 => n30094, Z => n22737);
   U28540 : NAND2_X1 port map( A1 => n23034, A2 => n4682, ZN => n22746);
   U28541 : XOR2_X1 port map( A1 => n38838, A2 => n29463, Z => n22751);
   U28542 : XOR2_X1 port map( A1 => n22752, A2 => n22751, Z => n22753);
   U28544 : XOR2_X1 port map( A1 => n22763, A2 => n19817, Z => n22764);
   U28545 : XOR2_X1 port map( A1 => n22766, A2 => n29476, Z => n22768);
   U28549 : XOR2_X1 port map( A1 => n39682, A2 => n19831, Z => n22782);
   U28552 : NAND2_X1 port map( A1 => n9050, A2 => n59, ZN => n22797);
   U28554 : OAI21_X1 port map( A1 => n22903, A2 => n906, B => n20872, ZN => 
                           n22815);
   U28555 : NAND2_X1 port map( A1 => n19307, A2 => n23028, ZN => n22817);
   U28560 : NAND3_X1 port map( A1 => n23149, A2 => n31838, A3 => n14556, ZN => 
                           n22831);
   U28563 : NAND3_X1 port map( A1 => n5702, A2 => n4573, A3 => n22931, ZN => 
                           n22846);
   U28564 : NAND2_X1 port map( A1 => n31906, A2 => n17090, ZN => n22852);
   U28566 : NOR2_X1 port map( A1 => n22875, A2 => n19840, ZN => n22876);
   U28567 : INV_X1 port map( I => n23123, ZN => n22877);
   U28568 : OAI21_X1 port map( A1 => n45, A2 => n23034, B => n35994, ZN => 
                           n22881);
   U28569 : NOR2_X1 port map( A1 => n38173, A2 => n1642, ZN => n22911);
   U28573 : NOR2_X1 port map( A1 => n23189, A2 => n23188, ZN => n22977);
   U28574 : NAND2_X1 port map( A1 => n34419, A2 => n23188, ZN => n22978);
   U28580 : NAND2_X1 port map( A1 => n36829, A2 => n23456, ZN => n22986);
   U28581 : NAND2_X1 port map( A1 => n18762, A2 => n30574, ZN => n22988);
   U28585 : MUX2_X1 port map( I0 => n23071, I1 => n23005, S => n5976, Z => 
                           n23006);
   U28587 : INV_X1 port map( I => n23479, ZN => n23017);
   U28590 : INV_X1 port map( I => n121, ZN => n23026);
   U28593 : NAND2_X1 port map( A1 => n18284, A2 => n23458, ZN => n23040);
   U28595 : NAND2_X1 port map( A1 => n23045, A2 => n11658, ZN => n23046);
   U28596 : NAND2_X1 port map( A1 => n9854, A2 => n38542, ZN => n23049);
   U28597 : NAND2_X1 port map( A1 => n33817, A2 => n23159, ZN => n23050);
   U28598 : INV_X1 port map( I => n23054, ZN => n23055);
   U28607 : NOR2_X1 port map( A1 => n14556, A2 => n31838, ZN => n23151);
   U28608 : NAND2_X1 port map( A1 => n16963, A2 => n36095, ZN => n23431);
   U28610 : AOI21_X1 port map( A1 => n38524, A2 => n23189, B => n23188, ZN => 
                           n23193);
   U28613 : XOR2_X1 port map( A1 => n19649, A2 => n23911, Z => n23220);
   U28615 : NAND3_X1 port map( A1 => n32351, A2 => n17556, A3 => n31644, ZN => 
                           n23218);
   U28617 : NAND2_X1 port map( A1 => n23277, A2 => n1629, ZN => n23228);
   U28620 : NAND3_X1 port map( A1 => n23462, A2 => n23458, A3 => n5083, ZN => 
                           n23240);
   U28621 : NAND2_X1 port map( A1 => n23420, A2 => n23602, ZN => n23252);
   U28624 : NAND2_X1 port map( A1 => n39001, A2 => n10024, ZN => n23267);
   U28625 : NAND2_X1 port map( A1 => n12093, A2 => n32158, ZN => n23271);
   U28626 : NAND2_X1 port map( A1 => n31332, A2 => n23539, ZN => n23276);
   U28627 : MUX2_X1 port map( I0 => n23534, I1 => n23276, S => n23538, Z => 
                           n23279);
   U28628 : XOR2_X1 port map( A1 => n23846, A2 => n29983, Z => n23280);
   U28633 : NAND3_X1 port map( A1 => n23450, A2 => n38173, A3 => n1642, ZN => 
                           n23291);
   U28635 : NAND2_X1 port map( A1 => n18762, A2 => n31586, ZN => n23295);
   U28636 : NAND2_X1 port map( A1 => n1135, A2 => n23293, ZN => n23294);
   U28639 : XOR2_X1 port map( A1 => n23783, A2 => n29879, Z => n23330);
   U28646 : OAI21_X1 port map( A1 => n39214, A2 => n7485, B => n23367, ZN => 
                           n23368);
   U28649 : NAND2_X1 port map( A1 => n39300, A2 => n23502, ZN => n23375);
   U28650 : XOR2_X1 port map( A1 => n33452, A2 => n19735, Z => n23378);
   U28651 : XOR2_X1 port map( A1 => n32122, A2 => n17462, Z => n23382);
   U28653 : INV_X1 port map( I => n23548, ZN => n23386);
   U28659 : NOR2_X1 port map( A1 => n30499, A2 => n23401, ZN => n23403);
   U28660 : XOR2_X1 port map( A1 => n23888, A2 => n29666, Z => n23409);
   U28661 : XOR2_X1 port map( A1 => n23734, A2 => n23409, Z => n23410);
   U28664 : XOR2_X1 port map( A1 => n23755, A2 => n29808, Z => n23428);
   U28665 : NAND3_X1 port map( A1 => n33287, A2 => n31661, A3 => n32930, ZN => 
                           n23427);
   U28666 : XOR2_X1 port map( A1 => n23717, A2 => n23428, Z => n23429);
   U28667 : AOI21_X1 port map( A1 => n1628, A2 => n3496, B => n23624, ZN => 
                           n23435);
   U28671 : NAND3_X1 port map( A1 => n23484, A2 => n23483, A3 => n9078, ZN => 
                           n23485);
   U28672 : NAND2_X1 port map( A1 => n23251, A2 => n23496, ZN => n23494);
   U28675 : NAND4_X1 port map( A1 => n23511, A2 => n11245, A3 => n23510, A4 => 
                           n23509, ZN => n23512);
   U28677 : XOR2_X1 port map( A1 => n19608, A2 => n30179, Z => n23549);
   U28678 : NAND2_X1 port map( A1 => n23583, A2 => n23582, ZN => n23584);
   U28680 : NOR2_X1 port map( A1 => n12597, A2 => n23602, ZN => n23603);
   U28683 : NAND2_X1 port map( A1 => n35506, A2 => n13305, ZN => n23630);
   U28685 : XOR2_X1 port map( A1 => n32122, A2 => n29831, Z => n23649);
   U28686 : XOR2_X1 port map( A1 => n24070, A2 => n19804, Z => n23653);
   U28687 : XOR2_X1 port map( A1 => n23886, A2 => n19527, Z => n23656);
   U28690 : XOR2_X1 port map( A1 => n24017, A2 => n23665, Z => n23666);
   U28691 : XOR2_X1 port map( A1 => n23955, A2 => n19913, Z => n23668);
   U28692 : XOR2_X1 port map( A1 => n24025, A2 => n19817, Z => n23672);
   U28694 : XOR2_X1 port map( A1 => n238, A2 => n29801, Z => n23687);
   U28695 : XOR2_X1 port map( A1 => n18279, A2 => n29325, Z => n23689);
   U28696 : XOR2_X1 port map( A1 => n18310, A2 => n23728, Z => n23692);
   U28698 : XOR2_X1 port map( A1 => n23698, A2 => n28910, Z => n23699);
   U28701 : XOR2_X1 port map( A1 => n24005, A2 => n19592, Z => n23713);
   U28702 : XOR2_X1 port map( A1 => n24077, A2 => n29474, Z => n23719);
   U28705 : XOR2_X1 port map( A1 => n35942, A2 => n29538, Z => n23727);
   U28706 : XOR2_X1 port map( A1 => n1617, A2 => n23728, Z => n23813);
   U28707 : INV_X1 port map( I => n24079, ZN => n23792);
   U28709 : XOR2_X1 port map( A1 => n23769, A2 => n19583, Z => n23733);
   U28710 : XOR2_X1 port map( A1 => n23884, A2 => n29707, Z => n23738);
   U28712 : INV_X1 port map( I => n23972, ZN => n23742);
   U28714 : INV_X1 port map( I => n23746, ZN => n23747);
   U28715 : INV_X1 port map( I => n23748, ZN => n23750);
   U28716 : NAND2_X1 port map( A1 => n23750, A2 => n23749, ZN => n23751);
   U28717 : XOR2_X1 port map( A1 => n23757, A2 => n23814, Z => n23758);
   U28718 : XOR2_X1 port map( A1 => n23850, A2 => n23759, Z => n23760);
   U28719 : XOR2_X1 port map( A1 => n23808, A2 => n19877, Z => n23763);
   U28720 : NAND4_X1 port map( A1 => n23767, A2 => n23766, A3 => n23796, A4 => 
                           n23765, ZN => n23768);
   U28721 : XOR2_X1 port map( A1 => n23769, A2 => n29442, Z => n23770);
   U28722 : XOR2_X1 port map( A1 => n23771, A2 => n23770, Z => n23772);
   U28723 : XOR2_X1 port map( A1 => n23933, A2 => n35942, Z => n23795);
   U28724 : MUX2_X1 port map( I0 => n9822, I1 => n23799, S => n1125, Z => 
                           n23800);
   U28725 : XOR2_X1 port map( A1 => n39209, A2 => n33866, Z => n23803);
   U28728 : NAND2_X1 port map( A1 => n9844, A2 => n12771, ZN => n23821);
   U28729 : OR2_X1 port map( A1 => n23821, A2 => n11265, Z => n23822);
   U28731 : NAND2_X1 port map( A1 => n545, A2 => n19915, ZN => n23828);
   U28732 : XOR2_X1 port map( A1 => n23851, A2 => n30016, Z => n23834);
   U28733 : XOR2_X1 port map( A1 => n35561, A2 => n19831, Z => n23836);
   U28734 : NOR2_X1 port map( A1 => n19880, A2 => n39467, ZN => n23845);
   U28735 : INV_X1 port map( I => n24061, ZN => n23838);
   U28736 : XOR2_X1 port map( A1 => n23866, A2 => n23842, Z => n23843);
   U28738 : XOR2_X1 port map( A1 => n23846, A2 => n29238, Z => n23847);
   U28739 : XOR2_X1 port map( A1 => n23890, A2 => n19952, Z => n23849);
   U28740 : XOR2_X1 port map( A1 => n19608, A2 => n29206, Z => n23853);
   U28742 : XOR2_X1 port map( A1 => n23861, A2 => n19839, Z => n23862);
   U28743 : XOR2_X1 port map( A1 => n23863, A2 => n23862, Z => n23864);
   U28744 : XOR2_X1 port map( A1 => n33452, A2 => n35702, Z => n23867);
   U28745 : XOR2_X1 port map( A1 => n24075, A2 => n29221, Z => n23870);
   U28748 : XOR2_X1 port map( A1 => n23970, A2 => n19866, Z => n23879);
   U28749 : XOR2_X1 port map( A1 => n24077, A2 => n33672, Z => n24014);
   U28751 : XOR2_X1 port map( A1 => n23988, A2 => n23893, Z => n23925);
   U28752 : XOR2_X1 port map( A1 => n23894, A2 => n19736, Z => n23895);
   U28753 : XOR2_X1 port map( A1 => n23925, A2 => n23895, Z => n23896);
   U28754 : XOR2_X1 port map( A1 => n23897, A2 => n23896, Z => n23907);
   U28756 : XOR2_X1 port map( A1 => n23900, A2 => n30170, Z => n23901);
   U28757 : XOR2_X1 port map( A1 => n23905, A2 => n29319, Z => n23906);
   U28760 : XOR2_X1 port map( A1 => n23609, A2 => n29689, Z => n23927);
   U28761 : XOR2_X1 port map( A1 => n23944, A2 => n23945, Z => n23949);
   U28762 : XOR2_X1 port map( A1 => n23609, A2 => n19780, Z => n23946);
   U28764 : XOR2_X1 port map( A1 => n23973, A2 => n19908, Z => n23974);
   U28765 : XOR2_X1 port map( A1 => n23976, A2 => n29602, Z => n23977);
   U28766 : MUX2_X1 port map( I0 => n24444, I1 => n23983, S => n24311, Z => 
                           n23994);
   U28769 : XOR2_X1 port map( A1 => n23988, A2 => n23987, Z => n23989);
   U28770 : XOR2_X1 port map( A1 => n23989, A2 => n20594, Z => n23990);
   U28771 : XOR2_X1 port map( A1 => n23991, A2 => n23990, Z => n24420);
   U28776 : XOR2_X1 port map( A1 => n24030, A2 => n19885, Z => n24032);
   U28777 : XOR2_X1 port map( A1 => n24036, A2 => n6561, Z => n24037);
   U28779 : XOR2_X1 port map( A1 => n30321, A2 => n19721, Z => n24042);
   U28780 : XOR2_X1 port map( A1 => n24047, A2 => n29295, Z => n24048);
   U28781 : XOR2_X1 port map( A1 => n24052, A2 => n19616, Z => n24054);
   U28782 : INV_X1 port map( I => n24133, ZN => n24072);
   U28783 : XOR2_X1 port map( A1 => n24076, A2 => n29363, Z => n24078);
   U28787 : NOR3_X1 port map( A1 => n16917, A2 => n24311, A3 => n253, ZN => 
                           n24091);
   U28790 : MUX2_X1 port map( I0 => n277, I1 => n24398, S => n24396, Z => 
                           n24105);
   U28791 : INV_X1 port map( I => n19880, ZN => n24170);
   U28792 : NAND2_X1 port map( A1 => n24105, A2 => n24170, ZN => n24109);
   U28794 : NOR2_X1 port map( A1 => n24168, A2 => n24395, ZN => n24107);
   U28797 : INV_X1 port map( I => n24410, ZN => n24111);
   U28798 : INV_X1 port map( I => n24161, ZN => n24117);
   U28802 : MUX2_X1 port map( I0 => n24129, I1 => n24157, S => n13653, Z => 
                           n24131);
   U28805 : NAND2_X1 port map( A1 => n24271, A2 => n18697, ZN => n24148);
   U28806 : XOR2_X1 port map( A1 => n38714, A2 => n19648, Z => n24150);
   U28807 : NOR2_X1 port map( A1 => n6849, A2 => n20537, ZN => n24163);
   U28808 : OAI21_X1 port map( A1 => n19942, A2 => n30897, B => n802, ZN => 
                           n24193);
   U28809 : NAND2_X1 port map( A1 => n35890, A2 => n31452, ZN => n24194);
   U28813 : NAND2_X1 port map( A1 => n24221, A2 => n6839, ZN => n24222);
   U28823 : NAND3_X1 port map( A1 => n19745, A2 => n24267, A3 => n24266, ZN => 
                           n24268);
   U28827 : NAND2_X1 port map( A1 => n24300, A2 => n37045, ZN => n24298);
   U28828 : NOR2_X1 port map( A1 => n37267, A2 => n24463, ZN => n24302);
   U28831 : NAND2_X1 port map( A1 => n24419, A2 => n24311, ZN => n24312);
   U28835 : XOR2_X1 port map( A1 => n19817, A2 => n25086, Z => n24325);
   U28836 : NAND4_X1 port map( A1 => n24342, A2 => n24341, A3 => n24339, A4 => 
                           n24340, ZN => n24343);
   U28838 : NOR2_X1 port map( A1 => n36082, A2 => n4008, ZN => n24363);
   U28840 : NAND3_X1 port map( A1 => n14167, A2 => n24818, A3 => n24824, ZN => 
                           n24388);
   U28841 : NAND2_X1 port map( A1 => n24392, A2 => n1283, ZN => n24393);
   U28845 : XOR2_X1 port map( A1 => n39756, A2 => n19761, Z => n24436);
   U28846 : NAND2_X1 port map( A1 => n24606, A2 => n20696, ZN => n24437);
   U28848 : NAND2_X1 port map( A1 => n14491, A2 => n24449, ZN => n24452);
   U28850 : MUX2_X1 port map( I0 => n24452, I1 => n24451, S => n17871, Z => 
                           n24456);
   U28856 : NAND2_X1 port map( A1 => n34123, A2 => n31684, ZN => n24498);
   U28858 : NOR2_X1 port map( A1 => n24876, A2 => n1580, ZN => n24504);
   U28862 : INV_X1 port map( I => n24530, ZN => n24531);
   U28866 : XOR2_X1 port map( A1 => n24944, A2 => n30248, Z => n24541);
   U28867 : XOR2_X1 port map( A1 => n24542, A2 => n24541, Z => n24543);
   U28868 : XOR2_X1 port map( A1 => n24544, A2 => n24543, Z => n25395);
   U28869 : XOR2_X1 port map( A1 => n9701, A2 => n24942, Z => n24551);
   U28871 : XOR2_X1 port map( A1 => n25218, A2 => n29689, Z => n24550);
   U28872 : XOR2_X1 port map( A1 => n24551, A2 => n24550, Z => n24552);
   U28875 : XOR2_X1 port map( A1 => n17184, A2 => n28910, Z => n24563);
   U28879 : NAND2_X1 port map( A1 => n18788, A2 => n24753, ZN => n24577);
   U28882 : NAND4_X1 port map( A1 => n24585, A2 => n24584, A3 => n24583, A4 => 
                           n24582, ZN => n24586);
   U28888 : INV_X1 port map( I => n24625, ZN => n24626);
   U28889 : XOR2_X1 port map( A1 => n1260, A2 => n19583, Z => n24632);
   U28891 : XOR2_X1 port map( A1 => n25247, A2 => n25280, Z => n24641);
   U28898 : XOR2_X1 port map( A1 => n24678, A2 => n19816, Z => n24679);
   U28899 : INV_X1 port map( I => n24687, ZN => n24690);
   U28900 : XOR2_X1 port map( A1 => n10792, A2 => n18991, Z => n24697);
   U28901 : NAND2_X1 port map( A1 => n16502, A2 => n7769, ZN => n24705);
   U28902 : AOI21_X1 port map( A1 => n24723, A2 => n5056, B => n24721, ZN => 
                           n24725);
   U28904 : XOR2_X1 port map( A1 => n38581, A2 => n25071, Z => n24801);
   U28905 : NOR2_X1 port map( A1 => n14939, A2 => n19868, ZN => n24815);
   U28906 : NOR3_X1 port map( A1 => n24821, A2 => n24820, A3 => n7529, ZN => 
                           n24822);
   U28910 : INV_X1 port map( I => n24843, ZN => n24844);
   U28911 : NAND2_X1 port map( A1 => n24844, A2 => n4973, ZN => n24845);
   U28915 : XOR2_X1 port map( A1 => n24857, A2 => n24858, Z => n24859);
   U28916 : XOR2_X1 port map( A1 => n25030, A2 => n18270, Z => n24860);
   U28917 : MUX2_X1 port map( I0 => n37477, I1 => n24869, S => n19901, Z => 
                           n24871);
   U28919 : NAND2_X1 port map( A1 => n24885, A2 => n24884, ZN => n24886);
   U28920 : XOR2_X1 port map( A1 => n25113, A2 => n19801, Z => n24891);
   U28922 : INV_X1 port map( I => n24904, ZN => n24905);
   U28923 : XOR2_X1 port map( A1 => n6727, A2 => n19763, Z => n24913);
   U28924 : XOR2_X1 port map( A1 => n24914, A2 => n24913, Z => n24915);
   U28925 : XOR2_X1 port map( A1 => n25085, A2 => n29978, Z => n24918);
   U28926 : XOR2_X1 port map( A1 => n38950, A2 => n19890, Z => n24919);
   U28927 : XOR2_X1 port map( A1 => n16627, A2 => n19732, Z => n24923);
   U28929 : XOR2_X1 port map( A1 => n16864, A2 => n29970, Z => n24940);
   U28930 : XOR2_X1 port map( A1 => n25232, A2 => n24940, Z => n24941);
   U28931 : XOR2_X1 port map( A1 => n25238, A2 => n29875, Z => n24945);
   U28933 : XOR2_X1 port map( A1 => n25226, A2 => n19774, Z => n24947);
   U28935 : XOR2_X1 port map( A1 => n24953, A2 => n24952, Z => n24954);
   U28936 : XOR2_X1 port map( A1 => n24955, A2 => n24954, Z => n25157);
   U28938 : XOR2_X1 port map( A1 => n25203, A2 => n29887, Z => n24960);
   U28939 : XOR2_X1 port map( A1 => n10792, A2 => n29363, Z => n24966);
   U28940 : OAI21_X2 port map( A1 => n24968, A2 => n24967, B => n19574, ZN => 
                           n26388);
   U28941 : XOR2_X1 port map( A1 => n25215, A2 => n19883, Z => n24971);
   U28942 : XOR2_X1 port map( A1 => n24972, A2 => n24971, Z => n24973);
   U28943 : XOR2_X1 port map( A1 => n25218, A2 => n29983, Z => n24975);
   U28944 : XOR2_X1 port map( A1 => n24976, A2 => n24975, Z => n24977);
   U28949 : XOR2_X1 port map( A1 => n25026, A2 => n30150, Z => n24988);
   U28950 : XOR2_X1 port map( A1 => n39146, A2 => n32195, Z => n24989);
   U28951 : XOR2_X1 port map( A1 => n25167, A2 => n24989, Z => n24990);
   U28952 : INV_X1 port map( I => n25546, ZN => n25482);
   U28953 : XOR2_X1 port map( A1 => n24991, A2 => n19721, Z => n24992);
   U28954 : XOR2_X1 port map( A1 => n25237, A2 => n5208, Z => n25004);
   U28955 : XOR2_X1 port map( A1 => n33208, A2 => n25090, Z => n25005);
   U28956 : MUX2_X1 port map( I0 => n31580, I1 => n12825, S => n18704, Z => 
                           n25012);
   U28957 : XOR2_X1 port map( A1 => n25014, A2 => n19903, Z => n25015);
   U28959 : INV_X1 port map( I => n25018, ZN => n25020);
   U28960 : NOR3_X1 port map( A1 => n25020, A2 => n38631, A3 => n25019, ZN => 
                           n25021);
   U28961 : XOR2_X1 port map( A1 => n25104, A2 => n30114, Z => n25023);
   U28962 : XOR2_X1 port map( A1 => n25024, A2 => n30104, Z => n25025);
   U28963 : XOR2_X1 port map( A1 => n25026, A2 => n19866, Z => n25027);
   U28964 : XOR2_X1 port map( A1 => n25226, A2 => n19839, Z => n25034);
   U28965 : NOR2_X1 port map( A1 => n34010, A2 => n25307, ZN => n25036);
   U28966 : XOR2_X1 port map( A1 => n39491, A2 => n29506, Z => n25041);
   U28967 : INV_X1 port map( I => n25047, ZN => n25051);
   U28968 : AOI22_X1 port map( A1 => n25051, A2 => n36634, B1 => n32488, B2 => 
                           n25049, ZN => n25056);
   U28969 : INV_X1 port map( I => n25052, ZN => n25054);
   U28970 : NAND2_X1 port map( A1 => n25054, A2 => n25053, ZN => n25055);
   U28972 : XOR2_X1 port map( A1 => n25259, A2 => n19407, Z => n25059);
   U28973 : XOR2_X1 port map( A1 => n25060, A2 => n25059, Z => n25061);
   U28976 : XOR2_X1 port map( A1 => n36075, A2 => n29514, Z => n25064);
   U28977 : XOR2_X1 port map( A1 => n25326, A2 => n25064, Z => n25065);
   U28979 : NOR2_X1 port map( A1 => n21302, A2 => n955, ZN => n25073);
   U28980 : XOR2_X1 port map( A1 => n6185, A2 => n25175, Z => n25078);
   U28981 : XOR2_X1 port map( A1 => n25076, A2 => n29371, Z => n25077);
   U28983 : XOR2_X1 port map( A1 => n10199, A2 => n25090, Z => n25092);
   U28984 : XOR2_X1 port map( A1 => n35900, A2 => n19825, Z => n25094);
   U28985 : XOR2_X1 port map( A1 => n39491, A2 => n29357, Z => n25098);
   U28986 : XOR2_X1 port map( A1 => n25098, A2 => n25099, Z => n25101);
   U28987 : INV_X1 port map( I => n25106, ZN => n25582);
   U28991 : XOR2_X1 port map( A1 => n29680, A2 => n38665, Z => n25119);
   U28992 : XOR2_X1 port map( A1 => n25120, A2 => n25119, Z => n25121);
   U28994 : INV_X1 port map( I => n25123, ZN => n25125);
   U28995 : XOR2_X1 port map( A1 => n25283, A2 => n25149, Z => n25129);
   U28996 : XOR2_X1 port map( A1 => n25127, A2 => n19877, Z => n25128);
   U28998 : XOR2_X1 port map( A1 => n25155, A2 => n35996, Z => n25135);
   U28999 : XOR2_X1 port map( A1 => n25135, A2 => n25134, Z => n25139);
   U29000 : XOR2_X1 port map( A1 => n39756, A2 => n19738, Z => n25137);
   U29002 : XOR2_X1 port map( A1 => n30865, A2 => n33216, Z => n25187);
   U29003 : XOR2_X1 port map( A1 => n25189, A2 => n1561, Z => n25190);
   U29005 : XOR2_X1 port map( A1 => n35707, A2 => n30169, Z => n25207);
   U29006 : XOR2_X1 port map( A1 => n39491, A2 => n30203, Z => n25213);
   U29009 : XOR2_X1 port map( A1 => n25231, A2 => n25232, Z => n25236);
   U29010 : XOR2_X1 port map( A1 => n24417, A2 => n19860, Z => n25233);
   U29011 : XOR2_X1 port map( A1 => n25234, A2 => n25233, Z => n25235);
   U29012 : XOR2_X1 port map( A1 => n16900, A2 => n28968, Z => n25276);
   U29013 : XOR2_X1 port map( A1 => n25280, A2 => n30120, Z => n25281);
   U29014 : XOR2_X1 port map( A1 => n38714, A2 => n29522, Z => n25304);
   U29015 : XOR2_X1 port map( A1 => n39491, A2 => n29647, Z => n25320);
   U29016 : OAI21_X1 port map( A1 => n25552, A2 => n19478, B => n18704, ZN => 
                           n25336);
   U29019 : NOR2_X1 port map( A1 => n12533, A2 => n31509, ZN => n25341);
   U29023 : NAND2_X1 port map( A1 => n25352, A2 => n25386, ZN => n25354);
   U29025 : NAND3_X1 port map( A1 => n14410, A2 => n6731, A3 => n9132, ZN => 
                           n25358);
   U29027 : MUX2_X1 port map( I0 => n25371, I1 => n25370, S => n25886, Z => 
                           n25377);
   U29030 : NAND2_X1 port map( A1 => n25394, A2 => n19398, ZN => n25397);
   U29032 : XOR2_X1 port map( A1 => n3413, A2 => n29920, Z => n25407);
   U29036 : NAND2_X1 port map( A1 => n38183, A2 => n20614, ZN => n25425);
   U29038 : NAND3_X1 port map( A1 => n952, A2 => n15406, A3 => n17029, ZN => 
                           n25428);
   U29039 : NAND2_X1 port map( A1 => n8070, A2 => n1252, ZN => n25776);
   U29040 : NAND2_X1 port map( A1 => n25429, A2 => n33946, ZN => n25431);
   U29042 : INV_X1 port map( I => n25717, ZN => n25437);
   U29043 : NAND2_X1 port map( A1 => n25869, A2 => n18162, ZN => n25440);
   U29045 : NAND3_X1 port map( A1 => n25614, A2 => n36816, A3 => n25575, ZN => 
                           n25451);
   U29047 : NOR2_X1 port map( A1 => n1109, A2 => n25577, ZN => n25456);
   U29048 : OAI21_X1 port map( A1 => n12404, A2 => n25381, B => n1109, ZN => 
                           n25457);
   U29050 : NOR2_X1 port map( A1 => n25469, A2 => n1257, ZN => n25471);
   U29057 : NAND2_X1 port map( A1 => n19548, A2 => n4603, ZN => n25503);
   U29058 : NOR2_X1 port map( A1 => n26015, A2 => n25899, ZN => n25507);
   U29059 : NAND2_X1 port map( A1 => n25507, A2 => n1522, ZN => n25508);
   U29060 : XOR2_X1 port map( A1 => n26418, A2 => n19820, Z => n25511);
   U29067 : NAND2_X1 port map( A1 => n12825, A2 => n14602, ZN => n25549);
   U29069 : AOI21_X1 port map( A1 => n25554, A2 => n19581, B => n12825, ZN => 
                           n25555);
   U29070 : NOR3_X1 port map( A1 => n14410, A2 => n6731, A3 => n9132, ZN => 
                           n25560);
   U29075 : NOR2_X1 port map( A1 => n37553, A2 => n1552, ZN => n25592);
   U29076 : XOR2_X1 port map( A1 => n26532, A2 => n19613, Z => n25594);
   U29084 : NAND3_X1 port map( A1 => n20856, A2 => n14082, A3 => n25642, ZN => 
                           n25643);
   U29087 : NAND2_X1 port map( A1 => n20456, A2 => n36226, ZN => n25657);
   U29088 : NAND2_X1 port map( A1 => n30436, A2 => n3356, ZN => n25658);
   U29091 : NOR2_X1 port map( A1 => n25677, A2 => n25674, ZN => n25675);
   U29095 : NAND2_X1 port map( A1 => n25712, A2 => n8304, ZN => n25713);
   U29098 : MUX2_X1 port map( I0 => n25730, I1 => n25729, S => n5166, Z => 
                           n25731);
   U29099 : XOR2_X1 port map( A1 => n25734, A2 => n25735, Z => n25736);
   U29100 : NAND2_X1 port map( A1 => n9530, A2 => n19793, ZN => n25741);
   U29104 : NAND2_X1 port map( A1 => n11807, A2 => n25760, ZN => n25762);
   U29105 : NAND3_X1 port map( A1 => n9855, A2 => n37683, A3 => n1012, ZN => 
                           n25761);
   U29106 : INV_X1 port map( I => n25775, ZN => n25780);
   U29107 : NAND3_X1 port map( A1 => n25778, A2 => n25777, A3 => n25776, ZN => 
                           n25779);
   U29109 : NAND2_X1 port map( A1 => n25747, A2 => n26020, ZN => n25787);
   U29113 : AOI21_X1 port map( A1 => n25966, A2 => n25804, B => n25803, ZN => 
                           n25805);
   U29114 : INV_X1 port map( I => n26186, ZN => n25810);
   U29115 : NOR2_X1 port map( A1 => n25814, A2 => n25813, ZN => n25815);
   U29119 : NAND2_X1 port map( A1 => n25830, A2 => n31340, ZN => n25831);
   U29123 : NOR2_X1 port map( A1 => n34898, A2 => n26075, ZN => n25840);
   U29128 : NAND2_X1 port map( A1 => n1522, A2 => n1098, ZN => n25902);
   U29129 : NAND2_X1 port map( A1 => n26015, A2 => n25899, ZN => n25901);
   U29130 : MUX2_X1 port map( I0 => n25902, I1 => n25901, S => n33327, Z => 
                           n25907);
   U29134 : MUX2_X1 port map( I0 => n25911, I1 => n25910, S => n26004, Z => 
                           n25914);
   U29135 : XOR2_X1 port map( A1 => n5084, A2 => n29661, Z => n25930);
   U29137 : NOR3_X1 port map( A1 => n25345, A2 => n26063, A3 => n25941, ZN => 
                           n25942);
   U29138 : NAND3_X1 port map( A1 => n11807, A2 => n15283, A3 => n9883, ZN => 
                           n25950);
   U29139 : NAND3_X1 port map( A1 => n37683, A2 => n34898, A3 => n15283, ZN => 
                           n25949);
   U29141 : NAND2_X1 port map( A1 => n25961, A2 => n25965, ZN => n25964);
   U29144 : NAND2_X1 port map( A1 => n25966, A2 => n26028, ZN => n25967);
   U29146 : INV_X1 port map( I => n26034, ZN => n25982);
   U29149 : NOR2_X1 port map( A1 => n26237, A2 => n30883, ZN => n26036);
   U29150 : NOR2_X1 port map( A1 => n1100, A2 => n26034, ZN => n26239);
   U29151 : XOR2_X1 port map( A1 => n26259, A2 => n26548, Z => n26085);
   U29154 : XOR2_X1 port map( A1 => n26319, A2 => n30253, Z => n26141);
   U29155 : NOR2_X1 port map( A1 => n37524, A2 => n12066, ZN => n26149);
   U29156 : XOR2_X1 port map( A1 => n1502, A2 => n19780, Z => n26144);
   U29157 : XOR2_X1 port map( A1 => n26411, A2 => n26144, Z => n26147);
   U29159 : AOI21_X1 port map( A1 => n36262, A2 => n10902, B => n26151, ZN => 
                           n26152);
   U29161 : XOR2_X1 port map( A1 => n4622, A2 => n19947, Z => n26156);
   U29162 : XOR2_X1 port map( A1 => n2150, A2 => n19860, Z => n26162);
   U29163 : INV_X1 port map( I => n26995, ZN => n26878);
   U29164 : NAND2_X1 port map( A1 => n20981, A2 => n27081, ZN => n26195);
   U29165 : XOR2_X1 port map( A1 => n26568, A2 => n35202, Z => n26168);
   U29166 : XOR2_X1 port map( A1 => n38279, A2 => n26168, Z => n26171);
   U29168 : XOR2_X1 port map( A1 => n26568, A2 => n26231, Z => n26192);
   U29169 : XOR2_X1 port map( A1 => n38896, A2 => n18270, Z => n26191);
   U29170 : NAND2_X1 port map( A1 => n33254, A2 => n37201, ZN => n26196);
   U29172 : XOR2_X1 port map( A1 => n26198, A2 => n26567, Z => n26200);
   U29176 : XOR2_X1 port map( A1 => n26291, A2 => n29319, Z => n26206);
   U29177 : XOR2_X1 port map( A1 => n26531, A2 => n19534, Z => n26209);
   U29178 : NAND2_X1 port map( A1 => n26212, A2 => n5908, ZN => n26217);
   U29179 : NAND3_X1 port map( A1 => n9868, A2 => n26214, A3 => n26213, ZN => 
                           n26216);
   U29182 : XOR2_X1 port map( A1 => n26388, A2 => n30120, Z => n26232);
   U29185 : XOR2_X1 port map( A1 => n39129, A2 => n19616, Z => n26243);
   U29186 : MUX2_X1 port map( I0 => n13181, I1 => n38483, S => n26876, Z => 
                           n26251);
   U29187 : XOR2_X1 port map( A1 => n26404, A2 => n19890, Z => n26260);
   U29188 : NOR2_X1 port map( A1 => n948, A2 => n26269, ZN => n26268);
   U29189 : XOR2_X1 port map( A1 => n36958, A2 => n29657, Z => n26277);
   U29190 : INV_X1 port map( I => n26379, ZN => n26280);
   U29191 : XOR2_X1 port map( A1 => n334, A2 => n26476, Z => n26282);
   U29192 : XOR2_X1 port map( A1 => n12839, A2 => n19770, Z => n26281);
   U29194 : XOR2_X1 port map( A1 => n2150, A2 => n19839, Z => n26289);
   U29195 : NAND2_X1 port map( A1 => n13392, A2 => n26764, ZN => n26299);
   U29196 : XOR2_X1 port map( A1 => n12649, A2 => n29394, Z => n26292);
   U29197 : XOR2_X1 port map( A1 => n26293, A2 => n26292, Z => n26294);
   U29200 : XOR2_X1 port map( A1 => n26386, A2 => n26465, Z => n26297);
   U29201 : XOR2_X1 port map( A1 => n26591, A2 => n19527, Z => n26301);
   U29205 : XOR2_X1 port map( A1 => n26510, A2 => n19950, Z => n26310);
   U29206 : XOR2_X1 port map( A1 => n26311, A2 => n26310, Z => n26312);
   U29208 : NAND2_X1 port map( A1 => n36424, A2 => n14377, ZN => n26316);
   U29210 : XOR2_X1 port map( A1 => n9989, A2 => n26504, Z => n26317);
   U29211 : XOR2_X1 port map( A1 => n26438, A2 => n26584, Z => n26574);
   U29212 : XOR2_X1 port map( A1 => n26319, A2 => n29295, Z => n26320);
   U29213 : XOR2_X1 port map( A1 => n26320, A2 => n26574, Z => n26321);
   U29215 : NAND2_X1 port map( A1 => n26331, A2 => n7460, ZN => n26327);
   U29216 : NAND4_X1 port map( A1 => n19574, A2 => n19775, A3 => n26327, A4 => 
                           n26326, ZN => n26333);
   U29217 : NAND3_X1 port map( A1 => n26331, A2 => n26330, A3 => n7460, ZN => 
                           n26332);
   U29218 : XOR2_X1 port map( A1 => n26441, A2 => n9085, Z => n26336);
   U29221 : XOR2_X1 port map( A1 => n29554, A2 => n1010, Z => n26343);
   U29222 : XOR2_X1 port map( A1 => n30090, A2 => n34148, Z => n26350);
   U29224 : NAND2_X1 port map( A1 => n1091, A2 => n26804, ZN => n26355);
   U29225 : XOR2_X1 port map( A1 => n26359, A2 => n29879, Z => n26360);
   U29229 : XOR2_X1 port map( A1 => n26456, A2 => n26404, Z => n26371);
   U29231 : XOR2_X1 port map( A1 => n26380, A2 => n26518, Z => n26383);
   U29232 : XOR2_X1 port map( A1 => n26381, A2 => n26542, Z => n26382);
   U29233 : XOR2_X1 port map( A1 => n26383, A2 => n26382, Z => n26384);
   U29234 : INV_X1 port map( I => n26389, ZN => n26390);
   U29235 : XOR2_X1 port map( A1 => n26391, A2 => n35702, Z => n26392);
   U29236 : XOR2_X1 port map( A1 => n26404, A2 => n19936, Z => n26405);
   U29238 : XOR2_X1 port map( A1 => n26456, A2 => n26407, Z => n26409);
   U29243 : NAND2_X1 port map( A1 => n26424, A2 => n19762, ZN => n26426);
   U29249 : XOR2_X1 port map( A1 => n35251, A2 => n26460, Z => n26461);
   U29250 : XOR2_X1 port map( A1 => n1238, A2 => n29538, Z => n26464);
   U29252 : XOR2_X1 port map( A1 => n34469, A2 => n19804, Z => n26473);
   U29253 : XOR2_X1 port map( A1 => n19450, A2 => n19622, Z => n26493);
   U29254 : XOR2_X1 port map( A1 => n35251, A2 => n19801, Z => n26496);
   U29256 : NAND2_X1 port map( A1 => n26936, A2 => n26937, ZN => n26515);
   U29257 : XOR2_X1 port map( A1 => n11105, A2 => n19774, Z => n26536);
   U29258 : XOR2_X1 port map( A1 => n39793, A2 => n26542, Z => n26544);
   U29260 : XOR2_X1 port map( A1 => n32464, A2 => n19732, Z => n26562);
   U29261 : INV_X1 port map( I => n26560, ZN => n26561);
   U29267 : XOR2_X1 port map( A1 => n26599, A2 => n19908, Z => n26600);
   U29268 : INV_X1 port map( I => n26989, ZN => n26607);
   U29270 : NAND2_X1 port map( A1 => n26692, A2 => n26879, ZN => n26610);
   U29274 : NOR2_X1 port map( A1 => n20223, A2 => n26780, ZN => n26621);
   U29280 : INV_X1 port map( I => n26929, ZN => n26636);
   U29288 : OAI21_X1 port map( A1 => n35197, A2 => n19442, B => n14488, ZN => 
                           n26675);
   U29289 : MUX2_X1 port map( I0 => n20021, I1 => n26675, S => n26674, Z => 
                           n26678);
   U29299 : NOR2_X1 port map( A1 => n33858, A2 => n26961, ZN => n26721);
   U29301 : NOR2_X1 port map( A1 => n26948, A2 => n39595, ZN => n26730);
   U29302 : NOR3_X1 port map( A1 => n26951, A2 => n26731, A3 => n26730, ZN => 
                           n26732);
   U29304 : NAND3_X1 port map( A1 => n17047, A2 => n26740, A3 => n1235, ZN => 
                           n26741);
   U29308 : OAI21_X1 port map( A1 => n12755, A2 => n19179, B => n26760, ZN => 
                           n26762);
   U29310 : NOR2_X1 port map( A1 => n26934, A2 => n17993, ZN => n26776);
   U29313 : NAND2_X1 port map( A1 => n866, A2 => n17712, ZN => n26783);
   U29314 : NAND2_X1 port map( A1 => n39564, A2 => n9147, ZN => n26793);
   U29318 : NAND2_X1 port map( A1 => n39823, A2 => n20321, ZN => n26842);
   U29320 : OAI21_X1 port map( A1 => n26849, A2 => n26945, B => n26848, ZN => 
                           n26850);
   U29321 : MUX2_X1 port map( I0 => n26851, I1 => n26850, S => n20660, Z => 
                           n26853);
   U29325 : NAND2_X1 port map( A1 => n30429, A2 => n27138, ZN => n26887);
   U29326 : NOR2_X1 port map( A1 => n26923, A2 => n26922, ZN => n26897);
   U29327 : XOR2_X1 port map( A1 => n19612, A2 => n29474, Z => n26916);
   U29330 : AOI21_X1 port map( A1 => n859, A2 => n26936, B => n26935, ZN => 
                           n26939);
   U29331 : NAND2_X1 port map( A1 => n36477, A2 => n26937, ZN => n26938);
   U29334 : INV_X1 port map( I => n26955, ZN => n26956);
   U29335 : NAND2_X1 port map( A1 => n26957, A2 => n8103, ZN => n26958);
   U29336 : NAND3_X1 port map( A1 => n27508, A2 => n31287, A3 => n19529, ZN => 
                           n26965);
   U29338 : NAND2_X1 port map( A1 => n26981, A2 => n26980, ZN => n26985);
   U29340 : NAND2_X1 port map( A1 => n26992, A2 => n13111, ZN => n26993);
   U29341 : NAND2_X1 port map( A1 => n27108, A2 => n18246, ZN => n26998);
   U29346 : NOR2_X1 port map( A1 => n27044, A2 => n27043, ZN => n27048);
   U29347 : INV_X1 port map( I => n27045, ZN => n27047);
   U29349 : NOR2_X1 port map( A1 => n27059, A2 => n38571, ZN => n27060);
   U29351 : XOR2_X1 port map( A1 => n38937, A2 => n16613, Z => n27080);
   U29354 : XOR2_X1 port map( A1 => n27362, A2 => n27087, Z => n27088);
   U29355 : XOR2_X1 port map( A1 => n27089, A2 => n27088, Z => n27481);
   U29357 : NAND2_X1 port map( A1 => n27092, A2 => n15276, ZN => n27094);
   U29358 : NAND3_X1 port map( A1 => n20092, A2 => n13992, A3 => n27098, ZN => 
                           n27099);
   U29362 : NAND3_X1 port map( A1 => n32697, A2 => n19334, A3 => n18717, ZN => 
                           n27106);
   U29363 : NAND3_X1 port map( A1 => n27180, A2 => n1085, A3 => n1478, ZN => 
                           n27109);
   U29364 : NAND2_X1 port map( A1 => n27430, A2 => n30986, ZN => n27121);
   U29366 : INV_X1 port map( I => n27124, ZN => n27127);
   U29367 : INV_X1 port map( I => n27125, ZN => n27126);
   U29368 : INV_X1 port map( I => n27139, ZN => n27143);
   U29369 : INV_X1 port map( I => n27140, ZN => n27142);
   U29370 : NAND4_X1 port map( A1 => n27144, A2 => n27143, A3 => n27142, A4 => 
                           n9593, ZN => n27145);
   U29374 : NAND2_X1 port map( A1 => n27175, A2 => n33369, ZN => n27176);
   U29380 : NAND3_X1 port map( A1 => n27391, A2 => n35895, A3 => n13699, ZN => 
                           n27203);
   U29383 : OAI21_X1 port map( A1 => n37, A2 => n38579, B => n1448, ZN => 
                           n27215);
   U29385 : AOI21_X1 port map( A1 => n28495, A2 => n1427, B => n7454, ZN => 
                           n27458);
   U29387 : INV_X1 port map( I => n27224, ZN => n27225);
   U29388 : XOR2_X1 port map( A1 => n27592, A2 => n19883, Z => n27229);
   U29394 : XOR2_X1 port map( A1 => n37812, A2 => n30065, Z => n27302);
   U29395 : NAND3_X1 port map( A1 => n14614, A2 => n4434, A3 => n27409, ZN => 
                           n27316);
   U29398 : INV_X1 port map( I => n27334, ZN => n27335);
   U29401 : NAND2_X1 port map( A1 => n19455, A2 => n38571, ZN => n27353);
   U29403 : NAND2_X1 port map( A1 => n33050, A2 => n35228, ZN => n27369);
   U29407 : NAND2_X1 port map( A1 => n27384, A2 => n33336, ZN => n27386);
   U29408 : NOR2_X1 port map( A1 => n27417, A2 => n27416, ZN => n27419);
   U29413 : NAND2_X1 port map( A1 => n4847, A2 => n27449, ZN => n27451);
   U29414 : NAND3_X1 port map( A1 => n27452, A2 => n2923, A3 => n27451, ZN => 
                           n27453);
   U29415 : XOR2_X1 port map( A1 => n13289, A2 => n27849, Z => n27461);
   U29416 : XOR2_X1 port map( A1 => n27594, A2 => n27766, Z => n27463);
   U29417 : XOR2_X1 port map( A1 => n27540, A2 => n29970, Z => n27467);
   U29418 : XNOR2_X1 port map( A1 => n27663, A2 => n29711, ZN => n27471);
   U29420 : XOR2_X1 port map( A1 => n29319, A2 => n27815, Z => n27479);
   U29421 : NAND2_X1 port map( A1 => n28124, A2 => n14404, ZN => n27482);
   U29422 : MUX2_X1 port map( I0 => n27486, I1 => n27485, S => n33335, Z => 
                           n27489);
   U29423 : INV_X1 port map( I => n27487, ZN => n27488);
   U29424 : XOR2_X1 port map( A1 => n4934, A2 => n29879, Z => n27491);
   U29425 : INV_X1 port map( I => Key(184), ZN => n29017);
   U29428 : XOR2_X1 port map( A1 => n38205, A2 => n27525, Z => n27514);
   U29429 : INV_X1 port map( I => n27592, ZN => n27517);
   U29430 : XOR2_X1 port map( A1 => n19612, A2 => n27517, Z => n27518);
   U29431 : XOR2_X1 port map( A1 => n27661, A2 => n29978, Z => n27521);
   U29432 : XOR2_X1 port map( A1 => n7549, A2 => n29432, Z => n27522);
   U29433 : XOR2_X1 port map( A1 => n38228, A2 => n29689, Z => n27529);
   U29435 : XOR2_X1 port map( A1 => n4934, A2 => n19929, Z => n27533);
   U29436 : XOR2_X1 port map( A1 => n27738, A2 => n19804, Z => n27536);
   U29438 : XOR2_X1 port map( A1 => n27661, A2 => n29371, Z => n27548);
   U29440 : XOR2_X1 port map( A1 => n16320, A2 => n4934, Z => n27551);
   U29441 : NAND2_X1 port map( A1 => n27553, A2 => n38860, ZN => n27572);
   U29442 : XOR2_X1 port map( A1 => n27786, A2 => n19721, Z => n27568);
   U29443 : XOR2_X1 port map( A1 => n37499, A2 => n19735, Z => n27577);
   U29444 : XOR2_X1 port map( A1 => n27735, A2 => n19498, Z => n27578);
   U29446 : NOR2_X1 port map( A1 => n27589, A2 => n27588, ZN => n27590);
   U29448 : XOR2_X1 port map( A1 => n29223, A2 => n27758, Z => n27600);
   U29449 : XOR2_X1 port map( A1 => n27601, A2 => n27600, Z => n27602);
   U29450 : XOR2_X1 port map( A1 => n27603, A2 => n27602, Z => n27604);
   U29451 : XOR2_X1 port map( A1 => n27609, A2 => n27608, Z => n27614);
   U29452 : XOR2_X1 port map( A1 => n34829, A2 => n29801, Z => n27611);
   U29453 : XOR2_X1 port map( A1 => n27612, A2 => n27611, Z => n27613);
   U29456 : XOR2_X1 port map( A1 => n35177, A2 => n30248, Z => n27627);
   U29457 : XOR2_X1 port map( A1 => n27633, A2 => n27828, Z => n27634);
   U29458 : XOR2_X1 port map( A1 => n17418, A2 => n27637, Z => n27639);
   U29459 : XOR2_X1 port map( A1 => n19355, A2 => n19613, Z => n27638);
   U29460 : XOR2_X1 port map( A1 => n27640, A2 => n29141, Z => n27641);
   U29461 : INV_X1 port map( I => n28074, ZN => n27652);
   U29462 : XOR2_X1 port map( A1 => n900, A2 => n27823, Z => n27649);
   U29463 : XOR2_X1 port map( A1 => n4934, A2 => n19738, Z => n27651);
   U29464 : XOR2_X1 port map( A1 => n19913, A2 => n27724, Z => n27658);
   U29466 : XOR2_X1 port map( A1 => n27679, A2 => n19612, Z => n27681);
   U29471 : XOR2_X1 port map( A1 => n27703, A2 => n31602, Z => n27704);
   U29472 : XOR2_X1 port map( A1 => n27754, A2 => n27705, Z => n27706);
   U29473 : XOR2_X1 port map( A1 => n27848, A2 => n19937, Z => n27720);
   U29474 : XOR2_X1 port map( A1 => n38207, A2 => n27739, Z => n27740);
   U29475 : INV_X1 port map( I => n27870, ZN => n27741);
   U29478 : XOR2_X1 port map( A1 => n27761, A2 => n29399, Z => n27762);
   U29479 : XOR2_X1 port map( A1 => n27860, A2 => n29363, Z => n27764);
   U29480 : XOR2_X1 port map( A1 => n27765, A2 => n27764, Z => n27771);
   U29481 : XOR2_X1 port map( A1 => n27767, A2 => n27766, Z => n27768);
   U29482 : XOR2_X1 port map( A1 => n27769, A2 => n27768, Z => n27770);
   U29484 : XOR2_X1 port map( A1 => n27786, A2 => n27787, Z => n27789);
   U29485 : XOR2_X1 port map( A1 => n27796, A2 => n19648, Z => n27797);
   U29486 : XOR2_X1 port map( A1 => n35190, A2 => n30068, Z => n27803);
   U29487 : XOR2_X1 port map( A1 => n31585, A2 => n29282, Z => n27812);
   U29489 : MUX2_X1 port map( I0 => n3989, I1 => n28255, S => n19601, Z => 
                           n27822);
   U29490 : XOR2_X1 port map( A1 => n37338, A2 => n27834, Z => n27836);
   U29491 : XOR2_X1 port map( A1 => n4934, A2 => n19833, Z => n27839);
   U29495 : NOR2_X1 port map( A1 => n28727, A2 => n38230, ZN => n27879);
   U29496 : XOR2_X1 port map( A1 => n28874, A2 => n19902, Z => n27880);
   U29499 : NAND3_X1 port map( A1 => n28103, A2 => n17314, A3 => n32352, ZN => 
                           n27889);
   U29500 : NAND2_X2 port map( A1 => n27890, A2 => n27889, ZN => n28696);
   U29501 : INV_X1 port map( I => n28066, ZN => n27892);
   U29505 : NAND3_X1 port map( A1 => n28224, A2 => n39112, A3 => n28229, ZN => 
                           n27913);
   U29507 : NOR2_X1 port map( A1 => n28715, A2 => n31015, ZN => n27927);
   U29509 : NOR2_X1 port map( A1 => n33460, A2 => n31015, ZN => n27926);
   U29511 : XOR2_X1 port map( A1 => n36913, A2 => n28827, Z => n27943);
   U29514 : XOR2_X1 port map( A1 => n19774, A2 => n29833, Z => n27942);
   U29522 : NAND2_X1 port map( A1 => n28256, A2 => n28260, ZN => n27982);
   U29523 : NAND2_X1 port map( A1 => n1420, A2 => n13379, ZN => n27984);
   U29524 : NAND3_X1 port map( A1 => n38365, A2 => n11375, A3 => n879, ZN => 
                           n27983);
   U29525 : NAND2_X1 port map( A1 => n8522, A2 => n5266, ZN => n27986);
   U29527 : NAND3_X1 port map( A1 => n28238, A2 => n28103, A3 => n1453, ZN => 
                           n27992);
   U29530 : NAND2_X1 port map( A1 => n32783, A2 => n1450, ZN => n28007);
   U29531 : NAND2_X1 port map( A1 => n34120, A2 => n13714, ZN => n28006);
   U29532 : NAND2_X1 port map( A1 => n28008, A2 => n1447, ZN => n28009);
   U29533 : NAND2_X1 port map( A1 => n28011, A2 => n28012, ZN => n28014);
   U29537 : NAND2_X1 port map( A1 => n20739, A2 => n4803, ZN => n28021);
   U29538 : NAND2_X1 port map( A1 => n28025, A2 => n28024, ZN => n28026);
   U29539 : NAND2_X1 port map( A1 => n28027, A2 => n28026, ZN => n28030);
   U29540 : OAI21_X1 port map( A1 => n28035, A2 => n28034, B => n36979, ZN => 
                           n28039);
   U29545 : NAND2_X1 port map( A1 => n19280, A2 => n1205, ZN => n28057);
   U29546 : NOR3_X1 port map( A1 => n1072, A2 => n34008, A3 => n28054, ZN => 
                           n28056);
   U29548 : NAND2_X1 port map( A1 => n28064, A2 => n28155, ZN => n28065);
   U29555 : XOR2_X1 port map( A1 => n29689, A2 => n28982, Z => n28100);
   U29556 : NAND2_X1 port map( A1 => n7325, A2 => n984, ZN => n28107);
   U29558 : NAND3_X1 port map( A1 => n19946, A2 => n28133, A3 => n28131, ZN => 
                           n28134);
   U29564 : MUX2_X1 port map( I0 => n28228, I1 => n28229, S => n28224, Z => 
                           n28226);
   U29568 : NAND2_X1 port map( A1 => n28257, A2 => n28256, ZN => n28259);
   U29570 : NAND2_X1 port map( A1 => n37329, A2 => n28157, ZN => n28270);
   U29573 : NAND2_X1 port map( A1 => n28307, A2 => n9599, ZN => n28308);
   U29574 : AOI21_X1 port map( A1 => n28632, A2 => n14209, B => n28635, ZN => 
                           n28317);
   U29575 : INV_X1 port map( I => n28634, ZN => n28316);
   U29576 : INV_X1 port map( I => n28633, ZN => n28315);
   U29577 : XOR2_X1 port map( A1 => n28319, A2 => n28318, Z => n28320);
   U29578 : NAND4_X1 port map( A1 => n28326, A2 => n19038, A3 => n28325, A4 => 
                           n30389, ZN => n28328);
   U29579 : XOR2_X1 port map( A1 => n4816, A2 => n19879, Z => n28332);
   U29581 : NAND2_X1 port map( A1 => n11413, A2 => n1433, ZN => n28337);
   U29583 : NAND2_X1 port map( A1 => n28350, A2 => n28349, ZN => n28354);
   U29586 : NAND2_X1 port map( A1 => n28509, A2 => n33460, ZN => n28364);
   U29595 : XOR2_X1 port map( A1 => n29221, A2 => n19035, Z => n28411);
   U29596 : XOR2_X1 port map( A1 => n29001, A2 => n28411, Z => n28412);
   U29598 : INV_X1 port map( I => n28418, ZN => n28421);
   U29599 : NAND3_X1 port map( A1 => n28421, A2 => n28420, A3 => n28419, ZN => 
                           n28424);
   U29600 : NAND2_X1 port map( A1 => n28422, A2 => n35694, ZN => n28423);
   U29601 : NOR3_X1 port map( A1 => n18871, A2 => n31045, A3 => n1429, ZN => 
                           n28426);
   U29602 : MUX2_X1 port map( I0 => n18875, I1 => n28437, S => n28554, Z => 
                           n28429);
   U29608 : NAND2_X1 port map( A1 => n17735, A2 => n32002, ZN => n28475);
   U29610 : MUX2_X1 port map( I0 => n28486, I1 => n28485, S => n28484, Z => 
                           n28487);
   U29611 : NAND2_X1 port map( A1 => n28487, A2 => n19893, ZN => n28488);
   U29618 : NAND2_X1 port map( A1 => n28745, A2 => n34244, ZN => n28524);
   U29620 : AOI21_X1 port map( A1 => n28530, A2 => n12527, B => n39435, ZN => 
                           n28531);
   U29622 : XOR2_X1 port map( A1 => n7288, A2 => n29832, Z => n28534);
   U29623 : XOR2_X1 port map( A1 => n29076, A2 => n28534, Z => n28542);
   U29624 : XOR2_X1 port map( A1 => n29247, A2 => n19860, Z => n28541);
   U29626 : XOR2_X1 port map( A1 => n28783, A2 => n10794, Z => n28540);
   U29627 : XOR2_X1 port map( A1 => n28791, A2 => n19770, Z => n28549);
   U29631 : NAND2_X1 port map( A1 => n1404, A2 => n29486, ZN => n28583);
   U29632 : AOI21_X1 port map( A1 => n29596, A2 => n33482, B => n28583, ZN => 
                           n28584);
   U29634 : NAND3_X1 port map( A1 => n9599, A2 => n35199, A3 => n35888, ZN => 
                           n28592);
   U29637 : XOR2_X1 port map( A1 => n28891, A2 => n28783, Z => n28630);
   U29646 : XOR2_X1 port map( A1 => n29303, A2 => n29145, Z => n28763);
   U29647 : XOR2_X1 port map( A1 => n29058, A2 => n19894, Z => n28762);
   U29649 : XOR2_X1 port map( A1 => n38189, A2 => n29647, Z => n28775);
   U29650 : INV_X1 port map( I => n19592, ZN => n28776);
   U29651 : XOR2_X1 port map( A1 => n18242, A2 => n29122, Z => n28779);
   U29652 : XOR2_X1 port map( A1 => n29121, A2 => n19936, Z => n28778);
   U29653 : XOR2_X1 port map( A1 => n28779, A2 => n28778, Z => n28782);
   U29654 : XOR2_X1 port map( A1 => n28991, A2 => n5130, Z => n28786);
   U29655 : XOR2_X1 port map( A1 => n28786, A2 => n28785, Z => n28787);
   U29656 : XOR2_X1 port map( A1 => n28842, A2 => n28794, Z => n28795);
   U29657 : NAND3_X1 port map( A1 => n28798, A2 => n28799, A3 => n15273, ZN => 
                           n28797);
   U29658 : OAI21_X1 port map( A1 => n28800, A2 => n28798, B => n28797, ZN => 
                           n28802);
   U29659 : NOR2_X1 port map( A1 => n28802, A2 => n28801, ZN => n28803);
   U29660 : XOR2_X1 port map( A1 => n28990, A2 => n28803, Z => n28804);
   U29661 : XOR2_X1 port map( A1 => n296, A2 => n30114, Z => n28806);
   U29662 : AOI21_X1 port map( A1 => n28808, A2 => n33577, B => n976, ZN => 
                           n28811);
   U29663 : XOR2_X1 port map( A1 => n28813, A2 => n30888, Z => n28814);
   U29664 : XOR2_X1 port map( A1 => n29824, A2 => n19760, Z => n28815);
   U29666 : XOR2_X1 port map( A1 => n28865, A2 => n27465, Z => n28820);
   U29668 : NAND2_X1 port map( A1 => n30161, A2 => n29185, ZN => n28825);
   U29669 : XOR2_X1 port map( A1 => n36913, A2 => n5130, Z => n28828);
   U29670 : XOR2_X1 port map( A1 => n29142, A2 => n29718, Z => n28844);
   U29673 : XOR2_X1 port map( A1 => n29837, A2 => n19780, Z => n28849);
   U29674 : XOR2_X1 port map( A1 => n28851, A2 => n28852, Z => n29099);
   U29675 : XOR2_X1 port map( A1 => n28855, A2 => n28854, Z => n28859);
   U29676 : XOR2_X1 port map( A1 => n29030, A2 => n28857, Z => n28858);
   U29677 : NAND3_X1 port map( A1 => n28962, A2 => n28862, A3 => n1178, ZN => 
                           n28863);
   U29678 : XOR2_X1 port map( A1 => n29063, A2 => n28865, Z => n28866);
   U29683 : INV_X1 port map( I => n28883, ZN => n29592);
   U29684 : INV_X1 port map( I => n29483, ZN => n29645);
   U29685 : NOR2_X1 port map( A1 => n29642, A2 => n29643, ZN => n29578);
   U29688 : XOR2_X1 port map( A1 => n19952, A2 => n28891, Z => n28892);
   U29689 : XOR2_X1 port map( A1 => n28893, A2 => n28892, Z => n28894);
   U29690 : XOR2_X1 port map( A1 => n39220, A2 => n19933, Z => n28898);
   U29693 : NAND2_X1 port map( A1 => n28901, A2 => n28900, ZN => n28903);
   U29694 : NAND2_X1 port map( A1 => n29548, A2 => n35176, ZN => n29556);
   U29695 : NAND2_X1 port map( A1 => n28904, A2 => n29556, ZN => n28905);
   U29696 : XOR2_X1 port map( A1 => n29058, A2 => n19732, Z => n28912);
   U29697 : XOR2_X1 port map( A1 => n34848, A2 => n31127, Z => n28915);
   U29698 : XOR2_X1 port map( A1 => n28916, A2 => n28915, Z => n28919);
   U29699 : XOR2_X1 port map( A1 => n16336, A2 => n28917, Z => n28918);
   U29700 : XOR2_X1 port map( A1 => n31396, A2 => n9930, Z => n28930);
   U29702 : XOR2_X1 port map( A1 => n29306, A2 => n35140, Z => n28935);
   U29704 : XOR2_X1 port map( A1 => n32022, A2 => n19943, Z => n28944);
   U29707 : XOR2_X1 port map( A1 => n29115, A2 => n29146, Z => n28951);
   U29711 : AND2_X1 port map( A1 => n28963, A2 => n28962, Z => n28964);
   U29712 : XOR2_X1 port map( A1 => n29023, A2 => n29123, Z => n28976);
   U29715 : OAI21_X1 port map( A1 => n9649, A2 => n29863, B => n19878, ZN => 
                           n28980);
   U29718 : XOR2_X1 port map( A1 => n9106, A2 => n10794, Z => n28993);
   U29719 : XOR2_X1 port map( A1 => n28991, A2 => n16320, Z => n28992);
   U29720 : XOR2_X1 port map( A1 => n28993, A2 => n28992, Z => n28994);
   U29721 : NAND2_X1 port map( A1 => n29940, A2 => n34179, ZN => n28996);
   U29722 : XOR2_X1 port map( A1 => n28997, A2 => n37112, Z => n28998);
   U29726 : NAND2_X1 port map( A1 => n30134, A2 => n37117, ZN => n29014);
   U29727 : NAND2_X1 port map( A1 => n29014, A2 => n30136, ZN => n29016);
   U29728 : XOR2_X1 port map( A1 => n29019, A2 => n31249, Z => Ciphertext(61));
   U29729 : XOR2_X1 port map( A1 => n29837, A2 => n29034, Z => n29035);
   U29730 : XOR2_X1 port map( A1 => n29824, A2 => n29320, Z => n29046);
   U29731 : XOR2_X1 port map( A1 => n29801, A2 => n6661, Z => n29055);
   U29732 : XOR2_X1 port map( A1 => n19513, A2 => n29063, Z => n29064);
   U29734 : XOR2_X1 port map( A1 => n17039, A2 => n29805, Z => n29075);
   U29735 : XOR2_X1 port map( A1 => n29076, A2 => n29075, Z => n29077);
   U29736 : XOR2_X1 port map( A1 => n29970, A2 => n29082, Z => n29083);
   U29738 : XOR2_X1 port map( A1 => n29088, A2 => n30253, Z => n29089);
   U29739 : XOR2_X1 port map( A1 => n29090, A2 => n29089, Z => n29091);
   U29740 : XOR2_X1 port map( A1 => n19622, A2 => n29096, Z => n29097);
   U29743 : XOR2_X1 port map( A1 => n19937, A2 => n16357, Z => n29107);
   U29744 : XOR2_X1 port map( A1 => n15581, A2 => n29109, Z => n29110);
   U29746 : XOR2_X1 port map( A1 => n29133, A2 => n29132, Z => n29134);
   U29747 : XOR2_X1 port map( A1 => n31522, A2 => n18242, Z => n29156);
   U29748 : XOR2_X1 port map( A1 => n29155, A2 => n29156, Z => n29157);
   U29751 : NOR2_X1 port map( A1 => n30093, A2 => n35175, ZN => n29176);
   U29756 : NAND2_X1 port map( A1 => n29843, A2 => n773, ZN => n29190);
   U29757 : MUX2_X1 port map( I0 => n29190, I1 => n29871, S => n29869, Z => 
                           n29193);
   U29758 : NAND2_X1 port map( A1 => n29692, A2 => n28, ZN => n29191);
   U29759 : NAND3_X1 port map( A1 => n29871, A2 => n37936, A3 => n29191, ZN => 
                           n29192);
   U29762 : NOR2_X1 port map( A1 => n29241, A2 => n29346, ZN => n29212);
   U29764 : INV_X1 port map( I => n30238, ZN => n29214);
   U29766 : XOR2_X1 port map( A1 => n29217, A2 => n30803, Z => Ciphertext(8));
   U29768 : NOR2_X1 port map( A1 => n29231, A2 => n29236, ZN => n29232);
   U29770 : XOR2_X1 port map( A1 => n1410, A2 => n29357, Z => n29244);
   U29773 : XOR2_X1 port map( A1 => n38221, A2 => n29290, Z => n29293);
   U29774 : XOR2_X1 port map( A1 => n29829, A2 => n1697, Z => n29291);
   U29776 : NOR2_X1 port map( A1 => n771, A2 => n37100, ZN => n29314);
   U29777 : NOR3_X1 port map( A1 => n14400, A2 => n29446, A3 => n29445, ZN => 
                           n29313);
   U29780 : XOR2_X1 port map( A1 => n29338, A2 => n1718, Z => n29323);
   U29781 : NAND3_X1 port map( A1 => n29323, A2 => n29335, A3 => n1391, ZN => 
                           n29332);
   U29782 : NAND3_X1 port map( A1 => n29324, A2 => n29338, A3 => n32790, ZN => 
                           n29331);
   U29783 : XOR2_X1 port map( A1 => n29325, A2 => n29339, Z => n29326);
   U29784 : NAND3_X1 port map( A1 => n29326, A2 => n20481, A3 => n38156, ZN => 
                           n29330);
   U29785 : XOR2_X1 port map( A1 => n16889, A2 => n1718, Z => n29327);
   U29786 : NAND2_X1 port map( A1 => n29328, A2 => n29327, ZN => n29329);
   U29787 : NAND4_X1 port map( A1 => n29332, A2 => n29331, A3 => n29330, A4 => 
                           n29329, ZN => Ciphertext(26));
   U29788 : INV_X1 port map( I => Key(81), ZN => n29337);
   U29790 : NAND2_X1 port map( A1 => n29361, A2 => n31307, ZN => n29356);
   U29793 : NOR2_X1 port map( A1 => n29373, A2 => n37096, ZN => n29359);
   U29794 : INV_X1 port map( I => n19933, ZN => n29360);
   U29798 : NAND3_X1 port map( A1 => n29410, A2 => n29413, A3 => n9790, ZN => 
                           n29393);
   U29803 : NAND3_X1 port map( A1 => n29390, A2 => n29413, A3 => n17849, ZN => 
                           n29391);
   U29805 : NAND2_X1 port map( A1 => n29413, A2 => n29409, ZN => n29396);
   U29807 : INV_X1 port map( I => n17849, ZN => n29407);
   U29808 : INV_X1 port map( I => n29413, ZN => n29408);
   U29809 : AOI21_X1 port map( A1 => n35272, A2 => n17849, B => n29412, ZN => 
                           n29415);
   U29810 : XOR2_X1 port map( A1 => n29417, A2 => n19732, Z => Ciphertext(41));
   U29812 : OAI21_X1 port map( A1 => n1392, A2 => n29438, B => n29434, ZN => 
                           n29431);
   U29813 : NOR3_X1 port map( A1 => n771, A2 => n14400, A3 => n29446, ZN => 
                           n29447);
   U29814 : INV_X1 port map( I => n29461, ZN => n29469);
   U29815 : XOR2_X1 port map( A1 => n29467, A2 => n19839, Z => Ciphertext(50));
   U29817 : OAI21_X1 port map( A1 => n9636, A2 => n39178, B => n29490, ZN => 
                           n29505);
   U29818 : NAND2_X1 port map( A1 => n29527, A2 => n33427, ZN => n29504);
   U29821 : XOR2_X1 port map( A1 => n29510, A2 => n29509, Z => Ciphertext(55));
   U29822 : MUX2_X1 port map( I0 => n19362, I1 => n35180, S => n18384, Z => 
                           n29513);
   U29824 : AOI21_X1 port map( A1 => n29513, A2 => n29517, B => n29512, ZN => 
                           n29515);
   U29825 : XOR2_X1 port map( A1 => n29515, A2 => n29514, Z => Ciphertext(56));
   U29828 : NAND2_X1 port map( A1 => n29519, A2 => n32317, ZN => n29520);
   U29829 : XOR2_X1 port map( A1 => n29523, A2 => n29522, Z => Ciphertext(57));
   U29830 : OAI21_X1 port map( A1 => n33427, A2 => n35180, B => n29524, ZN => 
                           n29526);
   U29831 : XOR2_X1 port map( A1 => n29529, A2 => n29528, Z => Ciphertext(58));
   U29832 : AOI21_X1 port map( A1 => n39178, A2 => n29531, B => n19362, ZN => 
                           n29533);
   U29835 : XOR2_X1 port map( A1 => n29539, A2 => n1698, Z => Ciphertext(60));
   U29837 : MUX2_X1 port map( I0 => n29548, I1 => n35176, S => n29555, Z => 
                           n29549);
   U29838 : NAND2_X1 port map( A1 => n29556, A2 => n29555, ZN => n29557);
   U29840 : NOR2_X1 port map( A1 => n29565, A2 => n29570, ZN => n29569);
   U29841 : XOR2_X1 port map( A1 => n29573, A2 => n35140, Z => Ciphertext(70));
   U29842 : NOR2_X1 port map( A1 => n20979, A2 => n19147, ZN => n29580);
   U29843 : INV_X1 port map( I => n29578, ZN => n29579);
   U29848 : NOR2_X1 port map( A1 => n29597, A2 => n29596, ZN => n29599);
   U29850 : AOI21_X1 port map( A1 => n35405, A2 => n29618, B => n29616, ZN => 
                           n29605);
   U29853 : OAI21_X1 port map( A1 => n29616, A2 => n31540, B => n29617, ZN => 
                           n29607);
   U29854 : XOR2_X1 port map( A1 => n29610, A2 => n1733, Z => Ciphertext(74));
   U29855 : MUX2_X1 port map( I0 => n29616, I1 => n29617, S => n29619, Z => 
                           n29613);
   U29856 : XOR2_X1 port map( A1 => n29615, A2 => n29614, Z => Ciphertext(75));
   U29857 : NAND2_X1 port map( A1 => n31540, A2 => n29619, ZN => n29621);
   U29858 : NAND2_X1 port map( A1 => n29624, A2 => n29623, ZN => n29628);
   U29859 : INV_X1 port map( I => n29630, ZN => n29631);
   U29862 : NOR3_X1 port map( A1 => n481, A2 => n29776, A3 => n34914, ZN => 
                           n29640);
   U29867 : NAND2_X1 port map( A1 => n19297, A2 => n29641, ZN => n29652);
   U29868 : OAI21_X1 port map( A1 => n29662, A2 => n19297, B => n17382, ZN => 
                           n29663);
   U29873 : NAND2_X1 port map( A1 => n29712, A2 => n29708, ZN => n29710);
   U29875 : NAND3_X1 port map( A1 => n14337, A2 => n29720, A3 => n29721, ZN => 
                           n29715);
   U29877 : AOI21_X1 port map( A1 => n29726, A2 => n19348, B => n29725, ZN => 
                           n29727);
   U29878 : XOR2_X1 port map( A1 => n29727, A2 => n1369, Z => Ciphertext(96));
   U29880 : NOR2_X1 port map( A1 => n29729, A2 => n29752, ZN => n29731);
   U29881 : XOR2_X1 port map( A1 => n29731, A2 => n29730, Z => Ciphertext(97));
   U29883 : NOR3_X1 port map( A1 => n38143, A2 => n29732, A3 => n29754, ZN => 
                           n29733);
   U29893 : XOR2_X1 port map( A1 => n29759, A2 => n19583, Z => Ciphertext(101))
                           ;
   U29896 : AOI21_X1 port map( A1 => n1407, A2 => n29815, B => n29902, ZN => 
                           n29775);
   U29898 : NAND2_X1 port map( A1 => n29788, A2 => n19716, ZN => n29784);
   U29901 : NOR2_X1 port map( A1 => n29794, A2 => n29792, ZN => n29793);
   U29902 : NAND2_X1 port map( A1 => n29795, A2 => n29794, ZN => n29796);
   U29904 : NAND3_X1 port map( A1 => n29811, A2 => n6652, A3 => n39018, ZN => 
                           n29807);
   U29905 : XOR2_X1 port map( A1 => n29809, A2 => n29808, Z => Ciphertext(111))
                           ;
   U29906 : INV_X1 port map( I => n14403, ZN => n29900);
   U29907 : XOR2_X1 port map( A1 => n11923, A2 => n19885, Z => n29821);
   U29908 : INV_X1 port map( I => n19890, ZN => n29825);
   U29909 : XOR2_X1 port map( A1 => n39348, A2 => n29825, Z => n29827);
   U29910 : XOR2_X1 port map( A1 => n29828, A2 => n5130, Z => n29830);
   U29911 : INV_X1 port map( I => n11861, ZN => n29842);
   U29914 : NAND2_X1 port map( A1 => n29883, A2 => n38217, ZN => n29874);
   U29915 : INV_X1 port map( I => n29883, ZN => n29888);
   U29919 : NOR2_X1 port map( A1 => n30057, A2 => n16353, ZN => n29896);
   U29920 : NAND2_X1 port map( A1 => n1407, A2 => n29900, ZN => n29901);
   U29922 : NOR2_X1 port map( A1 => n29905, A2 => n29954, ZN => n29910);
   U29923 : OAI21_X1 port map( A1 => n29908, A2 => n19878, B => n29906, ZN => 
                           n29909);
   U29925 : AOI21_X1 port map( A1 => n29922, A2 => n1174, B => n29912, ZN => 
                           n29914);
   U29926 : XOR2_X1 port map( A1 => n29915, A2 => n16320, Z => Ciphertext(128))
                           ;
   U29928 : INV_X1 port map( I => n29927, ZN => n29928);
   U29929 : OAI21_X1 port map( A1 => n29929, A2 => n31570, B => n29928, ZN => 
                           n29933);
   U29930 : NAND2_X1 port map( A1 => n21285, A2 => n17240, ZN => n29947);
   U29931 : OAI21_X1 port map( A1 => n29960, A2 => n29955, B => n29954, ZN => 
                           n29959);
   U29932 : OAI21_X1 port map( A1 => n29957, A2 => n18104, B => n29956, ZN => 
                           n29958);
   U29933 : NAND2_X1 port map( A1 => n18104, A2 => n29960, ZN => n29961);
   U29934 : AOI21_X1 port map( A1 => n13705, A2 => n29977, B => n31512, ZN => 
                           n29962);
   U29936 : OAI21_X1 port map( A1 => n29982, A2 => n29973, B => n29966, ZN => 
                           n29967);
   U29937 : XOR2_X1 port map( A1 => n29967, A2 => n19897, Z => Ciphertext(133))
                           ;
   U29939 : NAND2_X1 port map( A1 => n9918, A2 => n19909, ZN => n29985);
   U29940 : NAND2_X1 port map( A1 => n29986, A2 => n29985, ZN => n29988);
   U29943 : NOR3_X1 port map( A1 => n15643, A2 => n30038, A3 => n30024, ZN => 
                           n30004);
   U29944 : NAND3_X1 port map( A1 => n8529, A2 => n32628, A3 => n36850, ZN => 
                           n30002);
   U29946 : XOR2_X1 port map( A1 => n30008, A2 => n30007, Z => Ciphertext(138))
                           ;
   U29947 : AOI21_X1 port map( A1 => n30037, A2 => n30024, B => n30011, ZN => 
                           n30012);
   U29949 : AOI21_X1 port map( A1 => n30025, A2 => n39407, B => n33311, ZN => 
                           n30021);
   U29950 : INV_X1 port map( I => n30017, ZN => n30019);
   U29951 : NOR2_X1 port map( A1 => n30033, A2 => n30022, ZN => n30018);
   U29952 : OAI21_X1 port map( A1 => n30019, A2 => n30018, B => n30037, ZN => 
                           n30020);
   U29953 : NAND2_X1 port map( A1 => n30021, A2 => n30020, ZN => n30030);
   U29954 : OAI21_X1 port map( A1 => n30035, A2 => n30033, B => n33311, ZN => 
                           n30023);
   U29955 : AOI21_X1 port map( A1 => n30025, A2 => n30024, B => n30023, ZN => 
                           n30028);
   U29956 : NAND2_X1 port map( A1 => n30026, A2 => n15643, ZN => n30027);
   U29957 : OAI21_X1 port map( A1 => n30035, A2 => n30034, B => n30033, ZN => 
                           n30036);
   U29959 : XOR2_X1 port map( A1 => n30040, A2 => n16332, Z => Ciphertext(143))
                           ;
   U29964 : XOR2_X1 port map( A1 => n30091, A2 => n30090, Z => Ciphertext(153))
                           ;
   U29967 : NOR2_X1 port map( A1 => n10118, A2 => n30117, ZN => n30102);
   U29968 : XOR2_X1 port map( A1 => n30105, A2 => n1163, Z => Ciphertext(157));
   U29969 : MUX2_X1 port map( I0 => n10118, I1 => n35187, S => n30117, Z => 
                           n30113);
   U29970 : NAND2_X1 port map( A1 => n30109, A2 => n35186, ZN => n30110);
   U29971 : XOR2_X1 port map( A1 => n30116, A2 => n30115, Z => Ciphertext(159))
                           ;
   U29974 : INV_X1 port map( I => n19721, ZN => n30130);
   U29976 : XOR2_X1 port map( A1 => n30140, A2 => n17463, Z => Ciphertext(170))
                           ;
   U29977 : NAND2_X1 port map( A1 => n34177, A2 => n30141, ZN => n30143);
   U29980 : NAND3_X1 port map( A1 => n30183, A2 => n16676, A3 => n17997, ZN => 
                           n30168);
   U29981 : INV_X1 port map( I => n30162, ZN => n30163);
   U29982 : NAND2_X1 port map( A1 => n30193, A2 => n35210, ZN => n30194);
   U29984 : NOR2_X1 port map( A1 => n31549, A2 => n30210, ZN => n30204);
   U29986 : OAI21_X1 port map( A1 => n30215, A2 => n30214, B => n30213, ZN => 
                           n30216);
   U29987 : NOR2_X1 port map( A1 => n1399, A2 => n30220, ZN => n30223);
   U29988 : NAND3_X1 port map( A1 => n10590, A2 => n17238, A3 => n29210, ZN => 
                           n30231);
   U29990 : MUX2_X1 port map( I0 => n30260, I1 => n30259, S => n30257, Z => 
                           n30255);
   U29991 : XOR2_X1 port map( A1 => n30256, A2 => n965, Z => Ciphertext(190));
   U29993 : OAI21_X1 port map( A1 => n30260, A2 => n30259, B => n30258, ZN => 
                           n30261);
   U6354 : OAI21_X2 port map( A1 => n1042, A2 => n1320, B => n5111, ZN => 
                           n23056);
   U1533 : INV_X2 port map( I => n7304, ZN => n21900);
   U8697 : AOI21_X2 port map( A1 => n9809, A2 => n19397, B => n21588, ZN => 
                           n18559);
   U10139 : AOI21_X2 port map( A1 => n37216, A2 => n20238, B => n1840, ZN => 
                           n1839);
   U357 : INV_X4 port map( I => n18689, ZN => n1206);
   U1348 : INV_X2 port map( I => n17169, ZN => n13995);
   U478 : INV_X2 port map( I => n7757, ZN => n27378);
   U6816 : NAND2_X2 port map( A1 => n25819, A2 => n32924, ZN => n12252);
   U1322 : INV_X4 port map( I => n19586, ZN => n1314);
   U10040 : OAI21_X2 port map( A1 => n8720, A2 => n23095, B => n39356, ZN => 
                           n8719);
   U1540 : INV_X4 port map( I => n3562, ZN => n21599);
   U5940 : INV_X2 port map( I => n728, ZN => n9161);
   U2360 : NAND2_X2 port map( A1 => n29426, A2 => n29454, ZN => n29453);
   U2417 : AOI21_X2 port map( A1 => n38580, A2 => n28744, B => n10081, ZN => 
                           n13671);
   U578 : INV_X2 port map( I => n17217, ZN => n18534);
   U219 : NAND2_X2 port map( A1 => n28010, A2 => n28009, ZN => n28569);
   U625 : INV_X2 port map( I => n26278, ZN => n26456);
   U481 : INV_X2 port map( I => n27267, ZN => n27266);
   U801 : OAI21_X2 port map( A1 => n25753, A2 => n579, B => n38300, ZN => n2316
                           );
   U6553 : INV_X2 port map( I => n8919, ZN => n29421);
   U6099 : INV_X2 port map( I => n12055, ZN => n8919);
   U22329 : AOI21_X2 port map( A1 => n20308, A2 => n12077, B => n10242, ZN => 
                           n20961);
   U6566 : INV_X2 port map( I => n30186, ZN => n30159);
   U5570 : INV_X2 port map( I => n29341, ZN => n1391);
   U1446 : NAND2_X2 port map( A1 => n15382, A2 => n15380, ZN => n22132);
   U6323 : INV_X2 port map( I => n10635, ZN => n1613);
   U1346 : INV_X2 port map( I => n13694, ZN => n23142);
   U753 : INV_X2 port map( I => n18987, ZN => n25770);
   U1454 : INV_X2 port map( I => n9970, ZN => n1151);
   U10923 : NAND2_X2 port map( A1 => n3965, A2 => n6435, ZN => n3964);
   U13851 : AOI21_X2 port map( A1 => n21694, A2 => n15910, B => n15812, ZN => 
                           n15811);
   U8778 : BUF_X2 port map( I => Key(30), Z => n29509);
   U1300 : AOI21_X2 port map( A1 => n1043, A2 => n19000, B => n14556, ZN => 
                           n23155);
   U50 : NAND2_X2 port map( A1 => n29272, A2 => n29273, ZN => n29277);
   U8104 : AOI22_X2 port map( A1 => n25427, A2 => n19296, B1 => n15180, B2 => 
                           n14515, ZN => n4595);
   U785 : NAND2_X2 port map( A1 => n17471, A2 => n4046, ZN => n26019);
   U586 : INV_X2 port map( I => n19225, ZN => n7752);
   U414 : NAND2_X2 port map( A1 => n21248, A2 => n31287, ZN => n27507);
   U1074 : NOR2_X2 port map( A1 => n24184, A2 => n24300, ZN => n13881);
   U6076 : NAND2_X2 port map( A1 => n33404, A2 => n18720, ZN => n16074);
   U1244 : INV_X2 port map( I => n4618, ZN => n23569);
   U897 : INV_X2 port map( I => n7967, ZN => n25116);
   U3017 : NAND2_X1 port map( A1 => n22829, A2 => n23042, ZN => n20911);
   U10480 : BUF_X2 port map( I => Key(9), Z => n19498);
   U1124 : INV_X2 port map( I => n14709, ZN => n24266);
   U18608 : INV_X4 port map( I => n20793, ZN => n29869);
   U5813 : NOR2_X2 port map( A1 => n3293, A2 => n21895, ZN => n13421);
   U7500 : AOI21_X2 port map( A1 => n9017, A2 => n34915, B => n33841, ZN => 
                           n9016);
   U13839 : NAND2_X2 port map( A1 => n14920, A2 => n14919, ZN => n21370);
   U25076 : NAND2_X2 port map( A1 => n7613, A2 => n133, ZN => n22187);
   U2474 : INV_X2 port map( I => n19844, ZN => n28311);
   U26764 : AOI22_X2 port map( A1 => n31359, A2 => n25468, B1 => n25609, B2 => 
                           n17332, ZN => n17331);
   U1402 : AOI21_X2 port map( A1 => n11277, A2 => n15229, B => n11276, ZN => 
                           n11275);
   U8055 : NAND2_X2 port map( A1 => n5098, A2 => n4516, ZN => n19241);
   U2487 : NOR2_X2 port map( A1 => n28772, A2 => n17771, ZN => n28293);
   U9923 : NAND2_X2 port map( A1 => n4207, A2 => n31931, ZN => n10709);
   U9639 : NAND2_X2 port map( A1 => n24770, A2 => n8173, ZN => n24772);
   U100 : INV_X2 port map( I => n37060, ZN => n6851);
   U7065 : AOI21_X2 port map( A1 => n20998, A2 => n10709, B => n23444, ZN => 
                           n9347);
   U2467 : NOR2_X2 port map( A1 => n11658, A2 => n30443, ZN => n13642);
   U8623 : INV_X2 port map( I => n22178, ZN => n1148);
   U10677 : INV_X1 port map( I => n29437, ZN => n1389);
   U6137 : INV_X2 port map( I => n16327, ZN => n28191);
   U1441 : INV_X2 port map( I => n22155, ZN => n15004);
   U163 : NOR2_X2 port map( A1 => n20737, A2 => n20736, ZN => n20735);
   U1093 : INV_X2 port map( I => n802, ZN => n24221);
   U1104 : INV_X4 port map( I => n17911, ZN => n1125);
   U8455 : NAND2_X2 port map( A1 => n14305, A2 => n19614, ZN => n8721);
   U11632 : NOR2_X2 port map( A1 => n27270, A2 => n33050, ZN => n16479);
   U15569 : AOI21_X2 port map( A1 => n13337, A2 => n3119, B => n13336, ZN => 
                           n13335);
   U5680 : INV_X2 port map( I => n833, ZN => n18734);
   U1442 : INV_X2 port map( I => n8493, ZN => n15493);
   U5518 : NAND2_X2 port map( A1 => n1300, A2 => n6218, ZN => n23553);
   U3123 : INV_X1 port map( I => n26876, ZN => n4218);
   U346 : INV_X2 port map( I => n27910, ZN => n15704);
   U9998 : INV_X2 port map( I => n22923, ZN => n15770);
   U7213 : INV_X2 port map( I => n9422, ZN => n18999);
   U7110 : INV_X2 port map( I => n23390, ZN => n1644);
   U13228 : AOI21_X2 port map( A1 => n37196, A2 => n23355, B => n32158, ZN => 
                           n19006);
   U821 : AOI21_X2 port map( A1 => n25472, A2 => n31359, B => n25409, ZN => 
                           n15404);
   U5938 : INV_X4 port map( I => n18164, ZN => n25359);
   U356 : INV_X2 port map( I => n5525, ZN => n28286);
   U8930 : AOI22_X2 port map( A1 => n17115, A2 => n3532, B1 => n1419, B2 => 
                           n28683, ZN => n18191);
   U6933 : NAND2_X2 port map( A1 => n19678, A2 => n25261, ZN => n15459);
   U14233 : AOI22_X2 port map( A1 => n4697, A2 => n9141, B1 => n1881, B2 => 
                           n33591, ZN => n4076);
   U1769 : NAND2_X1 port map( A1 => n25396, A2 => n25397, ZN => n12995);
   U5449 : AND2_X1 port map( A1 => n27985, A2 => n34008, Z => n6050);
   U1391 : NOR2_X2 port map( A1 => n22126, A2 => n12077, ZN => n22255);
   U7111 : AOI21_X2 port map( A1 => n23027, A2 => n23026, B => n23025, ZN => 
                           n23542);
   U18300 : AOI22_X2 port map( A1 => n37146, A2 => n17225, B1 => n20508, B2 => 
                           n5384, ZN => n15710);
   U2260 : AOI21_X2 port map( A1 => n6045, A2 => n19693, B => n36225, ZN => 
                           n6044);
   U10043 : NAND2_X2 port map( A1 => n22928, A2 => n14817, ZN => n23066);
   U1461 : NAND2_X2 port map( A1 => n3618, A2 => n1990, ZN => n2190);
   U8251 : NAND2_X2 port map( A1 => n24696, A2 => n39196, ZN => n24695);
   U2025 : CLKBUF_X4 port map( I => n4179, Z => n26);
   U324 : INV_X2 port map( I => n27903, ZN => n28181);
   U13768 : OAI21_X2 port map( A1 => n20773, A2 => n21664, B => n1344, ZN => 
                           n4917);
   U16088 : OAI21_X2 port map( A1 => n1300, A2 => n6218, B => n31685, ZN => 
                           n4606);
   U8169 : INV_X2 port map( I => n25380, ZN => n10674);
   U12321 : NAND2_X2 port map( A1 => n25702, A2 => n19296, ZN => n11889);
   U1383 : NAND2_X2 port map( A1 => n1658, A2 => n10037, ZN => n3025);
   U279 : OAI21_X2 port map( A1 => n14585, A2 => n4306, B => n33612, ZN => 
                           n20201);
   U12783 : OAI21_X2 port map( A1 => n14154, A2 => n36757, B => n6298, ZN => 
                           n24277);
   U25154 : OAI22_X2 port map( A1 => n23262, A2 => n23263, B1 => n20867, B2 => 
                           n961, ZN => n16758);
   U841 : INV_X4 port map( I => n10414, ZN => n14410);
   U1833 : INV_X2 port map( I => n33263, ZN => n25939);
   U5849 : INV_X2 port map( I => n29307, ZN => n29389);
   U5862 : AOI22_X2 port map( A1 => n27887, A2 => n39789, B1 => n18687, B2 => 
                           n28175, ZN => n28595);
   U1094 : INV_X2 port map( I => n7319, ZN => n17871);
   U6005 : INV_X2 port map( I => n22599, ZN => n1656);
   U5959 : INV_X2 port map( I => n24696, ZN => n24806);
   U6930 : INV_X4 port map( I => n19863, ZN => n1117);
   U134 : INV_X2 port map( I => n39443, ZN => n29459);
   U6745 : NAND2_X2 port map( A1 => n18904, A2 => n18902, ZN => n26822);
   U9835 : NAND2_X2 port map( A1 => n7399, A2 => n11167, ZN => n23655);
   U9043 : OAI21_X2 port map( A1 => n28282, A2 => n16544, B => n10827, ZN => 
                           n28069);
   U16181 : NAND2_X2 port map( A1 => n13421, A2 => n3670, ZN => n14920);
   U12098 : NOR2_X2 port map( A1 => n25977, A2 => n7258, ZN => n11032);
   U6391 : NAND2_X2 port map( A1 => n22356, A2 => n22353, ZN => n22352);
   U24827 : AOI21_X2 port map( A1 => n22880, A2 => n23034, B => n23035, ZN => 
                           n22882);
   U25819 : NAND2_X2 port map( A1 => n21579, A2 => n11274, ZN => n21707);
   U5857 : INV_X2 port map( I => n28621, ZN => n974);
   U1497 : INV_X2 port map( I => n21506, ZN => n21551);
   U7221 : NOR2_X2 port map( A1 => n22267, A2 => n19515, ZN => n22071);
   U22122 : INV_X2 port map( I => n16500, ZN => n17114);
   U6501 : NAND2_X2 port map( A1 => n8147, A2 => n20720, ZN => n29472);
   U6283 : INV_X4 port map( I => n24874, ZN => n1580);
   U6061 : INV_X2 port map( I => n29475, ZN => n29478);
   U21805 : NAND2_X2 port map( A1 => n17485, A2 => n39666, ZN => n17484);
   U24501 : OAI22_X2 port map( A1 => n12144, A2 => n36887, B1 => n17938, B2 => 
                           n17233, ZN => n17485);
   U5588 : CLKBUF_X4 port map( I => n29495, Z => n18720);
   U558 : INV_X2 port map( I => n38591, ZN => n1500);
   U12741 : INV_X4 port map( I => n10667, ZN => n2731);
   U15485 : INV_X4 port map( I => n3158, ZN => n28246);
   U1728 : NOR2_X2 port map( A1 => n12540, A2 => n12538, ZN => n20642);
   U5892 : NAND2_X2 port map( A1 => n9240, A2 => n9239, ZN => n27131);
   U1382 : NAND2_X2 port map( A1 => n1663, A2 => n3236, ZN => n3237);
   U615 : INV_X2 port map( I => n302, ZN => n5960);
   U265 : NAND2_X2 port map( A1 => n28030, A2 => n28029, ZN => n28390);
   U25429 : INV_X2 port map( I => n21937, ZN => n21939);
   U18209 : OAI21_X2 port map( A1 => n23405, A2 => n5258, B => n9190, ZN => 
                           n23407);
   U1281 : OAI21_X2 port map( A1 => n16892, A2 => n32878, B => n21143, ZN => 
                           n22814);
   U2785 : NOR2_X2 port map( A1 => n4827, A2 => n4620, ZN => n6830);
   U8408 : NAND2_X2 port map( A1 => n23539, A2 => n23337, ZN => n23116);
   U915 : OAI21_X2 port map( A1 => n14168, A2 => n24740, B => n14165, ZN => 
                           n14164);
   U7261 : INV_X4 port map( I => n14493, ZN => n21702);
   U13356 : INV_X2 port map( I => n23592, ZN => n19232);
   U1245 : BUF_X4 port map( I => n23613, Z => n4525);
   U10885 : BUF_X2 port map( I => n29865, Z => n29937);
   U5566 : BUF_X4 port map( I => n20307, Z => n18588);
   U6624 : OAI21_X2 port map( A1 => n14103, A2 => n11876, B => n11875, ZN => 
                           n14760);
   U6333 : NAND2_X2 port map( A1 => n12154, A2 => n6159, ZN => n12153);
   U25235 : OAI21_X2 port map( A1 => n14952, A2 => n25855, B => n34961, ZN => 
                           n16117);
   U14043 : BUF_X2 port map( I => Key(5), Z => n29602);
   U2309 : NAND2_X2 port map( A1 => n10003, A2 => n32258, ZN => n8727);
   U7194 : OAI21_X2 port map( A1 => n18566, A2 => n21449, B => n3676, ZN => 
                           n9225);
   U1536 : INV_X2 port map( I => n20596, ZN => n18926);
   U5900 : OAI21_X2 port map( A1 => n30348, A2 => n2929, B => n36392, ZN => 
                           n7282);
   U6098 : INV_X2 port map( I => n30154, ZN => n30155);
   U28816 : OAI21_X2 port map( A1 => n1288, A2 => n1593, B => n32360, ZN => 
                           n24240);
   U616 : INV_X2 port map( I => n20389, ZN => n26992);
   U12259 : OAI21_X2 port map( A1 => n14589, A2 => n15924, B => n17029, ZN => 
                           n16896);
   U6538 : INV_X4 port map( I => n892, ZN => n9394);
   U7156 : NAND2_X2 port map( A1 => n14560, A2 => n783, ZN => n20518);
   U283 : AOI21_X2 port map( A1 => n2664, A2 => n1206, B => n2663, ZN => n3192)
                           ;
   U6371 : BUF_X2 port map( I => n8943, Z => n5581);
   U940 : NAND2_X2 port map( A1 => n24964, A2 => n3214, ZN => n25022);
   U126 : INV_X2 port map( I => n20524, ZN => n30242);
   U1123 : INV_X2 port map( I => n12758, ZN => n5985);
   U8546 : BUF_X2 port map( I => n22943, Z => n23167);
   U6023 : NAND2_X2 port map( A1 => n11329, A2 => n8519, ZN => n22288);
   U8559 : INV_X2 port map( I => n22676, ZN => n1667);
   U7476 : INV_X2 port map( I => n17225, ZN => n13762);
   U13428 : AOI22_X2 port map( A1 => n23185, A2 => n19538, B1 => n14396, B2 => 
                           n11328, ZN => n14017);
   U96 : INV_X2 port map( I => n20649, ZN => n29940);
   U7847 : AOI21_X2 port map( A1 => n12173, A2 => n31502, B => n12172, ZN => 
                           n12171);
   U3209 : INV_X1 port map( I => n27854, ZN => n1461);
   U7287 : NOR2_X2 port map( A1 => n18205, A2 => n21787, ZN => n21499);
   U8639 : NAND2_X2 port map( A1 => n22086, A2 => n36006, ZN => n22022);
   U393 : INV_X2 port map( I => n20976, ZN => n1077);
   U24537 : AOI22_X2 port map( A1 => n37152, A2 => n17112, B1 => n21508, B2 => 
                           n33852, ZN => n21513);
   U28865 : INV_X4 port map( I => n25048, ZN => n24909);
   U1350 : INV_X2 port map( I => n12471, ZN => n13650);
   U756 : NAND2_X2 port map( A1 => n1098, A2 => n25899, ZN => n10168);
   U8016 : NAND2_X2 port map( A1 => n26016, A2 => n25899, ZN => n26118);
   U7241 : INV_X4 port map( I => n11568, ZN => n19873);
   U11326 : NOR2_X2 port map( A1 => n4809, A2 => n14562, ZN => n2663);
   U13449 : OAI22_X2 port map( A1 => n22554, A2 => n19288, B1 => n22555, B2 => 
                           n22995, ZN => n6970);
   U475 : INV_X2 port map( I => n9037, ZN => n13471);
   U6008 : OAI21_X2 port map( A1 => n4765, A2 => n22136, B => n31412, ZN => 
                           n16347);
   U12289 : AOI21_X2 port map( A1 => n25471, A2 => n25472, B => n2962, ZN => 
                           n25473);
   U5946 : OAI21_X2 port map( A1 => n1118, A2 => n16547, B => n2747, ZN => 
                           n2745);
   U4157 : OAI21_X1 port map( A1 => n29918, A2 => n31570, B => n29916, ZN => 
                           n434);
   U5941 : NOR2_X2 port map( A1 => n39289, A2 => n16246, ZN => n10753);
   U10464 : BUF_X2 port map( I => Key(142), Z => n29838);
   U2266 : AOI21_X2 port map( A1 => n27031, A2 => n27318, B => n16101, ZN => 
                           n27032);
   U4597 : INV_X1 port map( I => n529, ZN => n528);
   U24771 : NAND2_X2 port map( A1 => n37152, A2 => n32544, ZN => n21596);
   U8523 : INV_X1 port map( I => n8628, ZN => n19319);
   U5943 : INV_X2 port map( I => n15883, ZN => n16246);
   U9416 : AOI21_X2 port map( A1 => n19241, A2 => n4602, B => n32979, ZN => 
                           n4400);
   U1352 : INV_X2 port map( I => n30443, ZN => n23045);
   U7055 : NAND2_X2 port map( A1 => n23373, A2 => n23374, ZN => n23376);
   U7113 : INV_X4 port map( I => n16528, ZN => n1302);
   U635 : INV_X2 port map( I => n26252, ZN => n26504);
   U9634 : AOI21_X2 port map( A1 => n6770, A2 => n1565, B => n11957, ZN => 
                           n23826);
   U112 : INV_X4 port map( I => n29455, ZN => n29426);
   U1134 : INV_X2 port map( I => n14290, ZN => n16832);
   U638 : INV_X2 port map( I => n19847, ZN => n1503);
   U16530 : INV_X4 port map( I => n4056, ZN => n5077);
   U12236 : INV_X1 port map( I => n11148, ZN => n1519);
   U10119 : NAND2_X2 port map( A1 => n8744, A2 => n8745, ZN => n9334);
   U5673 : INV_X4 port map( I => n9959, ZN => n910);
   U382 : INV_X2 port map( I => n27674, ZN => n18924);
   U20219 : NAND3_X2 port map( A1 => n1203, A2 => n28419, A3 => n33902, ZN => 
                           n28154);
   U6057 : BUF_X2 port map( I => Key(73), Z => n19937);
   U27638 : NOR2_X2 port map( A1 => n20930, A2 => n20929, ZN => n20928);
   U27690 : NOR2_X2 port map( A1 => n3293, A2 => n19699, ZN => n21489);
   U8511 : NOR2_X2 port map( A1 => n4846, A2 => n23101, ZN => n15638);
   U1456 : NAND2_X2 port map( A1 => n6419, A2 => n6417, ZN => n20351);
   U6440 : INV_X2 port map( I => n20703, ZN => n21550);
   U2045 : INV_X2 port map( I => n33417, ZN => n18374);
   U1537 : INV_X2 port map( I => n21575, ZN => n21594);
   U26110 : OAI21_X1 port map( A1 => n31412, A2 => n35771, B => n16364, ZN => 
                           n16621);
   U1523 : INV_X2 port map( I => n2533, ZN => n17102);
   U10142 : OAI22_X2 port map( A1 => n21985, A2 => n21986, B1 => n37216, B2 => 
                           n20238, ZN => n14754);
   U1043 : NOR2_X2 port map( A1 => n1606, A2 => n626, ZN => n4475);
   U7891 : INV_X2 port map( I => n26994, ZN => n19433);
   U7088 : INV_X4 port map( I => n37774, ZN => n12597);
   U6123 : INV_X2 port map( I => n28595, ZN => n28698);
   U2734 : NAND3_X2 port map( A1 => n22021, A2 => n22020, A3 => n14181, ZN => 
                           n22024);
   U1464 : AOI22_X2 port map( A1 => n1349, A2 => n2280, B1 => n2279, B2 => 
                           n21820, ZN => n237);
   U7102 : INV_X1 port map( I => n32616, ZN => n1291);
   U3833 : INV_X1 port map( I => n35373, ZN => n14939);
   U29291 : OAI22_X2 port map( A1 => n26831, A2 => n38928, B1 => n38852, B2 => 
                           n7752, ZN => n26682);
   U2271 : AOI21_X2 port map( A1 => n12398, A2 => n39037, B => n8036, ZN => 
                           n5287);
   U8644 : AOI22_X2 port map( A1 => n21719, A2 => n32704, B1 => n21720, B2 => 
                           n19647, ZN => n13241);
   U11769 : AOI22_X2 port map( A1 => n8815, A2 => n26951, B1 => n8816, B2 => 
                           n1236, ZN => n16700);
   U8378 : NOR2_X2 port map( A1 => n23508, A2 => n13150, ZN => n13149);
   U8451 : BUF_X4 port map( I => n14856, Z => n10174);
   U10747 : NAND2_X2 port map( A1 => n7749, A2 => n32415, ZN => n10731);
   U5933 : OAI21_X2 port map( A1 => n20216, A2 => n25514, B => n13129, ZN => 
                           n19209);
   U12551 : NAND3_X1 port map( A1 => n8648, A2 => n33412, A3 => n8647, ZN => 
                           n11906);
   U1127 : INV_X2 port map( I => n39814, ZN => n19895);
   U1498 : INV_X2 port map( I => n13473, ZN => n6241);
   U9758 : INV_X2 port map( I => n37934, ZN => n24411);
   U13974 : BUF_X2 port map( I => n21602, Z => n21784);
   U2342 : INV_X2 port map( I => n7993, ZN => n94);
   U6757 : NAND2_X2 port map( A1 => n33952, A2 => n31157, ZN => n26975);
   U8712 : NAND2_X2 port map( A1 => n20544, A2 => n17938, ZN => n21309);
   U24454 : AOI22_X2 port map( A1 => n16448, A2 => n14705, B1 => n16447, B2 => 
                           n12771, ZN => n16446);
   U9500 : INV_X2 port map( I => n31010, ZN => n7853);
   U19660 : INV_X4 port map( I => n23467, ZN => n6969);
   U24804 : NAND2_X2 port map( A1 => n10174, A2 => n23582, ZN => n23581);
   U1436 : NAND2_X2 port map( A1 => n14027, A2 => n2839, ZN => n14037);
   U1413 : OAI21_X2 port map( A1 => n14251, A2 => n19471, B => n22080, ZN => 
                           n16623);
   U8578 : NAND2_X2 port map( A1 => n36731, A2 => n4613, ZN => n22059);
   U5984 : BUF_X4 port map( I => n23296, Z => n23458);
   U6446 : INV_X2 port map( I => n21882, ZN => n21507);
   U394 : BUF_X4 port map( I => n3963, Z => n10653);
   U8708 : INV_X2 port map( I => n21640, ZN => n11411);
   U13358 : NAND2_X2 port map( A1 => n8144, A2 => n8143, ZN => n22927);
   U13597 : INV_X1 port map( I => n1323, ZN => n6473);
   U10435 : INV_X2 port map( I => n14418, ZN => n20544);
   U8030 : OAI21_X2 port map( A1 => n6543, A2 => n25835, B => n31954, ZN => 
                           n9461);
   U8059 : NAND2_X2 port map( A1 => n1522, A2 => n25900, ZN => n26119);
   U24300 : OAI22_X2 port map( A1 => n17333, A2 => n17334, B1 => n17335, B2 => 
                           n14196, ZN => n17942);
   U13963 : OR2_X2 port map( A1 => n21387, A2 => n21743, Z => n21749);
   U10143 : INV_X2 port map( I => n16487, ZN => n5246);
   U15522 : NAND3_X2 port map( A1 => n6345, A2 => n3077, A3 => n6346, ZN => 
                           n23561);
   U8034 : INV_X1 port map( I => n603, ZN => n21041);
   U2980 : NAND2_X2 port map( A1 => n126, A2 => n16495, ZN => n29249);
   U11246 : NOR2_X1 port map( A1 => n27621, A2 => n28149, ZN => n17753);
   U6542 : INV_X2 port map( I => n14179, ZN => n29348);
   U7222 : INV_X2 port map( I => n21961, ZN => n22190);
   U307 : INV_X1 port map( I => n11890, ZN => n27962);
   U5996 : INV_X2 port map( I => n23132, ZN => n23209);
   U2117 : NAND2_X1 port map( A1 => n13268, A2 => n7403, ZN => n13267);
   U10726 : AOI22_X2 port map( A1 => n34070, A2 => n29059, B1 => n30187, B2 => 
                           n7989, ZN => n8202);
   U24133 : OAI22_X2 port map( A1 => n15788, A2 => n25512, B1 => n36991, B2 => 
                           n13744, ZN => n15789);
   U1741 : INV_X1 port map( I => n21674, ZN => n21862);
   U24338 : NAND2_X2 port map( A1 => n14305, A2 => n16463, ZN => n18227);
   U2110 : NAND2_X1 port map( A1 => n22079, A2 => n16625, ZN => n16624);
   U2168 : INV_X4 port map( I => n20309, ZN => n1146);
   U12260 : AOI21_X2 port map( A1 => n21136, A2 => n9161, B => n21135, ZN => 
                           n11251);
   U7012 : NAND2_X2 port map( A1 => n1127, A2 => n24232, ZN => n24332);
   U17878 : NAND2_X1 port map( A1 => n12323, A2 => n11055, ZN => n9313);
   U1121 : INV_X2 port map( I => n15873, ZN => n16366);
   U7597 : INV_X2 port map( I => n28390, ZN => n28486);
   U22098 : INV_X2 port map( I => n15165, ZN => n13076);
   U9561 : INV_X2 port map( I => n30317, ZN => n25512);
   U11872 : INV_X4 port map( I => n19712, ZN => n2140);
   U243 : INV_X1 port map( I => n32535, ZN => n1189);
   U7282 : INV_X4 port map( I => n670, ZN => n21920);
   U12261 : AOI21_X2 port map( A1 => n25383, A2 => n1117, B => n25382, ZN => 
                           n25384);
   U9853 : AOI21_X2 port map( A1 => n23579, A2 => n23581, B => n13831, ZN => 
                           n20946);
   U2666 : OAI21_X2 port map( A1 => n14634, A2 => n15276, B => n40, ZN => 
                           n15772);
   U10000 : OAI21_X2 port map( A1 => n15638, A2 => n1824, B => n13734, ZN => 
                           n6469);
   U6952 : OAI21_X2 port map( A1 => n24824, A2 => n24494, B => n4351, ZN => 
                           n24496);
   U3177 : INV_X1 port map( I => n2799, ZN => n10104);
   U16523 : INV_X2 port map( I => n4048, ZN => n10158);
   U24440 : OAI22_X2 port map( A1 => n22839, A2 => n23103, B1 => n22838, B2 => 
                           n19788, ZN => n22842);
   U12095 : AOI21_X1 port map( A1 => n6783, A2 => n2349, B => n2621, ZN => 
                           n6785);
   U13015 : INV_X4 port map( I => n7834, ZN => n5953);
   U3171 : AOI21_X2 port map( A1 => n12387, A2 => n10019, B => n10193, ZN => 
                           n12364);
   U5820 : INV_X2 port map( I => n21668, ZN => n21845);
   U8445 : BUF_X4 port map( I => n23478, Z => n8692);
   U6667 : INV_X4 port map( I => n14389, ZN => n1074);
   U619 : INV_X2 port map( I => n10523, ZN => n26269);
   U10102 : INV_X4 port map( I => n6327, ZN => n23060);
   U949 : NAND2_X1 port map( A1 => n12385, A2 => n18110, ZN => n4608);
   U12055 : NAND2_X1 port map( A1 => n7677, A2 => n7678, ZN => n4431);
   U12846 : AOI21_X2 port map( A1 => n8360, A2 => n1279, B => n8359, ZN => 
                           n8358);
   U10168 : NAND2_X2 port map( A1 => n22070, A2 => n34452, ZN => n22381);
   U9594 : INV_X2 port map( I => n14164, ZN => n25014);
   U7836 : INV_X4 port map( I => n614, ZN => n15360);
   U957 : OAI21_X2 port map( A1 => n24518, A2 => n39817, B => n18114, ZN => 
                           n12914);
   U6565 : INV_X2 port map( I => n21116, ZN => n9918);
   U22955 : NAND3_X2 port map( A1 => n11378, A2 => n13805, A3 => n39672, ZN => 
                           n18594);
   U9981 : AOI22_X2 port map( A1 => n22893, A2 => n20590, B1 => n22793, B2 => 
                           n9975, ZN => n11671);
   U5869 : INV_X2 port map( I => n27523, ZN => n27674);
   U24388 : INV_X1 port map( I => n10029, ZN => n26672);
   U12466 : NAND2_X2 port map( A1 => n4603, A2 => n5050, ZN => n19965);
   U29860 : NAND2_X2 port map( A1 => n31517, A2 => n29636, ZN => n29638);
   U916 : NAND2_X2 port map( A1 => n14826, A2 => n24845, ZN => n25155);
   U28 : INV_X2 port map( I => n17996, ZN => n30177);
   U6121 : INV_X4 port map( I => n17751, ZN => n11164);
   U335 : INV_X2 port map( I => n34008, ZN => n984);
   U9740 : OAI21_X2 port map( A1 => n9386, A2 => n9519, B => n1606, ZN => n9381
                           );
   U9690 : AOI22_X2 port map( A1 => n24399, A2 => n1587, B1 => n35384, B2 => 
                           n24107, ZN => n24108);
   U11186 : AOI22_X2 port map( A1 => n12787, A2 => n38307, B1 => n12785, B2 => 
                           n12784, ZN => n6926);
   U6664 : INV_X1 port map( I => n9775, ZN => n18948);
   U13477 : NAND2_X2 port map( A1 => n20564, A2 => n23088, ZN => n17083);
   U11196 : NAND2_X1 port map( A1 => n13847, A2 => n7586, ZN => n10394);
   U14227 : OR2_X1 port map( A1 => n14967, A2 => n1874, Z => n2899);
   U23616 : INV_X4 port map( I => n17509, ZN => n24359);
   U2218 : AOI21_X2 port map( A1 => n18459, A2 => n31796, B => n4845, ZN => 
                           n18458);
   U839 : INV_X1 port map( I => n36019, ZN => n7265);
   U10135 : NAND2_X2 port map( A1 => n14036, A2 => n9843, ZN => n22044);
   U13806 : INV_X2 port map( I => n22250, ZN => n8496);
   U898 : INV_X2 port map( I => n25114, ZN => n25267);
   U7549 : INV_X2 port map( I => n7429, ZN => n28740);
   U18790 : INV_X2 port map( I => n5974, ZN => n17464);
   U9241 : INV_X1 port map( I => n27165, ZN => n1223);
   U12293 : NAND2_X2 port map( A1 => n25335, A2 => n31809, ZN => n20464);
   U1455 : INV_X4 port map( I => n7843, ZN => n11329);
   U20471 : NAND2_X1 port map( A1 => n13892, A2 => n38159, ZN => n8734);
   U7022 : OAI21_X2 port map( A1 => n13185, A2 => n12771, B => n14705, ZN => 
                           n12090);
   U6274 : NOR2_X2 port map( A1 => n37105, A2 => n12672, ZN => n12671);
   U12265 : AOI21_X2 port map( A1 => n25476, A2 => n25512, B => n16026, ZN => 
                           n16024);
   U24178 : INV_X1 port map( I => n19085, ZN => n29278);
   U11399 : INV_X1 port map( I => n31571, ZN => n21160);
   U23907 : INV_X4 port map( I => n13316, ZN => n16585);
   U14157 : INV_X2 port map( I => n20284, ZN => n29870);
   U1108 : INV_X4 port map( I => n24244, ZN => n959);
   U24953 : OAI21_X1 port map( A1 => n1235, A2 => n26743, B => n26741, ZN => 
                           n26745);
   U12154 : INV_X2 port map( I => n25876, ZN => n7079);
   U24400 : NAND2_X1 port map( A1 => n24096, A2 => n24478, ZN => n16430);
   U20896 : INV_X4 port map( I => n20359, ZN => n17029);
   U10678 : NAND2_X1 port map( A1 => n6803, A2 => n971, ZN => n29895);
   U13207 : AOI21_X2 port map( A1 => n23522, A2 => n34959, B => n23521, ZN => 
                           n17122);
   U10049 : NAND2_X2 port map( A1 => n32515, A2 => n14409, ZN => n18822);
   U29409 : OAI22_X2 port map( A1 => n27421, A2 => n27420, B1 => n30544, B2 => 
                           n31518, ZN => n27426);
   U21478 : AOI22_X2 port map( A1 => n16236, A2 => n7426, B1 => n23318, B2 => 
                           n23317, ZN => n16235);
   U2608 : INV_X2 port map( I => n19807, ZN => n25);
   U7001 : INV_X8 port map( I => n16585, ZN => n1029);
   U17237 : NAND2_X2 port map( A1 => n31004, A2 => n8304, ZN => n25400);
   U26387 : OR2_X1 port map( A1 => n24265, A2 => n24086, Z => n16311);
   U7114 : INV_X1 port map( I => n14856, ZN => n23506);
   U7127 : INV_X2 port map( I => n23587, ZN => n23325);
   U10974 : NOR2_X2 port map( A1 => n28598, A2 => n39425, ZN => n13718);
   U2267 : INV_X2 port map( I => n6285, ZN => n1211);
   U1467 : AOI22_X2 port map( A1 => n21760, A2 => n21759, B1 => n21758, B2 => 
                           n21757, ZN => n22177);
   U12661 : NOR2_X2 port map( A1 => n5431, A2 => n13495, ZN => n24568);
   U6316 : INV_X2 port map( I => n11449, ZN => n24403);
   U6000 : BUF_X2 port map( I => n23196, Z => n12029);
   U12080 : OAI21_X2 port map( A1 => n4248, A2 => n13885, B => n30937, ZN => 
                           n4247);
   U13124 : OAI21_X2 port map( A1 => n20066, A2 => n21118, B => n19665, ZN => 
                           n7399);
   U5555 : INV_X1 port map( I => n7696, ZN => n20535);
   U8029 : NAND2_X2 port map( A1 => n930, A2 => n7258, ZN => n9228);
   U4472 : INV_X1 port map( I => n29548, ZN => n1394);
   U8344 : NAND2_X2 port map( A1 => n17546, A2 => n19566, ZN => n24129);
   U12279 : OAI22_X2 port map( A1 => n8032, A2 => n12558, B1 => n8034, B2 => 
                           n12557, ZN => n3343);
   U29889 : INV_X1 port map( I => n29750, ZN => n29751);
   U8672 : AOI21_X2 port map( A1 => n17126, A2 => n34021, B => n21731, ZN => 
                           n12511);
   U6227 : INV_X2 port map( I => n25961, ZN => n8711);
   U5614 : INV_X2 port map( I => n19417, ZN => n985);
   U28730 : OAI21_X1 port map( A1 => n24819, A2 => n33412, B => n23824, ZN => 
                           n23825);
   U8783 : BUF_X2 port map( I => Key(180), Z => n30065);
   U6030 : NAND2_X2 port map( A1 => n4242, A2 => n4241, ZN => n22389);
   U5692 : INV_X2 port map( I => n25216, ZN => n13531);
   U8092 : AOI21_X2 port map( A1 => n37071, A2 => n39327, B => n14316, ZN => 
                           n16767);
   U1796 : NAND2_X2 port map( A1 => n13202, A2 => n21053, ZN => n13201);
   U1519 : INV_X2 port map( I => n21742, ZN => n21713);
   U11402 : BUF_X2 port map( I => n27875, Z => n28200);
   U16672 : NAND3_X1 port map( A1 => n28456, A2 => n28099, A3 => n6405, ZN => 
                           n4196);
   U17947 : INV_X1 port map( I => n9668, ZN => n15580);
   U6265 : NAND2_X2 port map( A1 => n1267, A2 => n19422, ZN => n18573);
   U13155 : INV_X1 port map( I => n24051, ZN => n1621);
   U5751 : INV_X1 port map( I => n39070, ZN => n1308);
   U11758 : INV_X2 port map( I => n21101, ZN => n1486);
   U914 : OAI21_X2 port map( A1 => n24580, A2 => n9997, B => n24885, ZN => 
                           n24984);
   U1194 : OAI21_X2 port map( A1 => n3363, A2 => n3366, B => n17122, ZN => 
                           n16488);
   U13459 : OAI21_X2 port map( A1 => n14628, A2 => n16604, B => n22996, ZN => 
                           n8144);
   U12568 : NAND2_X2 port map( A1 => n24568, A2 => n6822, ZN => n21053);
   U8404 : NAND2_X2 port map( A1 => n23488, A2 => n23487, ZN => n23599);
   U10451 : BUF_X2 port map( I => Key(8), Z => n29718);
   U12868 : NAND2_X2 port map( A1 => n11265, A2 => n10694, ZN => n10693);
   U18480 : INV_X2 port map( I => n8395, ZN => n28267);
   U10458 : BUF_X2 port map( I => Key(137), Z => n29394);
   U6454 : BUF_X2 port map( I => Key(108), Z => n29320);
   U14036 : BUF_X2 port map( I => Key(146), Z => n19648);
   U7319 : BUF_X2 port map( I => Key(151), Z => n29970);
   U10450 : BUF_X2 port map( I => Key(163), Z => n29325);
   U7311 : BUF_X2 port map( I => Key(96), Z => n19897);
   U6463 : BUF_X2 port map( I => Key(124), Z => n29983);
   U14047 : BUF_X2 port map( I => Key(110), Z => n19947);
   U5828 : BUF_X2 port map( I => Key(103), Z => n19908);
   U10476 : BUF_X2 port map( I => Key(154), Z => n19903);
   U8782 : BUF_X2 port map( I => Key(16), Z => n19407);
   U7321 : BUF_X2 port map( I => Key(160), Z => n19751);
   U8785 : BUF_X2 port map( I => Key(138), Z => n19890);
   U6472 : BUF_X2 port map( I => Key(70), Z => n19613);
   U6055 : BUF_X2 port map( I => Key(1), Z => n19758);
   U8786 : BUF_X2 port map( I => Key(42), Z => n30010);
   U20017 : BUF_X2 port map( I => Key(98), Z => n19866);
   U10456 : BUF_X2 port map( I => Key(165), Z => n29411);
   U6469 : BUF_X2 port map( I => Key(19), Z => n19860);
   U6457 : BUF_X2 port map( I => Key(82), Z => n19894);
   U6462 : BUF_X2 port map( I => Key(7), Z => n19952);
   U7322 : BUF_X2 port map( I => Key(162), Z => n19845);
   U8780 : BUF_X2 port map( I => Key(79), Z => n19681);
   U6470 : BUF_X2 port map( I => Key(190), Z => n19592);
   U14029 : BUF_X2 port map( I => Key(169), Z => n19820);
   U14027 : BUF_X2 port map( I => Key(13), Z => n19876);
   U14031 : BUF_X2 port map( I => Key(14), Z => n29974);
   U14040 : BUF_X2 port map( I => Key(127), Z => n19833);
   U10442 : BUF_X2 port map( I => Key(141), Z => n29554);
   U8791 : BUF_X2 port map( I => Key(120), Z => n19808);
   U8777 : BUF_X2 port map( I => Key(121), Z => n19774);
   U8788 : BUF_X2 port map( I => Key(50), Z => n29295);
   U6058 : BUF_X2 port map( I => Key(85), Z => n29514);
   U14033 : BUF_X2 port map( I => Key(170), Z => n19910);
   U10462 : BUF_X2 port map( I => Key(39), Z => n19874);
   U14026 : BUF_X2 port map( I => Key(84), Z => n19760);
   U14063 : BUF_X2 port map( I => Key(189), Z => n18270);
   U7316 : BUF_X2 port map( I => Key(46), Z => n19721);
   U8771 : BUF_X2 port map( I => Key(60), Z => n29003);
   U10468 : BUF_X2 port map( I => Key(76), Z => n19877);
   U14068 : BUF_X2 port map( I => Key(25), Z => n29269);
   U8770 : BUF_X2 port map( I => Key(88), Z => n19919);
   U8757 : BUF_X2 port map( I => Key(69), Z => n29978);
   U6455 : BUF_X2 port map( I => Key(130), Z => n19932);
   U10441 : BUF_X2 port map( I => Key(181), Z => n30085);
   U6471 : BUF_X2 port map( I => Key(40), Z => n19527);
   U13991 : INV_X1 port map( I => n29229, ZN => n17705);
   U6046 : BUF_X2 port map( I => n21880, Z => n17112);
   U8736 : INV_X1 port map( I => n19730, ZN => n1362);
   U4582 : CLKBUF_X2 port map( I => n688, Z => n526);
   U3061 : INV_X2 port map( I => n32370, ZN => n19202);
   U28713 : INV_X1 port map( I => n19749, ZN => n29934);
   U14055 : INV_X1 port map( I => n21791, ZN => n1722);
   U6445 : BUF_X2 port map( I => n21368, Z => n21892);
   U1507 : INV_X1 port map( I => n32820, ZN => n918);
   U4668 : CLKBUF_X2 port map( I => n17964, Z => n547);
   U7278 : INV_X2 port map( I => n21684, ZN => n21681);
   U24533 : NAND2_X1 port map( A1 => n21932, A2 => n21931, ZN => n21936);
   U10353 : NAND2_X1 port map( A1 => n6504, A2 => n21476, ZN => n21522);
   U28210 : NOR3_X1 port map( A1 => n21748, A2 => n21712, A3 => n21652, ZN => 
                           n21388);
   U13903 : INV_X1 port map( I => n21718, ZN => n5531);
   U1472 : OAI21_X1 port map( A1 => n3943, A2 => n10961, B => n261, ZN => n3913
                           );
   U8637 : CLKBUF_X4 port map( I => n22350, Z => n19837);
   U13670 : INV_X1 port map( I => n17308, ZN => n21996);
   U16609 : INV_X2 port map( I => n8882, ZN => n9252);
   U8596 : AOI21_X1 port map( A1 => n16266, A2 => n22356, B => n30315, ZN => 
                           n3971);
   U8541 : BUF_X2 port map( I => n22862, Z => n9472);
   U20559 : INV_X1 port map( I => n2046, ZN => n17131);
   U10085 : CLKBUF_X1 port map( I => n23131, Z => n19859);
   U13560 : CLKBUF_X1 port map( I => n19692, Z => n9975);
   U13529 : BUF_X2 port map( I => n18220, Z => n16963);
   U2720 : CLKBUF_X2 port map( I => n3952, Z => n59);
   U5239 : CLKBUF_X2 port map( I => n11643, Z => n3310);
   U2089 : OR2_X1 port map( A1 => n23100, A2 => n21094, Z => n13137);
   U13436 : INV_X1 port map( I => n23146, ZN => n5945);
   U28604 : NAND2_X1 port map( A1 => n23134, A2 => n23133, ZN => n23137);
   U23379 : NAND2_X1 port map( A1 => n23191, A2 => n12163, ZN => n18501);
   U13350 : NAND2_X1 port map( A1 => n5749, A2 => n17917, ZN => n5748);
   U13363 : NAND2_X1 port map( A1 => n5039, A2 => n5038, ZN => n6423);
   U5746 : INV_X2 port map( I => n30881, ZN => n1038);
   U22846 : NOR2_X1 port map( A1 => n23588, A2 => n1306, ZN => n11168);
   U3871 : CLKBUF_X2 port map( I => n23685, Z => n360);
   U1097 : INV_X2 port map( I => n37259, ZN => n13653);
   U13034 : BUF_X2 port map( I => n19341, Z => n9844);
   U13036 : CLKBUF_X2 port map( I => n24196, Z => n19402);
   U8332 : INV_X1 port map( I => n38702, ZN => n24357);
   U12975 : INV_X2 port map( I => n13453, ZN => n8463);
   U3744 : CLKBUF_X2 port map( I => n17844, Z => n326);
   U28824 : NOR2_X1 port map( A1 => n24275, A2 => n17709, ZN => n24278);
   U5711 : INV_X2 port map( I => n24764, ZN => n1269);
   U20984 : NOR2_X1 port map( A1 => n35813, A2 => n8430, ZN => n9257);
   U16273 : NOR2_X1 port map( A1 => n36955, A2 => n24638, ZN => n3751);
   U12525 : INV_X2 port map( I => n24961, ZN => n1555);
   U8199 : BUF_X2 port map( I => n11497, Z => n4664);
   U12473 : BUF_X2 port map( I => n25392, Z => n25689);
   U2696 : OAI21_X1 port map( A1 => n21233, A2 => n9241, B => n12675, ZN => 
                           n25628);
   U28874 : NAND2_X1 port map( A1 => n24553, A2 => n25394, ZN => n24554);
   U22764 : NAND2_X1 port map( A1 => n34583, A2 => n11018, ZN => n14669);
   U9437 : INV_X1 port map( I => n37378, ZN => n8883);
   U17452 : NOR2_X1 port map( A1 => n9380, A2 => n9379, ZN => n4776);
   U591 : INV_X2 port map( I => n861, ZN => n1492);
   U2119 : INV_X1 port map( I => n13854, ZN => n13952);
   U11697 : INV_X1 port map( I => n37245, ZN => n27098);
   U11491 : INV_X1 port map( I => n6818, ZN => n13270);
   U1711 : INV_X1 port map( I => n27407, ZN => n1483);
   U21027 : OR2_X1 port map( A1 => n26889, A2 => n36183, Z => n8485);
   U23096 : NAND2_X1 port map( A1 => n11638, A2 => n11637, ZN => n11639);
   U1651 : INV_X1 port map( I => n37639, ZN => n1459);
   U11456 : INV_X1 port map( I => n27537, ZN => n8865);
   U2863 : CLKBUF_X2 port map( I => n11459, Z => n99);
   U11392 : INV_X1 port map( I => n28101, ZN => n11732);
   U29493 : OAI22_X1 port map( A1 => n27996, A2 => n11461, B1 => n27876, B2 => 
                           n27998, ZN => n27877);
   U11280 : INV_X1 port map( I => n28197, ZN => n8880);
   U23674 : OAI21_X1 port map( A1 => n12807, A2 => n30846, B => n27980, ZN => 
                           n12808);
   U25498 : INV_X1 port map( I => n28324, ZN => n19038);
   U10977 : INV_X1 port map( I => n10305, ZN => n28697);
   U4165 : INV_X1 port map( I => n28382, ZN => n28457);
   U4685 : OAI21_X1 port map( A1 => n552, A2 => n551, B => n36775, ZN => n28477
                           );
   U10999 : NAND2_X1 port map( A1 => n11163, A2 => n28337, ZN => n28338);
   U15169 : INV_X1 port map( I => n3126, ZN => n3127);
   U26306 : INV_X1 port map( I => n14525, ZN => n29353);
   U25319 : INV_X1 port map( I => n35210, ZN => n19193);
   U10782 : NAND2_X1 port map( A1 => n29842, A2 => n21290, ZN => n21289);
   U6084 : CLKBUF_X4 port map( I => n8919, Z => n8918);
   U10735 : NOR2_X1 port map( A1 => n21324, A2 => n3379, ZN => n17877);
   U10716 : NAND2_X1 port map( A1 => n7899, A2 => n18043, ZN => n8228);
   U10439 : CLKBUF_X2 port map( I => Key(66), Z => n19763);
   U7314 : BUF_X2 port map( I => Key(147), Z => n19950);
   U10491 : BUF_X2 port map( I => Key(36), Z => n19817);
   U14054 : BUF_X2 port map( I => Key(176), Z => n29857);
   U6460 : BUF_X2 port map( I => Key(61), Z => n29051);
   U25528 : INV_X1 port map( I => n30253, ZN => n20483);
   U27951 : INV_X1 port map( I => n21628, ZN => n21435);
   U1506 : BUF_X2 port map( I => n18576, Z => n1990);
   U8533 : INV_X1 port map( I => n23196, ZN => n19645);
   U9985 : NOR2_X1 port map( A1 => n22922, A2 => n5838, ZN => n5749);
   U13175 : OAI21_X1 port map( A1 => n20841, A2 => n35506, B => n4968, ZN => 
                           n11530);
   U13121 : INV_X1 port map( I => n23764, ZN => n2044);
   U13047 : BUF_X2 port map( I => n16792, Z => n9963);
   U24173 : INV_X2 port map( I => n13872, ZN => n25261);
   U3643 : BUF_X2 port map( I => n33947, Z => n299);
   U12430 : INV_X2 port map( I => n25695, ZN => n13129);
   U28873 : OAI22_X1 port map( A1 => n19398, A2 => n25681, B1 => n33946, B2 => 
                           n25647, ZN => n24553);
   U29062 : NAND2_X1 port map( A1 => n25515, A2 => n19767, ZN => n25516);
   U29049 : NAND2_X1 port map( A1 => n5886, A2 => n31311, ZN => n25459);
   U27213 : NOR2_X1 port map( A1 => n39112, A2 => n19891, ZN => n20164);
   U8916 : CLKBUF_X2 port map( I => n9393, Z => n5414);
   U5585 : BUF_X2 port map( I => n11348, Z => n10590);
   U9229 : AOI22_X2 port map( A1 => n26710, A2 => n26179, B1 => n11305, B2 => 
                           n1493, ZN => n10595);
   U10997 : NOR2_X2 port map( A1 => n12541, A2 => n11438, ZN => n12540);
   U1730 : NAND2_X2 port map( A1 => n34171, A2 => n11490, ZN => n12541);
   U7990 : AOI21_X2 port map( A1 => n9228, A2 => n25925, B => n9227, ZN => 
                           n9226);
   U27135 : INV_X2 port map( I => n18157, ZN => n21111);
   U8498 : INV_X4 port map( I => n9677, ZN => n13734);
   U8663 : OAI21_X2 port map( A1 => n38438, A2 => n1355, B => n5601, ZN => 
                           n7964);
   U6421 : INV_X1 port map( I => n19387, ZN => n21887);
   U21688 : NOR2_X1 port map( A1 => n9552, A2 => n10629, ZN => n21710);
   U28360 : NAND2_X1 port map( A1 => n1692, A2 => n19337, ZN => n21877);
   U3733 : NOR2_X1 port map( A1 => n31604, A2 => n21667, ZN => n20468);
   U24722 : AOI21_X1 port map( A1 => n18417, A2 => n19542, B => n1157, ZN => 
                           n21533);
   U10359 : NAND2_X1 port map( A1 => n1692, A2 => n19395, ZN => n21874);
   U1500 : INV_X2 port map( I => n21436, ZN => n919);
   U10356 : NOR2_X1 port map( A1 => n21833, A2 => n19620, ZN => n8436);
   U13943 : AOI22_X1 port map( A1 => n19434, A2 => n21484, B1 => n21881, B2 => 
                           n17112, ZN => n13856);
   U28247 : AOI21_X1 port map( A1 => n21678, A2 => n21417, B => n36351, ZN => 
                           n21420);
   U22030 : NAND2_X1 port map( A1 => n17792, A2 => n9809, ZN => n19511);
   U26135 : AOI21_X1 port map( A1 => n15338, A2 => n13855, B => n21579, ZN => 
                           n21580);
   U26692 : NOR2_X1 port map( A1 => n21868, A2 => n15359, ZN => n17992);
   U22925 : NOR2_X1 port map( A1 => n21902, A2 => n35921, ZN => n21623);
   U24513 : AOI21_X1 port map( A1 => n15761, A2 => n21579, B => n36754, ZN => 
                           n15522);
   U26737 : NOR3_X1 port map( A1 => n9642, A2 => n20332, A3 => n21308, ZN => 
                           n20331);
   U1491 : NOR2_X1 port map( A1 => n31604, A2 => n21668, ZN => n21670);
   U10336 : AOI21_X1 port map( A1 => n1158, A2 => n21666, B => n8936, ZN => 
                           n9318);
   U2947 : AOI21_X1 port map( A1 => n3293, A2 => n21892, B => n21894, ZN => 
                           n119);
   U1468 : NAND2_X1 port map( A1 => n10961, A2 => n587, ZN => n6295);
   U2562 : NAND2_X1 port map( A1 => n21834, A2 => n21837, ZN => n9317);
   U24511 : NOR3_X1 port map( A1 => n18417, A2 => n21712, A3 => n1157, ZN => 
                           n19274);
   U26230 : NOR2_X1 port map( A1 => n16302, A2 => n21751, ZN => n15926);
   U28275 : NAND3_X1 port map( A1 => n36728, A2 => n21784, A3 => n32664, ZN => 
                           n21504);
   U10281 : NOR2_X1 port map( A1 => n19037, A2 => n9425, ZN => n21460);
   U24540 : AOI22_X1 port map( A1 => n21621, A2 => n21917, B1 => n33141, B2 => 
                           n18412, ZN => n18900);
   U8613 : INV_X1 port map( I => n22150, ZN => n22151);
   U14928 : INV_X2 port map( I => n8431, ZN => n18567);
   U16434 : INV_X2 port map( I => n39489, ZN => n22327);
   U5789 : NAND2_X1 port map( A1 => n38687, A2 => n22038, ZN => n3835);
   U4927 : NAND2_X1 port map( A1 => n18567, A2 => n8040, ZN => n3682);
   U18583 : NOR2_X1 port map( A1 => n33581, A2 => n915, ZN => n5734);
   U27848 : NOR2_X1 port map( A1 => n1335, A2 => n22310, ZN => n20282);
   U24538 : INV_X1 port map( I => n32675, ZN => n17411);
   U10152 : NOR2_X1 port map( A1 => n22065, A2 => n12077, ZN => n20299);
   U4174 : INV_X1 port map( I => n19773, ZN => n22268);
   U16723 : AOI21_X1 port map( A1 => n12230, A2 => n4240, B => n19873, ZN => 
                           n7815);
   U13668 : NAND2_X1 port map( A1 => n34282, A2 => n13519, ZN => n22309);
   U20323 : AOI21_X1 port map( A1 => n37089, A2 => n22143, B => n8029, ZN => 
                           n8028);
   U27346 : INV_X1 port map( I => n22342, ZN => n18766);
   U28146 : NAND3_X1 port map( A1 => n22307, A2 => n33359, A3 => n1335, ZN => 
                           n21335);
   U13653 : AOI21_X1 port map( A1 => n16499, A2 => n22256, B => n18567, ZN => 
                           n15967);
   U13601 : INV_X2 port map( I => n10488, ZN => n22668);
   U13725 : INV_X1 port map( I => n13704, ZN => n3239);
   U28349 : INV_X1 port map( I => n22572, ZN => n22559);
   U13585 : INV_X1 port map( I => n22508, ZN => n7162);
   U1699 : INV_X1 port map( I => n34073, ZN => n23005);
   U1364 : INV_X1 port map( I => n4997, ZN => n19000);
   U13546 : NOR2_X1 port map( A1 => n12925, A2 => n36369, ZN => n22467);
   U10064 : NAND2_X1 port map( A1 => n12315, A2 => n19645, ZN => n23199);
   U8487 : OAI21_X1 port map( A1 => n16963, A2 => n22915, B => n3310, ZN => 
                           n6712);
   U10021 : NOR2_X1 port map( A1 => n20372, A2 => n5515, ZN => n5785);
   U25742 : NAND2_X1 port map( A1 => n22467, A2 => n22899, ZN => n15201);
   U1299 : INV_X1 port map( I => n23190, ZN => n10828);
   U10024 : NAND2_X1 port map( A1 => n7960, A2 => n19293, ZN => n22917);
   U4706 : NOR2_X1 port map( A1 => n22709, A2 => n18415, ZN => n22861);
   U8524 : INV_X2 port map( I => n33934, ZN => n19538);
   U5987 : NAND3_X1 port map( A1 => n14396, A2 => n17968, A3 => n23186, ZN => 
                           n20302);
   U13439 : NAND3_X1 port map( A1 => n22979, A2 => n22978, A3 => n38524, ZN => 
                           n10471);
   U13420 : NOR2_X1 port map( A1 => n23030, A2 => n5380, ZN => n12509);
   U18105 : NAND2_X1 port map( A1 => n23161, A2 => n5111, ZN => n16887);
   U1259 : INV_X2 port map( I => n23607, ZN => n1637);
   U8394 : OAI21_X1 port map( A1 => n1302, A2 => n5492, B => n5487, ZN => n5491
                           );
   U7062 : AOI21_X1 port map( A1 => n10432, A2 => n13834, B => n1138, ZN => 
                           n9758);
   U27907 : NAND2_X1 port map( A1 => n23576, A2 => n23577, ZN => n20472);
   U28676 : NAND2_X1 port map( A1 => n23567, A2 => n23566, ZN => n23544);
   U20053 : NAND2_X1 port map( A1 => n23324, A2 => n19481, ZN => n7389);
   U23342 : NAND2_X1 port map( A1 => n37523, A2 => n31906, ZN => n12094);
   U13200 : NAND2_X1 port map( A1 => n23638, A2 => n23637, ZN => n3276);
   U8416 : INV_X1 port map( I => n31331, ZN => n1629);
   U13293 : AOI22_X1 port map( A1 => n14901, A2 => n34012, B1 => n23346, B2 => 
                           n35191, ZN => n2814);
   U28588 : NAND3_X1 port map( A1 => n23364, A2 => n9078, A3 => n23361, ZN => 
                           n23018);
   U28681 : AOI21_X1 port map( A1 => n23611, A2 => n23610, B => n38611, ZN => 
                           n23616);
   U3543 : NOR2_X1 port map( A1 => n18866, A2 => n34959, ZN => n3365);
   U5976 : INV_X2 port map( I => n2117, ZN => n14491);
   U6315 : INV_X1 port map( I => n24369, ZN => n24087);
   U5539 : INV_X1 port map( I => n24421, ZN => n24419);
   U1058 : NAND2_X1 port map( A1 => n24432, A2 => n24431, ZN => n21125);
   U9812 : INV_X1 port map( I => n30320, ZN => n24392);
   U24855 : OAI21_X1 port map( A1 => n17546, A2 => n24465, B => n24316, ZN => 
                           n18346);
   U5034 : AOI21_X1 port map( A1 => n1602, A2 => n16779, B => n9922, ZN => 
                           n14052);
   U25804 : NAND2_X1 port map( A1 => n15320, A2 => n20312, ZN => n15319);
   U3529 : AOI21_X1 port map( A1 => n13453, A2 => n9066, B => n12248, ZN => 
                           n9068);
   U5965 : NAND2_X1 port map( A1 => n24338, A2 => n12953, ZN => n10421);
   U5729 : NOR2_X1 port map( A1 => n18697, A2 => n20027, ZN => n24147);
   U1029 : NAND2_X1 port map( A1 => n24814, A2 => n24623, ZN => n24734);
   U970 : NOR2_X1 port map( A1 => n24529, A2 => n5897, ZN => n24530);
   U6278 : INV_X1 port map( I => n33230, ZN => n19431);
   U5285 : INV_X1 port map( I => n24735, ZN => n24852);
   U6982 : NAND2_X1 port map( A1 => n17618, A2 => n7529, ZN => n24494);
   U28884 : NOR2_X1 port map( A1 => n16238, A2 => n35981, ZN => n24596);
   U12611 : NAND2_X1 port map( A1 => n6822, A2 => n5431, ZN => n9478);
   U22153 : NAND2_X1 port map( A1 => n18845, A2 => n36376, ZN => n18844);
   U9660 : NAND2_X1 port map( A1 => n14267, A2 => n19431, ZN => n14266);
   U26524 : NOR2_X1 port map( A1 => n39681, A2 => n7552, ZN => n24715);
   U19083 : NAND2_X1 port map( A1 => n6337, A2 => n19484, ZN => n6336);
   U12642 : NAND2_X1 port map( A1 => n6186, A2 => n1026, ZN => n6184);
   U25204 : INV_X1 port map( I => n24532, ZN => n24618);
   U17943 : NAND3_X1 port map( A1 => n38674, A2 => n38668, A3 => n5124, ZN => 
                           n5122);
   U9655 : NOR2_X1 port map( A1 => n31845, A2 => n1026, ZN => n13583);
   U9619 : NAND2_X1 port map( A1 => n37106, A2 => n5431, ZN => n9500);
   U23403 : OAI22_X1 port map( A1 => n20301, A2 => n19886, B1 => n24566, B2 => 
                           n12159, ZN => n12208);
   U19609 : INV_X2 port map( I => n37052, ZN => n13943);
   U22529 : INV_X1 port map( I => n10584, ZN => n17774);
   U25559 : NOR2_X1 port map( A1 => n18880, A2 => n20359, ZN => n14778);
   U9572 : INV_X1 port map( I => n25631, ZN => n25728);
   U29068 : NAND2_X1 port map( A1 => n25550, A2 => n25549, ZN => n25556);
   U6896 : NOR2_X1 port map( A1 => n25550, A2 => n1537, ZN => n11066);
   U8118 : NOR2_X1 port map( A1 => n13943, A2 => n16264, ZN => n14100);
   U12385 : NOR2_X1 port map( A1 => n9800, A2 => n14460, ZN => n9482);
   U16100 : NAND2_X1 port map( A1 => n3602, A2 => n34755, ZN => n25346);
   U2599 : INV_X1 port map( I => n25157, ZN => n9915);
   U2179 : INV_X1 port map( I => n835, ZN => n1543);
   U2652 : NOR2_X1 port map( A1 => n33785, A2 => n25623, ZN => n17075);
   U1838 : NAND2_X1 port map( A1 => n7238, A2 => n19237, ZN => n7237);
   U21225 : NAND3_X1 port map( A1 => n20855, A2 => n1546, A3 => n19589, ZN => 
                           n14262);
   U757 : INV_X1 port map( I => n25836, ZN => n18375);
   U739 : INV_X1 port map( I => n21204, ZN => n1512);
   U15899 : INV_X1 port map( I => n33644, ZN => n25934);
   U27387 : NOR2_X1 port map( A1 => n1528, A2 => n1245, ZN => n20134);
   U20192 : INV_X1 port map( I => n25849, ZN => n25888);
   U744 : NAND2_X1 port map( A1 => n834, A2 => n1245, ZN => n4769);
   U9436 : NAND2_X1 port map( A1 => n1011, A2 => n6056, ZN => n3838);
   U6206 : OR2_X1 port map( A1 => n17008, A2 => n11533, Z => n9892);
   U19144 : NAND3_X1 port map( A1 => n25850, A2 => n25851, A3 => n928, ZN => 
                           n6398);
   U28988 : NAND2_X1 port map( A1 => n25996, A2 => n25994, ZN => n25112);
   U9421 : OAI21_X1 port map( A1 => n6056, A2 => n4382, B => n4381, ZN => n2124
                           );
   U26842 : NOR2_X1 port map( A1 => n7767, A2 => n33263, ZN => n20611);
   U4889 : AOI21_X1 port map( A1 => n26213, A2 => n9868, B => n26212, ZN => 
                           n14503);
   U9345 : INV_X1 port map( I => n26968, ZN => n19338);
   U2010 : NAND2_X1 port map( A1 => n36344, A2 => n860, ZN => n26622);
   U19421 : NOR3_X1 port map( A1 => n862, A2 => n26639, A3 => n17515, ZN => 
                           n12177);
   U24957 : NOR2_X1 port map( A1 => n26847, A2 => n10314, ZN => n20316);
   U570 : NOR2_X1 port map( A1 => n39823, A2 => n17237, ZN => n17323);
   U11851 : NAND2_X1 port map( A1 => n20699, A2 => n9179, ZN => n16177);
   U24962 : INV_X1 port map( I => n19371, ZN => n16222);
   U9328 : NOR2_X1 port map( A1 => n26830, A2 => n26959, ZN => n6909);
   U26161 : NAND2_X1 port map( A1 => n19332, A2 => n26740, ZN => n27014);
   U24922 : AOI21_X1 port map( A1 => n11616, A2 => n26751, B => n26752, ZN => 
                           n17229);
   U7852 : NOR2_X1 port map( A1 => n26898, A2 => n39287, ZN => n27043);
   U24997 : NAND2_X1 port map( A1 => n20575, A2 => n20576, ZN => n20574);
   U9290 : NOR2_X1 port map( A1 => n11707, A2 => n36391, ZN => n12987);
   U524 : OAI21_X1 port map( A1 => n11674, A2 => n16522, B => n19425, ZN => 
                           n10535);
   U7832 : INV_X1 port map( I => n8988, ZN => n8830);
   U3326 : OAI21_X1 port map( A1 => n31254, A2 => n20699, B => n212, ZN => 
                           n10796);
   U29230 : AOI21_X1 port map( A1 => n26724, A2 => n16970, B => n26627, ZN => 
                           n26372);
   U19038 : INV_X2 port map( I => n9369, ZN => n20133);
   U22471 : NAND2_X1 port map( A1 => n10461, A2 => n12156, ZN => n17720);
   U441 : INV_X1 port map( I => n18047, ZN => n1085);
   U2627 : INV_X1 port map( I => n17072, ZN => n27201);
   U517 : INV_X1 port map( I => n7424, ZN => n16946);
   U15504 : NAND2_X1 port map( A1 => n31518, A2 => n3059, ZN => n26953);
   U29411 : NAND2_X1 port map( A1 => n30412, A2 => n19719, ZN => n27445);
   U25318 : NOR2_X1 port map( A1 => n27092, A2 => n16043, ZN => n19077);
   U29112 : NOR2_X1 port map( A1 => n27069, A2 => n31433, ZN => n26074);
   U25259 : NAND2_X1 port map( A1 => n17720, A2 => n35427, ZN => n17719);
   U11731 : INV_X2 port map( I => n997, ZN => n1474);
   U29389 : OAI21_X1 port map( A1 => n27436, A2 => n27235, B => n27234, ZN => 
                           n27236);
   U11439 : INV_X1 port map( I => n27776, ZN => n27705);
   U23394 : INV_X2 port map( I => n12187, ZN => n28114);
   U26252 : INV_X1 port map( I => n32932, ZN => n28248);
   U7695 : NOR2_X1 port map( A1 => n28024, A2 => n20739, ZN => n28022);
   U9052 : NOR2_X1 port map( A1 => n7690, A2 => n2877, ZN => n2876);
   U342 : NAND3_X1 port map( A1 => n8523, A2 => n27901, A3 => n27996, ZN => 
                           n28403);
   U20312 : NAND3_X1 port map( A1 => n39574, A2 => n99, A3 => n19366, ZN => 
                           n7586);
   U6642 : NAND3_X1 port map( A1 => n11283, A2 => n36854, A3 => n3662, ZN => 
                           n2872);
   U1737 : AOI21_X1 port map( A1 => n19366, A2 => n28230, B => n12257, ZN => 
                           n28232);
   U9066 : NOR2_X1 port map( A1 => n28079, A2 => n1070, ZN => n7431);
   U9082 : NOR3_X1 port map( A1 => n3159, A2 => n28248, A3 => n28246, ZN => 
                           n3065);
   U24994 : NAND2_X1 port map( A1 => n28187, A2 => n16325, ZN => n16063);
   U11185 : NAND2_X1 port map( A1 => n33959, A2 => n6236, ZN => n3794);
   U29641 : NOR2_X1 port map( A1 => n30716, A2 => n180, ZN => n28664);
   U19163 : INV_X2 port map( I => n6426, ZN => n28759);
   U204 : INV_X2 port map( I => n28330, ZN => n1186);
   U2672 : INV_X1 port map( I => n28478, ZN => n3532);
   U6631 : INV_X1 port map( I => n36478, ZN => n1427);
   U11121 : INV_X1 port map( I => n28580, ZN => n13825);
   U24106 : NOR2_X1 port map( A1 => n39724, A2 => n18871, ZN => n14489);
   U259 : INV_X1 port map( I => n33100, ZN => n1415);
   U169 : AOI22_X1 port map( A1 => n17771, A2 => n31378, B1 => n12061, B2 => 
                           n9355, ZN => n309);
   U10973 : AOI22_X1 port map( A1 => n11488, A2 => n34007, B1 => n1189, B2 => 
                           n28528, ZN => n8853);
   U15257 : NAND3_X1 port map( A1 => n28501, A2 => n38145, A3 => n2790, ZN => 
                           n2789);
   U8961 : NAND2_X1 port map( A1 => n28515, A2 => n5093, ZN => n4429);
   U22712 : NAND2_X1 port map( A1 => n33318, A2 => n13508, ZN => n11869);
   U27685 : OAI21_X1 port map( A1 => n1420, A2 => n37204, B => n19668, ZN => 
                           n28568);
   U4486 : INV_X1 port map( I => n28463, ZN => n28641);
   U25301 : NAND3_X1 port map( A1 => n28495, A2 => n35173, A3 => n28356, ZN => 
                           n28357);
   U2247 : INV_X1 port map( I => n29042, ZN => n15480);
   U2236 : INV_X1 port map( I => n9393, ZN => n21299);
   U8921 : INV_X1 port map( I => n14076, ZN => n16116);
   U8911 : INV_X1 port map( I => n29344, ZN => n29481);
   U16871 : INV_X1 port map( I => n4392, ZN => n19693);
   U7439 : INV_X2 port map( I => n14400, ZN => n1401);
   U6572 : INV_X2 port map( I => n14559, ZN => n1181);
   U20669 : INV_X2 port map( I => n29195, ZN => n29702);
   U10828 : INV_X1 port map( I => n9716, ZN => n13136);
   U4263 : INV_X1 port map( I => n6163, ZN => n29182);
   U10789 : OAI21_X1 port map( A1 => n33784, A2 => n30241, B => n6443, ZN => 
                           n5306);
   U23491 : AOI21_X1 port map( A1 => n29287, A2 => n29286, B => n17225, ZN => 
                           n12372);
   U29742 : NAND2_X1 port map( A1 => n29102, A2 => n1175, ZN => n29103);
   U23554 : INV_X2 port map( I => n30178, ZN => n30183);
   U25 : INV_X1 port map( I => n18896, ZN => n18897);
   U8836 : INV_X1 port map( I => n30184, ZN => n16676);
   U32 : INV_X1 port map( I => n30097, ZN => n1380);
   U7379 : INV_X1 port map( I => n29855, ZN => n1171);
   U5838 : INV_X1 port map( I => n2858, ZN => n3725);
   U4996 : NOR3_X1 port map( A1 => n633, A2 => n1171, A3 => n32258, ZN => n9676
                           );
   U3 : AND2_X1 port map( A1 => n12979, A2 => n29220, Z => n9606);
   U19 : INV_X1 port map( I => n20538, ZN => n30822);
   U40 : INV_X1 port map( I => n30079, ZN => n30793);
   U43 : INV_X1 port map( I => n6205, ZN => n1054);
   U64 : NAND2_X1 port map( A1 => n31717, A2 => n14788, ZN => n31532);
   U82 : NOR2_X1 port map( A1 => n621, A2 => n20616, ZN => n4075);
   U88 : AND2_X1 port map( A1 => n29481, A2 => n29454, Z => n29425);
   U91 : OAI21_X1 port map( A1 => n39392, A2 => n12081, B => n29061, ZN => n400
                           );
   U92 : NAND3_X1 port map( A1 => n32894, A2 => n3986, A3 => n621, ZN => n31170
                           );
   U135 : NAND2_X1 port map( A1 => n29445, A2 => n29446, ZN => n5336);
   U137 : NAND2_X1 port map( A1 => n8726, A2 => n29346, ZN => n29349);
   U139 : NAND2_X1 port map( A1 => n29384, A2 => n11084, ZN => n31280);
   U162 : AOI21_X1 port map( A1 => n29591, A2 => n29592, B => n29598, ZN => 
                           n31374);
   U181 : NAND2_X1 port map( A1 => n11389, A2 => n9955, ZN => n31550);
   U191 : NAND2_X1 port map( A1 => n31313, A2 => n89, ZN => n5543);
   U269 : NAND2_X1 port map( A1 => n6405, A2 => n28434, ZN => n31389);
   U270 : NAND2_X1 port map( A1 => n7324, A2 => n28617, ZN => n30857);
   U274 : NOR2_X1 port map( A1 => n3014, A2 => n6426, ZN => n32274);
   U362 : AND2_X1 port map( A1 => n1446, A2 => n20577, Z => n30357);
   U364 : OR2_X1 port map( A1 => n28114, A2 => n28248, Z => n30293);
   U372 : NAND2_X1 port map( A1 => n32963, A2 => n33321, ZN => n18341);
   U391 : NAND3_X1 port map( A1 => n3983, A2 => n19996, A3 => n28279, ZN => 
                           n7186);
   U397 : NOR2_X1 port map( A1 => n5062, A2 => n28194, ZN => n5910);
   U398 : NAND2_X1 port map( A1 => n33669, A2 => n2877, ZN => n33959);
   U410 : NOR2_X1 port map( A1 => n28050, A2 => n11891, ZN => n32479);
   U422 : NAND3_X1 port map( A1 => n1453, A2 => n982, A3 => n2302, ZN => n3097)
                           ;
   U429 : NOR2_X1 port map( A1 => n28246, A2 => n28247, ZN => n32657);
   U447 : NAND2_X1 port map( A1 => n27888, A2 => n28238, ZN => n33199);
   U452 : NOR2_X1 port map( A1 => n1072, A2 => n34008, ZN => n14263);
   U455 : INV_X1 port map( I => n27948, ZN => n33321);
   U462 : NAND2_X1 port map( A1 => n1074, A2 => n28181, ZN => n30799);
   U466 : NOR2_X1 port map( A1 => n13081, A2 => n14399, ZN => n12475);
   U486 : NAND2_X1 port map( A1 => n1202, A2 => n11676, ZN => n33931);
   U500 : NAND2_X1 port map( A1 => n28102, A2 => n32352, ZN => n33201);
   U516 : INV_X1 port map( I => n9470, ZN => n8960);
   U528 : NOR2_X1 port map( A1 => n28238, A2 => n1453, ZN => n33202);
   U539 : BUF_X2 port map( I => n28153, Z => n33481);
   U563 : BUF_X2 port map( I => n10009, Z => n9534);
   U581 : INV_X1 port map( I => n27631, ZN => n31218);
   U654 : NAND2_X1 port map( A1 => n7606, A2 => n16520, ZN => n16514);
   U715 : NOR2_X1 port map( A1 => n31006, A2 => n17072, ZN => n31399);
   U723 : NOR2_X1 port map( A1 => n16482, A2 => n5772, ZN => n31680);
   U767 : AND2_X1 port map( A1 => n30986, A2 => n35427, Z => n3605);
   U810 : OR2_X1 port map( A1 => n26687, A2 => n17097, Z => n30335);
   U812 : OR2_X1 port map( A1 => n26979, A2 => n852, Z => n30352);
   U843 : OAI22_X1 port map( A1 => n27014, A2 => n11679, B1 => n27013, B2 => 
                           n38577, ZN => n32549);
   U846 : NAND2_X1 port map( A1 => n26815, A2 => n26973, ZN => n26816);
   U849 : AOI21_X1 port map( A1 => n20699, A2 => n849, B => n7516, ZN => n212);
   U854 : NOR2_X1 port map( A1 => n26718, A2 => n735, ZN => n33303);
   U855 : NOR2_X1 port map( A1 => n13393, A2 => n26764, ZN => n32669);
   U868 : NOR2_X1 port map( A1 => n16160, A2 => n866, ZN => n17279);
   U902 : AOI21_X1 port map( A1 => n18226, A2 => n26833, B => n26628, ZN => 
                           n30983);
   U942 : INV_X1 port map( I => n26899, ZN => n32016);
   U963 : NOR2_X1 port map( A1 => n875, A2 => n26937, ZN => n11325);
   U964 : NAND2_X1 port map( A1 => n26752, A2 => n26751, ZN => n33708);
   U979 : OR2_X1 port map( A1 => n26818, A2 => n4599, Z => n13219);
   U1022 : NAND2_X1 port map( A1 => n31919, A2 => n4769, ZN => n8295);
   U1032 : OAI21_X1 port map( A1 => n10179, A2 => n10180, B => n1101, ZN => 
                           n20116);
   U1049 : AOI21_X1 port map( A1 => n603, A2 => n34961, B => n26005, ZN => 
                           n33891);
   U1059 : NAND2_X2 port map( A1 => n20849, A2 => n5236, ZN => n2150);
   U1075 : NAND2_X1 port map( A1 => n7767, A2 => n8481, ZN => n31919);
   U1083 : NOR2_X1 port map( A1 => n15085, A2 => n15121, ZN => n10180);
   U1096 : NAND2_X1 port map( A1 => n36546, A2 => n31192, ZN => n30547);
   U1106 : NAND2_X1 port map( A1 => n26063, A2 => n25345, ZN => n25348);
   U1110 : NOR2_X1 port map( A1 => n26063, A2 => n26061, ZN => n33465);
   U1113 : NOR2_X1 port map( A1 => n17212, A2 => n7767, ZN => n25818);
   U1119 : NAND2_X1 port map( A1 => n16407, A2 => n18320, ZN => n25586);
   U1126 : NOR2_X1 port map( A1 => n36666, A2 => n5126, ZN => n4867);
   U1169 : NAND2_X1 port map( A1 => n35138, A2 => n33514, ZN => n2942);
   U1182 : NOR2_X1 port map( A1 => n603, A2 => n12548, ZN => n30695);
   U1198 : NAND2_X1 port map( A1 => n30625, A2 => n6939, ZN => n7136);
   U1199 : OAI21_X1 port map( A1 => n31388, A2 => n31386, B => n25755, ZN => 
                           n25758);
   U1207 : OAI21_X1 port map( A1 => n25008, A2 => n20052, B => n10082, ZN => 
                           n30625);
   U1211 : NOR2_X1 port map( A1 => n25753, A2 => n38338, ZN => n31388);
   U1222 : OAI21_X1 port map( A1 => n31809, A2 => n25460, B => n17183, ZN => 
                           n31843);
   U1233 : NOR2_X1 port map( A1 => n25337, A2 => n12828, ZN => n31842);
   U1263 : NAND2_X1 port map( A1 => n25469, A2 => n25468, ZN => n30936);
   U1266 : NAND2_X1 port map( A1 => n3568, A2 => n38661, ZN => n11243);
   U1280 : NOR2_X1 port map( A1 => n4384, A2 => n37795, ZN => n25536);
   U1307 : NOR2_X1 port map( A1 => n2250, A2 => n15515, ZN => n33250);
   U1308 : NOR2_X1 port map( A1 => n15422, A2 => n14779, ZN => n3319);
   U1329 : AND2_X1 port map( A1 => n3568, A2 => n5051, Z => n30388);
   U1373 : NAND2_X1 port map( A1 => n25615, A2 => n19264, ZN => n33648);
   U1493 : BUF_X2 port map( I => n25132, Z => n33208);
   U1528 : NAND2_X1 port map( A1 => n37852, A2 => n24866, ZN => n6934);
   U1545 : NOR2_X1 port map( A1 => n30843, A2 => n31861, ZN => n33125);
   U1553 : OAI21_X1 port map( A1 => n30948, A2 => n30947, B => n1271, ZN => 
                           n24502);
   U1557 : NOR2_X1 port map( A1 => n24759, A2 => n12633, ZN => n32971);
   U1559 : NAND2_X1 port map( A1 => n24621, A2 => n10116, ZN => n32062);
   U1561 : AND2_X1 port map( A1 => n8173, A2 => n30464, Z => n24771);
   U1563 : NAND2_X1 port map( A1 => n24824, A2 => n30845, ZN => n24387);
   U1569 : AND2_X1 port map( A1 => n36321, A2 => n7445, Z => n8804);
   U1584 : NOR2_X1 port map( A1 => n1581, A2 => n7770, ZN => n12681);
   U1593 : AND2_X1 port map( A1 => n31650, A2 => n17806, Z => n31530);
   U1594 : NAND2_X1 port map( A1 => n3076, A2 => n24668, ZN => n30915);
   U1595 : INV_X2 port map( I => n2341, ZN => n24664);
   U1602 : NOR2_X1 port map( A1 => n24680, A2 => n24883, ZN => n6707);
   U1616 : NAND2_X1 port map( A1 => n19828, A2 => n30464, ZN => n32618);
   U1617 : NAND3_X1 port map( A1 => n38194, A2 => n36471, A3 => n35901, ZN => 
                           n24574);
   U1685 : NAND2_X1 port map( A1 => n23817, A2 => n37134, ZN => n30766);
   U1692 : OAI21_X1 port map( A1 => n17709, A2 => n14378, B => n1586, ZN => 
                           n11317);
   U1701 : NAND2_X1 port map( A1 => n37732, A2 => n20083, ZN => n31044);
   U1702 : OAI21_X1 port map( A1 => n16366, A2 => n24406, B => n18920, ZN => 
                           n31175);
   U1715 : NAND2_X1 port map( A1 => n21043, A2 => n32899, ZN => n24424);
   U1732 : NAND2_X1 port map( A1 => n32742, A2 => n4986, ZN => n32741);
   U1735 : NAND2_X1 port map( A1 => n16918, A2 => n30927, ZN => n23993);
   U1743 : NAND2_X1 port map( A1 => n24478, A2 => n24479, ZN => n32784);
   U1744 : NAND2_X1 port map( A1 => n12975, A2 => n24433, ZN => n30646);
   U1749 : NOR2_X1 port map( A1 => n1282, A2 => n20404, ZN => n31921);
   U1752 : AOI21_X1 port map( A1 => n626, A2 => n24245, B => n959, ZN => n24094
                           );
   U1754 : NAND2_X1 port map( A1 => n17546, A2 => n24465, ZN => n33904);
   U1755 : NAND2_X1 port map( A1 => n30463, A2 => n30580, ZN => n31102);
   U1772 : AND2_X1 port map( A1 => n10477, A2 => n30311, Z => n32786);
   U1778 : BUF_X2 port map( I => n19295, Z => n32899);
   U1793 : INV_X1 port map( I => n30280, ZN => n30320);
   U1856 : OAI21_X1 port map( A1 => n21019, A2 => n23467, B => n31223, ZN => 
                           n23422);
   U1861 : NAND3_X1 port map( A1 => n1310, A2 => n35232, A3 => n14011, ZN => 
                           n13580);
   U1870 : NAND3_X1 port map( A1 => n35367, A2 => n23577, A3 => n20955, ZN => 
                           n20954);
   U1874 : AND2_X1 port map( A1 => n23631, A2 => n11342, Z => n20841);
   U1887 : NAND2_X1 port map( A1 => n23355, A2 => n31749, ZN => n14576);
   U1920 : OAI21_X1 port map( A1 => n32798, A2 => n23455, B => n33080, ZN => 
                           n20984);
   U1935 : AND2_X1 port map( A1 => n33496, A2 => n23619, Z => n30460);
   U1946 : OAI21_X1 port map( A1 => n23552, A2 => n37814, B => n14163, ZN => 
                           n30548);
   U1957 : AOI21_X1 port map( A1 => n22845, A2 => n22682, B => n15242, ZN => 
                           n15771);
   U1963 : INV_X1 port map( I => n3256, ZN => n5492);
   U1971 : INV_X1 port map( I => n23121, ZN => n9238);
   U1974 : NAND2_X1 port map( A1 => n31351, A2 => n33247, ZN => n19521);
   U1979 : NAND3_X1 port map( A1 => n23175, A2 => n121, A3 => n3803, ZN => 
                           n11472);
   U1984 : AOI22_X1 port map( A1 => n23149, A2 => n1146, B1 => n14234, B2 => 
                           n38604, ZN => n10699);
   U1989 : NAND2_X1 port map( A1 => n22709, A2 => n1651, ZN => n15344);
   U1991 : OAI21_X1 port map( A1 => n14409, A2 => n32677, B => n32676, ZN => 
                           n23207);
   U2016 : NOR2_X1 port map( A1 => n14396, A2 => n33745, ZN => n9770);
   U2017 : NOR2_X1 port map( A1 => n18515, A2 => n19945, ZN => n32216);
   U2018 : NOR2_X1 port map( A1 => n19698, A2 => n23101, ZN => n33074);
   U2035 : NOR2_X1 port map( A1 => n32636, A2 => n23149, ZN => n12239);
   U2036 : OAI21_X1 port map( A1 => n15033, A2 => n22932, B => n39527, ZN => 
                           n15032);
   U2050 : INV_X1 port map( I => n22559, ZN => n33694);
   U2051 : INV_X1 port map( I => n12437, ZN => n22575);
   U2068 : NOR2_X1 port map( A1 => n22676, A2 => n1670, ZN => n17341);
   U2084 : NAND3_X1 port map( A1 => n22299, A2 => n22301, A3 => n22300, ZN => 
                           n22302);
   U2103 : INV_X1 port map( I => n30818, ZN => n30817);
   U2108 : INV_X1 port map( I => n22262, ZN => n22125);
   U2123 : NOR2_X1 port map( A1 => n3003, A2 => n22229, ZN => n31859);
   U2124 : AOI21_X1 port map( A1 => n22234, A2 => n20351, B => n7497, ZN => 
                           n33859);
   U2130 : INV_X1 port map( I => n33678, ZN => n16635);
   U2139 : INV_X2 port map( I => n22234, ZN => n33860);
   U2164 : AOI21_X1 port map( A1 => n19377, A2 => n19376, B => n21894, ZN => 
                           n21369);
   U2166 : NOR2_X1 port map( A1 => n21670, A2 => n6198, ZN => n33636);
   U2167 : AND2_X1 port map( A1 => n35921, A2 => n21903, Z => n30397);
   U2171 : NOR2_X1 port map( A1 => n14424, A2 => n21788, ZN => n32857);
   U2181 : NOR2_X1 port map( A1 => n18417, A2 => n30731, ZN => n31975);
   U2188 : NOR2_X1 port map( A1 => n31335, A2 => n21888, ZN => n21333);
   U2197 : NAND2_X1 port map( A1 => n35921, A2 => n18152, ZN => n33731);
   U2211 : NOR2_X2 port map( A1 => n38782, A2 => n16677, ZN => n17816);
   U2220 : INV_X2 port map( I => n5871, ZN => n24738);
   U2230 : NAND2_X2 port map( A1 => n16990, A2 => n5871, ZN => n7847);
   U2232 : INV_X2 port map( I => n15350, ZN => n21987);
   U2262 : NAND2_X2 port map( A1 => n18831, A2 => n25557, ZN => n13988);
   U2265 : NOR2_X2 port map( A1 => n30851, A2 => n35904, ZN => n19569);
   U2270 : INV_X2 port map( I => n25718, ZN => n25563);
   U2281 : INV_X2 port map( I => n14350, ZN => n25009);
   U2308 : BUF_X4 port map( I => n21445, Z => n21847);
   U2317 : OAI21_X2 port map( A1 => n10374, A2 => n12671, B => n25048, ZN => 
                           n10373);
   U2330 : CLKBUF_X4 port map( I => n30095, Z => n6147);
   U2377 : NAND2_X1 port map( A1 => n14076, A2 => n29493, ZN => n29451);
   U2387 : NAND2_X1 port map( A1 => n4083, A2 => n30195, ZN => n1757);
   U2405 : AOI21_X1 port map( A1 => n12320, A2 => n29441, B => n12317, ZN => 
                           n12316);
   U2422 : NOR2_X1 port map( A1 => n28089, A2 => n288, ZN => n8206);
   U2431 : AOI22_X1 port map( A1 => n26826, A2 => n26825, B1 => n19442, B2 => 
                           n19762, ZN => n20022);
   U2435 : OAI21_X1 port map( A1 => n31283, A2 => n9249, B => n3700, ZN => 
                           n9248);
   U2445 : NAND2_X1 port map( A1 => n9716, A2 => n1061, ZN => n32649);
   U2453 : NAND3_X1 port map( A1 => n6818, A2 => n1798, A3 => n33803, ZN => 
                           n13292);
   U2485 : AOI21_X1 port map( A1 => n3860, A2 => n29927, B => n19097, ZN => 
                           n29925);
   U2490 : NAND2_X1 port map( A1 => n14949, A2 => n17072, ZN => n17298);
   U2499 : AOI21_X1 port map( A1 => n16917, A2 => n24443, B => n1596, ZN => 
                           n30927);
   U2516 : AOI21_X1 port map( A1 => n6684, A2 => n6421, B => n1637, ZN => 
                           n23216);
   U2524 : BUF_X2 port map( I => Key(41), Z => n29964);
   U2536 : OAI21_X1 port map( A1 => n31516, A2 => n29761, B => n19599, ZN => 
                           n7001);
   U2592 : NAND2_X1 port map( A1 => n31889, A2 => n31888, ZN => n31887);
   U2601 : CLKBUF_X2 port map( I => n15153, Z => n31788);
   U2611 : AOI21_X1 port map( A1 => n12303, A2 => n12302, B => n9534, ZN => 
                           n18497);
   U2623 : NOR2_X1 port map( A1 => n982, A2 => n28236, ZN => n27991);
   U2629 : OAI21_X1 port map( A1 => n6181, A2 => n19318, B => n39689, ZN => 
                           n29646);
   U2645 : AND2_X1 port map( A1 => n37085, A2 => n25421, Z => n25612);
   U2647 : OR2_X1 port map( A1 => n28962, A2 => n19599, Z => n30391);
   U2669 : NAND2_X1 port map( A1 => n25540, A2 => n30317, ZN => n25474);
   U2674 : NOR2_X1 port map( A1 => n14418, A2 => n19202, ZN => n21536);
   U2675 : NOR2_X1 port map( A1 => n19202, A2 => n13285, ZN => n32372);
   U2701 : OR2_X1 port map( A1 => n5348, A2 => n19458, Z => n4169);
   U2705 : INV_X1 port map( I => n38584, ZN => n1502);
   U2721 : INV_X1 port map( I => n7335, ZN => n1628);
   U2757 : NAND2_X1 port map( A1 => n33307, A2 => n28021, ZN => n32963);
   U2760 : INV_X1 port map( I => n28676, ZN => n28671);
   U2771 : CLKBUF_X4 port map( I => n17876, Z => n14337);
   U2804 : NAND2_X1 port map( A1 => n2717, A2 => n15925, ZN => n30955);
   U2808 : NAND2_X1 port map( A1 => n11125, A2 => n30165, ZN => n30166);
   U2840 : NOR2_X1 port map( A1 => n30716, A2 => n28454, ZN => n32236);
   U2850 : NAND2_X1 port map( A1 => n31307, A2 => n29367, ZN => n29368);
   U2857 : NAND2_X1 port map( A1 => n29412, A2 => n17849, ZN => n15043);
   U2886 : NAND3_X1 port map( A1 => n15345, A2 => n15344, A3 => n39034, ZN => 
                           n15343);
   U2898 : NAND2_X1 port map( A1 => n982, A2 => n17314, ZN => n16851);
   U2902 : INV_X2 port map( I => n29660, ZN => n1390);
   U2907 : INV_X1 port map( I => n2296, ZN => n29593);
   U2921 : AOI21_X1 port map( A1 => n27292, A2 => n27221, B => n39546, ZN => 
                           n27018);
   U2926 : NOR2_X1 port map( A1 => n13981, A2 => n12943, ZN => n12942);
   U2934 : AOI21_X1 port map( A1 => n6036, A2 => n22156, B => n37199, ZN => 
                           n667);
   U2936 : OAI22_X1 port map( A1 => n22048, A2 => n16935, B1 => n36151, B2 => 
                           n6036, ZN => n14957);
   U2945 : NOR2_X1 port map( A1 => n1178, A2 => n17105, ZN => n7002);
   U2946 : AOI22_X1 port map( A1 => n29762, A2 => n29764, B1 => n29696, B2 => 
                           n17105, ZN => n7003);
   U2949 : NAND3_X1 port map( A1 => n30793, A2 => n30078, A3 => n30077, ZN => 
                           n30075);
   U3046 : OAI22_X1 port map( A1 => n19945, A2 => n17080, B1 => n17918, B2 => 
                           n17021, ZN => n22845);
   U3065 : NOR2_X1 port map( A1 => n9329, A2 => n38162, ZN => n9352);
   U3074 : NAND2_X1 port map( A1 => n32601, A2 => n23473, ZN => n32630);
   U3079 : CLKBUF_X1 port map( I => n37632, Z => n31160);
   U3080 : INV_X2 port map( I => n13799, ZN => n14400);
   U3089 : INV_X1 port map( I => n26713, ZN => n26849);
   U3092 : INV_X1 port map( I => n18711, ZN => n22245);
   U3100 : INV_X1 port map( I => n36798, ZN => n18801);
   U3129 : NAND2_X1 port map( A1 => n22204, A2 => n16265, ZN => n22206);
   U3130 : NAND2_X1 port map( A1 => n22204, A2 => n16265, ZN => n16262);
   U3151 : NOR2_X1 port map( A1 => n36340, A2 => n19901, ZN => n7154);
   U3155 : INV_X2 port map( I => n35443, ZN => n24792);
   U3160 : NAND2_X1 port map( A1 => n14400, A2 => n9733, ZN => n18140);
   U3161 : OAI21_X1 port map( A1 => n30144, A2 => n30132, B => n35234, ZN => 
                           n30133);
   U3168 : NOR2_X1 port map( A1 => n29975, A2 => n29980, ZN => n19041);
   U3176 : INV_X2 port map( I => n10907, ZN => n10906);
   U3199 : INV_X1 port map( I => n7485, ZN => n10494);
   U3200 : NOR2_X1 port map( A1 => n35367, A2 => n7485, ZN => n32363);
   U3203 : AOI21_X1 port map( A1 => n23572, A2 => n7485, B => n23571, ZN => 
                           n23367);
   U3220 : OAI21_X1 port map( A1 => n13805, A2 => n21684, B => n21431, ZN => 
                           n21416);
   U3229 : NAND2_X1 port map( A1 => n26702, A2 => n6190, ZN => n32261);
   U3244 : NAND2_X1 port map( A1 => n24759, A2 => n10054, ZN => n24762);
   U3248 : NAND2_X1 port map( A1 => n14404, A2 => n11891, ZN => n32059);
   U3272 : NAND2_X1 port map( A1 => n28237, A2 => n14462, ZN => n3779);
   U3282 : NAND2_X1 port map( A1 => n306, A2 => n28677, ZN => n28575);
   U3298 : OR2_X1 port map( A1 => n27919, A2 => n20860, Z => n27920);
   U3305 : NOR2_X1 port map( A1 => n17989, A2 => n35755, ZN => n7108);
   U3332 : INV_X1 port map( I => n3760, ZN => n24685);
   U3348 : NAND2_X1 port map( A1 => n25727, A2 => n16264, ZN => n25730);
   U3365 : NOR2_X1 port map( A1 => n4524, A2 => n37088, ZN => n23253);
   U3420 : NOR2_X1 port map( A1 => n18415, A2 => n18707, ZN => n5437);
   U3437 : AOI22_X1 port map( A1 => n12115, A2 => n1527, B1 => n31263, B2 => 
                           n38185, ZN => n13280);
   U3438 : INV_X1 port map( I => n32243, ZN => n13065);
   U3450 : AND2_X1 port map( A1 => n36369, A2 => n2350, Z => n30272);
   U3453 : INV_X2 port map( I => n8452, ZN => n9854);
   U3456 : OR2_X1 port map( A1 => n23531, A2 => n36539, Z => n30275);
   U3461 : NOR2_X2 port map( A1 => n23078, A2 => n23076, ZN => n32878);
   U3472 : INV_X2 port map( I => n38749, ZN => n32391);
   U3474 : XNOR2_X1 port map( A1 => n23773, A2 => n23772, ZN => n30280);
   U3493 : AND2_X1 port map( A1 => n27181, A2 => n27180, Z => n30288);
   U3533 : OR2_X1 port map( A1 => n29641, A2 => n29660, Z => n30295);
   U3539 : OR2_X2 port map( A1 => n2047, A2 => n17169, Z => n9651);
   U3561 : INV_X1 port map( I => n734, ZN => n2366);
   U3565 : NAND2_X1 port map( A1 => n28431, A2 => n28728, ZN => n31889);
   U3575 : NAND2_X1 port map( A1 => n8537, A2 => n19998, ZN => n19997);
   U3602 : AND2_X2 port map( A1 => n7666, A2 => n13794, Z => n14525);
   U3611 : NAND2_X1 port map( A1 => n36569, A2 => n11729, ZN => n27415);
   U3614 : NOR2_X1 port map( A1 => n6686, A2 => n11729, ZN => n11728);
   U3617 : NOR2_X1 port map( A1 => n9290, A2 => n38162, ZN => n9353);
   U3638 : NAND3_X1 port map( A1 => n28671, A2 => n36685, A3 => n1068, ZN => 
                           n28678);
   U3645 : NOR2_X1 port map( A1 => n3992, A2 => n2451, ZN => n30825);
   U3689 : INV_X1 port map( I => n10621, ZN => n10622);
   U3700 : INV_X2 port map( I => n4803, ZN => n27951);
   U3709 : NOR2_X1 port map( A1 => n11020, A2 => n27306, ZN => n12214);
   U3714 : NAND2_X1 port map( A1 => n9751, A2 => n19746, ZN => n18880);
   U3749 : INV_X1 port map( I => n26115, ZN => n25927);
   U3750 : NOR2_X1 port map( A1 => n2561, A2 => n26115, ZN => n2423);
   U3781 : AND2_X2 port map( A1 => n8628, A2 => n16174, Z => n17226);
   U3805 : NAND2_X1 port map( A1 => n3313, A2 => n35198, ZN => n27067);
   U3808 : NAND2_X1 port map( A1 => n8173, A2 => n5957, ZN => n14838);
   U3840 : AOI21_X1 port map( A1 => n12952, A2 => n1145, B => n35994, ZN => 
                           n4895);
   U3844 : NAND2_X1 port map( A1 => n257, A2 => n7810, ZN => n24669);
   U3895 : CLKBUF_X1 port map( I => n34175, Z => n33358);
   U3896 : BUF_X2 port map( I => n1418, Z => n32014);
   U3902 : NAND2_X1 port map( A1 => n274, A2 => n28278, ZN => n31116);
   U3905 : OR2_X1 port map( A1 => n33553, A2 => n10817, Z => n10827);
   U3910 : CLKBUF_X1 port map( I => n19982, Z => n30846);
   U3937 : NAND2_X1 port map( A1 => n1008, A2 => n36873, ZN => n32006);
   U3938 : NOR2_X1 port map( A1 => n32170, A2 => n19338, ZN => n32169);
   U3943 : OAI21_X1 port map( A1 => n21041, A2 => n25912, B => n32689, ZN => 
                           n16952);
   U3949 : INV_X2 port map( I => n5356, ZN => n1514);
   U3959 : NAND2_X1 port map( A1 => n826, A2 => n9893, ZN => n5860);
   U3960 : BUF_X2 port map( I => n15883, Z => n10882);
   U4004 : INV_X1 port map( I => n23199, ZN => n32872);
   U4013 : INV_X1 port map( I => n4846, ZN => n33075);
   U4016 : BUF_X2 port map( I => n22925, Z => n19535);
   U4028 : NAND2_X1 port map( A1 => n1683, A2 => n17781, ZN => n32803);
   U4043 : NOR2_X1 port map( A1 => n11149, A2 => n17307, ZN => n30826);
   U4046 : CLKBUF_X4 port map( I => n133, Z => n32640);
   U4047 : NAND2_X1 port map( A1 => n21751, A2 => n33876, ZN => n31365);
   U4059 : NAND2_X1 port map( A1 => n21676, A2 => n33053, ZN => n33052);
   U4062 : NOR2_X1 port map( A1 => n19641, A2 => n18143, ZN => n31034);
   U4066 : INV_X1 port map( I => n29964, ZN => n30324);
   U4067 : BUF_X2 port map( I => Key(58), Z => n19624);
   U4076 : NAND2_X1 port map( A1 => n3465, A2 => n31160, ZN => n31495);
   U4084 : INV_X2 port map( I => n29754, ZN => n30555);
   U4085 : NAND2_X1 port map( A1 => n31549, A2 => n30210, ZN => n33520);
   U4086 : NAND2_X1 port map( A1 => n20078, A2 => n30793, ZN => n20949);
   U4087 : NAND2_X1 port map( A1 => n20437, A2 => n29568, ZN => n30496);
   U4089 : AOI22_X1 port map( A1 => n4445, A2 => n5471, B1 => n19508, B2 => 
                           n2121, ZN => n32192);
   U4095 : NOR2_X1 port map( A1 => n34175, A2 => n19994, ZN => n5001);
   U4103 : OR2_X1 port map( A1 => n30160, A2 => n29185, Z => n3958);
   U4110 : NAND2_X1 port map( A1 => n29768, A2 => n29769, ZN => n5762);
   U4118 : CLKBUF_X2 port map( I => n29941, Z => n31629);
   U4128 : INV_X1 port map( I => n29249, ZN => n31173);
   U4149 : NOR2_X1 port map( A1 => n11028, A2 => n9141, ZN => n30714);
   U4158 : NOR2_X1 port map( A1 => n28749, A2 => n28748, ZN => n33123);
   U4166 : NOR2_X1 port map( A1 => n4228, A2 => n28356, ZN => n5926);
   U4172 : NAND2_X1 port map( A1 => n28443, A2 => n28444, ZN => n33472);
   U4176 : NOR2_X1 port map( A1 => n10305, A2 => n1418, ZN => n32314);
   U4179 : INV_X1 port map( I => n20621, ZN => n33555);
   U4198 : INV_X1 port map( I => n4232, ZN => n33353);
   U4200 : OR2_X1 port map( A1 => n11413, A2 => n20662, Z => n11613);
   U4205 : CLKBUF_X2 port map( I => n28689, Z => n31418);
   U4207 : NAND2_X1 port map( A1 => n31118, A2 => n31116, ZN => n13179);
   U4219 : NAND2_X1 port map( A1 => n35827, A2 => n30955, ZN => n5938);
   U4234 : NAND2_X1 port map( A1 => n13623, A2 => n1069, ZN => n31002);
   U4238 : INV_X1 port map( I => n31119, ZN => n31118);
   U4246 : INV_X1 port map( I => n28247, ZN => n31616);
   U4248 : NOR2_X1 port map( A1 => n28123, A2 => n10836, ZN => n32480);
   U4260 : CLKBUF_X2 port map( I => n28017, Z => n18150);
   U4284 : CLKBUF_X2 port map( I => n15287, Z => n31438);
   U4285 : CLKBUF_X4 port map( I => n27755, Z => n33587);
   U4295 : AND3_X2 port map( A1 => n17151, A2 => n15277, A3 => n15275, Z => 
                           n31602);
   U4304 : NAND2_X1 port map( A1 => n15748, A2 => n33017, ZN => n33016);
   U4314 : NAND2_X1 port map( A1 => n27113, A2 => n1481, ZN => n32756);
   U4324 : INV_X1 port map( I => n26889, ZN => n11432);
   U4340 : CLKBUF_X2 port map( I => n7632, Z => n32020);
   U4349 : BUF_X2 port map( I => n37245, Z => n5035);
   U4365 : NAND2_X1 port map( A1 => n32006, A2 => n32005, ZN => n9654);
   U4372 : NOR2_X1 port map( A1 => n33802, A2 => n10754, ZN => n21317);
   U4374 : NAND2_X1 port map( A1 => n17449, A2 => n8010, ZN => n17448);
   U4377 : INV_X1 port map( I => n26149, ZN => n33026);
   U4388 : AND2_X1 port map( A1 => n26918, A2 => n13393, Z => n30363);
   U4396 : BUF_X2 port map( I => n10029, Z => n15411);
   U4417 : CLKBUF_X2 port map( I => n755, Z => n30942);
   U4419 : CLKBUF_X2 port map( I => n18210, Z => n32009);
   U4447 : NAND2_X1 port map( A1 => n25905, A2 => n25904, ZN => n33630);
   U4459 : OR2_X1 port map( A1 => n26005, A2 => n25856, Z => n30468);
   U4462 : NOR2_X1 port map( A1 => n17791, A2 => n31133, ZN => n14680);
   U4464 : OR2_X1 port map( A1 => n38548, A2 => n34217, Z => n30425);
   U4481 : NOR2_X1 port map( A1 => n26019, A2 => n5859, ZN => n26022);
   U4495 : INV_X1 port map( I => n25108, ZN => n31416);
   U4498 : NAND2_X1 port map( A1 => n3278, A2 => n34087, ZN => n31963);
   U4503 : NAND2_X1 port map( A1 => n18145, A2 => n32355, ZN => n20007);
   U4505 : OAI21_X1 port map( A1 => n32291, A2 => n32279, B => n32278, ZN => 
                           n19501);
   U4507 : OR2_X1 port map( A1 => n21254, A2 => n33242, Z => n25724);
   U4513 : OR2_X1 port map( A1 => n31895, A2 => n31587, Z => n25444);
   U4520 : BUF_X2 port map( I => n25683, Z => n30633);
   U4531 : OR2_X1 port map( A1 => n10563, A2 => n25754, Z => n30399);
   U4550 : BUF_X2 port map( I => n10686, Z => n4467);
   U4555 : INV_X1 port map( I => n25239, ZN => n32613);
   U4562 : CLKBUF_X4 port map( I => n25292, Z => n30865);
   U4565 : BUF_X1 port map( I => n15186, Z => n33439);
   U4584 : CLKBUF_X2 port map( I => n19691, Z => n30733);
   U4586 : NAND2_X1 port map( A1 => n7830, A2 => n5607, ZN => n32368);
   U4587 : NAND2_X1 port map( A1 => n31361, A2 => n31360, ZN => n6081);
   U4595 : NAND2_X1 port map( A1 => n32641, A2 => n24800, ZN => n32644);
   U4596 : INV_X1 port map( I => n32641, ZN => n24656);
   U4620 : INV_X1 port map( I => n8173, ZN => n31713);
   U4622 : INV_X2 port map( I => n10931, ZN => n33409);
   U4624 : CLKBUF_X2 port map( I => n24673, Z => n33042);
   U4631 : NAND2_X1 port map( A1 => n14283, A2 => n1028, ZN => n16854);
   U4656 : OR2_X1 port map( A1 => n37732, A2 => n21125, Z => n30414);
   U4672 : INV_X1 port map( I => n7406, ZN => n30647);
   U4687 : INV_X1 port map( I => n24483, ZN => n33442);
   U4691 : NAND2_X1 port map( A1 => n24100, A2 => n37467, ZN => n24101);
   U4704 : CLKBUF_X2 port map( I => n19846, Z => n32973);
   U4709 : INV_X1 port map( I => n23724, ZN => n31178);
   U4711 : CLKBUF_X4 port map( I => n10638, Z => n32776);
   U4715 : INV_X1 port map( I => n23911, ZN => n1619);
   U4716 : INV_X1 port map( I => n2656, ZN => n31927);
   U4725 : OR2_X1 port map( A1 => n20817, A2 => n23516, Z => n23265);
   U4727 : NAND2_X1 port map( A1 => n2601, A2 => n17556, ZN => n2598);
   U4728 : NAND2_X1 port map( A1 => n33721, A2 => n23571, ZN => n33720);
   U4736 : AND2_X1 port map( A1 => n31586, A2 => n23456, Z => n30440);
   U4741 : NOR2_X1 port map( A1 => n20972, A2 => n23483, ZN => n20991);
   U4742 : AND2_X1 port map( A1 => n38535, A2 => n23516, Z => n14649);
   U4743 : CLKBUF_X2 port map( I => n33703, Z => n30499);
   U4751 : AND2_X1 port map( A1 => n18199, A2 => n31906, Z => n31949);
   U4752 : CLKBUF_X2 port map( I => n23607, Z => n32246);
   U4753 : BUF_X2 port map( I => n23568, Z => n31644);
   U4756 : OR2_X1 port map( A1 => n16197, A2 => n14429, Z => n30340);
   U4768 : NAND2_X1 port map( A1 => n21292, A2 => n33414, ZN => n22984);
   U4770 : OR2_X1 port map( A1 => n23022, A2 => n1655, Z => n7751);
   U4774 : CLKBUF_X2 port map( I => n4862, Z => n32270);
   U4778 : INV_X1 port map( I => n22932, ZN => n33554);
   U4783 : AND2_X1 port map( A1 => n19134, A2 => n23124, Z => n30360);
   U4788 : INV_X1 port map( I => n22990, ZN => n17930);
   U4792 : CLKBUF_X2 port map( I => n17464, Z => n31019);
   U4793 : CLKBUF_X2 port map( I => n782, Z => n31093);
   U4800 : CLKBUF_X2 port map( I => n4997, Z => n31838);
   U4806 : CLKBUF_X2 port map( I => n4291, Z => n32796);
   U4809 : BUF_X2 port map( I => n23129, Z => n19621);
   U4818 : INV_X1 port map( I => n10382, ZN => n33273);
   U4826 : NOR2_X1 port map( A1 => n16453, A2 => n16452, ZN => n30798);
   U4831 : INV_X2 port map( I => n17942, ZN => n30323);
   U4832 : INV_X1 port map( I => n33781, ZN => n33780);
   U4834 : AOI21_X1 port map( A1 => n31458, A2 => n17529, B => n22289, ZN => 
                           n2384);
   U4837 : NAND2_X1 port map( A1 => n22266, A2 => n33282, ZN => n21458);
   U4840 : NAND2_X1 port map( A1 => n22050, A2 => n4200, ZN => n30615);
   U4844 : INV_X2 port map( I => n22274, ZN => n1676);
   U4846 : CLKBUF_X2 port map( I => n22219, Z => n32408);
   U4854 : CLKBUF_X2 port map( I => n19518, Z => n33489);
   U4856 : NOR2_X1 port map( A1 => n21671, A2 => n6197, ZN => n31972);
   U4862 : NAND2_X1 port map( A1 => n33363, A2 => n21545, ZN => n33700);
   U4863 : NAND2_X1 port map( A1 => n21675, A2 => n19641, ZN => n33054);
   U4865 : OAI21_X1 port map( A1 => n18174, A2 => n36351, B => n31034, ZN => 
                           n6269);
   U4869 : CLKBUF_X2 port map( I => n21818, Z => n19388);
   U4873 : CLKBUF_X2 port map( I => n18027, Z => n32525);
   U4877 : CLKBUF_X2 port map( I => n21740, Z => n19287);
   U4878 : INV_X1 port map( I => n19932, ZN => n33515);
   U4885 : CLKBUF_X2 port map( I => n20887, Z => n32138);
   U4886 : CLKBUF_X2 port map( I => n21823, Z => n18143);
   U4887 : CLKBUF_X2 port map( I => n16333, Z => n33280);
   U4903 : NAND2_X1 port map( A1 => n15891, A2 => n21887, ZN => n33876);
   U4905 : NOR2_X1 port map( A1 => n14493, A2 => n19709, ZN => n19708);
   U4908 : NOR2_X1 port map( A1 => n19287, A2 => n38546, ZN => n21391);
   U4912 : INV_X1 port map( I => n21814, ZN => n21429);
   U4921 : NOR2_X1 port map( A1 => n17265, A2 => n19274, ZN => n12025);
   U4928 : NOR3_X1 port map( A1 => n21681, A2 => n19262, A3 => n19768, ZN => 
                           n18593);
   U4937 : NOR2_X1 port map( A1 => n10961, A2 => n21810, ZN => n36);
   U4945 : INV_X1 port map( I => n20368, ZN => n15053);
   U4955 : NAND2_X1 port map( A1 => n20996, A2 => n22047, ZN => n21971);
   U4960 : INV_X1 port map( I => n19655, ZN => n3001);
   U4998 : OR2_X1 port map( A1 => n22298, A2 => n19778, Z => n4280);
   U5015 : INV_X2 port map( I => n22067, ZN => n10242);
   U5018 : INV_X1 port map( I => n22569, ZN => n31012);
   U5028 : INV_X1 port map( I => n22463, ZN => n9187);
   U5045 : CLKBUF_X1 port map( I => n33990, Z => n32993);
   U5055 : NAND2_X1 port map( A1 => n17021, A2 => n22682, ZN => n18515);
   U5068 : INV_X1 port map( I => n23106, ZN => n31947);
   U5077 : CLKBUF_X2 port map( I => n22837, Z => n19788);
   U5078 : NOR2_X1 port map( A1 => n12163, A2 => n23188, ZN => n12699);
   U5082 : AOI21_X1 port map( A1 => n11307, A2 => n23107, B => n23111, ZN => 
                           n33414);
   U5104 : NAND2_X1 port map( A1 => n32042, A2 => n23060, ZN => n32041);
   U5109 : NAND2_X1 port map( A1 => n12083, A2 => n12028, ZN => n31611);
   U5188 : NOR2_X1 port map( A1 => n35689, A2 => n1642, ZN => n21250);
   U5190 : AND3_X1 port map( A1 => n1138, A2 => n10174, A3 => n23582, Z => 
                           n30445);
   U5235 : AND3_X1 port map( A1 => n17931, A2 => n23352, A3 => n13217, Z => 
                           n30456);
   U5249 : OAI22_X1 port map( A1 => n13150, A2 => n23578, B1 => n23506, B2 => 
                           n23580, ZN => n20947);
   U5250 : AND3_X1 port map( A1 => n15981, A2 => n17556, A3 => n1137, Z => n789
                           );
   U5256 : OAI21_X1 port map( A1 => n13602, A2 => n23390, B => n23452, ZN => 
                           n4543);
   U5262 : AND2_X1 port map( A1 => n18747, A2 => n23531, Z => n30457);
   U5268 : AOI22_X1 port map( A1 => n16716, A2 => n8692, B1 => n6176, B2 => 
                           n22513, ZN => n6139);
   U5276 : INV_X1 port map( I => n20777, ZN => n33573);
   U5284 : INV_X1 port map( I => n23841, ZN => n23788);
   U5286 : INV_X1 port map( I => n23812, ZN => n32097);
   U5304 : NAND2_X1 port map( A1 => n24114, A2 => n30320, ZN => n32742);
   U5310 : NOR2_X1 port map( A1 => n24371, A2 => n18466, ZN => n4784);
   U5316 : INV_X1 port map( I => n12975, ZN => n20339);
   U5353 : INV_X1 port map( I => n24863, ZN => n1566);
   U5376 : NAND2_X1 port map( A1 => n1909, A2 => n38626, ZN => n30635);
   U5384 : NOR2_X1 port map( A1 => n24692, A2 => n24576, ZN => n30642);
   U5390 : NAND2_X1 port map( A1 => n16196, A2 => n30699, ZN => n30698);
   U5404 : NAND2_X1 port map( A1 => n12633, A2 => n24759, ZN => n14267);
   U5410 : NOR2_X1 port map( A1 => n8127, A2 => n12124, ZN => n13638);
   U5419 : NAND2_X1 port map( A1 => n958, A2 => n30642, ZN => n6837);
   U5433 : INV_X1 port map( I => n33439, ZN => n30649);
   U5476 : CLKBUF_X2 port map( I => n21254, Z => n560);
   U5482 : INV_X2 port map( I => n13943, ZN => n18294);
   U5485 : NOR2_X1 port map( A1 => n31780, A2 => n19696, ZN => n11268);
   U5487 : NOR2_X1 port map( A1 => n25409, A2 => n25470, ZN => n25410);
   U5491 : NAND2_X1 port map( A1 => n4603, A2 => n31557, ZN => n32355);
   U5500 : NAND3_X1 port map( A1 => n9161, A2 => n17353, A3 => n32085, ZN => 
                           n11847);
   U5515 : INV_X2 port map( I => n35828, ZN => n26056);
   U5596 : INV_X1 port map( I => n19498, ZN => n33216);
   U5611 : INV_X1 port map( I => n21098, ZN => n17360);
   U5619 : INV_X1 port map( I => n33486, ZN => n26308);
   U5622 : OAI21_X1 port map( A1 => n31473, A2 => n1852, B => n18801, ZN => 
                           n1851);
   U5632 : NAND2_X1 port map( A1 => n26708, A2 => n36355, ZN => n32005);
   U5636 : NAND2_X1 port map( A1 => n26700, A2 => n14636, ZN => n17449);
   U5639 : NAND2_X1 port map( A1 => n26645, A2 => n34005, ZN => n19673);
   U5643 : NAND2_X1 port map( A1 => n14412, A2 => n17158, ZN => n32280);
   U5645 : INV_X1 port map( I => n26987, ZN => n13949);
   U5647 : AND3_X1 port map( A1 => n11864, A2 => n852, A3 => n26978, Z => 
                           n30356);
   U5660 : NAND2_X1 port map( A1 => n26831, A2 => n2882, ZN => n3091);
   U5712 : INV_X1 port map( I => n15433, ZN => n30811);
   U5720 : AOI21_X1 port map( A1 => n31518, A2 => n21248, B => n35265, ZN => 
                           n27422);
   U5731 : NAND2_X1 port map( A1 => n32169, A2 => n32167, ZN => n32166);
   U5737 : NOR2_X1 port map( A1 => n27372, A2 => n27269, ZN => n3469);
   U5797 : INV_X1 port map( I => n3604, ZN => n32021);
   U5840 : INV_X1 port map( I => n38213, ZN => n31304);
   U5851 : INV_X1 port map( I => n33584, ZN => n11947);
   U5863 : OAI21_X1 port map( A1 => n37418, A2 => n36197, B => n1076, ZN => 
                           n31119);
   U5875 : NAND2_X1 port map( A1 => n27877, A2 => n28001, ZN => n27878);
   U5904 : INV_X1 port map( I => n28739, ZN => n30581);
   U5909 : NAND2_X1 port map( A1 => n30370, A2 => n28138, ZN => n27966);
   U5932 : AOI21_X1 port map( A1 => n4284, A2 => n1196, B => n32575, ZN => 
                           n30741);
   U5947 : NAND2_X1 port map( A1 => n37204, A2 => n9668, ZN => n19668);
   U5983 : NAND2_X1 port map( A1 => n30741, A2 => n28682, ZN => n33610);
   U6016 : INV_X1 port map( I => n28888, ZN => n31398);
   U6019 : INV_X1 port map( I => n29099, ZN => n31692);
   U6025 : NAND2_X1 port map( A1 => n31699, A2 => n30380, ZN => n7030);
   U6068 : NAND2_X1 port map( A1 => n6443, A2 => n30242, ZN => n29009);
   U6070 : AOI21_X1 port map( A1 => n1175, A2 => n10590, B => n29210, ZN => 
                           n7899);
   U6082 : NAND2_X1 port map( A1 => n9508, A2 => n5570, ZN => n2861);
   U6083 : NOR2_X1 port map( A1 => n7141, A2 => n3986, ZN => n3170);
   U6086 : INV_X1 port map( I => n4169, ZN => n18413);
   U6090 : OAI21_X1 port map( A1 => n29699, A2 => n29701, B => n29700, ZN => 
                           n8345);
   U6093 : NAND2_X1 port map( A1 => n775, A2 => n34652, ZN => n33071);
   U6101 : CLKBUF_X1 port map( I => n29885, Z => n31598);
   U6103 : INV_X1 port map( I => n10848, ZN => n32706);
   U6106 : INV_X1 port map( I => n31532, ZN => n31211);
   U6109 : NOR2_X1 port map( A1 => n35176, A2 => n6252, ZN => n29540);
   U6114 : OAI21_X1 port map( A1 => n29732, A2 => n29755, B => n29756, ZN => 
                           n33766);
   U6134 : NAND2_X1 port map( A1 => n6622, A2 => n29968, ZN => n30709);
   U6166 : XNOR2_X1 port map( A1 => n36750, A2 => n19908, ZN => n30329);
   U6169 : XNOR2_X1 port map( A1 => n35241, A2 => n27576, ZN => n30333);
   U6173 : NOR2_X1 port map( A1 => n26687, A2 => n26978, ZN => n30336);
   U6179 : AND2_X1 port map( A1 => n18186, A2 => n17598, Z => n30339);
   U6191 : AND2_X1 port map( A1 => n18197, A2 => n18198, Z => n30342);
   U6194 : AND2_X1 port map( A1 => n31594, A2 => n23380, Z => n30345);
   U6207 : OR2_X1 port map( A1 => n22051, A2 => n35755, Z => n30354);
   U6215 : AND2_X1 port map( A1 => n26973, A2 => n26974, Z => n30355);
   U6234 : AND2_X1 port map( A1 => n1212, A2 => n15357, Z => n30369);
   U6236 : XNOR2_X1 port map( A1 => n9611, A2 => n1358, ZN => n30371);
   U6244 : AND2_X1 port map( A1 => n19415, A2 => n12235, Z => n30378);
   U6264 : NOR2_X1 port map( A1 => n37067, A2 => n9197, ZN => n30385);
   U6284 : OR2_X1 port map( A1 => n18417, A2 => n19287, Z => n30393);
   U6285 : AND2_X1 port map( A1 => n14880, A2 => n33925, Z => n30394);
   U6297 : XNOR2_X1 port map( A1 => n22665, A2 => n28968, ZN => n30402);
   U6302 : XNOR2_X1 port map( A1 => n23880, A2 => n30120, ZN => n30403);
   U6307 : XNOR2_X1 port map( A1 => n13569, A2 => n37109, ZN => n30404);
   U6309 : XNOR2_X1 port map( A1 => n29831, A2 => n25160, ZN => n30405);
   U6310 : XNOR2_X1 port map( A1 => n22651, A2 => n29298, ZN => n30406);
   U6322 : XNOR2_X1 port map( A1 => n11923, A2 => n28831, ZN => n30408);
   U6327 : XNOR2_X1 port map( A1 => n19221, A2 => n965, ZN => n30409);
   U6342 : AND3_X1 port map( A1 => n1472, A2 => n32926, A3 => n27447, Z => 
                           n30416);
   U6359 : OR2_X1 port map( A1 => n23570, A2 => n17556, Z => n30420);
   U6364 : INV_X1 port map( I => n21818, ZN => n21817);
   U6370 : XOR2_X1 port map( A1 => n20340, A2 => n20016, Z => n30423);
   U6375 : INV_X1 port map( I => n30629, ZN => n21039);
   U6380 : AND3_X2 port map( A1 => n19470, A2 => n34016, A3 => n20694, Z => 
                           n30427);
   U6384 : INV_X1 port map( I => n31473, ZN => n9320);
   U6386 : INV_X2 port map( I => n23542, ZN => n12154);
   U6393 : INV_X2 port map( I => n13442, ZN => n15209);
   U6400 : AND2_X1 port map( A1 => n28708, A2 => n28716, Z => n30431);
   U6403 : AND2_X1 port map( A1 => n16224, A2 => n29935, Z => n30432);
   U6410 : NAND2_X1 port map( A1 => n18077, A2 => n9781, ZN => n31358);
   U6431 : XOR2_X1 port map( A1 => n25279, A2 => n25281, Z => n30433);
   U6434 : INV_X1 port map( I => n30117, ZN => n30100);
   U6448 : XNOR2_X1 port map( A1 => n25189, A2 => n35379, ZN => n30435);
   U6450 : INV_X1 port map( I => n8745, ZN => n3109);
   U6486 : INV_X1 port map( I => n21571, ZN => n19271);
   U6496 : XNOR2_X1 port map( A1 => n22630, A2 => n36362, ZN => n30442);
   U6499 : INV_X2 port map( I => n5891, ZN => n12952);
   U6506 : XNOR2_X1 port map( A1 => n9982, A2 => n19902, ZN => n30444);
   U6508 : XNOR2_X1 port map( A1 => n23720, A2 => n23719, ZN => n30446);
   U6511 : XNOR2_X1 port map( A1 => n18582, A2 => n16893, ZN => n30447);
   U6512 : INV_X1 port map( I => n4291, ZN => n19698);
   U6514 : XNOR2_X1 port map( A1 => n15608, A2 => n15607, ZN => n30448);
   U6519 : XOR2_X1 port map( A1 => n22479, A2 => n22478, Z => n30450);
   U6521 : XOR2_X1 port map( A1 => n23739, A2 => n23738, Z => n30451);
   U6522 : XNOR2_X1 port map( A1 => n23915, A2 => n23914, ZN => n30452);
   U6523 : INV_X1 port map( I => n25683, ZN => n25649);
   U6527 : OR3_X1 port map( A1 => n4525, A2 => n20788, A3 => n37088, Z => 
                           n30453);
   U6534 : INV_X1 port map( I => n23610, ZN => n23292);
   U6541 : XNOR2_X1 port map( A1 => n23715, A2 => n14220, ZN => n30458);
   U6549 : XOR2_X1 port map( A1 => n19775, A2 => n6185, Z => n30459);
   U6552 : XOR2_X1 port map( A1 => n15679, A2 => n19875, Z => n30461);
   U6568 : INV_X1 port map( I => n25553, ZN => n18704);
   U6573 : XNOR2_X1 port map( A1 => n26520, A2 => n26551, ZN => n30469);
   U6584 : XNOR2_X1 port map( A1 => n8833, A2 => n30101, ZN => n30471);
   U6592 : XNOR2_X1 port map( A1 => n18399, A2 => n29238, ZN => n30473);
   U6599 : XNOR2_X1 port map( A1 => n35227, A2 => n15700, ZN => n30478);
   U6600 : XNOR2_X1 port map( A1 => n34332, A2 => n11994, ZN => n30479);
   U6602 : XNOR2_X1 port map( A1 => n1358, A2 => n9757, ZN => n30480);
   U6605 : XNOR2_X1 port map( A1 => n14566, A2 => n27578, ZN => n30481);
   U6606 : XNOR2_X1 port map( A1 => n27683, A2 => n19624, ZN => n30482);
   U6610 : XNOR2_X1 port map( A1 => n27683, A2 => n19583, ZN => n30483);
   U6632 : XNOR2_X1 port map( A1 => n38153, A2 => n31017, ZN => n30487);
   U6635 : XNOR2_X1 port map( A1 => n12430, A2 => n30094, ZN => n30488);
   U6636 : INV_X2 port map( I => n20010, ZN => n28149);
   U6641 : XNOR2_X1 port map( A1 => n29087, A2 => n28834, ZN => n30489);
   U6659 : OAI22_X1 port map( A1 => n14075, A2 => n29571, B1 => n31899, B2 => 
                           n30496, ZN => n14072);
   U6676 : NAND2_X2 port map( A1 => n5424, A2 => n19771, ZN => n28739);
   U6683 : XOR2_X1 port map( A1 => n31370, A2 => n30433, Z => n19582);
   U6686 : NAND2_X1 port map( A1 => n6181, A2 => n19318, ZN => n29648);
   U6720 : INV_X2 port map( I => n30503, ZN => n12682);
   U6734 : AND2_X1 port map( A1 => n2882, A2 => n7527, Z => n26726);
   U6737 : INV_X2 port map( I => n33966, ZN => n11898);
   U6739 : AOI21_X2 port map( A1 => n37138, A2 => n22890, B => n33361, ZN => 
                           n30701);
   U6789 : NAND3_X2 port map( A1 => n4484, A2 => n4483, A3 => n26547, ZN => 
                           n4034);
   U6791 : AOI22_X2 port map( A1 => n1746, A2 => n17530, B1 => n18303, B2 => 
                           n22042, ZN => n22182);
   U6797 : XNOR2_X1 port map( A1 => n3521, A2 => n30207, ZN => n31830);
   U6802 : NAND2_X1 port map( A1 => n3581, A2 => n7921, ZN => n31302);
   U6814 : XOR2_X1 port map( A1 => n30509, A2 => n12016, Z => n10162);
   U6815 : XOR2_X1 port map( A1 => n7582, A2 => n10163, Z => n30509);
   U6832 : XOR2_X1 port map( A1 => n23661, A2 => n31247, Z => n722);
   U6841 : XOR2_X1 port map( A1 => n30512, A2 => n19866, Z => Ciphertext(147));
   U6880 : OAI21_X2 port map( A1 => n13398, A2 => n19670, B => n30520, ZN => 
                           n19807);
   U6903 : NAND2_X2 port map( A1 => n24666, A2 => n24665, ZN => n2653);
   U6914 : NOR2_X1 port map( A1 => n12625, A2 => n16933, ZN => n33251);
   U6928 : INV_X2 port map( I => n23352, ZN => n31906);
   U6934 : XOR2_X1 port map( A1 => n27524, A2 => n27204, Z => n7061);
   U6951 : OR2_X1 port map( A1 => n27969, A2 => n876, Z => n18440);
   U6958 : XOR2_X1 port map( A1 => n29095, A2 => n17880, Z => n29835);
   U6961 : AOI21_X2 port map( A1 => n28059, A2 => n28548, B => n19354, ZN => 
                           n29095);
   U6964 : NOR2_X1 port map( A1 => n19891, A2 => n19605, ZN => n15569);
   U6967 : OAI21_X2 port map( A1 => n10626, A2 => n1588, B => n30529, ZN => 
                           n20326);
   U7015 : NAND2_X2 port map( A1 => n10254, A2 => n19750, ZN => n28052);
   U7024 : NAND2_X1 port map( A1 => n38198, A2 => n39140, ZN => n30611);
   U7025 : XOR2_X1 port map( A1 => n26253, A2 => n26026, Z => n26154);
   U7064 : OR2_X1 port map( A1 => n29346, A2 => n29241, Z => n13738);
   U7122 : XOR2_X1 port map( A1 => n18642, A2 => n30541, Z => n13410);
   U7124 : XOR2_X1 port map( A1 => n25028, A2 => n25029, Z => n30541);
   U7165 : XOR2_X1 port map( A1 => n27651, A2 => n27649, Z => n8281);
   U7216 : AOI21_X2 port map( A1 => n30547, A2 => n30546, B => n33795, ZN => 
                           n20491);
   U7240 : XOR2_X1 port map( A1 => n26227, A2 => n7602, Z => n26145);
   U7285 : AND2_X1 port map( A1 => n33147, A2 => n114, Z => n3784);
   U7326 : XOR2_X1 port map( A1 => n30551, A2 => n1980, Z => n1978);
   U7330 : XOR2_X1 port map( A1 => n31565, A2 => n10558, Z => n13383);
   U7338 : AND2_X1 port map( A1 => n23404, A2 => n2273, Z => n2274);
   U7343 : XOR2_X1 port map( A1 => n27769, A2 => n2582, Z => n20341);
   U7364 : NOR2_X2 port map( A1 => n33135, A2 => n13335, ZN => n31944);
   U7367 : OR2_X1 port map( A1 => n19941, A2 => n25581, Z => n32172);
   U7393 : NAND2_X1 port map( A1 => n4240, A2 => n32107, ZN => n30558);
   U7395 : AOI21_X2 port map( A1 => n18603, A2 => n20896, B => n19242, ZN => 
                           n15014);
   U7397 : XOR2_X1 port map( A1 => n20586, A2 => n19936, Z => n6768);
   U7403 : OAI21_X2 port map( A1 => n31825, A2 => n30457, B => n6611, ZN => 
                           n20586);
   U7425 : XOR2_X1 port map( A1 => n4476, A2 => n27847, Z => n30560);
   U7427 : XOR2_X1 port map( A1 => n30561, A2 => n14221, Z => n2372);
   U7428 : XOR2_X1 port map( A1 => n12741, A2 => n7489, Z => n30561);
   U7440 : XOR2_X1 port map( A1 => n30562, A2 => n13575, Z => n24741);
   U7462 : XOR2_X1 port map( A1 => n1504, A2 => n2150, Z => n8075);
   U7498 : NOR3_X2 port map( A1 => n19042, A2 => n31416, A3 => n18407, ZN => 
                           n25111);
   U7521 : NAND2_X2 port map( A1 => n10787, A2 => n10785, ZN => n33440);
   U7525 : NAND2_X1 port map( A1 => n24903, A2 => n37097, ZN => n24906);
   U7534 : NOR2_X2 port map( A1 => n2260, A2 => n2258, ZN => n27828);
   U7543 : OAI21_X2 port map( A1 => n5834, A2 => n9928, B => n4713, ZN => 
                           n11588);
   U7556 : XOR2_X1 port map( A1 => n7089, A2 => n29246, Z => n30578);
   U7561 : NAND2_X2 port map( A1 => n18257, A2 => n3096, ZN => n29789);
   U7562 : OAI22_X2 port map( A1 => n3245, A2 => n3246, B1 => n3247, B2 => 
                           n19508, ZN => n3096);
   U7614 : NOR2_X1 port map( A1 => n32046, A2 => n32566, ZN => n30582);
   U7616 : XOR2_X1 port map( A1 => n29021, A2 => n18931, Z => n29000);
   U7655 : AND2_X1 port map( A1 => n21822, A2 => n21857, Z => n21676);
   U7656 : INV_X2 port map( I => n19945, ZN => n33361);
   U7658 : NOR3_X1 port map( A1 => n1211, A2 => n31571, A3 => n30484, ZN => 
                           n31808);
   U7665 : NAND2_X2 port map( A1 => n17745, A2 => n17742, ZN => n24011);
   U7677 : NAND2_X2 port map( A1 => n24476, A2 => n24475, ZN => n24784);
   U7678 : XOR2_X1 port map( A1 => n3748, A2 => n3747, Z => n13124);
   U7682 : NAND3_X1 port map( A1 => n2861, A2 => n2859, A3 => n2860, ZN => 
                           n30664);
   U7691 : OR2_X1 port map( A1 => n840, A2 => n35828, Z => n5680);
   U7697 : NAND3_X1 port map( A1 => n25056, A2 => n37215, A3 => n25055, ZN => 
                           n33176);
   U7701 : NAND2_X2 port map( A1 => n32077, A2 => n6264, ZN => n28695);
   U7709 : XOR2_X1 port map( A1 => n30727, A2 => n29301, Z => n30602);
   U7711 : XOR2_X1 port map( A1 => n17567, A2 => n29054, Z => n29301);
   U7718 : INV_X2 port map( I => n28660, ZN => n28551);
   U7744 : AOI21_X2 port map( A1 => n28743, A2 => n28742, B => n30596, ZN => 
                           n12430);
   U7745 : OAI22_X2 port map( A1 => n30949, A2 => n31269, B1 => n28740, B2 => 
                           n28739, ZN => n30596);
   U7752 : AOI22_X2 port map( A1 => n13843, A2 => n24912, B1 => n30598, B2 => 
                           n36752, ZN => n25026);
   U7763 : AOI21_X2 port map( A1 => n8576, A2 => n17351, B => n8575, ZN => 
                           n12233);
   U7764 : AOI22_X2 port map( A1 => n30599, A2 => n22882, B1 => n22881, B2 => 
                           n14402, ZN => n23237);
   U7770 : XOR2_X1 port map( A1 => n31535, A2 => n1365, Z => n9164);
   U7785 : XOR2_X1 port map( A1 => n30602, A2 => n18405, Z => n4850);
   U7801 : NOR2_X2 port map( A1 => n9178, A2 => n9188, ZN => n18773);
   U7805 : NAND3_X1 port map( A1 => n6569, A2 => n24381, A3 => n6570, ZN => 
                           n30603);
   U7834 : XOR2_X1 port map( A1 => n3557, A2 => n31304, Z => n2159);
   U7842 : XOR2_X1 port map( A1 => n32646, A2 => n29522, Z => n33037);
   U7870 : OR2_X1 port map( A1 => n31164, A2 => n31661, Z => n11286);
   U7872 : XOR2_X1 port map( A1 => n35053, A2 => n14374, Z => n16190);
   U7877 : INV_X2 port map( I => n30607, ZN => n31809);
   U7914 : NAND2_X2 port map( A1 => n17214, A2 => n30608, ZN => n7063);
   U7921 : XOR2_X1 port map( A1 => n26523, A2 => n26526, Z => n30609);
   U7922 : XOR2_X1 port map( A1 => n38177, A2 => n16665, Z => n30610);
   U7932 : AOI22_X1 port map( A1 => n29577, A2 => n29565, B1 => n29566, B2 => 
                           n29563, ZN => n31197);
   U7933 : OR2_X1 port map( A1 => n13038, A2 => n39070, Z => n31235);
   U7949 : XOR2_X1 port map( A1 => n9947, A2 => n30482, Z => n30781);
   U7966 : NAND3_X1 port map( A1 => n29965, A2 => n1170, A3 => n29975, ZN => 
                           n29966);
   U7975 : NAND2_X1 port map( A1 => n31310, A2 => n1242, ZN => n25454);
   U7982 : OAI21_X1 port map( A1 => n29852, A2 => n11898, B => n11897, ZN => 
                           n30616);
   U8002 : XOR2_X1 port map( A1 => n2825, A2 => n20446, Z => n2824);
   U8006 : NAND2_X2 port map( A1 => n15023, A2 => n14513, ZN => n30894);
   U8021 : XOR2_X1 port map( A1 => n22774, A2 => n706, Z => n10237);
   U8024 : INV_X4 port map( I => n19828, ZN => n24770);
   U8032 : XOR2_X1 port map( A1 => n30619, A2 => n4616, Z => n1794);
   U8075 : OAI21_X2 port map( A1 => n13666, A2 => n8139, B => n13664, ZN => 
                           n25296);
   U8084 : XOR2_X1 port map( A1 => n27835, A2 => n27836, Z => n30626);
   U8093 : XNOR2_X1 port map( A1 => n27697, A2 => n12999, ZN => n32137);
   U8152 : OAI21_X2 port map( A1 => n30353, A2 => n30886, B => n29342, ZN => 
                           n15768);
   U8156 : INV_X1 port map( I => n792, ZN => n30632);
   U8164 : OAI22_X2 port map( A1 => n8446, A2 => n8445, B1 => n32548, B2 => 
                           n39828, ZN => n29885);
   U8176 : AND2_X1 port map( A1 => n27198, A2 => n13973, Z => n27031);
   U8226 : NAND2_X1 port map( A1 => n32670, A2 => n29375, ZN => n29315);
   U8230 : NAND3_X1 port map( A1 => n30643, A2 => n26643, A3 => n6606, ZN => 
                           n4484);
   U8235 : INV_X1 port map( I => n16466, ZN => n30988);
   U8245 : XOR2_X1 port map( A1 => n30645, A2 => n19624, Z => Ciphertext(59));
   U8259 : OAI21_X2 port map( A1 => n33422, A2 => n29973, B => n29971, ZN => 
                           n32570);
   U8272 : OR2_X1 port map( A1 => n23071, A2 => n14390, Z => n32626);
   U8278 : XOR2_X1 port map( A1 => n25009, A2 => n30649, Z => n30648);
   U8308 : NOR2_X2 port map( A1 => n30652, A2 => n16744, ZN => n17101);
   U8314 : XOR2_X1 port map( A1 => n28839, A2 => n28871, Z => n27944);
   U8334 : NAND2_X2 port map( A1 => n19661, A2 => n19360, ZN => n18682);
   U8359 : NAND2_X1 port map( A1 => n3218, A2 => n3217, ZN => n30653);
   U8401 : XOR2_X1 port map( A1 => n30657, A2 => n1365, Z => Ciphertext(73));
   U8424 : XOR2_X1 port map( A1 => n24933, A2 => n25197, Z => n25314);
   U8425 : NAND2_X2 port map( A1 => n17962, A2 => n17963, ZN => n24933);
   U8462 : XOR2_X1 port map( A1 => n19374, A2 => n14221, Z => n10156);
   U8478 : AOI21_X2 port map( A1 => n30360, A2 => n272, B => n30663, ZN => 
                           n3047);
   U8483 : NAND2_X2 port map( A1 => n30664, A2 => n2856, ZN => n2858);
   U8528 : OAI21_X2 port map( A1 => n27445, A2 => n27444, B => n30667, ZN => 
                           n27852);
   U8531 : XNOR2_X1 port map( A1 => n23658, A2 => n23910, ZN => n23740);
   U8539 : OAI21_X2 port map( A1 => n13776, A2 => n5427, B => n28269, ZN => 
                           n30668);
   U8572 : NOR2_X1 port map( A1 => n1470, A2 => n34279, ZN => n7922);
   U8577 : NAND2_X2 port map( A1 => n8506, A2 => n12510, ZN => n27288);
   U8611 : XOR2_X1 port map( A1 => n31782, A2 => n29022, Z => n32604);
   U8748 : NOR2_X1 port map( A1 => n29578, A2 => n28885, ZN => n30675);
   U8749 : AND2_X1 port map( A1 => n22407, A2 => n30676, Z => n18166);
   U8755 : NAND2_X2 port map( A1 => n4952, A2 => n30677, ZN => n15085);
   U8799 : OR2_X1 port map( A1 => n18519, A2 => n12162, Z => n7235);
   U8803 : XNOR2_X1 port map( A1 => n7247, A2 => n38184, ZN => n30819);
   U8820 : NAND2_X1 port map( A1 => n30454, A2 => n33734, ZN => n24216);
   U8840 : INV_X1 port map( I => n16657, ZN => n16655);
   U8842 : XOR2_X1 port map( A1 => n31778, A2 => n19213, Z => n31777);
   U8846 : XOR2_X1 port map( A1 => n29257, A2 => n29031, Z => n28041);
   U8858 : XOR2_X1 port map( A1 => n12399, A2 => n12402, Z => n12414);
   U8862 : XOR2_X1 port map( A1 => n32795, A2 => n30682, Z => n679);
   U8892 : AOI21_X2 port map( A1 => n20863, A2 => n31270, B => n30684, ZN => 
                           n4670);
   U8913 : XOR2_X1 port map( A1 => n8400, A2 => n30688, Z => n30687);
   U8918 : XOR2_X1 port map( A1 => n25156, A2 => n25043, Z => n8702);
   U8922 : NAND2_X2 port map( A1 => n3654, A2 => n3653, ZN => n25043);
   U8960 : INV_X2 port map( I => n18480, ZN => n2639);
   U8962 : INV_X1 port map( I => n32620, ZN => n17426);
   U8978 : NAND2_X2 port map( A1 => n19873, A2 => n34813, ZN => n7768);
   U8979 : INV_X2 port map( I => n30701, ZN => n71);
   U8981 : NOR2_X1 port map( A1 => n2868, A2 => n19888, ZN => n30702);
   U8989 : NAND2_X2 port map( A1 => n30704, A2 => n11847, ZN => n17212);
   U8991 : OAI21_X2 port map( A1 => n16317, A2 => n16316, B => n16315, ZN => 
                           n30704);
   U8992 : INV_X1 port map( I => n31984, ZN => n25362);
   U8995 : INV_X2 port map( I => n1666, ZN => n22459);
   U8998 : XOR2_X1 port map( A1 => n1666, A2 => n22503, Z => n20753);
   U8999 : NOR2_X2 port map( A1 => n30424, A2 => n30706, ZN => n1666);
   U9024 : XOR2_X1 port map( A1 => n27817, A2 => n18182, Z => n32698);
   U9038 : XOR2_X1 port map( A1 => n32621, A2 => n14872, Z => n29500);
   U9046 : NOR2_X2 port map( A1 => n20533, A2 => n30980, ZN => n28715);
   U9050 : OAI22_X1 port map( A1 => n5677, A2 => n19143, B1 => n30711, B2 => 
                           n30709, ZN => n17030);
   U9051 : NOR2_X1 port map( A1 => n1170, A2 => n6623, ZN => n30711);
   U9055 : NAND3_X1 port map( A1 => n5019, A2 => n13705, A3 => n5018, ZN => 
                           n19252);
   U9056 : NOR2_X1 port map( A1 => n35265, A2 => n27424, ZN => n30712);
   U9070 : NOR2_X1 port map( A1 => n19294, A2 => n24812, ZN => n24615);
   U9074 : XOR2_X1 port map( A1 => n22732, A2 => n4819, Z => n4896);
   U9079 : OR2_X2 port map( A1 => n9501, A2 => n9338, Z => n9441);
   U9080 : XOR2_X1 port map( A1 => n3028, A2 => n3029, Z => n9501);
   U9107 : XNOR2_X1 port map( A1 => n38181, A2 => n35249, ZN => n10183);
   U9125 : OAI21_X1 port map( A1 => n25469, A2 => n10004, B => n25606, ZN => 
                           n18249);
   U9143 : OR2_X1 port map( A1 => n39489, A2 => n22250, Z => n21090);
   U9178 : OR2_X1 port map( A1 => n3369, A2 => n26691, Z => n30726);
   U9198 : XOR2_X1 port map( A1 => n15271, A2 => n29300, Z => n30727);
   U9217 : XOR2_X1 port map( A1 => n30730, A2 => n30065, Z => Ciphertext(145));
   U9219 : NAND2_X1 port map( A1 => n33677, A2 => n33679, ZN => n31379);
   U9226 : INV_X1 port map( I => n21387, ZN => n21652);
   U9232 : NAND2_X1 port map( A1 => n30731, A2 => n18417, ZN => n14587);
   U9233 : XOR2_X1 port map( A1 => n21386, A2 => Key(125), Z => n21387);
   U9238 : AOI21_X2 port map( A1 => n30392, A2 => n18298, B => n17182, ZN => 
                           n2167);
   U9240 : NAND2_X2 port map( A1 => n16289, A2 => n16290, ZN => n22274);
   U9262 : INV_X2 port map( I => n2457, ZN => n20749);
   U9266 : NAND2_X2 port map( A1 => n27895, A2 => n28290, ZN => n2457);
   U9267 : NAND2_X1 port map( A1 => n231, A2 => n26268, ZN => n33142);
   U9270 : XOR2_X1 port map( A1 => n16334, A2 => n30734, Z => n19639);
   U9272 : XOR2_X1 port map( A1 => n19405, A2 => n29131, Z => n30734);
   U9284 : NAND2_X2 port map( A1 => n37245, A2 => n27211, ZN => n27259);
   U9289 : INV_X2 port map( I => n30736, ZN => n18721);
   U9299 : NAND2_X2 port map( A1 => n30738, A2 => n16137, ZN => n26009);
   U9305 : NAND2_X1 port map( A1 => n25740, A2 => n12624, ZN => n30738);
   U9317 : AND2_X1 port map( A1 => n1131, A2 => n12064, Z => n9460);
   U9329 : XOR2_X1 port map( A1 => n5434, A2 => n11321, Z => n32349);
   U9358 : NAND2_X1 port map( A1 => n29762, A2 => n29761, ZN => n30745);
   U9404 : XOR2_X1 port map( A1 => Plaintext(89), A2 => Key(89), Z => n21883);
   U9428 : NAND2_X2 port map( A1 => n11148, A2 => n15575, ZN => n25829);
   U9444 : INV_X4 port map( I => n33955, ZN => n1446);
   U9504 : OAI21_X2 port map( A1 => n1551, A2 => n15180, B => n16234, ZN => 
                           n25702);
   U9512 : XOR2_X1 port map( A1 => n25285, A2 => n13530, Z => n30756);
   U9559 : NAND2_X2 port map( A1 => n17118, A2 => n1151, ZN => n22178);
   U9563 : NAND2_X2 port map( A1 => n19907, A2 => n19906, ZN => n17118);
   U9577 : NOR2_X2 port map( A1 => n24833, A2 => n31385, ZN => n24755);
   U9618 : AOI21_X1 port map( A1 => n39065, A2 => n27069, B => n39417, ZN => 
                           n3581);
   U9657 : INV_X1 port map( I => n34166, ZN => n33842);
   U9675 : NAND2_X2 port map( A1 => n1951, A2 => n4416, ZN => n23931);
   U9691 : XOR2_X1 port map( A1 => n24064, A2 => n23658, Z => n23598);
   U9700 : XOR2_X1 port map( A1 => n4896, A2 => n15311, Z => n5540);
   U9704 : NAND2_X2 port map( A1 => n3025, A2 => n3024, ZN => n15311);
   U9736 : NAND2_X2 port map( A1 => n12523, A2 => n12524, ZN => n17455);
   U9746 : OAI21_X2 port map( A1 => n28377, A2 => n28665, B => n4002, ZN => 
                           n9112);
   U9747 : XOR2_X1 port map( A1 => n27759, A2 => n30771, Z => n33373);
   U9748 : XOR2_X1 port map( A1 => n27537, A2 => n37443, Z => n30771);
   U9769 : NAND2_X2 port map( A1 => n11083, A2 => n33662, ZN => n27273);
   U9777 : AOI21_X2 port map( A1 => n31130, A2 => n32725, B => n13159, ZN => 
                           n33662);
   U9818 : XOR2_X1 port map( A1 => n26167, A2 => n19798, Z => n30776);
   U9827 : XOR2_X1 port map( A1 => n39723, A2 => n19676, Z => n28958);
   U9840 : AOI21_X2 port map( A1 => n6065, A2 => n13033, B => n24963, ZN => 
                           n30778);
   U9856 : OAI21_X2 port map( A1 => n13469, A2 => n12475, B => n28165, ZN => 
                           n30780);
   U9895 : NAND2_X1 port map( A1 => n26706, A2 => n26705, ZN => n32347);
   U9900 : NAND2_X2 port map( A1 => n3319, A2 => n30945, ZN => n26115);
   U9904 : XOR2_X1 port map( A1 => n10483, A2 => n31983, Z => n4841);
   U9920 : NOR2_X1 port map( A1 => n31755, A2 => n36623, ZN => n30952);
   U9934 : OR2_X1 port map( A1 => n29236, A2 => n8728, Z => n14198);
   U9942 : AOI21_X1 port map( A1 => n23467, A2 => n3256, B => n18682, ZN => 
                           n31223);
   U9946 : OAI22_X1 port map( A1 => n5418, A2 => n28209, B1 => n28210, B2 => 
                           n28313, ZN => n30785);
   U9969 : OR2_X1 port map( A1 => n30764, A2 => n24719, Z => n6540);
   U9986 : BUF_X4 port map( I => n20326, Z => n6822);
   U9990 : OAI21_X2 port map( A1 => n3600, A2 => n3671, B => n3599, ZN => 
                           n20078);
   U9997 : NAND2_X2 port map( A1 => n30794, A2 => n10263, ZN => n12892);
   U10008 : NAND2_X2 port map( A1 => n17126, A2 => n13959, ZN => n30794);
   U10016 : NOR2_X2 port map( A1 => n30808, A2 => n5325, ZN => n12667);
   U10039 : NOR2_X2 port map( A1 => n30798, A2 => n16454, ZN => n17605);
   U10042 : NAND2_X2 port map( A1 => n21705, A2 => n21704, ZN => n22204);
   U10057 : INV_X4 port map( I => n30800, ZN => n22287);
   U10112 : XOR2_X1 port map( A1 => n27464, A2 => n30803, Z => n27029);
   U10116 : INV_X1 port map( I => n19816, ZN => n30803);
   U10125 : NAND2_X2 port map( A1 => n28539, A2 => n28495, ZN => n11129);
   U10145 : XOR2_X1 port map( A1 => n30806, A2 => n27816, Z => n31996);
   U10151 : NAND2_X2 port map( A1 => n26264, A2 => n15429, ZN => n15434);
   U10192 : NAND2_X1 port map( A1 => n19173, A2 => n29565, ZN => n31284);
   U10228 : OAI22_X2 port map( A1 => n15771, A2 => n15770, B1 => n18518, B2 => 
                           n22923, ZN => n23354);
   U10274 : OAI21_X2 port map( A1 => n32335, A2 => n2559, B => n29583, ZN => 
                           n2557);
   U10300 : XOR2_X1 port map( A1 => n26274, A2 => n26223, Z => n31627);
   U10301 : NOR2_X2 port map( A1 => n16344, A2 => n19048, ZN => n26274);
   U10363 : INV_X2 port map( I => n19746, ZN => n15443);
   U10398 : XOR2_X1 port map( A1 => n22625, A2 => n15610, Z => n15609);
   U10495 : AOI22_X1 port map( A1 => n29625, A2 => n29626, B1 => n29628, B2 => 
                           n29627, ZN => n31366);
   U10500 : NAND2_X2 port map( A1 => n1350, A2 => n39716, ZN => n11378);
   U10507 : INV_X2 port map( I => n32474, ZN => n19601);
   U10514 : NOR2_X2 port map( A1 => n24495, A2 => n24496, ZN => n24931);
   U10572 : XOR2_X1 port map( A1 => n5252, A2 => n5251, Z => n30831);
   U10613 : OAI21_X2 port map( A1 => n12062, A2 => n19452, B => n11860, ZN => 
                           n26070);
   U10639 : NOR2_X1 port map( A1 => n29498, A2 => n37614, ZN => n29302);
   U10646 : XOR2_X1 port map( A1 => n30318, A2 => n1260, Z => n30838);
   U10650 : OAI21_X2 port map( A1 => n27360, A2 => n32557, B => n30840, ZN => 
                           n2260);
   U10668 : XOR2_X1 port map( A1 => n23917, A2 => n23953, Z => n2120);
   U10680 : AOI21_X2 port map( A1 => n29633, A2 => n20816, B => n30847, ZN => 
                           n19297);
   U10682 : OAI22_X2 port map( A1 => n34089, A2 => n29632, B1 => n16385, B2 => 
                           n20982, ZN => n30847);
   U10683 : XOR2_X1 port map( A1 => n37699, A2 => n963, Z => n10163);
   U10759 : OR2_X1 port map( A1 => n23983, A2 => n16917, Z => n12646);
   U10761 : OAI21_X1 port map( A1 => n16502, A2 => n37640, B => n30854, ZN => 
                           n5123);
   U10767 : NAND2_X2 port map( A1 => n22227, A2 => n7357, ZN => n4316);
   U10801 : INV_X2 port map( I => n17984, ZN => n30859);
   U10803 : INV_X4 port map( I => n22238, ZN => n9546);
   U10869 : XOR2_X1 port map( A1 => n4592, A2 => n9518, Z => n16858);
   U10898 : OR2_X1 port map( A1 => n12302, A2 => n4803, Z => n11353);
   U10908 : INV_X1 port map( I => n36371, ZN => n1334);
   U10931 : XOR2_X1 port map( A1 => n16897, A2 => n18395, Z => n15450);
   U10932 : NOR2_X2 port map( A1 => n14935, A2 => n14934, ZN => n18395);
   U10943 : XOR2_X1 port map( A1 => n8775, A2 => n8773, Z => n28843);
   U10954 : OR2_X1 port map( A1 => n12331, A2 => n20449, Z => n22554);
   U10971 : NAND2_X1 port map( A1 => n15928, A2 => n21029, ZN => n32663);
   U10979 : NAND2_X2 port map( A1 => n20387, A2 => n20386, ZN => n22776);
   U10998 : AOI21_X2 port map( A1 => n29503, A2 => n29502, B => n37374, ZN => 
                           n29530);
   U11000 : NOR2_X1 port map( A1 => n29501, A2 => n18190, ZN => n30886);
   U11012 : XOR2_X1 port map( A1 => n1259, A2 => n19359, Z => n14639);
   U11024 : INV_X2 port map( I => n30890, ZN => n826);
   U11025 : XOR2_X1 port map( A1 => n13936, A2 => n13937, Z => n30890);
   U11028 : NAND2_X2 port map( A1 => n30323, A2 => n17943, ZN => n22772);
   U11031 : XOR2_X1 port map( A1 => n30891, A2 => n8631, Z => n8824);
   U11049 : XOR2_X1 port map( A1 => n33272, A2 => n30895, Z => n33244);
   U11050 : XOR2_X1 port map( A1 => n22321, A2 => n16531, Z => n30895);
   U11052 : BUF_X2 port map( I => n24192, Z => n30897);
   U11078 : NAND2_X1 port map( A1 => n27411, A2 => n6355, ZN => n10359);
   U11117 : INV_X2 port map( I => n30905, ZN => n10817);
   U11119 : XOR2_X1 port map( A1 => n10818, A2 => n10819, Z => n30905);
   U11123 : NOR2_X1 port map( A1 => n28396, A2 => n9848, ZN => n28298);
   U11162 : XOR2_X1 port map( A1 => n27675, A2 => n5697, Z => n30907);
   U11164 : OAI21_X1 port map( A1 => n1028, A2 => n24782, B => n24545, ZN => 
                           n16948);
   U11172 : NAND2_X2 port map( A1 => n30908, A2 => n4568, ZN => n11694);
   U11180 : INV_X1 port map( I => n13155, ZN => n26509);
   U11181 : XOR2_X1 port map( A1 => n19289, A2 => n13155, Z => n12860);
   U11190 : XOR2_X1 port map( A1 => n25144, A2 => n25299, Z => n30910);
   U11212 : NAND2_X2 port map( A1 => n30914, A2 => n24131, ZN => n24887);
   U11248 : XOR2_X1 port map( A1 => n1462, A2 => n17418, Z => n18633);
   U11315 : NAND2_X2 port map( A1 => n28573, A2 => n30928, ZN => n29837);
   U11318 : NAND3_X1 port map( A1 => n19321, A2 => n19322, A3 => n28666, ZN => 
                           n30928);
   U11334 : OR2_X1 port map( A1 => n691, A2 => n29548, Z => n15174);
   U11348 : AOI21_X2 port map( A1 => n27328, A2 => n27325, B => n32555, ZN => 
                           n30933);
   U11373 : XOR2_X1 port map( A1 => n13969, A2 => n12775, Z => n13332);
   U11376 : XOR2_X1 port map( A1 => n11358, A2 => n30938, Z => n9958);
   U11378 : XOR2_X1 port map( A1 => n17621, A2 => n30487, Z => n30938);
   U11383 : NAND2_X2 port map( A1 => n30939, A2 => n27324, ZN => n27735);
   U11397 : INV_X2 port map( I => n29441, ZN => n29435);
   U11398 : NAND2_X2 port map( A1 => n12261, A2 => n18494, ZN => n29441);
   U11435 : AOI21_X1 port map( A1 => n18518, A2 => n7537, B => n33361, ZN => 
                           n18516);
   U11444 : INV_X2 port map( I => n30946, ZN => n875);
   U11458 : NOR2_X1 port map( A1 => n1579, A2 => n19420, ZN => n30948);
   U11473 : XOR2_X1 port map( A1 => n28373, A2 => n28372, Z => n30956);
   U11520 : XOR2_X1 port map( A1 => n24013, A2 => n17725, Z => n16109);
   U11533 : XOR2_X1 port map( A1 => n23755, A2 => n18301, Z => n23736);
   U11535 : OAI22_X2 port map( A1 => n10612, A2 => n13560, B1 => n10614, B2 => 
                           n10613, ZN => n18301);
   U11550 : NAND2_X2 port map( A1 => n30962, A2 => n27925, ZN => n5418);
   U11555 : XOR2_X1 port map( A1 => n24068, A2 => n5842, Z => n30963);
   U11583 : NAND2_X2 port map( A1 => n30965, A2 => n28477, ZN => n29093);
   U11584 : OAI21_X2 port map( A1 => n9674, A2 => n31088, B => n9673, ZN => 
                           n30965);
   U11594 : OAI21_X2 port map( A1 => n31452, A2 => n24283, B => n24284, ZN => 
                           n24120);
   U11601 : NOR2_X1 port map( A1 => n38367, A2 => n32472, ZN => n17867);
   U11622 : XOR2_X1 port map( A1 => n23813, A2 => n34851, Z => n30976);
   U11630 : AOI22_X2 port map( A1 => n1673, A2 => n30306, B1 => n12077, B2 => 
                           n22126, ZN => n32667);
   U11631 : XOR2_X1 port map( A1 => n27731, A2 => n19943, Z => n27079);
   U11639 : XOR2_X1 port map( A1 => n30971, A2 => n30169, Z => Ciphertext(174))
                           ;
   U11647 : AOI21_X2 port map( A1 => n20947, A2 => n14855, B => n20946, ZN => 
                           n23762);
   U11650 : XOR2_X1 port map( A1 => n30972, A2 => n27518, Z => n7729);
   U11651 : XOR2_X1 port map( A1 => n27640, A2 => n30973, Z => n30972);
   U11656 : INV_X1 port map( I => n29718, ZN => n30973);
   U11657 : NOR2_X2 port map( A1 => n8385, A2 => n14261, ZN => n10508);
   U11662 : XNOR2_X1 port map( A1 => n5688, A2 => n34513, ZN => n33486);
   U11663 : XOR2_X1 port map( A1 => n26369, A2 => n26371, Z => n19021);
   U11672 : NOR2_X1 port map( A1 => n21445, A2 => n16496, ZN => n21671);
   U11686 : OR2_X1 port map( A1 => n7424, A2 => n14949, Z => n27321);
   U11699 : NAND2_X1 port map( A1 => n1382, A2 => n35175, ZN => n2490);
   U11730 : OR2_X2 port map( A1 => n17767, A2 => n7281, Z => n6777);
   U11748 : INV_X2 port map( I => n30982, ZN => n33949);
   U11763 : NOR2_X1 port map( A1 => n23435, A2 => n34494, ZN => n31798);
   U11785 : OR2_X1 port map( A1 => n30986, A2 => n9369, Z => n9415);
   U11796 : XOR2_X1 port map( A1 => n30990, A2 => n8975, Z => n13595);
   U11798 : XOR2_X1 port map( A1 => n27727, A2 => n8974, Z => n30990);
   U11814 : OAI21_X2 port map( A1 => n10467, A2 => n10468, B => n9683, ZN => 
                           n31181);
   U11819 : XOR2_X1 port map( A1 => n26530, A2 => n26559, Z => n32386);
   U11827 : AND3_X1 port map( A1 => n1755, A2 => n4083, A3 => n20405, Z => 
                           n30197);
   U11842 : XOR2_X1 port map( A1 => n34091, A2 => n8283, Z => n30994);
   U11845 : NAND2_X2 port map( A1 => n10261, A2 => n12892, ZN => n22194);
   U11854 : NAND2_X2 port map( A1 => n16024, A2 => n13743, ZN => n25860);
   U11876 : OR2_X1 port map( A1 => n7424, A2 => n31006, Z => n20725);
   U11887 : XOR2_X1 port map( A1 => n10860, A2 => n10858, Z => n17169);
   U11891 : NAND2_X1 port map( A1 => n31002, A2 => n31001, ZN => n13621);
   U11902 : NOR2_X1 port map( A1 => n20655, A2 => n24433, ZN => n20654);
   U11903 : NOR2_X1 port map( A1 => n24444, A2 => n24443, ZN => n31003);
   U11908 : NAND2_X1 port map( A1 => n20873, A2 => n22813, ZN => n23075);
   U11909 : NOR2_X1 port map( A1 => n12790, A2 => n17887, ZN => n22967);
   U11918 : AOI22_X2 port map( A1 => n31475, A2 => n33864, B1 => n3884, B2 => 
                           n8757, ZN => n32506);
   U11953 : OR3_X1 port map( A1 => n9790, A2 => n35272, A3 => n16260, Z => 
                           n31997);
   U11985 : INV_X2 port map( I => n14949, ZN => n31006);
   U12011 : NAND2_X2 port map( A1 => n20663, A2 => n14232, ZN => n11875);
   U12020 : AOI22_X2 port map( A1 => n18645, A2 => n21469, B1 => n2628, B2 => 
                           n12314, ZN => n2736);
   U12031 : OAI21_X2 port map( A1 => n23571, A2 => n23577, B => n12153, ZN => 
                           n23540);
   U12088 : NAND2_X1 port map( A1 => n33905, A2 => n33904, ZN => n32057);
   U12090 : XOR2_X1 port map( A1 => n19428, A2 => n31016, Z => n32621);
   U12104 : XOR2_X1 port map( A1 => n29303, A2 => n31017, Z => n31016);
   U12110 : INV_X1 port map( I => n19534, ZN => n31017);
   U12123 : AOI21_X2 port map( A1 => n14103, A2 => n11875, B => n11876, ZN => 
                           n7428);
   U12152 : XOR2_X1 port map( A1 => n15450, A2 => n21259, Z => n13936);
   U12159 : XOR2_X1 port map( A1 => n19072, A2 => n3589, Z => n437);
   U12166 : XOR2_X1 port map( A1 => n17486, A2 => n17487, Z => n7371);
   U12172 : NAND3_X1 port map( A1 => n4864, A2 => n4865, A3 => n1047, ZN => 
                           n6032);
   U12185 : NAND2_X2 port map( A1 => n28557, A2 => n28558, ZN => n9930);
   U12199 : OAI21_X1 port map( A1 => n24784, A2 => n37411, B => n31023, ZN => 
                           n15878);
   U12222 : XOR2_X1 port map( A1 => n32646, A2 => n19800, Z => n22532);
   U12253 : AND2_X1 port map( A1 => n29361, A2 => n13804, Z => n32767);
   U12263 : AOI22_X1 port map( A1 => n21618, A2 => n3907, B1 => n38673, B2 => 
                           n38448, ZN => n3909);
   U12277 : XOR2_X1 port map( A1 => n31031, A2 => n33434, Z => n20284);
   U12329 : XOR2_X1 port map( A1 => n25077, A2 => n25078, Z => n33044);
   U12331 : NAND2_X1 port map( A1 => n21282, A2 => n21283, ZN => n31726);
   U12393 : INV_X2 port map( I => n28025, ZN => n27948);
   U12406 : OR2_X1 port map( A1 => n19863, A2 => n19153, Z => n12463);
   U12439 : XOR2_X1 port map( A1 => n447, A2 => n31046, Z => n3852);
   U12451 : XOR2_X1 port map( A1 => n3855, A2 => n29029, Z => n31046);
   U12454 : OR2_X1 port map( A1 => n31278, A2 => n13144, Z => n24114);
   U12462 : INV_X2 port map( I => n31507, ZN => n21401);
   U12464 : NAND3_X2 port map( A1 => n18341, A2 => n19038, A3 => n19039, ZN => 
                           n28434);
   U12470 : XOR2_X1 port map( A1 => n3645, A2 => n31047, Z => n25669);
   U12489 : XOR2_X1 port map( A1 => n25202, A2 => n30459, Z => n31047);
   U12494 : XOR2_X1 port map( A1 => n26155, A2 => n25947, Z => n5965);
   U12510 : NOR2_X2 port map( A1 => n30131, A2 => n18588, ZN => n12350);
   U12535 : XOR2_X1 port map( A1 => n8132, A2 => n14102, Z => n14101);
   U12559 : NOR2_X2 port map( A1 => n10420, A2 => n37056, ZN => n28418);
   U12563 : AOI21_X1 port map( A1 => n28546, A2 => n3944, B => n36623, ZN => 
                           n31699);
   U12596 : XNOR2_X1 port map( A1 => n15671, A2 => n11253, ZN => n31352);
   U12624 : NAND3_X1 port map( A1 => n29763, A2 => n29764, A3 => n19599, ZN => 
                           n31059);
   U12630 : INV_X4 port map( I => n2242, ZN => n9105);
   U12633 : AOI21_X2 port map( A1 => n6332, A2 => n19147, B => n2243, ZN => 
                           n2242);
   U12638 : NAND3_X1 port map( A1 => n15737, A2 => n35224, A3 => n15224, ZN => 
                           n28466);
   U12643 : XOR2_X1 port map( A1 => n269, A2 => n31062, Z => n31061);
   U12645 : INV_X1 port map( I => n19843, ZN => n31062);
   U12682 : XOR2_X1 port map( A1 => n24959, A2 => n30682, Z => n1819);
   U12696 : XOR2_X1 port map( A1 => n31070, A2 => n31585, Z => n27473);
   U12710 : NOR2_X1 port map( A1 => n32318, A2 => n17685, ZN => n22253);
   U12730 : NAND2_X1 port map( A1 => n4889, A2 => n5938, ZN => n3193);
   U12742 : AOI21_X2 port map( A1 => n11056, A2 => n29422, B => n907, ZN => 
                           n29354);
   U12747 : NAND2_X2 port map( A1 => n18550, A2 => n18552, ZN => n18148);
   U12752 : XOR2_X1 port map( A1 => n8110, A2 => n11935, Z => n26225);
   U12754 : NOR2_X1 port map( A1 => n21747, A2 => n38546, ZN => n32808);
   U12775 : NAND3_X1 port map( A1 => n29384, A2 => n10422, A3 => n11084, ZN => 
                           n6262);
   U12786 : XOR2_X1 port map( A1 => n11074, A2 => n11076, Z => n13417);
   U12819 : AOI21_X2 port map( A1 => n23331, A2 => n32226, B => n20118, ZN => 
                           n24070);
   U12821 : AOI21_X2 port map( A1 => n20438, A2 => n4601, B => n5245, ZN => 
                           n25247);
   U12825 : INV_X2 port map( I => n31078, ZN => n12064);
   U12832 : OAI21_X2 port map( A1 => n16224, A2 => n29935, B => n8593, ZN => 
                           n8592);
   U12833 : INV_X2 port map( I => n18910, ZN => n18972);
   U12864 : NAND2_X2 port map( A1 => n31082, A2 => n25628, ZN => n11033);
   U12881 : NAND2_X2 port map( A1 => n35618, A2 => n8275, ZN => n5527);
   U12892 : NOR2_X2 port map( A1 => n3685, A2 => n38886, ZN => n12665);
   U12910 : XOR2_X1 port map( A1 => n31086, A2 => n29934, Z => Ciphertext(131))
                           ;
   U12930 : AOI22_X1 port map( A1 => n29931, A2 => n9591, B1 => n29933, B2 => 
                           n29932, ZN => n31086);
   U12944 : NAND2_X2 port map( A1 => n24243, A2 => n17591, ZN => n7520);
   U12964 : OAI22_X2 port map( A1 => n13762, A2 => n34064, B1 => n29287, B2 => 
                           n29348, ZN => n12371);
   U12972 : XOR2_X1 port map( A1 => n31089, A2 => n7382, Z => n10816);
   U13005 : NAND2_X2 port map( A1 => n14017, A2 => n31090, ZN => n23619);
   U13009 : OR2_X1 port map( A1 => n23186, A2 => n11197, Z => n31090);
   U13011 : NAND2_X1 port map( A1 => n20835, A2 => n23390, ZN => n31091);
   U13013 : BUF_X2 port map( I => n14349, Z => n31092);
   U13017 : XOR2_X1 port map( A1 => n7358, A2 => n22614, Z => n4279);
   U13037 : NAND2_X2 port map( A1 => n31094, A2 => n16543, ZN => n33707);
   U13042 : AOI21_X2 port map( A1 => n28699, A2 => n16494, B => n13718, ZN => 
                           n126);
   U13059 : NAND2_X2 port map( A1 => n2725, A2 => n32918, ZN => n20276);
   U13064 : XOR2_X1 port map( A1 => n22748, A2 => n7200, Z => n7199);
   U13079 : XOR2_X1 port map( A1 => n13871, A2 => n14104, Z => n24369);
   U13086 : XOR2_X1 port map( A1 => n2135, A2 => n2136, Z => n2134);
   U13131 : NAND2_X2 port map( A1 => n22043, A2 => n22044, ZN => n22634);
   U13134 : NOR2_X2 port map( A1 => n9667, A2 => n26008, ZN => n33892);
   U13151 : NOR2_X2 port map( A1 => n32183, A2 => n31102, ZN => n33286);
   U13156 : AND2_X2 port map( A1 => n32838, A2 => n16832, Z => n13884);
   U13157 : XOR2_X1 port map( A1 => n3240, A2 => n31103, Z => n11643);
   U13158 : XOR2_X1 port map( A1 => n22530, A2 => n18969, Z => n31103);
   U13163 : XOR2_X1 port map( A1 => n31628, A2 => n25271, Z => n21154);
   U13172 : INV_X4 port map( I => n12064, ZN => n15049);
   U13189 : XOR2_X1 port map( A1 => n6388, A2 => n31108, Z => n10810);
   U13196 : XOR2_X1 port map( A1 => n20695, A2 => n6387, Z => n31108);
   U13220 : OR2_X1 port map( A1 => n27009, A2 => n12156, Z => n31110);
   U13224 : NAND2_X2 port map( A1 => n4988, A2 => n4989, ZN => n33293);
   U13225 : NAND2_X2 port map( A1 => n31115, A2 => n31114, ZN => n18987);
   U13236 : XOR2_X1 port map( A1 => n25226, A2 => n14385, Z => n25289);
   U13245 : OR2_X1 port map( A1 => n12408, A2 => n16547, Z => n32430);
   U13247 : INV_X2 port map( I => n31121, ZN => n28152);
   U13255 : NOR3_X2 port map( A1 => n4578, A2 => n31123, A3 => n31122, ZN => 
                           n24961);
   U13259 : NAND2_X2 port map( A1 => n31124, A2 => n33042, ZN => n3214);
   U13265 : AOI22_X1 port map( A1 => n29665, A2 => n30295, B1 => n29648, B2 => 
                           n29654, ZN => n32288);
   U13279 : INV_X2 port map( I => n9113, ZN => n9114);
   U13302 : XOR2_X1 port map( A1 => n31129, A2 => n33466, Z => n12315);
   U13306 : XOR2_X1 port map( A1 => n19118, A2 => n22602, Z => n31129);
   U13309 : XOR2_X1 port map( A1 => n20668, A2 => n22532, Z => n11750);
   U13319 : XOR2_X1 port map( A1 => n9121, A2 => n9123, Z => n9458);
   U13335 : XOR2_X1 port map( A1 => n15164, A2 => n27719, Z => n17138);
   U13378 : NAND2_X2 port map( A1 => n24120, A2 => n32891, ZN => n23766);
   U13382 : XOR2_X1 port map( A1 => n26420, A2 => n3710, Z => n33751);
   U13406 : XOR2_X1 port map( A1 => n31138, A2 => n27229, Z => n342);
   U13410 : XOR2_X1 port map( A1 => n24994, A2 => n31139, Z => n14350);
   U13415 : INV_X2 port map( I => n36992, ZN => n4880);
   U13430 : INV_X4 port map( I => n23523, ZN => n23522);
   U13432 : XOR2_X1 port map( A1 => n4305, A2 => n1819, Z => n33188);
   U13435 : XOR2_X1 port map( A1 => n31149, A2 => n1361, Z => Ciphertext(83));
   U13445 : AOI22_X1 port map( A1 => n29665, A2 => n29664, B1 => n29663, B2 => 
                           n1390, ZN => n31149);
   U13454 : NAND2_X2 port map( A1 => n992, A2 => n32557, ZN => n31150);
   U13458 : NAND2_X2 port map( A1 => n13228, A2 => n13227, ZN => n24250);
   U13491 : XOR2_X1 port map( A1 => n16587, A2 => n31152, Z => n6834);
   U13493 : XOR2_X1 port map( A1 => n29071, A2 => n19814, Z => n31152);
   U13500 : XOR2_X1 port map( A1 => n2864, A2 => n39172, Z => n31154);
   U13562 : NAND2_X1 port map( A1 => n35828, A2 => n9743, ZN => n5681);
   U13578 : XOR2_X1 port map( A1 => n21197, A2 => n22614, Z => n5703);
   U13581 : XOR2_X1 port map( A1 => n22711, A2 => n22475, Z => n22614);
   U13646 : XOR2_X1 port map( A1 => n29111, A2 => n13933, Z => n31162);
   U13704 : XOR2_X1 port map( A1 => n27714, A2 => n7345, Z => n4783);
   U13790 : XOR2_X1 port map( A1 => n35529, A2 => n31173, Z => n20006);
   U13803 : NAND2_X2 port map( A1 => n18281, A2 => n7905, ZN => n28516);
   U13810 : AND2_X1 port map( A1 => n39504, A2 => n8735, Z => n31177);
   U13819 : XOR2_X1 port map( A1 => n9122, A2 => n31178, Z => n8300);
   U13828 : OR2_X1 port map( A1 => n15854, A2 => n10959, Z => n29892);
   U13836 : XOR2_X1 port map( A1 => n2161, A2 => n2162, Z => n29865);
   U13841 : XOR2_X1 port map( A1 => n12850, A2 => n33165, Z => n11562);
   U13876 : NAND2_X2 port map( A1 => n1102, A2 => n25966, ZN => n19340);
   U13902 : OAI22_X2 port map( A1 => n20287, A2 => n29634, B1 => n20286, B2 => 
                           n20289, ZN => n29660);
   U13982 : XOR2_X1 port map( A1 => n31191, A2 => n27695, Z => n27696);
   U13983 : XOR2_X1 port map( A1 => n13569, A2 => n34963, Z => n31191);
   U14073 : NAND2_X1 port map( A1 => n16778, A2 => n9405, ZN => n9404);
   U14076 : NAND2_X1 port map( A1 => n16778, A2 => n13880, ZN => n31194);
   U14094 : INV_X2 port map( I => n31196, ZN => n2799);
   U14096 : XOR2_X1 port map( A1 => n2800, A2 => n4129, Z => n31196);
   U14102 : XOR2_X1 port map( A1 => n31197, A2 => n33661, Z => Ciphertext(67));
   U14104 : XOR2_X1 port map( A1 => n27777, A2 => n27707, Z => n27204);
   U14124 : NOR3_X1 port map( A1 => n30859, A2 => n37104, A3 => n33561, ZN => 
                           n5481);
   U14139 : INV_X2 port map( I => n31204, ZN => n27790);
   U14141 : XOR2_X1 port map( A1 => n22447, A2 => n700, Z => n7932);
   U14149 : INV_X2 port map( I => n31207, ZN => n10383);
   U14156 : NAND2_X2 port map( A1 => n31132, A2 => n24416, ZN => n17496);
   U14173 : AOI21_X1 port map( A1 => n31212, A2 => n31211, B => n29338, ZN => 
                           n3285);
   U14174 : NAND2_X1 port map( A1 => n29339, A2 => n29336, ZN => n31212);
   U14175 : INV_X4 port map( I => n10383, ZN => n33745);
   U14196 : XOR2_X1 port map( A1 => n11374, A2 => n746, Z => n31215);
   U14211 : NAND2_X2 port map( A1 => n32813, A2 => n2363, ZN => n27408);
   U14217 : OAI21_X1 port map( A1 => n19972, A2 => n1234, B => n31220, ZN => 
                           n2364);
   U14246 : XOR2_X1 port map( A1 => n6470, A2 => n31230, Z => n9516);
   U14247 : XOR2_X1 port map( A1 => n27555, A2 => n18709, Z => n31230);
   U14248 : OR2_X1 port map( A1 => n29810, A2 => n13192, Z => n31231);
   U14265 : XOR2_X1 port map( A1 => n8908, A2 => n38225, Z => n31233);
   U14273 : AOI22_X2 port map( A1 => n13259, A2 => n13019, B1 => n25204, B2 => 
                           n24944, ZN => n25299);
   U14278 : NAND2_X2 port map( A1 => n31236, A2 => n5299, ZN => n30178);
   U14305 : AND2_X1 port map( A1 => n39814, A2 => n17509, Z => n2975);
   U14318 : INV_X1 port map( I => n23768, ZN => n31245);
   U14319 : NOR2_X1 port map( A1 => n31245, A2 => n5897, ZN => n31360);
   U14320 : XOR2_X1 port map( A1 => n15930, A2 => n25275, Z => n25007);
   U14330 : NOR2_X1 port map( A1 => n24283, A2 => n24284, ZN => n20732);
   U14338 : BUF_X2 port map( I => n23775, Z => n31247);
   U14344 : XOR2_X1 port map( A1 => n37812, A2 => n31249, Z => n31248);
   U14347 : XOR2_X1 port map( A1 => n17245, A2 => n31689, Z => n31688);
   U14353 : INV_X2 port map( I => n31250, ZN => n733);
   U14354 : XOR2_X1 port map( A1 => n3579, A2 => n3577, Z => n31250);
   U14357 : AND2_X1 port map( A1 => n32146, A2 => n28620, Z => n13404);
   U14361 : AOI21_X2 port map( A1 => n25433, A2 => n36086, B => n18565, ZN => 
                           n26106);
   U14367 : AOI22_X2 port map( A1 => n31252, A2 => n14371, B1 => n4128, B2 => 
                           n32899, ZN => n20728);
   U14369 : INV_X2 port map( I => n14422, ZN => n1055);
   U14383 : NAND2_X1 port map( A1 => n31258, A2 => n19098, ZN => n10031);
   U14391 : NAND2_X2 port map( A1 => n33317, A2 => n20158, ZN => n24713);
   U14406 : AND2_X1 port map( A1 => n21671, A2 => n21672, Z => n6046);
   U14407 : AND2_X1 port map( A1 => n38886, A2 => n17509, Z => n2971);
   U14422 : NAND2_X1 port map( A1 => n10590, A2 => n16786, ZN => n30228);
   U14425 : NOR2_X1 port map( A1 => n15794, A2 => n10383, ZN => n11197);
   U14443 : NAND2_X2 port map( A1 => n31447, A2 => n10186, ZN => n27275);
   U14444 : NAND2_X2 port map( A1 => n30193, A2 => n35870, ZN => n15267);
   U14447 : XOR2_X1 port map( A1 => n12903, A2 => n1902, Z => n12850);
   U14468 : OAI21_X1 port map( A1 => n14968, A2 => n31269, B => n31268, ZN => 
                           n7478);
   U14470 : NAND2_X1 port map( A1 => n14968, A2 => n1186, ZN => n31268);
   U14472 : INV_X2 port map( I => n14987, ZN => n31269);
   U14479 : XOR2_X1 port map( A1 => n26521, A2 => n9301, Z => n9300);
   U14485 : INV_X2 port map( I => n20864, ZN => n31270);
   U14504 : INV_X2 port map( I => n31272, ZN => n31494);
   U14511 : NAND2_X2 port map( A1 => n31274, A2 => n16220, ZN => n27292);
   U14520 : BUF_X2 port map( I => n37661, Z => n31275);
   U14560 : NAND2_X2 port map( A1 => n2955, A2 => n13466, ZN => n17008);
   U14561 : XNOR2_X1 port map( A1 => n28997, A2 => n38222, ZN => n29139);
   U14565 : INV_X2 port map( I => n31278, ZN => n14704);
   U14567 : XOR2_X1 port map( A1 => n25296, A2 => n30761, Z => n24976);
   U14582 : XOR2_X1 port map( A1 => n2959, A2 => n24920, Z => n15195);
   U14583 : XOR2_X1 port map( A1 => n31281, A2 => n24977, Z => n20514);
   U14601 : OR2_X1 port map( A1 => n28114, A2 => n13457, Z => n32485);
   U14603 : AOI21_X2 port map( A1 => n3527, A2 => n19476, B => n6044, ZN => 
                           n9828);
   U14619 : OR2_X1 port map( A1 => n19085, A2 => n5530, Z => n11398);
   U14639 : NOR2_X2 port map( A1 => n26001, A2 => n5753, ZN => n25897);
   U14658 : XOR2_X1 port map( A1 => n25159, A2 => n30405, Z => n31289);
   U14661 : NAND2_X2 port map( A1 => n16883, A2 => n16031, ZN => n23808);
   U14673 : INV_X2 port map( I => n31294, ZN => n17509);
   U14680 : NOR2_X1 port map( A1 => n8165, A2 => n993, ZN => n31806);
   U14681 : XOR2_X1 port map( A1 => n33041, A2 => n31295, Z => n32306);
   U14683 : INV_X1 port map( I => n29051, ZN => n31295);
   U14688 : INV_X2 port map( I => n32536, ZN => n13744);
   U14693 : AND2_X1 port map( A1 => n19233, A2 => n17509, Z => n4053);
   U14695 : XOR2_X1 port map( A1 => n35350, A2 => n1215, Z => n7345);
   U14709 : XOR2_X1 port map( A1 => n25146, A2 => n24928, Z => n25172);
   U14722 : NAND2_X2 port map( A1 => n6019, A2 => n30052, ZN => n30054);
   U14729 : XOR2_X1 port map( A1 => n129, A2 => n11661, Z => n11663);
   U14747 : NAND2_X2 port map( A1 => n21445, A2 => n21845, ZN => n14868);
   U14751 : NAND2_X2 port map( A1 => n2765, A2 => n21864, ZN => n13055);
   U14755 : NOR2_X1 port map( A1 => n14635, A2 => n19955, ZN => n18234);
   U14756 : XOR2_X1 port map( A1 => n9154, A2 => n38291, Z => n599);
   U14774 : AND2_X1 port map( A1 => n23516, A2 => n23518, Z => n18388);
   U14775 : AND2_X2 port map( A1 => n24285, A2 => n24287, Z => n9922);
   U14786 : XOR2_X1 port map( A1 => n26357, A2 => n38219, Z => n16082);
   U14804 : NAND2_X2 port map( A1 => n5474, A2 => n25787, ZN => n26520);
   U14813 : NAND2_X2 port map( A1 => n9125, A2 => n9124, ZN => n22492);
   U14834 : XOR2_X1 port map( A1 => n1463, A2 => n19860, Z => n31314);
   U14856 : NAND2_X1 port map( A1 => n26093, A2 => n33258, ZN => n31318);
   U14867 : NAND2_X2 port map( A1 => n20236, A2 => n20237, ZN => n33644);
   U14873 : OR2_X1 port map( A1 => n1676, A2 => n36214, Z => n33679);
   U14878 : XOR2_X1 port map( A1 => n19103, A2 => n19100, Z => n24463);
   U14879 : NAND2_X2 port map( A1 => n7323, A2 => n31322, ZN => n25867);
   U14880 : NOR2_X1 port map( A1 => n7528, A2 => n12673, ZN => n12785);
   U14892 : NOR2_X2 port map( A1 => n36752, A2 => n37105, ZN => n5653);
   U14906 : INV_X4 port map( I => n2765, ZN => n12080);
   U14912 : XOR2_X1 port map( A1 => n10129, A2 => n31327, Z => n10132);
   U14917 : XOR2_X1 port map( A1 => n27819, A2 => n1938, Z => n31327);
   U14924 : NAND2_X2 port map( A1 => n4329, A2 => n11912, ZN => n33316);
   U14925 : INV_X2 port map( I => n31329, ZN => n5112);
   U14947 : NOR2_X2 port map( A1 => n31871, A2 => n6713, ZN => n11413);
   U14948 : INV_X2 port map( I => n29591, ZN => n29597);
   U14954 : AOI21_X1 port map( A1 => n20041, A2 => n20517, B => n11449, ZN => 
                           n33264);
   U14966 : XOR2_X1 port map( A1 => n17879, A2 => n31334, Z => n17878);
   U14968 : XOR2_X1 port map( A1 => n24927, A2 => n33311, Z => n31334);
   U14975 : INV_X2 port map( I => n31335, ZN => n2532);
   U14976 : XOR2_X1 port map( A1 => Plaintext(104), A2 => Key(104), Z => n31335
                           );
   U14985 : NAND2_X2 port map( A1 => n12130, A2 => n31343, ZN => n2553);
   U14991 : AND2_X1 port map( A1 => n775, A2 => n20616, Z => n14127);
   U14992 : INV_X2 port map( I => n31341, ZN => n10314);
   U14993 : XOR2_X1 port map( A1 => n10316, A2 => n10315, Z => n31341);
   U15008 : AND2_X1 port map( A1 => n26031, A2 => n35903, Z => n5981);
   U15028 : OR2_X2 port map( A1 => n20171, A2 => n14000, Z => n26674);
   U15029 : XOR2_X1 port map( A1 => n17957, A2 => n29248, Z => n13800);
   U15050 : NOR2_X1 port map( A1 => n7445, A2 => n35981, ZN => n31346);
   U15069 : AOI22_X2 port map( A1 => n24374, A2 => n31349, B1 => n13070, B2 => 
                           n24430, ZN => n24864);
   U15074 : NAND2_X1 port map( A1 => n38609, A2 => n16081, ZN => n31349);
   U15084 : NAND2_X2 port map( A1 => n14553, A2 => n138, ZN => n31984);
   U15087 : NAND2_X1 port map( A1 => n31350, A2 => n1192, ZN => n20487);
   U15115 : NAND2_X1 port map( A1 => n9821, A2 => n9822, ZN => n14169);
   U15123 : XOR2_X1 port map( A1 => n11899, A2 => n25293, Z => n9007);
   U15127 : XOR2_X1 port map( A1 => n20333, A2 => n13342, Z => n25293);
   U15146 : OAI21_X2 port map( A1 => n6491, A2 => n24710, B => n13046, ZN => 
                           n24701);
   U15150 : OR2_X1 port map( A1 => n14404, A2 => n28123, Z => n27107);
   U15154 : XOR2_X1 port map( A1 => n7137, A2 => n22587, Z => n22605);
   U15157 : INV_X2 port map( I => n20541, ZN => n19050);
   U15168 : NOR2_X1 port map( A1 => n23958, A2 => n24469, ZN => n17789);
   U15185 : NAND2_X2 port map( A1 => n11065, A2 => n11064, ZN => n17400);
   U15186 : NOR2_X2 port map( A1 => n11066, A2 => n10719, ZN => n11065);
   U15199 : NAND3_X2 port map( A1 => n31735, A2 => n27135, A3 => n31734, ZN => 
                           n12551);
   U15206 : XOR2_X1 port map( A1 => n19536, A2 => n23939, Z => n23972);
   U15222 : INV_X1 port map( I => n30095, ZN => n30086);
   U15223 : AND2_X1 port map( A1 => n15085, A2 => n5753, Z => n10179);
   U15240 : NAND2_X2 port map( A1 => n31365, A2 => n7551, ZN => n10632);
   U15242 : XOR2_X1 port map( A1 => n31366, A2 => n38962, Z => Ciphertext(77));
   U15252 : NOR2_X2 port map( A1 => n31369, A2 => n9904, ZN => n12661);
   U15296 : XOR2_X1 port map( A1 => n31377, A2 => n893, Z => n32251);
   U15299 : XOR2_X1 port map( A1 => n29242, A2 => n12707, Z => n12939);
   U15303 : AND2_X1 port map( A1 => n28559, A2 => n31353, Z => n7615);
   U15305 : NOR2_X1 port map( A1 => n31378, A2 => n28402, ZN => n9355);
   U15307 : AOI21_X1 port map( A1 => n36827, A2 => n10544, B => n37804, ZN => 
                           n11680);
   U15308 : OAI22_X1 port map( A1 => n24162, A2 => n914, B1 => n124, B2 => 
                           n10152, ZN => n2674);
   U15309 : OR2_X1 port map( A1 => n28152, A2 => n28153, Z => n9168);
   U15322 : XOR2_X1 port map( A1 => Plaintext(16), A2 => Key(16), Z => n31381);
   U15323 : AND2_X1 port map( A1 => n25460, A2 => n31809, Z => n25008);
   U15336 : XOR2_X1 port map( A1 => n16062, A2 => n8482, Z => n32165);
   U15337 : OAI22_X2 port map( A1 => n15706, A2 => n6670, B1 => n6671, B2 => 
                           n6672, ZN => n33678);
   U15345 : XOR2_X1 port map( A1 => n27579, A2 => n3891, Z => n3887);
   U15353 : XOR2_X1 port map( A1 => n3953, A2 => n39804, Z => n17910);
   U15359 : OAI21_X1 port map( A1 => n37748, A2 => n39226, B => n38300, ZN => 
                           n31386);
   U15401 : INV_X4 port map( I => n5112, ZN => n14472);
   U15411 : AND2_X1 port map( A1 => n25820, A2 => n17791, Z => n11633);
   U15414 : NOR3_X1 port map( A1 => n39083, A2 => n31549, A3 => n30213, ZN => 
                           n7792);
   U15419 : NAND2_X2 port map( A1 => n12617, A2 => n1630, ZN => n23397);
   U15427 : OAI21_X2 port map( A1 => n31400, A2 => n31399, B => n27391, ZN => 
                           n18171);
   U15436 : XOR2_X1 port map( A1 => n507, A2 => n25298, Z => n13919);
   U15443 : XOR2_X1 port map( A1 => n10385, A2 => n34126, Z => n31401);
   U15453 : XOR2_X1 port map( A1 => n6641, A2 => n27696, Z => n20531);
   U15459 : NAND2_X2 port map( A1 => n18289, A2 => n7660, ZN => n25991);
   U15463 : AND2_X1 port map( A1 => n22320, A2 => n22319, Z => n33594);
   U15470 : NOR2_X1 port map( A1 => n23173, A2 => n34757, ZN => n22939);
   U15494 : NAND2_X2 port map( A1 => n1454, A2 => n18689, ZN => n4809);
   U15520 : XOR2_X1 port map( A1 => n33083, A2 => n26158, Z => n31414);
   U15526 : NAND2_X2 port map( A1 => n32091, A2 => n24753, ZN => n5888);
   U15543 : OAI21_X2 port map( A1 => n18456, A2 => n18455, B => n18454, ZN => 
                           n24694);
   U15544 : INV_X2 port map( I => n20512, ZN => n28023);
   U15547 : XOR2_X1 port map( A1 => n20511, A2 => n14641, Z => n20512);
   U15548 : NAND2_X1 port map( A1 => n33291, A2 => n8745, ZN => n3107);
   U15553 : NAND2_X1 port map( A1 => n38762, A2 => n4649, ZN => n13769);
   U15578 : XOR2_X1 port map( A1 => n12244, A2 => n29144, Z => n29037);
   U15584 : NAND3_X2 port map( A1 => n28359, A2 => n28357, A3 => n28358, ZN => 
                           n12244);
   U15595 : NOR2_X1 port map( A1 => n5926, A2 => n5927, ZN => n31424);
   U15596 : INV_X2 port map( I => n31426, ZN => n28231);
   U15605 : NAND2_X1 port map( A1 => n30311, A2 => n3869, ZN => n7773);
   U15609 : XOR2_X1 port map( A1 => n31427, A2 => n28412, Z => n28414);
   U15610 : XOR2_X1 port map( A1 => n28406, A2 => n28959, Z => n31427);
   U15611 : OAI22_X2 port map( A1 => n39706, A2 => n10477, B1 => n1609, B2 => 
                           n15751, ZN => n24353);
   U15612 : XNOR2_X1 port map( A1 => n1659, A2 => n15513, ZN => n32331);
   U15620 : AOI22_X2 port map( A1 => n21336, A2 => n21599, B1 => n20535, B2 => 
                           n17992, ZN => n17991);
   U15643 : NOR2_X2 port map( A1 => n29909, A2 => n29910, ZN => n29929);
   U15645 : OAI21_X2 port map( A1 => n17145, A2 => n18656, B => n31407, ZN => 
                           n17154);
   U15660 : AOI22_X1 port map( A1 => n30119, A2 => n16275, B1 => n16277, B2 => 
                           n30107, ZN => n31430);
   U15668 : XOR2_X1 port map( A1 => n11791, A2 => n33622, Z => n17021);
   U15669 : NAND3_X1 port map( A1 => n4986, A2 => n24393, A3 => n15018, ZN => 
                           n16450);
   U15676 : NAND2_X2 port map( A1 => n32404, A2 => n18050, ZN => n27773);
   U15687 : AOI21_X2 port map( A1 => n23441, A2 => n1290, B => n17960, ZN => 
                           n23442);
   U15726 : NAND2_X2 port map( A1 => n16932, A2 => n11026, ZN => n29144);
   U15738 : XOR2_X1 port map( A1 => n25039, A2 => n25318, Z => n4501);
   U15762 : AOI21_X2 port map( A1 => n5490, A2 => n1302, B => n31441, ZN => 
                           n5488);
   U15763 : NOR2_X2 port map( A1 => n18989, A2 => n23468, ZN => n31441);
   U15768 : OAI21_X1 port map( A1 => n31912, A2 => n31911, B => n968, ZN => 
                           n2569);
   U15770 : XOR2_X1 port map( A1 => n31442, A2 => n870, Z => n15774);
   U15772 : INV_X1 port map( I => n29903, ZN => n31444);
   U15779 : OR2_X1 port map( A1 => n35207, A2 => n18827, Z => n16071);
   U15780 : NAND2_X2 port map( A1 => n1295, A2 => n33840, ZN => n11453);
   U15816 : XOR2_X1 port map( A1 => n27722, A2 => n27753, Z => n19231);
   U15837 : NAND2_X2 port map( A1 => n1597, A2 => n37377, ZN => n6298);
   U15843 : XOR2_X1 port map( A1 => n29094, A2 => n29164, Z => n6537);
   U15844 : XOR2_X1 port map( A1 => n29058, A2 => n17880, Z => n29164);
   U15861 : NAND2_X2 port map( A1 => n14027, A2 => n1338, ZN => n2841);
   U15885 : NOR2_X2 port map( A1 => n19700, A2 => n26879, ZN => n26994);
   U15905 : NOR2_X2 port map( A1 => n32575, A2 => n38629, ZN => n28683);
   U15910 : NOR2_X1 port map( A1 => n24146, A2 => n1123, ZN => n31464);
   U15912 : INV_X2 port map( I => n1230, ZN => n20399);
   U15936 : XOR2_X1 port map( A1 => n24079, A2 => n20340, Z => n31466);
   U15937 : XOR2_X1 port map( A1 => n14309, A2 => n31576, Z => n2988);
   U15951 : NAND2_X2 port map( A1 => n1418, A2 => n28695, ZN => n28598);
   U15973 : OR2_X1 port map( A1 => n33786, A2 => n20276, Z => n23054);
   U16028 : NAND3_X2 port map( A1 => n3746, A2 => n23385, A3 => n3743, ZN => 
                           n9518);
   U16037 : NAND3_X1 port map( A1 => n33608, A2 => n33607, A3 => n29732, ZN => 
                           n31477);
   U16067 : NAND2_X2 port map( A1 => n3681, A2 => n3682, ZN => n22064);
   U16070 : NOR2_X1 port map( A1 => n3452, A2 => n31019, ZN => n19660);
   U16076 : NAND2_X2 port map( A1 => n31484, A2 => n20250, ZN => n19828);
   U16082 : NAND2_X2 port map( A1 => n6089, A2 => n6088, ZN => n9395);
   U16084 : XOR2_X1 port map( A1 => n5241, A2 => n19833, Z => n1880);
   U16086 : INV_X2 port map( I => n22350, ZN => n21288);
   U16093 : NAND2_X1 port map( A1 => n22350, A2 => n30315, ZN => n16267);
   U16094 : NAND2_X2 port map( A1 => n21716, A2 => n21717, ZN => n22350);
   U16095 : XOR2_X1 port map( A1 => n22570, A2 => n29657, Z => n644);
   U16130 : NAND2_X2 port map( A1 => n3513, A2 => n4034, ZN => n27299);
   U16142 : NAND3_X2 port map( A1 => n34117, A2 => n25790, A3 => n1019, ZN => 
                           n18463);
   U16144 : INV_X1 port map( I => n33267, ZN => n33266);
   U16165 : XOR2_X1 port map( A1 => n19221, A2 => n29285, Z => n31492);
   U16176 : AOI21_X2 port map( A1 => n34064, A2 => n13349, B => n29348, ZN => 
                           n13000);
   U16183 : AND2_X1 port map( A1 => n9775, A2 => n9791, Z => n28101);
   U16201 : XOR2_X1 port map( A1 => n31500, A2 => n29130, Z => n13052);
   U16202 : XOR2_X1 port map( A1 => n29124, A2 => n35255, Z => n31500);
   U16208 : NAND3_X2 port map( A1 => n15881, A2 => n15882, A3 => n37238, ZN => 
                           n25778);
   U16226 : AOI21_X2 port map( A1 => n3912, A2 => n2690, B => n30427, ZN => n32
                           );
   U16240 : XOR2_X1 port map( A1 => n31505, A2 => n30452, Z => n32310);
   U16272 : OAI21_X2 port map( A1 => n16252, A2 => n29421, B => n13153, ZN => 
                           n1820);
   U16276 : NAND2_X2 port map( A1 => n9914, A2 => n6002, ZN => n29218);
   U16294 : NAND2_X2 port map( A1 => n38143, A2 => n29756, ZN => n29737);
   U16305 : BUF_X2 port map( I => n28848, Z => n31516);
   U16318 : CLKBUF_X4 port map( I => n12410, Z => n11658);
   U16323 : INV_X1 port map( I => n32477, ZN => n24270);
   U16344 : OAI21_X1 port map( A1 => n14093, A2 => n4640, B => n19435, ZN => 
                           n13726);
   U16347 : AOI22_X1 port map( A1 => n28773, A2 => n5662, B1 => n32286, B2 => 
                           n9353, ZN => n20430);
   U16361 : XOR2_X1 port map( A1 => Plaintext(185), A2 => Key(185), Z => n31507
                           );
   U16363 : XOR2_X1 port map( A1 => n22754, A2 => n31508, Z => n31559);
   U16367 : XOR2_X1 port map( A1 => n22570, A2 => n29221, Z => n31508);
   U16368 : XNOR2_X1 port map( A1 => n5816, A2 => n5815, ZN => n31509);
   U16374 : INV_X1 port map( I => n8475, ZN => n1409);
   U16379 : OR2_X1 port map( A1 => n33368, A2 => n31511, Z => n19111);
   U16385 : AND2_X1 port map( A1 => n17983, A2 => n29961, Z => n31512);
   U16386 : OAI21_X1 port map( A1 => n32480, A2 => n32479, B => n19750, ZN => 
                           n5665);
   U16416 : NAND2_X1 port map( A1 => n2823, A2 => n14209, ZN => n2774);
   U16420 : NAND2_X1 port map( A1 => n252, A2 => n6657, ZN => n6656);
   U16422 : INV_X2 port map( I => n15853, ZN => n16510);
   U16426 : NAND2_X1 port map( A1 => n16510, A2 => n21285, ZN => n10147);
   U16450 : NOR2_X1 port map( A1 => n20491, A2 => n20490, ZN => n26349);
   U16459 : AOI21_X1 port map( A1 => n13004, A2 => n10355, B => n37955, ZN => 
                           n32388);
   U16467 : NAND2_X2 port map( A1 => n31516, A2 => n29760, ZN => n31517);
   U16493 : NAND2_X1 port map( A1 => n2364, A2 => n735, ZN => n2363);
   U16509 : NAND3_X1 port map( A1 => n29416, A2 => n29408, A3 => n29409, ZN => 
                           n15042);
   U16535 : NOR2_X1 port map( A1 => n27404, A2 => n27390, ZN => n33888);
   U16539 : AOI22_X1 port map( A1 => n10293, A2 => n31968, B1 => n10292, B2 => 
                           n29888, ZN => n32470);
   U16556 : NAND2_X1 port map( A1 => n3538, A2 => n28330, ZN => n17522);
   U16557 : AND2_X2 port map( A1 => n16700, A2 => n31638, Z => n31518);
   U16579 : NAND3_X1 port map( A1 => n29997, A2 => n30042, A3 => n16328, ZN => 
                           n19196);
   U16583 : NOR2_X1 port map( A1 => n7583, A2 => n33346, ZN => n31660);
   U16610 : NOR2_X1 port map( A1 => n35023, A2 => n28366, ZN => n32315);
   U16616 : NAND2_X1 port map( A1 => n30129, A2 => n17192, ZN => n31693);
   U16623 : INV_X1 port map( I => n33324, ZN => n938);
   U16631 : AND2_X1 port map( A1 => n16542, A2 => n9528, Z => n31520);
   U16640 : NAND2_X1 port map( A1 => n9534, A2 => n12302, ZN => n10351);
   U16665 : INV_X2 port map( I => n13054, ZN => n27557);
   U16666 : AND2_X1 port map( A1 => n30260, A2 => n30259, Z => n14512);
   U16670 : NAND2_X1 port map( A1 => n8659, A2 => n14237, ZN => n31522);
   U16675 : BUF_X2 port map( I => n20207, Z => n7949);
   U16679 : INV_X2 port map( I => n28578, ZN => n3598);
   U16684 : NAND3_X1 port map( A1 => n26972, A2 => n15980, A3 => n26973, ZN => 
                           n15979);
   U16686 : NAND3_X1 port map( A1 => n26974, A2 => n26972, A3 => n32427, ZN => 
                           n16573);
   U16705 : NAND2_X1 port map( A1 => n29338, A2 => n38151, ZN => n3288);
   U16712 : NOR2_X1 port map( A1 => n1173, A2 => n18042, ZN => n29670);
   U16727 : OAI21_X1 port map( A1 => n1178, A2 => n29763, B => n17105, ZN => 
                           n17539);
   U16728 : NAND2_X1 port map( A1 => n13196, A2 => n13194, ZN => n31523);
   U16754 : NOR2_X1 port map( A1 => n28733, A2 => n13151, ZN => n8036);
   U16758 : NOR2_X1 port map( A1 => n16123, A2 => n18667, ZN => n18616);
   U16763 : AND2_X1 port map( A1 => n29403, A2 => n20159, Z => n13850);
   U16774 : INV_X2 port map( I => n20522, ZN => n1059);
   U16780 : AND2_X1 port map( A1 => n15601, A2 => n3462, Z => n3465);
   U16781 : NAND3_X1 port map( A1 => n5525, A2 => n19541, A3 => n11375, ZN => 
                           n28162);
   U16799 : OAI21_X2 port map( A1 => n28419, A2 => n8960, B => n7365, ZN => 
                           n7483);
   U16807 : NAND2_X1 port map( A1 => n33207, A2 => n13384, ZN => n32079);
   U16811 : NOR2_X1 port map( A1 => n1055, A2 => n771, ZN => n13263);
   U16822 : NOR2_X2 port map( A1 => n33548, A2 => n33547, ZN => n33546);
   U16825 : XOR2_X1 port map( A1 => n6536, A2 => n31525, Z => n33674);
   U16827 : XOR2_X1 port map( A1 => n19735, A2 => n29058, Z => n31525);
   U16834 : XOR2_X1 port map( A1 => n15077, A2 => n15453, Z => n31526);
   U16837 : NOR2_X1 port map( A1 => n139, A2 => n32925, ZN => n31527);
   U16844 : INV_X1 port map( I => n17347, ZN => n29546);
   U16852 : NAND2_X1 port map( A1 => n28577, A2 => n28578, ZN => n33195);
   U16859 : CLKBUF_X4 port map( I => n18806, Z => n3631);
   U16876 : AOI21_X2 port map( A1 => n4528, A2 => n1132, B => n4526, ZN => 
                           n31528);
   U16905 : NAND2_X1 port map( A1 => n26876, A2 => n32168, ZN => n32167);
   U16906 : NOR2_X1 port map( A1 => n26876, A2 => n36801, ZN => n32170);
   U16928 : OR2_X1 port map( A1 => n12428, A2 => n18720, Z => n29470);
   U16935 : NOR2_X1 port map( A1 => n28220, A2 => n4649, ZN => n31774);
   U16936 : NAND2_X1 port map( A1 => n31774, A2 => n1436, ZN => n9236);
   U16943 : NAND2_X1 port map( A1 => n15981, A2 => n17017, ZN => n23570);
   U16966 : NOR2_X1 port map( A1 => n11334, A2 => n26935, ZN => n32958);
   U16992 : NAND3_X1 port map( A1 => n30051, A2 => n9918, A3 => n1057, ZN => 
                           n20170);
   U16996 : INV_X1 port map( I => n9918, ZN => n30053);
   U16998 : OAI21_X1 port map( A1 => n12156, A2 => n27009, B => n5983, ZN => 
                           n27558);
   U17000 : XNOR2_X1 port map( A1 => n33243, A2 => n26448, ZN => n31537);
   U17005 : CLKBUF_X2 port map( I => n27737, Z => n32795);
   U17006 : OAI21_X1 port map( A1 => n33006, A2 => n26974, B => n5935, ZN => 
                           n15708);
   U17027 : AND2_X1 port map( A1 => n29600, A2 => n33746, Z => n31540);
   U17032 : NAND2_X1 port map( A1 => n20427, A2 => n19896, ZN => n20426);
   U17035 : NAND2_X1 port map( A1 => n29511, A2 => n29516, ZN => n33428);
   U17039 : NAND2_X1 port map( A1 => n19260, A2 => n29535, ZN => n29511);
   U17047 : NAND4_X1 port map( A1 => n2450, A2 => n2448, A3 => n9104, A4 => 
                           n29479, ZN => n33463);
   U17054 : AOI21_X2 port map( A1 => n23024, A2 => n23177, B => n14130, ZN => 
                           n23025);
   U17055 : XNOR2_X1 port map( A1 => n34545, A2 => n22615, ZN => n31541);
   U17060 : INV_X1 port map( I => n4604, ZN => n32185);
   U17062 : NAND2_X1 port map( A1 => n20288, A2 => n33358, ZN => n20287);
   U17067 : INV_X2 port map( I => n6287, ZN => n28453);
   U17079 : NAND2_X1 port map( A1 => n1052, A2 => n18829, ZN => n33565);
   U17091 : INV_X1 port map( I => n30432, ZN => n31545);
   U17092 : INV_X1 port map( I => n8275, ZN => n20623);
   U17093 : NOR2_X1 port map( A1 => n22364, A2 => n8275, ZN => n22226);
   U17094 : NAND2_X1 port map( A1 => n29870, A2 => n773, ZN => n18477);
   U17100 : NAND3_X1 port map( A1 => n31624, A2 => n2029, A3 => n25927, ZN => 
                           n11771);
   U17103 : INV_X1 port map( I => n2029, ZN => n3277);
   U17107 : INV_X2 port map( I => n22264, ZN => n14251);
   U17109 : NAND2_X1 port map( A1 => n32759, A2 => n16108, ZN => n11028);
   U17110 : NOR2_X1 port map( A1 => n8166, A2 => n8798, ZN => n31805);
   U17120 : NAND2_X1 port map( A1 => n38749, A2 => n24515, ZN => n32389);
   U17127 : INV_X1 port map( I => n5880, ZN => n32467);
   U17136 : NAND2_X1 port map( A1 => n8253, A2 => n5675, ZN => n8251);
   U17153 : XOR2_X1 port map( A1 => n18738, A2 => n18735, Z => n31546);
   U17160 : NAND2_X1 port map( A1 => n29413, A2 => n29410, ZN => n32234);
   U17169 : OAI21_X1 port map( A1 => n2335, A2 => n2334, B => n33649, ZN => 
                           n31548);
   U17170 : NAND2_X2 port map( A1 => n21300, A2 => n33651, ZN => n31549);
   U17178 : NAND3_X2 port map( A1 => n10998, A2 => n10999, A3 => n27059, ZN => 
                           n31551);
   U17200 : INV_X2 port map( I => n37632, ZN => n18039);
   U17202 : AOI22_X1 port map( A1 => n16596, A2 => n16597, B1 => n16595, B2 => 
                           n17369, ZN => n32353);
   U17208 : AOI21_X1 port map( A1 => n19272, A2 => n29555, B => n29546, ZN => 
                           n28904);
   U17209 : AND3_X2 port map( A1 => n6408, A2 => n9500, A3 => n6409, Z => 
                           n31552);
   U17216 : AND2_X1 port map( A1 => n19700, A2 => n14459, Z => n31555);
   U17218 : NOR2_X1 port map( A1 => n10764, A2 => n26098, ZN => n10765);
   U17224 : OAI22_X1 port map( A1 => n33023, A2 => n18140, B1 => n14400, B2 => 
                           n29445, ZN => n29448);
   U17225 : NAND2_X1 port map( A1 => n32671, A2 => n29445, ZN => n32670);
   U17226 : NOR2_X1 port map( A1 => n16295, A2 => n33707, ZN => n16494);
   U17244 : NAND2_X1 port map( A1 => n14891, A2 => n18667, ZN => n29262);
   U17254 : NAND2_X1 port map( A1 => n33555, A2 => n28738, ZN => n5968);
   U17294 : NAND2_X1 port map( A1 => n7529, A2 => n8646, ZN => n251);
   U17303 : NAND2_X1 port map( A1 => n15649, A2 => n5028, ZN => n31755);
   U17309 : NAND2_X1 port map( A1 => n13730, A2 => n1226, ZN => n6818);
   U17314 : NOR2_X1 port map( A1 => n29980, A2 => n29968, ZN => n32130);
   U17330 : INV_X1 port map( I => n9939, ZN => n10385);
   U17363 : XOR2_X1 port map( A1 => n16942, A2 => n20767, Z => n31564);
   U17366 : NAND3_X2 port map( A1 => n34116, A2 => n1781, A3 => n1777, ZN => 
                           n31566);
   U17374 : INV_X1 port map( I => n29033, ZN => n31720);
   U17376 : NAND2_X2 port map( A1 => n16050, A2 => n16051, ZN => n31568);
   U17391 : NOR2_X1 port map( A1 => n5921, A2 => n29721, ZN => n566);
   U17413 : XNOR2_X1 port map( A1 => n8502, A2 => n26570, ZN => n33165);
   U17415 : NAND2_X1 port map( A1 => n1036, A2 => n12966, ZN => n3048);
   U17423 : AND3_X2 port map( A1 => n8591, A2 => n8590, A3 => n31980, Z => 
                           n31569);
   U17424 : AND3_X2 port map( A1 => n8591, A2 => n8590, A3 => n31980, Z => 
                           n31570);
   U17426 : NAND2_X1 port map( A1 => n13094, A2 => n13414, ZN => n23440);
   U17428 : XOR2_X1 port map( A1 => n5566, A2 => n5565, Z => n31571);
   U17432 : INV_X1 port map( I => n13055, ZN => n22399);
   U17437 : AOI21_X2 port map( A1 => n1799, A2 => n4225, B => n24862, ZN => 
                           n1802);
   U17443 : XNOR2_X1 port map( A1 => n9151, A2 => n33504, ZN => n31575);
   U17444 : INV_X1 port map( I => n22968, ZN => n23035);
   U17454 : INV_X1 port map( I => n27697, ZN => n32811);
   U17459 : AND2_X2 port map( A1 => n16699, A2 => n11092, Z => n14947);
   U17466 : INV_X2 port map( I => n12892, ZN => n9987);
   U17469 : NOR2_X1 port map( A1 => n24432, A2 => n24431, ZN => n15828);
   U17486 : OAI22_X2 port map( A1 => n2842, A2 => n2841, B1 => n1671, B2 => 
                           n22182, ZN => n31576);
   U17504 : INV_X1 port map( I => n22490, ZN => n7118);
   U17518 : NAND2_X1 port map( A1 => n9329, A2 => n15540, ZN => n32284);
   U17531 : XOR2_X1 port map( A1 => n20303, A2 => n24949, Z => n31587);
   U17543 : AOI21_X1 port map( A1 => n13952, A2 => n17022, B => n13951, ZN => 
                           n13950);
   U17573 : NOR2_X2 port map( A1 => n12772, A2 => n24394, ZN => n11213);
   U17577 : NOR2_X1 port map( A1 => n29220, A2 => n10429, ZN => n13106);
   U17578 : XOR2_X1 port map( A1 => n4898, A2 => n6158, Z => n31595);
   U17580 : XOR2_X1 port map( A1 => n11017, A2 => n33850, Z => n31596);
   U17604 : NAND2_X1 port map( A1 => n23516, A2 => n19671, ZN => n4737);
   U17612 : AOI21_X1 port map( A1 => n23356, A2 => n39534, B => n33696, ZN => 
                           n24051);
   U17630 : OAI21_X1 port map( A1 => n25860, A2 => n33997, B => n33558, ZN => 
                           n3807);
   U17646 : INV_X1 port map( I => n9862, ZN => n15123);
   U17648 : XOR2_X1 port map( A1 => n21346, A2 => Key(25), Z => n31604);
   U17653 : XOR2_X1 port map( A1 => n10225, A2 => n10221, Z => n31605);
   U17664 : NOR2_X1 port map( A1 => n37632, A2 => n3462, ZN => n31911);
   U17667 : AND2_X2 port map( A1 => n17833, A2 => n6484, Z => n21475);
   U17669 : INV_X1 port map( I => n17833, ZN => n21476);
   U17692 : NAND2_X2 port map( A1 => n28749, A2 => n28622, ZN => n18990);
   U17709 : INV_X1 port map( I => n19478, ZN => n14602);
   U17714 : NAND2_X1 port map( A1 => n27936, A2 => n28109, ZN => n33613);
   U17721 : NOR2_X1 port map( A1 => n19768, A2 => n35973, ZN => n21414);
   U17736 : XOR2_X1 port map( A1 => n22200, A2 => n22201, Z => n31617);
   U17743 : XOR2_X1 port map( A1 => n31618, A2 => n18296, Z => Ciphertext(186))
                           ;
   U17746 : AOI22_X1 port map( A1 => n20074, A2 => n11701, B1 => n30247, B2 => 
                           n19663, ZN => n31618);
   U17747 : NOR2_X1 port map( A1 => n13258, A2 => n1722, ZN => n21659);
   U17748 : XOR2_X1 port map( A1 => n6447, A2 => Plaintext(134), Z => n13258);
   U17756 : INV_X1 port map( I => n29120, ZN => n1061);
   U17757 : OAI21_X2 port map( A1 => n24263, A2 => n31621, B => n16645, ZN => 
                           n24634);
   U17764 : NAND2_X2 port map( A1 => n14766, A2 => n33552, ZN => n28330);
   U17767 : XOR2_X1 port map( A1 => n15114, A2 => n31622, Z => n24247);
   U17768 : XOR2_X1 port map( A1 => n23870, A2 => n23871, Z => n31622);
   U17789 : NOR2_X2 port map( A1 => n7324, A2 => n15792, ZN => n28442);
   U17791 : NAND2_X2 port map( A1 => n24672, A2 => n12418, ZN => n25271);
   U17839 : XOR2_X1 port map( A1 => n31636, A2 => n672, Z => n4118);
   U17844 : NAND2_X2 port map( A1 => n31637, A2 => n12124, ZN => n15943);
   U17852 : XOR2_X1 port map( A1 => n27579, A2 => n18650, Z => n7829);
   U17855 : XOR2_X1 port map( A1 => n1938, A2 => n27557, Z => n27579);
   U17874 : OR2_X1 port map( A1 => n7847, A2 => n24538, Z => n32699);
   U17879 : OAI22_X1 port map( A1 => n29552, A2 => n29551, B1 => n29549, B2 => 
                           n29550, ZN => n29553);
   U17888 : NAND2_X1 port map( A1 => n3979, A2 => n27401, ZN => n31812);
   U17889 : AND2_X1 port map( A1 => n16252, A2 => n32946, Z => n31958);
   U17899 : AOI21_X2 port map( A1 => n5686, A2 => n1103, B => n5684, ZN => 
                           n9576);
   U17908 : OR2_X1 port map( A1 => n22499, A2 => n31649, Z => n31648);
   U17912 : OAI21_X2 port map( A1 => n16615, A2 => n7130, B => n23154, ZN => 
                           n23434);
   U17927 : BUF_X2 port map( I => n17499, Z => n31651);
   U17942 : XOR2_X1 port map( A1 => n31655, A2 => n23790, Z => n19577);
   U17949 : NAND2_X2 port map( A1 => n31656, A2 => n7799, ZN => n29045);
   U17952 : XOR2_X1 port map( A1 => n17417, A2 => n38228, Z => n27807);
   U17971 : NOR3_X1 port map( A1 => n15172, A2 => n14553, A3 => n9751, ZN => 
                           n14779);
   U17982 : NAND2_X2 port map( A1 => n6810, A2 => n17732, ZN => n18785);
   U17991 : XNOR2_X1 port map( A1 => n25181, A2 => n25086, ZN => n15779);
   U17999 : NAND2_X2 port map( A1 => n31665, A2 => n25889, ZN => n17309);
   U18024 : OR2_X1 port map( A1 => n27252, A2 => n36840, Z => n31668);
   U18030 : OR2_X1 port map( A1 => n2257, A2 => n22085, Z => n5345);
   U18032 : NOR2_X2 port map( A1 => n21481, A2 => n21480, ZN => n2257);
   U18042 : NAND2_X2 port map( A1 => n18591, A2 => n18594, ZN => n22263);
   U18047 : XOR2_X1 port map( A1 => n3655, A2 => n12233, Z => n4556);
   U18101 : AOI22_X2 port map( A1 => n29427, A2 => n1176, B1 => n15864, B2 => 
                           n357, ZN => n29284);
   U18102 : OAI22_X2 port map( A1 => n32671, A2 => n29445, B1 => n29446, B2 => 
                           n14422, ZN => n29427);
   U18106 : NAND2_X2 port map( A1 => n24646, A2 => n16238, ZN => n24793);
   U18116 : XOR2_X1 port map( A1 => n27001, A2 => n21176, Z => n31682);
   U18126 : XOR2_X1 port map( A1 => n31688, A2 => n16010, Z => n16009);
   U18150 : NAND2_X1 port map( A1 => n31693, A2 => n30127, ZN => n11446);
   U18170 : NAND3_X1 port map( A1 => n25756, A2 => n10563, A3 => n25754, ZN => 
                           n31695);
   U18179 : XOR2_X1 port map( A1 => n16336, A2 => n8654, Z => n13189);
   U18195 : XOR2_X1 port map( A1 => n29139, A2 => n28834, Z => n10365);
   U18206 : NAND2_X1 port map( A1 => n344, A2 => n21023, ZN => n20290);
   U18213 : NAND2_X2 port map( A1 => n16777, A2 => n30894, ZN => n15015);
   U18217 : OR2_X1 port map( A1 => n39815, A2 => n37045, Z => n33217);
   U18230 : AOI21_X2 port map( A1 => n31713, A2 => n31711, B => n13428, ZN => 
                           n7968);
   U18233 : AND2_X1 port map( A1 => n29925, A2 => n29924, Z => n31727);
   U18241 : NAND2_X2 port map( A1 => n45, A2 => n23034, ZN => n23119);
   U18243 : XOR2_X1 port map( A1 => n8873, A2 => n31718, Z => n31824);
   U18244 : XOR2_X1 port map( A1 => n27678, A2 => n30404, Z => n31718);
   U18247 : NAND2_X2 port map( A1 => n5458, A2 => n5459, ZN => n27687);
   U18250 : AOI22_X2 port map( A1 => n2971, A2 => n1031, B1 => n2972, B2 => 
                           n2439, ZN => n33730);
   U18262 : XOR2_X1 port map( A1 => n27592, A2 => n12613, Z => n27813);
   U18263 : NAND2_X2 port map( A1 => n53, A2 => n9739, ZN => n12613);
   U18272 : NAND2_X1 port map( A1 => n31595, A2 => n30000, ZN => n15328);
   U18276 : OAI21_X2 port map( A1 => n12706, A2 => n2340, B => n31723, ZN => 
                           n16050);
   U18280 : XOR2_X1 port map( A1 => n31725, A2 => n3666, Z => n21235);
   U18293 : NOR2_X2 port map( A1 => n5093, A2 => n16108, ZN => n4697);
   U18310 : INV_X2 port map( I => n31731, ZN => n4201);
   U18319 : XOR2_X1 port map( A1 => n25255, A2 => n25001, Z => n7958);
   U18320 : XOR2_X1 port map( A1 => n25278, A2 => n6759, Z => n25255);
   U18342 : NAND2_X2 port map( A1 => n31736, A2 => n22526, ZN => n23484);
   U18346 : NAND2_X2 port map( A1 => n31737, A2 => n18608, ZN => n24883);
   U18348 : NAND2_X1 port map( A1 => n24125, A2 => n38812, ZN => n31737);
   U18352 : XOR2_X1 port map( A1 => n7958, A2 => n7957, Z => n25683);
   U18353 : XOR2_X1 port map( A1 => n27779, A2 => n4709, Z => n11564);
   U18398 : NOR2_X1 port map( A1 => n19893, A2 => n35172, ZN => n31743);
   U18415 : XNOR2_X1 port map( A1 => n16565, A2 => n27715, ZN => n32181);
   U18420 : NOR2_X1 port map( A1 => n13217, A2 => n13029, ZN => n31749);
   U18439 : XOR2_X1 port map( A1 => n31752, A2 => n10955, Z => n14395);
   U18445 : INV_X2 port map( I => n39484, ZN => n1222);
   U18451 : AOI22_X2 port map( A1 => n5374, A2 => n27037, B1 => n13895, B2 => 
                           n5035, ZN => n27566);
   U18458 : AOI22_X2 port map( A1 => n23652, A2 => n36556, B1 => n32937, B2 => 
                           n31759, ZN => n18983);
   U18472 : NAND2_X2 port map( A1 => n9342, A2 => n9343, ZN => n8026);
   U18482 : INV_X2 port map( I => n31760, ZN => n32989);
   U18485 : XOR2_X1 port map( A1 => n2695, A2 => n31762, Z => n7993);
   U18486 : XOR2_X1 port map( A1 => n18655, A2 => n23689, Z => n31762);
   U18487 : OAI22_X1 port map( A1 => n8691, A2 => n11701, B1 => n30250, B2 => 
                           n11700, ZN => n32204);
   U18490 : NAND2_X2 port map( A1 => n11700, A2 => n30262, ZN => n8691);
   U18515 : XOR2_X1 port map( A1 => n10430, A2 => n3140, Z => n10390);
   U18523 : XOR2_X1 port map( A1 => n16898, A2 => n31771, Z => n22450);
   U18525 : INV_X2 port map( I => n10429, ZN => n31772);
   U18550 : NAND2_X2 port map( A1 => n32482, A2 => n17448, ZN => n27284);
   U18572 : NAND2_X1 port map( A1 => n7317, A2 => n692, ZN => n11257);
   U18585 : XOR2_X1 port map( A1 => n31779, A2 => n19407, Z => Ciphertext(149))
                           ;
   U18586 : OAI22_X1 port map( A1 => n30080, A2 => n30081, B1 => n19551, B2 => 
                           n19550, ZN => n31779);
   U18598 : XOR2_X1 port map( A1 => n19642, A2 => n35318, Z => n11612);
   U18625 : OAI22_X2 port map( A1 => n11639, A2 => n7494, B1 => n8411, B2 => 
                           n26623, ZN => n10301);
   U18626 : INV_X2 port map( I => n31784, ZN => n28279);
   U18662 : XOR2_X1 port map( A1 => n13931, A2 => n26280, Z => n31790);
   U18673 : NAND2_X2 port map( A1 => n28387, A2 => n18259, ZN => n28891);
   U18686 : XOR2_X1 port map( A1 => n27861, A2 => n2138, Z => n31794);
   U18700 : OAI21_X2 port map( A1 => n25563, A2 => n25716, B => n9132, ZN => 
                           n25564);
   U18707 : NOR2_X2 port map( A1 => n8693, A2 => n22468, ZN => n23478);
   U18714 : NAND2_X1 port map( A1 => n33457, A2 => n33456, ZN => n3593);
   U18717 : XOR2_X1 port map( A1 => n31801, A2 => n29321, Z => Ciphertext(25));
   U18719 : NAND2_X2 port map( A1 => n13947, A2 => n13950, ZN => n27404);
   U18721 : XOR2_X1 port map( A1 => n828, A2 => n14644, Z => n19830);
   U18731 : NOR3_X2 port map( A1 => n31806, A2 => n31805, A3 => n37241, ZN => 
                           n8169);
   U18737 : INV_X2 port map( I => n27810, ZN => n31807);
   U18754 : OAI22_X2 port map( A1 => n1183, A2 => n29815, B1 => n18222, B2 => 
                           n8677, ZN => n14216);
   U18759 : NAND2_X1 port map( A1 => n7173, A2 => n25379, ZN => n32826);
   U18773 : XOR2_X1 port map( A1 => n17627, A2 => n29092, Z => n31811);
   U18775 : OR2_X1 port map( A1 => n17032, A2 => n8604, Z => n28042);
   U18782 : NAND3_X2 port map( A1 => n11877, A2 => n22998, A3 => n20214, ZN => 
                           n3256);
   U18787 : XOR2_X1 port map( A1 => n7942, A2 => n22476, Z => n31815);
   U18803 : NAND3_X2 port map( A1 => n3070, A2 => n28134, A3 => n3069, ZN => 
                           n28685);
   U18818 : XOR2_X1 port map( A1 => n27501, A2 => n17349, Z => n27678);
   U18823 : XOR2_X1 port map( A1 => n31823, A2 => n38176, Z => n12824);
   U18824 : INV_X2 port map( I => n26582, ZN => n31823);
   U18839 : NOR3_X1 port map( A1 => n28105, A2 => n1205, A3 => n5352, ZN => 
                           n28106);
   U18846 : INV_X2 port map( I => n31824, ZN => n20056);
   U18866 : NAND2_X2 port map( A1 => n3861, A2 => n5579, ZN => n29855);
   U18867 : NOR2_X2 port map( A1 => n2346, A2 => n11830, ZN => n3861);
   U18869 : XOR2_X1 port map( A1 => n10371, A2 => n23743, Z => n6388);
   U18876 : XOR2_X1 port map( A1 => n19188, A2 => n31830, Z => n33809);
   U18879 : NAND2_X2 port map( A1 => n23219, A2 => n23218, ZN => n23899);
   U18889 : NAND2_X1 port map( A1 => n30041, A2 => n5348, ZN => n7208);
   U18908 : XOR2_X1 port map( A1 => n27687, A2 => n27736, Z => n15548);
   U18910 : NAND2_X2 port map( A1 => n6875, A2 => n6874, ZN => n27736);
   U18922 : NAND2_X2 port map( A1 => n31835, A2 => n23158, ZN => n23430);
   U18927 : AND2_X1 port map( A1 => n19768, A2 => n35973, Z => n18592);
   U18930 : NOR2_X1 port map( A1 => n2688, A2 => n9321, ZN => n31836);
   U18932 : XOR2_X1 port map( A1 => n1666, A2 => n1323, Z => n6546);
   U18951 : NAND2_X2 port map( A1 => n32851, A2 => n8019, ZN => n27153);
   U18952 : OAI22_X2 port map( A1 => n27350, A2 => n8830, B1 => n993, B2 => 
                           n19477, ZN => n26749);
   U18953 : INV_X2 port map( I => n31840, ZN => n26459);
   U18954 : XOR2_X1 port map( A1 => n31841, A2 => n29152, Z => n4354);
   U18972 : AOI22_X2 port map( A1 => n17856, A2 => n14176, B1 => n31848, B2 => 
                           n31847, ZN => n17751);
   U18978 : XOR2_X1 port map( A1 => n31851, A2 => n23565, Z => n18811);
   U18979 : NAND2_X2 port map( A1 => n31852, A2 => n9280, ZN => n24623);
   U18981 : XOR2_X1 port map( A1 => n19807, A2 => n25171, Z => n317);
   U18985 : NAND2_X2 port map( A1 => n13161, A2 => n19158, ZN => n22624);
   U18998 : AND2_X1 port map( A1 => n8688, A2 => n8679, Z => n31857);
   U19001 : NAND2_X2 port map( A1 => n33163, A2 => n16301, ZN => n32471);
   U19004 : XOR2_X1 port map( A1 => n32528, A2 => n26517, Z => n9301);
   U19084 : XOR2_X1 port map( A1 => Plaintext(142), A2 => Key(142), Z => n32370
                           );
   U19089 : OAI22_X2 port map( A1 => n6217, A2 => n23531, B1 => n23528, B2 => 
                           n6218, ZN => n23554);
   U19090 : XOR2_X1 port map( A1 => n17659, A2 => n31867, Z => n14254);
   U19097 : XOR2_X1 port map( A1 => n5520, A2 => n27733, Z => n32361);
   U19103 : XOR2_X1 port map( A1 => n23835, A2 => n7919, Z => n31869);
   U19109 : INV_X1 port map( I => n21249, ZN => n33547);
   U19122 : XOR2_X1 port map( A1 => n19081, A2 => n26542, Z => n26369);
   U19125 : NAND2_X2 port map( A1 => n25972, A2 => n9811, ZN => n26542);
   U19129 : XOR2_X1 port map( A1 => n22457, A2 => n3622, Z => n3621);
   U19145 : OAI22_X2 port map( A1 => n1440, A2 => n27940, B1 => n11732, B2 => 
                           n2717, ZN => n31876);
   U19158 : XOR2_X1 port map( A1 => n31880, A2 => n32842, Z => n2264);
   U19190 : AND2_X1 port map( A1 => n16224, A2 => n14557, Z => n12276);
   U19211 : XOR2_X1 port map( A1 => n5177, A2 => n5176, Z => n11617);
   U19230 : NAND2_X2 port map( A1 => n16006, A2 => n16007, ZN => n7485);
   U19258 : OAI21_X2 port map( A1 => n37169, A2 => n31893, B => n38317, ZN => 
                           n19356);
   U19271 : XOR2_X1 port map( A1 => n29090, A2 => n14099, Z => n6164);
   U19282 : XOR2_X1 port map( A1 => n1669, A2 => n22371, Z => n22597);
   U19297 : INV_X2 port map( I => n31897, ZN => n852);
   U19302 : XOR2_X1 port map( A1 => n26373, A2 => n5444, Z => n31897);
   U19308 : XNOR2_X1 port map( A1 => n10811, A2 => n15384, ZN => n29696);
   U19318 : XOR2_X1 port map( A1 => n14039, A2 => n31898, Z => n3552);
   U19324 : XOR2_X1 port map( A1 => n32092, A2 => n2996, Z => n29942);
   U19325 : NAND2_X2 port map( A1 => n9197, A2 => n24879, ZN => n18744);
   U19329 : AOI21_X2 port map( A1 => n39321, A2 => n3101, B => n31900, ZN => 
                           n3175);
   U19346 : INV_X2 port map( I => n37105, ZN => n32488);
   U19369 : XOR2_X1 port map( A1 => n33178, A2 => n18577, Z => n31909);
   U19377 : NOR2_X2 port map( A1 => n5817, A2 => n10713, ZN => n5871);
   U19380 : XOR2_X1 port map( A1 => n2229, A2 => n33676, Z => n33734);
   U19394 : XOR2_X1 port map( A1 => n31914, A2 => n29690, Z => Ciphertext(89));
   U19407 : AOI22_X2 port map( A1 => n32247, A2 => n1126, B1 => n31916, B2 => 
                           n17076, ZN => n32956);
   U19408 : XOR2_X1 port map( A1 => n8183, A2 => n25274, Z => n4238);
   U19420 : NAND2_X2 port map( A1 => n32089, A2 => n20972, ZN => n6141);
   U19436 : XOR2_X1 port map( A1 => n10225, A2 => n10221, Z => n26494);
   U19446 : NAND2_X2 port map( A1 => n20264, A2 => n31918, ZN => n31948);
   U19456 : INV_X2 port map( I => n31920, ZN => n12729);
   U19481 : NOR2_X1 port map( A1 => n27278, A2 => n27279, ZN => n31925);
   U19485 : NOR2_X1 port map( A1 => n35217, A2 => n12049, ZN => n10451);
   U19492 : AND2_X1 port map( A1 => n23515, A2 => n38292, Z => n2853);
   U19498 : XOR2_X1 port map( A1 => n31927, A2 => n23888, Z => n2806);
   U19539 : NAND3_X1 port map( A1 => n33656, A2 => n21160, A3 => n30484, ZN => 
                           n31932);
   U19560 : XOR2_X1 port map( A1 => n27466, A2 => n27858, Z => n12971);
   U19564 : INV_X1 port map( I => n23928, ZN => n32383);
   U19574 : XOR2_X1 port map( A1 => n22778, A2 => n31933, Z => n22780);
   U19604 : OAI21_X2 port map( A1 => n33281, A2 => n18962, B => n12232, ZN => 
                           n30184);
   U19621 : AOI22_X2 port map( A1 => n21925, A2 => n21469, B1 => n4057, B2 => 
                           n11411, ZN => n4056);
   U19646 : INV_X1 port map( I => n16610, ZN => n1510);
   U19655 : NAND2_X2 port map( A1 => n31940, A2 => n31939, ZN => n22161);
   U19658 : INV_X2 port map( I => n22008, ZN => n31939);
   U19661 : XOR2_X1 port map( A1 => n26588, A2 => n16294, Z => n26296);
   U19662 : XOR2_X1 port map( A1 => n22687, A2 => n12730, Z => n22490);
   U19686 : NAND2_X2 port map( A1 => n4903, A2 => n31946, ZN => n17094);
   U19693 : AOI21_X2 port map( A1 => n13774, A2 => n18244, B => n31947, ZN => 
                           n31946);
   U19696 : INV_X4 port map( I => n21099, ZN => n32168);
   U19709 : XOR2_X1 port map( A1 => n22391, A2 => n22510, Z => n8547);
   U19713 : AND3_X1 port map( A1 => n13233, A2 => n12924, A3 => n21270, Z => 
                           n13722);
   U19732 : XOR2_X1 port map( A1 => n4624, A2 => n22598, Z => n22392);
   U19733 : OAI22_X2 port map( A1 => n7132, A2 => n20375, B1 => n22499, B2 => 
                           n7131, ZN => n22598);
   U19740 : AND2_X1 port map( A1 => n29365, A2 => n37096, Z => n13274);
   U19749 : INV_X4 port map( I => n33140, ZN => n14423);
   U19751 : AOI21_X1 port map( A1 => n1473, A2 => n17142, B => n35500, ZN => 
                           n4089);
   U19756 : NOR2_X1 port map( A1 => n85, A2 => n2242, ZN => n12148);
   U19776 : NAND2_X2 port map( A1 => n13500, A2 => n13498, ZN => n27959);
   U19788 : NAND2_X1 port map( A1 => n21446, A2 => n21445, ZN => n21349);
   U19802 : NAND2_X1 port map( A1 => n31967, A2 => n19252, ZN => n33484);
   U19805 : OAI21_X1 port map( A1 => n32129, A2 => n32130, B => n18897, ZN => 
                           n31967);
   U19838 : XOR2_X1 port map( A1 => n27774, A2 => n27570, Z => n27539);
   U19843 : XNOR2_X1 port map( A1 => n12494, A2 => n12491, ZN => n31971);
   U19845 : OAI21_X2 port map( A1 => n31972, A2 => n33636, B => n21673, ZN => 
                           n11044);
   U19847 : XOR2_X1 port map( A1 => n32106, A2 => n19897, Z => n32766);
   U19850 : OR2_X1 port map( A1 => n25114, A2 => n25097, Z => n33896);
   U19851 : OAI21_X2 port map( A1 => n20927, A2 => n20928, B => n20925, ZN => 
                           n25114);
   U19855 : INV_X2 port map( I => n31976, ZN => n8529);
   U19856 : INV_X2 port map( I => n20960, ZN => n10231);
   U19859 : INV_X2 port map( I => n31978, ZN => n876);
   U19885 : XOR2_X1 port map( A1 => n13954, A2 => n32022, Z => n32678);
   U19894 : NOR2_X1 port map( A1 => n17412, A2 => n32304, ZN => n11677);
   U19895 : XOR2_X1 port map( A1 => n8516, A2 => n8514, Z => n32304);
   U19913 : INV_X2 port map( I => n3873, ZN => n31982);
   U19919 : XOR2_X1 port map( A1 => n17272, A2 => n30480, Z => n31983);
   U19920 : NAND3_X2 port map( A1 => n31985, A2 => n26659, A3 => n30352, ZN => 
                           n27249);
   U19922 : NAND2_X1 port map( A1 => n32142, A2 => n11864, ZN => n31985);
   U19929 : OR2_X1 port map( A1 => n2147, A2 => n28745, Z => n18201);
   U19935 : NOR2_X2 port map( A1 => n2347, A2 => n3861, ZN => n29858);
   U19951 : INV_X2 port map( I => n27919, ZN => n28215);
   U19961 : NOR2_X1 port map( A1 => n6217, A2 => n23532, ZN => n8269);
   U19971 : XOR2_X1 port map( A1 => n23910, A2 => n23884, Z => n23979);
   U19989 : OAI22_X2 port map( A1 => n23200, A2 => n11354, B1 => n13527, B2 => 
                           n33247, ZN => n33453);
   U19990 : NAND2_X1 port map( A1 => n13181, A2 => n26876, ZN => n13182);
   U19994 : AND2_X1 port map( A1 => n4947, A2 => n5112, Z => n32076);
   U20005 : AOI21_X1 port map( A1 => n5681, A2 => n5680, B => n927, ZN => n4677
                           );
   U20010 : XOR2_X1 port map( A1 => n33812, A2 => n1510, Z => n31999);
   U20011 : OR2_X1 port map( A1 => n24597, A2 => n36321, Z => n10056);
   U20012 : INV_X2 port map( I => n32001, ZN => n167);
   U20018 : NAND3_X2 port map( A1 => n18859, A2 => n32004, A3 => n33841, ZN => 
                           n11534);
   U20021 : XOR2_X1 port map( A1 => n12341, A2 => n29649, Z => n2997);
   U20026 : XOR2_X1 port map( A1 => n26518, A2 => n32003, Z => n5765);
   U20038 : NAND2_X2 port map( A1 => n28666, A2 => n33995, ZN => n4120);
   U20039 : AOI21_X2 port map( A1 => n10753, A2 => n953, B => n32011, ZN => 
                           n6965);
   U20043 : NAND2_X2 port map( A1 => n32926, A2 => n36496, ZN => n27244);
   U20067 : AND2_X1 port map( A1 => n32881, A2 => n15257, Z => n32018);
   U20071 : NAND2_X2 port map( A1 => n28184, A2 => n28185, ZN => n17397);
   U20076 : XOR2_X1 port map( A1 => n8742, A2 => n27558, Z => n3604);
   U20090 : XOR2_X1 port map( A1 => n11919, A2 => n30483, Z => n18580);
   U20091 : XOR2_X1 port map( A1 => n27786, A2 => n15401, Z => n11919);
   U20094 : XOR2_X1 port map( A1 => n23784, A2 => n6091, Z => n6090);
   U20095 : XOR2_X1 port map( A1 => n24070, A2 => n23903, Z => n23784);
   U20102 : OR2_X1 port map( A1 => n38822, A2 => n20566, Z => n13739);
   U20108 : XOR2_X1 port map( A1 => n25222, A2 => n32033, Z => n821);
   U20111 : XOR2_X1 port map( A1 => n25076, A2 => n31552, Z => n32033);
   U20114 : OR2_X1 port map( A1 => n15350, A2 => n10632, Z => n22340);
   U20130 : OR2_X1 port map( A1 => n5282, A2 => n32391, Z => n12946);
   U20144 : XOR2_X1 port map( A1 => n23722, A2 => n30446, Z => n24279);
   U20156 : XOR2_X1 port map( A1 => n14359, A2 => n32049, Z => n33958);
   U20161 : OR2_X1 port map( A1 => n28463, A2 => n28464, Z => n15709);
   U20181 : AOI21_X2 port map( A1 => n32916, A2 => n6469, B => n14578, ZN => 
                           n3116);
   U20182 : XOR2_X1 port map( A1 => n7944, A2 => n30775, Z => n6142);
   U20183 : NAND2_X2 port map( A1 => n7150, A2 => n7149, ZN => n7944);
   U20194 : OAI21_X2 port map( A1 => n4868, A2 => n4867, B => n32052, ZN => 
                           n32051);
   U20196 : XOR2_X1 port map( A1 => n16356, A2 => n29514, Z => n3299);
   U20197 : NAND2_X2 port map( A1 => n16256, A2 => n16272, ZN => n16356);
   U20200 : OAI22_X2 port map( A1 => n15952, A2 => n919, B1 => n15951, B2 => 
                           n32412, ZN => n22264);
   U20226 : XOR2_X1 port map( A1 => n32387, A2 => n9976, Z => n18345);
   U20227 : XOR2_X1 port map( A1 => n4587, A2 => n4588, Z => n21152);
   U20269 : XOR2_X1 port map( A1 => n32071, A2 => n13327, Z => n15598);
   U20275 : XOR2_X1 port map( A1 => n27547, A2 => n15548, Z => n32071);
   U20276 : OR2_X1 port map( A1 => n32535, A2 => n28621, Z => n9107);
   U20282 : XOR2_X1 port map( A1 => n8559, A2 => n8558, Z => n8557);
   U20283 : XOR2_X1 port map( A1 => n26544, A2 => n17051, Z => n33357);
   U20292 : NAND2_X2 port map( A1 => n26948, A2 => n20223, ZN => n26950);
   U20295 : NAND2_X2 port map( A1 => n16896, A2 => n13210, ZN => n10834);
   U20297 : XOR2_X1 port map( A1 => n36595, A2 => n29602, Z => n32073);
   U20313 : XOR2_X1 port map( A1 => n11571, A2 => n5002, Z => n11569);
   U20315 : XOR2_X1 port map( A1 => n13630, A2 => n13234, Z => n4671);
   U20322 : XOR2_X1 port map( A1 => n22760, A2 => n30329, Z => n32083);
   U20332 : INV_X2 port map( I => n7090, ZN => n20774);
   U20334 : NAND2_X1 port map( A1 => n18651, A2 => n18652, ZN => n18420);
   U20338 : NAND2_X2 port map( A1 => n32087, A2 => n15846, ZN => n25136);
   U20355 : XOR2_X1 port map( A1 => n24024, A2 => n12972, Z => n32090);
   U20383 : XOR2_X1 port map( A1 => n2995, A2 => n29161, Z => n32092);
   U20403 : XOR2_X1 port map( A1 => n23982, A2 => n13978, Z => n23801);
   U20408 : NAND3_X1 port map( A1 => n23161, A2 => n7071, A3 => n10436, ZN => 
                           n10438);
   U20415 : AND2_X1 port map( A1 => n13029, A2 => n23352, Z => n16456);
   U20423 : XOR2_X1 port map( A1 => n32097, A2 => n713, Z => n32096);
   U20431 : AND3_X1 port map( A1 => n13584, A2 => n1285, A3 => n32838, Z => 
                           n14291);
   U20432 : NAND2_X1 port map( A1 => n25068, A2 => n32101, ZN => n25070);
   U20451 : XOR2_X1 port map( A1 => n32103, A2 => n17402, Z => n10375);
   U20452 : XOR2_X1 port map( A1 => n13844, A2 => n22278, Z => n17402);
   U20458 : NAND2_X1 port map( A1 => n7955, A2 => n14423, ZN => n20869);
   U20466 : NAND2_X1 port map( A1 => n7778, A2 => n32388, ZN => n2239);
   U20468 : XOR2_X1 port map( A1 => n3638, A2 => n32110, Z => n11784);
   U20469 : XOR2_X1 port map( A1 => n3641, A2 => n20886, Z => n32110);
   U20482 : XOR2_X1 port map( A1 => n26205, A2 => n13324, Z => n33039);
   U20491 : XOR2_X1 port map( A1 => n32118, A2 => n12132, Z => n32486);
   U20501 : XOR2_X1 port map( A1 => n29071, A2 => n32120, Z => n18159);
   U20502 : INV_X1 port map( I => n29371, ZN => n32120);
   U20511 : XOR2_X1 port map( A1 => n38226, A2 => n19845, Z => n18510);
   U20520 : BUF_X2 port map( I => n33073, Z => n32123);
   U20530 : OAI21_X1 port map( A1 => n28049, A2 => n19410, B => n19435, ZN => 
                           n7409);
   U20540 : XOR2_X1 port map( A1 => n32126, A2 => n32125, Z => n8219);
   U20541 : XOR2_X1 port map( A1 => n8199, A2 => n20678, Z => n32125);
   U20547 : XOR2_X1 port map( A1 => n27648, A2 => n27819, Z => n32127);
   U20555 : XOR2_X1 port map( A1 => n32128, A2 => n30442, Z => n22887);
   U20592 : OAI22_X2 port map( A1 => n34459, A2 => n28669, B1 => n33337, B2 => 
                           n14209, ZN => n28798);
   U20593 : XOR2_X1 port map( A1 => n27698, A2 => n32137, Z => n17110);
   U20597 : INV_X2 port map( I => n755, ZN => n14458);
   U20605 : XOR2_X1 port map( A1 => n6124, A2 => n22670, Z => n32972);
   U20618 : INV_X4 port map( I => n32141, ZN => n9197);
   U20621 : NOR2_X2 port map( A1 => n15069, A2 => n298, ZN => n32141);
   U20643 : XOR2_X1 port map( A1 => n6930, A2 => n14307, Z => n28373);
   U20652 : XOR2_X1 port map( A1 => n32149, A2 => n27721, Z => n18447);
   U20660 : OAI22_X2 port map( A1 => n8017, A2 => n32039, B1 => n8792, B2 => 
                           n11044, ZN => n32151);
   U20679 : AOI22_X2 port map( A1 => n32152, A2 => n19007, B1 => n24403, B2 => 
                           n13412, ZN => n12307);
   U20686 : NAND2_X2 port map( A1 => n25767, A2 => n9379, ZN => n11293);
   U20688 : NAND2_X2 port map( A1 => n35015, A2 => n5753, ZN => n25767);
   U20689 : XOR2_X1 port map( A1 => n32154, A2 => n15400, Z => n32446);
   U20694 : XOR2_X1 port map( A1 => n27636, A2 => n5650, Z => n5649);
   U20697 : NOR2_X1 port map( A1 => n29267, A2 => n29276, ZN => n29268);
   U20699 : INV_X1 port map( I => n32176, ZN => n33668);
   U20700 : NOR2_X1 port map( A1 => n25585, A2 => n16867, ZN => n32156);
   U20703 : NOR2_X1 port map( A1 => n19609, A2 => n21823, ZN => n21675);
   U20712 : XNOR2_X1 port map( A1 => n23884, A2 => n1725, ZN => n33232);
   U20713 : AOI21_X1 port map( A1 => n15597, A2 => n18383, B => n15598, ZN => 
                           n17248);
   U20742 : INV_X2 port map( I => n32161, ZN => n15359);
   U20746 : XOR2_X1 port map( A1 => Plaintext(98), A2 => Key(98), Z => n32161);
   U20750 : AOI21_X2 port map( A1 => n21797, A2 => n1354, B => n32162, ZN => 
                           n16659);
   U20752 : NOR2_X2 port map( A1 => n1354, A2 => n32163, ZN => n32162);
   U20754 : INV_X2 port map( I => n15619, ZN => n32164);
   U20755 : AOI21_X1 port map( A1 => n34166, A2 => n27895, B => n28290, ZN => 
                           n14176);
   U20770 : NAND2_X2 port map( A1 => n19687, A2 => n32166, ZN => n27108);
   U20799 : XOR2_X1 port map( A1 => n33243, A2 => n26448, Z => n5639);
   U20809 : XOR2_X1 port map( A1 => n183, A2 => n32181, Z => n6285);
   U20810 : XOR2_X1 port map( A1 => n3393, A2 => n3392, Z => n15187);
   U20819 : NAND2_X1 port map( A1 => n32234, A2 => n32423, ZN => n32303);
   U20845 : XOR2_X1 port map( A1 => n18310, A2 => n7113, Z => n7112);
   U20846 : NAND2_X2 port map( A1 => n7114, A2 => n8023, ZN => n18310);
   U20850 : NAND2_X2 port map( A1 => n4297, A2 => n4296, ZN => n14139);
   U20852 : XOR2_X1 port map( A1 => n25105, A2 => n5058, Z => n25351);
   U20865 : BUF_X2 port map( I => n9470, Z => n32186);
   U20874 : XOR2_X1 port map( A1 => n32188, A2 => n20479, Z => Ciphertext(28));
   U20875 : AOI21_X1 port map( A1 => n32303, A2 => n29406, B => n32302, ZN => 
                           n13329);
   U20880 : NAND3_X1 port map( A1 => n18071, A2 => n17578, A3 => n14524, ZN => 
                           n23133);
   U20882 : XOR2_X1 port map( A1 => n33718, A2 => n8900, Z => n15913);
   U20894 : XOR2_X1 port map( A1 => n8163, A2 => n19932, Z => n25150);
   U20913 : OR2_X2 port map( A1 => n19226, A2 => n26921, Z => n26920);
   U20914 : NAND2_X1 port map( A1 => n4957, A2 => n14558, ZN => n2675);
   U20924 : XOR2_X1 port map( A1 => n29835, A2 => n29305, Z => n32203);
   U20929 : INV_X4 port map( I => n32956, ZN => n25048);
   U20939 : NOR2_X2 port map( A1 => n28532, A2 => n11413, ZN => n11412);
   U20944 : OAI21_X2 port map( A1 => n32208, A2 => n11008, B => n3438, ZN => 
                           n8519);
   U20954 : XOR2_X1 port map( A1 => n32308, A2 => n2529, Z => n2527);
   U20959 : XOR2_X1 port map( A1 => n32210, A2 => n2025, Z => n15907);
   U20963 : OAI22_X2 port map( A1 => n6517, A2 => n33864, B1 => n6519, B2 => 
                           n6518, ZN => n32230);
   U20973 : XOR2_X1 port map( A1 => n32211, A2 => n9446, Z => n2297);
   U20974 : XOR2_X1 port map( A1 => n23382, A2 => n23387, Z => n32211);
   U20998 : NAND2_X2 port map( A1 => n6506, A2 => n8683, ZN => n8120);
   U20999 : NAND2_X2 port map( A1 => n6171, A2 => n8121, ZN => n6506);
   U21001 : XOR2_X1 port map( A1 => n27782, A2 => n32217, Z => n9401);
   U21007 : XOR2_X1 port map( A1 => n27542, A2 => n32218, Z => n32217);
   U21024 : XOR2_X1 port map( A1 => n11880, A2 => n15010, Z => n32219);
   U21046 : BUF_X2 port map( I => n23639, Z => n32226);
   U21053 : XOR2_X1 port map( A1 => n32227, A2 => n25201, Z => n3645);
   U21056 : XOR2_X1 port map( A1 => n3647, A2 => n25203, Z => n32227);
   U21059 : INV_X1 port map( I => n28188, ZN => n14376);
   U21064 : MUX2_X1 port map( I0 => n13492, I1 => n28036, S => n28188, Z => 
                           n16567);
   U21101 : XOR2_X1 port map( A1 => n27617, A2 => n31163, Z => n27619);
   U21106 : NAND2_X1 port map( A1 => n30793, A2 => n20078, ZN => n6453);
   U21109 : NAND2_X2 port map( A1 => n11676, A2 => n27910, ZN => n15727);
   U21125 : XNOR2_X1 port map( A1 => n36075, A2 => n16864, ZN => n25264);
   U21148 : XOR2_X1 port map( A1 => n8336, A2 => n8333, Z => n13989);
   U21168 : MUX2_X1 port map( I0 => n30210, I1 => n14387, S => n30213, Z => 
                           n15420);
   U21172 : XOR2_X1 port map( A1 => n32354, A2 => n27710, Z => n8335);
   U21173 : XNOR2_X1 port map( A1 => n26538, A2 => n26339, ZN => n5176);
   U21183 : NOR2_X1 port map( A1 => n38732, A2 => n36991, ZN => n25538);
   U21208 : AND2_X1 port map( A1 => n5042, A2 => n32536, Z => n13301);
   U21233 : XNOR2_X1 port map( A1 => n14039, A2 => n29165, ZN => n29022);
   U21240 : NAND3_X2 port map( A1 => n12413, A2 => n3194, A3 => n3195, ZN => 
                           n20509);
   U21253 : NOR2_X1 port map( A1 => n23467, A2 => n23634, ZN => n23421);
   U21258 : BUF_X2 port map( I => n6205, Z => n32258);
   U21259 : OR2_X1 port map( A1 => n25990, A2 => n38548, Z => n32586);
   U21270 : OAI22_X1 port map( A1 => n30214, A2 => n31549, B1 => n14869, B2 => 
                           n30211, ZN => n32263);
   U21272 : NAND2_X1 port map( A1 => n9445, A2 => n1379, ZN => n11395);
   U21301 : INV_X4 port map( I => n12729, ZN => n14409);
   U21313 : NAND2_X1 port map( A1 => n32280, A2 => n26672, ZN => n11220);
   U21328 : XOR2_X1 port map( A1 => n14364, A2 => n32275, Z => n10134);
   U21329 : XOR2_X1 port map( A1 => n8940, A2 => n28500, Z => n32275);
   U21331 : XOR2_X1 port map( A1 => n39231, A2 => n30248, Z => n13115);
   U21333 : XOR2_X1 port map( A1 => n20609, A2 => n32276, Z => n22904);
   U21334 : XOR2_X1 port map( A1 => n20607, A2 => n22379, Z => n32276);
   U21337 : NOR2_X1 port map( A1 => n29654, A2 => n32290, ZN => n19412);
   U21349 : XOR2_X1 port map( A1 => n32106, A2 => n26402, Z => n26433);
   U21351 : INV_X2 port map( I => n27417, ZN => n1478);
   U21353 : XOR2_X1 port map( A1 => n25079, A2 => n25283, Z => n13596);
   U21367 : XOR2_X1 port map( A1 => n7829, A2 => n30481, Z => n7828);
   U21375 : NOR2_X1 port map( A1 => n19563, A2 => n27180, ZN => n32837);
   U21382 : NAND3_X1 port map( A1 => n18832, A2 => n19743, A3 => n18144, ZN => 
                           n20431);
   U21413 : XOR2_X1 port map( A1 => n32288, A2 => n1708, Z => Ciphertext(79));
   U21418 : XOR2_X1 port map( A1 => n635, A2 => n3241, Z => n11219);
   U21441 : XOR2_X1 port map( A1 => n32293, A2 => n6549, Z => n6548);
   U21445 : AND3_X1 port map( A1 => n14271, A2 => n1236, A3 => n26862, Z => 
                           n32563);
   U21451 : XOR2_X1 port map( A1 => n31591, A2 => n29411, Z => n28950);
   U21453 : NAND2_X2 port map( A1 => n9842, A2 => n32301, ZN => n24782);
   U21456 : OAI21_X1 port map( A1 => n32297, A2 => n11757, B => n36272, ZN => 
                           n32301);
   U21474 : INV_X2 port map( I => n26598, ZN => n1504);
   U21475 : NAND2_X2 port map( A1 => n26052, A2 => n26051, ZN => n26598);
   U21481 : AND2_X1 port map( A1 => n29405, A2 => n35272, Z => n32302);
   U21521 : XOR2_X1 port map( A1 => n38370, A2 => n35215, Z => n32308);
   U21540 : INV_X1 port map( I => n22419, ZN => n33806);
   U21553 : XOR2_X1 port map( A1 => n32312, A2 => n15273, Z => Ciphertext(104))
                           ;
   U21554 : OAI22_X1 port map( A1 => n5468, A2 => n32050, B1 => n5467, B2 => 
                           n3377, ZN => n32312);
   U21556 : INV_X2 port map( I => n33738, ZN => n32313);
   U21558 : XOR2_X1 port map( A1 => n15838, A2 => Plaintext(94), Z => n21885);
   U21606 : NOR2_X1 port map( A1 => n25576, A2 => n25577, ZN => n32325);
   U21608 : NOR2_X1 port map( A1 => n23003, A2 => n19823, ZN => n32327);
   U21633 : NAND2_X2 port map( A1 => n32332, A2 => n13462, ZN => n8059);
   U21645 : OR2_X1 port map( A1 => n14500, A2 => n14426, Z => n19290);
   U21646 : XOR2_X1 port map( A1 => n25093, A2 => n25132, Z => n20304);
   U21647 : NOR2_X2 port map( A1 => n12208, A2 => n30410, ZN => n25093);
   U21662 : XOR2_X1 port map( A1 => n1324, A2 => n22615, Z => n10797);
   U21663 : XOR2_X1 port map( A1 => n32339, A2 => n850, Z => n32986);
   U21665 : XOR2_X1 port map( A1 => n32340, A2 => n19801, Z => Ciphertext(18));
   U21667 : OAI22_X1 port map( A1 => n29268, A2 => n16233, B1 => n16232, B2 => 
                           n29278, ZN => n32340);
   U21679 : NAND2_X2 port map( A1 => n13741, A2 => n13742, ZN => n24759);
   U21680 : XOR2_X1 port map( A1 => n13383, A2 => n33037, Z => n709);
   U21690 : OAI21_X2 port map( A1 => n6270, A2 => n6271, B => n21809, ZN => 
                           n22238);
   U21704 : NOR3_X1 port map( A1 => n32796, A2 => n13042, A3 => n23101, ZN => 
                           n14578);
   U21739 : XOR2_X1 port map( A1 => n32353, A2 => n29051, Z => Ciphertext(80));
   U21748 : XOR2_X1 port map( A1 => n18004, A2 => n7028, Z => n26442);
   U21761 : NAND2_X2 port map( A1 => n2238, A2 => n2239, ZN => n8537);
   U21762 : XOR2_X1 port map( A1 => n32361, A2 => n5522, Z => n12909);
   U21771 : OAI21_X2 port map( A1 => n32584, A2 => n32585, B => n28181, ZN => 
                           n8087);
   U21775 : XOR2_X1 port map( A1 => n32369, A2 => n27569, Z => n11137);
   U21776 : XOR2_X1 port map( A1 => n33587, A2 => n27676, Z => n32369);
   U21778 : AOI21_X2 port map( A1 => n17484, A2 => n17483, B => n17482, ZN => 
                           n32675);
   U21781 : INV_X4 port map( I => n3662, ZN => n33669);
   U21782 : XOR2_X1 port map( A1 => n25214, A2 => n35268, Z => n3163);
   U21788 : XOR2_X1 port map( A1 => n29044, A2 => n14820, Z => n13177);
   U21796 : XOR2_X1 port map( A1 => n32375, A2 => n16440, Z => n16160);
   U21815 : XOR2_X1 port map( A1 => n32382, A2 => n2474, Z => n33193);
   U21822 : AOI22_X2 port map( A1 => n20749, A2 => n33842, B1 => n28291, B2 => 
                           n5469, ZN => n33059);
   U21824 : XOR2_X1 port map( A1 => n24001, A2 => n24000, Z => n32387);
   U21825 : XOR2_X1 port map( A1 => n3525, A2 => n3522, Z => n4352);
   U21826 : NOR2_X1 port map( A1 => n7361, A2 => n13653, ZN => n33905);
   U21829 : XOR2_X1 port map( A1 => n32239, A2 => n4117, Z => n23723);
   U21838 : NAND2_X1 port map( A1 => n32390, A2 => n32389, ZN => n12518);
   U21850 : AND2_X1 port map( A1 => n23619, A2 => n10480, Z => n15458);
   U21854 : NAND2_X2 port map( A1 => n19537, A2 => n32394, ZN => n13300);
   U21867 : XOR2_X1 port map( A1 => n32396, A2 => n5719, Z => n5012);
   U21868 : XOR2_X1 port map( A1 => n23745, A2 => n30371, Z => n32396);
   U21869 : XOR2_X1 port map( A1 => n17006, A2 => n16004, Z => n32890);
   U21878 : NAND2_X2 port map( A1 => n4280, A2 => n17841, ZN => n22711);
   U21913 : XNOR2_X1 port map( A1 => n14888, A2 => n14887, ZN => n32661);
   U21914 : AND2_X1 port map( A1 => n23574, A2 => n12154, Z => n5049);
   U21915 : XOR2_X1 port map( A1 => n1923, A2 => n32402, Z => n1921);
   U21916 : XOR2_X1 port map( A1 => n14386, A2 => n30403, Z => n32402);
   U21919 : NAND2_X2 port map( A1 => n2701, A2 => n15959, ZN => n15960);
   U21925 : AOI21_X1 port map( A1 => n1654, A2 => n9472, B => n39155, ZN => 
                           n5436);
   U21935 : XOR2_X1 port map( A1 => n1745, A2 => n29509, Z => n9497);
   U21940 : XOR2_X1 port map( A1 => n2651, A2 => n22616, Z => n2650);
   U21944 : XOR2_X1 port map( A1 => n12839, A2 => n35200, Z => n18737);
   U21946 : INV_X2 port map( I => n1921, ZN => n15461);
   U21955 : NAND2_X1 port map( A1 => n21435, A2 => n21358, ZN => n21665);
   U21974 : XOR2_X1 port map( A1 => n20608, A2 => n33990, Z => n20607);
   U21983 : NAND2_X1 port map( A1 => n11515, A2 => n37098, ZN => n8822);
   U21994 : NOR2_X2 port map( A1 => n12443, A2 => n17314, ZN => n9688);
   U22016 : XOR2_X1 port map( A1 => n35196, A2 => n19805, Z => n2119);
   U22025 : XOR2_X1 port map( A1 => n6363, A2 => n22565, Z => n32420);
   U22034 : XOR2_X1 port map( A1 => n22608, A2 => n18446, Z => n353);
   U22043 : AND2_X1 port map( A1 => n32666, A2 => n29409, Z => n32423);
   U22046 : INV_X1 port map( I => n37064, ZN => n33926);
   U22070 : XOR2_X1 port map( A1 => n17758, A2 => n26253, Z => n26457);
   U22076 : NOR3_X2 port map( A1 => n26035, A2 => n26036, A3 => n26239, ZN => 
                           n17758);
   U22081 : XOR2_X1 port map( A1 => n22609, A2 => n22733, Z => n32431);
   U22092 : NOR2_X2 port map( A1 => n25920, A2 => n25919, ZN => n18862);
   U22128 : OAI21_X2 port map( A1 => n1991, A2 => n1992, B => n25332, ZN => 
                           n4382);
   U22146 : NOR2_X2 port map( A1 => n28551, A2 => n37758, ZN => n8800);
   U22156 : XOR2_X1 port map( A1 => n33559, A2 => n32440, Z => n8116);
   U22160 : XOR2_X1 port map( A1 => n33420, A2 => n30461, Z => n32440);
   U22161 : XOR2_X1 port map( A1 => n11887, A2 => n32441, Z => n129);
   U22166 : XOR2_X1 port map( A1 => n295, A2 => n32464, Z => n32442);
   U22168 : XOR2_X1 port map( A1 => n29151, A2 => n30488, Z => n6158);
   U22176 : XOR2_X1 port map( A1 => n12988, A2 => n32443, Z => n11284);
   U22180 : XOR2_X1 port map( A1 => n4419, A2 => n27754, Z => n32443);
   U22198 : INV_X2 port map( I => n32446, ZN => n33955);
   U22200 : XOR2_X1 port map( A1 => n13791, A2 => n32447, Z => n18688);
   U22201 : XOR2_X1 port map( A1 => n27841, A2 => n18893, Z => n32447);
   U22208 : NAND3_X1 port map( A1 => n12259, A2 => n28147, A3 => n12258, ZN => 
                           n17214);
   U22225 : BUF_X2 port map( I => n1722, Z => n32456);
   U22232 : AOI21_X1 port map( A1 => n19017, A2 => n9422, B => n32457, ZN => 
                           n21365);
   U22250 : XOR2_X1 port map( A1 => n32460, A2 => n21294, Z => Ciphertext(146))
                           ;
   U22259 : AOI21_X1 port map( A1 => n20131, A2 => n20132, B => n32462, ZN => 
                           n20129);
   U22263 : OR2_X1 port map( A1 => n27395, A2 => n9037, Z => n32463);
   U22274 : XOR2_X1 port map( A1 => n29023, A2 => n32465, Z => n3938);
   U22283 : NOR2_X1 port map( A1 => n38141, A2 => n39018, ZN => n32466);
   U22288 : AOI22_X2 port map( A1 => n4887, A2 => n18575, B1 => n9764, B2 => 
                           n9763, ZN => n4886);
   U22295 : XOR2_X1 port map( A1 => n32470, A2 => n29875, Z => Ciphertext(120))
                           ;
   U22299 : OR3_X1 port map( A1 => n17072, A2 => n14881, A3 => n31006, Z => 
                           n26868);
   U22311 : NAND2_X1 port map( A1 => n1403, A2 => n20102, ZN => n15327);
   U22312 : NAND2_X2 port map( A1 => n18113, A2 => n32481, ZN => n26128);
   U22317 : XOR2_X1 port map( A1 => n13439, A2 => n11098, Z => n23852);
   U22320 : XOR2_X1 port map( A1 => n24050, A2 => n39038, Z => n33055);
   U22365 : INV_X2 port map( I => n32486, ZN => n25639);
   U22377 : XOR2_X1 port map( A1 => n32490, A2 => n19805, Z => n3560);
   U22378 : OAI21_X2 port map( A1 => n32495, A2 => n32494, B => n39321, ZN => 
                           n32871);
   U22379 : NOR2_X1 port map( A1 => n1116, A2 => n21042, ZN => n32494);
   U22404 : NAND2_X2 port map( A1 => n17055, A2 => n18019, ZN => n32535);
   U22411 : XOR2_X1 port map( A1 => n16427, A2 => n25848, Z => n32505);
   U22418 : INV_X2 port map( I => n20514, ZN => n33491);
   U22429 : AOI21_X2 port map( A1 => n17023, A2 => n17025, B => n8989, ZN => 
                           n8988);
   U22441 : XOR2_X1 port map( A1 => n32512, A2 => n28631, Z => n28899);
   U22454 : XOR2_X1 port map( A1 => n8732, A2 => n32516, Z => n19446);
   U22459 : XOR2_X1 port map( A1 => n29039, A2 => n29159, Z => n4223);
   U22463 : XOR2_X1 port map( A1 => n10256, A2 => n7564, Z => n28125);
   U22466 : XOR2_X1 port map( A1 => n32519, A2 => n29711, Z => Ciphertext(91));
   U22472 : NAND3_X2 port map( A1 => n20169, A2 => n10435, A3 => n20170, ZN => 
                           n30079);
   U22514 : XOR2_X1 port map( A1 => n23905, A2 => n16055, Z => n8113);
   U22517 : AND2_X1 port map( A1 => n15325, A2 => n23440, Z => n32526);
   U22526 : MUX2_X1 port map( I0 => n15867, I1 => n29797, S => n3096, Z => 
                           n5468);
   U22562 : XOR2_X1 port map( A1 => n32532, A2 => n10447, Z => n25700);
   U22572 : INV_X2 port map( I => n32534, ZN => n33948);
   U22581 : XOR2_X1 port map( A1 => n25243, A2 => n25218, Z => n17606);
   U22591 : NAND2_X1 port map( A1 => n19307, A2 => n15290, ZN => n22791);
   U22592 : INV_X2 port map( I => n32537, ZN => n15289);
   U22610 : XOR2_X1 port map( A1 => n6211, A2 => n32540, Z => n6550);
   U22619 : BUF_X2 port map( I => n21594, Z => n32544);
   U22631 : AOI22_X2 port map( A1 => n32546, A2 => n30544, B1 => n9268, B2 => 
                           n30768, ZN => n27470);
   U22639 : XOR2_X1 port map( A1 => n27767, A2 => n8059, Z => n15736);
   U22645 : NOR2_X2 port map( A1 => n27015, A2 => n32549, ZN => n27221);
   U22651 : OR2_X1 port map( A1 => n23234, A2 => n20788, Z => n2953);
   U22701 : NOR2_X2 port map( A1 => n14394, A2 => n26786, ZN => n26720);
   U22723 : NAND2_X2 port map( A1 => n3099, A2 => n3098, ZN => n26194);
   U22724 : OR2_X1 port map( A1 => n10338, A2 => n26695, Z => n231);
   U22725 : NAND2_X2 port map( A1 => n33142, A2 => n26270, ZN => n18549);
   U22745 : INV_X2 port map( I => n32556, ZN => n18077);
   U22761 : INV_X1 port map( I => n7742, ZN => n32559);
   U22769 : XOR2_X1 port map( A1 => n23911, A2 => n32562, Z => n10771);
   U22771 : NAND2_X2 port map( A1 => n18382, A2 => n18381, ZN => n23911);
   U22811 : XOR2_X1 port map( A1 => n32567, A2 => n4022, Z => n14347);
   U22813 : XOR2_X1 port map( A1 => n26324, A2 => n4021, Z => n32567);
   U22822 : XOR2_X1 port map( A1 => n19967, A2 => n34096, Z => n13116);
   U22826 : XOR2_X1 port map( A1 => n33176, A2 => n1262, Z => n19967);
   U22829 : NAND2_X2 port map( A1 => n16879, A2 => n14431, ZN => n6180);
   U22839 : NAND3_X1 port map( A1 => n29947, A2 => n29946, A3 => n39745, ZN => 
                           n29948);
   U22842 : NAND3_X1 port map( A1 => n11181, A2 => n17286, A3 => n31598, ZN => 
                           n32572);
   U22851 : NAND2_X2 port map( A1 => n4529, A2 => n6797, ZN => n6795);
   U22863 : XOR2_X1 port map( A1 => n19254, A2 => n29970, Z => n33862);
   U22870 : NAND2_X2 port map( A1 => n6808, A2 => n4917, ZN => n19254);
   U22875 : INV_X4 port map( I => n25639, ZN => n33130);
   U22923 : INV_X2 port map( I => n32579, ZN => n9242);
   U22927 : XOR2_X1 port map( A1 => n9400, A2 => n9401, Z => n32579);
   U22928 : INV_X1 port map( I => n11353, ZN => n28027);
   U22938 : XOR2_X1 port map( A1 => n25193, A2 => n24932, Z => n6306);
   U22939 : NAND2_X2 port map( A1 => n15877, A2 => n24491, ZN => n25193);
   U22946 : NOR2_X2 port map( A1 => n33249, A2 => n34016, ZN => n11703);
   U22947 : XOR2_X1 port map( A1 => n32581, A2 => n8059, Z => n13283);
   U22949 : INV_X2 port map( I => n33470, ZN => n32581);
   U22966 : NAND2_X2 port map( A1 => n4193, A2 => n3809, ZN => n4192);
   U22967 : NOR2_X2 port map( A1 => n18832, A2 => n12406, ZN => n32584);
   U22970 : NAND2_X2 port map( A1 => n8697, A2 => n32588, ZN => n8742);
   U22997 : AND2_X1 port map( A1 => n1627, A2 => n37088, Z => n32594);
   U22998 : INV_X2 port map( I => n32599, ZN => n9797);
   U23021 : INV_X2 port map( I => n22887, ZN => n22804);
   U23036 : OAI21_X1 port map( A1 => n29658, A2 => n29662, B => n30295, ZN => 
                           n17368);
   U23139 : XOR2_X1 port map( A1 => n22642, A2 => n22441, Z => n6610);
   U23162 : NAND2_X2 port map( A1 => n17436, A2 => n17435, ZN => n4613);
   U23176 : INV_X2 port map( I => n11702, ZN => n32617);
   U23178 : NOR2_X1 port map( A1 => n1816, A2 => n15839, ZN => n21574);
   U23179 : NAND2_X2 port map( A1 => n24339, A2 => n24340, ZN => n8173);
   U23183 : NAND2_X1 port map( A1 => n17424, A2 => n29500, ZN => n32620);
   U23203 : NAND2_X1 port map( A1 => n3452, A2 => n23071, ZN => n32625);
   U23233 : OR2_X1 port map( A1 => n5044, A2 => n6159, Z => n11214);
   U23246 : XOR2_X1 port map( A1 => n8281, A2 => n33158, Z => n32638);
   U23247 : XOR2_X1 port map( A1 => n32639, A2 => n32910, Z => n20152);
   U23252 : NAND2_X2 port map( A1 => n19694, A2 => n26977, ZN => n27417);
   U23257 : OAI21_X2 port map( A1 => n26250, A2 => n26251, B => n20912, ZN => 
                           n27361);
   U23290 : NAND3_X2 port map( A1 => n32644, A2 => n17979, A3 => n32643, ZN => 
                           n25218);
   U23298 : XOR2_X1 port map( A1 => n30322, A2 => n4210, Z => n17988);
   U23325 : AOI22_X2 port map( A1 => n6058, A2 => n16363, B1 => n27979, B2 => 
                           n885, ZN => n32650);
   U23334 : OAI21_X2 port map( A1 => n17669, A2 => n17668, B => n12243, ZN => 
                           n12242);
   U23374 : NOR2_X1 port map( A1 => n27213, A2 => n4847, ZN => n11767);
   U23380 : NAND2_X2 port map( A1 => n10723, A2 => n25728, ZN => n32658);
   U23388 : INV_X2 port map( I => n17533, ZN => n11283);
   U23410 : XOR2_X1 port map( A1 => n9643, A2 => n36068, Z => n32660);
   U23416 : XOR2_X1 port map( A1 => n32662, A2 => n32661, Z => n32708);
   U23424 : BUF_X2 port map( I => n21951, Z => n32664);
   U23455 : NAND4_X1 port map( A1 => n29403, A2 => n29401, A3 => n29402, A4 => 
                           n29400, ZN => n32666);
   U23456 : NAND2_X2 port map( A1 => n33468, A2 => n32667, ZN => n22741);
   U23462 : AOI22_X2 port map( A1 => n6081, A2 => n6083, B1 => n32477, B2 => 
                           n33986, ZN => n24944);
   U23470 : OR2_X1 port map( A1 => n1755, A2 => n20405, Z => n33206);
   U23510 : XOR2_X1 port map( A1 => n28780, A2 => n32678, Z => n266);
   U23525 : OR2_X1 port map( A1 => n24712, A2 => n7506, Z => n24902);
   U23537 : XOR2_X1 port map( A1 => n5836, A2 => n22735, Z => n5835);
   U23556 : XOR2_X1 port map( A1 => n25126, A2 => n606, Z => n32685);
   U23560 : XOR2_X1 port map( A1 => n33690, A2 => n27689, Z => n32686);
   U23571 : NOR2_X2 port map( A1 => n16945, A2 => n7062, ZN => n6381);
   U23572 : XOR2_X1 port map( A1 => n20706, A2 => n27745, Z => n27791);
   U23581 : XOR2_X1 port map( A1 => n27713, A2 => n27548, Z => n13327);
   U23604 : NOR2_X1 port map( A1 => n15280, A2 => n33678, ZN => n33677);
   U23610 : XOR2_X1 port map( A1 => n32698, A2 => n20166, Z => n19605);
   U23649 : NAND2_X2 port map( A1 => n4531, A2 => n28453, ZN => n32702);
   U23650 : XOR2_X1 port map( A1 => n27859, A2 => n11919, Z => n12775);
   U23652 : INV_X2 port map( I => n32708, ZN => n33431);
   U23668 : NAND2_X1 port map( A1 => n17527, A2 => n17526, ZN => n17525);
   U23678 : NOR2_X1 port map( A1 => n22274, A2 => n15868, ZN => n16364);
   U23694 : NOR2_X2 port map( A1 => n5590, A2 => n5589, ZN => n5588);
   U23716 : XOR2_X1 port map( A1 => n32718, A2 => n19444, Z => n21184);
   U23728 : NAND3_X1 port map( A1 => n20597, A2 => n28758, A3 => n2022, ZN => 
                           n104);
   U23730 : NOR2_X1 port map( A1 => n18719, A2 => n37188, ZN => n32719);
   U23734 : NAND2_X1 port map( A1 => n6137, A2 => n26354, ZN => n6136);
   U23737 : XOR2_X1 port map( A1 => n17110, A2 => n9026, Z => n17767);
   U23811 : OAI21_X1 port map( A1 => n19398, A2 => n25429, B => n25679, ZN => 
                           n25396);
   U23812 : XOR2_X1 port map( A1 => n39723, A2 => n29920, Z => n14098);
   U23834 : XNOR2_X1 port map( A1 => n4341, A2 => n28891, ZN => n28838);
   U23840 : AOI21_X2 port map( A1 => n37622, A2 => n1293, B => n37064, ZN => 
                           n2369);
   U23845 : NAND2_X1 port map( A1 => n27137, A2 => n27347, ZN => n8166);
   U23877 : NAND2_X2 port map( A1 => n12077, A2 => n32675, ZN => n22066);
   U23883 : XOR2_X1 port map( A1 => n3117, A2 => n32746, Z => n33967);
   U23886 : XOR2_X1 port map( A1 => n29251, A2 => n29250, Z => n32746);
   U23890 : INV_X2 port map( I => n32750, ZN => n33963);
   U23923 : NAND2_X1 port map( A1 => n902, A2 => n28772, ZN => n515);
   U23948 : NAND2_X2 port map( A1 => n17228, A2 => n17229, ZN => n27046);
   U23958 : INV_X2 port map( I => n32760, ZN => n293);
   U23962 : XOR2_X1 port map( A1 => Key(3), A2 => Plaintext(3), Z => n32760);
   U23974 : NOR2_X1 port map( A1 => n24650, A2 => n36340, ZN => n32761);
   U24006 : XOR2_X1 port map( A1 => n3490, A2 => n3489, Z => n13365);
   U24009 : XOR2_X1 port map( A1 => Plaintext(150), A2 => Key(150), Z => n33073
                           );
   U24026 : NOR2_X1 port map( A1 => n4631, A2 => n19059, ZN => n32768);
   U24033 : XOR2_X1 port map( A1 => n26489, A2 => n26338, Z => n26538);
   U24052 : XOR2_X1 port map( A1 => n16431, A2 => n13326, Z => n32773);
   U24069 : NOR2_X2 port map( A1 => n26863, A2 => n15037, ZN => n14065);
   U24071 : NAND3_X2 port map( A1 => n15137, A2 => n18771, A3 => n24663, ZN => 
                           n24665);
   U24073 : NAND3_X2 port map( A1 => n12646, A2 => n11104, A3 => n5066, ZN => 
                           n32825);
   U24075 : XOR2_X1 port map( A1 => n20107, A2 => n32779, Z => n18183);
   U24078 : XOR2_X1 port map( A1 => n26346, A2 => n15078, Z => n32779);
   U24079 : XOR2_X1 port map( A1 => n14393, A2 => n27739, Z => n26169);
   U24090 : OR2_X1 port map( A1 => n22256, A2 => n1342, Z => n22258);
   U24114 : NAND2_X2 port map( A1 => n14139, A2 => n22262, ZN => n22080);
   U24150 : NAND2_X2 port map( A1 => n22086, A2 => n2696, ZN => n12964);
   U24160 : XOR2_X1 port map( A1 => Plaintext(190), A2 => Key(190), Z => n20685
                           );
   U24164 : NOR2_X1 port map( A1 => n20835, A2 => n33496, ZN => n32798);
   U24166 : NAND2_X2 port map( A1 => n32799, A2 => n2077, ZN => n3540);
   U24184 : INV_X2 port map( I => n32805, ZN => n19697);
   U24187 : XOR2_X1 port map( A1 => n21218, A2 => n21216, Z => n32805);
   U24188 : XOR2_X1 port map( A1 => n23866, A2 => n23867, Z => n2511);
   U24192 : INV_X2 port map( I => n32806, ZN => n735);
   U24194 : XOR2_X1 port map( A1 => n32807, A2 => n11947, Z => n5103);
   U24202 : NAND3_X1 port map( A1 => n22128, A2 => n3678, A3 => n15663, ZN => 
                           n3677);
   U24205 : XOR2_X1 port map( A1 => n7247, A2 => n24928, Z => n9390);
   U24210 : XOR2_X1 port map( A1 => n38816, A2 => n32811, Z => n767);
   U24214 : NOR2_X2 port map( A1 => n2362, A2 => n32814, ZN => n32813);
   U24217 : AND2_X1 port map( A1 => n26787, A2 => n26470, Z => n32814);
   U24224 : XOR2_X1 port map( A1 => n13193, A2 => n6561, Z => n17680);
   U24235 : INV_X2 port map( I => n32821, ZN => n33939);
   U24240 : INV_X2 port map( I => n32822, ZN => n281);
   U24251 : NAND3_X1 port map( A1 => n14132, A2 => n26134, A3 => n33909, ZN => 
                           n14131);
   U24263 : OR2_X2 port map( A1 => n37052, A2 => n13873, Z => n25566);
   U24268 : OAI22_X2 port map( A1 => n33586, A2 => n1591, B1 => n24244, B2 => 
                           n18329, ZN => n15955);
   U24272 : OAI21_X2 port map( A1 => n2333, A2 => n7539, B => n28530, ZN => 
                           n33649);
   U24278 : NAND2_X1 port map( A1 => n34016, A2 => n7900, ZN => n9287);
   U24285 : NAND2_X2 port map( A1 => n7253, A2 => n7252, ZN => n20156);
   U24317 : NOR2_X2 port map( A1 => n17602, A2 => n17600, ZN => n32829);
   U24327 : OR2_X1 port map( A1 => n37093, A2 => n11678, Z => n20808);
   U24330 : INV_X2 port map( I => n37086, ZN => n19978);
   U24356 : OR2_X1 port map( A1 => n8818, A2 => n33955, Z => n8370);
   U24361 : OR2_X1 port map( A1 => n29890, A2 => n6885, Z => n17526);
   U24366 : AND2_X1 port map( A1 => n17630, A2 => n23078, Z => n32877);
   U24368 : NAND2_X1 port map( A1 => n1424, A2 => n38860, ZN => n32833);
   U24383 : OAI21_X2 port map( A1 => n22275, A2 => n16351, B => n17576, ZN => 
                           n22761);
   U24399 : NAND2_X2 port map( A1 => n19503, A2 => n19501, ZN => n25900);
   U24403 : XOR2_X1 port map( A1 => n35220, A2 => n32836, Z => n14643);
   U24405 : INV_X1 port map( I => n29711, ZN => n32836);
   U24412 : AOI22_X2 port map( A1 => n17444, A2 => n16828, B1 => n14525, B2 => 
                           n29266, ZN => n29271);
   U24417 : XOR2_X1 port map( A1 => n35936, A2 => n38468, Z => n24000);
   U24435 : XOR2_X1 port map( A1 => n15450, A2 => n15220, Z => n3028);
   U24438 : XOR2_X1 port map( A1 => n6710, A2 => n33220, Z => n8151);
   U24453 : AOI21_X1 port map( A1 => n11181, A2 => n31533, B => n15773, ZN => 
                           n10831);
   U24455 : XOR2_X1 port map( A1 => n29260, A2 => n28948, Z => n28949);
   U24496 : NOR2_X1 port map( A1 => n27964, A2 => n20157, ZN => n14093);
   U24515 : NAND2_X1 port map( A1 => n37064, A2 => n23256, ZN => n2368);
   U24519 : AND2_X1 port map( A1 => n15627, A2 => n31049, Z => n32850);
   U24531 : OAI21_X1 port map( A1 => n28380, A2 => n20494, B => n37776, ZN => 
                           n28381);
   U24565 : NAND2_X1 port map( A1 => n18667, A2 => n30233, ZN => n14789);
   U24576 : INV_X2 port map( I => n32855, ZN => n14424);
   U24580 : XOR2_X1 port map( A1 => Plaintext(133), A2 => Key(133), Z => n32855
                           );
   U24589 : INV_X2 port map( I => n32856, ZN => n23125);
   U24612 : OAI21_X2 port map( A1 => n32857, A2 => n21528, B => n35071, ZN => 
                           n2991);
   U24615 : NAND2_X2 port map( A1 => n32860, A2 => n20629, ZN => n24049);
   U24616 : AOI22_X2 port map( A1 => n9621, A2 => n2692, B1 => n32616, B2 => 
                           n19119, ZN => n32860);
   U24629 : OAI21_X2 port map( A1 => n25497, A2 => n32867, B => n14490, ZN => 
                           n25899);
   U24643 : XOR2_X1 port map( A1 => n29158, A2 => n17452, Z => n6774);
   U24645 : NOR2_X1 port map( A1 => n30069, A2 => n30071, ZN => n30067);
   U24649 : XOR2_X1 port map( A1 => n28971, A2 => n19904, Z => n13954);
   U24654 : AOI21_X2 port map( A1 => n33829, A2 => n33472, B => n28445, ZN => 
                           n28971);
   U24666 : NAND2_X2 port map( A1 => n28140, A2 => n28119, ZN => n28345);
   U24740 : OAI21_X2 port map( A1 => n32878, A2 => n32877, B => n23183, ZN => 
                           n23349);
   U24760 : OAI21_X2 port map( A1 => n23504, A2 => n1133, B => n23505, ZN => 
                           n32883);
   U24762 : XOR2_X1 port map( A1 => n359, A2 => n22285, Z => n18291);
   U24785 : XOR2_X1 port map( A1 => n32884, A2 => n30122, Z => Ciphertext(162))
                           ;
   U24834 : INV_X2 port map( I => n22131, ZN => n32889);
   U24843 : INV_X2 port map( I => n1627, ZN => n1132);
   U24856 : XOR2_X1 port map( A1 => n36516, A2 => n10370, Z => n16153);
   U24868 : INV_X2 port map( I => n32893, ZN => n33933);
   U24891 : XOR2_X1 port map( A1 => n33660, A2 => n26453, Z => n17657);
   U24903 : XOR2_X1 port map( A1 => n28979, A2 => n18522, Z => n32895);
   U24919 : XOR2_X1 port map( A1 => n38560, A2 => n32896, Z => n3657);
   U24920 : XOR2_X1 port map( A1 => n26537, A2 => n748, Z => n8187);
   U24942 : OR2_X1 port map( A1 => n20517, A2 => n35242, Z => n15899);
   U24951 : XOR2_X1 port map( A1 => n6477, A2 => n8409, Z => n8408);
   U24954 : XOR2_X1 port map( A1 => n32903, A2 => n37112, Z => Ciphertext(183))
                           ;
   U24970 : XOR2_X1 port map( A1 => n33399, A2 => n17134, Z => n816);
   U24980 : AOI21_X2 port map( A1 => n23546, A2 => n31644, B => n23545, ZN => 
                           n23880);
   U25017 : OAI22_X2 port map( A1 => n21297, A2 => n1138, B1 => n21296, B2 => 
                           n23579, ZN => n33698);
   U25024 : INV_X2 port map( I => n8372, ZN => n27174);
   U25035 : XOR2_X1 port map( A1 => n17493, A2 => n30408, Z => n447);
   U25039 : XOR2_X1 port map( A1 => n24038, A2 => n23808, Z => n16030);
   U25059 : XOR2_X1 port map( A1 => n23904, A2 => n24067, Z => n19103);
   U25071 : NAND2_X2 port map( A1 => n16636, A2 => n22868, ZN => n33703);
   U25077 : XOR2_X1 port map( A1 => n10012, A2 => n25323, Z => n32910);
   U25078 : AOI21_X2 port map( A1 => n32911, A2 => n25537, B => n25536, ZN => 
                           n17803);
   U25095 : AOI21_X2 port map( A1 => n13149, A2 => n23578, B => n23257, ZN => 
                           n6054);
   U25104 : NAND3_X1 port map( A1 => n1224, A2 => n27379, A3 => n27378, ZN => 
                           n32913);
   U25117 : XOR2_X1 port map( A1 => n20448, A2 => n33837, Z => n14456);
   U25119 : XOR2_X1 port map( A1 => n26528, A2 => n646, Z => n32915);
   U25149 : MUX2_X1 port map( I0 => n4306, I1 => n38419, S => n33955, Z => 
                           n8369);
   U25176 : OAI21_X2 port map( A1 => n20469, A2 => n20468, B => n21668, ZN => 
                           n33929);
   U25199 : XOR2_X1 port map( A1 => n7936, A2 => n680, Z => n1986);
   U25215 : XOR2_X1 port map( A1 => n12431, A2 => n12432, Z => n6493);
   U25229 : NAND2_X2 port map( A1 => n17502, A2 => n30595, ZN => n33816);
   U25255 : NAND2_X2 port map( A1 => n946, A2 => n948, ZN => n32929);
   U25267 : AOI22_X2 port map( A1 => n3543, A2 => n5380, B1 => n3542, B2 => 
                           n23032, ZN => n3544);
   U25276 : XOR2_X1 port map( A1 => n17129, A2 => n19198, Z => n19955);
   U25288 : NAND2_X1 port map( A1 => n30111, A2 => n35186, ZN => n32933);
   U25299 : XOR2_X1 port map( A1 => n26334, A2 => n16830, Z => n32934);
   U25317 : AOI22_X2 port map( A1 => n12080, A2 => n37089, B1 => n22244, B2 => 
                           n8679, ZN => n2589);
   U25334 : OR3_X1 port map( A1 => n21042, A2 => n25639, A3 => n841, Z => 
                           n25360);
   U25351 : AOI21_X2 port map( A1 => n22064, A2 => n1341, B => n4045, ZN => 
                           n4441);
   U25370 : NOR3_X2 port map( A1 => n30340, A2 => n33453, A3 => n14606, ZN => 
                           n18747);
   U25381 : NAND2_X2 port map( A1 => n3993, A2 => n4324, ZN => n9037);
   U25393 : AOI21_X1 port map( A1 => n2211, A2 => n11344, B => n22324, ZN => 
                           n4619);
   U25397 : NAND2_X2 port map( A1 => n18855, A2 => n4116, ZN => n2008);
   U25426 : INV_X2 port map( I => n32951, ZN => n14553);
   U25427 : OAI21_X2 port map( A1 => n32953, A2 => n32952, B => n28415, ZN => 
                           n2270);
   U25435 : NOR2_X2 port map( A1 => n9599, A2 => n1068, ZN => n32953);
   U25440 : XOR2_X1 port map( A1 => n33865, A2 => n17223, Z => n8629);
   U25448 : NOR2_X1 port map( A1 => n4682, A2 => n12952, ZN => n9928);
   U25450 : XOR2_X1 port map( A1 => n31822, A2 => n32955, Z => n33372);
   U25452 : XOR2_X1 port map( A1 => n15481, A2 => n15480, Z => n32955);
   U25477 : AND2_X1 port map( A1 => n29740, A2 => n29739, Z => n33767);
   U25508 : XOR2_X1 port map( A1 => n16296, A2 => n29269, Z => n11525);
   U25533 : NAND2_X2 port map( A1 => n28385, A2 => n28384, ZN => n1775);
   U25581 : XOR2_X1 port map( A1 => n33129, A2 => n22492, Z => n11437);
   U25597 : NAND2_X2 port map( A1 => n21534, A2 => n16930, ZN => n133);
   U25599 : XNOR2_X1 port map( A1 => n9858, A2 => n30085, ZN => n33121);
   U25614 : NAND2_X1 port map( A1 => n36548, A2 => n35273, ZN => n32980);
   U25617 : XOR2_X1 port map( A1 => n28837, A2 => n29301, Z => n21084);
   U25622 : NAND3_X2 port map( A1 => n37776, A2 => n6405, A3 => n28458, ZN => 
                           n32983);
   U25624 : INV_X4 port map( I => n32984, ZN => n27235);
   U25625 : INV_X2 port map( I => n32985, ZN => n4083);
   U25628 : NAND2_X2 port map( A1 => n20823, A2 => n27236, ZN => n27829);
   U25711 : NAND2_X1 port map( A1 => n25327, A2 => n25484, ZN => n25374);
   U25726 : XOR2_X1 port map( A1 => n27080, A2 => n27079, Z => n7564);
   U25727 : OAI21_X2 port map( A1 => n16283, A2 => n33004, B => n584, ZN => 
                           n20387);
   U25728 : NOR2_X1 port map( A1 => n1151, A2 => n17118, ZN => n33004);
   U25739 : XOR2_X1 port map( A1 => n35404, A2 => n37112, Z => n33005);
   U25755 : AND2_X1 port map( A1 => n38198, A2 => n26055, Z => n13731);
   U25773 : XOR2_X1 port map( A1 => n5534, A2 => n20232, Z => n33007);
   U25778 : NAND2_X1 port map( A1 => n13522, A2 => n13521, ZN => n33028);
   U25784 : INV_X2 port map( I => n33008, ZN => n17097);
   U25805 : INV_X4 port map( I => n21308, ZN => n33771);
   U25810 : OR2_X1 port map( A1 => n10223, A2 => n3669, Z => n33011);
   U25821 : NAND2_X2 port map( A1 => n24630, A2 => n11271, ZN => n24526);
   U25829 : XOR2_X1 port map( A1 => n33013, A2 => n6049, Z => n5350);
   U25833 : XOR2_X1 port map( A1 => n10036, A2 => n30333, Z => n33013);
   U25856 : OR2_X1 port map( A1 => n16042, A2 => n27267, Z => n33017);
   U25881 : INV_X2 port map( I => n33023, ZN => n771);
   U25886 : NAND2_X1 port map( A1 => n18439, A2 => n18440, ZN => n20920);
   U25905 : NAND2_X2 port map( A1 => n33028, A2 => n33700, ZN => n13519);
   U25914 : XOR2_X1 port map( A1 => n26146, A2 => n26147, Z => n33029);
   U25925 : OAI21_X2 port map( A1 => n11386, A2 => n7260, B => n33030, ZN => 
                           n26596);
   U25929 : NAND2_X2 port map( A1 => n9111, A2 => n9112, ZN => n9106);
   U25930 : NOR2_X2 port map( A1 => n33034, A2 => n5810, ZN => n5807);
   U25931 : OAI22_X1 port map( A1 => n10747, A2 => n14379, B1 => n13584, B2 => 
                           n10659, ZN => n11134);
   U25941 : XOR2_X1 port map( A1 => n25267, A2 => n6411, Z => n6410);
   U25945 : NOR2_X2 port map( A1 => n37198, A2 => n7606, ZN => n27010);
   U25975 : NAND2_X1 port map( A1 => n28222, A2 => n200, ZN => n33048);
   U25978 : XOR2_X1 port map( A1 => n10957, A2 => n33049, Z => n11266);
   U25995 : XOR2_X1 port map( A1 => n24030, A2 => n19770, Z => n33049);
   U25996 : INV_X1 port map( I => n26286, ZN => n8558);
   U25998 : XOR2_X1 port map( A1 => n26286, A2 => n26228, Z => n26230);
   U26005 : NAND3_X2 port map( A1 => n26869, A2 => n27393, A3 => n26868, ZN => 
                           n27617);
   U26006 : BUF_X2 port map( I => n27365, Z => n33050);
   U26013 : INV_X2 port map( I => n19605, ZN => n28133);
   U26018 : NOR2_X1 port map( A1 => n11013, A2 => n11044, ZN => n11012);
   U26027 : INV_X2 port map( I => n33055, ZN => n16523);
   U26032 : NAND2_X2 port map( A1 => n24554, A2 => n33056, ZN => n26075);
   U26038 : INV_X2 port map( I => n33057, ZN => n2395);
   U26077 : NAND2_X2 port map( A1 => n33092, A2 => n12879, ZN => n10429);
   U26093 : XOR2_X1 port map( A1 => n33067, A2 => n6057, Z => n2000);
   U26099 : OAI21_X2 port map( A1 => n13263, A2 => n17089, B => n19244, ZN => 
                           n29403);
   U26103 : NAND2_X2 port map( A1 => n12684, A2 => n15708, ZN => n6686);
   U26105 : AND2_X1 port map( A1 => n26837, A2 => n13758, Z => n15512);
   U26116 : XOR2_X1 port map( A1 => n6307, A2 => n6304, Z => n835);
   U26128 : OAI22_X2 port map( A1 => n25510, A2 => n11834, B1 => n16247, B2 => 
                           n34574, ZN => n26338);
   U26157 : OR2_X1 port map( A1 => n33782, A2 => n22268, Z => n33072);
   U26160 : OR2_X1 port map( A1 => n12403, A2 => n8517, Z => n17848);
   U26184 : OAI21_X2 port map( A1 => n4473, A2 => n9155, B => n15743, ZN => 
                           n4159);
   U26190 : NAND2_X2 port map( A1 => n3006, A2 => n23502, ZN => n12822);
   U26198 : NAND2_X1 port map( A1 => n2429, A2 => n5630, ZN => n2428);
   U26219 : XOR2_X1 port map( A1 => n28954, A2 => n29304, Z => n28955);
   U26228 : XOR2_X1 port map( A1 => n2511, A2 => n2510, Z => n16816);
   U26231 : AND2_X1 port map( A1 => n6652, A2 => n5970, Z => n3612);
   U26241 : INV_X2 port map( I => n14318, ZN => n26833);
   U26247 : XOR2_X1 port map( A1 => n6007, A2 => n14319, Z => n14318);
   U26263 : XOR2_X1 port map( A1 => n21007, A2 => n2431, Z => n20622);
   U26265 : INV_X2 port map( I => n4498, ZN => n16328);
   U26270 : XNOR2_X1 port map( A1 => n29134, A2 => n29135, ZN => n4498);
   U26273 : XOR2_X1 port map( A1 => n33385, A2 => n20117, Z => n26747);
   U26276 : NOR2_X2 port map( A1 => n33156, A2 => n3691, ZN => n5449);
   U26280 : XOR2_X1 port map( A1 => n9091, A2 => n7346, Z => n13994);
   U26287 : NAND2_X2 port map( A1 => n6669, A2 => n15707, ZN => n22150);
   U26294 : XOR2_X1 port map( A1 => n28867, A2 => n19160, Z => n11017);
   U26308 : XOR2_X1 port map( A1 => n18001, A2 => n30402, Z => n22424);
   U26319 : XOR2_X1 port map( A1 => n22174, A2 => n22567, Z => n18597);
   U26331 : XOR2_X1 port map( A1 => n7475, A2 => n17423, Z => n23777);
   U26334 : NAND2_X2 port map( A1 => n22914, A2 => n22913, ZN => n17423);
   U26345 : OR2_X1 port map( A1 => n13728, A2 => n21805, Z => n10875);
   U26346 : XOR2_X1 port map( A1 => n10929, A2 => Key(59), Z => n13728);
   U26381 : OR2_X1 port map( A1 => n27854, A2 => n27498, Z => n5695);
   U26399 : OAI21_X2 port map( A1 => n18464, A2 => n14504, B => n18463, ZN => 
                           n11935);
   U26400 : NOR2_X1 port map( A1 => n14011, A2 => n23637, ZN => n7598);
   U26404 : XOR2_X1 port map( A1 => Plaintext(57), A2 => Key(57), Z => n7654);
   U26405 : XOR2_X1 port map( A1 => n27765, A2 => n682, Z => n33111);
   U26438 : XOR2_X1 port map( A1 => n33118, A2 => n4589, Z => n4588);
   U26444 : XOR2_X1 port map( A1 => n7603, A2 => n20843, Z => n33118);
   U26459 : OAI21_X1 port map( A1 => n14708, A2 => n21302, B => n15541, ZN => 
                           n15542);
   U26466 : XOR2_X1 port map( A1 => n13171, A2 => n33121, Z => n33120);
   U26467 : XNOR2_X1 port map( A1 => n26182, A2 => n25407, ZN => n33131);
   U26470 : NOR2_X1 port map( A1 => n33123, A2 => n30953, ZN => n7384);
   U26494 : INV_X1 port map( I => n4306, ZN => n898);
   U26496 : AND2_X1 port map( A1 => n18261, A2 => n4306, Z => n19139);
   U26501 : INV_X2 port map( I => n22566, ZN => n33129);
   U26503 : NOR2_X2 port map( A1 => n23600, A2 => n23601, ZN => n23605);
   U26530 : XOR2_X1 port map( A1 => n27840, A2 => n8896, Z => n33133);
   U26536 : XNOR2_X1 port map( A1 => n23661, A2 => n38350, ZN => n33524);
   U26545 : XOR2_X1 port map( A1 => n12411, A2 => n31575, Z => n11903);
   U26581 : NAND2_X2 port map( A1 => n7812, A2 => n7811, ZN => n7810);
   U26596 : AOI22_X2 port map( A1 => n10731, A2 => n19480, B1 => n30246, B2 => 
                           n39187, ZN => n30257);
   U26599 : AND2_X1 port map( A1 => n19341, A2 => n24394, Z => n16448);
   U26600 : NOR2_X1 port map( A1 => n38151, A2 => n14858, ZN => n33139);
   U26628 : INV_X2 port map( I => n33144, ZN => n862);
   U26632 : XOR2_X1 port map( A1 => n29111, A2 => n8285, Z => n8284);
   U26633 : NAND2_X2 port map( A1 => n33145, A2 => n15817, ZN => n22307);
   U26634 : NAND2_X2 port map( A1 => n33413, A2 => n15816, ZN => n33145);
   U26635 : NOR2_X1 port map( A1 => n8165, A2 => n33146, ZN => n12626);
   U26640 : NOR2_X2 port map( A1 => n26744, A2 => n26745, ZN => n27347);
   U26642 : INV_X2 port map( I => n33147, ZN => n1816);
   U26645 : OAI22_X2 port map( A1 => n1059, A2 => n20525, B1 => n30243, B2 => 
                           n30242, ZN => n30191);
   U26648 : NAND2_X2 port map( A1 => n17187, A2 => n17188, ZN => n26559);
   U26652 : XOR2_X1 port map( A1 => n23979, A2 => n11938, Z => n11117);
   U26665 : NOR2_X2 port map( A1 => n18087, A2 => n16934, ZN => n22676);
   U26672 : NAND2_X2 port map( A1 => n26833, A2 => n7527, ZN => n26831);
   U26674 : NAND2_X2 port map( A1 => n15184, A2 => n12923, ZN => n4604);
   U26706 : XOR2_X1 port map( A1 => n25193, A2 => n25090, Z => n25265);
   U26711 : XOR2_X1 port map( A1 => Plaintext(174), A2 => Key(174), Z => n695);
   U26715 : XOR2_X1 port map( A1 => n33153, A2 => n25150, Z => n9557);
   U26716 : XOR2_X1 port map( A1 => n24933, A2 => n16422, Z => n33153);
   U26720 : OAI21_X1 port map( A1 => n9668, A2 => n6287, B => n38155, ZN => 
                           n7296);
   U26721 : NOR2_X1 port map( A1 => n6414, A2 => n6416, ZN => n6776);
   U26733 : AND2_X1 port map( A1 => n17249, A2 => n37351, Z => n33156);
   U26736 : AND2_X1 port map( A1 => n20026, A2 => n12829, Z => n29385);
   U26753 : XOR2_X1 port map( A1 => n28805, A2 => n28804, Z => n30243);
   U26755 : XOR2_X1 port map( A1 => n27650, A2 => n8280, Z => n33158);
   U26758 : INV_X2 port map( I => n15718, ZN => n20102);
   U26759 : XOR2_X1 port map( A1 => n4898, A2 => n6158, Z => n15718);
   U26792 : XOR2_X1 port map( A1 => n16019, A2 => n29060, Z => n8516);
   U26824 : XOR2_X1 port map( A1 => n20618, A2 => n648, Z => n33166);
   U26839 : INV_X2 port map( I => n33170, ZN => n21546);
   U26851 : XOR2_X1 port map( A1 => Key(109), A2 => Plaintext(109), Z => n33170
                           );
   U26871 : OR2_X1 port map( A1 => n27385, A2 => n27064, Z => n33340);
   U26896 : XOR2_X1 port map( A1 => n20353, A2 => n20352, Z => n22603);
   U26912 : XOR2_X1 port map( A1 => n13634, A2 => n33400, Z => n14191);
   U26938 : XOR2_X1 port map( A1 => n23730, A2 => n23788, Z => n33179);
   U26942 : XOR2_X1 port map( A1 => Plaintext(7), A2 => Key(7), Z => n33324);
   U26945 : NAND2_X2 port map( A1 => n33180, A2 => n14572, ZN => n1326);
   U26958 : NAND2_X2 port map( A1 => n29473, A2 => n29470, ZN => n7303);
   U26969 : XOR2_X1 port map( A1 => n29168, A2 => n33183, Z => n9707);
   U26976 : XOR2_X1 port map( A1 => n15581, A2 => n33184, Z => n33183);
   U27006 : NAND2_X1 port map( A1 => n14946, A2 => n2189, ZN => n33186);
   U27011 : XOR2_X1 port map( A1 => n1817, A2 => n33188, Z => n25569);
   U27030 : NOR3_X1 port map( A1 => n1414, A2 => n28478, A3 => n38629, ZN => 
                           n3056);
   U27031 : AOI22_X2 port map( A1 => n21514, A2 => n21568, B1 => n15528, B2 => 
                           n33885, ZN => n16961);
   U27032 : NOR2_X2 port map( A1 => n3293, A2 => n3294, ZN => n15528);
   U27033 : XOR2_X1 port map( A1 => n38209, A2 => n26460, Z => n11050);
   U27057 : XOR2_X1 port map( A1 => n33192, A2 => n19775, Z => Ciphertext(172))
                           ;
   U27065 : INV_X2 port map( I => n33193, ZN => n2741);
   U27069 : XOR2_X1 port map( A1 => n25166, A2 => n33198, Z => n10971);
   U27079 : XOR2_X1 port map( A1 => n25165, A2 => n25275, Z => n33198);
   U27127 : XOR2_X1 port map( A1 => n12988, A2 => n5744, Z => n5743);
   U27128 : XOR2_X1 port map( A1 => n2867, A2 => n27511, Z => n12988);
   U27133 : XOR2_X1 port map( A1 => n22458, A2 => n33215, Z => n33936);
   U27141 : XOR2_X1 port map( A1 => n22648, A2 => n33216, Z => n33215);
   U27148 : NAND3_X2 port map( A1 => n14206, A2 => n33217, A3 => n14392, ZN => 
                           n14205);
   U27158 : XOR2_X1 port map( A1 => n29822, A2 => n33219, Z => n27881);
   U27167 : XOR2_X1 port map( A1 => n31522, A2 => n15745, Z => n33219);
   U27172 : XOR2_X1 port map( A1 => n6709, A2 => n18604, Z => n33220);
   U27181 : XOR2_X1 port map( A1 => n26570, A2 => n33223, Z => n14144);
   U27183 : XOR2_X1 port map( A1 => n33812, A2 => n19432, Z => n33223);
   U27184 : XNOR2_X1 port map( A1 => n14272, A2 => n4117, ZN => n792);
   U27186 : AND2_X1 port map( A1 => n19978, A2 => n33384, Z => n3011);
   U27199 : INV_X2 port map( I => n33227, ZN => n22567);
   U27202 : OAI21_X2 port map( A1 => n5576, A2 => n5577, B => n33228, ZN => 
                           n33227);
   U27216 : XOR2_X1 port map( A1 => n18359, A2 => n17528, Z => n12464);
   U27225 : XOR2_X1 port map( A1 => n9932, A2 => n1509, Z => n33233);
   U27250 : NAND2_X2 port map( A1 => n23754, A2 => n5740, ZN => n5897);
   U27257 : XOR2_X1 port map( A1 => n5571, A2 => n30450, Z => n2309);
   U27264 : XOR2_X1 port map( A1 => n33239, A2 => n3346, Z => n16284);
   U27268 : XOR2_X1 port map( A1 => n34498, A2 => n23957, Z => n33239);
   U27271 : XOR2_X1 port map( A1 => n22697, A2 => n22698, Z => n21163);
   U27281 : XOR2_X1 port map( A1 => n4091, A2 => n4090, Z => n33242);
   U27309 : NAND3_X2 port map( A1 => n24608, A2 => n31161, A3 => n19255, ZN => 
                           n18563);
   U27377 : NAND2_X2 port map( A1 => n33246, A2 => n29697, ZN => n29721);
   U27386 : XOR2_X1 port map( A1 => n23890, A2 => n7833, Z => n33248);
   U27391 : AND2_X1 port map( A1 => n19349, A2 => n38669, Z => n552);
   U27392 : BUF_X2 port map( I => n33506, Z => n33249);
   U27400 : NAND2_X1 port map( A1 => n4737, A2 => n7049, ZN => n13005);
   U27406 : NAND3_X1 port map( A1 => n15822, A2 => n15823, A3 => n20423, ZN => 
                           n33567);
   U27460 : OAI22_X2 port map( A1 => n33257, A2 => n2102, B1 => n23096, B2 => 
                           n1144, ZN => n23516);
   U27475 : NAND2_X2 port map( A1 => n9225, A2 => n9222, ZN => n22542);
   U27477 : XOR2_X1 port map( A1 => n21376, A2 => Key(68), Z => n33506);
   U27508 : NAND2_X1 port map( A1 => n27158, A2 => n27159, ZN => n33262);
   U27517 : OR2_X1 port map( A1 => n23473, A2 => n32601, Z => n15462);
   U27545 : BUF_X2 port map( I => n19644, Z => n33268);
   U27566 : XOR2_X1 port map( A1 => n15339, A2 => n33273, Z => n33272);
   U27570 : OR2_X1 port map( A1 => n13055, A2 => n22243, Z => n2588);
   U27593 : AND2_X1 port map( A1 => n22118, A2 => n22117, Z => n33282);
   U27616 : NAND2_X2 port map( A1 => n18216, A2 => n2954, ZN => n33284);
   U27623 : INV_X4 port map( I => n33286, ZN => n2341);
   U27639 : OR2_X1 port map( A1 => n22035, A2 => n33288, Z => n18953);
   U27644 : NOR2_X1 port map( A1 => n9486, A2 => n9484, ZN => n33291);
   U27660 : XOR2_X1 port map( A1 => n28913, A2 => n33295, Z => n17906);
   U27661 : XOR2_X1 port map( A1 => n36905, A2 => n5862, Z => n33295);
   U27663 : XOR2_X1 port map( A1 => n29065, A2 => n33296, Z => n17326);
   U27671 : XOR2_X1 port map( A1 => n29144, A2 => n19624, Z => n33296);
   U27675 : AOI21_X2 port map( A1 => n29873, A2 => n29869, B => n33297, ZN => 
                           n29890);
   U27680 : AND2_X1 port map( A1 => n15463, A2 => n16593, Z => n22871);
   U27715 : XOR2_X1 port map( A1 => n33300, A2 => n33299, Z => n846);
   U27721 : INV_X1 port map( I => n9989, ZN => n33299);
   U27723 : XOR2_X1 port map( A1 => n19879, A2 => n1009, Z => n33300);
   U27731 : NAND2_X2 port map( A1 => n25874, A2 => n36546, ZN => n25876);
   U27735 : OAI22_X2 port map( A1 => n33303, A2 => n9156, B1 => n26788, B2 => 
                           n26720, ZN => n27365);
   U27739 : OAI21_X2 port map( A1 => n14002, A2 => n14003, B => n14001, ZN => 
                           n14941);
   U27744 : XOR2_X1 port map( A1 => n22610, A2 => n32836, Z => n14610);
   U27758 : NAND2_X2 port map( A1 => n8662, A2 => n22398, ZN => n22610);
   U27769 : XOR2_X1 port map( A1 => n27645, A2 => n33310, Z => n33309);
   U27781 : INV_X2 port map( I => n20829, ZN => n33310);
   U27787 : XOR2_X1 port map( A1 => n33398, A2 => n33311, Z => n8748);
   U27798 : XOR2_X1 port map( A1 => n27598, A2 => n16972, Z => n33313);
   U27805 : XOR2_X1 port map( A1 => n33315, A2 => n22550, Z => n7120);
   U27808 : OR2_X1 port map( A1 => n37043, A2 => n10334, Z => n15230);
   U27841 : BUF_X2 port map( I => n6426, Z => n33318);
   U27845 : OR2_X1 port map( A1 => n25537, A2 => n25484, Z => n25464);
   U27851 : XOR2_X1 port map( A1 => n15056, A2 => n33319, Z => n881);
   U27854 : XOR2_X1 port map( A1 => n27672, A2 => n33320, Z => n33319);
   U27867 : INV_X1 port map( I => n29562, ZN => n33320);
   U27887 : XOR2_X1 port map( A1 => n5553, A2 => n26605, Z => n13544);
   U27890 : XOR2_X1 port map( A1 => n15609, A2 => n30448, Z => n407);
   U27901 : INV_X2 port map( I => n28456, ZN => n33325);
   U27913 : NAND2_X2 port map( A1 => n1823, A2 => n28434, ZN => n28456);
   U27932 : INV_X2 port map( I => n33326, ZN => n892);
   U27940 : INV_X1 port map( I => n1010, ZN => n26142);
   U27991 : XOR2_X1 port map( A1 => n18733, A2 => n17884, Z => n33334);
   U27994 : XOR2_X1 port map( A1 => n8920, A2 => n25329, Z => n13012);
   U28003 : XOR2_X1 port map( A1 => n39756, A2 => n38993, Z => n24981);
   U28004 : MUX2_X1 port map( I0 => n29662, I1 => n29659, S => n19297, Z => 
                           n16595);
   U28022 : XOR2_X1 port map( A1 => n11137, A2 => n7353, Z => n11136);
   U28030 : OR2_X1 port map( A1 => n15281, A2 => n10667, Z => n5934);
   U28070 : INV_X2 port map( I => n28596, ZN => n1418);
   U28071 : NAND2_X2 port map( A1 => n10150, A2 => n10151, ZN => n28596);
   U28109 : INV_X1 port map( I => n8365, ZN => n33346);
   U28119 : XOR2_X1 port map( A1 => n33350, A2 => n37109, Z => Ciphertext(7));
   U28166 : OAI21_X1 port map( A1 => n33946, A2 => n7705, B => n25429, ZN => 
                           n7956);
   U28168 : AOI21_X2 port map( A1 => n4423, A2 => n10408, B => n33355, ZN => 
                           n12198);
   U28172 : OAI21_X2 port map( A1 => n30225, A2 => n33963, B => n33362, ZN => 
                           n33355);
   U28173 : NOR2_X1 port map( A1 => n19157, A2 => n29409, ZN => n29397);
   U28199 : XOR2_X1 port map( A1 => n24632, A2 => n24631, Z => n24633);
   U28227 : NAND2_X1 port map( A1 => n29980, A2 => n33360, ZN => n7271);
   U28245 : NOR2_X1 port map( A1 => n29979, A2 => n29968, ZN => n33360);
   U28268 : INV_X1 port map( I => n21331, ZN => n33363);
   U28313 : XOR2_X1 port map( A1 => n27751, A2 => n18122, Z => n33364);
   U28390 : OAI22_X2 port map( A1 => n33366, A2 => n33365, B1 => n6220, B2 => 
                           n32974, ZN => n2915);
   U28426 : XOR2_X1 port map( A1 => n25122, A2 => n25121, Z => n25490);
   U28452 : XNOR2_X1 port map( A1 => n6527, A2 => n24025, ZN => n10413);
   U28461 : XOR2_X1 port map( A1 => n22571, A2 => n33371, Z => n11498);
   U28470 : XOR2_X1 port map( A1 => n22588, A2 => n11500, Z => n33371);
   U28475 : XOR2_X1 port map( A1 => n15118, A2 => n30455, Z => n23214);
   U28525 : OAI21_X2 port map( A1 => n31550, A2 => n8473, B => n33375, ZN => 
                           n14221);
   U28551 : NAND2_X2 port map( A1 => n20910, A2 => n20911, ZN => n23523);
   U28571 : AOI21_X1 port map( A1 => n2846, A2 => n27167, B => n6908, ZN => 
                           n33380);
   U28622 : NAND3_X2 port map( A1 => n23291, A2 => n23289, A3 => n23290, ZN => 
                           n24047);
   U28629 : XOR2_X1 port map( A1 => n11190, A2 => n19848, Z => n22607);
   U28643 : XOR2_X1 port map( A1 => n12613, A2 => n29334, Z => n10057);
   U28656 : XOR2_X1 port map( A1 => n36958, A2 => n26504, Z => n33388);
   U28657 : OAI21_X2 port map( A1 => n21639, A2 => n21638, B => n33389, ZN => 
                           n22362);
   U28658 : XOR2_X1 port map( A1 => n25102, A2 => n25103, Z => n25105);
   U28668 : XOR2_X1 port map( A1 => n9036, A2 => n19648, Z => n3668);
   U28708 : BUF_X2 port map( I => n26018, Z => n33395);
   U28750 : NAND3_X2 port map( A1 => n25530, A2 => n25528, A3 => n25529, ZN => 
                           n25797);
   U28758 : BUF_X2 port map( I => n9185, Z => n33398);
   U28825 : XOR2_X1 port map( A1 => n10427, A2 => n10426, Z => n10282);
   U28830 : AOI21_X2 port map( A1 => n21543, A2 => n19822, B => n33402, ZN => 
                           n16760);
   U28834 : NOR2_X1 port map( A1 => n16762, A2 => n21702, ZN => n33402);
   U28851 : XOR2_X1 port map( A1 => n11667, A2 => n7603, Z => n26276);
   U28864 : XOR2_X1 port map( A1 => n27810, A2 => n19649, Z => n11997);
   U28909 : XOR2_X1 port map( A1 => n5635, A2 => n33410, Z => n13725);
   U28912 : XOR2_X1 port map( A1 => n11883, A2 => n11882, Z => n33410);
   U28932 : NAND2_X2 port map( A1 => n18938, A2 => n18936, ZN => n5056);
   U28978 : NAND2_X2 port map( A1 => n21886, A2 => n547, ZN => n1847);
   U28993 : XOR2_X1 port map( A1 => n17310, A2 => n33415, Z => n22693);
   U29004 : AOI21_X1 port map( A1 => n29739, A2 => n29755, B => n29756, ZN => 
                           n33416);
   U29007 : OAI21_X2 port map( A1 => n3199, A2 => n7635, B => n33418, ZN => 
                           n28620);
   U29017 : XOR2_X1 port map( A1 => n33419, A2 => n29399, Z => Ciphertext(37));
   U29020 : AOI22_X1 port map( A1 => n29398, A2 => n29414, B1 => n29397, B2 => 
                           n29410, ZN => n33419);
   U29022 : XOR2_X1 port map( A1 => n5841, A2 => n7917, Z => n33420);
   U29028 : INV_X2 port map( I => n11136, ZN => n12406);
   U29037 : XOR2_X1 port map( A1 => n14385, A2 => n14374, Z => n9567);
   U29046 : XOR2_X1 port map( A1 => n18363, A2 => n18317, Z => n18316);
   U29052 : XOR2_X1 port map( A1 => n33426, A2 => n10823, Z => n2196);
   U29053 : XOR2_X1 port map( A1 => n9989, A2 => n26440, Z => n33426);
   U29078 : OR2_X1 port map( A1 => n2741, A2 => n12519, Z => n13114);
   U29083 : XOR2_X1 port map( A1 => n26227, A2 => n18399, Z => n26492);
   U29101 : NAND2_X2 port map( A1 => n25477, A2 => n25479, ZN => n25335);
   U29131 : XOR2_X1 port map( A1 => n3790, A2 => n3791, Z => n33429);
   U29132 : INV_X2 port map( I => n37117, ZN => n30145);
   U29158 : NOR2_X2 port map( A1 => n23245, A2 => n23244, ZN => n23695);
   U29278 : INV_X4 port map( I => n33512, ZN => n15643);
   U29300 : INV_X2 port map( I => n33446, ZN => n33950);
   U29332 : NAND2_X2 port map( A1 => n21247, A2 => n11970, ZN => n21246);
   U29393 : NAND2_X1 port map( A1 => n1596, A2 => n30833, ZN => n33456);
   U29396 : NAND2_X2 port map( A1 => n10937, A2 => n24172, ZN => n33459);
   U29410 : OR2_X1 port map( A1 => n15044, A2 => n29409, Z => n14517);
   U29465 : NAND2_X2 port map( A1 => n33911, A2 => n33462, ZN => n3601);
   U29469 : XOR2_X1 port map( A1 => n33463, A2 => n19760, Z => Ciphertext(49));
   U29477 : INV_X1 port map( I => n26060, ZN => n33464);
   U29508 : XOR2_X1 port map( A1 => n27689, A2 => n29206, Z => n3114);
   U29519 : XOR2_X1 port map( A1 => n8037, A2 => n8038, Z => n33466);
   U29544 : XOR2_X1 port map( A1 => n762, A2 => n30478, Z => n11814);
   U29562 : NAND2_X2 port map( A1 => n29181, A2 => n33476, ZN => n18829);
   U29565 : XOR2_X1 port map( A1 => n21055, A2 => n29143, Z => n33478);
   U29566 : NAND2_X1 port map( A1 => n20184, A2 => n13499, ZN => n13498);
   U29567 : INV_X2 port map( I => n33479, ZN => n21099);
   U29593 : AOI22_X1 port map( A1 => n30263, A2 => n13786, B1 => n30261, B2 => 
                           n31529, ZN => n7681);
   U29606 : XOR2_X1 port map( A1 => n33484, A2 => n1162, Z => Ciphertext(134));
   U29639 : NAND2_X2 port map( A1 => n33487, A2 => n22163, ZN => n16667);
   U29642 : NOR2_X2 port map( A1 => n19195, A2 => n19197, ZN => n29981);
   U29709 : NOR3_X2 port map( A1 => n7610, A2 => n12388, A3 => n24850, ZN => 
                           n14385);
   U29723 : CLKBUF_X12 port map( I => n15159, Z => n33495);
   U29765 : OAI22_X1 port map( A1 => n29007, A2 => n17192, B1 => n38164, B2 => 
                           n29008, ZN => n29012);
   U29792 : XOR2_X1 port map( A1 => n27770, A2 => n27771, Z => n27772);
   U29795 : OAI21_X1 port map( A1 => n21339, A2 => n1693, B => n7962, ZN => 
                           n6690);
   U29827 : XOR2_X1 port map( A1 => n33659, A2 => n16149, Z => n24421);
   U29836 : XOR2_X1 port map( A1 => n12437, A2 => n33515, Z => n22410);
   U29864 : OAI21_X1 port map( A1 => n31549, A2 => n33521, B => n33520, ZN => 
                           n8231);
   U29871 : XOR2_X1 port map( A1 => n25180, A2 => n25198, Z => n2959);
   U29886 : NAND3_X2 port map( A1 => n5895, A2 => n7130, A3 => n31019, ZN => 
                           n33526);
   U29887 : XOR2_X1 port map( A1 => n33527, A2 => n9557, Z => n7492);
   U29913 : NOR2_X2 port map( A1 => n13976, A2 => n33528, ZN => n15540);
   U29935 : INV_X1 port map( I => n30454, ZN => n33531);
   U29962 : OAI21_X2 port map( A1 => n9286, A2 => n9102, B => n33534, ZN => 
                           n474);
   U30002 : XOR2_X1 port map( A1 => n22412, A2 => n22413, Z => n22946);
   U30003 : OAI22_X2 port map( A1 => n7003, A2 => n19599, B1 => n7001, B2 => 
                           n7002, ZN => n29756);
   U30007 : OAI21_X1 port map( A1 => n33767, A2 => n29756, B => n33766, ZN => 
                           n29749);
   U30010 : OR2_X1 port map( A1 => n22287, A2 => n8519, Z => n33549);
   U30011 : INV_X2 port map( I => n33550, ZN => n670);
   U30012 : XOR2_X1 port map( A1 => Plaintext(2), A2 => Key(2), Z => n33550);
   U30013 : NAND2_X1 port map( A1 => n30959, A2 => n28069, ZN => n33552);
   U30015 : INV_X2 port map( I => n33553, ZN => n33957);
   U30018 : OAI22_X2 port map( A1 => n124, A2 => n11004, B1 => n12953, B2 => 
                           n15320, ZN => n24337);
   U30021 : NAND2_X2 port map( A1 => n12206, A2 => n24502, ZN => n25132);
   U30028 : OAI21_X1 port map( A1 => n20147, A2 => n22226, B => n20643, ZN => 
                           n20146);
   U30042 : XOR2_X1 port map( A1 => n26308, A2 => n33566, Z => n11975);
   U30043 : XOR2_X1 port map( A1 => n5690, A2 => n26307, Z => n33566);
   U30046 : XOR2_X1 port map( A1 => n33568, A2 => n21076, Z => n4856);
   U30047 : XOR2_X1 port map( A1 => n29127, A2 => n33569, Z => n33568);
   U30048 : INV_X1 port map( I => n19908, ZN => n33569);
   U30051 : XOR2_X1 port map( A1 => n10549, A2 => n33572, Z => n19341);
   U30052 : XOR2_X1 port map( A1 => n33573, A2 => n10548, Z => n33572);
   U30053 : XNOR2_X1 port map( A1 => n26551, A2 => n26541, ZN => n15819);
   U30060 : NAND2_X2 port map( A1 => n20969, A2 => n7831, ZN => n16542);
   U30061 : NAND3_X1 port map( A1 => n38156, A2 => n29339, A3 => n1391, ZN => 
                           n20480);
   U30065 : NAND2_X2 port map( A1 => n9250, A2 => n9248, ZN => n29678);
   U30073 : XOR2_X1 port map( A1 => n23959, A2 => n17404, Z => n9446);
   U30074 : BUF_X2 port map( I => n12341, Z => n33584);
   U30075 : OAI21_X1 port map( A1 => n18294, A2 => n5166, B => n25725, ZN => 
                           n25726);
   U30077 : NOR2_X2 port map( A1 => n948, A2 => n12844, ZN => n8963);
   U30082 : XOR2_X1 port map( A1 => n23662, A2 => n7129, Z => n7128);
   U30086 : XOR2_X1 port map( A1 => n28988, A2 => n28989, Z => n6835);
   U30090 : INV_X2 port map( I => n27932, ZN => n1072);
   U30091 : XOR2_X1 port map( A1 => n11154, A2 => n11152, Z => n27932);
   U30096 : XOR2_X1 port map( A1 => n33595, A2 => n1938, Z => n1936);
   U30099 : NAND2_X1 port map( A1 => n2488, A2 => n2490, ZN => n2487);
   U30101 : OR2_X1 port map( A1 => n30494, A2 => n30833, Z => n24269);
   U30104 : NAND2_X1 port map( A1 => n10314, A2 => n26852, ZN => n21249);
   U30107 : XOR2_X1 port map( A1 => n26585, A2 => n4622, Z => n10319);
   U30109 : INV_X2 port map( I => n33604, ZN => n8193);
   U30110 : XNOR2_X1 port map( A1 => n11575, A2 => n5600, ZN => n33604);
   U30113 : XOR2_X1 port map( A1 => n3696, A2 => n3695, Z => n8889);
   U30115 : OR2_X1 port map( A1 => n30555, A2 => n38143, Z => n33608);
   U30117 : AOI21_X2 port map( A1 => n33610, A2 => n4665, B => n28309, ZN => 
                           n2269);
   U30118 : OAI21_X1 port map( A1 => n898, A2 => n20577, B => n33612, ZN => 
                           n33611);
   U30120 : XOR2_X1 port map( A1 => n29074, A2 => n33614, Z => n20325);
   U30121 : XOR2_X1 port map( A1 => n29131, A2 => n18430, Z => n33614);
   U30130 : INV_X2 port map( I => n33621, ZN => n4603);
   U30131 : XOR2_X1 port map( A1 => n22516, A2 => n11793, Z => n33622);
   U30134 : NAND2_X1 port map( A1 => n29175, A2 => n18134, ZN => n30089);
   U30137 : INV_X2 port map( I => n33625, ZN => n12478);
   U30138 : XNOR2_X1 port map( A1 => n317, A2 => n9094, ZN => n33625);
   U30141 : NAND2_X2 port map( A1 => n15634, A2 => n33628, ZN => n18062);
   U30142 : NAND3_X2 port map( A1 => n37184, A2 => n25503, A3 => n35611, ZN => 
                           n33628);
   U30144 : NAND3_X1 port map( A1 => n29365, A2 => n12943, A3 => n37096, ZN => 
                           n29370);
   U30145 : INV_X2 port map( I => n17179, ZN => n10140);
   U30149 : XOR2_X1 port map( A1 => n26433, A2 => n8625, Z => n33733);
   U30150 : XOR2_X1 port map( A1 => n21346, A2 => Key(25), Z => n21669);
   U30155 : XOR2_X1 port map( A1 => n16689, A2 => n16687, Z => n22798);
   U30156 : XOR2_X1 port map( A1 => n33777, A2 => n19066, Z => n29456);
   U30158 : XOR2_X1 port map( A1 => n33642, A2 => n9159, Z => n14462);
   U30159 : AOI21_X2 port map( A1 => n33643, A2 => n12167, B => n17383, ZN => 
                           n29659);
   U30161 : XOR2_X1 port map( A1 => n14039, A2 => n19035, Z => n28999);
   U30162 : OR2_X1 port map( A1 => n8479, A2 => n2752, Z => n6137);
   U30163 : INV_X2 port map( I => n25966, ZN => n26030);
   U30164 : NAND2_X2 port map( A1 => n20187, A2 => n20186, ZN => n25966);
   U30167 : NAND2_X2 port map( A1 => n11910, A2 => n17132, ZN => n27326);
   U30168 : NAND2_X2 port map( A1 => n17415, A2 => n17416, ZN => n12327);
   U30170 : XOR2_X1 port map( A1 => n9230, A2 => n12989, Z => n33650);
   U30173 : AOI22_X2 port map( A1 => n30190, A2 => n5414, B1 => n10628, B2 => 
                           n30238, ZN => n33651);
   U30174 : OAI22_X2 port map( A1 => n11213, A2 => n15237, B1 => n12090, B2 => 
                           n13186, ZN => n10931);
   U30179 : NAND3_X2 port map( A1 => n7013, A2 => n7012, A3 => n7014, ZN => 
                           n7712);
   U30181 : XOR2_X1 port map( A1 => n26387, A2 => n10878, Z => n33653);
   U30184 : XOR2_X1 port map( A1 => n22778, A2 => n22687, Z => n22546);
   U30187 : NOR2_X2 port map( A1 => n29488, A2 => n29489, ZN => n29535);
   U30191 : XOR2_X1 port map( A1 => n23966, A2 => n16153, Z => n33659);
   U30192 : XOR2_X1 port map( A1 => n7152, A2 => n7153, Z => n25553);
   U30193 : XOR2_X1 port map( A1 => n26602, A2 => n33661, Z => n33660);
   U30195 : XOR2_X1 port map( A1 => n32885, A2 => n6634, Z => n6633);
   U30196 : AOI22_X1 port map( A1 => n8062, A2 => n33664, B1 => n8064, B2 => 
                           n21147, ZN => n8060);
   U30197 : NAND2_X1 port map( A1 => n19348, A2 => n29756, ZN => n33664);
   U30198 : INV_X2 port map( I => n33665, ZN => n4879);
   U30199 : XOR2_X1 port map( A1 => n5782, A2 => n5781, Z => n33665);
   U30200 : INV_X2 port map( I => n30249, ZN => n30260);
   U30210 : NAND3_X2 port map( A1 => n33671, A2 => n18101, A3 => n17584, ZN => 
                           n24805);
   U30211 : NAND3_X1 port map( A1 => n17586, A2 => n37122, A3 => n19880, ZN => 
                           n33671);
   U30220 : OR2_X1 port map( A1 => n12218, A2 => n15038, Z => n28271);
   U30223 : XOR2_X1 port map( A1 => n28850, A2 => n16017, Z => n29152);
   U30225 : XOR2_X1 port map( A1 => n25271, A2 => n25155, Z => n24948);
   U30229 : NOR2_X1 port map( A1 => n1450, A2 => n15357, ZN => n13053);
   U30234 : XOR2_X1 port map( A1 => n19254, A2 => n22598, Z => n18446);
   U30235 : XOR2_X1 port map( A1 => n15673, A2 => n33687, Z => n15672);
   U30236 : XOR2_X1 port map( A1 => n26590, A2 => n19736, Z => n33687);
   U30237 : XOR2_X1 port map( A1 => n16216, A2 => n7854, Z => n7780);
   U30241 : XOR2_X1 port map( A1 => n15824, A2 => n33694, Z => n33693);
   U30246 : NAND2_X2 port map( A1 => n2766, A2 => n25650, ZN => n18661);
   U30247 : XOR2_X1 port map( A1 => n25011, A2 => n13596, Z => n2896);
   U30248 : OAI22_X2 port map( A1 => n37196, A2 => n36564, B1 => n23351, B2 => 
                           n32158, ZN => n33696);
   U30255 : NAND2_X2 port map( A1 => n19337, A2 => n19395, ZN => n21545);
   U30262 : XOR2_X1 port map( A1 => n26531, A2 => n26341, Z => n26342);
   U30264 : NAND3_X1 port map( A1 => n39425, A2 => n1418, A3 => n37081, ZN => 
                           n12947);
   U30265 : NAND2_X2 port map( A1 => n33760, A2 => n21038, ZN => n29755);
   U30266 : XOR2_X1 port map( A1 => n1456, A2 => n27828, Z => n18662);
   U30269 : MUX2_X1 port map( I0 => n36226, I1 => n378, S => n4604, Z => n15183
                           );
   U30273 : NOR2_X1 port map( A1 => n15880, A2 => n17194, ZN => n33709);
   U30276 : NOR2_X2 port map( A1 => n6977, A2 => n35560, ZN => n10468);
   U30280 : NOR2_X2 port map( A1 => n15981, A2 => n1137, ZN => n2601);
   U30283 : XOR2_X1 port map( A1 => n33716, A2 => n29169, Z => n29897);
   U30284 : NAND2_X2 port map( A1 => n37105, A2 => n12672, ZN => n24728);
   U30285 : XOR2_X1 port map( A1 => n28935, A2 => n33717, Z => n33965);
   U30286 : XOR2_X1 port map( A1 => n28500, A2 => n38195, Z => n33717);
   U30290 : XOR2_X1 port map( A1 => n26194, A2 => n20539, Z => n33718);
   U30292 : XOR2_X1 port map( A1 => n1825, A2 => n11559, Z => n33722);
   U30298 : OAI21_X1 port map( A1 => n35921, A2 => n9942, B => n33731, ZN => 
                           n21443);
   U30300 : XOR2_X1 port map( A1 => n33733, A2 => n8626, Z => n860);
   U30308 : OAI21_X2 port map( A1 => n8175, A2 => n24338, B => n8174, ZN => 
                           n24339);
   U30310 : NAND2_X2 port map( A1 => n33944, A2 => n370, ZN => n33743);
   U30314 : MUX2_X1 port map( I0 => n28555, I1 => n28556, S => n37758, Z => 
                           n28557);
   U30315 : XOR2_X1 port map( A1 => n29130, A2 => n29129, Z => n29135);
   U30316 : XNOR2_X1 port map( A1 => n29121, A2 => n29122, ZN => n29130);
   U30317 : NAND2_X2 port map( A1 => n29600, A2 => n33746, ZN => n29623);
   U30319 : NAND3_X1 port map( A1 => n37213, A2 => n19259, A3 => n26103, ZN => 
                           n26104);
   U30320 : XOR2_X1 port map( A1 => n29147, A2 => n15960, Z => n29086);
   U30321 : XOR2_X1 port map( A1 => n33749, A2 => n33751, Z => n2819);
   U30322 : XOR2_X1 port map( A1 => n12145, A2 => n26417, Z => n5849);
   U30326 : XOR2_X1 port map( A1 => n33750, A2 => n3712, Z => n33749);
   U30327 : INV_X1 port map( I => n24744, ZN => n33754);
   U30328 : XOR2_X1 port map( A1 => n33756, A2 => n22476, Z => n6329);
   U30331 : XOR2_X1 port map( A1 => n12480, A2 => n33757, Z => n12840);
   U30332 : XOR2_X1 port map( A1 => n1621, A2 => n12842, Z => n33757);
   U30333 : XOR2_X1 port map( A1 => n27490, A2 => n1936, Z => n33758);
   U30334 : XOR2_X1 port map( A1 => n33759, A2 => n10070, Z => n11727);
   U30341 : OAI21_X2 port map( A1 => n20330, A2 => n20331, B => n7601, ZN => 
                           n22067);
   U30346 : INV_X1 port map( I => n6732, ZN => n11146);
   U30349 : BUF_X2 port map( I => n18047, Z => n33773);
   U30356 : XOR2_X1 port map( A1 => n5382, A2 => n33776, Z => n855);
   U30357 : XOR2_X1 port map( A1 => n12860, A2 => n12859, Z => n33776);
   U30359 : XOR2_X1 port map( A1 => n12736, A2 => n12735, Z => n12788);
   U30360 : NAND2_X2 port map( A1 => n6036, A2 => n22277, ZN => n22048);
   U30366 : XOR2_X1 port map( A1 => n16650, A2 => n494, Z => n33789);
   U30382 : XOR2_X1 port map( A1 => n23783, A2 => n23938, Z => n8671);
   U30383 : NAND2_X2 port map( A1 => n33799, A2 => n27426, ZN => n13054);
   U30391 : NOR2_X1 port map( A1 => n33561, A2 => n26606, ZN => n33802);
   U30396 : XOR2_X1 port map( A1 => n6741, A2 => n4883, Z => n18209);
   U30398 : XOR2_X1 port map( A1 => n38148, A2 => n5261, Z => n33807);
   U30399 : INV_X2 port map( I => n33808, ZN => n20793);
   U30410 : XOR2_X1 port map( A1 => n727, A2 => n33810, Z => n354);
   U30411 : XOR2_X1 port map( A1 => n8163, A2 => n33811, Z => n33810);
   U30412 : INV_X1 port map( I => n19735, ZN => n33811);
   U30414 : NOR2_X2 port map( A1 => n33813, A2 => n10832, ZN => n6885);
   U30422 : AOI22_X2 port map( A1 => n8928, A2 => n20978, B1 => n23554, B2 => 
                           n35039, ZN => n13617);
   U30425 : INV_X4 port map( I => n18519, ZN => n33826);
   U30429 : XOR2_X1 port map( A1 => n6893, A2 => n20483, Z => n33824);
   U30430 : OAI21_X2 port map( A1 => n19237, A2 => n25557, B => n33825, ZN => 
                           n25777);
   U30439 : XOR2_X1 port map( A1 => n4059, A2 => n4061, Z => n4300);
   U30447 : XOR2_X1 port map( A1 => n18662, A2 => n27832, Z => n33831);
   U30449 : NAND2_X1 port map( A1 => n20743, A2 => n23211, ZN => n33832);
   U30453 : XOR2_X1 port map( A1 => n27552, A2 => n27551, Z => n33837);
   U30454 : XOR2_X1 port map( A1 => n33839, A2 => n36529, Z => n3257);
   U30455 : XOR2_X1 port map( A1 => n3261, A2 => n9184, Z => n33839);
   U30456 : INV_X1 port map( I => n7194, ZN => n30230);
   U30460 : OAI21_X2 port map( A1 => n2294, A2 => n2378, B => n29592, ZN => 
                           n33844);
   U30464 : BUF_X2 port map( I => n7090, Z => n33845);
   U30470 : XOR2_X1 port map( A1 => n14264, A2 => n20454, Z => n9038);
   U30472 : XOR2_X1 port map( A1 => n33848, A2 => n3872, Z => n15754);
   U30475 : XOR2_X1 port map( A1 => n11015, A2 => n11016, Z => n33850);
   U30479 : XOR2_X1 port map( A1 => n13102, A2 => n13101, Z => n33851);
   U30488 : NAND2_X1 port map( A1 => n16693, A2 => n19823, ZN => n19661);
   U30489 : NAND2_X2 port map( A1 => n29870, A2 => n10096, ZN => n29871);
   U30490 : OR2_X1 port map( A1 => n15852, A2 => n36661, Z => n21979);
   U30491 : OAI21_X2 port map( A1 => n19320, A2 => n1813, B => n532, ZN => 
                           n11344);
   U30492 : AOI22_X2 port map( A1 => n26728, A2 => n14380, B1 => n26777, B2 => 
                           n31982, ZN => n33853);
   U30502 : XOR2_X1 port map( A1 => n22594, A2 => n33866, Z => n33865);
   U30505 : XOR2_X1 port map( A1 => n10413, A2 => n3316, Z => n33868);
   U30506 : NAND3_X1 port map( A1 => n1623, A2 => n38535, A3 => n10024, ZN => 
                           n33869);
   U30510 : XOR2_X1 port map( A1 => n27526, A2 => n27473, Z => n33870);
   U30511 : INV_X1 port map( I => n2940, ZN => n25844);
   U30514 : XOR2_X1 port map( A1 => n26399, A2 => n26398, Z => n7689);
   U30520 : NAND2_X2 port map( A1 => n2932, A2 => n30420, ZN => n23996);
   U30523 : INV_X2 port map( I => n31378, ZN => n10618);
   U30526 : INV_X2 port map( I => n33890, ZN => n773);
   U30530 : NAND2_X2 port map( A1 => n14080, A2 => n5960, ZN => n26794);
   U30531 : XOR2_X1 port map( A1 => n14563, A2 => n24950, Z => n3029);
   U30534 : NAND2_X2 port map( A1 => n14822, A2 => n21739, ZN => n7560);
   U30536 : XOR2_X1 port map( A1 => n33906, A2 => n1725, Z => Ciphertext(78));
   U30537 : AOI22_X1 port map( A1 => n17368, A2 => n19318, B1 => n29646, B2 => 
                           n29658, ZN => n33906);
   U30539 : NAND2_X2 port map( A1 => n6208, A2 => n6206, ZN => n6205);
   U30547 : XOR2_X1 port map( A1 => n5246, A2 => n22562, Z => n22419);
   U30548 : OAI22_X1 port map( A1 => n18070, A2 => n1387, B1 => n29228, B2 => 
                           n14933, ZN => n14200);
   U30550 : BUF_X2 port map( I => n16487, Z => n33916);
   U30569 : NAND2_X2 port map( A1 => n25778, A2 => n25776, ZN => n2830);
   U30572 : XOR2_X1 port map( A1 => n11903, A2 => n7573, Z => n26818);
   U30577 : INV_X2 port map( I => n7273, ZN => n24142);
   U30579 : NOR2_X2 port map( A1 => n5015, A2 => n5014, ZN => n9276);
   U30583 : OAI22_X2 port map( A1 => n16411, A2 => n16810, B1 => n16410, B2 => 
                           n16809, ZN => n25962);
   U30585 : CLKBUF_X4 port map( I => n26995, Z => n19364);
   U30588 : XOR2_X1 port map( A1 => n16551, A2 => n16550, Z => n33954);
   U30590 : XOR2_X1 port map( A1 => n13751, A2 => n13749, Z => n33956);
   U30591 : INV_X4 port map( I => n12685, ZN => n18246);
   U30592 : XNOR2_X1 port map( A1 => n8909, A2 => n29083, ZN => n33962);
   U30595 : INV_X2 port map( I => n11896, ZN => n14557);
   U30597 : OR2_X2 port map( A1 => n10097, A2 => n18445, Z => n33966);
   U30598 : AND2_X1 port map( A1 => n29721, A2 => n14337, Z => n33968);
   U30599 : INV_X2 port map( I => n28817, ZN => n28925);
   U3421 : BUF_X2 port map( I => n12519, Z => n3226);
   U15475 : INV_X2 port map( I => n3462, ZN => n8955);
   U9227 : INV_X4 port map( I => n27403, ZN => n1220);
   U3911 : INV_X2 port map( I => n2561, ZN => n9175);
   U5822 : INV_X4 port map( I => n18293, ZN => n917);
   U5706 : INV_X2 port map( I => n24912, ZN => n1273);
   U12087 : OAI21_X2 port map( A1 => n25792, A2 => n25975, B => n17002, ZN => 
                           n25795);
   U1188 : INV_X2 port map( I => n19580, ZN => n25835);
   U6510 : INV_X2 port map( I => n15535, ZN => n968);
   U16873 : INV_X2 port map( I => n3861, ZN => n2944);
   U10138 : NOR2_X2 port map( A1 => n14270, A2 => n4902, ZN => n9392);
   U6809 : INV_X2 port map( I => n26274, ZN => n1509);
   U22777 : INV_X2 port map( I => n11048, ZN => n11890);
   U380 : OAI21_X2 port map( A1 => n27959, A2 => n20185, B => n10721, ZN => 
                           n10720);
   U5871 : NAND2_X2 port map( A1 => n17114, A2 => n33405, ZN => n13500);
   U25694 : INV_X2 port map( I => n13457, ZN => n21223);
   U5048 : NAND2_X2 port map( A1 => n26134, A2 => n25936, ZN => n26024);
   U1221 : AOI21_X2 port map( A1 => n32654, A2 => n10753, B => n20683, ZN => 
                           n11860);
   U7339 : OAI22_X2 port map( A1 => n36764, A2 => n11898, B1 => n2858, B2 => 
                           n5579, ZN => n29860);
   U3258 : NAND2_X2 port map( A1 => n2625, A2 => n17400, ZN => n21040);
   U10896 : INV_X2 port map( I => n11406, ZN => n16252);
   U23384 : INV_X2 port map( I => n19147, ZN => n12167);
   U16469 : NAND2_X2 port map( A1 => n29354, A2 => n12994, ZN => n12993);
   U1098 : INV_X2 port map( I => n17790, ZN => n20864);
   U17113 : INV_X2 port map( I => n16692, ZN => n23071);
   U1040 : OAI21_X2 port map( A1 => n9384, A2 => n4475, B => n1591, ZN => n9382
                           );
   U842 : INV_X4 port map( I => n16836, ZN => n953);
   U16551 : AOI21_X2 port map( A1 => n24392, A2 => n11265, B => n12771, ZN => 
                           n15237);
   U2358 : INV_X2 port map( I => n28692, ZN => n18453);
   U3582 : NAND2_X2 port map( A1 => n15176, A2 => n36442, ZN => n23338);
   U27370 : NAND2_X2 port map( A1 => n18838, A2 => n25108, ZN => n25993);
   U13068 : INV_X2 port map( I => n16524, ZN => n16368);
   U9696 : OAI21_X2 port map( A1 => n24209, A2 => n24207, B => n24208, ZN => 
                           n18938);
   U1938 : INV_X2 port map( I => n13370, ZN => n23578);
   U580 : INV_X2 port map( I => n866, ZN => n26862);
   U5776 : NAND2_X2 port map( A1 => n20403, A2 => n9295, ZN => n9726);
   U15038 : NAND2_X1 port map( A1 => n22807, A2 => n23119, ZN => n31345);
   U1485 : NAND2_X2 port map( A1 => n18715, A2 => n24882, ZN => n25211);
   U27483 : INV_X2 port map( I => n28651, ZN => n28490);
   U763 : NAND2_X2 port map( A1 => n8137, A2 => n27379, ZN => n27300);
   U22306 : INV_X2 port map( I => n37045, ZN => n24184);
   U246 : INV_X2 port map( I => n6932, ZN => n28386);
   U13 : NAND2_X2 port map( A1 => n15773, A2 => n29890, ZN => n29881);
   U1777 : OAI21_X2 port map( A1 => n30900, A2 => n31827, B => n5276, ZN => 
                           n5508);
   U10705 : OAI21_X2 port map( A1 => n9818, A2 => n9817, B => n1056, ZN => 
                           n4916);
   U13467 : NOR2_X2 port map( A1 => n22812, A2 => n22811, ZN => n23587);
   U2155 : INV_X4 port map( I => n5077, ZN => n31940);
   U6320 : BUF_X4 port map( I => n23761, Z => n24300);
   U5290 : NAND2_X2 port map( A1 => n37319, A2 => n37107, ZN => n11796);
   U5569 : INV_X2 port map( I => n26403, ZN => n10491);
   U10669 : AOI21_X2 port map( A1 => n3156, A2 => n3155, B => n3154, ZN => 
                           n3153);
   U2350 : OAI21_X2 port map( A1 => n1997, A2 => n7591, B => n1440, ZN => n7252
                           );
   U349 : INV_X2 port map( I => n6640, ZN => n1069);
   U3916 : BUF_X4 port map( I => n33533, Z => n33178);
   U300 : INV_X2 port map( I => n16067, ZN => n28485);
   U9745 : NAND2_X2 port map( A1 => n24209, A2 => n18937, ZN => n18936);
   U9838 : NAND2_X2 port map( A1 => n3382, A2 => n1629, ZN => n5186);
   U3630 : INV_X2 port map( I => n26779, ZN => n26945);
   U1412 : INV_X2 port map( I => n25569, ZN => n15180);
   U2047 : INV_X2 port map( I => n20679, ZN => n1341);
   U991 : INV_X2 port map( I => n24864, ZN => n1030);
   U2472 : INV_X2 port map( I => n36996, ZN => n23166);
   U732 : INV_X4 port map( I => n16867, ZN => n10062);
   U6294 : AND2_X1 port map( A1 => n35216, A2 => n220, Z => n30400);
   U1386 : INV_X2 port map( I => n34134, ZN => n7075);
   U1825 : BUF_X4 port map( I => n14272, Z => n32190);
   U7190 : OAI21_X2 port map( A1 => n18566, A2 => n21451, B => n18567, ZN => 
                           n21452);
   U14730 : AOI21_X2 port map( A1 => n2300, A2 => n21672, B => n21847, ZN => 
                           n8073);
   U1648 : AOI22_X2 port map( A1 => n18376, A2 => n1520, B1 => n31954, B2 => 
                           n362, ZN => n25837);
   U327 : NAND2_X2 port map( A1 => n28742, A2 => n5424, ZN => n16530);
   U448 : NOR2_X2 port map( A1 => n11375, A2 => n28159, ZN => n28287);
   U131 : NAND2_X2 port map( A1 => n9708, A2 => n30159, ZN => n33362);
   U22212 : NAND2_X2 port map( A1 => n17329, A2 => n17331, ZN => n17458);
   U3138 : OAI21_X2 port map( A1 => n4225, A2 => n32093, B => n35952, ZN => 
                           n2164);
   U1908 : INV_X4 port map( I => n10736, ZN => n946);
   U11661 : OAI21_X2 port map( A1 => n23350, A2 => n37523, B => n30974, ZN => 
                           n23356);
   U12678 : NAND2_X2 port map( A1 => n9578, A2 => n9583, ZN => n15282);
   U30416 : NAND3_X2 port map( A1 => n33816, A2 => n10224, A3 => n33815, ZN => 
                           n9499);
   U4514 : NOR2_X2 port map( A1 => n24649, A2 => n31796, ZN => n4845);
   U3141 : NAND2_X2 port map( A1 => n24648, A2 => n36340, ZN => n24649);
   U6036 : NOR2_X2 port map( A1 => n15149, A2 => n33771, ZN => n15148);
   U2777 : NAND2_X2 port map( A1 => n30024, A2 => n30038, ZN => n30015);
   U5927 : OAI21_X2 port map( A1 => n27946, A2 => n12406, B => n20431, ZN => 
                           n33528);
   U3921 : BUF_X4 port map( I => n16692, Z => n9954);
   U1141 : INV_X2 port map( I => n16296, ZN => n16342);
   U1956 : BUF_X2 port map( I => n8668, Z => n605);
   U81 : OAI21_X2 port map( A1 => n29302, A2 => n29461, B => n38051, ZN => 
                           n21195);
   U17554 : NAND2_X2 port map( A1 => n33190, A2 => n5287, ZN => n31591);
   U3433 : INV_X2 port map( I => n21126, ZN => n18603);
   U3794 : INV_X4 port map( I => n38220, ZN => n7905);
   U12600 : AOI22_X2 port map( A1 => n6229, A2 => n24910, B1 => n12671, B2 => 
                           n24909, ZN => n6228);
   U27338 : INV_X2 port map( I => n18739, ZN => n19091);
   U15360 : INV_X2 port map( I => n3713, ZN => n17556);
   U8386 : NAND2_X2 port map( A1 => n8757, A2 => n33864, ZN => n23360);
   U9389 : AOI21_X2 port map( A1 => n9962, A2 => n9961, B => n1527, ZN => 
                           n16344);
   U5654 : INV_X2 port map( I => n35543, ZN => n20578);
   U1551 : NAND2_X2 port map( A1 => n8139, A2 => n18654, ZN => n30929);
   U14862 : OAI21_X2 port map( A1 => n1823, A2 => n7555, B => n28378, ZN => 
                           n20496);
   U6836 : NOR2_X2 port map( A1 => n3013, A2 => n35855, ZN => n26190);
   U2879 : NAND2_X2 port map( A1 => n28704, A2 => n38220, ZN => n28700);
   U1068 : INV_X2 port map( I => n31917, ZN => n9568);
   U3240 : NAND2_X2 port map( A1 => n32338, A2 => n34559, ZN => n28765);
   U5561 : INV_X4 port map( I => n15575, ZN => n1021);
   U12634 : INV_X2 port map( I => n24724, ZN => n6542);
   U3693 : NOR3_X1 port map( A1 => n33925, A2 => n36422, A3 => n8809, ZN => 
                           n14879);
   U10098 : INV_X4 port map( I => n23142, ZN => n1652);
   U7266 : NOR2_X2 port map( A1 => n5391, A2 => n36912, ZN => n5551);
   U2976 : NAND2_X2 port map( A1 => n16619, A2 => n11120, ZN => n28650);
   U7466 : OAI21_X1 port map( A1 => n28283, A2 => n27980, B => n30565, ZN => 
                           n16543);
   U9288 : NAND2_X1 port map( A1 => n11968, A2 => n30180, ZN => n30185);
   U2099 : INV_X2 port map( I => n22066, ZN => n1673);
   U17989 : OAI21_X2 port map( A1 => n30400, A2 => n31660, B => n38013, ZN => 
                           n31904);
   U16704 : INV_X2 port map( I => n26516, ZN => n19081);
   U18292 : INV_X2 port map( I => n29532, ZN => n29517);
   U2657 : NOR2_X2 port map( A1 => n19546, A2 => n20923, ZN => n4373);
   U2703 : NOR2_X2 port map( A1 => n34114, A2 => n54, ZN => n53);
   U4988 : AOI21_X2 port map( A1 => n502, A2 => n34128, B => n36443, ZN => 
                           n32551);
   U11773 : NAND2_X2 port map( A1 => n37074, A2 => n106, ZN => n9239);
   U7874 : INV_X4 port map( I => n1006, ZN => n3388);
   U574 : INV_X2 port map( I => n10314, ZN => n20660);
   U22525 : NAND3_X2 port map( A1 => n25534, A2 => n25535, A3 => n37795, ZN => 
                           n32911);
   U1814 : INV_X2 port map( I => n33483, ZN => n802);
   U6604 : INV_X2 port map( I => n28376, ZN => n28377);
   U13721 : AOI21_X2 port map( A1 => n9903, A2 => n22238, B => n13632, ZN => 
                           n9838);
   U3196 : NOR2_X2 port map( A1 => n35580, A2 => n26354, ZN => n14521);
   U407 : OAI21_X2 port map( A1 => n19456, A2 => n16127, B => n20561, ZN => 
                           n27061);
   U7168 : BUF_X4 port map( I => n14395, Z => n14396);
   U542 : INV_X2 port map( I => n31682, ZN => n14480);
   U17177 : NAND2_X2 port map( A1 => n38448, A2 => n1049, ZN => n21983);
   U1997 : NAND2_X2 port map( A1 => n23099, A2 => n13650, ZN => n8337);
   U12502 : NAND2_X2 port map( A1 => n2848, A2 => n2847, ZN => n10646);
   U2064 : NAND2_X2 port map( A1 => n12079, A2 => n22131, ZN => n13615);
   U252 : NOR2_X2 port map( A1 => n33424, A2 => n36165, ZN => n14398);
   U435 : NAND2_X2 port map( A1 => n33957, A2 => n10817, ZN => n30959);
   U119 : NOR2_X2 port map( A1 => n39322, A2 => n18667, ZN => n14773);
   U4989 : INV_X2 port map( I => n9987, ZN => n21001);
   U5695 : NAND3_X2 port map( A1 => n18115, A2 => n24161, A3 => n13128, ZN => 
                           n11768);
   U337 : NOR2_X2 port map( A1 => n1190, A2 => n14209, ZN => n2822);
   U3109 : INV_X4 port map( I => n14553, ZN => n1108);
   U3859 : INV_X2 port map( I => n5888, ZN => n355);
   U8441 : INV_X2 port map( I => n18762, ZN => n20620);
   U9367 : OAI21_X1 port map( A1 => n13971, A2 => n26000, B => n2310, ZN => 
                           n13387);
   U5520 : NAND2_X1 port map( A1 => n2311, A2 => n25998, ZN => n2310);
   U24518 : INV_X2 port map( I => n36728, ZN => n21950);
   U14186 : NAND2_X2 port map( A1 => n34485, A2 => n15677, ZN => n21266);
   U21593 : OAI21_X1 port map( A1 => n10345, A2 => n21783, B => n21504, ZN => 
                           n32319);
   U16969 : NAND2_X2 port map( A1 => n4508, A2 => n4506, ZN => n6932);
   U16548 : OAI21_X2 port map( A1 => n14680, A2 => n15449, B => n1018, ZN => 
                           n25707);
   U2158 : OAI21_X2 port map( A1 => n18372, A2 => n35822, B => n6200, ZN => 
                           n6199);
   U12383 : AOI21_X2 port map( A1 => n30366, A2 => n21223, B => n15087, ZN => 
                           n31042);
   U863 : INV_X4 port map( I => n37051, ZN => n1024);
   U3797 : INV_X2 port map( I => n17813, ZN => n22055);
   U1875 : NAND2_X2 port map( A1 => n32260, A2 => n23569, ZN => n23365);
   U21830 : NOR2_X2 port map( A1 => n22330, A2 => n22329, ZN => n22671);
   U4193 : NAND2_X2 port map( A1 => n13044, A2 => n19483, ZN => n439);
   U27166 : NAND2_X1 port map( A1 => n18214, A2 => n1015, ZN => n18213);
   U2427 : INV_X2 port map( I => n13794, ZN => n29384);
   U13970 : BUF_X2 port map( I => n21352, Z => n21683);
   U10685 : AOI21_X2 port map( A1 => n29991, A2 => n29992, B => n29990, ZN => 
                           n9233);
   U26348 : INV_X2 port map( I => n33980, ZN => n28115);
   U10350 : NAND2_X2 port map( A1 => n21920, A2 => n19323, ZN => n7587);
   U5772 : INV_X2 port map( I => n22671, ZN => n1662);
   U23299 : INV_X2 port map( I => n12012, ZN => n20936);
   U1273 : OAI21_X2 port map( A1 => n17930, A2 => n39518, B => n39500, ZN => 
                           n17929);
   U16271 : INV_X2 port map( I => n24637, ZN => n11712);
   U12302 : NAND2_X2 port map( A1 => n17271, A2 => n12500, ZN => n14300);
   U5409 : NOR2_X2 port map( A1 => n33042, A2 => n2731, ZN => n16541);
   U1872 : NAND2_X2 port map( A1 => n1301, A2 => n35915, ZN => n2084);
   U9732 : INV_X4 port map( I => n17810, ZN => n8041);
   U5734 : INV_X2 port map( I => n16271, ZN => n18302);
   U17205 : OR2_X2 port map( A1 => n24280, A2 => n19959, Z => n24284);
   U966 : NOR2_X2 port map( A1 => n13588, A2 => n14065, ZN => n32948);
   U29 : INV_X2 port map( I => n29747, ZN => n29739);
   U9180 : NAND2_X2 port map( A1 => n26965, A2 => n27507, ZN => n11462);
   U1636 : INV_X4 port map( I => n37097, ZN => n20158);
   U4415 : BUF_X4 port map( I => n13543, Z => n13393);
   U582 : INV_X2 port map( I => n26863, ZN => n1089);
   U6091 : AOI21_X2 port map( A1 => n14592, A2 => n39745, B => n17633, ZN => 
                           n6920);
   U7080 : INV_X2 port map( I => n13150, ZN => n13831);
   U9379 : OAI21_X2 port map( A1 => n26190, A2 => n32243, B => n39507, ZN => 
                           n19573);
   U1556 : AOI21_X2 port map( A1 => n25674, A2 => n19589, B => n6592, ZN => 
                           n18058);
   U5999 : INV_X2 port map( I => n19692, ZN => n16104);
   U10329 : OAI21_X2 port map( A1 => n21423, A2 => n21667, B => n21672, ZN => 
                           n21424);
   U978 : NAND2_X1 port map( A1 => n5389, A2 => n24852, ZN => n199);
   U6077 : NAND2_X2 port map( A1 => n13441, A2 => n29586, ZN => n28864);
   U11765 : NAND2_X1 port map( A1 => n3103, A2 => n30983, ZN => n3102);
   U4913 : INV_X2 port map( I => n2008, ZN => n2405);
   U10314 : AOI21_X2 port map( A1 => n13956, A2 => n13044, B => n18496, ZN => 
                           n11174);
   U3027 : BUF_X2 port map( I => n32165, Z => n138);
   U5870 : NAND2_X1 port map( A1 => n28048, A2 => n28260, ZN => n4975);
   U8490 : OAI21_X2 port map( A1 => n1652, A2 => n1313, B => n3906, ZN => n8766
                           );
   U6043 : NAND2_X2 port map( A1 => n9863, A2 => n39495, ZN => n13044);
   U1378 : INV_X4 port map( I => n2576, ZN => n33114);
   U13858 : OAI21_X2 port map( A1 => n21920, A2 => n21621, B => n7587, ZN => 
                           n6800);
   U5593 : NOR2_X2 port map( A1 => n25934, A2 => n38185, ZN => n25800);
   U27627 : NAND2_X2 port map( A1 => n25556, A2 => n1537, ZN => n20236);
   U10365 : AOI22_X2 port map( A1 => n21455, A2 => n21695, B1 => n21454, B2 => 
                           n19395, ZN => n13788);
   U2774 : NAND2_X2 port map( A1 => n22891, A2 => n5838, ZN => n70);
   U5761 : NAND2_X2 port map( A1 => n33745, A2 => n31093, ZN => n17968);
   U10292 : OAI21_X1 port map( A1 => n15436, A2 => n15493, B => n15435, ZN => 
                           n30818);
   U3829 : NAND2_X2 port map( A1 => n21101, A2 => n34001, ZN => n27272);
   U17108 : NOR2_X2 port map( A1 => n22264, A2 => n33738, ZN => n14249);
   U15764 : INV_X2 port map( I => n39680, ZN => n3294);
   U1101 : INV_X2 port map( I => n19341, ZN => n16449);
   U2929 : BUF_X2 port map( I => n4392, Z => n33861);
   U13968 : BUF_X4 port map( I => n21358, Z => n21666);
   U5392 : INV_X2 port map( I => n24713, ZN => n15193);
   U6748 : NOR2_X1 port map( A1 => n26772, A2 => n18225, ZN => n3103);
   U4604 : NAND2_X2 port map( A1 => n10168, A2 => n25751, ZN => n26014);
   U27443 : INV_X2 port map( I => n19016, ZN => n19609);
   U15765 : INV_X1 port map( I => n39680, ZN => n3670);
   U1161 : INV_X2 port map( I => n6302, ZN => n32497);
   U6001 : INV_X1 port map( I => n22925, ZN => n23058);
   U24711 : INV_X2 port map( I => n22137, ZN => n16283);
   U4892 : NAND2_X2 port map( A1 => n18417, A2 => n21712, ZN => n21747);
   U7184 : INV_X2 port map( I => n22491, ZN => n22025);
   U25396 : OAI22_X2 port map( A1 => n2008, A2 => n21924, B1 => n11852, B2 => 
                           n9316, ZN => n4913);
   U19016 : OAI22_X2 port map( A1 => n1156, A2 => n21853, B1 => n1355, B2 => 
                           n21808, ZN => n6271);
   U201 : OAI21_X1 port map( A1 => n32274, A2 => n13508, B => n32273, ZN => 
                           n11536);
   U27174 : INV_X4 port map( I => n23089, ZN => n23169);
   U7996 : NOR2_X2 port map( A1 => n15021, A2 => n25898, ZN => n10475);
   U9771 : INV_X4 port map( I => n24359, ZN => n3685);
   U6834 : NOR2_X2 port map( A1 => n34577, A2 => n26001, ZN => n25898);
   U1178 : OAI21_X2 port map( A1 => n23611, A2 => n4525, B => n4527, ZN => 
                           n4526);
   U26636 : NOR2_X2 port map( A1 => n21266, A2 => n30900, ZN => n16903);
   U7724 : OAI21_X2 port map( A1 => n1442, A2 => n886, B => n5239, ZN => n7945)
                           ;
   U5825 : INV_X4 port map( I => n7982, ZN => n21339);
   U2563 : NOR2_X2 port map( A1 => n13, A2 => n12, ZN => n18454);
   U8083 : NAND2_X2 port map( A1 => n7853, A2 => n38178, ZN => n16373);
   U1489 : AOI21_X2 port map( A1 => n18339, A2 => n20367, B => n21950, ZN => 
                           n18338);
   U1659 : INV_X4 port map( I => n17501, ZN => n17502);
   U5760 : NAND2_X2 port map( A1 => n7494, A2 => n27259, ZN => n8411);
   U10031 : NAND2_X2 port map( A1 => n121, A2 => n33045, ZN => n23024);
   U1621 : OAI21_X2 port map( A1 => n22246, A2 => n33571, B => n37938, ZN => 
                           n22247);
   U11387 : INV_X2 port map( I => n18148, ZN => n24608);
   U719 : INV_X2 port map( I => n2830, ZN => n26101);
   U3742 : INV_X2 port map( I => n36549, ZN => n26866);
   U865 : INV_X2 port map( I => n733, ZN => n25690);
   U13656 : NOR2_X2 port map( A1 => n9838, A2 => n13633, ZN => n13631);
   U1530 : OAI21_X2 port map( A1 => n34040, A2 => n32761, B => n31796, ZN => 
                           n471);
   U3792 : OAI21_X2 port map( A1 => n30475, A2 => n30712, B => n27189, ZN => 
                           n31421);
   U9873 : AOI21_X2 port map( A1 => n10709, A2 => n35963, B => n38894, ZN => 
                           n10708);
   U7390 : AOI22_X2 port map( A1 => n2907, A2 => n30558, B1 => n2909, B2 => 
                           n2910, ZN => n8649);
   U4055 : NOR2_X2 port map( A1 => n6864, A2 => n8892, ZN => n29272);
   U12347 : NAND2_X2 port map( A1 => n11589, A2 => n33268, ZN => n4018);
   U21346 : INV_X4 port map( I => n7536, ZN => n8971);
   U17344 : AOI22_X2 port map( A1 => n22103, A2 => n20234, B1 => n22102, B2 => 
                           n22335, ZN => n22104);
   U18946 : INV_X4 port map( I => n27153, ZN => n5311);
   U12109 : NAND2_X1 port map( A1 => n3837, A2 => n30629, ZN => n11269);
   U6042 : INV_X4 port map( I => n19587, ZN => n5391);
   U13644 : NAND2_X2 port map( A1 => n15347, A2 => n36443, ZN => n2587);
   U19288 : INV_X2 port map( I => n6581, ZN => n19588);
   U17467 : INV_X2 port map( I => n8293, ZN => n21692);
   U5739 : INV_X2 port map( I => n23623, ZN => n23780);
   U3314 : NOR2_X2 port map( A1 => n7485, A2 => n33747, ZN => n23576);
   U7262 : NOR2_X1 port map( A1 => n7962, A2 => n9964, ZN => n5601);
   U4665 : INV_X2 port map( I => n15738, ZN => n20321);
   U336 : NAND2_X2 port map( A1 => n18144, A2 => n11136, ZN => n28180);
   U3963 : OAI21_X2 port map( A1 => n5215, A2 => n5214, B => n36453, ZN => 
                           n9504);
   U2624 : OAI21_X2 port map( A1 => n16395, A2 => n16394, B => n31331, ZN => 
                           n16393);
   U7155 : INV_X4 port map( I => n23107, ZN => n20782);
   U9578 : BUF_X2 port map( I => n25488, Z => n6696);
   U20510 : NOR2_X2 port map( A1 => n18174, A2 => n455, ZN => n14541);
   U6753 : INV_X2 port map( I => n26269, ZN => n26696);
   U10185 : AOI22_X2 port map( A1 => n20374, A2 => n36245, B1 => n20375, B2 => 
                           n1154, ZN => n9125);
   U2071 : NAND2_X2 port map( A1 => n14027, A2 => n36428, ZN => n31458);
   U10170 : OAI21_X2 port map( A1 => n4110, A2 => n1681, B => n6361, ZN => 
                           n4109);
   U3404 : AOI22_X2 port map( A1 => n16484, A2 => n23468, B1 => n21019, B2 => 
                           n32858, ZN => n3194);
   U13961 : OR3_X2 port map( A1 => n19549, A2 => n21870, A3 => n3562, Z => 
                           n17665);
   U1842 : NAND2_X2 port map( A1 => n18478, A2 => n23635, ZN => n3195);
   U8549 : AND2_X2 port map( A1 => n23080, A2 => n10962, Z => n1824);
   U7976 : NAND2_X1 port map( A1 => n8295, A2 => n34417, ZN => n8294);
   U14793 : NAND2_X1 port map( A1 => n9404, A2 => n13880, ZN => n31313);
   U6044 : NAND2_X2 port map( A1 => n21928, A2 => n19372, ZN => n21727);
   U27637 : INV_X2 port map( I => n35290, ZN => n33288);
   U4841 : OR2_X1 port map( A1 => n22035, A2 => n35290, Z => n20388);
   U25129 : INV_X2 port map( I => n23468, ZN => n21019);
   U15832 : INV_X2 port map( I => n30897, ZN => n6839);
   U699 : AOI21_X2 port map( A1 => n8384, A2 => n26807, B => n8382, ZN => n8381
                           );
   U14590 : AOI22_X2 port map( A1 => n21379, A2 => n9102, B1 => n11703, B2 => 
                           n1346, ZN => n5930);
   U15138 : AOI21_X2 port map( A1 => n34016, A2 => n587, B => n2690, ZN => 
                           n21379);
   U5246 : AOI21_X2 port map( A1 => n15462, A2 => n34823, B => n9835, ZN => 
                           n11560);
   U6245 : NAND2_X2 port map( A1 => n5519, A2 => n14436, ZN => n5672);
   U408 : AOI21_X2 port map( A1 => n34387, A2 => n8642, B => n1474, ZN => n8641
                           );
   U16972 : INV_X2 port map( I => n19891, ZN => n28131);
   U8655 : INV_X2 port map( I => n22497, ZN => n1154);
   U534 : NAND2_X2 port map( A1 => n26708, A2 => n17034, ZN => n15825);
   U2723 : BUF_X4 port map( I => n27392, Z => n14881);
   U3439 : NAND2_X2 port map( A1 => n7512, A2 => n33879, ZN => n25799);
   U13689 : NAND2_X2 port map( A1 => n7578, A2 => n22296, ZN => n11144);
   U409 : NAND2_X2 port map( A1 => n5239, A2 => n5352, ZN => n7719);
   U13056 : INV_X1 port map( I => n12973, ZN => n4563);
   U1577 : OAI21_X2 port map( A1 => n933, A2 => n1271, B => n13221, ZN => 
                           n13220);
   U6151 : NOR2_X2 port map( A1 => n34360, A2 => n37075, ZN => n8383);
   U5834 : INV_X2 port map( I => n29720, ZN => n29708);
   U10399 : BUF_X2 port map( I => n21937, Z => n19375);
   U17659 : NOR2_X2 port map( A1 => n3158, A2 => n3159, ZN => n33292);
   U1847 : NAND2_X2 port map( A1 => n23334, A2 => n23635, ZN => n32573);
   U8267 : NAND2_X1 port map( A1 => n12809, A2 => n12808, ZN => n31094);
   U10162 : AOI21_X2 port map( A1 => n14622, A2 => n22229, B => n22230, ZN => 
                           n20551);
   U3346 : OAI21_X1 port map( A1 => n14100, A2 => n25727, B => n19678, ZN => 
                           n17740);
   U836 : INV_X2 port map( I => n37048, ZN => n25337);
   U12666 : AOI21_X2 port map( A1 => n18468, A2 => n15333, B => n19630, ZN => 
                           n7610);
   U22344 : NOR3_X2 port map( A1 => n32938, A2 => n32937, A3 => n34044, ZN => 
                           n32483);
   U15178 : AOI21_X2 port map( A1 => n12407, A2 => n16547, B => n2730, ZN => 
                           n3253);
   U1977 : NAND2_X2 port map( A1 => n14343, A2 => n14188, ZN => n19168);
   U4855 : AOI22_X2 port map( A1 => n21637, A2 => n21636, B1 => n21942, B2 => 
                           n19133, ZN => n33389);
   U20145 : INV_X2 port map( I => n24733, ZN => n24841);
   U1505 : INV_X2 port map( I => n16897, ZN => n33400);
   U2799 : INV_X2 port map( I => n7225, ZN => n15122);
   U10686 : NOR2_X1 port map( A1 => n7363, A2 => n6372, ZN => n10943);
   U11710 : INV_X1 port map( I => n19203, ZN => n1471);
   U16708 : OAI21_X2 port map( A1 => n18063, A2 => n24862, B => n31684, ZN => 
                           n4227);
   U11109 : NOR2_X1 port map( A1 => n24424, A2 => n7658, ZN => n7657);
   U28579 : AOI22_X2 port map( A1 => n33196, A2 => n20782, B1 => n22982, B2 => 
                           n23111, ZN => n22983);
   U2460 : INV_X2 port map( I => n6314, ZN => n16580);
   U16437 : INV_X4 port map( I => n26837, ZN => n20211);
   U30293 : NAND3_X2 port map( A1 => n33724, A2 => n19591, A3 => n32014, ZN => 
                           n16473);
   U17082 : OAI22_X2 port map( A1 => n2746, A2 => n37202, B1 => n16541, B2 => 
                           n2745, ZN => n16539);
   U1046 : NOR2_X2 port map( A1 => n3228, A2 => n3227, ZN => n10798);
   U6464 : CLKBUF_X2 port map( I => Key(164), Z => n29363);
   U6439 : INV_X2 port map( I => n10212, ZN => n10211);
   U4632 : INV_X4 port map( I => n11710, ZN => n19630);
   U16536 : NAND2_X2 port map( A1 => n20634, A2 => n26219, ZN => n13156);
   U1458 : AOI21_X2 port map( A1 => n21936, A2 => n21935, B => n21934, ZN => 
                           n22130);
   U26980 : INV_X4 port map( I => n23567, ZN => n15981);
   U11225 : NAND3_X2 port map( A1 => n17647, A2 => n13955, A3 => n28276, ZN => 
                           n11005);
   U6956 : OAI21_X2 port map( A1 => n30528, A2 => n1490, B => n26670, ZN => 
                           n18879);
   U6957 : AOI22_X2 port map( A1 => n19331, A2 => n26972, B1 => n32427, B2 => 
                           n5935, ZN => n30528);
   U12225 : AOI21_X2 port map( A1 => n15355, A2 => n8907, B => n8905, ZN => 
                           n16879);
   U8543 : INV_X1 port map( I => n8943, ZN => n15911);
   U3839 : AOI22_X2 port map( A1 => n5555, A2 => n12952, B1 => n23035, B2 => 
                           n7575, ZN => n4972);
   U2581 : NOR2_X2 port map( A1 => n26014, A2 => n26013, ZN => n7517);
   U249 : INV_X2 port map( I => n16303, ZN => n28756);
   U6498 : INV_X1 port map( I => n12952, ZN => n14402);
   U2338 : INV_X4 port map( I => n29595, ZN => n31667);
   U9821 : CLKBUF_X4 port map( I => n24318, Z => n19566);
   U5069 : INV_X2 port map( I => n27884, ZN => n28256);
   U24679 : OAI21_X2 port map( A1 => n13081, A2 => n1437, B => n28274, ZN => 
                           n17647);
   U7588 : INV_X2 port map( I => n28659, ZN => n28427);
   U8366 : NAND2_X2 port map( A1 => n2087, A2 => n9011, ZN => n2086);
   U965 : INV_X2 port map( I => n37235, ZN => n6606);
   U25997 : NAND2_X2 port map( A1 => n31595, A2 => n36166, ZN => n30058);
   U1038 : OAI21_X2 port map( A1 => n12984, A2 => n25989, B => n30571, ZN => 
                           n11423);
   U17505 : INV_X4 port map( I => n29885, ZN => n15773);
   U3676 : NOR2_X2 port map( A1 => n17013, A2 => n25410, ZN => n9788);
   U21744 : INV_X2 port map( I => n3120, ZN => n24592);
   U18479 : AOI21_X2 port map( A1 => n23470, A2 => n1292, B => n1310, ZN => 
                           n15564);
   U16639 : NAND2_X2 port map( A1 => n27370, A2 => n27369, ZN => n32332);
   U11586 : AOI21_X2 port map( A1 => n27366, A2 => n27364, B => n16482, ZN => 
                           n27370);
   U2964 : INV_X4 port map( I => n12430, ZN => n29260);
   U4361 : NAND2_X2 port map( A1 => n26822, A2 => n26823, ZN => n4098);
   U16237 : NAND2_X1 port map( A1 => n3723, A2 => n39418, ZN => n3722);
   U12614 : NAND2_X1 port map( A1 => n7806, A2 => n5167, ZN => n7805);
   U874 : INV_X2 port map( I => n18966, ZN => n25487);
   U7072 : AOI21_X2 port map( A1 => n23493, A2 => n35130, B => n23315, ZN => 
                           n14129);
   U29965 : OAI22_X2 port map( A1 => n5597, A2 => n25517, B1 => n5596, B2 => 
                           n25620, ZN => n33535);
   U15045 : INV_X4 port map( I => n2597, ZN => n10220);
   U5824 : BUF_X2 port map( I => n21927, Z => n19372);
   U10279 : BUF_X4 port map( I => n18711, Z => n9265);
   U15546 : OAI21_X2 port map( A1 => n3377, A2 => n29793, B => n36096, ZN => 
                           n9456);
   U24755 : NAND2_X2 port map( A1 => n1354, A2 => n18028, ZN => n18026);
   U5601 : NOR2_X2 port map( A1 => n33995, A2 => n39020, ZN => n3389);
   U13431 : NAND2_X2 port map( A1 => n8337, A2 => n11582, ZN => n18499);
   U22608 : OAI21_X2 port map( A1 => n18193, A2 => n2348, B => n10747, ZN => 
                           n24341);
   U4384 : INV_X4 port map( I => n20404, ZN => n1593);
   U9425 : NAND2_X2 port map( A1 => n2625, A2 => n6056, ZN => n7292);
   U3164 : INV_X2 port map( I => n4209, ZN => n22757);
   U18075 : INV_X2 port map( I => n18467, ZN => n6604);
   U14091 : NAND2_X1 port map( A1 => n17323, A2 => n1002, ZN => n20575);
   U1213 : INV_X2 port map( I => n6263, ZN => n23552);
   U3303 : NAND2_X2 port map( A1 => n17989, A2 => n22310, ZN => n22051);
   U4619 : BUF_X2 port map( I => n24694, Z => n32398);
   U10103 : BUF_X2 port map( I => n23202, Z => n2350);
   U12942 : INV_X4 port map( I => n35960, ZN => n20411);
   U5321 : OAI21_X2 port map( A1 => n7949, A2 => n24119, B => n232, ZN => n5853
                           );
   U647 : INV_X2 port map( I => n38149, ZN => n26568);
   U1788 : INV_X4 port map( I => n24432, ZN => n1608);
   U21795 : NAND2_X1 port map( A1 => n14876, A2 => n22804, ZN => n14875);
   U790 : INV_X4 port map( I => n17029, ZN => n19095);
   U710 : NAND2_X2 port map( A1 => n9633, A2 => n27253, ZN => n31716);
   U5718 : NAND2_X2 port map( A1 => n12360, A2 => n13555, ZN => n24098);
   U12644 : OAI21_X1 port map( A1 => n957, A2 => n31845, B => n10403, ZN => 
                           n23858);
   U1440 : INV_X2 port map( I => n2696, ZN => n18360);
   U24648 : INV_X1 port map( I => n26740, ZN => n17786);
   U5899 : INV_X2 port map( I => n15371, ZN => n1489);
   U3300 : BUF_X2 port map( I => n27919, Z => n28079);
   U8666 : OAI21_X2 port map( A1 => n6381, A2 => n21766, B => n9759, ZN => 
                           n5006);
   U2579 : NAND2_X2 port map( A1 => n31038, A2 => n18809, ZN => n6075);
   U3642 : OAI22_X2 port map( A1 => n2451, A2 => n37289, B1 => n10479, B2 => 
                           n12373, ZN => n31038);
   U12240 : INV_X2 port map( I => n19240, ZN => n1522);
   U9919 : NAND2_X2 port map( A1 => n14845, A2 => n35192, ZN => n17521);
   U1109 : INV_X2 port map( I => n94, ZN => n24235);
   U8246 : NAND2_X1 port map( A1 => n11609, A2 => n5224, ZN => n5223);
   U23573 : AOI21_X2 port map( A1 => n13626, A2 => n34920, B => n12628, ZN => 
                           n13571);
   U4950 : INV_X1 port map( I => n4472, ZN => n1312);
   U6022 : NOR2_X2 port map( A1 => n22196, A2 => n38976, ZN => n22286);
   U2239 : INV_X1 port map( I => n14784, ZN => n6960);
   U7179 : INV_X2 port map( I => n14381, ZN => n1046);
   U7738 : INV_X2 port map( I => n5350, ZN => n5352);
   U10250 : NAND2_X2 port map( A1 => n18360, A2 => n36006, ZN => n5693);
   U2833 : BUF_X2 port map( I => n26795, Z => n106);
   U2337 : AOI21_X2 port map( A1 => n9688, A2 => n32352, B => n17085, ZN => 
                           n3945);
   U3593 : AOI21_X2 port map( A1 => n5908, A2 => n35059, B => n26039, ZN => 
                           n9882);
   U8454 : AOI21_X2 port map( A1 => n4890, A2 => n22905, B => n23045, ZN => 
                           n22906);
   U9710 : NAND2_X1 port map( A1 => n24132, A2 => n39309, ZN => n17259);
   U5365 : INV_X1 port map( I => n20891, ZN => n26786);
   U10778 : OAI21_X2 port map( A1 => n11410, A2 => n11409, B => n17225, ZN => 
                           n13134);
   U3306 : BUF_X4 port map( I => n13904, Z => n13555);
   U2127 : AOI22_X2 port map( A1 => n1340, A2 => n32478, B1 => n4200, B2 => 
                           n17499, ZN => n7107);
   U4362 : NAND2_X2 port map( A1 => n12162, A2 => n18519, ZN => n13218);
   U7774 : OAI21_X2 port map( A1 => n27115, A2 => n19334, B => n9633, ZN => 
                           n12744);
   U18780 : NOR2_X2 port map( A1 => n9347, A2 => n9349, ZN => n9344);
   U22282 : INV_X4 port map( I => n36422, ZN => n14994);
   U23214 : INV_X4 port map( I => n11823, ZN => n16576);
   U12591 : OAI21_X2 port map( A1 => n12518, A2 => n37421, B => n9826, ZN => 
                           n24438);
   U11544 : INV_X2 port map( I => n27570, ZN => n1468);
   U25460 : INV_X2 port map( I => n2348, ZN => n24326);
   U4226 : NAND2_X1 port map( A1 => n30991, A2 => n7409, ZN => n27967);
   U23288 : INV_X2 port map( I => n32776, ZN => n17580);
   U12662 : OAI21_X2 port map( A1 => n18744, A2 => n35049, B => n19643, ZN => 
                           n15554);
   U4292 : INV_X4 port map( I => n28114, ZN => n28249);
   U6407 : BUF_X2 port map( I => n33678, Z => n2458);
   U10041 : AOI21_X2 port map( A1 => n3119, A2 => n23110, B => n33196, ZN => 
                           n12121);
   U27912 : INV_X2 port map( I => n34013, ZN => n23174);
   U5777 : INV_X2 port map( I => n32135, ZN => n18568);
   U2981 : NOR2_X2 port map( A1 => n27081, A2 => n35750, ZN => n27163);
   U1177 : AOI21_X2 port map( A1 => n23748, A2 => n13752, B => n10763, ZN => 
                           n6911);
   U17298 : NOR2_X2 port map( A1 => n29426, A2 => n29454, ZN => n29482);
   U7144 : OAI22_X2 port map( A1 => n12123, A2 => n19697, B1 => n1142, B2 => 
                           n20230, ZN => n12122);
   U2537 : OAI22_X2 port map( A1 => n28525, A2 => n28736, B1 => n8050, B2 => 
                           n28735, ZN => n19354);
   U10095 : INV_X2 port map( I => n22921, ZN => n5838);
   U5024 : NAND2_X2 port map( A1 => n9321, A2 => n23548, ZN => n23229);
   U26974 : INV_X2 port map( I => n39830, ZN => n29704);
   U22555 : NAND4_X2 port map( A1 => n11065, A2 => n11064, A3 => n17331, A4 => 
                           n17329, ZN => n25959);
   U25909 : INV_X2 port map( I => n33029, ZN => n33952);
   U4797 : NAND2_X1 port map( A1 => n20790, A2 => n35282, ZN => n583);
   U18711 : BUF_X4 port map( I => n15426, Z => n31796);
   U1947 : AOI21_X2 port map( A1 => n35689, A2 => n30506, B => n21130, ZN => 
                           n15940);
   U25817 : NAND2_X2 port map( A1 => n22344, A2 => n15350, ZN => n21984);
   U1306 : AOI21_X2 port map( A1 => n33826, A2 => n25557, B => n19367, ZN => 
                           n33825);
   U3186 : INV_X4 port map( I => n21822, ZN => n18174);
   U12014 : INV_X2 port map( I => n31791, ZN => n1879);
   U13139 : OAI22_X2 port map( A1 => n5759, A2 => n23017, B1 => n8692, B2 => 
                           n9078, ZN => n23019);
   U21871 : NAND2_X2 port map( A1 => n11144, A2 => n22248, ZN => n11143);
   U11568 : BUF_X2 port map( I => n7611, Z => n4964);
   U3599 : AND2_X1 port map( A1 => n27385, A2 => n18549, Z => n5220);
   U30384 : INV_X4 port map( I => n9876, ZN => n22344);
   U18791 : INV_X1 port map( I => n17464, ZN => n18679);
   U17549 : INV_X2 port map( I => n17775, ZN => n32441);
   U5850 : INV_X2 port map( I => n16116, ZN => n29494);
   U2595 : OAI22_X2 port map( A1 => n5669, A2 => n33081, B1 => n32777, B2 => 
                           n31788, ZN => n30239);
   U16617 : OAI22_X2 port map( A1 => n6720, A2 => n15773, B1 => n967, B2 => 
                           n38217, ZN => n29889);
   U44 : NOR2_X2 port map( A1 => n33813, A2 => n10832, ZN => n31533);
   U28432 : AOI21_X2 port map( A1 => n22345, A2 => n22344, B => n22343, ZN => 
                           n22346);
   U21082 : INV_X2 port map( I => n8544, ZN => n9677);
   U8721 : INV_X2 port map( I => n21872, ZN => n21695);
   U5043 : INV_X2 port map( I => n10705, ZN => n22541);
   U25106 : NOR2_X2 port map( A1 => n36227, A2 => n35685, ZN => n16027);
   U6444 : INV_X2 port map( I => n21740, ZN => n21748);
   U8434 : INV_X4 port map( I => n31931, ZN => n1301);
   U2183 : OR2_X1 port map( A1 => n21822, A2 => n19016, Z => n21678);
   U16378 : INV_X4 port map( I => n31511, ZN => n29587);
   U13050 : INV_X2 port map( I => n24318, ZN => n18348);
   U26149 : NAND2_X2 port map( A1 => n27959, A2 => n37671, ZN => n18036);
   U6149 : NOR2_X2 port map( A1 => n38900, A2 => n37075, ZN => n27560);
   U2032 : AOI21_X2 port map( A1 => n24390, A2 => n14292, B => n14291, ZN => 
                           n16068);
   U10255 : INV_X2 port map( I => n22223, ZN => n22165);
   U24504 : NAND2_X1 port map( A1 => n9670, A2 => n21576, ZN => n20588);
   U26286 : AOI21_X2 port map( A1 => n30306, A2 => n17685, B => n22067, ZN => 
                           n22068);
   U651 : NAND3_X2 port map( A1 => n36528, A2 => n27244, A3 => n991, ZN => 
                           n30678);
   U4578 : INV_X2 port map( I => n1326, ZN => n8679);
   U12763 : INV_X2 port map( I => n19294, ZN => n24811);
   U22330 : AOI21_X2 port map( A1 => n937, A2 => n10242, B => n17723, ZN => 
                           n22127);
   U9744 : OAI21_X2 port map( A1 => n24251, A2 => n24466, B => n33379, ZN => 
                           n13264);
   U30004 : AOI21_X2 port map( A1 => n21482, A2 => n21483, B => n5751, ZN => 
                           n14125);
   U1414 : NAND2_X2 port map( A1 => n7916, A2 => n22239, ZN => n9903);
   U2478 : INV_X4 port map( I => n34016, ZN => n5751);
   U10429 : CLKBUF_X4 port map( I => n21933, Z => n20003);
   U12459 : INV_X2 port map( I => n18909, ZN => n6894);
   U3509 : INV_X2 port map( I => n3014, ZN => n1416);
   U4984 : INV_X2 port map( I => n22239, ZN => n3181);
   U6430 : INV_X4 port map( I => n20266, ZN => n1349);
   U8036 : OAI21_X2 port map( A1 => n1521, A2 => n11033, B => n7258, ZN => 
                           n7260);
   U3988 : NAND2_X2 port map( A1 => n4536, A2 => n36720, ZN => n31446);
   U2466 : BUF_X2 port map( I => n29641, Z => n6181);
   U23304 : OAI21_X2 port map( A1 => n4600, A2 => n35525, B => n12027, ZN => 
                           n18123);
   U28817 : OAI21_X2 port map( A1 => n33379, A2 => n19566, B => n24467, ZN => 
                           n24253);
   U244 : INV_X4 port map( I => n18875, ZN => n1431);
   U12820 : NAND2_X1 port map( A1 => n18532, A2 => n12146, ZN => n2091);
   U19566 : INV_X4 port map( I => n12289, ZN => n23533);
   U19162 : INV_X2 port map( I => n29937, ZN => n16060);
   U26468 : INV_X2 port map( I => n19982, ZN => n16544);
   U8365 : OAI22_X2 port map( A1 => n1953, A2 => n2601, B1 => n31829, B2 => 
                           n1298, ZN => n1951);
   U11716 : AOI22_X2 port map( A1 => n10891, A2 => n10890, B1 => n7912, B2 => 
                           n35580, ZN => n8506);
   U16624 : INV_X2 port map( I => n16186, ZN => n4914);
   U3204 : INV_X1 port map( I => n25367, ZN => n15791);
   U8467 : AOI22_X2 port map( A1 => n22803, A2 => n12029, B1 => n10552, B2 => 
                           n1646, ZN => n10551);
   U1430 : NAND2_X2 port map( A1 => n2257, A2 => n6347, ZN => n5894);
   U1170 : NAND3_X2 port map( A1 => n6514, A2 => n36630, A3 => n4147, ZN => 
                           n22971);
   U975 : NAND2_X1 port map( A1 => n5387, A2 => n24853, ZN => n198);
   U5026 : AOI21_X2 port map( A1 => n17638, A2 => n22187, B => n39607, ZN => 
                           n17637);
   U6547 : NAND2_X2 port map( A1 => n29937, A2 => n30049, ZN => n2160);
   U7270 : CLKBUF_X4 port map( I => n21441, Z => n21840);
   U24420 : OAI21_X2 port map( A1 => n18253, A2 => n22322, B => n22323, ZN => 
                           n17970);
   U11788 : OAI21_X2 port map( A1 => n20103, A2 => n18773, B => n26734, ZN => 
                           n21008);
   U21247 : INV_X4 port map( I => n15248, ZN => n15389);
   U341 : NOR2_X2 port map( A1 => n6115, A2 => n6114, ZN => n30993);
   U10409 : INV_X1 port map( I => n21933, ZN => n15696);
   U8040 : NAND2_X2 port map( A1 => n29080, A2 => n1822, ZN => n1821);
   U18098 : NAND2_X1 port map( A1 => n20419, A2 => n35115, ZN => n27333);
   U16311 : INV_X2 port map( I => n22765, ZN => n19014);
   U2993 : NAND2_X2 port map( A1 => n28115, A2 => n28246, ZN => n21238);
   U10502 : OAI21_X1 port map( A1 => n39656, A2 => n3562, B => n31035, ZN => 
                           n30824);
   U1689 : INV_X2 port map( I => n27895, ZN => n981);
   U1663 : NOR2_X1 port map( A1 => n815, A2 => n10089, ZN => n8106);
   U1230 : NAND2_X2 port map( A1 => n23533, A2 => n23535, ZN => n5184);
   U10268 : INV_X2 port map( I => n22196, ZN => n1327);
   U12075 : NAND2_X2 port map( A1 => n9378, A2 => n7135, ZN => n9377);
   U14142 : NAND2_X2 port map( A1 => n31206, A2 => n14239, ZN => n8659);
   U25138 : INV_X2 port map( I => n23955, ZN => n21030);
   U27678 : NAND2_X2 port map( A1 => n30396, A2 => n29871, ZN => n33297);
   U12917 : AOI21_X2 port map( A1 => n15899, A2 => n15968, B => n13555, ZN => 
                           n15898);
   U26448 : INV_X4 port map( I => n21137, ZN => n28193);
   U5259 : INV_X2 port map( I => n24076, ZN => n24075);
   U1693 : OAI21_X2 port map( A1 => n37733, A2 => n5572, B => n32507, ZN => 
                           n2464);
   U4551 : BUF_X2 port map( I => n25553, Z => n19581);
   U7463 : OAI22_X1 port map( A1 => n3372, A2 => n12350, B1 => n3897, B2 => 
                           n3898, ZN => n33192);
   U3823 : INV_X2 port map( I => n13728, ZN => n7536);
   U20477 : INV_X2 port map( I => n22135, ZN => n8017);
   U9741 : OAI21_X2 port map( A1 => n35300, A2 => n24373, B => n33937, ZN => 
                           n12579);
   U20083 : NOR2_X2 port map( A1 => n19530, A2 => n23085, ZN => n19281);
   U4183 : NOR2_X1 port map( A1 => n7615, A2 => n28442, ZN => n33829);
   U17937 : INV_X2 port map( I => n19496, ZN => n21587);
   U12617 : OAI21_X2 port map( A1 => n1268, A2 => n20155, B => n24712, ZN => 
                           n1907);
   U13267 : OAI21_X2 port map( A1 => n19119, A2 => n23281, B => n1291, ZN => 
                           n17443);
   U5174 : INV_X2 port map( I => n37218, ZN => n23034);
   U1933 : INV_X2 port map( I => n23502, ZN => n1294);
   U3835 : NOR2_X2 port map( A1 => n24707, A2 => n34526, ZN => n32477);
   U2819 : NAND3_X2 port map( A1 => n25988, A2 => n25990, A3 => n38548, ZN => 
                           n25766);
   U20728 : OR3_X1 port map( A1 => n35586, A2 => n22996, A3 => n3310, Z => 
                           n32159);
   U14044 : BUF_X2 port map( I => Key(156), Z => n19904);
   U3002 : OAI21_X2 port map( A1 => n12392, A2 => n23111, B => n23108, ZN => 
                           n18527);
   U4790 : BUF_X4 port map( I => n19938, Z => n15330);
   U6251 : INV_X2 port map( I => n32026, ZN => n25545);
   U945 : INV_X2 port map( I => n12159, ZN => n1843);
   U23778 : INV_X2 port map( I => n37084, ZN => n14601);
   U17359 : AOI21_X1 port map( A1 => n10846, A2 => n17885, B => n10845, ZN => 
                           n4739);
   U1757 : AOI22_X2 port map( A1 => n12579, A2 => n24118, B1 => n12580, B2 => 
                           n14478, ZN => n5139);
   U11587 : NAND2_X2 port map( A1 => n27587, A2 => n12074, ZN => n27039);
   U1684 : OAI22_X2 port map( A1 => n21080, A2 => n9547, B1 => n21081, B2 => 
                           n18329, ZN => n23908);
   U17040 : INV_X2 port map( I => n21152, ZN => n10736);
   U6986 : INV_X2 port map( I => n24529, ZN => n24710);
   U6707 : NOR2_X2 port map( A1 => n9201, A2 => n13471, ZN => n27319);
   U21641 : AOI22_X2 port map( A1 => n11687, A2 => n34452, B1 => n33623, B2 => 
                           n13899, ZN => n32337);
   U4707 : INV_X1 port map( I => n23944, ZN => n30849);
   U10309 : AOI21_X2 port map( A1 => n587, A2 => n13472, B => n21565, ZN => 
                           n3270);
   U29789 : INV_X2 port map( I => n29456, ZN => n29377);
   U1102 : INV_X4 port map( I => n626, ZN => n11673);
   U7491 : INV_X4 port map( I => n1962, ZN => n29776);
   U13988 : INV_X4 port map( I => n14424, ZN => n21787);
   U16397 : OAI21_X2 port map( A1 => n38537, A2 => n28570, B => n979, ZN => 
                           n33663);
   U10713 : NOR2_X2 port map( A1 => n16392, A2 => n16391, ZN => n16390);
   U3242 : BUF_X4 port map( I => n10820, Z => n196);
   U1062 : NAND2_X2 port map( A1 => n26118, A2 => n1098, ZN => n33485);
   U13564 : BUF_X2 port map( I => n22853, Z => n22995);
   U2843 : INV_X2 port map( I => n9668, ZN => n30716);
   U4659 : NAND2_X1 port map( A1 => n24380, A2 => n32937, ZN => n4178);
   U12629 : OAI21_X2 port map( A1 => n35968, A2 => n35088, B => n4176, ZN => 
                           n17961);
   U13357 : NOR2_X2 port map( A1 => n15373, A2 => n20076, ZN => n7011);
   U6940 : AOI22_X1 port map( A1 => n20030, A2 => n7445, B1 => n24794, B2 => 
                           n20029, ZN => n20028);
   U23583 : INV_X2 port map( I => n17412, ZN => n30240);
   U7727 : INV_X1 port map( I => n19667, ZN => n28138);
   U29551 : INV_X4 port map( I => n39020, ZN => n979);
   U2818 : INV_X2 port map( I => n20830, ZN => n29378);
   U2305 : INV_X1 port map( I => n21445, ZN => n21844);
   U25212 : NOR2_X2 port map( A1 => n26118, A2 => n1098, ZN => n20061);
   U12287 : NOR2_X2 port map( A1 => n25506, A2 => n15635, ZN => n15634);
   U16759 : NAND2_X2 port map( A1 => n37544, A2 => n18667, ZN => n11634);
   U4030 : OAI21_X2 port map( A1 => n21954, A2 => n30996, B => n22190, ZN => 
                           n21956);
   U1867 : OAI21_X2 port map( A1 => n25456, A2 => n25455, B => n10674, ZN => 
                           n25458);
   U28118 : NOR2_X2 port map( A1 => n1117, A2 => n25379, ZN => n25455);
   U1745 : INV_X1 port map( I => n9520, ZN => n18329);
   U14621 : NAND2_X1 port map( A1 => n29911, A2 => n7457, ZN => n29931);
   U5896 : BUF_X2 port map( I => n20896, Z => n31832);
   U18046 : INV_X1 port map( I => n5078, ZN => n9899);
   U5659 : NAND2_X2 port map( A1 => n26743, A2 => n11679, ZN => n30722);
   U22131 : NOR2_X1 port map( A1 => n23425, A2 => n10633, ZN => n13579);
   U5558 : INV_X2 port map( I => n11834, ZN => n25995);
   U24808 : NOR2_X2 port map( A1 => n22833, A2 => n22937, ZN => n15555);
   U8779 : BUF_X2 port map( I => Key(93), Z => n19804);
   U15457 : AOI21_X1 port map( A1 => n22088, A2 => n31407, B => n3002, ZN => 
                           n22090);
   U8576 : NOR2_X2 port map( A1 => n8749, A2 => n8679, ZN => n22402);
   U8602 : BUF_X4 port map( I => n10463, Z => n8749);
   U8565 : NAND2_X2 port map( A1 => n21984, A2 => n20238, ZN => n21985);
   U8339 : NOR2_X2 port map( A1 => n3869, A2 => n24477, ZN => n24234);
   U7474 : INV_X2 port map( I => n775, ZN => n1058);
   U13762 : NOR2_X2 port map( A1 => n4283, A2 => n6036, ZN => n9904);
   U6615 : AND2_X1 port map( A1 => n27066, A2 => n1000, Z => n30485);
   U12540 : OAI21_X1 port map( A1 => n24814, A2 => n9277, B => n11121, ZN => 
                           n12832);
   U21094 : INV_X1 port map( I => n3433, ZN => n32232);
   U12772 : OAI22_X2 port map( A1 => n11760, A2 => n7344, B1 => n17947, B2 => 
                           n14705, ZN => n11759);
   U5847 : INV_X2 port map( I => n16252, ZN => n29422);
   U4847 : BUF_X2 port map( I => n32675, Z => n32318);
   U20691 : NOR2_X2 port map( A1 => n8070, A2 => n7986, ZN => n7987);
   U6116 : INV_X2 port map( I => n28473, ZN => n9586);
   U9708 : AOI21_X2 port map( A1 => n24332, A2 => n24336, B => n19382, ZN => 
                           n6955);
   U4229 : NAND2_X1 port map( A1 => n8370, A2 => n8819, ZN => n31781);
   U18414 : AOI21_X1 port map( A1 => n5711, A2 => n5541, B => n5710, ZN => 
                           n6424);
   U10167 : NAND2_X2 port map( A1 => n1671, A2 => n22289, ZN => n1781);
   U10454 : CLKBUF_X2 port map( I => Key(20), Z => n19676);
   U24457 : NOR2_X1 port map( A1 => n32843, A2 => n25815, ZN => n193);
   U29378 : NOR2_X2 port map( A1 => n25783, A2 => n10807, ZN => n15552);
   U16742 : INV_X1 port map( I => n10071, ZN => n17080);
   U2935 : NOR2_X2 port map( A1 => n19136, A2 => n6036, ZN => n15134);
   U15164 : NAND2_X1 port map( A1 => n31353, A2 => n28656, ZN => n10369);
   U3528 : INV_X1 port map( I => n29755, ZN => n29741);
   U22139 : NAND3_X2 port map( A1 => n1491, A2 => n19575, A3 => n14382, ZN => 
                           n12220);
   U8872 : INV_X2 port map( I => n20113, ZN => n29420);
   U3412 : OAI21_X2 port map( A1 => n33442, A2 => n23704, B => n24484, ZN => 
                           n346);
   U521 : NOR2_X2 port map( A1 => n7627, A2 => n7628, ZN => n7397);
   U4864 : INV_X2 port map( I => n31664, ZN => n17735);
   U25446 : NAND2_X2 port map( A1 => n9288, A2 => n9287, ZN => n33534);
   U13506 : NAND3_X2 port map( A1 => n22746, A2 => n12032, A3 => n35040, ZN => 
                           n11822);
   U4670 : NOR2_X1 port map( A1 => n32787, A2 => n32786, ZN => n32785);
   U6398 : NOR2_X2 port map( A1 => n10418, A2 => n10417, ZN => n22040);
   U10811 : NAND2_X2 port map( A1 => n30166, A2 => n1181, ZN => n30172);
   U15604 : INV_X2 port map( I => n319, ZN => n16114);
   U358 : CLKBUF_X4 port map( I => n27772, Z => n28282);
   U16967 : OAI21_X2 port map( A1 => n24516, A2 => n38749, B => n35801, ZN => 
                           n24517);
   U8117 : OAI21_X2 port map( A1 => n12629, A2 => n10055, B => n1541, ZN => 
                           n14025);
   U19037 : CLKBUF_X4 port map( I => n24878, Z => n31861);
   U17761 : INV_X1 port map( I => n39112, ZN => n8232);
   U14769 : INV_X2 port map( I => n19525, ZN => n2338);
   U29071 : NAND2_X2 port map( A1 => n25691, A2 => n18894, ZN => n25568);
   U14317 : NAND3_X1 port map( A1 => n14540, A2 => n17525, A3 => n32572, ZN => 
                           n9953);
   U20915 : NAND2_X2 port map( A1 => n7286, A2 => n19420, ZN => n8318);
   U10086 : INV_X4 port map( I => n23028, ZN => n1315);
   U9350 : INV_X2 port map( I => n26630, ZN => n26761);
   U4573 : OAI21_X2 port map( A1 => n38293, A2 => n24595, B => n30960, ZN => 
                           n25140);
   U24510 : NAND2_X2 port map( A1 => n18412, A2 => n21920, ZN => n21921);
   U30287 : NOR2_X2 port map( A1 => n16107, A2 => n15112, ZN => n5244);
   U11882 : OAI21_X2 port map( A1 => n26922, A2 => n26764, B => n26920, ZN => 
                           n26737);
   U2903 : NAND2_X2 port map( A1 => n2457, A2 => n5469, ZN => n31847);
   U8211 : NAND2_X1 port map( A1 => n7176, A2 => n9614, ZN => n20030);
   U16052 : AOI22_X2 port map( A1 => n32318, A2 => n17723, B1 => n12077, B2 => 
                           n30306, ZN => n31481);
   U9138 : BUF_X2 port map( I => n27882, Z => n28260);
   U12158 : AOI22_X2 port map( A1 => n1243, A2 => n8377, B1 => n8376, B2 => 
                           n36404, ZN => n11270);
   U5886 : OAI21_X2 port map( A1 => n28034, A2 => n9969, B => n7310, ZN => 
                           n7309);
   U2605 : INV_X4 port map( I => n28191, ZN => n28034);
   U20503 : OAI21_X1 port map( A1 => n19017, A2 => n20376, B => n21977, ZN => 
                           n21978);
   U6136 : NAND2_X2 port map( A1 => n1396, A2 => n9105, ZN => n29479);
   U17260 : NAND2_X1 port map( A1 => n16173, A2 => n27435, ZN => n5998);
   U16471 : INV_X2 port map( I => n3974, ZN => n14488);
   U11795 : NOR2_X1 port map( A1 => n16402, A2 => n33396, ZN => n16401);
   U11306 : AOI21_X1 port map( A1 => n28272, A2 => n28012, B => n8308, ZN => 
                           n8307);
   U2937 : NOR2_X2 port map( A1 => n6036, A2 => n4935, ZN => n14925);
   U7878 : NAND2_X2 port map( A1 => n26817, A2 => n20635, ZN => n20634);
   U10988 : NOR2_X2 port map( A1 => n5244, A2 => n5243, ZN => n20845);
   U12694 : NAND2_X2 port map( A1 => n24692, A2 => n30764, ZN => n24693);
   U8137 : INV_X2 port map( I => n730, ZN => n1530);
   U24456 : NAND3_X1 port map( A1 => n24181, A2 => n277, A3 => n24398, ZN => 
                           n18632);
   U20015 : NAND2_X1 port map( A1 => n19028, A2 => n37377, ZN => n11316);
   U22904 : NOR3_X2 port map( A1 => n33843, A2 => n14209, A3 => n31597, ZN => 
                           n12651);
   U16532 : INV_X1 port map( I => n14837, ZN => n12314);
   U11197 : NAND2_X1 port map( A1 => n20920, A2 => n39574, ZN => n19414);
   U6376 : INV_X2 port map( I => n12015, ZN => n963);
   U23731 : OAI22_X2 port map( A1 => n29316, A2 => n38328, B1 => n29203, B2 => 
                           n39585, ZN => n19706);
   U1645 : BUF_X2 port map( I => n18860, Z => n8368);
   U1496 : INV_X2 port map( I => n20887, ZN => n19133);
   U9122 : OAI21_X2 port map( A1 => n10288, A2 => n16869, B => n16950, ZN => 
                           n10287);
   U4929 : INV_X2 port map( I => n13166, ZN => n25422);
   U7730 : INV_X2 port map( I => n17410, ZN => n1437);
   U1534 : INV_X2 port map( I => n4116, ZN => n18657);
   U27797 : INV_X2 port map( I => n20070, ZN => n28089);
   U18036 : NAND3_X2 port map( A1 => n9456, A2 => n20962, A3 => n9457, ZN => 
                           n5073);
   U25153 : AOI21_X2 port map( A1 => n23262, A2 => n16047, B => n23401, ZN => 
                           n16757);
   U11448 : BUF_X2 port map( I => n27700, Z => n19612);
   U6578 : NAND2_X2 port map( A1 => n35248, A2 => n319, ZN => n30470);
   U13368 : AOI21_X2 port map( A1 => n23157, A2 => n23158, B => n23156, ZN => 
                           n6345);
   U24061 : NAND2_X1 port map( A1 => n18814, A2 => n38145, ZN => n20737);
   U4874 : BUF_X2 port map( I => n33324, Z => n33154);
   U10673 : INV_X4 port map( I => n30844, ZN => n6300);
   U11422 : INV_X4 port map( I => n988, ZN => n28274);
   U7053 : NAND3_X2 port map( A1 => n11214, A2 => n1134, A3 => n23383, ZN => 
                           n3746);
   U13862 : NAND2_X1 port map( A1 => n18954, A2 => n20003, ZN => n3484);
   U8661 : AOI21_X1 port map( A1 => n21522, A2 => n19511, B => n21587, ZN => 
                           n5104);
   U1987 : NAND3_X2 port map( A1 => n32626, A2 => n7130, A3 => n32625, ZN => 
                           n20907);
   U23802 : INV_X2 port map( I => n13091, ZN => n28153);
   U4630 : BUF_X4 port map( I => n24759, Z => n10019);
   U12988 : NOR2_X2 port map( A1 => n914, A2 => n12953, ZN => n4957);
   U9950 : INV_X2 port map( I => n19481, ZN => n23588);
   U2328 : AOI21_X2 port map( A1 => n28034, A2 => n36979, B => n7309, ZN => 
                           n11470);
   U7568 : INV_X1 port map( I => n1190, ZN => n18098);
   U1776 : BUF_X4 port map( I => n14491, Z => n32507);
   U4337 : INV_X2 port map( I => n21050, ZN => n1218);
   U6319 : INV_X2 port map( I => n20484, ZN => n24470);
   U13723 : AOI22_X2 port map( A1 => n20280, A2 => n13519, B1 => n20282, B2 => 
                           n1340, ZN => n19460);
   U2770 : INV_X2 port map( I => n38395, ZN => n13632);
   U10423 : BUF_X2 port map( I => n21805, Z => n19545);
   U8775 : BUF_X2 port map( I => Key(95), Z => n19885);
   U8796 : NAND2_X1 port map( A1 => n20964, A2 => n29468, ZN => n6343);
   U10394 : INV_X2 port map( I => n21111, ZN => n8468);
   U10045 : AOI21_X2 port map( A1 => n2350, A2 => n23201, B => n33697, ZN => 
                           n13527);
   U6838 : NAND2_X2 port map( A1 => n4606, A2 => n30275, ZN => n31825);
   U3083 : NOR2_X1 port map( A1 => n6203, A2 => n6201, ZN => n6208);
   U10111 : INV_X2 port map( I => n8197, ZN => n23094);
   U2779 : NOR2_X2 port map( A1 => n11090, A2 => n20528, ZN => n11089);
   U18543 : INV_X2 port map( I => n27580, ZN => n27532);
   U24621 : NAND2_X1 port map( A1 => n25919, A2 => n16814, ZN => n16813);
   U7033 : INV_X4 port map( I => n24461, ZN => n1126);
   U30560 : BUF_X2 port map( I => n9861, Z => n33921);
   U22227 : OAI21_X2 port map( A1 => n31875, A2 => n997, B => n13364, ZN => 
                           n16248);
   U3872 : INV_X2 port map( I => n261, ZN => n21565);
   U20097 : NAND2_X1 port map( A1 => n18251, A2 => n18250, ZN => n27324);
   U17462 : INV_X1 port map( I => n15159, ZN => n1541);
   U8904 : INV_X2 port map( I => n8184, ZN => n29497);
   U2384 : NAND3_X1 port map( A1 => n26686, A2 => n18357, A3 => n33301, ZN => 
                           n113);
   U2737 : INV_X4 port map( I => n15320, ZN => n914);
   U14061 : BUF_X2 port map( I => Key(175), Z => n29805);
   U8774 : BUF_X2 port map( I => Key(4), Z => n19736);
   U6456 : BUF_X2 port map( I => Key(52), Z => n29238);
   U7315 : BUF_X2 port map( I => Key(0), Z => n29399);
   U6465 : BUF_X2 port map( I => Key(31), Z => n19843);
   U10465 : BUF_X2 port map( I => Key(45), Z => n30120);
   U14041 : BUF_X2 port map( I => Key(43), Z => n30068);
   U10407 : CLKBUF_X4 port map( I => n21743, Z => n19542);
   U6451 : INV_X2 port map( I => n15354, ZN => n13855);
   U7289 : BUF_X2 port map( I => n13679, Z => n8597);
   U14021 : CLKBUF_X1 port map( I => n21722, Z => n18855);
   U14345 : INV_X1 port map( I => n19902, ZN => n31249);
   U21020 : INV_X1 port map( I => n19736, ZN => n32218);
   U13990 : BUF_X2 port map( I => n21835, Z => n19620);
   U26614 : INV_X1 port map( I => n33141, ZN => n21620);
   U13871 : NOR2_X1 port map( A1 => n21388, A2 => n21715, ZN => n16290);
   U13868 : OAI21_X1 port map( A1 => n21842, A2 => n21900, B => n15031, ZN => 
                           n12119);
   U10345 : NAND2_X1 port map( A1 => n34021, A2 => n21554, ZN => n10893);
   U1476 : NAND2_X1 port map( A1 => n21622, A2 => n8467, ZN => n2403);
   U5794 : INV_X2 port map( I => n22042, ZN => n1338);
   U27114 : INV_X2 port map( I => n21980, ZN => n22301);
   U24738 : NOR2_X1 port map( A1 => n34488, A2 => n36303, ZN => n19159);
   U6396 : INV_X2 port map( I => n22040, ZN => n22289);
   U10266 : CLKBUF_X4 port map( I => n22294, Z => n18854);
   U10155 : AOI22_X1 port map( A1 => n21262, A2 => n22268, B1 => n21261, B2 => 
                           n32259, ZN => n21260);
   U13685 : NOR2_X1 port map( A1 => n20043, A2 => n21960, ZN => n10025);
   U13701 : INV_X1 port map( I => n22213, ZN => n12030);
   U10134 : NAND2_X1 port map( A1 => n20146, A2 => n20148, ZN => n19328);
   U2097 : INV_X1 port map( I => n17943, ZN => n1670);
   U2594 : CLKBUF_X4 port map( I => n9873, Z => n3475);
   U2932 : CLKBUF_X2 port map( I => n22744, Z => n32863);
   U13594 : INV_X1 port map( I => n22604, ZN => n11254);
   U4391 : INV_X1 port map( I => n1661, ZN => n7158);
   U5050 : CLKBUF_X2 port map( I => n10962, Z => n903);
   U2015 : BUF_X2 port map( I => n12925, Z => n33247);
   U14225 : INV_X1 port map( I => n22974, ZN => n1872);
   U4785 : BUF_X2 port map( I => n20840, Z => n32032);
   U19962 : INV_X2 port map( I => n7327, ZN => n14556);
   U25722 : NOR2_X1 port map( A1 => n22974, A2 => n15163, ZN => n16733);
   U5992 : INV_X2 port map( I => n14556, ZN => n23114);
   U16021 : NOR2_X1 port map( A1 => n18071, A2 => n20408, ZN => n20743);
   U12862 : INV_X1 port map( I => n6827, ZN => n31081);
   U5100 : OAI21_X1 port map( A1 => n5786, A2 => n5785, B => n19865, ZN => 
                           n14352);
   U21855 : NAND2_X1 port map( A1 => n23033, A2 => n16967, ZN => n11435);
   U21607 : NOR2_X1 port map( A1 => n23004, A2 => n23070, ZN => n32326);
   U13452 : INV_X2 port map( I => n22512, ZN => n4473);
   U18343 : AOI21_X1 port map( A1 => n18516, A2 => n22924, B => n32216, ZN => 
                           n31736);
   U1719 : NAND2_X1 port map( A1 => n11435, A2 => n23127, ZN => n4597);
   U13444 : OAI21_X1 port map( A1 => n22995, A2 => n23067, B => n20024, ZN => 
                           n8012);
   U13399 : AOI22_X1 port map( A1 => n23112, A2 => n1142, B1 => n23113, B2 => 
                           n33196, ZN => n18702);
   U24392 : NAND2_X1 port map( A1 => n19361, A2 => n15503, ZN => n15502);
   U4217 : INV_X2 port map( I => n17094, ZN => n14845);
   U6339 : CLKBUF_X4 port map( I => n18682, Z => n5487);
   U5750 : BUF_X2 port map( I => n34959, Z => n3363);
   U3997 : CLKBUF_X4 port map( I => n31944, Z => n30506);
   U15838 : INV_X2 port map( I => n33609, ZN => n15787);
   U1857 : NAND2_X1 port map( A1 => n18199, A2 => n37523, ZN => n23274);
   U5252 : OAI21_X1 port map( A1 => n22912, A2 => n22911, B => n36191, ZN => 
                           n22914);
   U25263 : INV_X1 port map( I => n23903, ZN => n8704);
   U1150 : INV_X1 port map( I => n6527, ZN => n5071);
   U5279 : INV_X1 port map( I => n23904, ZN => n6051);
   U13027 : CLKBUF_X2 port map( I => n801, Z => n7730);
   U13048 : CLKBUF_X4 port map( I => n23907, Z => n24245);
   U10602 : CLKBUF_X2 port map( I => n24421, Z => n30833);
   U3722 : CLKBUF_X4 port map( I => n36552, Z => n6849);
   U9810 : CLKBUF_X4 port map( I => n10734, Z => n2348);
   U6562 : OR2_X1 port map( A1 => n15775, A2 => n16792, Z => n30463);
   U8340 : NOR2_X1 port map( A1 => n24446, A2 => n24445, ZN => n13708);
   U14495 : OAI21_X1 port map( A1 => n24426, A2 => n24258, B => n2089, ZN => 
                           n2088);
   U8319 : OR2_X1 port map( A1 => n23958, A2 => n8193, Z => n8194);
   U1706 : INV_X1 port map( I => n15018, ZN => n16447);
   U24881 : NAND2_X1 port map( A1 => n24474, A2 => n37916, ZN => n24475);
   U26417 : NAND2_X1 port map( A1 => n24386, A2 => n16375, ZN => n16374);
   U1005 : BUF_X2 port map( I => n20728, Z => n524);
   U3237 : BUF_X4 port map( I => n15266, Z => n3120);
   U4637 : INV_X1 port map( I => n30530, ZN => n30529);
   U3664 : OAI21_X1 port map( A1 => n24794, A2 => n36321, B => n24596, ZN => 
                           n24598);
   U1666 : NAND2_X1 port map( A1 => n31519, A2 => n32898, ZN => n31328);
   U5356 : INV_X2 port map( I => n24623, ZN => n21231);
   U4612 : BUF_X2 port map( I => n24614, Z => n33821);
   U4621 : CLKBUF_X2 port map( I => n13966, Z => n33480);
   U6992 : CLKBUF_X4 port map( I => n24623, Z => n9277);
   U3784 : OAI21_X1 port map( A1 => n15664, A2 => n34354, B => n36471, ZN => 
                           n13746);
   U1658 : NAND2_X1 port map( A1 => n9277, A2 => n33818, ZN => n14936);
   U6963 : INV_X1 port map( I => n24752, ZN => n12706);
   U951 : NAND2_X1 port map( A1 => n7342, A2 => n24659, ZN => n24178);
   U28785 : INV_X1 port map( I => n24620, ZN => n24084);
   U20218 : NAND2_X1 port map( A1 => n24622, A2 => n32064, ZN => n32063);
   U12487 : NOR2_X1 port map( A1 => n16421, A2 => n16420, ZN => n13398);
   U2662 : NOR2_X1 port map( A1 => n9438, A2 => n2931, ZN => n2930);
   U1958 : INV_X1 port map( I => n33038, ZN => n6411);
   U24864 : INV_X1 port map( I => n24935, ZN => n25024);
   U24468 : INV_X1 port map( I => n19418, ZN => n25394);
   U9564 : INV_X1 port map( I => n39289, ZN => n8879);
   U12447 : CLKBUF_X2 port map( I => n19418, Z => n18298);
   U6681 : INV_X2 port map( I => n19582, ZN => n6731);
   U4506 : CLKBUF_X4 port map( I => n11496, Z => n32419);
   U4501 : OAI21_X1 port map( A1 => n30377, A2 => n25341, B => n1543, ZN => 
                           n25344);
   U12399 : NAND2_X1 port map( A1 => n25066, A2 => n35887, ZN => n25067);
   U1240 : OAI21_X1 port map( A1 => n5483, A2 => n7853, B => n18810, ZN => 
                           n31322);
   U26900 : OAI21_X1 port map( A1 => n32419, A2 => n36249, B => n17472, ZN => 
                           n17471);
   U21851 : INV_X2 port map( I => n39140, ZN => n1244);
   U4497 : NAND2_X1 port map( A1 => n2958, A2 => n13465, ZN => n32044);
   U22287 : INV_X2 port map( I => n26041, ZN => n32469);
   U25210 : NAND2_X1 port map( A1 => n18838, A2 => n25509, ZN => n19042);
   U15042 : NAND2_X1 port map( A1 => n6221, A2 => n3575, ZN => n6220);
   U12119 : NAND2_X1 port map( A1 => n25737, A2 => n9859, ZN => n6153);
   U17155 : INV_X2 port map( I => n17212, ZN => n8481);
   U12175 : INV_X1 port map( I => n26129, ZN => n8543);
   U9384 : NAND2_X1 port map( A1 => n6152, A2 => n6153, ZN => n6150);
   U25236 : INV_X1 port map( I => n25854, ZN => n14952);
   U7985 : NAND2_X1 port map( A1 => n6478, A2 => n8255, ZN => n6219);
   U3446 : INV_X1 port map( I => n35238, ZN => n13147);
   U12047 : NAND2_X1 port map( A1 => n25739, A2 => n30621, ZN => n10509);
   U18448 : CLKBUF_X2 port map( I => n26520, Z => n32528);
   U20616 : OR2_X1 port map( A1 => n35269, A2 => n36392, Z => n32693);
   U17930 : INV_X2 port map( I => n9081, ZN => n8155);
   U2795 : INV_X2 port map( I => n14080, ZN => n26708);
   U7936 : INV_X1 port map( I => n9899, ZN => n9269);
   U27161 : NAND2_X1 port map( A1 => n26266, A2 => n26655, ZN => n19204);
   U588 : INV_X2 port map( I => n26688, ZN => n26980);
   U11750 : NAND2_X1 port map( A1 => n14485, A2 => n5405, ZN => n4483);
   U27574 : INV_X1 port map( I => n26865, ZN => n26775);
   U20162 : NAND2_X1 port map( A1 => n20547, A2 => n20754, ZN => n7469);
   U29339 : OAI21_X1 port map( A1 => n26983, A2 => n852, B => n17097, ZN => 
                           n26984);
   U23438 : NAND2_X1 port map( A1 => n26985, A2 => n26984, ZN => n18047);
   U25589 : CLKBUF_X4 port map( I => n7974, Z => n32976);
   U22767 : INV_X2 port map( I => n11020, ZN => n17166);
   U509 : INV_X2 port map( I => n14153, ZN => n27274);
   U9186 : INV_X1 port map( I => n10461, ZN => n27429);
   U5736 : INV_X1 port map( I => n19061, ZN => n32771);
   U6711 : NOR2_X1 port map( A1 => n27084, A2 => n27274, ZN => n5664);
   U24035 : OAI21_X1 port map( A1 => n10677, A2 => n27410, B => n32771, ZN => 
                           n399);
   U19671 : OAI21_X1 port map( A1 => n31943, A2 => n35299, B => n9680, ZN => 
                           n26447);
   U3690 : BUF_X4 port map( I => n10621, Z => n33690);
   U2088 : INV_X1 port map( I => n12971, ZN => n11502);
   U29865 : INV_X2 port map( I => n33522, ZN => n3158);
   U19902 : INV_X2 port map( I => n7281, ZN => n16065);
   U17161 : BUF_X4 port map( I => n27671, Z => n28024);
   U4268 : BUF_X2 port map( I => n1455, Z => n33405);
   U5484 : INV_X2 port map( I => n12218, ZN => n14500);
   U9044 : NAND2_X1 port map( A1 => n28257, A2 => n28258, ZN => n11025);
   U4259 : CLKBUF_X2 port map( I => n12909, Z => n33002);
   U11388 : NOR2_X1 port map( A1 => n438, A2 => n28205, ZN => n1753);
   U9041 : NAND2_X1 port map( A1 => n20639, A2 => n27974, ZN => n8265);
   U11301 : INV_X1 port map( I => n28004, ZN => n7984);
   U415 : NOR2_X1 port map( A1 => n3198, A2 => n32150, ZN => n33418);
   U11284 : OAI22_X1 port map( A1 => n8327, A2 => n4347, B1 => n8149, B2 => 
                           n8326, ZN => n8325);
   U27299 : INV_X2 port map( I => n28685, ZN => n1429);
   U20101 : INV_X2 port map( I => n7428, ZN => n16778);
   U11155 : INV_X2 port map( I => n10544, ZN => n3252);
   U355 : INV_X2 port map( I => n15792, ZN => n17978);
   U18074 : NOR2_X1 port map( A1 => n14516, A2 => n15631, ZN => n15630);
   U11074 : NOR2_X1 port map( A1 => n32315, A2 => n32314, ZN => n10304);
   U11072 : OAI21_X1 port map( A1 => n17073, A2 => n32595, B => n3191, ZN => 
                           n15323);
   U16924 : NAND2_X1 port map( A1 => n28718, A2 => n16505, ZN => n31608);
   U6038 : CLKBUF_X1 port map( I => n29146, Z => n30888);
   U20087 : CLKBUF_X2 port map( I => n29121, Z => n32022);
   U18785 : INV_X2 port map( I => n20460, ZN => n29081);
   U8903 : INV_X2 port map( I => n771, ZN => n1176);
   U10848 : CLKBUF_X2 port map( I => n29483, Z => n19734);
   U28063 : INV_X2 port map( I => n29196, ZN => n29701);
   U1919 : INV_X2 port map( I => n8529, ZN => n14437);
   U2471 : NAND2_X1 port map( A1 => n29702, A2 => n8941, ZN => n7502);
   U21889 : OAI21_X1 port map( A1 => n30051, A2 => n19909, B => n10671, ZN => 
                           n10670);
   U27385 : NAND2_X1 port map( A1 => n17540, A2 => n17539, ZN => n33246);
   U8868 : OAI21_X1 port map( A1 => n1060, A2 => n29702, B => n14511, ZN => 
                           n16389);
   U10734 : NAND2_X1 port map( A1 => n6207, A2 => n13573, ZN => n6206);
   U8787 : CLKBUF_X2 port map( I => Key(166), Z => n29442);
   U14034 : CLKBUF_X2 port map( I => Key(107), Z => n19801);
   U8769 : CLKBUF_X2 port map( I => Key(167), Z => n29506);
   U14065 : BUF_X2 port map( I => Key(132), Z => n19887);
   U7318 : CLKBUF_X2 port map( I => Key(91), Z => n29831);
   U5826 : CLKBUF_X2 port map( I => Key(150), Z => n9981);
   U10489 : BUF_X2 port map( I => Key(92), Z => n19851);
   U6453 : BUF_X2 port map( I => Key(106), Z => n19780);
   U7317 : BUF_X2 port map( I => Key(33), Z => n19805);
   U8766 : BUF_X2 port map( I => Key(129), Z => n19775);
   U14016 : BUF_X2 port map( I => n21674, Z => n19641);
   U7293 : INV_X1 port map( I => n29285, ZN => n1160);
   U13918 : INV_X1 port map( I => n21749, ZN => n21715);
   U5786 : INV_X2 port map( I => n22301, ZN => n20357);
   U2895 : NAND2_X1 port map( A1 => n10762, A2 => n11327, ZN => n22213);
   U19488 : OAI22_X1 port map( A1 => n11171, A2 => n35754, B1 => n34246, B2 => 
                           n22360, ZN => n15488);
   U4021 : BUF_X2 port map( I => n11778, Z => n33697);
   U13573 : BUF_X2 port map( I => n23089, Z => n19488);
   U19289 : INV_X2 port map( I => n19588, ZN => n22512);
   U1262 : BUF_X4 port map( I => n8660, Z => n6684);
   U2896 : INV_X1 port map( I => n13217, ZN => n17090);
   U1904 : INV_X1 port map( I => n23272, ZN => n18939);
   U13297 : CLKBUF_X2 port map( I => n21068, Z => n10024);
   U24906 : NOR2_X1 port map( A1 => n18762, A2 => n1039, ZN => n20997);
   U29938 : NOR2_X1 port map( A1 => n4183, A2 => n37319, ZN => n33532);
   U12822 : OAI21_X1 port map( A1 => n12120, A2 => n24469, B => n8200, ZN => 
                           n10751);
   U6970 : AOI21_X1 port map( A1 => n4666, A2 => n24132, B => n1128, ZN => 
                           n30530);
   U5357 : NAND2_X1 port map( A1 => n24591, A2 => n24694, ZN => n16079);
   U17378 : NAND2_X1 port map( A1 => n16050, A2 => n16051, ZN => n2931);
   U12522 : INV_X1 port map( I => n25040, ZN => n11964);
   U9554 : NAND2_X1 port map( A1 => n5541, A2 => n5519, ZN => n8033);
   U27774 : INV_X2 port map( I => n33948, ZN => n19963);
   U5453 : NOR2_X1 port map( A1 => n299, A2 => n19495, ZN => n25066);
   U23372 : CLKBUF_X4 port map( I => n16836, Z => n32654);
   U9476 : OAI21_X1 port map( A1 => n7956, A2 => n30633, B => n19490, ZN => 
                           n2766);
   U12114 : INV_X1 port map( I => n25933, ZN => n12721);
   U3763 : OAI21_X1 port map( A1 => n25737, A2 => n25887, B => n26070, ZN => 
                           n6152);
   U1697 : OAI21_X1 port map( A1 => n8543, A2 => n34745, B => n31827, ZN => 
                           n25405);
   U3893 : NOR2_X1 port map( A1 => n4138, A2 => n26797, ZN => n9179);
   U11800 : NAND2_X1 port map( A1 => n9731, A2 => n26951, ZN => n4689);
   U2126 : INV_X2 port map( I => n12755, ZN => n6891);
   U3928 : BUF_X1 port map( I => n31014, Z => n30871);
   U606 : NAND3_X1 port map( A1 => n1474, A2 => n16237, A3 => n16263, ZN => 
                           n27312);
   U29412 : NAND2_X1 port map( A1 => n4782, A2 => n3531, ZN => n1939);
   U9146 : NAND2_X1 port map( A1 => n10574, A2 => n16966, ZN => n10580);
   U26744 : CLKBUF_X1 port map( I => n27779, Z => n20772);
   U16281 : BUF_X2 port map( I => n5402, Z => n4347);
   U30535 : BUF_X2 port map( I => n37056, Z => n33902);
   U7705 : INV_X1 port map( I => n6990, ZN => n8522);
   U256 : INV_X2 port map( I => n5237, ZN => n9141);
   U11131 : INV_X1 port map( I => n14760, ZN => n12717);
   U7925 : INV_X1 port map( I => n28301, ZN => n21025);
   U11122 : INV_X1 port map( I => n28370, ZN => n13824);
   U158 : NAND2_X2 port map( A1 => n11665, A2 => n11664, ZN => n28840);
   U10850 : AND2_X1 port map( A1 => n21299, A2 => n15153, Z => n10628);
   U5832 : CLKBUF_X2 port map( I => n29684, Z => n19497);
   U4433 : NOR2_X2 port map( A1 => n25939, A2 => n17915, ZN => n20612);
   U2963 : BUF_X2 port map( I => n9001, Z => n32309);
   U28079 : INV_X2 port map( I => n21184, ZN => n29454);
   U9636 : INV_X2 port map( I => n24635, ZN => n3125);
   U4533 : INV_X4 port map( I => n12246, ZN => n13366);
   U13985 : BUF_X2 port map( I => n15370, Z => n14783);
   U4228 : BUF_X2 port map( I => n18450, Z => n452);
   U6424 : BUF_X2 port map( I => n19387, Z => n4759);
   U10412 : INV_X1 port map( I => n21777, ZN => n21465);
   U4894 : NOR2_X1 port map( A1 => n35921, A2 => n1348, ZN => n15456);
   U8723 : NAND2_X1 port map( A1 => n10120, A2 => n8799, ZN => n13701);
   U6156 : INV_X1 port map( I => n19641, ZN => n33053);
   U12309 : NAND2_X1 port map( A1 => n3562, A2 => n10629, ZN => n31035);
   U27471 : NOR2_X1 port map( A1 => n19479, A2 => n19091, ZN => n21632);
   U1517 : INV_X1 port map( I => n35921, ZN => n21440);
   U2191 : NOR2_X1 port map( A1 => n35921, A2 => n18152, ZN => n21842);
   U24751 : AOI21_X1 port map( A1 => n21656, A2 => n17938, B => n21780, ZN => 
                           n18877);
   U13916 : OAI21_X1 port map( A1 => n21465, A2 => n19091, B => n21939, ZN => 
                           n15437);
   U30373 : NAND2_X1 port map( A1 => n8700, A2 => n21775, ZN => n19075);
   U10406 : BUF_X2 port map( I => n13473, Z => n13472);
   U2200 : NAND2_X1 port map( A1 => n15696, A2 => n32164, ZN => n32163);
   U2007 : NOR2_X1 port map( A1 => n37111, A2 => n32123, ZN => n20368);
   U21947 : NOR2_X1 port map( A1 => n18412, A2 => n21111, ZN => n21621);
   U6418 : INV_X1 port map( I => n18926, ZN => n21557);
   U20666 : INV_X1 port map( I => n7935, ZN => n14837);
   U27340 : NOR2_X1 port map( A1 => n8700, A2 => n18710, ZN => n21940);
   U24532 : NAND3_X1 port map( A1 => n19517, A2 => n21672, A3 => n18219, ZN => 
                           n16654);
   U17769 : AOI22_X1 port map( A1 => n8700, A2 => n19479, B1 => n19350, B2 => 
                           n21775, ZN => n18712);
   U28253 : NAND2_X1 port map( A1 => n21666, A2 => n32412, ZN => n21437);
   U13874 : AOI21_X1 port map( A1 => n17679, A2 => n21309, B => n17678, ZN => 
                           n6669);
   U24733 : NOR2_X1 port map( A1 => n15097, A2 => n21822, ZN => n15096);
   U24754 : INV_X1 port map( I => n21932, ZN => n21607);
   U13932 : OAI21_X1 port map( A1 => n21333, A2 => n2531, B => n21889, ZN => 
                           n15814);
   U1492 : NOR2_X1 port map( A1 => n13472, A2 => n5751, ZN => n21377);
   U5008 : NOR2_X1 port map( A1 => n20328, A2 => n21551, ZN => n21653);
   U25953 : AOI21_X1 port map( A1 => n21498, A2 => n20003, B => n32164, ZN => 
                           n16287);
   U27341 : OAI21_X1 port map( A1 => n21775, A2 => n18710, B => n8700, ZN => 
                           n21609);
   U26070 : OAI22_X1 port map( A1 => n21437, A2 => n19620, B1 => n20682, B2 => 
                           n21666, ZN => n15490);
   U13863 : OAI21_X1 port map( A1 => n21467, A2 => n21468, B => n11411, ZN => 
                           n2737);
   U1976 : INV_X2 port map( I => n21587, ZN => n21588);
   U8653 : NOR2_X1 port map( A1 => n16901, A2 => n3865, ZN => n3864);
   U6401 : BUF_X2 port map( I => n22389, Z => n4239);
   U13759 : NAND2_X1 port map( A1 => n14027, A2 => n17086, ZN => n17664);
   U16601 : NAND2_X1 port map( A1 => n8496, A2 => n19373, ZN => n22069);
   U6395 : NOR2_X1 port map( A1 => n18303, A2 => n1746, ZN => n3086);
   U10273 : INV_X1 port map( I => n11044, ZN => n22220);
   U14165 : INV_X1 port map( I => n11344, ZN => n22325);
   U6394 : INV_X1 port map( I => n22362, ZN => n1672);
   U6402 : INV_X1 port map( I => n22389, ZN => n4240);
   U17243 : NOR2_X1 port map( A1 => n17074, A2 => n10632, ZN => n10631);
   U18844 : NAND2_X1 port map( A1 => n6036, A2 => n22315, ZN => n18674);
   U10275 : INV_X1 port map( I => n19373, ZN => n1681);
   U26031 : NAND2_X1 port map( A1 => n7613, A2 => n22184, ZN => n21974);
   U10236 : AOI21_X1 port map( A1 => n6451, A2 => n1151, B => n22177, ZN => 
                           n16282);
   U28377 : NAND2_X1 port map( A1 => n1048, A2 => n21973, ZN => n21975);
   U21861 : NAND2_X1 port map( A1 => n36563, A2 => n22332, ZN => n22065);
   U4979 : INV_X1 port map( I => n22364, ZN => n22366);
   U4803 : INV_X1 port map( I => n22315, ZN => n22156);
   U1408 : INV_X1 port map( I => n3269, ZN => n3268);
   U5788 : INV_X2 port map( I => n12077, ZN => n17723);
   U8581 : INV_X1 port map( I => n22289, ZN => n17531);
   U18481 : INV_X1 port map( I => n22215, ZN => n22361);
   U3131 : INV_X1 port map( I => n20889, ZN => n22140);
   U20604 : AOI21_X1 port map( A1 => n164, A2 => n22293, B => n22140, ZN => 
                           n33792);
   U9006 : NOR2_X1 port map( A1 => n8118, A2 => n22148, ZN => n30706);
   U1764 : NAND2_X1 port map( A1 => n22064, A2 => n3680, ZN => n3679);
   U5450 : INV_X1 port map( I => n22332, ZN => n22252);
   U15641 : NAND3_X1 port map( A1 => n3181, A2 => n34407, A3 => n13632, ZN => 
                           n21926);
   U1406 : NAND2_X1 port map( A1 => n8348, A2 => n7613, ZN => n20256);
   U26544 : AOI21_X1 port map( A1 => n22140, A2 => n33713, B => n18854, ZN => 
                           n20354);
   U17907 : OAI21_X1 port map( A1 => n22498, A2 => n1154, B => n31648, ZN => 
                           n18635);
   U4982 : INV_X1 port map( I => n22741, ZN => n11500);
   U6372 : INV_X1 port map( I => n20353, ZN => n22583);
   U10122 : INV_X1 port map( I => n22529, ZN => n22515);
   U26666 : INV_X1 port map( I => n22699, ZN => n17223);
   U16458 : INV_X1 port map( I => n22789, ZN => n22601);
   U2042 : NOR2_X1 port map( A1 => n1142, A2 => n12392, ZN => n33763);
   U2038 : INV_X2 port map( I => n22929, ZN => n22865);
   U1318 : INV_X1 port map( I => n3952, ZN => n23032);
   U17563 : INV_X2 port map( I => n23078, ZN => n23182);
   U24005 : INV_X1 port map( I => n782, ZN => n23084);
   U24829 : NAND2_X1 port map( A1 => n23169, A2 => n531, ZN => n18147);
   U13473 : NAND2_X1 port map( A1 => n1042, A2 => n1320, ZN => n3200);
   U25972 : BUF_X2 port map( I => n21132, Z => n33045);
   U23498 : INV_X1 port map( I => n301, ZN => n32677);
   U10106 : INV_X1 port map( I => n23131, ZN => n23211);
   U5995 : NAND2_X1 port map( A1 => n23181, A2 => n23078, ZN => n8673);
   U27322 : NOR2_X1 port map( A1 => n9954, A2 => n18679, ZN => n19659);
   U28565 : NOR2_X1 port map( A1 => n22866, A2 => n22865, ZN => n22867);
   U8751 : NAND3_X1 port map( A1 => n18244, A2 => n13042, A3 => n23101, ZN => 
                           n30676);
   U8551 : INV_X2 port map( I => n23125, ZN => n23197);
   U10052 : NOR2_X1 port map( A1 => n14396, A2 => n13719, ZN => n14724);
   U16597 : INV_X1 port map( I => n23067, ZN => n4107);
   U1319 : INV_X1 port map( I => n3273, ZN => n22955);
   U20186 : NOR2_X1 port map( A1 => n13734, A2 => n903, ZN => n13775);
   U13541 : OR2_X1 port map( A1 => n34014, A2 => n59, Z => n23127);
   U5110 : OAI21_X1 port map( A1 => n22867, A2 => n22991, B => n39500, ZN => 
                           n22868);
   U8471 : AOI21_X1 port map( A1 => n272, A2 => n19351, B => n9238, ZN => 
                           n14189);
   U10009 : AOI21_X1 port map( A1 => n36839, A2 => n23214, B => n5569, ZN => 
                           n2254);
   U24432 : AOI21_X1 port map( A1 => n1316, A2 => n20174, B => n1648, ZN => 
                           n15503);
   U15096 : NAND2_X1 port map( A1 => n22899, A2 => n36369, ZN => n31351);
   U13537 : NOR2_X1 port map( A1 => n3273, A2 => n19621, ZN => n3542);
   U21415 : NAND2_X1 port map( A1 => n23023, A2 => n9080, ZN => n23027);
   U4210 : OAI21_X1 port map( A1 => n13775, A2 => n23105, B => n23104, ZN => 
                           n4903);
   U2752 : NOR2_X1 port map( A1 => n14882, A2 => n13408, ZN => n13407);
   U28609 : NAND3_X1 port map( A1 => n33045, A2 => n17691, A3 => n23178, ZN => 
                           n23180);
   U13370 : OAI21_X1 port map( A1 => n3547, A2 => n3546, B => n19621, ZN => 
                           n3545);
   U15031 : AOI21_X1 port map( A1 => n6500, A2 => n1650, B => n6498, ZN => 
                           n6497);
   U27628 : INV_X2 port map( I => n32024, ZN => n33287);
   U3451 : INV_X1 port map( I => n5357, ZN => n12790);
   U2100 : CLKBUF_X2 port map( I => n17094, Z => n14901);
   U7118 : INV_X1 port map( I => n23566, ZN => n1643);
   U13340 : INV_X2 port map( I => n23496, ZN => n23315);
   U3863 : AOI21_X1 port map( A1 => n35068, A2 => n13305, B => n35501, ZN => 
                           n13304);
   U18449 : NAND2_X1 port map( A1 => n33496, A2 => n10480, ZN => n23284);
   U2978 : INV_X1 port map( I => n23308, ZN => n1631);
   U2552 : NAND2_X1 port map( A1 => n23307, A2 => n16182, ZN => n23479);
   U20667 : INV_X1 port map( I => n23250, ZN => n7939);
   U1180 : INV_X1 port map( I => n12154, ZN => n20955);
   U17529 : AND2_X1 port map( A1 => n71, A2 => n70, Z => n31586);
   U8379 : NAND2_X1 port map( A1 => n1290, A2 => n9862, ZN => n23439);
   U13130 : NAND2_X1 port map( A1 => n23439, A2 => n23440, ZN => n9971);
   U6326 : NAND2_X1 port map( A1 => n23575, A2 => n1134, ZN => n3583);
   U28619 : NAND3_X1 port map( A1 => n1134, A2 => n23571, A3 => n7485, ZN => 
                           n23232);
   U9964 : INV_X1 port map( I => n17511, ZN => n23474);
   U13146 : OAI21_X1 port map( A1 => n22967, A2 => n23493, B => n22966, ZN => 
                           n22972);
   U7115 : NAND4_X1 port map( A1 => n23432, A2 => n23433, A3 => n23434, A4 => 
                           n23431, ZN => n23559);
   U7094 : NOR2_X1 port map( A1 => n23624, A2 => n33894, ZN => n23625);
   U6674 : NOR2_X1 port map( A1 => n4600, A2 => n1310, ZN => n21156);
   U23776 : NOR2_X1 port map( A1 => n13305, A2 => n33349, ZN => n23281);
   U28647 : AOI21_X1 port map( A1 => n18284, A2 => n5083, B => n23458, ZN => 
                           n23372);
   U13308 : INV_X1 port map( I => n18989, ZN => n16484);
   U2517 : AOI21_X1 port map( A1 => n23312, A2 => n6421, B => n1637, ZN => 
                           n23313);
   U5243 : NAND3_X1 port map( A1 => n33720, A2 => n33719, A3 => n12154, ZN => 
                           n15495);
   U9874 : NAND2_X1 port map( A1 => n35545, A2 => n36965, ZN => n8054);
   U21764 : OAI21_X1 port map( A1 => n32363, A2 => n33721, B => n32362, ZN => 
                           n23369);
   U20233 : OAI21_X1 port map( A1 => n23282, A2 => n39194, B => n32068, ZN => 
                           n16883);
   U28623 : NAND2_X1 port map( A1 => n36564, A2 => n36027, ZN => n23259);
   U25160 : OAI21_X1 port map( A1 => n12093, A2 => n36027, B => n36564, ZN => 
                           n14721);
   U17484 : NAND2_X1 port map( A1 => n10989, A2 => n8054, ZN => n8053);
   U8364 : INV_X1 port map( I => n23774, ZN => n2221);
   U9833 : NAND3_X1 port map( A1 => n36701, A2 => n36011, A3 => n1160, ZN => 
                           n12819);
   U1152 : INV_X1 port map( I => n23899, ZN => n20340);
   U28795 : INV_X1 port map( I => n24300, ZN => n24110);
   U18174 : NAND2_X1 port map( A1 => n12235, A2 => n16081, ZN => n31697);
   U14451 : INV_X1 port map( I => n2052, ZN => n24383);
   U6321 : INV_X1 port map( I => n16792, ZN => n11585);
   U9791 : OAI21_X1 port map( A1 => n19402, A2 => n37848, B => n6515, ZN => 
                           n24198);
   U24276 : NAND2_X1 port map( A1 => n1597, A2 => n24143, ZN => n14156);
   U9766 : NAND2_X1 port map( A1 => n24359, A2 => n19895, ZN => n4051);
   U21506 : NAND2_X1 port map( A1 => n39605, A2 => n24282, ZN => n32492);
   U12895 : INV_X1 port map( I => n19864, ZN => n20396);
   U9768 : NAND2_X1 port map( A1 => n17871, A2 => n33450, ZN => n24152);
   U1729 : NAND2_X1 port map( A1 => n24194, A2 => n6515, ZN => n32491);
   U1787 : OAI21_X1 port map( A1 => n1128, A2 => n1130, B => n32069, ZN => 
                           n24474);
   U12849 : NAND2_X1 port map( A1 => n24473, A2 => n39309, ZN => n2579);
   U8328 : NOR2_X1 port map( A1 => n2348, A2 => n1285, ZN => n14292);
   U28812 : NAND2_X1 port map( A1 => n1599, A2 => n13453, ZN => n24217);
   U8299 : NOR2_X1 port map( A1 => n24390, A2 => n2348, ZN => n16829);
   U1712 : NAND2_X1 port map( A1 => n12481, A2 => n12202, ZN => n32183);
   U22917 : NOR2_X1 port map( A1 => n32891, A2 => n17911, ZN => n5855);
   U13004 : INV_X1 port map( I => n33450, ZN => n24449);
   U3360 : NOR2_X1 port map( A1 => n10008, A2 => n17810, ZN => n32938);
   U9717 : NOR2_X1 port map( A1 => n24411, A2 => n37651, ZN => n12423);
   U17758 : AOI21_X1 port map( A1 => n18116, A2 => n33240, B => n39373, ZN => 
                           n31621);
   U6999 : OAI21_X1 port map( A1 => n13881, A2 => n8581, B => n14392, ZN => 
                           n13742);
   U9698 : OAI21_X1 port map( A1 => n24472, A2 => n24471, B => n1130, ZN => 
                           n24476);
   U12965 : NOR2_X1 port map( A1 => n6839, A2 => n19942, ZN => n9722);
   U12959 : NOR2_X1 port map( A1 => n801, A2 => n24266, ZN => n11194);
   U6969 : NAND2_X1 port map( A1 => n10116, A2 => n17087, ZN => n5388);
   U12395 : NAND2_X1 port map( A1 => n31044, A2 => n24434, ZN => n24511);
   U24749 : INV_X2 port map( I => n15467, ZN => n32882);
   U5964 : AOI22_X1 port map( A1 => n5358, A2 => n37264, B1 => n24147, B2 => 
                           n1604, ZN => n5359);
   U8253 : INV_X1 port map( I => n35981, ZN => n1583);
   U26820 : INV_X2 port map( I => n15426, ZN => n19901);
   U20158 : NAND2_X1 port map( A1 => n24620, A2 => n19868, ZN => n24622);
   U5379 : NOR2_X1 port map( A1 => n16210, A2 => n24782, ZN => n7342);
   U3832 : NAND4_X1 port map( A1 => n13045, A2 => n23796, A3 => n13048, A4 => 
                           n13047, ZN => n13046);
   U25202 : AOI21_X1 port map( A1 => n5056, A2 => n958, B => n16077, ZN => 
                           n16076);
   U12524 : NOR2_X1 port map( A1 => n18168, A2 => n6037, ZN => n8578);
   U25206 : NAND2_X1 port map( A1 => n24695, A2 => n19565, ZN => n24619);
   U6990 : INV_X1 port map( I => n24782, ZN => n24660);
   U981 : NAND2_X1 port map( A1 => n24698, A2 => n37097, ZN => n24581);
   U3667 : AOI21_X1 port map( A1 => n24794, A2 => n7445, B => n36321, ZN => 
                           n10141);
   U12723 : NAND2_X1 port map( A1 => n31796, A2 => n37477, ZN => n1948);
   U20024 : NAND2_X1 port map( A1 => n24619, A2 => n11126, ZN => n11258);
   U20036 : NOR2_X1 port map( A1 => n24732, A2 => n24639, ZN => n12782);
   U1578 : OAI21_X1 port map( A1 => n14999, A2 => n1566, B => n33480, ZN => 
                           n30941);
   U9651 : NAND2_X1 port map( A1 => n11712, A2 => n24592, ZN => n3750);
   U27708 : INV_X1 port map( I => n39196, ZN => n1574);
   U28700 : NAND2_X1 port map( A1 => n35901, A2 => n34354, ZN => n23705);
   U28097 : NAND2_X1 port map( A1 => n33344, A2 => n7520, ZN => n18468);
   U972 : INV_X2 port map( I => n1580, ZN => n7831);
   U2659 : OR2_X1 port map( A1 => n15266, A2 => n7520, Z => n24849);
   U3057 : NOR2_X1 port map( A1 => n11712, A2 => n24849, ZN => n24850);
   U1661 : NAND2_X1 port map( A1 => n37983, A2 => n39279, ZN => n30700);
   U10348 : OAI21_X1 port map( A1 => n7286, A2 => n8314, B => n30554, ZN => 
                           n24834);
   U28883 : OAI21_X1 port map( A1 => n37396, A2 => n4973, B => n24733, ZN => 
                           n24595);
   U3831 : NOR2_X1 port map( A1 => n5871, A2 => n31722, ZN => n18504);
   U12555 : NAND3_X1 port map( A1 => n24747, A2 => n24887, A3 => n13735, ZN => 
                           n16195);
   U9608 : OAI21_X1 port map( A1 => n4909, A2 => n24608, B => n4908, ZN => 
                           n7064);
   U28855 : NAND3_X1 port map( A1 => n24691, A2 => n24765, A3 => n18324, ZN => 
                           n24493);
   U28847 : NAND2_X1 port map( A1 => n34138, A2 => n24795, ZN => n24439);
   U26131 : NAND2_X1 port map( A1 => n34138, A2 => n35981, ZN => n17267);
   U2012 : NAND2_X1 port map( A1 => n30764, A2 => n24717, ZN => n24720);
   U28886 : NAND2_X1 port map( A1 => n19886, A2 => n33821, ZN => n24616);
   U3967 : AOI22_X1 port map( A1 => n24671, A2 => n1119, B1 => n24670, B2 => 
                           n30843, ZN => n12418);
   U1554 : NOR3_X1 port map( A1 => n18570, A2 => n31346, A3 => n35521, ZN => 
                           n18569);
   U4601 : NAND2_X1 port map( A1 => n12672, A2 => n12654, ZN => n30598);
   U923 : NAND2_X1 port map( A1 => n6335, A2 => n442, ZN => n11738);
   U17496 : OAI21_X1 port map( A1 => n13340, A2 => n32019, B => n17453, ZN => 
                           n13342);
   U869 : INV_X1 port map( I => n25598, ZN => n20515);
   U5312 : BUF_X2 port map( I => n20627, Z => n16677);
   U1395 : INV_X1 port map( I => n2799, ZN => n32085);
   U21048 : INV_X1 port map( I => n31669, ZN => n14413);
   U12377 : NOR2_X1 port map( A1 => n4664, A2 => n833, ZN => n17472);
   U6913 : INV_X2 port map( I => n6300, ZN => n12629);
   U9584 : INV_X1 port map( I => n11496, ZN => n1256);
   U14638 : NAND2_X1 port map( A1 => n3602, A2 => n33491, ZN => n20746);
   U30114 : OAI21_X1 port map( A1 => n34755, A2 => n3602, B => n9815, ZN => 
                           n17305);
   U16478 : NAND3_X1 port map( A1 => n4467, A2 => n33268, A3 => n25361, ZN => 
                           n4464);
   U24878 : NAND2_X1 port map( A1 => n12309, A2 => n25574, ZN => n18029);
   U23218 : OAI21_X1 port map( A1 => n1543, A2 => n38178, B => n7853, ZN => 
                           n25342);
   U12317 : NAND2_X1 port map( A1 => n11873, A2 => n1249, ZN => n11549);
   U786 : OAI21_X1 port map( A1 => n16316, A2 => n5455, B => n6894, ZN => n5454
                           );
   U16343 : NAND2_X1 port map( A1 => n541, A2 => n25620, ZN => n11550);
   U21721 : NOR2_X1 port map( A1 => n25620, A2 => n541, ZN => n9602);
   U6887 : INV_X1 port map( I => n6448, ZN => n20121);
   U6559 : INV_X1 port map( I => n4603, ZN => n25688);
   U6580 : INV_X1 port map( I => n19589, ZN => n20856);
   U9498 : AOI22_X1 port map( A1 => n4664, A2 => n4047, B1 => n19637, B2 => 
                           n32419, ZN => n4046);
   U29066 : NOR2_X1 port map( A1 => n517, A2 => n16933, ZN => n25547);
   U18223 : NAND2_X1 port map( A1 => n9915, A2 => n25699, ZN => n31707);
   U14835 : NAND3_X1 port map( A1 => n14443, A2 => n25489, A3 => n38245, ZN => 
                           n31820);
   U29021 : NAND2_X1 port map( A1 => n25342, A2 => n12533, ZN => n25343);
   U12408 : NAND2_X1 port map( A1 => n25617, A2 => n25616, ZN => n5248);
   U9487 : NAND2_X1 port map( A1 => n7284, A2 => n7876, ZN => n7875);
   U12400 : NAND2_X1 port map( A1 => n12131, A2 => n32868, ZN => n10313);
   U8109 : OAI21_X1 port map( A1 => n25638, A2 => n25716, B => n25637, ZN => 
                           n18108);
   U1223 : NOR2_X1 port map( A1 => n33491, A2 => n3602, ZN => n31457);
   U8132 : NOR2_X1 port map( A1 => n6573, A2 => n25416, ZN => n14915);
   U12358 : AOI21_X1 port map( A1 => n7875, A2 => n11495, B => n1255, ZN => 
                           n7874);
   U8793 : OAI21_X1 port map( A1 => n25045, A2 => n17480, B => n25467, ZN => 
                           n30677);
   U5597 : INV_X2 port map( I => n4699, ZN => n32747);
   U1187 : INV_X1 port map( I => n26020, ZN => n31311);
   U14300 : INV_X2 port map( I => n31242, ZN => n11834);
   U9443 : INV_X1 port map( I => n36922, ZN => n26058);
   U24887 : NAND2_X1 port map( A1 => n14793, A2 => n36226, ZN => n18283);
   U3475 : NOR2_X1 port map( A1 => n31192, A2 => n36546, ZN => n2892);
   U759 : CLKBUF_X2 port map( I => n25956, Z => n318);
   U12202 : INV_X2 port map( I => n25814, ZN => n26131);
   U5544 : INV_X1 port map( I => n7660, ZN => n11762);
   U9402 : OAI21_X1 port map( A1 => n4602, A2 => n4516, B => n929, ZN => n12002
                           );
   U17281 : OAI21_X1 port map( A1 => n25928, A2 => n5356, B => n30302, ZN => 
                           n14774);
   U12192 : NAND2_X1 port map( A1 => n1106, A2 => n14793, ZN => n16432);
   U1133 : NOR2_X1 port map( A1 => n25747, A2 => n1524, ZN => n32782);
   U8304 : OAI21_X1 port map( A1 => n2892, A2 => n2891, B => n6390, ZN => 
                           n30651);
   U29102 : NAND2_X1 port map( A1 => n33348, A2 => n26020, ZN => n25748);
   U6837 : OAI21_X1 port map( A1 => n4382, A2 => n2625, B => n25334, ZN => 
                           n6105);
   U2210 : NAND2_X1 port map( A1 => n16867, A2 => n25966, ZN => n32333);
   U2635 : NAND2_X1 port map( A1 => n6222, A2 => n6390, ZN => n30546);
   U2707 : INV_X1 port map( I => n33909, ZN => n26133);
   U20195 : INV_X2 port map( I => n15677, ZN => n32052);
   U23088 : NOR2_X1 port map( A1 => n19740, A2 => n11834, ZN => n11624);
   U9430 : NOR2_X1 port map( A1 => n25940, A2 => n1528, ZN => n13524);
   U8042 : CLKBUF_X2 port map( I => n18176, Z => n6578);
   U662 : NAND2_X1 port map( A1 => n603, A2 => n25797, ZN => n25911);
   U6946 : INV_X1 port map( I => n26093, ZN => n931);
   U15268 : OAI22_X1 port map( A1 => n10321, A2 => n25447, B1 => n17700, B2 => 
                           n31367, ZN => n31831);
   U12128 : OAI21_X1 port map( A1 => n13119, A2 => n25869, B => n1017, ZN => 
                           n13118);
   U16062 : NAND2_X1 port map( A1 => n7961, A2 => n3575, ZN => n25879);
   U6824 : OAI21_X1 port map( A1 => n14573, A2 => n1106, B => n25768, ZN => 
                           n6103);
   U17724 : NOR2_X1 port map( A1 => n13869, A2 => n446, ZN => n12895);
   U6843 : AOI21_X1 port map( A1 => n25993, A2 => n19740, B => n12234, ZN => 
                           n16397);
   U4448 : NAND2_X1 port map( A1 => n3838, A2 => n21040, ZN => n3837);
   U669 : NAND2_X1 port map( A1 => n26065, A2 => n9530, ZN => n26066);
   U1028 : NAND2_X1 port map( A1 => n32109, A2 => n13732, ZN => n5552);
   U26122 : INV_X1 port map( I => n9743, ZN => n18002);
   U7512 : NOR2_X1 port map( A1 => n32721, A2 => n30568, ZN => n14286);
   U12030 : INV_X1 port map( I => n20600, ZN => n7439);
   U14563 : NAND2_X1 port map( A1 => n31654, A2 => n13391, ZN => n13068);
   U5664 : INV_X1 port map( I => n26594, ZN => n26484);
   U7964 : INV_X1 port map( I => n5848, ZN => n26499);
   U16652 : INV_X1 port map( I => n7018, ZN => n7028);
   U3035 : INV_X1 port map( I => n3781, ZN => n19024);
   U27261 : INV_X1 port map( I => n18490, ZN => n19217);
   U637 : INV_X1 port map( I => n5084, ZN => n26588);
   U12008 : INV_X1 port map( I => n26334, ZN => n8310);
   U529 : INV_X2 port map( I => n19951, ZN => n1088);
   U20239 : BUF_X2 port map( I => n14347, Z => n7527);
   U6185 : INV_X2 port map( I => n14962, ZN => n13588);
   U11805 : NAND2_X1 port map( A1 => n32168, A2 => n26970, ZN => n17575);
   U4526 : INV_X1 port map( I => n37524, ZN => n12549);
   U2612 : AOI21_X1 port map( A1 => n14377, A2 => n19179, B => n26811, ZN => 
                           n26632);
   U567 : INV_X1 port map( I => n26665, ZN => n26978);
   U2763 : NAND2_X1 port map( A1 => n3369, A2 => n3368, ZN => n30725);
   U29296 : NAND3_X1 port map( A1 => n7978, A2 => n26703, A3 => n26702, ZN => 
                           n26705);
   U15959 : NOR2_X1 port map( A1 => n26934, A2 => n32745, ZN => n4970);
   U24655 : NAND2_X1 port map( A1 => n26952, A2 => n37055, ZN => n15251);
   U20942 : OAI21_X1 port map( A1 => n4138, A2 => n20699, B => n26797, ZN => 
                           n18792);
   U27600 : NOR2_X1 port map( A1 => n7527, A2 => n35967, ZN => n26628);
   U18949 : NAND2_X1 port map( A1 => n6190, A2 => n26265, ZN => n26266);
   U9261 : NOR2_X1 port map( A1 => n14382, A2 => n10355, ZN => n7392);
   U29309 : NOR2_X1 port map( A1 => n13393, A2 => n26918, ZN => n26766);
   U30166 : NOR2_X1 port map( A1 => n26841, A2 => n20578, ZN => n11708);
   U2616 : NAND2_X1 port map( A1 => n19179, A2 => n12755, ZN => n31647);
   U7954 : INV_X2 port map( I => n14355, ZN => n26722);
   U4394 : BUF_X2 port map( I => n14459, Z => n32797);
   U15824 : NAND2_X1 port map( A1 => n19700, A2 => n14459, ZN => n26691);
   U856 : NAND2_X1 port map( A1 => n20575, A2 => n26612, ZN => n11387);
   U6766 : AOI21_X1 port map( A1 => n4138, A2 => n7516, B => n26797, ZN => 
                           n9764);
   U24647 : NOR2_X1 port map( A1 => n38577, A2 => n6615, ZN => n17785);
   U11853 : NAND2_X1 port map( A1 => n26663, A2 => n15825, ZN => n7005);
   U9271 : NAND2_X1 port map( A1 => n33333, A2 => n26932, ZN => n6605);
   U6758 : OAI21_X1 port map( A1 => n20882, A2 => n26815, B => n1497, ZN => 
                           n18311);
   U24956 : NOR2_X1 port map( A1 => n26803, A2 => n15594, ZN => n19505);
   U21006 : NAND2_X1 port map( A1 => n17237, A2 => n31526, ZN => n8465);
   U6833 : NOR2_X1 port map( A1 => n5480, A2 => n5481, ZN => n5479);
   U6171 : NAND2_X1 port map( A1 => n15763, A2 => n26975, ZN => n19694);
   U29262 : OR2_X1 port map( A1 => n26930, A2 => n26564, Z => n26581);
   U749 : INV_X2 port map( I => n9956, ZN => n27198);
   U489 : INV_X2 port map( I => n1487, ZN => n27406);
   U5884 : INV_X1 port map( I => n3092, ZN => n27401);
   U7828 : INV_X1 port map( I => n27449, ZN => n27263);
   U27417 : INV_X1 port map( I => n27283, ZN => n33254);
   U7126 : AOI21_X1 port map( A1 => n27387, A2 => n35299, B => n39826, ZN => 
                           n30542);
   U27373 : INV_X1 port map( I => n27211, ZN => n20092);
   U1560 : INV_X1 port map( I => n27397, ZN => n2520);
   U4348 : BUF_X2 port map( I => n9956, Z => n9201);
   U9216 : NAND2_X1 port map( A1 => n27395, A2 => n9956, ZN => n11805);
   U29373 : NAND2_X1 port map( A1 => n27298, A2 => n27378, ZN => n27171);
   U24965 : OAI21_X1 port map( A1 => n27391, A2 => n35895, B => n13699, ZN => 
                           n18250);
   U24381 : NOR2_X1 port map( A1 => n27438, A2 => n34977, ZN => n14764);
   U9172 : OAI21_X1 port map( A1 => n30986, A2 => n10051, B => n12156, ZN => 
                           n9454);
   U10657 : NAND2_X1 port map( A1 => n15360, A2 => n1000, ZN => n30840);
   U425 : INV_X1 port map( I => n27181, ZN => n7418);
   U6162 : INV_X2 port map( I => n27484, ZN => n11039);
   U29344 : NAND2_X1 port map( A1 => n27358, A2 => n15360, ZN => n27020);
   U24563 : NOR2_X1 port map( A1 => n2949, A2 => n7606, ZN => n32852);
   U9203 : NAND2_X1 port map( A1 => n38060, A2 => n12485, ZN => n27207);
   U25253 : NAND3_X1 port map( A1 => n13471, A2 => n27199, A3 => n27198, ZN => 
                           n26914);
   U11507 : NAND2_X1 port map( A1 => n13793, A2 => n35897, ZN => n13792);
   U27576 : NAND2_X1 port map( A1 => n26999, A2 => n27054, ZN => n19802);
   U29361 : NOR2_X1 port map( A1 => n36911, A2 => n27455, ZN => n27103);
   U15938 : AOI22_X1 port map( A1 => n27055, A2 => n31672, B1 => n1475, B2 => 
                           n3466, ZN => n3467);
   U7762 : NAND2_X1 port map( A1 => n19077, A2 => n27265, ZN => n18986);
   U26138 : NAND3_X1 port map( A1 => n27154, A2 => n5311, A3 => n27406, ZN => 
                           n26789);
   U6733 : INV_X2 port map( I => n2760, ZN => n27388);
   U17194 : NAND2_X1 port map( A1 => n7231, A2 => n27181, ZN => n7230);
   U14825 : NAND2_X1 port map( A1 => n14261, A2 => n38900, ZN => n27559);
   U15365 : NAND2_X1 port map( A1 => n15276, A2 => n36969, ZN => n15275);
   U5525 : AOI22_X1 port map( A1 => n11039, A2 => n11038, B1 => n27401, B2 => 
                           n11043, ZN => n11037);
   U2607 : INV_X1 port map( I => n27735, ZN => n27596);
   U3501 : INV_X1 port map( I => n5899, ZN => n6990);
   U16402 : INV_X1 port map( I => n1455, ZN => n20184);
   U298 : NAND3_X1 port map( A1 => n28032, A2 => n8149, A3 => n1204, ZN => 
                           n9663);
   U25464 : NAND2_X1 port map( A1 => n989, A2 => n1069, ZN => n14640);
   U15718 : INV_X2 port map( I => n11512, ZN => n31942);
   U14315 : INV_X1 port map( I => n28093, ZN => n16950);
   U12457 : AND2_X1 port map( A1 => n33958, A2 => n19764, Z => n28148);
   U9092 : NOR2_X1 port map( A1 => n17032, A2 => n28267, ZN => n3231);
   U310 : NAND2_X1 port map( A1 => n3158, A2 => n28248, ZN => n28251);
   U3904 : OAI21_X1 port map( A1 => n33185, A2 => n16987, B => n1071, ZN => 
                           n30991);
   U24111 : NAND3_X1 port map( A1 => n1442, A2 => n28054, A3 => n1205, ZN => 
                           n13696);
   U11286 : NAND2_X1 port map( A1 => n28035, A2 => n7310, ZN => n13599);
   U7625 : NOR2_X1 port map( A1 => n27934, A2 => n19435, ZN => n10228);
   U24995 : OAI21_X1 port map( A1 => n28193, A2 => n28194, B => n27866, ZN => 
                           n27906);
   U24673 : NAND2_X1 port map( A1 => n17197, A2 => n17598, ZN => n27930);
   U30544 : NOR2_X1 port map( A1 => n18665, A2 => n28266, ZN => n33912);
   U11339 : NAND2_X1 port map( A1 => n17390, A2 => n28290, ZN => n7190);
   U7685 : INV_X1 port map( I => n28267, ZN => n20519);
   U5395 : INV_X1 port map( I => n14562, ZN => n28265);
   U21482 : INV_X1 port map( I => n28152, ZN => n9169);
   U4015 : AOI21_X1 port map( A1 => n36844, A2 => n28248, B => n37451, ZN => 
                           n12531);
   U15473 : NOR2_X1 port map( A1 => n33307, A2 => n28025, ZN => n20967);
   U7661 : NAND2_X1 port map( A1 => n5403, A2 => n21160, ZN => n3843);
   U7633 : NAND3_X1 port map( A1 => n28085, A2 => n6643, A3 => n989, ZN => 
                           n28086);
   U23235 : NAND3_X1 port map( A1 => n28283, A2 => n28067, A3 => n7528, ZN => 
                           n32778);
   U11250 : OAI22_X1 port map( A1 => n27929, A2 => n3511, B1 => n28193, B2 => 
                           n27930, ZN => n5706);
   U16910 : NAND2_X1 port map( A1 => n28024, A2 => n4803, ZN => n27666);
   U17699 : NAND3_X1 port map( A1 => n28251, A2 => n21223, A3 => n28249, ZN => 
                           n31606);
   U3569 : OR2_X1 port map( A1 => n15727, A2 => n28220, Z => n11648);
   U19496 : OAI21_X1 port map( A1 => n6643, A2 => n18841, B => n6777, ZN => 
                           n27917);
   U6198 : OR2_X1 port map( A1 => n28047, A2 => n3990, Z => n30350);
   U9068 : OAI22_X1 port map( A1 => n15694, A2 => n21137, B1 => n15695, B2 => 
                           n28193, ZN => n4504);
   U14109 : AOI21_X1 port map( A1 => n28266, A2 => n14562, B => n28267, ZN => 
                           n28176);
   U6649 : NAND2_X1 port map( A1 => n28223, A2 => n2868, ZN => n3069);
   U5926 : NOR2_X1 port map( A1 => n10166, A2 => n33185, ZN => n3533);
   U8521 : NOR2_X1 port map( A1 => n27917, A2 => n1069, ZN => n30980);
   U254 : INV_X1 port map( I => n27908, ZN => n28299);
   U6621 : INV_X1 port map( I => n28713, ZN => n1425);
   U4209 : CLKBUF_X2 port map( I => n5237, Z => n33591);
   U6117 : INV_X1 port map( I => n11296, ZN => n15022);
   U5855 : INV_X1 port map( I => n28537, ZN => n28495);
   U3239 : INV_X1 port map( I => n34559, ZN => n1187);
   U11142 : NAND2_X1 port map( A1 => n10618, A2 => n5662, ZN => n18089);
   U11079 : AOI21_X1 port map( A1 => n8800, A2 => n28553, B => n18984, ZN => 
                           n2327);
   U11064 : INV_X1 port map( I => n13598, ZN => n16308);
   U25306 : INV_X1 port map( I => n32575, ZN => n16038);
   U11015 : NOR2_X1 port map( A1 => n18018, A2 => n13563, ZN => n28693);
   U4164 : INV_X1 port map( I => n18990, ZN => n33107);
   U7501 : OAI21_X1 port map( A1 => n8759, A2 => n39147, B => n28440, ZN => 
                           n9783);
   U21119 : NAND3_X1 port map( A1 => n16398, A2 => n8714, A3 => n13151, ZN => 
                           n33190);
   U222 : INV_X1 port map( I => n16107, ZN => n28499);
   U29633 : OAI21_X1 port map( A1 => n28685, A2 => n18871, B => n39724, ZN => 
                           n28586);
   U10982 : NAND2_X1 port map( A1 => n28428, A2 => n28661, ZN => n12797);
   U6550 : INV_X2 port map( I => n30055, ZN => n1057);
   U10844 : NAND2_X1 port map( A1 => n29937, A2 => n14557, ZN => n6692);
   U2380 : BUF_X2 port map( I => n28414, Z => n29699);
   U101 : INV_X1 port map( I => n29769, ZN => n1063);
   U8874 : NAND2_X1 port map( A1 => n29815, A2 => n14600, ZN => n13573);
   U10843 : INV_X1 port map( I => n29581, ZN => n20085);
   U2910 : NAND2_X1 port map( A1 => n2296, A2 => n31667, ZN => n894);
   U26264 : OAI21_X1 port map( A1 => n12878, A2 => n14525, B => n16828, ZN => 
                           n33092);
   U29800 : INV_X1 port map( I => n16828, ZN => n29382);
   U2359 : INV_X2 port map( I => n29454, ZN => n17295);
   U2574 : NOR2_X1 port map( A1 => n8919, A2 => n37060, ZN => n14755);
   U104 : INV_X1 port map( I => n30195, ZN => n33394);
   U1843 : NOR2_X1 port map( A1 => n1182, A2 => n29195, ZN => n8346);
   U25863 : NAND2_X1 port map( A1 => n29776, A2 => n29781, ZN => n16790);
   U5582 : INV_X1 port map( I => n30153, ZN => n19480);
   U78 : NAND2_X1 port map( A1 => n29211, A2 => n17225, ZN => n30655);
   U14718 : NAND2_X1 port map( A1 => n31296, A2 => n19909, ZN => n10435);
   U25333 : INV_X1 port map( I => n14773, ZN => n29316);
   U5578 : OAI21_X1 port map( A1 => n32671, A2 => n14400, B => n31095, ZN => 
                           n15864);
   U20647 : NOR2_X1 port map( A1 => n29892, A2 => n971, ZN => n10832);
   U15237 : NOR2_X1 port map( A1 => n36207, A2 => n30198, ZN => n2768);
   U68 : NAND3_X1 port map( A1 => n1401, A2 => n37100, A3 => n9733, ZN => 
                           n29400);
   U5575 : NAND2_X1 port map( A1 => n7164, A2 => n7163, ZN => n13384);
   U7373 : INV_X1 port map( I => n29339, ZN => n29318);
   U2381 : NOR2_X1 port map( A1 => n30071, A2 => n4377, ZN => n30070);
   U27745 : INV_X2 port map( I => n15643, ZN => n30037);
   U12 : INV_X1 port map( I => n1391, ZN => n20481);
   U16973 : AND2_X1 port map( A1 => n8399, A2 => n18457, Z => n31534);
   U22922 : OAI21_X1 port map( A1 => n30107, A2 => n35186, B => n12203, ZN => 
                           n18483);
   U5 : NOR2_X1 port map( A1 => n30127, A2 => n17193, ZN => n34706);
   U17 : NAND2_X1 port map( A1 => n30022, A2 => n30034, ZN => n30003);
   U35 : OR2_X1 port map( A1 => n4377, A2 => n4378, Z => n6489);
   U53 : INV_X1 port map( I => n30259, ZN => n32865);
   U63 : NOR2_X1 port map( A1 => n11596, A2 => n11594, ZN => n35185);
   U90 : NOR2_X1 port map( A1 => n1400, A2 => n30161, ZN => n36607);
   U98 : OAI21_X1 port map( A1 => n19050, A2 => n6938, B => n34344, ZN => 
                           n34589);
   U106 : NAND2_X1 port map( A1 => n29896, A2 => n21167, ZN => n36402);
   U114 : NAND2_X1 port map( A1 => n482, A2 => n1181, ZN => n36022);
   U121 : NAND3_X1 port map( A1 => n7207, A2 => n12940, A3 => n29262, ZN => 
                           n32189);
   U132 : NOR2_X1 port map( A1 => n21287, A2 => n105, ZN => n32498);
   U147 : NAND2_X1 port map( A1 => n21270, A2 => n29586, ZN => n34805);
   U160 : NOR2_X1 port map( A1 => n37060, A2 => n20018, ZN => n34761);
   U182 : AND2_X1 port map( A1 => n16353, A2 => n20102, Z => n34082);
   U193 : INV_X1 port map( I => n29643, ZN => n34006);
   U212 : INV_X1 port map( I => n5289, ZN => n36990);
   U239 : AOI22_X1 port map( A1 => n2822, A2 => n30894, B1 => n16777, B2 => 
                           n28633, ZN => n14929);
   U240 : INV_X1 port map( I => n34893, ZN => n13422);
   U248 : AND2_X1 port map( A1 => n11330, A2 => n39435, Z => n12605);
   U261 : OAI21_X1 port map( A1 => n36814, A2 => n16303, B => n16304, ZN => 
                           n28399);
   U264 : NAND2_X1 port map( A1 => n36671, A2 => n1193, ZN => n36567);
   U273 : AND2_X1 port map( A1 => n35173, A2 => n28496, Z => n34172);
   U280 : NOR3_X1 port map( A1 => n36791, A2 => n15224, A3 => n13151, ZN => 
                           n34893);
   U289 : NAND2_X1 port map( A1 => n30894, A2 => n1190, ZN => n28632);
   U292 : OR2_X1 port map( A1 => n5418, A2 => n31015, Z => n31077);
   U295 : NAND2_X1 port map( A1 => n28505, A2 => n11164, ZN => n34794);
   U301 : NAND2_X1 port map( A1 => n31643, A2 => n34539, ZN => n28467);
   U308 : OR2_X1 port map( A1 => n17583, A2 => n5424, Z => n30949);
   U311 : NOR2_X1 port map( A1 => n28650, A2 => n18960, ZN => n11469);
   U320 : AOI21_X1 port map( A1 => n36993, A2 => n12653, B => n15022, ZN => 
                           n35935);
   U323 : NAND3_X1 port map( A1 => n30716, A2 => n1420, A3 => n314, ZN => 
                           n36124);
   U350 : OR2_X1 port map( A1 => n31871, A2 => n6713, Z => n35182);
   U363 : BUF_X2 port map( I => n28713, Z => n36671);
   U367 : NAND2_X1 port map( A1 => n30894, A2 => n28669, ZN => n36993);
   U388 : NAND2_X1 port map( A1 => n28544, A2 => n13133, ZN => n34539);
   U389 : NAND2_X1 port map( A1 => n32575, A2 => n36320, ZN => n6819);
   U402 : NAND2_X1 port map( A1 => n33707, A2 => n28695, ZN => n10305);
   U423 : NAND2_X1 port map( A1 => n1424, A2 => n36791, ZN => n15235);
   U431 : NAND2_X1 port map( A1 => n28724, A2 => n28723, ZN => n18814);
   U444 : NAND3_X1 port map( A1 => n33002, A2 => n889, A3 => n16325, ZN => 
                           n34832);
   U451 : NAND3_X1 port map( A1 => n35659, A2 => n35658, A3 => n35657, ZN => 
                           n36236);
   U458 : OAI21_X1 port map( A1 => n34442, A2 => n34441, B => n20519, ZN => 
                           n35570);
   U472 : NAND2_X1 port map( A1 => n8232, A2 => n28224, ZN => n35658);
   U480 : AOI22_X1 port map( A1 => n12723, A2 => n3990, B1 => n28256, B2 => 
                           n28172, ZN => n36936);
   U483 : NAND2_X1 port map( A1 => n28151, A2 => n28152, ZN => n37015);
   U488 : INV_X1 port map( I => n5239, ZN => n19280);
   U491 : OAI21_X1 port map( A1 => n28165, A2 => n37057, B => n28274, ZN => 
                           n36052);
   U493 : NOR2_X1 port map( A1 => n15704, A2 => n33931, ZN => n36689);
   U494 : AND2_X1 port map( A1 => n17410, A2 => n28165, Z => n34028);
   U496 : NAND2_X1 port map( A1 => n34948, A2 => n34949, ZN => n34470);
   U499 : INV_X1 port map( I => n4809, ZN => n34442);
   U520 : NOR2_X1 port map( A1 => n9514, A2 => n1438, ZN => n28206);
   U531 : AOI21_X1 port map( A1 => n28163, A2 => n7690, B => n27979, ZN => 
                           n6236);
   U556 : NAND2_X1 port map( A1 => n28156, A2 => n28290, ZN => n34186);
   U564 : NOR2_X1 port map( A1 => n28290, A2 => n877, ZN => n16513);
   U583 : OR2_X1 port map( A1 => n988, A2 => n14399, Z => n34069);
   U597 : NAND2_X1 port map( A1 => n28260, A2 => n34410, ZN => n34948);
   U602 : BUF_X2 port map( I => n21126, Z => n13714);
   U617 : AND2_X1 port map( A1 => n1445, A2 => n35225, Z => n20188);
   U630 : NOR2_X1 port map( A1 => n1204, A2 => n33656, ZN => n18044);
   U632 : NAND2_X1 port map( A1 => n4457, A2 => n14389, ZN => n18530);
   U661 : INV_X1 port map( I => n27792, ZN => n34812);
   U670 : INV_X1 port map( I => n27657, ZN => n35853);
   U673 : INV_X1 port map( I => n27829, ZN => n34531);
   U681 : INV_X1 port map( I => n9013, ZN => n1464);
   U683 : NOR2_X1 port map( A1 => n36234, A2 => n20740, ZN => n15984);
   U685 : NAND2_X1 port map( A1 => n4105, A2 => n4104, ZN => n9739);
   U688 : AND2_X1 port map( A1 => n34769, A2 => n27165, Z => n18768);
   U690 : OR2_X1 port map( A1 => n27403, A2 => n36865, Z => n34111);
   U692 : OR2_X1 port map( A1 => n27372, A2 => n37890, Z => n27373);
   U697 : NOR2_X1 port map( A1 => n35825, A2 => n33146, ZN => n34777);
   U702 : NAND2_X1 port map( A1 => n2306, A2 => n1891, ZN => n34811);
   U703 : AND2_X1 port map( A1 => n35904, A2 => n27284, Z => n19570);
   U726 : INV_X1 port map( I => n36200, ZN => n27311);
   U740 : AND2_X1 port map( A1 => n9369, A2 => n30986, Z => n18489);
   U741 : CLKBUF_X1 port map( I => n27383, Z => n33336);
   U742 : AND2_X1 port map( A1 => n6686, A2 => n11729, Z => n27231);
   U745 : NAND2_X1 port map( A1 => n27364, A2 => n5772, ZN => n36073);
   U751 : NAND3_X1 port map( A1 => n27131, A2 => n27343, A3 => n36183, ZN => 
                           n26999);
   U758 : AOI21_X1 port map( A1 => n39305, A2 => n33893, B => n16043, ZN => 
                           n34705);
   U779 : AND2_X1 port map( A1 => n19477, A2 => n27349, Z => n30429);
   U795 : NOR2_X1 port map( A1 => n995, A2 => n1226, ZN => n13266);
   U820 : AOI21_X1 port map( A1 => n18246, A2 => n33773, B => n27416, ZN => 
                           n33235);
   U831 : AND2_X1 port map( A1 => n10171, A2 => n27583, Z => n8698);
   U834 : INV_X1 port map( I => n27284, ZN => n1084);
   U837 : NOR2_X1 port map( A1 => n27137, A2 => n8798, ZN => n18652);
   U859 : NAND2_X1 port map( A1 => n32602, A2 => n7978, ZN => n36243);
   U917 : NAND3_X1 port map( A1 => n35489, A2 => n34058, A3 => n1088, ZN => 
                           n26657);
   U920 : OR2_X1 port map( A1 => n26961, A2 => n20936, Z => n8650);
   U921 : AND2_X1 port map( A1 => n13111, A2 => n19364, Z => n34071);
   U935 : NAND2_X1 port map( A1 => n33302, A2 => n26619, ZN => n36589);
   U944 : NAND2_X1 port map( A1 => n3825, A2 => n11226, ZN => n4195);
   U961 : NAND3_X1 port map( A1 => n2100, A2 => n2101, A3 => n4211, ZN => 
                           n30715);
   U982 : NOR2_X1 port map( A1 => n20573, A2 => n17237, ZN => n11709);
   U983 : OR2_X1 port map( A1 => n26703, A2 => n10440, Z => n34058);
   U995 : NOR2_X1 port map( A1 => n3825, A2 => n11138, ZN => n15314);
   U1000 : OAI21_X1 port map( A1 => n26852, A2 => n14453, B => n5537, ZN => 
                           n35612);
   U1002 : AND2_X1 port map( A1 => n26876, A2 => n14455, Z => n2081);
   U1009 : INV_X1 port map( I => n26824, ZN => n26424);
   U1010 : NAND2_X1 port map( A1 => n18903, A2 => n19615, ZN => n18902);
   U1012 : NOR2_X1 port map( A1 => n26878, A2 => n26879, ZN => n3369);
   U1013 : INV_X2 port map( I => n26619, ZN => n26951);
   U1019 : CLKBUF_X2 port map( I => n26666, Z => n19449);
   U1026 : NAND2_X1 port map( A1 => n26849, A2 => n10314, ZN => n34908);
   U1027 : OR2_X1 port map( A1 => n13605, A2 => n5869, Z => n4410);
   U1031 : AND2_X1 port map( A1 => n26961, A2 => n35259, Z => n34075);
   U1067 : CLKBUF_X2 port map( I => n26931, Z => n19222);
   U1069 : OR2_X1 port map( A1 => n32623, A2 => n15386, Z => n26671);
   U1084 : BUF_X2 port map( I => n19436, Z => n13111);
   U1091 : INV_X1 port map( I => n18012, ZN => n33551);
   U1103 : OAI21_X1 port map( A1 => n11386, A2 => n7260, B => n33030, ZN => 
                           n35240);
   U1142 : NAND2_X1 port map( A1 => n16397, A2 => n25994, ZN => n36951);
   U1153 : AND2_X1 port map( A1 => n2561, A2 => n2029, Z => n25846);
   U1157 : NAND2_X1 port map( A1 => n15677, A2 => n36666, ZN => n36665);
   U1160 : NAND2_X1 port map( A1 => n18176, A2 => n25348, ZN => n35891);
   U1167 : AND2_X1 port map( A1 => n25742, A2 => n25770, Z => n34018);
   U1173 : OR2_X1 port map( A1 => n2865, A2 => n3642, Z => n25926);
   U1183 : NAND3_X1 port map( A1 => n586, A2 => n1020, A3 => n26018, ZN => 
                           n15966);
   U1201 : NAND3_X1 port map( A1 => n26121, A2 => n26123, A3 => n26122, ZN => 
                           n8133);
   U1202 : NOR2_X1 port map( A1 => n25945, A2 => n31523, ZN => n26331);
   U1203 : NOR2_X1 port map( A1 => n11834, A2 => n25956, ZN => n34573);
   U1204 : OR2_X1 port map( A1 => n26015, A2 => n31719, Z => n12457);
   U1235 : NAND3_X1 port map( A1 => n18283, A2 => n18282, A3 => n3356, ZN => 
                           n18426);
   U1246 : AND2_X1 port map( A1 => n33258, A2 => n26093, Z => n8005);
   U1250 : NAND2_X1 port map( A1 => n26070, A2 => n34685, ZN => n15795);
   U1278 : OR2_X1 port map( A1 => n9916, A2 => n26134, Z => n32843);
   U1298 : INV_X1 port map( I => n834, ZN => n36906);
   U1315 : NAND2_X1 port map( A1 => n36451, A2 => n36449, ZN => n17372);
   U1335 : NOR3_X1 port map( A1 => n17915, A2 => n8481, A3 => n7767, ZN => 
                           n8480);
   U1357 : CLKBUF_X4 port map( I => n35138, Z => n365);
   U1385 : BUF_X4 port map( I => n25951, Z => n34217);
   U1398 : OAI21_X1 port map( A1 => n25525, A2 => n25526, B => n517, ZN => 
                           n25530);
   U1411 : OAI21_X1 port map( A1 => n36941, A2 => n36940, B => n19095, ZN => 
                           n13210);
   U1431 : OAI21_X1 port map( A1 => n35171, A2 => n25699, B => n31721, ZN => 
                           n24957);
   U1437 : NOR2_X1 port map( A1 => n1536, A2 => n12368, ZN => n35660);
   U1438 : NAND2_X1 port map( A1 => n35763, A2 => n11550, ZN => n11544);
   U1459 : INV_X1 port map( I => n7391, ZN => n36411);
   U1462 : AND2_X1 port map( A1 => n611, A2 => n25328, Z => n14631);
   U1494 : OR2_X1 port map( A1 => n14410, A2 => n6731, Z => n34078);
   U1501 : NOR2_X1 port map( A1 => n6300, A2 => n33495, ZN => n34487);
   U1503 : NOR2_X1 port map( A1 => n39599, A2 => n37993, ZN => n25638);
   U1510 : NAND2_X1 port map( A1 => n6731, A2 => n37051, ZN => n35349);
   U1515 : NAND2_X1 port map( A1 => n25603, A2 => n21302, ZN => n25605);
   U1543 : NAND2_X1 port map( A1 => n25462, A2 => n36133, ZN => n36132);
   U1588 : CLKBUF_X2 port map( I => n25631, Z => n5051);
   U1589 : NOR2_X1 port map( A1 => n19548, A2 => n5050, ZN => n25393);
   U1590 : AND2_X1 port map( A1 => n13460, A2 => n25422, Z => n34081);
   U1596 : NOR2_X1 port map( A1 => n14708, A2 => n15541, ZN => n36487);
   U1601 : OR2_X1 port map( A1 => n33950, A2 => n25692, Z => n12780);
   U1603 : INV_X1 port map( I => n15172, ZN => n36524);
   U1607 : NOR2_X1 port map( A1 => n25484, A2 => n3985, ZN => n36135);
   U1609 : INV_X1 port map( I => n25486, ZN => n19829);
   U1622 : OAI21_X1 port map( A1 => n12533, A2 => n31010, B => n14436, ZN => 
                           n8034);
   U1624 : NAND2_X1 port map( A1 => n841, A2 => n18164, ZN => n9800);
   U1626 : NOR2_X1 port map( A1 => n20888, A2 => n25614, ZN => n10034);
   U1630 : CLKBUF_X1 port map( I => n14481, Z => n36086);
   U1634 : NOR2_X1 port map( A1 => n20515, A2 => n3602, ZN => n25068);
   U1635 : AND2_X1 port map( A1 => n252, A2 => n16931, Z => n25495);
   U1670 : CLKBUF_X1 port map( I => n20153, Z => n32904);
   U1674 : BUF_X2 port map( I => n25490, Z => n25620);
   U1723 : INV_X1 port map( I => n8542, ZN => n5434);
   U1771 : NOR2_X1 port map( A1 => n13518, A2 => n8264, ZN => n36786);
   U1774 : AND2_X1 port map( A1 => n24728, A2 => n3510, Z => n20180);
   U1783 : OR2_X1 port map( A1 => n24900, A2 => n19279, Z => n30419);
   U1795 : NOR2_X1 port map( A1 => n24646, A2 => n24794, ZN => n18570);
   U1798 : NOR2_X1 port map( A1 => n24605, A2 => n24774, ZN => n31122);
   U1804 : NOR2_X1 port map( A1 => n24669, A2 => n24668, ZN => n36787);
   U1807 : INV_X1 port map( I => n24749, ZN => n24751);
   U1809 : AND2_X1 port map( A1 => n24683, A2 => n36058, Z => n18056);
   U1813 : CLKBUF_X2 port map( I => n36058, Z => n35801);
   U1823 : OR2_X1 port map( A1 => n16841, A2 => n24799, Z => n11942);
   U1828 : NAND3_X1 port map( A1 => n259, A2 => n24630, A3 => n24826, ZN => 
                           n37017);
   U1836 : NOR2_X1 port map( A1 => n24828, A2 => n9218, ZN => n24816);
   U1853 : AND2_X1 port map( A1 => n24416, A2 => n17351, Z => n24507);
   U1869 : NAND2_X1 port map( A1 => n9478, A2 => n34796, ZN => n34904);
   U1877 : INV_X2 port map( I => n15332, ZN => n33344);
   U1878 : OAI21_X1 port map( A1 => n34039, A2 => n19566, B => n34384, ZN => 
                           n24324);
   U1882 : NAND2_X1 port map( A1 => n31519, A2 => n24784, ZN => n24613);
   U1895 : AND2_X1 port map( A1 => n1600, A2 => n19782, Z => n34039);
   U1898 : OAI21_X1 port map( A1 => n33379, A2 => n13653, B => n19566, ZN => 
                           n34384);
   U1899 : OR2_X1 port map( A1 => n39196, A2 => n24805, Z => n24532);
   U1901 : INV_X1 port map( I => n24819, ZN => n1565);
   U1902 : OAI21_X1 port map( A1 => n24630, A2 => n9218, B => n24826, ZN => 
                           n34796);
   U1903 : NOR2_X1 port map( A1 => n9197, A2 => n24879, ZN => n35048);
   U1926 : NAND2_X1 port map( A1 => n24819, A2 => n8646, ZN => n14166);
   U1929 : NOR2_X1 port map( A1 => n39818, A2 => n34758, ZN => n34420);
   U1937 : NOR2_X1 port map( A1 => n19653, A2 => n35712, ZN => n35840);
   U1950 : NOR2_X1 port map( A1 => n3133, A2 => n12953, ZN => n36273);
   U1953 : NOR2_X1 port map( A1 => n35150, A2 => n5855, ZN => n5854);
   U1964 : NOR3_X1 port map( A1 => n1125, A2 => n31452, A3 => n6515, ZN => 
                           n35086);
   U1983 : NAND2_X1 port map( A1 => n24459, A2 => n24457, ZN => n36157);
   U1993 : NOR2_X1 port map( A1 => n19782, A2 => n1600, ZN => n35872);
   U2001 : CLKBUF_X1 port map( I => n23819, Z => n35712);
   U2002 : CLKBUF_X2 port map( I => n16459, Z => n609);
   U2004 : BUF_X2 port map( I => n24142, Z => n36757);
   U2013 : NAND2_X1 port map( A1 => n14491, A2 => n1605, ZN => n35004);
   U2014 : NOR3_X1 port map( A1 => n24443, A2 => n253, A3 => n30833, ZN => 
                           n35815);
   U2053 : NAND2_X1 port map( A1 => n24158, A2 => n1280, ZN => n31852);
   U2060 : AND2_X1 port map( A1 => n32899, A2 => n9193, Z => n31490);
   U2069 : NOR2_X1 port map( A1 => n6465, A2 => n1275, ZN => n36622);
   U2073 : NOR2_X1 port map( A1 => n19584, A2 => n24419, ZN => n35814);
   U2091 : CLKBUF_X2 port map( I => n36500, Z => n35761);
   U2095 : AND2_X1 port map( A1 => n18302, A2 => n14378, Z => n34074);
   U2101 : NAND2_X1 port map( A1 => n1606, A2 => n24245, ZN => n14662);
   U2113 : AND2_X1 port map( A1 => n33057, A2 => n24104, Z => n24331);
   U2121 : NOR2_X1 port map( A1 => n24169, A2 => n277, ZN => n34655);
   U2125 : BUF_X2 port map( I => n24308, Z => n19745);
   U2128 : BUF_X2 port map( I => n24317, Z => n19782);
   U2147 : INV_X1 port map( I => n23912, ZN => n23957);
   U2154 : OAI21_X1 port map( A1 => n34337, A2 => n34336, B => n23560, ZN => 
                           n14354);
   U2160 : AOI21_X1 port map( A1 => n1301, A2 => n33316, B => n23444, ZN => 
                           n10989);
   U2162 : OR2_X1 port map( A1 => n10143, A2 => n39401, Z => n7819);
   U2175 : NAND2_X1 port map( A1 => n34602, A2 => n36129, ZN => n35355);
   U2176 : NAND3_X1 port map( A1 => n37774, A2 => n23602, A3 => n35664, ZN => 
                           n30276);
   U2190 : NAND2_X1 port map( A1 => n35974, A2 => n35536, ZN => n430);
   U2202 : AOI21_X1 port map( A1 => n23522, A2 => n23521, B => n36219, ZN => 
                           n19227);
   U2203 : OAI21_X1 port map( A1 => n3309, A2 => n5591, B => n34635, ZN => 
                           n3745);
   U2205 : OAI21_X1 port map( A1 => n11468, A2 => n12851, B => n15122, ZN => 
                           n12982);
   U2207 : NOR2_X1 port map( A1 => n35938, A2 => n7335, ZN => n34337);
   U2223 : NAND3_X1 port map( A1 => n35892, A2 => n23641, A3 => n1310, ZN => 
                           n9609);
   U2225 : AOI21_X1 port map( A1 => n11453, A2 => n23746, B => n960, ZN => 
                           n6910);
   U2243 : INV_X2 port map( I => n35331, ZN => n23444);
   U2261 : NOR2_X1 port map( A1 => n33840, A2 => n34506, ZN => n2681);
   U2263 : NAND2_X1 port map( A1 => n23494, A2 => n4147, ZN => n36129);
   U2299 : OR2_X1 port map( A1 => n33747, A2 => n35367, Z => n23383);
   U2301 : BUF_X2 port map( I => n3496, Z => n35938);
   U2321 : INV_X1 port map( I => n13038, ZN => n35501);
   U2327 : OR2_X1 port map( A1 => n8757, A2 => n19005, Z => n34068);
   U2334 : NAND3_X1 port map( A1 => n32032, A2 => n36185, A3 => n36184, ZN => 
                           n11473);
   U2336 : NOR2_X1 port map( A1 => n36422, A2 => n32515, ZN => n34696);
   U2341 : INV_X1 port map( I => n33544, ZN => n35955);
   U2344 : NAND2_X1 port map( A1 => n34713, A2 => n1044, ZN => n10553);
   U2364 : NOR2_X1 port map( A1 => n19524, A2 => n22900, ZN => n34401);
   U2372 : NAND2_X1 port map( A1 => n19586, A2 => n23084, ZN => n23186);
   U2382 : NOR2_X1 port map( A1 => n1314, A2 => n23084, ZN => n9769);
   U2396 : NOR3_X1 port map( A1 => n14089, A2 => n1046, A3 => n20267, ZN => 
                           n4773);
   U2400 : NAND2_X1 port map( A1 => n22899, A2 => n23201, ZN => n36638);
   U2402 : NAND2_X1 port map( A1 => n32515, A2 => n33925, ZN => n13945);
   U2408 : INV_X1 port map( I => n1831, ZN => n35288);
   U2410 : INV_X1 port map( I => n5581, ZN => n35591);
   U2412 : CLKBUF_X2 port map( I => n19966, Z => n35918);
   U2415 : CLKBUF_X2 port map( I => n23122, Z => n19351);
   U2434 : BUF_X2 port map( I => n13587, Z => n1763);
   U2440 : NOR2_X1 port map( A1 => n23165, A2 => n36554, ZN => n36553);
   U2456 : INV_X1 port map( I => n12961, ZN => n14439);
   U2464 : INV_X1 port map( I => n22443, ZN => n35848);
   U2473 : NAND2_X1 port map( A1 => n36466, A2 => n1329, ZN => n7867);
   U2476 : INV_X1 port map( I => n19328, ZN => n22687);
   U2481 : INV_X1 port map( I => n22665, ZN => n34545);
   U2489 : AND2_X1 port map( A1 => n2765, A2 => n34808, Z => n2435);
   U2495 : INV_X1 port map( I => n37217, ZN => n34015);
   U2502 : NAND2_X1 port map( A1 => n22390, A2 => n19873, ZN => n13778);
   U2506 : OR2_X1 port map( A1 => n19655, A2 => n22160, Z => n34023);
   U2510 : NAND3_X1 port map( A1 => n22246, A2 => n33571, A3 => n20889, ZN => 
                           n19080);
   U2511 : OAI21_X1 port map( A1 => n22344, A2 => n21987, B => n22341, ZN => 
                           n1838);
   U2521 : INV_X1 port map( I => n3863, ZN => n35822);
   U2528 : NAND2_X1 port map( A1 => n22282, A2 => n22130, ZN => n21963);
   U2535 : INV_X2 port map( I => n20376, ZN => n36661);
   U2542 : AND2_X1 port map( A1 => n9387, A2 => n22222, Z => n19253);
   U2543 : INV_X1 port map( I => n15229, ZN => n34925);
   U2546 : OR2_X1 port map( A1 => n2765, A2 => n22243, Z => n4864);
   U2548 : NAND2_X1 port map( A1 => n22091, A2 => n19837, ZN => n22097);
   U2551 : NOR2_X1 port map( A1 => n22271, A2 => n22316, ZN => n36139);
   U2565 : NAND2_X1 port map( A1 => n1333, A2 => n18656, ZN => n18730);
   U2572 : INV_X1 port map( I => n22067, ZN => n36563);
   U2575 : NAND2_X1 port map( A1 => n39489, A2 => n6947, ZN => n6946);
   U2582 : NOR2_X2 port map( A1 => n8442, A2 => n8440, ZN => n22400);
   U2588 : NAND2_X1 port map( A1 => n12927, A2 => n21932, ZN => n16660);
   U2593 : AOI22_X1 port map( A1 => n18742, A2 => n36519, B1 => n4084, B2 => 
                           n18710, ZN => n35833);
   U2596 : OAI21_X1 port map( A1 => n16163, A2 => n21601, B => n17102, ZN => 
                           n7551);
   U2622 : INV_X1 port map( I => n21743, ZN => n17266);
   U2632 : AND2_X1 port map( A1 => n12144, A2 => n1351, Z => n12142);
   U2634 : NAND2_X1 port map( A1 => n12332, A2 => n16305, ZN => n35999);
   U2636 : INV_X1 port map( I => n21410, ZN => n35043);
   U2639 : OAI22_X1 port map( A1 => n21556, A2 => n19323, B1 => n21620, B2 => 
                           n18412, ZN => n36353);
   U2644 : INV_X1 port map( I => n36062, ZN => n14450);
   U2649 : NOR2_X1 port map( A1 => n18710, A2 => n21630, ZN => n21631);
   U2653 : INV_X1 port map( I => n21576, ZN => n36781);
   U2661 : NOR2_X1 port map( A1 => n21484, A2 => n21880, ZN => n36780);
   U2673 : AND2_X1 port map( A1 => n1454, A2 => n1206, Z => n33981);
   U2681 : INV_X2 port map( I => n19658, ZN => n24373);
   U2685 : BUF_X2 port map( I => n8219, Z => n7866);
   U2687 : NAND2_X2 port map( A1 => n19573, A2 => n4292, ZN => n35454);
   U2691 : INV_X2 port map( I => n27882, ZN => n28255);
   U2704 : NAND2_X2 port map( A1 => n36685, A2 => n28677, ZN => n28577);
   U2708 : NAND2_X2 port map( A1 => n6075, A2 => n6077, ZN => n32870);
   U2711 : BUF_X4 port map( I => n37378, Z => n31626);
   U2713 : INV_X2 port map( I => n24759, ZN => n14265);
   U2722 : NOR2_X2 port map( A1 => n21583, A2 => n21893, ZN => n21514);
   U2724 : OAI22_X2 port map( A1 => n36673, A2 => n1578, B1 => n31213, B2 => 
                           n24799, ZN => n8576);
   U2726 : OR2_X1 port map( A1 => n33840, A2 => n14477, Z => n2682);
   U2741 : OAI21_X1 port map( A1 => n37783, A2 => n8149, B => n28089, ZN => 
                           n5403);
   U2758 : INV_X2 port map( I => n13151, ZN => n1417);
   U2772 : AND2_X1 port map( A1 => n8413, A2 => n11636, Z => n11651);
   U2783 : NAND2_X1 port map( A1 => n36348, A2 => n27974, ZN => n27978);
   U2793 : AOI21_X1 port map( A1 => n13081, A2 => n28273, B => n10642, ZN => 
                           n36348);
   U2794 : AOI21_X1 port map( A1 => n29219, A2 => n31772, B => n32209, ZN => 
                           n122);
   U2803 : NAND2_X1 port map( A1 => n6019, A2 => n9918, ZN => n16490);
   U2811 : NAND3_X1 port map( A1 => n18883, A2 => n28591, A3 => n306, ZN => 
                           n15629);
   U2837 : NAND2_X1 port map( A1 => n20274, A2 => n36421, ZN => n36420);
   U2841 : NAND3_X1 port map( A1 => n31120, A2 => n3818, A3 => n30076, ZN => 
                           n34292);
   U2848 : NOR2_X1 port map( A1 => n34592, A2 => n7637, ZN => n9967);
   U2849 : NAND2_X1 port map( A1 => n19884, A2 => n16874, ZN => n29181);
   U2856 : OAI21_X1 port map( A1 => n22149, A2 => n5821, B => n18999, ZN => 
                           n9124);
   U2860 : AOI22_X1 port map( A1 => n32457, A2 => n8071, B1 => n20376, B2 => 
                           n1154, ZN => n7212);
   U2861 : OR2_X1 port map( A1 => n29884, A2 => n29883, Z => n14540);
   U2865 : NAND2_X1 port map( A1 => n8089, A2 => n14323, ZN => n13616);
   U2868 : NOR2_X1 port map( A1 => n20572, A2 => n38365, ZN => n33725);
   U2870 : NOR2_X1 port map( A1 => n38365, A2 => n20572, ZN => n18013);
   U2874 : OAI21_X1 port map( A1 => n15922, A2 => n20572, B => n11166, ZN => 
                           n11368);
   U2882 : NOR2_X1 port map( A1 => n37040, A2 => n12685, ZN => n14588);
   U2887 : NAND2_X1 port map( A1 => n29635, A2 => n20290, ZN => n20286);
   U2892 : NAND2_X1 port map( A1 => n6001, A2 => n31772, ZN => n36977);
   U2905 : NAND3_X1 port map( A1 => n3818, A2 => n31120, A3 => n30077, ZN => 
                           n30072);
   U2913 : NAND3_X1 port map( A1 => n28723, A2 => n28724, A3 => n28722, ZN => 
                           n18187);
   U2957 : INV_X2 port map( I => n20159, ZN => n29409);
   U2958 : CLKBUF_X2 port map( I => n20159, Z => n9790);
   U2962 : INV_X2 port map( I => n13545, ZN => n2803);
   U2972 : NOR3_X1 port map( A1 => n13446, A2 => n19007, A3 => n24403, ZN => 
                           n7084);
   U2973 : NAND2_X1 port map( A1 => n13446, A2 => n13555, ZN => n34598);
   U2975 : AOI22_X1 port map( A1 => n29400, A2 => n13850, B1 => n17849, B2 => 
                           n16260, ZN => n29414);
   U2982 : NOR2_X1 port map( A1 => n25481, A2 => n32026, ZN => n25526);
   U2984 : NOR2_X1 port map( A1 => n27887, A2 => n1454, ZN => n33913);
   U2986 : NOR2_X1 port map( A1 => n2989, A2 => n11361, ZN => n3336);
   U2998 : NAND2_X1 port map( A1 => n26780, A2 => n20223, ZN => n32743);
   U3001 : NAND2_X1 port map( A1 => n26780, A2 => n17712, ZN => n35410);
   U3009 : CLKBUF_X4 port map( I => n23682, Z => n1607);
   U3010 : NOR2_X1 port map( A1 => n30003, A2 => n35103, ZN => n35588);
   U3011 : AND2_X1 port map( A1 => n19844, A2 => n28713, Z => n8218);
   U3028 : NOR2_X1 port map( A1 => n20274, A2 => n4768, ZN => n34707);
   U3029 : NAND2_X1 port map( A1 => n5270, A2 => n30032, ZN => n30039);
   U3030 : OAI21_X1 port map( A1 => n19458, A2 => n30042, B => n30041, ZN => 
                           n19884);
   U3033 : AOI21_X1 port map( A1 => n24779, A2 => n16210, B => n30421, ZN => 
                           n3016);
   U3071 : NAND2_X1 port map( A1 => n26578, A2 => n26564, ZN => n26580);
   U3085 : NOR2_X1 port map( A1 => n16889, A2 => n31532, ZN => n12370);
   U3102 : AOI21_X1 port map( A1 => n13014, A2 => n11981, B => n29209, ZN => 
                           n34592);
   U3108 : OR2_X1 port map( A1 => n1404, A2 => n29592, Z => n14433);
   U3118 : INV_X2 port map( I => n4945, ZN => n27979);
   U3137 : NOR2_X1 port map( A1 => n9751, A2 => n20359, ZN => n14619);
   U3143 : NOR2_X1 port map( A1 => n12829, A2 => n12876, ZN => n29383);
   U3144 : NAND3_X1 port map( A1 => n10422, A2 => n12876, A3 => n29310, ZN => 
                           n29079);
   U3167 : NAND2_X1 port map( A1 => n29367, A2 => n37095, ZN => n19060);
   U3173 : NAND2_X1 port map( A1 => n30117, A2 => n18829, ZN => n12203);
   U3179 : OAI21_X1 port map( A1 => n259, A2 => n33012, B => n11081, ZN => 
                           n11054);
   U3184 : NOR2_X1 port map( A1 => n11081, A2 => n17986, ZN => n11053);
   U3185 : NAND2_X1 port map( A1 => n24826, A2 => n11081, ZN => n14519);
   U3189 : NAND2_X1 port map( A1 => n18743, A2 => n35051, ZN => n12189);
   U3194 : NOR2_X1 port map( A1 => n31557, A2 => n25689, ZN => n36309);
   U3202 : NOR2_X1 port map( A1 => n31557, A2 => n6448, ZN => n25686);
   U3206 : NAND3_X1 port map( A1 => n15038, A2 => n11628, A3 => n12218, ZN => 
                           n27620);
   U3215 : NOR2_X1 port map( A1 => n28012, A2 => n11628, ZN => n15269);
   U3219 : OAI21_X1 port map( A1 => n30128, A2 => n1385, B => n10813, ZN => 
                           n13298);
   U3221 : NAND2_X1 port map( A1 => n1407, A2 => n31444, ZN => n6202);
   U3231 : NOR2_X1 port map( A1 => n1061, A2 => n14179, ZN => n11410);
   U3235 : NAND2_X1 port map( A1 => n9242, A2 => n20010, ZN => n28150);
   U3250 : NOR2_X1 port map( A1 => n14783, A2 => n20277, ZN => n21472);
   U3255 : INV_X1 port map( I => n8605, ZN => n14970);
   U3263 : NOR2_X1 port map( A1 => n12717, A2 => n12718, ZN => n33337);
   U3268 : INV_X1 port map( I => n19096, ZN => n12442);
   U3273 : AOI21_X1 port map( A1 => n2050, A2 => n14640, B => n28222, ZN => 
                           n436);
   U3280 : OAI22_X1 port map( A1 => n16213, A2 => n21051, B1 => n7939, B2 => 
                           n23379, ZN => n15969);
   U3281 : INV_X1 port map( I => n16213, ZN => n35974);
   U3283 : CLKBUF_X1 port map( I => n18908, Z => n34847);
   U3285 : OR2_X1 port map( A1 => n25483, A2 => n25328, Z => n18787);
   U3335 : AND2_X1 port map( A1 => n19398, A2 => n25681, Z => n30392);
   U3336 : BUF_X2 port map( I => n25395, Z => n25681);
   U3339 : AOI21_X1 port map( A1 => n31120, A2 => n30069, B => n3815, ZN => 
                           n19551);
   U3340 : NAND2_X1 port map( A1 => n20535, A2 => n21869, ZN => n9592);
   U3341 : NAND2_X1 port map( A1 => n13594, A2 => n28680, ZN => n28719);
   U3369 : NAND2_X1 port map( A1 => n36996, A2 => n23165, ZN => n22810);
   U3383 : NOR2_X1 port map( A1 => n24473, A2 => n39074, ZN => n24471);
   U3386 : AOI21_X1 port map( A1 => n31494, A2 => n30484, B => n288, ZN => 
                           n5158);
   U3397 : NAND2_X1 port map( A1 => n19366, A2 => n27969, ZN => n18439);
   U3406 : NAND2_X1 port map( A1 => n28048, A2 => n28255, ZN => n34949);
   U3413 : NOR2_X1 port map( A1 => n15518, A2 => n17477, ZN => n36591);
   U3415 : INV_X1 port map( I => n15267, ZN => n34618);
   U3430 : NOR3_X1 port map( A1 => n5001, A2 => n21023, A3 => n8762, ZN => 
                           n19747);
   U3435 : NAND3_X1 port map( A1 => n32527, A2 => n15825, A3 => n31502, ZN => 
                           n35436);
   U3445 : NOR3_X1 port map( A1 => n31444, A2 => n14158, A3 => n19424, ZN => 
                           n10605);
   U3449 : OR3_X2 port map( A1 => n987, A2 => n1070, A3 => n7872, Z => n16632);
   U3477 : INV_X2 port map( I => n29700, ZN => n1060);
   U3478 : AOI21_X1 port map( A1 => n1182, A2 => n5977, B => n29700, ZN => 
                           n20816);
   U3480 : CLKBUF_X2 port map( I => n29865, Z => n33256);
   U3504 : AOI22_X1 port map( A1 => n1398, A2 => n29701, B1 => n8941, B2 => 
                           n5977, ZN => n8347);
   U3510 : NAND2_X1 port map( A1 => n29430, A2 => n38051, ZN => n29342);
   U3517 : NOR2_X1 port map( A1 => n9677, A2 => n903, ZN => n3410);
   U3518 : NAND2_X1 port map( A1 => n35528, A2 => n9677, ZN => n32916);
   U3521 : NOR2_X1 port map( A1 => n9677, A2 => n19788, ZN => n13774);
   U3531 : INV_X1 port map( I => n30054, ZN => n31296);
   U3534 : NAND3_X1 port map( A1 => n30054, A2 => n30053, A3 => n16468, ZN => 
                           n20169);
   U3551 : NOR3_X1 port map( A1 => n28222, A2 => n18841, A3 => n16065, ZN => 
                           n35368);
   U3556 : OAI22_X1 port map( A1 => n10803, A2 => n29222, B1 => n31772, B2 => 
                           n6002, ZN => n12691);
   U3572 : NOR2_X1 port map( A1 => n22245, A2 => n7046, ZN => n22034);
   U3573 : NAND2_X1 port map( A1 => n22245, A2 => n20889, ZN => n22035);
   U3588 : NAND3_X1 port map( A1 => n26234, A2 => n26066, A3 => n26067, ZN => 
                           n8248);
   U3594 : NOR2_X1 port map( A1 => n9020, A2 => n24309, ZN => n13547);
   U3597 : OR2_X1 port map( A1 => n29532, A2 => n29531, Z => n17104);
   U3615 : NAND3_X1 port map( A1 => n2348, A2 => n1285, A3 => n14379, ZN => 
                           n12202);
   U3624 : AND2_X1 port map( A1 => n33086, A2 => n14139, Z => n34090);
   U3627 : AOI22_X1 port map( A1 => n35526, A2 => n33086, B1 => n22263, B2 => 
                           n22262, ZN => n14252);
   U3637 : AOI21_X1 port map( A1 => n28615, A2 => n13379, B => n37204, ZN => 
                           n28455);
   U3639 : NOR3_X1 port map( A1 => n28453, A2 => n13379, A3 => n180, ZN => 
                           n2573);
   U3644 : NOR2_X1 port map( A1 => n12626, A2 => n34777, ZN => n18124);
   U3673 : NAND2_X1 port map( A1 => n31263, A2 => n37502, ZN => n9961);
   U3677 : NAND2_X1 port map( A1 => n28578, A2 => n28591, ZN => n34670);
   U3683 : NAND3_X1 port map( A1 => n585, A2 => n1605, A3 => n33450, ZN => 
                           n1875);
   U3692 : NOR2_X1 port map( A1 => n36385, A2 => n24866, ZN => n8315);
   U3703 : NAND2_X1 port map( A1 => n26695, A2 => n10524, ZN => n26699);
   U3730 : NAND2_X1 port map( A1 => n13642, A2 => n21094, ZN => n10123);
   U3731 : AOI22_X1 port map( A1 => n13642, A2 => n11582, B1 => n38986, B2 => 
                           n2658, ZN => n14066);
   U3734 : INV_X1 port map( I => n13642, ZN => n34185);
   U3736 : INV_X1 port map( I => n19680, ZN => n22129);
   U3738 : INV_X1 port map( I => n21291, ZN => n21094);
   U3739 : NOR2_X1 port map( A1 => n22161, A2 => n6576, ZN => n36188);
   U3740 : NAND2_X1 port map( A1 => n17066, A2 => n24382, ZN => n16375);
   U3760 : NOR2_X1 port map( A1 => n32537, A2 => n13124, ZN => n33969);
   U3771 : INV_X2 port map( I => n17918, ZN => n19945);
   U3772 : AND2_X1 port map( A1 => n35955, A2 => n30326, Z => n33973);
   U3778 : INV_X1 port map( I => n38173, ZN => n1641);
   U3789 : INV_X2 port map( I => n8069, ZN => n32450);
   U3795 : AND2_X1 port map( A1 => n25484, A2 => n36162, Z => n33976);
   U3809 : BUF_X4 port map( I => n38416, Z => n3356);
   U3810 : INV_X4 port map( I => n3343, ZN => n34265);
   U3814 : AND3_X1 port map( A1 => n25931, A2 => n37378, A3 => n26135, Z => 
                           n33978);
   U3818 : NAND2_X2 port map( A1 => n6075, A2 => n6077, ZN => n35228);
   U3825 : OR2_X1 port map( A1 => n5675, A2 => n32191, Z => n33979);
   U3827 : INV_X2 port map( I => n28179, ZN => n36573);
   U3848 : AOI21_X2 port map( A1 => n30786, A2 => n28311, B => n30785, ZN => 
                           n35249);
   U3854 : NAND2_X1 port map( A1 => n28355, A2 => n28611, ZN => n28358);
   U3864 : AND3_X1 port map( A1 => n19886, A2 => n12159, A3 => n36296, Z => 
                           n30410);
   U3865 : INV_X1 port map( I => n28186, ZN => n15597);
   U3867 : AOI21_X1 port map( A1 => n37209, A2 => n38724, B => n11168, ZN => 
                           n11167);
   U3870 : NAND2_X1 port map( A1 => n38244, A2 => n38724, ZN => n22822);
   U3876 : CLKBUF_X12 port map( I => n31558, Z => n33817);
   U3886 : NAND2_X1 port map( A1 => n3059, A2 => n31287, ZN => n31744);
   U3889 : AOI21_X1 port map( A1 => n35004, A2 => n7883, B => n24314, ZN => 
                           n7036);
   U3891 : OAI21_X1 port map( A1 => n11512, A2 => n17447, B => n28128, ZN => 
                           n14118);
   U3901 : OR2_X2 port map( A1 => n8824, A2 => n35233, Z => n8825);
   U3903 : AOI21_X1 port map( A1 => n1205, A2 => n5352, B => n984, ZN => n13251
                           );
   U3912 : NAND2_X1 port map( A1 => n37378, A2 => n18142, ZN => n11888);
   U3925 : AOI22_X1 port map( A1 => n4195, A2 => n17217, B1 => n36480, B2 => 
                           n4194, ZN => n4193);
   U3926 : NAND2_X1 port map( A1 => n15411, A2 => n17217, ZN => n9060);
   U3932 : NOR2_X1 port map( A1 => n23484, A2 => n6303, ZN => n16716);
   U3951 : AOI21_X1 port map( A1 => n924, A2 => n19449, B => n1006, ZN => n9099
                           );
   U3965 : NAND2_X1 port map( A1 => n27180, A2 => n6686, ZN => n7231);
   U3968 : INV_X1 port map( I => n6686, ZN => n36569);
   U3994 : NAND2_X1 port map( A1 => n9956, A2 => n4353, ZN => n2306);
   U4000 : INV_X1 port map( I => n25395, ZN => n25429);
   U4003 : INV_X1 port map( I => n24753, ZN => n24126);
   U4006 : NOR2_X2 port map( A1 => n24404, A2 => n13904, ZN => n13412);
   U4009 : INV_X2 port map( I => n16619, ZN => n28653);
   U4019 : NAND2_X1 port map( A1 => n2292, A2 => n26961, ZN => n26962);
   U4020 : INV_X2 port map( I => n26961, ZN => n4211);
   U4038 : INV_X1 port map( I => n24933, ZN => n9324);
   U4051 : NAND2_X1 port map( A1 => n26131, A2 => n9916, ZN => n20771);
   U4092 : CLKBUF_X1 port map( I => n24761, Z => n34458);
   U4109 : INV_X1 port map( I => n22517, ZN => n36265);
   U4113 : INV_X1 port map( I => n22620, ZN => n22724);
   U4117 : AND2_X2 port map( A1 => n26668, A2 => n19867, Z => n14922);
   U4145 : BUF_X4 port map( I => n22767, Z => n33990);
   U4148 : INV_X2 port map( I => n21150, ZN => n19637);
   U4163 : NOR3_X1 port map( A1 => n9379, A2 => n33440, A3 => n5753, ZN => 
                           n7111);
   U4169 : AOI22_X1 port map( A1 => n21991, A2 => n22264, B1 => n22262, B2 => 
                           n22261, ZN => n21992);
   U4180 : CLKBUF_X12 port map( I => n15261, Z => n35248);
   U4182 : AOI21_X1 port map( A1 => n38487, A2 => n24381, B => n7210, ZN => 
                           n24386);
   U4184 : NAND3_X2 port map( A1 => n11328, A2 => n35567, A3 => n19586, ZN => 
                           n7683);
   U4187 : NOR2_X1 port map( A1 => n26041, A2 => n8407, ZN => n25869);
   U4191 : NOR2_X1 port map( A1 => n22154, A2 => n9824, ZN => n35194);
   U4192 : NAND3_X1 port map( A1 => n12814, A2 => n9824, A3 => n12793, ZN => 
                           n6200);
   U4202 : NAND2_X1 port map( A1 => n9824, A2 => n3863, ZN => n22271);
   U4214 : AND3_X2 port map( A1 => n1574, A2 => n24806, A3 => n7552, Z => 
                           n18541);
   U4216 : INV_X2 port map( I => n7552, ZN => n957);
   U4231 : OAI21_X1 port map( A1 => n1643, A2 => n17017, B => n23569, ZN => 
                           n23217);
   U4242 : AND2_X2 port map( A1 => n23132, A2 => n22674, Z => n36783);
   U4262 : OAI22_X1 port map( A1 => n6451, A2 => n33860, B1 => n22177, B2 => 
                           n17118, ZN => n36466);
   U4269 : AND2_X2 port map( A1 => n35859, A2 => n13745, Z => n23085);
   U4272 : CLKBUF_X1 port map( I => n9876, Z => n35685);
   U4273 : NAND2_X1 port map( A1 => n22341, A2 => n9876, ZN => n36176);
   U4274 : NOR2_X1 port map( A1 => n22228, A2 => n22229, ZN => n34256);
   U4300 : AND2_X2 port map( A1 => n13572, A2 => n37218, Z => n7575);
   U4301 : NAND2_X1 port map( A1 => n35855, A2 => n7901, ZN => n25933);
   U4308 : INV_X1 port map( I => n10792, ZN => n6461);
   U4313 : NAND2_X1 port map( A1 => n11081, A2 => n24817, ZN => n24527);
   U4335 : NOR2_X1 port map( A1 => n38996, A2 => n17032, ZN => n34441);
   U4382 : NAND2_X1 port map( A1 => n13872, A2 => n25631, ZN => n5100);
   U4402 : INV_X1 port map( I => n23963, ZN => n1622);
   U4418 : NOR2_X1 port map( A1 => n11834, A2 => n9413, ZN => n11833);
   U4423 : CLKBUF_X12 port map( I => n33645, Z => n32003);
   U4429 : CLKBUF_X12 port map( I => n19658, Z => n19415);
   U4431 : BUF_X4 port map( I => n3900, Z => n33995);
   U4434 : OR2_X2 port map( A1 => n5871, A2 => n31679, Z => n18509);
   U4440 : NAND3_X1 port map( A1 => n4192, A2 => n32926, A3 => n32566, ZN => 
                           n4014);
   U4451 : NAND2_X1 port map( A1 => n4232, A2 => n36827, ZN => n10543);
   U4452 : NAND2_X2 port map( A1 => n22326, A2 => n9165, ZN => n22328);
   U4484 : INV_X1 port map( I => n5929, ZN => n8204);
   U4491 : NOR2_X1 port map( A1 => n20494, A2 => n39423, ZN => n20495);
   U4524 : NAND2_X1 port map( A1 => n18044, A2 => n28089, ZN => n32182);
   U4529 : NAND2_X1 port map( A1 => n33656, A2 => n28089, ZN => n8326);
   U4535 : OR2_X2 port map( A1 => n10379, A2 => n10375, Z => n11913);
   U4538 : INV_X1 port map( I => n24070, ZN => n19646);
   U4549 : NAND2_X1 port map( A1 => n27098, A2 => n8412, ZN => n13896);
   U4569 : NOR3_X1 port map( A1 => n378, A2 => n1106, A3 => n36226, ZN => n195)
                           ;
   U4591 : OAI22_X1 port map( A1 => n37213, A2 => n17624, B1 => n25866, B2 => 
                           n35207, ZN => n30656);
   U4606 : INV_X1 port map( I => n9757, ZN => n1462);
   U4615 : INV_X1 port map( I => n15540, ZN => n32286);
   U4616 : NOR2_X1 port map( A1 => n31418, A2 => n15540, ZN => n36835);
   U4625 : INV_X1 port map( I => n16445, ZN => n4986);
   U4641 : NOR2_X1 port map( A1 => n25933, A2 => n38168, ZN => n17954);
   U4643 : OR2_X2 port map( A1 => n3092, A2 => n17095, Z => n20419);
   U4650 : NAND3_X1 port map( A1 => n33871, A2 => n25999, A3 => n9833, ZN => 
                           n17994);
   U4673 : NAND2_X1 port map( A1 => n26, A2 => n22317, ZN => n18372);
   U4675 : INV_X1 port map( I => n22317, ZN => n1679);
   U4676 : INV_X1 port map( I => n384, ZN => n5405);
   U4682 : NOR2_X1 port map( A1 => n15573, A2 => n33046, ZN => n35789);
   U4690 : AOI21_X1 port map( A1 => n19351, A2 => n1645, B => n23124, ZN => 
                           n23022);
   U4714 : NOR2_X1 port map( A1 => n25769, A2 => n25943, ZN => n6579);
   U4744 : INV_X1 port map( I => n35138, ZN => n35098);
   U4759 : INV_X1 port map( I => n26092, ZN => n25945);
   U4794 : NAND3_X1 port map( A1 => n29266, A2 => n20026, A3 => n29384, ZN => 
                           n30863);
   U4795 : AOI22_X1 port map( A1 => n20099, A2 => n13559, B1 => n30087, B2 => 
                           n30093, ZN => n36699);
   U4796 : NAND2_X1 port map( A1 => n11940, A2 => n31534, ZN => n34621);
   U4823 : CLKBUF_X2 port map( I => n29768, Z => n10096);
   U4829 : INV_X1 port map( I => n28380, ZN => n34638);
   U4830 : INV_X1 port map( I => n28679, ZN => n34286);
   U4842 : CLKBUF_X2 port map( I => n16778, Z => n34459);
   U4851 : INV_X2 port map( I => n28656, ZN => n28617);
   U4853 : NOR2_X1 port map( A1 => n36029, A2 => n10393, ZN => n36478);
   U4861 : AOI21_X1 port map( A1 => n14361, A2 => n9089, B => n156, ZN => 
                           n34212);
   U4867 : CLKBUF_X1 port map( I => n32474, Z => n34410);
   U4896 : INV_X1 port map( I => n35617, ZN => n34770);
   U4907 : CLKBUF_X1 port map( I => n27424, Z => n35897);
   U4914 : CLKBUF_X2 port map( I => n12485, Z => n36159);
   U4951 : CLKBUF_X2 port map( I => n9899, Z => n36078);
   U4962 : AND2_X1 port map( A1 => n30883, A2 => n25978, Z => n25979);
   U4967 : NAND2_X1 port map( A1 => n34745, A2 => n5126, ZN => n34743);
   U4993 : CLKBUF_X2 port map( I => n34692, Z => n34485);
   U4997 : BUF_X2 port map( I => n5859, Z => n33348);
   U5010 : NAND2_X1 port map( A1 => n15791, A2 => n34076, ZN => n13743);
   U5014 : NAND2_X1 port map( A1 => n12866, A2 => n34027, ZN => n20337);
   U5035 : OR2_X1 port map( A1 => n25637, A2 => n25716, Z => n34027);
   U5057 : CLKBUF_X2 port map( I => n25581, Z => n36794);
   U5058 : INV_X1 port map( I => n25290, ZN => n35894);
   U5061 : OAI21_X1 port map( A1 => n24793, A2 => n35981, B => n35519, ZN => 
                           n24647);
   U5064 : INV_X1 port map( I => n24869, ZN => n36821);
   U5071 : NAND2_X1 port map( A1 => n35521, A2 => n35520, ZN => n35519);
   U5073 : INV_X1 port map( I => n35952, ZN => n34694);
   U5075 : INV_X2 port map( I => n24745, ZN => n16999);
   U5116 : BUF_X4 port map( I => n13045, Z => n34526);
   U5173 : OR2_X1 port map( A1 => n38886, A2 => n1129, Z => n34077);
   U5214 : CLKBUF_X4 port map( I => n12822, Z => n36701);
   U5263 : INV_X1 port map( I => n22836, ZN => n34726);
   U5265 : INV_X1 port map( I => n12245, ZN => n34772);
   U5272 : NOR2_X1 port map( A1 => n8197, A2 => n31183, ZN => n34727);
   U5275 : CLKBUF_X1 port map( I => n10375, Z => n34190);
   U5297 : BUF_X4 port map( I => n22085, Z => n36006);
   U5299 : AOI21_X1 port map( A1 => n21947, A2 => n32123, B => n21946, ZN => 
                           n21953);
   U5303 : INV_X1 port map( I => n19780, ZN => n34017);
   U5306 : BUF_X2 port map( I => Key(145), Z => n19738);
   U5308 : OAI21_X1 port map( A1 => n30089, A2 => n1380, B => n36699, ZN => 
                           n30091);
   U5328 : NAND3_X1 port map( A1 => n29559, A2 => n6252, A3 => n35176, ZN => 
                           n35141);
   U5333 : NAND2_X1 port map( A1 => n32865, A2 => n30260, ZN => n36674);
   U5338 : INV_X1 port map( I => n3378, ZN => n36676);
   U5344 : NOR2_X1 port map( A1 => n36268, A2 => n34082, ZN => n36172);
   U5351 : AND2_X1 port map( A1 => n29531, A2 => n29535, Z => n9636);
   U5361 : NAND2_X1 port map( A1 => n20433, A2 => n21023, ZN => n36126);
   U5366 : NAND2_X1 port map( A1 => n29079, A2 => n18457, ZN => n36997);
   U5367 : NAND2_X1 port map( A1 => n29214, A2 => n10628, ZN => n36694);
   U5377 : BUF_X2 port map( I => n16388, Z => n5977);
   U5380 : OR2_X1 port map( A1 => n16599, A2 => n16388, Z => n29698);
   U5394 : INV_X1 port map( I => n29500, ZN => n14873);
   U5397 : CLKBUF_X2 port map( I => n29943, Z => n36166);
   U5431 : INV_X1 port map( I => n36742, ZN => n30292);
   U5445 : INV_X1 port map( I => n28604, ZN => n36248);
   U5448 : AND2_X1 port map( A1 => n19893, A2 => n28484, Z => n34047);
   U5452 : NAND2_X1 port map( A1 => n2469, A2 => n19759, ZN => n35805);
   U5463 : INV_X1 port map( I => n10680, ZN => n34462);
   U5470 : CLKBUF_X1 port map( I => n13690, Z => n36165);
   U5493 : NAND2_X1 port map( A1 => n30293, A2 => n12531, ZN => n36525);
   U5495 : NOR2_X1 port map( A1 => n28164, A2 => n7690, ZN => n34596);
   U5506 : INV_X1 port map( I => n34212, ZN => n4978);
   U5511 : INV_X1 port map( I => n4155, ZN => n28126);
   U5517 : NOR2_X1 port map( A1 => n35469, A2 => n9242, ZN => n27622);
   U5527 : BUF_X2 port map( I => n7828, Z => n5469);
   U5528 : CLKBUF_X2 port map( I => n13332, Z => n36877);
   U5530 : BUF_X4 port map( I => n8057, Z => n34008);
   U5532 : INV_X1 port map( I => n32581, ZN => n34313);
   U5535 : INV_X4 port map( I => n6847, ZN => n900);
   U5536 : INV_X1 port map( I => n11487, ZN => n11486);
   U5542 : NAND2_X1 port map( A1 => n35107, A2 => n36679, ZN => n27356);
   U5545 : NAND2_X1 port map( A1 => n2563, A2 => n35730, ZN => n35729);
   U5559 : INV_X1 port map( I => n30542, ZN => n34889);
   U5563 : NAND2_X1 port map( A1 => n27353, A2 => n7291, ZN => n35107);
   U5571 : AND2_X1 port map( A1 => n1481, A2 => n7716, Z => n34114);
   U5572 : NAND2_X1 port map( A1 => n19300, A2 => n36073, ZN => n27057);
   U5574 : NOR2_X1 port map( A1 => n35258, A2 => n13266, ZN => n13268);
   U5579 : BUF_X4 port map( I => n5218, Z => n34562);
   U5589 : NAND2_X1 port map( A1 => n11765, A2 => n27449, ZN => n34704);
   U5595 : CLKBUF_X1 port map( I => n13278, Z => n35473);
   U5613 : NOR2_X1 port map( A1 => n15616, A2 => n36984, ZN => n26140);
   U5623 : BUF_X2 port map( I => n2722, Z => n34853);
   U5633 : OAI21_X1 port map( A1 => n26895, A2 => n16222, B => n16221, ZN => 
                           n16220);
   U5635 : NAND2_X1 port map( A1 => n34003, A2 => n35410, ZN => n35409);
   U5638 : AND2_X1 port map( A1 => n8556, A2 => n20936, Z => n34034);
   U5646 : OAI21_X2 port map( A1 => n14485, A2 => n17394, B => n26933, ZN => 
                           n17393);
   U5650 : AND2_X1 port map( A1 => n26707, A2 => n19951, Z => n32348);
   U5663 : CLKBUF_X1 port map( I => n740, Z => n35259);
   U5676 : INV_X1 port map( I => n26490, ZN => n35637);
   U5679 : INV_X1 port map( I => n26233, ZN => n35471);
   U5685 : INV_X1 port map( I => n26166, ZN => n35639);
   U5694 : CLKBUF_X2 port map( I => n6130, Z => n36544);
   U5717 : NOR2_X1 port map( A1 => n4553, A2 => n34265, ZN => n14564);
   U5723 : AOI21_X1 port map( A1 => n26071, A2 => n11858, B => n36896, ZN => 
                           n36900);
   U5730 : NAND2_X1 port map( A1 => n25970, A2 => n39015, ZN => n34645);
   U5735 : NAND2_X1 port map( A1 => n26058, A2 => n33293, ZN => n36658);
   U5756 : CLKBUF_X4 port map( I => n8375, Z => n36404);
   U5762 : BUF_X2 port map( I => n14212, Z => n30937);
   U5774 : NAND2_X1 port map( A1 => n36324, A2 => n35632, ZN => n36163);
   U5775 : OAI21_X1 port map( A1 => n611, A2 => n32904, B => n36142, ZN => 
                           n7488);
   U5803 : INV_X1 port map( I => n25068, ZN => n36324);
   U5805 : AND2_X1 port map( A1 => n6300, A2 => n9526, Z => n34083);
   U5836 : BUF_X2 port map( I => n25481, Z => n36083);
   U5848 : CLKBUF_X4 port map( I => n21031, Z => n20052);
   U5856 : CLKBUF_X2 port map( I => n36075, Z => n35996);
   U5859 : CLKBUF_X2 port map( I => n35900, Z => n35053);
   U5865 : CLKBUF_X2 port map( I => n25040, Z => n35379);
   U5882 : NOR2_X1 port map( A1 => n24539, A2 => n16990, ZN => n35118);
   U5890 : AOI21_X1 port map( A1 => n24786, A2 => n7831, B => n36697, ZN => 
                           n30413);
   U5902 : NAND2_X1 port map( A1 => n14275, A2 => n1565, ZN => n35784);
   U5919 : OAI21_X1 port map( A1 => n34694, A2 => n3697, B => n2231, ZN => 
                           n35886);
   U5920 : NAND2_X1 port map( A1 => n24613, A2 => n37411, ZN => n36697);
   U5921 : NAND2_X1 port map( A1 => n24659, A2 => n19, ZN => n36560);
   U5929 : INV_X1 port map( I => n21018, ZN => n1799);
   U5948 : CLKBUF_X2 port map( I => n24732, Z => n34662);
   U5958 : OAI21_X1 port map( A1 => n17546, A2 => n24467, B => n35774, ZN => 
                           n24323);
   U5968 : BUF_X2 port map( I => n14999, Z => n31684);
   U5975 : NAND2_X1 port map( A1 => n24818, A2 => n24821, ZN => n8647);
   U5980 : INV_X1 port map( I => n24821, ZN => n36180);
   U5993 : NAND2_X1 port map( A1 => n35503, A2 => n34043, ZN => n35056);
   U5998 : INV_X2 port map( I => n8646, ZN => n24824);
   U6003 : CLKBUF_X4 port map( I => n15467, Z => n34011);
   U6004 : OR2_X1 port map( A1 => n10065, A2 => n10439, Z => n36542);
   U6006 : INV_X1 port map( I => n35504, ZN => n35503);
   U6017 : NAND2_X2 port map( A1 => n33743, A2 => n36740, ZN => n30572);
   U6035 : CLKBUF_X2 port map( I => n24247, Z => n19818);
   U6047 : OR2_X1 port map( A1 => n24245, A2 => n24244, Z => n21080);
   U6059 : CLKBUF_X2 port map( I => n16832, Z => n36378);
   U6065 : CLKBUF_X1 port map( I => n24279, Z => n35890);
   U6078 : CLKBUF_X2 port map( I => n24307, Z => n305);
   U6088 : INV_X1 port map( I => n23960, ZN => n36541);
   U6094 : NOR2_X1 port map( A1 => n35812, A2 => n35811, ZN => n11452);
   U6107 : INV_X1 port map( I => n9349, ZN => n35278);
   U6108 : INV_X1 port map( I => n23752, ZN => n35812);
   U6111 : NAND2_X1 port map( A1 => n2274, A2 => n3363, ZN => n23408);
   U6113 : NAND2_X1 port map( A1 => n35007, A2 => n23229, ZN => n21014);
   U6115 : INV_X1 port map( I => n10633, ZN => n35892);
   U6120 : INV_X1 port map( I => n36888, ZN => n23593);
   U6122 : NOR2_X1 port map( A1 => n35068, A2 => n35501, ZN => n13767);
   U6153 : CLKBUF_X4 port map( I => n32366, Z => n36720);
   U6180 : CLKBUF_X2 port map( I => n11342, Z => n35068);
   U6183 : NOR2_X1 port map( A1 => n14429, A2 => n16197, ZN => n32583);
   U6186 : INV_X1 port map( I => n34448, ZN => n14606);
   U6193 : NAND2_X1 port map( A1 => n16198, A2 => n23212, ZN => n34448);
   U6196 : INV_X2 port map( I => n23423, ZN => n34012);
   U6202 : NAND2_X1 port map( A1 => n35806, A2 => n23211, ZN => n20744);
   U6217 : CLKBUF_X2 port map( I => n33934, Z => n35567);
   U6243 : INV_X1 port map( I => n18941, ZN => n35148);
   U6248 : INV_X1 port map( I => n22616, ZN => n34698);
   U6269 : INV_X1 port map( I => n22744, ZN => n33863);
   U6279 : NAND2_X1 port map( A1 => n34023, A2 => n34256, ZN => n12568);
   U6280 : NOR2_X1 port map( A1 => n22069, A2 => n4114, ZN => n36084);
   U6290 : BUF_X2 port map( I => n22150, Z => n31412);
   U6295 : CLKBUF_X2 port map( I => n16880, Z => n34920);
   U6317 : CLKBUF_X4 port map( I => n36214, Z => n35771);
   U6329 : CLKBUF_X1 port map( I => n16265, Z => n35060);
   U6330 : NOR2_X1 port map( A1 => n5733, A2 => n17242, ZN => n3865);
   U6337 : INV_X1 port map( I => n28934, ZN => n35140);
   U6338 : CLKBUF_X2 port map( I => n21428, Z => n35973);
   U6340 : BUF_X4 port map( I => n21518, Z => n34016);
   U6347 : NOR2_X1 port map( A1 => n18293, A2 => n19372, ZN => n37032);
   U6355 : INV_X1 port map( I => n32525, ZN => n35651);
   U6378 : OAI21_X1 port map( A1 => n17948, A2 => n21710, B => n21868, ZN => 
                           n21);
   U6383 : INV_X2 port map( I => n33249, ZN => n2690);
   U6389 : NOR2_X1 port map( A1 => n3484, A2 => n32410, ZN => n34932);
   U6406 : AOI21_X1 port map( A1 => n36781, A2 => n21484, B => n36780, ZN => 
                           n36779);
   U6414 : NAND2_X1 port map( A1 => n10893, A2 => n36490, ZN => n4242);
   U6415 : CLKBUF_X2 port map( I => n21791, Z => n9759);
   U6417 : NAND2_X1 port map( A1 => n17763, A2 => n21707, ZN => n15817);
   U6422 : CLKBUF_X2 port map( I => n21484, Z => n33852);
   U6428 : CLKBUF_X4 port map( I => n21741, Z => n1157);
   U6443 : OAI22_X1 port map( A1 => n21778, A2 => n34922, B1 => n21612, B2 => 
                           n36519, ZN => n21614);
   U6473 : INV_X1 port map( I => n36397, ZN => n10762);
   U6474 : OAI21_X1 port map( A1 => n16536, A2 => n32164, B => n15125, ZN => 
                           n21658);
   U6480 : INV_X1 port map( I => n14139, ZN => n22259);
   U6484 : INV_X1 port map( I => n22341, ZN => n18558);
   U6487 : AOI21_X1 port map( A1 => n21702, A2 => n19709, B => n1353, ZN => 
                           n21703);
   U6490 : AOI21_X1 port map( A1 => n7357, A2 => n20646, B => n20643, ZN => 
                           n35943);
   U6494 : CLKBUF_X4 port map( I => n8899, Z => n4388);
   U6502 : CLKBUF_X1 port map( I => n22250, Z => n34488);
   U6513 : INV_X1 port map( I => n22214, ZN => n22216);
   U6528 : INV_X2 port map( I => n1333, ZN => n17359);
   U6529 : NOR2_X1 port map( A1 => n22160, A2 => n18656, ZN => n14622);
   U6537 : CLKBUF_X2 port map( I => n19373, Z => n36303);
   U6544 : NAND3_X1 port map( A1 => n21845, A2 => n21844, A3 => n21672, ZN => 
                           n21673);
   U6557 : NAND2_X1 port map( A1 => n30828, A2 => n30826, ZN => n35675);
   U6560 : CLKBUF_X2 port map( I => n19515, Z => n34452);
   U6581 : NOR2_X1 port map( A1 => n22399, A2 => n31857, ZN => n8662);
   U6613 : INV_X1 port map( I => n22702, ZN => n22701);
   U6614 : INV_X1 port map( I => n22607, ZN => n35078);
   U6628 : NAND2_X1 port map( A1 => n3273, A2 => n23032, ZN => n23033);
   U6638 : INV_X1 port map( I => n20449, ZN => n22866);
   U6639 : NAND2_X1 port map( A1 => n11582, A2 => n20570, ZN => n4890);
   U6640 : NAND2_X1 port map( A1 => n9954, A2 => n14390, ZN => n23004);
   U6662 : NAND2_X1 port map( A1 => n30594, A2 => n20372, ZN => n3811);
   U6663 : NAND2_X1 port map( A1 => n23013, A2 => n23012, ZN => n5039);
   U6665 : INV_X1 port map( I => n14560, ZN => n23000);
   U6666 : NOR2_X1 port map( A1 => n12925, A2 => n36369, ZN => n36368);
   U6671 : NAND2_X1 port map( A1 => n13734, A2 => n19788, ZN => n22839);
   U6673 : INV_X1 port map( I => n5337, ZN => n15045);
   U6699 : AOI22_X1 port map( A1 => n15885, A2 => n23128, B1 => n19621, B2 => 
                           n34014, ZN => n15884);
   U6700 : NAND2_X1 port map( A1 => n12621, A2 => n36763, ZN => n12620);
   U6702 : NAND3_X1 port map( A1 => n15163, A2 => n22810, A3 => n22809, ZN => 
                           n16731);
   U6708 : NAND2_X1 port map( A1 => n11108, A2 => n23423, ZN => n1893);
   U6716 : NAND2_X1 port map( A1 => n23358, A2 => n30299, ZN => n36035);
   U6724 : NAND2_X1 port map( A1 => n35130, A2 => n23315, ZN => n33638);
   U6742 : NAND2_X1 port map( A1 => n23749, A2 => n9321, ZN => n35007);
   U6768 : OAI21_X1 port map( A1 => n16094, A2 => n15176, B => n35569, ZN => 
                           n36785);
   U6773 : INV_X1 port map( I => n18849, ZN => n13224);
   U6781 : INV_X1 port map( I => n7475, ZN => n7185);
   U6785 : INV_X1 port map( I => n13395, ZN => n23789);
   U6799 : NOR2_X1 port map( A1 => n35253, A2 => n18907, ZN => n31488);
   U6801 : INV_X1 port map( I => n23073, ZN => n34900);
   U6817 : INV_X1 port map( I => n24457, ZN => n2972);
   U6831 : NAND3_X1 port map( A1 => n17711, A2 => n36757, A3 => n17709, ZN => 
                           n17710);
   U6839 : NOR3_X1 port map( A1 => n11361, A2 => n19895, A3 => n24359, ZN => 
                           n23941);
   U6846 : AOI21_X1 port map( A1 => n24087, A2 => n24433, B => n1608, ZN => 
                           n10023);
   U6851 : NAND3_X1 port map( A1 => n1282, A2 => n20404, A3 => n24346, ZN => 
                           n24347);
   U6852 : INV_X1 port map( I => n5955, ZN => n24348);
   U6856 : NOR2_X1 port map( A1 => n14704, A2 => n1283, ZN => n13186);
   U6861 : NAND2_X1 port map( A1 => n17259, A2 => n7240, ZN => n3307);
   U6874 : OAI21_X1 port map( A1 => n12423, A2 => n18920, B => n1594, ZN => 
                           n12422);
   U6875 : OR2_X1 port map( A1 => n7693, A2 => n17087, Z => n34115);
   U6884 : CLKBUF_X2 port map( I => n24492, Z => n36090);
   U6894 : NAND2_X1 port map( A1 => n18324, A2 => n24764, ZN => n18325);
   U6901 : OR2_X1 port map( A1 => n36471, A2 => n2018, Z => n20064);
   U6905 : AOI21_X1 port map( A1 => n11846, A2 => n19828, B => n5957, ZN => 
                           n7930);
   U6919 : NOR3_X1 port map( A1 => n13128, A2 => n2747, A3 => n2731, ZN => 
                           n2730);
   U6922 : NOR2_X1 port map( A1 => n34935, A2 => n34934, ZN => n34821);
   U6931 : INV_X1 port map( I => n38171, ZN => n24978);
   U6939 : NOR3_X1 port map( A1 => n35952, A2 => n3697, A3 => n14999, ZN => 
                           n33945);
   U6953 : NAND2_X1 port map( A1 => n11642, A2 => n31530, ZN => n24882);
   U6977 : CLKBUF_X2 port map( I => n6759, Z => n61);
   U6980 : INV_X1 port map( I => n25225, ZN => n35511);
   U6989 : NOR2_X1 port map( A1 => n4048, A2 => n18734, ZN => n15356);
   U6995 : NOR2_X1 port map( A1 => n36708, A2 => n36707, ZN => n30705);
   U6998 : NAND2_X1 port map( A1 => n33491, A2 => n20515, ZN => n36323);
   U7003 : NAND2_X1 port map( A1 => n36794, A2 => n25390, ZN => n24894);
   U7005 : NAND2_X1 port map( A1 => n1253, A2 => n16677, ZN => n25388);
   U7006 : NOR2_X1 port map( A1 => n15356, A2 => n19637, ZN => n15355);
   U7018 : NAND2_X1 port map( A1 => n1253, A2 => n19941, ZN => n36793);
   U7020 : OR2_X1 port map( A1 => n25261, A2 => n32989, Z => n34103);
   U7029 : NOR2_X1 port map( A1 => n25545, A2 => n25481, ZN => n2247);
   U7032 : OR2_X1 port map( A1 => n25680, A2 => n30633, Z => n7540);
   U7037 : NAND2_X1 port map( A1 => n25402, A2 => n5314, ZN => n18113);
   U7043 : INV_X1 port map( I => n19264, ZN => n12381);
   U7046 : NAND2_X1 port map( A1 => n25547, A2 => n19701, ZN => n18599);
   U7048 : NAND2_X1 port map( A1 => n25416, A2 => n30377, ZN => n14914);
   U7049 : OAI21_X1 port map( A1 => n37049, A2 => n31457, B => n32101, ZN => 
                           n36277);
   U7068 : INV_X1 port map( I => n25111, ZN => n25994);
   U7070 : NAND2_X1 port map( A1 => n1101, A2 => n9380, ZN => n8860);
   U7089 : INV_X2 port map( I => n16250, ZN => n12199);
   U7095 : NAND2_X1 port map( A1 => n34692, A2 => n36532, ZN => n26129);
   U7121 : INV_X1 port map( I => n26340, ZN => n26341);
   U7125 : NOR2_X1 port map( A1 => n37073, A2 => n11858, ZN => n17311);
   U7130 : INV_X1 port map( I => n26601, ZN => n34478);
   U7132 : INV_X1 port map( I => n2594, ZN => n5381);
   U7142 : NAND3_X1 port map( A1 => n13391, A2 => n35744, A3 => n17008, ZN => 
                           n26096);
   U7158 : INV_X1 port map( I => n26492, ZN => n159);
   U7163 : INV_X1 port map( I => n5078, ZN => n35967);
   U7178 : NAND2_X1 port map( A1 => n30942, A2 => n1006, ZN => n4651);
   U7189 : NAND3_X1 port map( A1 => n1088, A2 => n26701, A3 => n26700, ZN => 
                           n26706);
   U7211 : NAND2_X1 port map( A1 => n3449, A2 => n13588, ZN => n31226);
   U7212 : NAND2_X1 port map( A1 => n21277, A2 => n20936, ZN => n2101);
   U7217 : CLKBUF_X4 port map( I => n26747, Z => n15594);
   U7225 : NAND2_X1 port map( A1 => n34003, A2 => n34426, ZN => n26785);
   U7227 : NAND2_X1 port map( A1 => n6190, A2 => n10440, ZN => n35489);
   U7236 : OAI21_X1 port map( A1 => n14412, A2 => n15411, B => n32892, ZN => 
                           n36445);
   U7242 : NOR2_X1 port map( A1 => n26632, A2 => n12755, ZN => n19250);
   U7249 : NAND2_X1 port map( A1 => n862, A2 => n2451, ZN => n26892);
   U7260 : AOI21_X1 port map( A1 => n925, A2 => n1008, B => n15825, ZN => n7007
                           );
   U7264 : INV_X1 port map( I => n26264, ZN => n34228);
   U7273 : NAND2_X1 port map( A1 => n6605, A2 => n5720, ZN => n7585);
   U7276 : NAND3_X1 port map( A1 => n26722, A2 => n16970, A3 => n19225, ZN => 
                           n8685);
   U7299 : NAND2_X1 port map( A1 => n27214, A2 => n11765, ZN => n27093);
   U7337 : INV_X1 port map( I => n27259, ZN => n5365);
   U7348 : AOI21_X1 port map( A1 => n10946, A2 => n27403, B => n35258, ZN => 
                           n31185);
   U7365 : NAND3_X1 port map( A1 => n11805, A2 => n32463, A3 => n38907, ZN => 
                           n576);
   U7368 : AOI22_X1 port map( A1 => n27388, A2 => n14327, B1 => n39826, B2 => 
                           n2761, ZN => n31943);
   U7369 : NAND2_X1 port map( A1 => n34705, A2 => n34704, ZN => n34493);
   U7385 : NAND2_X1 port map( A1 => n27335, A2 => n2035, ZN => n27487);
   U7404 : INV_X1 port map( I => n14808, ZN => n35889);
   U7418 : NAND3_X1 port map( A1 => n1086, A2 => n17166, A3 => n4781, ZN => 
                           n12075);
   U7420 : INV_X1 port map( I => n27707, ZN => n34708);
   U7422 : INV_X1 port map( I => n27678, ZN => n34409);
   U7426 : INV_X1 port map( I => n886, ZN => n36325);
   U7429 : INV_X1 port map( I => n4266, ZN => n35089);
   U7437 : NOR2_X1 port map( A1 => n28194, A2 => n17197, ZN => n27928);
   U7445 : NOR2_X1 port map( A1 => n27970, A2 => n28148, ZN => n19969);
   U7448 : NAND2_X1 port map( A1 => n28114, A2 => n28115, ZN => n3066);
   U7451 : NOR2_X1 port map( A1 => n580, A2 => n39571, ZN => n7223);
   U7458 : NAND2_X1 port map( A1 => n8207, A2 => n1204, ZN => n8327);
   U7472 : NAND2_X1 port map( A1 => n28172, A2 => n28258, ZN => n18192);
   U7477 : OR2_X1 port map( A1 => n28278, A2 => n19995, Z => n27543);
   U7484 : NAND2_X1 port map( A1 => n12260, A2 => n9845, ZN => n13876);
   U7511 : NOR2_X1 port map( A1 => n6819, A2 => n35911, ZN => n3055);
   U7516 : NOR3_X1 port map( A1 => n1195, A2 => n31542, A3 => n8131, ZN => 
                           n32800);
   U7523 : NAND2_X1 port map( A1 => n33046, A2 => n1815, ZN => n28640);
   U7536 : NAND2_X1 port map( A1 => n28409, A2 => n1426, ZN => n28410);
   U7538 : INV_X1 port map( I => n5645, ZN => n31615);
   U7540 : INV_X1 port map( I => n28997, ZN => n1412);
   U7541 : INV_X1 port map( I => n28966, ZN => n15682);
   U7544 : INV_X1 port map( I => n29152, ZN => n36828);
   U7547 : CLKBUF_X2 port map( I => n28840, Z => n7667);
   U7553 : CLKBUF_X2 port map( I => n29381, Z => n32906);
   U7570 : CLKBUF_X1 port map( I => n29769, Z => n28);
   U7578 : NAND2_X1 port map( A1 => n5335, A2 => n1055, ZN => n4790);
   U7583 : NOR2_X1 port map( A1 => n18104, A2 => n29956, ZN => n29905);
   U7584 : OR2_X1 port map( A1 => n20524, A2 => n19224, Z => n30152);
   U7585 : NAND2_X1 port map( A1 => n38051, A2 => n2954, ZN => n29502);
   U7589 : INV_X1 port map( I => n3430, ZN => n35975);
   U7593 : AOI21_X1 port map( A1 => n36550, A2 => n16828, B => n29385, ZN => 
                           n31180);
   U7594 : NAND2_X1 port map( A1 => n28880, A2 => n31511, ZN => n34806);
   U7596 : NAND3_X1 port map( A1 => n29770, A2 => n29843, A3 => n29844, ZN => 
                           n29771);
   U7602 : NAND3_X1 port map( A1 => n30720, A2 => n1757, A3 => n11826, ZN => 
                           n33557);
   U7605 : INV_X1 port map( I => n5530, ZN => n3378);
   U7606 : INV_X1 port map( I => n15841, ZN => n29440);
   U7611 : OAI22_X1 port map( A1 => n29369, A2 => n11067, B1 => n13981, B2 => 
                           n16683, ZN => n13277);
   U7619 : CLKBUF_X2 port map( I => n18257, Z => n32050);
   U7620 : OAI22_X1 port map( A1 => n10942, A2 => n30033, B1 => n30014, B2 => 
                           n15643, ZN => n32531);
   U7623 : INV_X1 port map( I => n30203, ZN => n1050);
   U7624 : AOI22_X1 port map( A1 => n30039, A2 => n35103, B1 => n30036, B2 => 
                           n30037, ZN => n30040);
   U7629 : OR2_X1 port map( A1 => n22282, A2 => n22130, Z => n34019);
   U7631 : XNOR2_X1 port map( A1 => n4441, A2 => n10213, ZN => n34020);
   U7632 : NAND2_X1 port map( A1 => n9737, A2 => n12535, ZN => n34021);
   U7634 : XNOR2_X1 port map( A1 => n15413, A2 => n13356, ZN => n34022);
   U7636 : XNOR2_X1 port map( A1 => n26296, A2 => n26295, ZN => n34024);
   U7644 : AND2_X1 port map( A1 => n34014, A2 => n3273, Z => n34030);
   U7645 : AND2_X1 port map( A1 => n34080, A2 => n959, Z => n34031);
   U7647 : XNOR2_X1 port map( A1 => n25298, A2 => n30101, ZN => n34032);
   U7649 : AND2_X1 port map( A1 => n38163, A2 => n30128, Z => n34033);
   U7654 : OR2_X1 port map( A1 => n33888, A2 => n994, Z => n34037);
   U7657 : XNOR2_X1 port map( A1 => n28931, A2 => n28930, ZN => n34038);
   U7659 : AND2_X1 port map( A1 => n1432, A2 => n8349, Z => n34041);
   U7663 : AND2_X1 port map( A1 => n38317, A2 => n38668, Z => n34042);
   U7667 : OR2_X1 port map( A1 => n38303, A2 => n6849, Z => n34043);
   U7676 : OR2_X1 port map( A1 => n21860, A2 => n19641, Z => n34048);
   U7681 : AND2_X1 port map( A1 => n10120, A2 => n21839, Z => n34049);
   U7683 : XOR2_X1 port map( A1 => n18270, A2 => n32931, Z => n34050);
   U7686 : XNOR2_X1 port map( A1 => n3610, A2 => n19751, ZN => n34052);
   U7688 : XNOR2_X1 port map( A1 => n35376, A2 => n19613, ZN => n34053);
   U7689 : XNOR2_X1 port map( A1 => n13617, A2 => n29371, ZN => n34054);
   U7693 : XNOR2_X1 port map( A1 => n14907, A2 => n1459, ZN => n34056);
   U7694 : AND2_X1 port map( A1 => n32262, A2 => n32261, Z => n34057);
   U7696 : AND2_X1 port map( A1 => n14734, A2 => n14527, Z => n34059);
   U7710 : XNOR2_X1 port map( A1 => n7161, A2 => n7158, ZN => n34062);
   U7715 : AND3_X1 port map( A1 => n26764, A2 => n3606, A3 => n13393, Z => 
                           n34063);
   U7721 : AND2_X1 port map( A1 => n19647, A2 => n668, Z => n34066);
   U7723 : OR2_X1 port map( A1 => n13998, A2 => n13997, Z => n34067);
   U7735 : AND2_X1 port map( A1 => n9954, A2 => n19823, Z => n34072);
   U7739 : INV_X1 port map( I => n8071, ZN => n1339);
   U7740 : BUF_X2 port map( I => n8071, Z => n5821);
   U7757 : AND2_X1 port map( A1 => n25361, A2 => n12896, Z => n34085);
   U7759 : OR2_X2 port map( A1 => n16080, A2 => n14473, Z => n34087);
   U7761 : XNOR2_X1 port map( A1 => n17048, A2 => n33551, ZN => n34088);
   U7766 : OR2_X1 port map( A1 => n29701, A2 => n28414, Z => n34089);
   U7769 : XNOR2_X1 port map( A1 => n25256, A2 => n4556, ZN => n34092);
   U7771 : XNOR2_X1 port map( A1 => n29463, A2 => n27815, ZN => n34094);
   U7776 : XNOR2_X1 port map( A1 => n25229, A2 => n1710, ZN => n34096);
   U7779 : OR2_X1 port map( A1 => n34180, A2 => n29700, Z => n34097);
   U7790 : XNOR2_X1 port map( A1 => n22486, A2 => n22426, ZN => n34104);
   U7793 : AND2_X1 port map( A1 => n30843, A2 => n8264, Z => n34105);
   U7804 : AND2_X1 port map( A1 => n25677, A2 => n19589, Z => n34112);
   U7807 : INV_X1 port map( I => n23792, ZN => n34851);
   U7809 : INV_X1 port map( I => n29474, ZN => n36040);
   U7810 : INV_X1 port map( I => n28807, ZN => n28764);
   U7818 : INV_X1 port map( I => n29732, ZN => n29753);
   U7824 : INV_X1 port map( I => n38217, ZN => n11181);
   U7839 : XNOR2_X1 port map( A1 => Key(189), A2 => Plaintext(189), ZN => 
                           n34122);
   U7859 : AND2_X1 port map( A1 => n3628, A2 => n16967, Z => n34124);
   U7861 : INV_X2 port map( I => n4886, ZN => n27069);
   U7863 : XNOR2_X1 port map( A1 => n14374, A2 => n25193, ZN => n34126);
   U7875 : OR2_X2 port map( A1 => n22100, A2 => n22058, Z => n34128);
   U7884 : AND2_X1 port map( A1 => n23478, A2 => n23479, Z => n34129);
   U7888 : INV_X1 port map( I => n37815, ZN => n23159);
   U7892 : XNOR2_X1 port map( A1 => n7475, A2 => n23880, ZN => n34132);
   U7913 : XNOR2_X1 port map( A1 => n39797, A2 => n29562, ZN => n34135);
   U7916 : XOR2_X1 port map( A1 => n33271, A2 => n25194, Z => n34136);
   U7919 : XNOR2_X1 port map( A1 => n25284, A2 => n25283, ZN => n34137);
   U7935 : XNOR2_X1 port map( A1 => n25006, A2 => n34945, ZN => n34139);
   U7944 : XNOR2_X1 port map( A1 => n25215, A2 => n29857, ZN => n34142);
   U7947 : XNOR2_X1 port map( A1 => n29707, A2 => n7481, ZN => n34144);
   U7950 : XNOR2_X1 port map( A1 => n19729, A2 => n26514, ZN => n34145);
   U7951 : XNOR2_X1 port map( A1 => n24985, A2 => n24984, ZN => n34147);
   U7952 : OR2_X2 port map( A1 => n20491, A2 => n20490, Z => n34148);
   U7953 : XNOR2_X1 port map( A1 => n37498, A2 => n35702, ZN => n34149);
   U7961 : XNOR2_X1 port map( A1 => n8340, A2 => n25853, ZN => n34151);
   U7965 : XNOR2_X1 port map( A1 => n26403, A2 => n15530, ZN => n34152);
   U7967 : AND2_X2 port map( A1 => n31362, A2 => n9833, Z => n34154);
   U7971 : XNOR2_X1 port map( A1 => n37476, A2 => n39559, ZN => n34157);
   U7977 : INV_X1 port map( I => n18135, ZN => n26220);
   U7983 : XNOR2_X1 port map( A1 => n19450, A2 => n19733, ZN => n34161);
   U7984 : INV_X1 port map( I => n7959, ZN => n26702);
   U7988 : XOR2_X1 port map( A1 => n27746, A2 => n19733, Z => n34162);
   U7991 : NOR2_X1 port map( A1 => n1093, A2 => n11334, ZN => n34163);
   U8031 : XNOR2_X1 port map( A1 => n21084, A2 => n30956, ZN => n34175);
   U8035 : XNOR2_X1 port map( A1 => n9786, A2 => n28994, ZN => n34179);
   U8043 : XNOR2_X1 port map( A1 => n29153, A2 => n14195, ZN => n34181);
   U8044 : AND2_X1 port map( A1 => n29755, A2 => n29754, Z => n34182);
   U8045 : XNOR2_X1 port map( A1 => n3941, A2 => n632, ZN => n34183);
   U8050 : NAND2_X1 port map( A1 => n34186, A2 => n5469, ZN => n20306);
   U8076 : NAND2_X2 port map( A1 => n36972, A2 => n28065, ZN => n7429);
   U8080 : NAND2_X1 port map( A1 => n6118, A2 => n6119, ZN => n6117);
   U8086 : NOR2_X2 port map( A1 => n34261, A2 => n25602, ZN => n34260);
   U8087 : NAND2_X1 port map( A1 => n36902, A2 => n26, ZN => n20986);
   U8102 : XOR2_X1 port map( A1 => n20025, A2 => n29072, Z => n4616);
   U8107 : OAI21_X2 port map( A1 => n28317, A2 => n28316, B => n28315, ZN => 
                           n29072);
   U8120 : NOR2_X2 port map( A1 => n20319, A2 => n27879, ZN => n28874);
   U8124 : AOI22_X2 port map( A1 => n34193, A2 => n2603, B1 => n15623, B2 => 
                           n1076, ZN => n15023);
   U8125 : AND2_X1 port map( A1 => n28149, A2 => n2604, Z => n34193);
   U8130 : XOR2_X1 port map( A1 => n25210, A2 => n14214, Z => n5721);
   U8139 : XOR2_X1 port map( A1 => n135, A2 => n34196, Z => n8365);
   U8140 : XOR2_X1 port map( A1 => n6283, A2 => n650, Z => n34196);
   U8141 : AOI21_X2 port map( A1 => n16670, A2 => n16669, B => n34197, ZN => 
                           n16668);
   U8150 : XOR2_X1 port map( A1 => n34178, A2 => n3082, Z => n6316);
   U8158 : BUF_X4 port map( I => n35399, Z => n35290);
   U8159 : OR2_X1 port map( A1 => n12260, A2 => n12257, Z => n12259);
   U8161 : INV_X2 port map( I => n16699, ZN => n36105);
   U8162 : AOI21_X2 port map( A1 => n7058, A2 => n12080, B => n34201, ZN => 
                           n22549);
   U8163 : OAI21_X2 port map( A1 => n12080, A2 => n21865, B => n36680, ZN => 
                           n34201);
   U8166 : XOR2_X1 port map( A1 => n3476, A2 => n34202, Z => n7518);
   U8173 : NOR2_X1 port map( A1 => n38487, A2 => n33314, ZN => n6567);
   U8182 : INV_X1 port map( I => n25302, ZN => n34208);
   U8189 : INV_X2 port map( I => n34203, ZN => n30844);
   U8191 : XOR2_X1 port map( A1 => n3185, A2 => n3186, Z => n34203);
   U8193 : INV_X1 port map( I => n9059, ZN => n34205);
   U8206 : AND2_X1 port map( A1 => n15172, A2 => n11150, Z => n14589);
   U8217 : NAND3_X2 port map( A1 => n14748, A2 => n14747, A3 => n15238, ZN => 
                           n4524);
   U8219 : NAND2_X1 port map( A1 => n37003, A2 => n34521, ZN => n10814);
   U8221 : AOI22_X2 port map( A1 => n16016, A2 => n17102, B1 => n21029, B2 => 
                           n21601, ZN => n16015);
   U8222 : NOR2_X2 port map( A1 => n16302, A2 => n33280, ZN => n16016);
   U8223 : XOR2_X1 port map( A1 => n30632, A2 => n23850, Z => n311);
   U8227 : XOR2_X1 port map( A1 => n34208, A2 => n25329, Z => n34414);
   U8228 : XOR2_X1 port map( A1 => n17908, A2 => n19014, Z => n17907);
   U8241 : NAND3_X2 port map( A1 => n31704, A2 => n30863, A3 => n29353, ZN => 
                           n29367);
   U8268 : XOR2_X1 port map( A1 => n11563, A2 => n34213, Z => n7090);
   U8270 : AND2_X1 port map( A1 => n22229, A2 => n22228, Z => n17145);
   U8275 : NAND2_X1 port map( A1 => n13166, A2 => n34576, ZN => n4726);
   U8280 : XOR2_X1 port map( A1 => n17455, A2 => n26596, Z => n34214);
   U8303 : XOR2_X1 port map( A1 => Plaintext(66), A2 => Key(66), Z => n261);
   U8305 : AOI22_X1 port map( A1 => n29860, A2 => n29859, B1 => n34215, B2 => 
                           n36764, ZN => n2070);
   U8306 : OR2_X1 port map( A1 => n2073, A2 => n2858, Z => n34215);
   U8316 : OAI22_X2 port map( A1 => n21566, A2 => n7183, B1 => n35, B2 => n36, 
                           ZN => n22038);
   U8318 : INV_X2 port map( I => n34218, ZN => n889);
   U8336 : XOR2_X1 port map( A1 => n34221, A2 => n12205, Z => n36831);
   U8337 : XOR2_X1 port map( A1 => n21866, A2 => n13591, Z => n34221);
   U8349 : NOR2_X1 port map( A1 => n29336, A2 => n14858, ZN => n4520);
   U8363 : XOR2_X1 port map( A1 => n9205, A2 => n22618, Z => n12016);
   U8374 : AND2_X1 port map( A1 => n24244, A2 => n9520, Z => n9386);
   U8392 : NOR2_X2 port map( A1 => n20211, A2 => n13757, ZN => n34224);
   U8402 : NAND2_X1 port map( A1 => n15430, A2 => n34225, ZN => n35033);
   U8403 : NAND2_X1 port map( A1 => n30811, A2 => n34226, ZN => n34225);
   U8405 : NOR2_X1 port map( A1 => n34228, A2 => n34227, ZN => n34226);
   U8406 : NAND2_X1 port map( A1 => n15429, A2 => n29602, ZN => n34227);
   U8413 : MUX2_X1 port map( I0 => n12527, I1 => n36588, S => n5383, Z => n2334
                           );
   U8417 : NAND3_X2 port map( A1 => n36460, A2 => n34501, A3 => n36459, ZN => 
                           n3213);
   U8444 : OR2_X1 port map( A1 => n25829, A2 => n32193, Z => n1956);
   U8446 : OAI21_X2 port map( A1 => n20222, A2 => n35230, B => n20221, ZN => 
                           n23829);
   U8448 : XOR2_X1 port map( A1 => n21284, A2 => n34231, Z => n8554);
   U8456 : XOR2_X1 port map( A1 => n269, A2 => n35464, Z => n34231);
   U8463 : XOR2_X1 port map( A1 => n15871, A2 => n22621, Z => n22714);
   U8485 : NAND2_X2 port map( A1 => n6012, A2 => n35436, ZN => n34279);
   U8493 : NAND2_X2 port map( A1 => n34233, A2 => n12883, ZN => n16309);
   U8495 : OAI21_X2 port map( A1 => n12882, A2 => n32236, B => n21073, ZN => 
                           n34233);
   U8505 : INV_X2 port map( I => n34235, ZN => n33964);
   U8507 : XOR2_X1 port map( A1 => n12560, A2 => n12563, Z => n34235);
   U8515 : NAND3_X1 port map( A1 => n26217, A2 => n26216, A3 => n26218, ZN => 
                           n34237);
   U8516 : NAND2_X1 port map( A1 => n5670, A2 => n5525, ZN => n34515);
   U8522 : AOI21_X1 port map( A1 => n14928, A2 => n8493, B => n19604, ZN => 
                           n14927);
   U8525 : XOR2_X1 port map( A1 => n10117, A2 => n34238, Z => n32540);
   U8529 : XOR2_X1 port map( A1 => n38207, A2 => n34239, Z => n34238);
   U8556 : XOR2_X1 port map( A1 => n22552, A2 => n14309, Z => n7039);
   U8558 : NAND2_X2 port map( A1 => n13766, A2 => n13765, ZN => n14309);
   U8600 : BUF_X2 port map( I => n6263, Z => n34245);
   U8601 : NAND2_X1 port map( A1 => n30252, A2 => n30250, ZN => n16167);
   U8604 : NAND2_X2 port map( A1 => n19663, A2 => n30259, ZN => n30252);
   U8607 : NOR2_X1 port map( A1 => n21662, A2 => n36728, ZN => n21946);
   U8617 : NAND2_X2 port map( A1 => n35644, A2 => n32552, ZN => n23548);
   U8633 : NAND2_X2 port map( A1 => n18227, A2 => n21229, ZN => n34962);
   U8642 : OR2_X1 port map( A1 => n12078, A2 => n19371, Z => n9204);
   U8645 : OAI21_X2 port map( A1 => n26922, A2 => n19371, B => n26764, ZN => 
                           n12078);
   U8648 : XNOR2_X1 port map( A1 => n11201, A2 => n30065, ZN => n34274);
   U8664 : XOR2_X1 port map( A1 => Plaintext(157), A2 => Key(157), Z => n34247)
                           ;
   U8682 : XOR2_X1 port map( A1 => n12195, A2 => n18778, Z => n15413);
   U8684 : NAND2_X2 port map( A1 => n4630, A2 => n4629, ZN => n12195);
   U8695 : XOR2_X1 port map( A1 => n22747, A2 => n12194, Z => n34250);
   U8698 : NAND3_X2 port map( A1 => n7722, A2 => n18660, A3 => n22168, ZN => 
                           n23472);
   U8705 : INV_X4 port map( I => n25328, ZN => n36133);
   U8711 : XOR2_X1 port map( A1 => n8181, A2 => n34251, Z => n34594);
   U8729 : XOR2_X1 port map( A1 => n12935, A2 => n12934, Z => n12933);
   U8743 : XOR2_X1 port map( A1 => n30831, A2 => n17043, Z => n36034);
   U8813 : XOR2_X1 port map( A1 => n25249, A2 => n25100, Z => n24544);
   U8817 : NAND2_X2 port map( A1 => n33896, A2 => n8606, ZN => n25249);
   U8824 : XOR2_X1 port map( A1 => n23928, A2 => n23965, Z => n31851);
   U8855 : NAND2_X2 port map( A1 => n34984, A2 => n12499, ZN => n34559);
   U8877 : NOR2_X2 port map( A1 => n14091, A2 => n28426, ZN => n29167);
   U8879 : AOI21_X2 port map( A1 => n35525, A2 => n12083, B => n1292, ZN => 
                           n12027);
   U8880 : INV_X2 port map( I => n14011, ZN => n1292);
   U8884 : NAND2_X2 port map( A1 => n7011, A2 => n15375, ZN => n14011);
   U8900 : AOI21_X2 port map( A1 => n11379, A2 => n34246, B => n34259, ZN => 
                           n22623);
   U8915 : OAI22_X2 port map( A1 => n16580, A2 => n18290, B1 => n29482, B2 => 
                           n12479, ZN => n29531);
   U8925 : AOI22_X2 port map( A1 => n34868, A2 => n34262, B1 => n12590, B2 => 
                           n30335, ZN => n27064);
   U8933 : NOR2_X1 port map( A1 => n29841, A2 => n105, ZN => n21236);
   U8942 : NAND2_X2 port map( A1 => n33255, A2 => n13267, ZN => n20706);
   U8946 : XOR2_X1 port map( A1 => n7967, A2 => n24927, Z => n25156);
   U8949 : NAND2_X2 port map( A1 => n4224, A2 => n4227, ZN => n24927);
   U8957 : NAND3_X2 port map( A1 => n10003, A2 => n29851, A3 => n32258, ZN => 
                           n34267);
   U8970 : XOR2_X1 port map( A1 => n8702, A2 => n14507, Z => n20627);
   U8972 : NOR2_X2 port map( A1 => n7658, A2 => n9193, ZN => n34268);
   U8976 : INV_X2 port map( I => n17095, ZN => n13753);
   U8977 : NAND2_X2 port map( A1 => n33631, A2 => n3095, ZN => n17095);
   U8985 : XOR2_X1 port map( A1 => n32433, A2 => n25175, Z => n25254);
   U8987 : AOI21_X2 port map( A1 => n33755, A2 => n33754, B => n30385, ZN => 
                           n32433);
   U8988 : INV_X2 port map( I => n33539, ZN => n34857);
   U8996 : XOR2_X1 port map( A1 => n26342, A2 => n26494, Z => n10233);
   U9010 : NAND2_X2 port map( A1 => n34270, A2 => n13134, ZN => n5530);
   U9011 : OAI21_X2 port map( A1 => n13136, A2 => n37146, B => n13762, ZN => 
                           n34270);
   U9012 : NAND2_X2 port map( A1 => n34272, A2 => n39821, ZN => n36535);
   U9017 : NAND3_X1 port map( A1 => n17508, A2 => n32601, A3 => n17511, ZN => 
                           n22680);
   U9018 : XOR2_X1 port map( A1 => n20753, A2 => n34274, Z => n10501);
   U9035 : NAND2_X2 port map( A1 => n34275, A2 => n15795, ZN => n2542);
   U9040 : OAI21_X2 port map( A1 => n945, A2 => n15984, B => n34276, ZN => 
                           n15982);
   U9042 : NAND2_X2 port map( A1 => n15983, A2 => n945, ZN => n34276);
   U9057 : XOR2_X1 port map( A1 => n14941, A2 => n28991, Z => n29039);
   U9059 : NAND3_X2 port map( A1 => n28471, A2 => n28470, A3 => n28730, ZN => 
                           n28991);
   U9062 : XOR2_X1 port map( A1 => n11541, A2 => n22761, Z => n22543);
   U9065 : NAND2_X1 port map( A1 => n25544, A2 => n15515, ZN => n19702);
   U9067 : AOI21_X2 port map( A1 => n28107, A2 => n28108, B => n28106, ZN => 
                           n34695);
   U9076 : AOI21_X2 port map( A1 => n18312, A2 => n23333, B => n12191, ZN => 
                           n23245);
   U9078 : NAND2_X2 port map( A1 => n6969, A2 => n3256, ZN => n23333);
   U9081 : NOR2_X2 port map( A1 => n37171, A2 => n34277, ZN => n3112);
   U9088 : NAND2_X1 port map( A1 => n24577, A2 => n19484, ZN => n24578);
   U9099 : NAND2_X2 port map( A1 => n8262, A2 => n27240, ZN => n27102);
   U9105 : OR2_X1 port map( A1 => n21111, A2 => n18926, Z => n21558);
   U9124 : NAND2_X2 port map( A1 => n17299, A2 => n17301, ZN => n33230);
   U9135 : XOR2_X1 port map( A1 => n10492, A2 => n10491, Z => n9984);
   U9139 : XOR2_X1 port map( A1 => n34284, A2 => n17428, Z => Ciphertext(188));
   U9140 : AOI22_X1 port map( A1 => n16167, A2 => n11700, B1 => n13990, B2 => 
                           n13991, ZN => n34284);
   U9145 : INV_X2 port map( I => n28036, ZN => n28189);
   U9150 : XOR2_X1 port map( A1 => n34287, A2 => n20483, Z => Ciphertext(189));
   U9153 : XOR2_X1 port map( A1 => n36746, A2 => n34288, Z => n404);
   U9154 : XOR2_X1 port map( A1 => n3703, A2 => n4816, Z => n34288);
   U9162 : INV_X2 port map( I => n26075, ZN => n25992);
   U9167 : XOR2_X1 port map( A1 => n34289, A2 => n34703, Z => n9509);
   U9175 : XOR2_X1 port map( A1 => n33058, A2 => n19220, Z => n19418);
   U9177 : NOR2_X1 port map( A1 => n3815, A2 => n20078, ZN => n4379);
   U9187 : NAND2_X2 port map( A1 => n6116, A2 => n30993, ZN => n16559);
   U9188 : OAI22_X1 port map( A1 => n1218, A2 => n17095, B1 => n21050, B2 => 
                           n3977, ZN => n3979);
   U9190 : XOR2_X1 port map( A1 => n27735, A2 => n34290, Z => n27841);
   U9192 : NAND2_X1 port map( A1 => n27336, A2 => n27487, ZN => n34290);
   U9193 : NAND2_X2 port map( A1 => n36709, A2 => n34291, ZN => n29070);
   U9195 : XOR2_X1 port map( A1 => n2627, A2 => n27504, Z => n34986);
   U9204 : AND2_X1 port map( A1 => n29810, A2 => n29803, Z => n29812);
   U9253 : NAND2_X1 port map( A1 => n8529, A2 => n30049, ZN => n19108);
   U9254 : AND2_X1 port map( A1 => n11453, A2 => n34506, Z => n4960);
   U9255 : OAI21_X1 port map( A1 => n1340, A2 => n32478, B => n34296, ZN => 
                           n22308);
   U9260 : NAND2_X1 port map( A1 => n32478, A2 => n22307, ZN => n34296);
   U9273 : NOR2_X2 port map( A1 => n35660, A2 => n35117, ZN => n34297);
   U9283 : NOR2_X2 port map( A1 => n1432, A2 => n28690, ZN => n34298);
   U9293 : NAND2_X1 port map( A1 => n27137, A2 => n8798, ZN => n34299);
   U9309 : AOI21_X2 port map( A1 => n13403, A2 => n11488, B => n13401, ZN => 
                           n34301);
   U9319 : NAND2_X1 port map( A1 => n1340, A2 => n4200, ZN => n21337);
   U9321 : NOR2_X2 port map( A1 => n20740, A2 => n12306, ZN => n15986);
   U9324 : NOR2_X2 port map( A1 => n18879, A2 => n18956, ZN => n20740);
   U9351 : OAI21_X2 port map( A1 => n34303, A2 => n1564, B => n24630, ZN => 
                           n14768);
   U9394 : XOR2_X1 port map( A1 => n34306, A2 => n3802, Z => n26265);
   U9395 : XOR2_X1 port map( A1 => n26528, A2 => n36644, Z => n34306);
   U9396 : OAI22_X2 port map( A1 => n19364, A2 => n26992, B1 => n13110, B2 => 
                           n14459, ZN => n26877);
   U9417 : NOR2_X1 port map( A1 => n14502, A2 => n11778, ZN => n6018);
   U9435 : NAND3_X1 port map( A1 => n4171, A2 => n12328, A3 => n32168, ZN => 
                           n34461);
   U9446 : NAND3_X1 port map( A1 => n9913, A2 => n969, A3 => n29477, ZN => 
                           n9104);
   U9447 : NAND2_X2 port map( A1 => n34559, A2 => n35203, ZN => n13170);
   U9469 : NOR2_X2 port map( A1 => n30356, A2 => n30336, ZN => n34311);
   U9473 : NAND2_X2 port map( A1 => n36526, A2 => n27356, ZN => n27766);
   U9474 : NAND2_X2 port map( A1 => n34953, A2 => n36436, ZN => n12437);
   U9477 : BUF_X2 port map( I => n19113, Z => n34312);
   U9483 : INV_X4 port map( I => n16853, ZN => n1424);
   U9491 : NOR2_X2 port map( A1 => n32450, A2 => n5112, ZN => n2149);
   U9502 : OR2_X1 port map( A1 => n38395, A2 => n17864, Z => n22148);
   U9507 : XOR2_X1 port map( A1 => n26221, A2 => n16497, Z => n15821);
   U9508 : OR2_X1 port map( A1 => n858, A2 => n33895, Z => n26872);
   U9515 : XOR2_X1 port map( A1 => n34314, A2 => n34313, Z => n36602);
   U9518 : XOR2_X1 port map( A1 => n31585, A2 => n29857, Z => n34314);
   U9527 : OAI21_X2 port map( A1 => n15992, A2 => n37184, B => n15991, ZN => 
                           n34898);
   U9531 : NOR2_X2 port map( A1 => n25433, A2 => n25685, ZN => n15992);
   U9537 : XOR2_X1 port map( A1 => n17478, A2 => n34315, Z => n24039);
   U9544 : OAI21_X2 port map( A1 => n16227, A2 => n16228, B => n20943, ZN => 
                           n34317);
   U9549 : OAI21_X2 port map( A1 => n16306, A2 => n8933, B => n8932, ZN => 
                           n17417);
   U9556 : OAI21_X1 port map( A1 => n30118, A2 => n30119, B => n34319, ZN => 
                           n19031);
   U9557 : AOI22_X1 port map( A1 => n19032, A2 => n10118, B1 => n19033, B2 => 
                           n16180, ZN => n34319);
   U9560 : XOR2_X1 port map( A1 => n29063, A2 => n29115, Z => n14388);
   U9565 : OAI21_X2 port map( A1 => n36031, A2 => n36032, B => n28587, ZN => 
                           n29063);
   U9567 : NAND2_X2 port map( A1 => n24639, A2 => n24732, ZN => n24843);
   U9579 : NAND2_X2 port map( A1 => n20378, A2 => n36267, ZN => n24639);
   U9585 : OAI21_X1 port map( A1 => n16060, A2 => n30047, B => n8529, ZN => 
                           n16059);
   U9593 : XOR2_X1 port map( A1 => n27469, A2 => n10866, Z => n35834);
   U9613 : NOR2_X2 port map( A1 => n31205, A2 => n26131, ZN => n26132);
   U9629 : INV_X2 port map( I => n17618, ZN => n14167);
   U9630 : NAND2_X2 port map( A1 => n36229, A2 => n23822, ZN => n17618);
   U9632 : XOR2_X1 port map( A1 => n34323, A2 => n19432, Z => Ciphertext(84));
   U9644 : NAND2_X2 port map( A1 => n34324, A2 => n25678, ZN => n33909);
   U9648 : OAI22_X2 port map( A1 => n25676, A2 => n14273, B1 => n25675, B2 => 
                           n19589, ZN => n34324);
   U9650 : OAI21_X2 port map( A1 => n15110, A2 => n28756, B => n15109, ZN => 
                           n15270);
   U9656 : XOR2_X1 port map( A1 => n13189, A2 => n13187, Z => n34325);
   U9661 : NAND2_X1 port map( A1 => n8014, A2 => n5227, ZN => n24943);
   U9680 : AOI22_X1 port map( A1 => n6629, A2 => n8082, B1 => n35172, B2 => 
                           n19893, ZN => n34326);
   U9693 : OAI21_X2 port map( A1 => n35514, A2 => n38337, B => n35513, ZN => 
                           n19976);
   U9701 : INV_X2 port map( I => n27499, ZN => n34332);
   U9729 : AOI21_X2 port map( A1 => n5751, A2 => n19470, B => n34329, ZN => 
                           n3271);
   U9730 : INV_X2 port map( I => n7900, ZN => n34329);
   U9733 : NAND2_X2 port map( A1 => n21517, A2 => n261, ZN => n7900);
   U9770 : AND2_X1 port map( A1 => n14793, A2 => n36922, Z => n36575);
   U9785 : NAND2_X2 port map( A1 => n34335, A2 => n32036, ZN => n4771);
   U9790 : AND2_X1 port map( A1 => n20359, A2 => n32951, Z => n36707);
   U9792 : XOR2_X1 port map( A1 => n5694, A2 => n30907, Z => n15047);
   U9793 : INV_X2 port map( I => n23561, ZN => n34336);
   U9800 : NOR2_X1 port map( A1 => n31078, A2 => n36380, ZN => n19140);
   U9814 : AOI21_X2 port map( A1 => n28195, A2 => n9897, B => n34342, ZN => 
                           n15473);
   U9822 : NAND2_X2 port map( A1 => n34343, A2 => n20665, ZN => n25175);
   U9824 : NAND3_X2 port map( A1 => n30419, A2 => n17377, A3 => n20158, ZN => 
                           n34343);
   U9830 : AOI22_X2 port map( A1 => n21915, A2 => n5391, B1 => n21913, B2 => 
                           n938, ZN => n5303);
   U9842 : XNOR2_X1 port map( A1 => n16526, A2 => n14164, ZN => n25285);
   U9849 : NAND2_X2 port map( A1 => n1898, A2 => n30572, ZN => n19979);
   U9850 : NOR2_X2 port map( A1 => n32633, A2 => n19465, ZN => n35452);
   U9852 : NAND2_X2 port map( A1 => n7305, A2 => n2140, ZN => n32633);
   U9854 : INV_X2 port map( I => n34347, ZN => n15592);
   U9862 : XOR2_X1 port map( A1 => n26207, A2 => n20213, Z => n26529);
   U9864 : AOI21_X2 port map( A1 => n10139, A2 => n10138, B => n10137, ZN => 
                           n26207);
   U9867 : XOR2_X1 port map( A1 => n7060, A2 => n12988, Z => n7059);
   U9871 : OR2_X1 port map( A1 => n1190, A2 => n11296, Z => n28634);
   U9888 : XOR2_X1 port map( A1 => n34352, A2 => n5279, Z => n33856);
   U9894 : XOR2_X1 port map( A1 => n22586, A2 => n33824, Z => n34352);
   U9909 : NAND2_X2 port map( A1 => n15618, A2 => n26099, ZN => n26421);
   U9910 : NAND2_X2 port map( A1 => n16118, A2 => n16117, ZN => n26234);
   U9911 : OR2_X1 port map( A1 => n38194, A2 => n34354, Z => n18196);
   U9932 : NAND3_X2 port map( A1 => n13571, A2 => n4662, A3 => n4661, ZN => 
                           n9873);
   U9939 : XOR2_X1 port map( A1 => n4783, A2 => n14174, Z => n27575);
   U9947 : XOR2_X1 port map( A1 => n22599, A2 => n12730, Z => n6311);
   U9952 : NAND2_X2 port map( A1 => n13480, A2 => n15487, ZN => n12730);
   U9959 : NAND2_X1 port map( A1 => n30304, A2 => n13601, ZN => n28431);
   U9961 : XOR2_X1 port map( A1 => n7068, A2 => n27820, Z => n35871);
   U9965 : OR2_X1 port map( A1 => n5112, A2 => n8069, Z => n13033);
   U9973 : XOR2_X1 port map( A1 => n34358, A2 => n30839, Z => n31121);
   U10015 : XOR2_X1 port map( A1 => n9085, A2 => n38176, Z => n26397);
   U10026 : NAND2_X2 port map( A1 => n31098, A2 => n3846, ZN => n3845);
   U10028 : XOR2_X1 port map( A1 => n1884, A2 => n1885, Z => n1883);
   U10054 : NAND2_X2 port map( A1 => n28264, A2 => n28263, ZN => n28745);
   U10055 : XOR2_X1 port map( A1 => n35209, A2 => n7402, Z => n26537);
   U10080 : INV_X2 port map( I => n34365, ZN => n871);
   U10089 : OR2_X1 port map( A1 => n30859, A2 => n4599, Z => n26882);
   U10092 : NOR2_X2 port map( A1 => n34366, A2 => n17789, ZN => n21242);
   U10093 : XOR2_X1 port map( A1 => n3292, A2 => n25065, Z => n9781);
   U10120 : INV_X2 port map( I => n34370, ZN => n33960);
   U10121 : XOR2_X1 port map( A1 => n20693, A2 => n10169, Z => n34370);
   U10123 : NAND2_X2 port map( A1 => n34371, A2 => n13334, ZN => n17132);
   U10124 : NOR2_X2 port map( A1 => n34372, A2 => n34123, ZN => n2288);
   U10126 : NAND3_X1 port map( A1 => n31280, A2 => n31279, A3 => n12876, ZN => 
                           n31704);
   U10130 : NAND2_X2 port map( A1 => n34904, A2 => n34905, ZN => n11950);
   U10140 : NAND2_X2 port map( A1 => n966, A2 => n13192, ZN => n13986);
   U10147 : XOR2_X1 port map( A1 => n467, A2 => n29025, Z => n34375);
   U10166 : XOR2_X1 port map( A1 => n34377, A2 => n23744, Z => n36952);
   U10172 : XOR2_X1 port map( A1 => n23846, A2 => n23987, Z => n34377);
   U10177 : NAND2_X2 port map( A1 => n10553, A2 => n10551, ZN => n36442);
   U10186 : INV_X2 port map( I => n17864, ZN => n34379);
   U10187 : OR2_X1 port map( A1 => n22238, A2 => n34379, Z => n9524);
   U10215 : NAND2_X2 port map( A1 => n34383, A2 => n9993, ZN => n36857);
   U10217 : OAI21_X2 port map( A1 => n18720, A2 => n29491, B => n29418, ZN => 
                           n34383);
   U10221 : NOR2_X1 port map( A1 => n19985, A2 => n32164, ZN => n34931);
   U10223 : NAND3_X2 port map( A1 => n1956, A2 => n1743, A3 => n1954, ZN => 
                           n7402);
   U10235 : NAND2_X2 port map( A1 => n30929, A2 => n30930, ZN => n33271);
   U10240 : XOR2_X1 port map( A1 => n23776, A2 => n16138, Z => n4562);
   U10242 : AND2_X1 port map( A1 => n15626, A2 => n12144, Z => n13345);
   U10248 : NAND2_X2 port map( A1 => n2191, A2 => n38629, ZN => n28580);
   U10259 : XOR2_X1 port map( A1 => n33921, A2 => n34017, Z => n824);
   U10260 : INV_X2 port map( I => n31872, ZN => n25214);
   U10262 : XOR2_X1 port map( A1 => n31872, A2 => n34391, Z => n17834);
   U10263 : INV_X1 port map( I => n29974, ZN => n34391);
   U10265 : NAND2_X2 port map( A1 => n35785, A2 => n35784, ZN => n31872);
   U10267 : NOR2_X2 port map( A1 => n193, A2 => n20451, ZN => n34469);
   U10269 : NAND2_X2 port map( A1 => n34392, A2 => n13589, ZN => n26134);
   U10277 : XOR2_X1 port map( A1 => n34394, A2 => n30207, Z => Ciphertext(181))
                           ;
   U10282 : NAND3_X2 port map( A1 => n30205, A2 => n16548, A3 => n30206, ZN => 
                           n34394);
   U10310 : XOR2_X1 port map( A1 => n34397, A2 => n354, Z => n32951);
   U10315 : XOR2_X1 port map( A1 => n34398, A2 => n391, Z => n36292);
   U10317 : XOR2_X1 port map( A1 => n4673, A2 => n34088, Z => n34398);
   U10333 : INV_X4 port map( I => n11628, ZN => n1198);
   U10383 : NAND2_X2 port map( A1 => n17865, A2 => n6269, ZN => n17864);
   U10413 : NAND2_X2 port map( A1 => n34405, A2 => n34404, ZN => n30424);
   U10420 : INV_X2 port map( I => n22145, ZN => n34404);
   U10496 : NOR2_X2 port map( A1 => n7916, A2 => n22238, ZN => n34406);
   U10501 : XOR2_X1 port map( A1 => n34408, A2 => n16103, Z => n16102);
   U10504 : NAND3_X2 port map( A1 => n36403, A2 => n32668, A3 => n36402, ZN => 
                           n29930);
   U10505 : XOR2_X1 port map( A1 => n10343, A2 => n14307, Z => n5728);
   U10537 : NAND2_X2 port map( A1 => n24364, A2 => n24365, ZN => n25181);
   U10547 : XOR2_X1 port map( A1 => n19072, A2 => n20618, Z => n32210);
   U10558 : NAND2_X1 port map( A1 => n15751, A2 => n24477, ZN => n24479);
   U10560 : NOR2_X2 port map( A1 => n31159, A2 => n31158, ZN => n35828);
   U10568 : XOR2_X1 port map( A1 => n8894, A2 => n31620, Z => n18498);
   U10570 : OR2_X1 port map( A1 => n20056, A2 => n35149, Z => n28197);
   U10573 : AND2_X1 port map( A1 => n5457, A2 => n14858, Z => n5456);
   U10578 : AOI21_X2 port map( A1 => n9135, A2 => n2192, B => n33580, ZN => 
                           n35924);
   U10587 : AOI22_X2 port map( A1 => n34857, A2 => n26055, B1 => n26054, B2 => 
                           n25424, ZN => n6784);
   U10595 : NAND2_X2 port map( A1 => n34415, A2 => n27994, ZN => n28659);
   U10596 : AND2_X1 port map( A1 => n27993, A2 => n27992, Z => n34415);
   U10614 : XOR2_X1 port map( A1 => n15050, A2 => n34418, Z => n15052);
   U10617 : XOR2_X1 port map( A1 => n24987, A2 => n34147, Z => n34418);
   U10625 : NAND2_X2 port map( A1 => n34420, A2 => n16374, ZN => n35952);
   U10663 : OAI22_X2 port map( A1 => n18559, A2 => n21589, B1 => n18560, B2 => 
                           n18561, ZN => n22341);
   U10666 : XOR2_X1 port map( A1 => n14144, A2 => n34428, Z => n26861);
   U10671 : XOR2_X1 port map( A1 => n19051, A2 => n14143, Z => n34428);
   U10676 : XOR2_X1 port map( A1 => n2218, A2 => n2217, Z => n20686);
   U10688 : NAND2_X1 port map( A1 => n4986, A2 => n16449, ZN => n34430);
   U10696 : XOR2_X1 port map( A1 => n36041, A2 => n8100, Z => n9374);
   U10717 : XOR2_X1 port map( A1 => n24049, A2 => n23757, Z => n34435);
   U10732 : XOR2_X1 port map( A1 => n19989, A2 => n19987, Z => n28174);
   U10739 : OR2_X1 port map( A1 => n24470, A2 => n15461, Z => n36789);
   U10745 : XOR2_X1 port map( A1 => n22082, A2 => n696, Z => n18434);
   U10750 : NAND2_X2 port map( A1 => n34438, A2 => n34437, ZN => n33919);
   U10753 : NAND2_X1 port map( A1 => n32760, A2 => n18926, ZN => n21559);
   U10756 : XOR2_X1 port map( A1 => n34439, A2 => n4070, Z => n31294);
   U10768 : INV_X2 port map( I => n22588, ZN => n34440);
   U10777 : NAND3_X2 port map( A1 => n28547, A2 => n14278, A3 => n28735, ZN => 
                           n28627);
   U10781 : NOR2_X2 port map( A1 => n1752, A2 => n34446, ZN => n34503);
   U10790 : AOI21_X1 port map( A1 => n36678, A2 => n1551, B => n371, ZN => 
                           n3278);
   U10798 : BUF_X2 port map( I => n19417, Z => n34447);
   U10804 : NAND2_X2 port map( A1 => n32132, A2 => n32413, ZN => n32575);
   U10812 : NOR2_X2 port map( A1 => n19373, A2 => n9165, ZN => n11364);
   U10819 : NAND2_X2 port map( A1 => n32583, A2 => n34448, ZN => n23532);
   U10825 : XOR2_X1 port map( A1 => n10771, A2 => n34450, Z => n10770);
   U10827 : XOR2_X1 port map( A1 => n23968, A2 => n34451, Z => n34450);
   U10838 : XOR2_X1 port map( A1 => n34453, A2 => n12912, Z => n12951);
   U10855 : XOR2_X1 port map( A1 => n4326, A2 => n22957, Z => n34453);
   U10857 : XOR2_X1 port map( A1 => n5724, A2 => n34454, Z => n11896);
   U10858 : XOR2_X1 port map( A1 => n29821, A2 => n5728, Z => n34454);
   U10871 : OR2_X1 port map( A1 => n17917, A2 => n22921, Z => n32133);
   U10920 : NAND2_X2 port map( A1 => n35453, A2 => n20644, ZN => n8407);
   U10930 : NAND3_X2 port map( A1 => n32752, A2 => n32650, A3 => n31882, ZN => 
                           n15855);
   U10937 : AOI21_X2 port map( A1 => n36850, A2 => n12273, B => n12272, ZN => 
                           n34460);
   U10940 : NAND2_X2 port map( A1 => n34995, A2 => n20172, ZN => n7044);
   U10950 : AOI22_X2 port map( A1 => n11713, A2 => n11712, B1 => n11711, B2 => 
                           n10013, ZN => n19156);
   U10958 : XOR2_X1 port map( A1 => n25127, A2 => n25177, Z => n25217);
   U10964 : OAI21_X1 port map( A1 => n22975, A2 => n34467, B => n34466, ZN => 
                           n23087);
   U10966 : NAND2_X1 port map( A1 => n34467, A2 => n23167, ZN => n34466);
   U10967 : XOR2_X1 port map( A1 => n34468, A2 => n34104, Z => n35687);
   U10985 : AOI21_X2 port map( A1 => n37279, A2 => n23559, B => n34336, ZN => 
                           n34472);
   U10990 : INV_X2 port map( I => n34473, ZN => n33579);
   U11005 : INV_X2 port map( I => n17597, ZN => n12940);
   U11013 : NAND3_X1 port map( A1 => n15080, A2 => n15081, A3 => n19538, ZN => 
                           n15079);
   U11017 : XOR2_X1 port map( A1 => n17430, A2 => n34474, Z => n17830);
   U11018 : XOR2_X1 port map( A1 => n12125, A2 => n17429, Z => n34474);
   U11020 : NAND2_X1 port map( A1 => n19631, A2 => n1195, ZN => n12336);
   U11021 : NAND2_X2 port map( A1 => n11280, A2 => n11279, ZN => n1195);
   U11022 : INV_X4 port map( I => n33579, ZN => n35314);
   U11023 : INV_X4 port map( I => n34475, ZN => n22324);
   U11040 : NAND2_X1 port map( A1 => n20948, A2 => n20949, ZN => n34476);
   U11045 : OAI22_X1 port map( A1 => n21302, A2 => n17246, B1 => n955, B2 => 
                           n826, ZN => n15543);
   U11046 : AND2_X1 port map( A1 => n4377, A2 => n4378, Z => n4168);
   U11047 : XOR2_X1 port map( A1 => n34477, A2 => n32604, Z => n28848);
   U11058 : XOR2_X1 port map( A1 => n17797, A2 => n34478, Z => n31261);
   U11066 : NAND2_X2 port map( A1 => n34480, A2 => n4504, ZN => n16619);
   U11070 : NAND2_X2 port map( A1 => n6747, A2 => n20441, ZN => n25435);
   U11073 : XNOR2_X1 port map( A1 => n5816, A2 => n5815, ZN => n34483);
   U11076 : XOR2_X1 port map( A1 => n23926, A2 => n23925, Z => n1929);
   U11088 : NAND3_X1 port map( A1 => n32497, A2 => n6578, A3 => n9530, ZN => 
                           n34486);
   U11094 : XOR2_X1 port map( A1 => n21284, A2 => n27720, Z => n18049);
   U11096 : XOR2_X1 port map( A1 => n27773, A2 => n27503, Z => n21284);
   U11101 : XOR2_X1 port map( A1 => n26364, A2 => n26336, Z => n9555);
   U11104 : XOR2_X1 port map( A1 => n1009, A2 => n7133, Z => n26364);
   U11135 : NAND2_X2 port map( A1 => n28299, A2 => n16303, ZN => n28301);
   U11137 : NOR2_X2 port map( A1 => n13323, A2 => n13321, ZN => n16303);
   U11139 : NOR2_X1 port map( A1 => n34561, A2 => n24287, ZN => n14684);
   U11146 : XOR2_X1 port map( A1 => n5610, A2 => n26514, Z => n34489);
   U11149 : OAI22_X1 port map( A1 => n19564, A2 => n1478, B1 => n18246, B2 => 
                           n1085, ZN => n7232);
   U11150 : NAND2_X1 port map( A1 => n35881, A2 => n19587, ZN => n5533);
   U11154 : NOR2_X2 port map( A1 => n4317, A2 => n22157, ZN => n6582);
   U11168 : XOR2_X1 port map( A1 => n3376, A2 => n3375, Z => n24192);
   U11171 : INV_X2 port map( I => n34490, ZN => n30454);
   U11173 : XOR2_X1 port map( A1 => n15860, A2 => n15859, Z => n34490);
   U11175 : NAND2_X2 port map( A1 => n36947, A2 => n28964, ZN => n13192);
   U11176 : XOR2_X1 port map( A1 => n15220, A2 => n25198, Z => n3185);
   U11177 : AOI22_X2 port map( A1 => n2930, A2 => n20168, B1 => n31568, B2 => 
                           n25242, ZN => n15220);
   U11191 : XOR2_X1 port map( A1 => n5347, A2 => n33478, Z => n5348);
   U11193 : BUF_X2 port map( I => n33609, Z => n34494);
   U11194 : XOR2_X1 port map( A1 => n26335, A2 => n34495, Z => n19533);
   U11198 : XOR2_X1 port map( A1 => n26585, A2 => n34768, Z => n26335);
   U11203 : NOR2_X2 port map( A1 => n32853, A2 => n32852, ZN => n27574);
   U11207 : NOR3_X1 port map( A1 => n35588, A2 => n34622, A3 => n30004, ZN => 
                           n30008);
   U11217 : INV_X2 port map( I => n34496, ZN => n19891);
   U11219 : XNOR2_X1 port map( A1 => n9039, A2 => n8781, ZN => n34496);
   U11221 : XOR2_X1 port map( A1 => n3773, A2 => n34497, Z => n10620);
   U11222 : XOR2_X1 port map( A1 => n33672, A2 => n34498, Z => n34497);
   U11228 : NAND2_X2 port map( A1 => n29237, A2 => n3263, ZN => n29228);
   U11231 : NAND2_X2 port map( A1 => n16839, A2 => n29079, ZN => n29237);
   U11238 : XOR2_X1 port map( A1 => n8474, A2 => n2371, Z => n2370);
   U11241 : NAND2_X1 port map( A1 => n6248, A2 => n25328, ZN => n34501);
   U11256 : NAND2_X2 port map( A1 => n34503, A2 => n14790, ZN => n13151);
   U11264 : NAND2_X2 port map( A1 => n13970, A2 => n1123, ZN => n34504);
   U11265 : NOR2_X2 port map( A1 => n36683, A2 => n26, ZN => n16578);
   U11267 : NOR2_X2 port map( A1 => n16407, A2 => n25961, ZN => n25923);
   U11282 : INV_X2 port map( I => n9920, ZN => n34506);
   U11294 : AOI22_X2 port map( A1 => n38011, A2 => n5451, B1 => n17249, B2 => 
                           n938, ZN => n5776);
   U11298 : NAND2_X2 port map( A1 => n2566, A2 => n28693, ZN => n31127);
   U11305 : XOR2_X1 port map( A1 => n19766, A2 => n16362, Z => n3890);
   U11322 : NAND2_X2 port map( A1 => n35899, A2 => n17997, ZN => n11968);
   U11323 : XOR2_X1 port map( A1 => n476, A2 => n39575, Z => n20016);
   U11328 : NAND2_X2 port map( A1 => n35012, A2 => n23485, ZN => n476);
   U11332 : XOR2_X1 port map( A1 => n35227, A2 => n27845, Z => n27605);
   U11333 : NAND2_X2 port map( A1 => n22493, A2 => n6176, ZN => n23480);
   U11338 : NOR2_X2 port map( A1 => n28207, A2 => n7541, ZN => n28720);
   U11343 : AOI22_X2 port map( A1 => n16308, A2 => n19754, B1 => n5396, B2 => 
                           n34510, ZN => n20319);
   U11344 : OAI21_X1 port map( A1 => n1222, A2 => n15284, B => n27197, ZN => 
                           n6508);
   U11349 : XOR2_X1 port map( A1 => n25310, A2 => n6232, Z => n6231);
   U11350 : XOR2_X1 port map( A1 => n34091, A2 => n3776, Z => n35129);
   U11357 : AOI21_X2 port map( A1 => n34512, A2 => n32333, B => n37008, ZN => 
                           n37007);
   U11370 : AOI21_X2 port map( A1 => n16201, A2 => n36722, B => n11668, ZN => 
                           n26556);
   U11372 : XOR2_X1 port map( A1 => n34514, A2 => n17707, Z => n10039);
   U11379 : XOR2_X1 port map( A1 => n30318, A2 => n24873, Z => n34514);
   U11390 : XOR2_X1 port map( A1 => n8284, A2 => n30994, Z => n11782);
   U11401 : XOR2_X1 port map( A1 => n34518, A2 => n30423, Z => n32838);
   U11404 : NOR2_X1 port map( A1 => n25957, A2 => n18406, ZN => n34519);
   U11407 : OAI22_X2 port map( A1 => n29782, A2 => n16682, B1 => n19716, B2 => 
                           n3096, ZN => n29798);
   U11421 : XOR2_X1 port map( A1 => n20065, A2 => n215, Z => n35269);
   U11426 : XOR2_X1 port map( A1 => n20540, A2 => n7474, Z => n215);
   U11436 : INV_X2 port map( I => n34521, ZN => n37050);
   U11437 : XNOR2_X1 port map( A1 => n35510, A2 => n13938, ZN => n34521);
   U11440 : NAND2_X2 port map( A1 => n25593, A2 => n19401, ZN => n25961);
   U11461 : NAND2_X2 port map( A1 => n22919, A2 => n23072, ZN => n34557);
   U11464 : NAND3_X2 port map( A1 => n15836, A2 => n6450, A3 => n16259, ZN => 
                           n9719);
   U11466 : INV_X1 port map( I => n34522, ZN => n23143);
   U11468 : NOR2_X1 port map( A1 => n8765, A2 => n34522, ZN => n5628);
   U11470 : AOI21_X2 port map( A1 => n32248, A2 => n12263, B => n12427, ZN => 
                           n8894);
   U11472 : NOR2_X2 port map( A1 => n826, A2 => n37050, ZN => n25602);
   U11479 : OAI21_X2 port map( A1 => n33892, A2 => n33891, B => n25911, ZN => 
                           n34768);
   U11480 : AOI21_X1 port map( A1 => n10479, A2 => n17515, B => n9690, ZN => 
                           n17514);
   U11509 : NOR2_X2 port map( A1 => n32358, A2 => n31465, ZN => n2600);
   U11523 : INV_X2 port map( I => n34532, ZN => n26724);
   U11527 : XOR2_X1 port map( A1 => n19021, A2 => n19018, Z => n34532);
   U11528 : AOI22_X2 port map( A1 => n34533, A2 => n1523, B1 => n5475, B2 => 
                           n5886, ZN => n5474);
   U11546 : OAI22_X1 port map( A1 => n29511, A2 => n35180, B1 => n29524, B2 => 
                           n29531, ZN => n29512);
   U11564 : XOR2_X1 port map( A1 => n35227, A2 => n14808, Z => n27806);
   U11565 : AOI21_X2 port map( A1 => n27073, A2 => n18228, B => n30933, ZN => 
                           n35227);
   U11574 : NAND2_X2 port map( A1 => n6554, A2 => n34540, ZN => n10461);
   U11576 : AOI22_X2 port map( A1 => n6312, A2 => n441, B1 => n6313, B2 => 
                           n18809, ZN => n34540);
   U11607 : INV_X2 port map( I => n34546, ZN => n16692);
   U11608 : XNOR2_X1 port map( A1 => n22605, A2 => n33856, ZN => n34546);
   U11610 : INV_X4 port map( I => n9193, ZN => n1034);
   U11618 : NAND2_X1 port map( A1 => n692, A2 => n9833, ZN => n16240);
   U11623 : BUF_X2 port map( I => n35233, Z => n34547);
   U11638 : XOR2_X1 port map( A1 => n18490, A2 => n26519, Z => n12429);
   U11648 : INV_X2 port map( I => n34549, ZN => n36197);
   U11655 : XOR2_X1 port map( A1 => n33112, A2 => n33111, Z => n34549);
   U11667 : AOI21_X1 port map( A1 => n11111, A2 => n19108, B => n29935, ZN => 
                           n10097);
   U11668 : XOR2_X1 port map( A1 => n34552, A2 => n29849, Z => Ciphertext(114))
                           ;
   U11673 : NAND2_X2 port map( A1 => n36555, A2 => n34554, ZN => n7481);
   U11676 : XOR2_X1 port map( A1 => n27847, A2 => n35678, Z => n16607);
   U11690 : INV_X4 port map( I => n33952, ZN => n36262);
   U11691 : OAI21_X2 port map( A1 => n34072, A2 => n22919, B => n34557, ZN => 
                           n22828);
   U11701 : AOI21_X2 port map( A1 => n6654, A2 => n13685, B => n13684, ZN => 
                           n13683);
   U11703 : XOR2_X1 port map( A1 => n23830, A2 => n23804, Z => n6530);
   U11709 : XOR2_X1 port map( A1 => n26396, A2 => n3781, Z => n26205);
   U11717 : NOR2_X1 port map( A1 => n32682, A2 => n36935, ZN => n34568);
   U11718 : AND2_X1 port map( A1 => n36323, A2 => n25601, Z => n35632);
   U11728 : NOR2_X1 port map( A1 => n32059, A2 => n10254, ZN => n34569);
   U11738 : XOR2_X1 port map( A1 => n4223, A2 => n4221, Z => n30233);
   U11745 : NAND2_X2 port map( A1 => n31028, A2 => n34571, ZN => n9413);
   U11752 : INV_X2 port map( I => n12234, ZN => n34574);
   U11755 : XOR2_X1 port map( A1 => n17593, A2 => n25087, Z => n12311);
   U11757 : INV_X2 port map( I => n34957, ZN => n26905);
   U11767 : AOI21_X2 port map( A1 => n34575, A2 => n19402, B => n9371, ZN => 
                           n33108);
   U11770 : NAND2_X2 port map( A1 => n6515, A2 => n33599, ZN => n34575);
   U11786 : INV_X2 port map( I => n37085, ZN => n13166);
   U11787 : NAND2_X1 port map( A1 => n37085, A2 => n34576, ZN => n19463);
   U11790 : XOR2_X1 port map( A1 => n35645, A2 => n12293, Z => n18507);
   U11794 : XNOR2_X1 port map( A1 => n26566, A2 => n20139, ZN => n34593);
   U11797 : AND2_X1 port map( A1 => n26905, A2 => n39477, Z => n9423);
   U11806 : NAND2_X1 port map( A1 => n6415, A2 => n9267, ZN => n6414);
   U11808 : NAND2_X2 port map( A1 => n3918, A2 => n12887, ZN => n9267);
   U11820 : XOR2_X1 port map( A1 => n34580, A2 => n18852, Z => n13127);
   U11823 : OAI21_X2 port map( A1 => n14695, A2 => n3783, B => n38305, ZN => 
                           n21139);
   U11828 : XOR2_X1 port map( A1 => n2431, A2 => n38167, Z => n32512);
   U11831 : NOR3_X2 port map( A1 => n1541, A2 => n6300, A3 => n34010, ZN => 
                           n34581);
   U11837 : XOR2_X1 port map( A1 => n32298, A2 => n35243, Z => n4815);
   U11870 : NOR2_X2 port map( A1 => n34801, A2 => n12651, ZN => n12650);
   U11885 : XOR2_X1 port map( A1 => n27864, A2 => n10653, Z => n9160);
   U11888 : XOR2_X1 port map( A1 => n34586, A2 => n23755, Z => n12520);
   U11922 : INV_X2 port map( I => n34587, ZN => n15922);
   U11950 : NAND2_X2 port map( A1 => n13911, A2 => n13909, ZN => n22511);
   U11957 : XOR2_X1 port map( A1 => n3705, A2 => n3707, Z => n4386);
   U11958 : XOR2_X1 port map( A1 => n23734, A2 => n23662, Z => n11724);
   U11961 : AOI22_X2 port map( A1 => n34589, A2 => n30225, B1 => n30222, B2 => 
                           n30223, ZN => n30259);
   U11978 : XOR2_X1 port map( A1 => n23419, A2 => n9344, Z => n23830);
   U11989 : OR2_X1 port map( A1 => n10375, A2 => n10334, Z => n10377);
   U11994 : NAND2_X1 port map( A1 => n30647, A2 => n30646, ZN => n34750);
   U11996 : XOR2_X1 port map( A1 => n32844, A2 => n34593, Z => n30989);
   U11998 : OR2_X1 port map( A1 => n25923, A2 => n25922, Z => n15378);
   U11999 : XOR2_X1 port map( A1 => n16085, A2 => n27161, Z => n4364);
   U12004 : AND2_X1 port map( A1 => n24538, A2 => n35893, Z => n35119);
   U12035 : NOR2_X2 port map( A1 => n17476, A2 => n34596, ZN => n28578);
   U12044 : INV_X2 port map( I => n34597, ZN => n31010);
   U12050 : XNOR2_X1 port map( A1 => n33044, A2 => n11103, ZN => n34597);
   U12057 : NOR2_X1 port map( A1 => n31010, A2 => n9740, ZN => n8494);
   U12058 : INV_X2 port map( I => n36226, ZN => n1097);
   U12068 : NAND2_X1 port map( A1 => n8158, A2 => n8159, ZN => n8157);
   U12072 : NAND2_X1 port map( A1 => n35745, A2 => n34279, ZN => n20143);
   U12081 : XOR2_X1 port map( A1 => n33400, A2 => n39320, Z => n33399);
   U12103 : OAI21_X2 port map( A1 => n4466, A2 => n4465, B => n4464, ZN => 
                           n26090);
   U12112 : NOR2_X2 port map( A1 => n34599, A2 => n35935, ZN => n29166);
   U12126 : NAND2_X1 port map( A1 => n13082, A2 => n32638, ZN => n27974);
   U12132 : BUF_X2 port map( I => Key(67), Z => n29879);
   U12144 : AOI22_X1 port map( A1 => n29890, A2 => n32706, B1 => n17286, B2 => 
                           n11182, ZN => n11785);
   U12149 : AOI22_X2 port map( A1 => n6703, A2 => n11412, B1 => n9443, B2 => 
                           n5890, ZN => n9442);
   U12155 : BUF_X2 port map( I => n28616, Z => n314);
   U12164 : XOR2_X1 port map( A1 => n20447, A2 => n2824, Z => n29120);
   U12197 : NAND2_X2 port map( A1 => n36131, A2 => n36130, ZN => n34602);
   U12200 : NAND2_X2 port map( A1 => n11907, A2 => n20657, ZN => n24938);
   U12214 : OR2_X2 port map( A1 => n30853, A2 => n26832, Z => n26835);
   U12223 : NAND2_X2 port map( A1 => n25867, A2 => n26048, ZN => n26021);
   U12226 : XOR2_X1 port map( A1 => n6379, A2 => n34604, Z => n2394);
   U12227 : XOR2_X1 port map( A1 => n23669, A2 => n23668, Z => n34604);
   U12239 : NOR2_X2 port map( A1 => n27389, A2 => n21272, ZN => n20871);
   U12248 : NAND2_X1 port map( A1 => n20018, A2 => n35217, ZN => n15712);
   U12255 : XOR2_X1 port map( A1 => n27714, A2 => n184, Z => n183);
   U12256 : XOR2_X1 port map( A1 => n27525, A2 => n27834, Z => n27714);
   U12290 : NAND3_X2 port map( A1 => n7483, A2 => n28154, A3 => n17818, ZN => 
                           n31597);
   U12295 : NAND2_X2 port map( A1 => n33481, A2 => n18770, ZN => n17818);
   U12303 : NOR2_X1 port map( A1 => n35608, A2 => n39628, ZN => n34608);
   U12304 : NAND2_X2 port map( A1 => n10176, A2 => n399, ZN => n27724);
   U12332 : INV_X2 port map( I => n34610, ZN => n32080);
   U12346 : XOR2_X1 port map( A1 => n13116, A2 => n34611, Z => n19223);
   U12363 : NAND2_X1 port map( A1 => n30588, A2 => n19334, ZN => n30587);
   U12379 : NAND2_X2 port map( A1 => n34615, A2 => n4690, ZN => n23577);
   U12387 : XOR2_X1 port map( A1 => n34616, A2 => n11503, Z => n17210);
   U12404 : OAI22_X1 port map( A1 => n30257, A2 => n30259, B1 => n30262, B2 => 
                           n38204, ZN => n30263);
   U12407 : NAND2_X1 port map( A1 => n28543, A2 => n28739, ZN => n5969);
   U12416 : NAND2_X2 port map( A1 => n16530, A2 => n17522, ZN => n28543);
   U12421 : BUF_X2 port map( I => n18619, Z => n34620);
   U12426 : XOR2_X1 port map( A1 => n27527, A2 => n27567, Z => n15400);
   U12431 : XOR2_X1 port map( A1 => n15401, A2 => n8364, Z => n27567);
   U12453 : NAND2_X2 port map( A1 => n7469, A2 => n7468, ZN => n36200);
   U12463 : NAND2_X2 port map( A1 => n20768, A2 => n20770, ZN => n26585);
   U12479 : AOI21_X1 port map( A1 => n18780, A2 => n30014, B => n30034, ZN => 
                           n34622);
   U12491 : OAI22_X2 port map( A1 => n33234, A2 => n33235, B1 => n35495, B2 => 
                           n27419, ZN => n27737);
   U12504 : NOR2_X1 port map( A1 => n17632, A2 => n17240, ZN => n35063);
   U12507 : NAND2_X1 port map( A1 => n19312, A2 => n35063, ZN => n6921);
   U12516 : NAND2_X1 port map( A1 => n21897, A2 => n11576, ZN => n5733);
   U12520 : NOR2_X2 port map( A1 => n34627, A2 => n8635, ZN => n29044);
   U12541 : NAND2_X2 port map( A1 => n8399, A2 => n18457, ZN => n3263);
   U12542 : AOI22_X2 port map( A1 => n1820, A2 => n15712, B1 => n8918, B2 => 
                           n34761, ZN => n8399);
   U12552 : NAND3_X2 port map( A1 => n9237, A2 => n9236, A3 => n15727, ZN => 
                           n20445);
   U12554 : XOR2_X1 port map( A1 => n254, A2 => n39691, Z => n34630);
   U12557 : AND2_X1 port map( A1 => n20056, A2 => n18186, Z => n15694);
   U12565 : NAND2_X2 port map( A1 => n12852, A2 => n11007, ZN => n32208);
   U12566 : NAND2_X2 port map( A1 => n1159, A2 => n17242, ZN => n12852);
   U12589 : XOR2_X1 port map( A1 => n27827, A2 => n34634, Z => n19467);
   U12593 : XOR2_X1 port map( A1 => n27826, A2 => n11031, Z => n34634);
   U12599 : NOR2_X2 port map( A1 => n34357, A2 => n39194, ZN => n11468);
   U12605 : AOI22_X2 port map( A1 => n34639, A2 => n34638, B1 => n28378, B2 => 
                           n28098, ZN => n4197);
   U12608 : NAND2_X2 port map( A1 => n29011, A2 => n20219, ZN => n8287);
   U12610 : NOR2_X2 port map( A1 => n7855, A2 => n34641, ZN => n4847);
   U12618 : INV_X1 port map( I => n34642, ZN => n34641);
   U12622 : NOR2_X2 port map( A1 => n32326, A2 => n32327, ZN => n35715);
   U12625 : NAND3_X1 port map( A1 => n28246, A2 => n39399, A3 => n28115, ZN => 
                           n32413);
   U12627 : XOR2_X1 port map( A1 => n36379, A2 => n24009, Z => n24316);
   U12650 : NAND2_X2 port map( A1 => n6647, A2 => n1315, ZN => n14006);
   U12656 : XOR2_X1 port map( A1 => n29258, A2 => n34649, Z => n13288);
   U12664 : XOR2_X1 port map( A1 => n34650, A2 => n33313, Z => n10255);
   U12670 : OR2_X1 port map( A1 => n24383, A2 => n18402, Z => n6569);
   U12676 : NAND3_X2 port map( A1 => n18095, A2 => n1494, A3 => n20211, ZN => 
                           n20217);
   U12683 : OAI21_X2 port map( A1 => n979, A2 => n38075, B => n28570, ZN => 
                           n34651);
   U12687 : NAND2_X2 port map( A1 => n3253, A2 => n32430, ZN => n14374);
   U12691 : OAI22_X2 port map( A1 => n5075, A2 => n36457, B1 => n8204, B2 => 
                           n32889, ZN => n34654);
   U12692 : NOR2_X2 port map( A1 => n37187, A2 => n34655, ZN => n9581);
   U12693 : XOR2_X1 port map( A1 => n15532, A2 => n8671, Z => n8670);
   U12695 : XOR2_X1 port map( A1 => n22588, A2 => n5242, Z => n7137);
   U12699 : NAND2_X2 port map( A1 => n4497, A2 => n35193, ZN => n5242);
   U12700 : INV_X2 port map( I => n12718, ZN => n1190);
   U12701 : OAI21_X2 port map( A1 => n9850, A2 => n9684, B => n12420, ZN => 
                           n12718);
   U12709 : NAND2_X2 port map( A1 => n23308, A2 => n23607, ZN => n23413);
   U12711 : NAND2_X2 port map( A1 => n35715, A2 => n23007, ZN => n23308);
   U12716 : BUF_X2 port map( I => n11950, Z => n35404);
   U12731 : NAND2_X2 port map( A1 => n28427, A2 => n1194, ZN => n28394);
   U12746 : OR2_X1 port map( A1 => n1414, A2 => n2191, Z => n30740);
   U12749 : XOR2_X1 port map( A1 => n22723, A2 => n34663, Z => n4738);
   U12751 : XOR2_X1 port map( A1 => n15765, A2 => n22762, Z => n34663);
   U12769 : NAND2_X2 port map( A1 => n14924, A2 => n14926, ZN => n36750);
   U12776 : AOI22_X1 port map( A1 => n11022, A2 => n14512, B1 => n30263, B2 => 
                           n8691, ZN => n34778);
   U12789 : BUF_X2 port map( I => n2052, Z => n35253);
   U12793 : INV_X1 port map( I => n20865, ZN => n35879);
   U12804 : NAND2_X2 port map( A1 => n30689, A2 => n4485, ZN => n34717);
   U12808 : NAND2_X2 port map( A1 => n29885, A2 => n6720, ZN => n29880);
   U12823 : INV_X4 port map( I => n28033, ZN => n987);
   U12826 : AOI21_X2 port map( A1 => n30285, A2 => n26882, B => n37104, ZN => 
                           n34669);
   U12828 : OAI21_X2 port map( A1 => n34671, A2 => n34667, B => n34670, ZN => 
                           n28416);
   U12829 : INV_X1 port map( I => n28577, ZN => n34671);
   U12831 : XOR2_X1 port map( A1 => n20452, A2 => n34672, Z => n35633);
   U12835 : INV_X1 port map( I => n29399, ZN => n34672);
   U12856 : OR2_X1 port map( A1 => n18619, A2 => n12138, Z => n12801);
   U12866 : OAI22_X1 port map( A1 => n16513, A2 => n5469, B1 => n5470, B2 => 
                           n21239, ZN => n6588);
   U12869 : XOR2_X1 port map( A1 => n5289, A2 => n8473, Z => n12401);
   U12874 : OAI22_X2 port map( A1 => n19588, A2 => n14561, B1 => n15388, B2 => 
                           n4472, ZN => n15743);
   U12877 : XOR2_X1 port map( A1 => n11383, A2 => n23829, Z => n23943);
   U12885 : BUF_X2 port map( I => n22491, Z => n34678);
   U12886 : XOR2_X1 port map( A1 => n15448, A2 => n19717, Z => n22466);
   U12894 : XOR2_X1 port map( A1 => n30560, A2 => n34680, Z => n5351);
   U12896 : XOR2_X1 port map( A1 => n4266, A2 => n27825, Z => n34680);
   U12897 : OR2_X1 port map( A1 => n27624, A2 => n28153, Z => n9721);
   U12899 : OAI21_X2 port map( A1 => n16589, A2 => n30052, B => n34681, ZN => 
                           n18896);
   U12913 : XNOR2_X1 port map( A1 => n1859, A2 => n27701, ZN => n27089);
   U12918 : XOR2_X1 port map( A1 => n27633, A2 => n27799, Z => n27701);
   U12922 : NOR2_X2 port map( A1 => n1220, A2 => n31683, ZN => n34682);
   U12932 : AOI22_X1 port map( A1 => n31326, A2 => n29990, B1 => n4011, B2 => 
                           n30045, ZN => n30141);
   U12941 : NOR2_X2 port map( A1 => n8423, A2 => n28740, ZN => n1874);
   U12947 : XOR2_X1 port map( A1 => n27605, A2 => n31248, Z => n34686);
   U12949 : NAND2_X2 port map( A1 => n29189, A2 => n34688, ZN => n29754);
   U12951 : NAND2_X2 port map( A1 => n3248, A2 => n3250, ZN => n36913);
   U12954 : NOR2_X2 port map( A1 => n36246, A2 => n13820, ZN => n3248);
   U12966 : XOR2_X1 port map( A1 => n34691, A2 => n9719, Z => n22416);
   U12979 : OAI21_X2 port map( A1 => n11735, A2 => n4463, B => n4462, ZN => 
                           n27710);
   U12986 : XOR2_X1 port map( A1 => n23760, A2 => n16337, Z => n23761);
   U13010 : INV_X2 port map( I => n10986, ZN => n10724);
   U13022 : OAI21_X2 port map( A1 => n33973, A2 => n34696, B => n8806, ZN => 
                           n7577);
   U13028 : XOR2_X1 port map( A1 => n13840, A2 => n34697, Z => n12961);
   U13029 : XOR2_X1 port map( A1 => n13842, A2 => n34698, Z => n34697);
   U13041 : OR2_X1 port map( A1 => n690, A2 => n8736, Z => n20682);
   U13045 : INV_X2 port map( I => n34699, ZN => n15839);
   U13046 : XOR2_X1 port map( A1 => Plaintext(92), A2 => Key(92), Z => n34699);
   U13049 : NAND3_X2 port map( A1 => n13137, A2 => n12473, A3 => n12472, ZN => 
                           n23423);
   U13054 : OR2_X1 port map( A1 => n22354, A2 => n22353, Z => n22209);
   U13062 : NAND2_X2 port map( A1 => n27004, A2 => n35914, ZN => n27834);
   U13072 : NOR2_X1 port map( A1 => n19364, A2 => n26879, ZN => n26609);
   U13082 : NAND2_X2 port map( A1 => n19413, A2 => n35124, ZN => n4232);
   U13094 : NAND2_X1 port map( A1 => n22051, A2 => n22307, ZN => n30613);
   U13101 : XOR2_X1 port map( A1 => n19355, A2 => n27729, Z => n31204);
   U13106 : NAND2_X2 port map( A1 => n18073, A2 => n18075, ZN => n27729);
   U13108 : XOR2_X1 port map( A1 => n9511, A2 => n22641, Z => n34703);
   U13109 : INV_X1 port map( I => n39194, ZN => n9924);
   U13110 : OR2_X1 port map( A1 => n39194, A2 => n12966, Z => n17958);
   U13114 : XOR2_X1 port map( A1 => n10812, A2 => n10811, Z => n29174);
   U13115 : XOR2_X1 port map( A1 => n7004, A2 => n29082, Z => n10811);
   U13123 : XOR2_X1 port map( A1 => n34709, A2 => n34708, Z => n14641);
   U13125 : XOR2_X1 port map( A1 => n31438, A2 => n27815, Z => n34709);
   U13136 : NAND2_X2 port map( A1 => n34711, A2 => n34210, ZN => n34820);
   U13142 : NAND2_X2 port map( A1 => n23596, A2 => n23595, ZN => n3006);
   U13145 : AOI21_X2 port map( A1 => n36701, A2 => n36011, B => n1160, ZN => 
                           n12821);
   U13148 : XOR2_X1 port map( A1 => n34712, A2 => n26417, Z => n33473);
   U13181 : AOI21_X2 port map( A1 => n22956, A2 => n34457, B => n34716, ZN => 
                           n5619);
   U13188 : BUF_X2 port map( I => n22561, Z => n34718);
   U13197 : AOI22_X2 port map( A1 => n11528, A2 => n1038, B1 => n17454, B2 => 
                           n23515, ZN => n13978);
   U13213 : XOR2_X1 port map( A1 => n14986, A2 => n8182, Z => n8181);
   U13227 : XOR2_X1 port map( A1 => n7402, A2 => n31791, Z => n8902);
   U13244 : XOR2_X1 port map( A1 => n26356, A2 => n18004, Z => n14784);
   U13248 : OAI21_X2 port map( A1 => n5508, A2 => n32052, B => n32051, ZN => 
                           n18004);
   U13254 : XOR2_X1 port map( A1 => n6943, A2 => n6940, Z => n35242);
   U13257 : NOR2_X2 port map( A1 => n7423, A2 => n26120, ZN => n26013);
   U13262 : XOR2_X1 port map( A1 => n12383, A2 => n8310, Z => n34722);
   U13268 : INV_X1 port map( I => n34723, ZN => n24786);
   U13270 : NOR2_X1 port map( A1 => n35686, A2 => n37016, ZN => n34723);
   U13290 : XOR2_X1 port map( A1 => n19342, A2 => n34724, Z => n13694);
   U13296 : XOR2_X1 port map( A1 => n13844, A2 => n32420, Z => n34724);
   U13321 : XOR2_X1 port map( A1 => n35554, A2 => n20684, Z => n170);
   U13322 : NAND2_X2 port map( A1 => n25900, A2 => n25801, ZN => n25751);
   U13324 : XOR2_X1 port map( A1 => n34728, A2 => n37129, Z => n5520);
   U13326 : XOR2_X1 port map( A1 => n27554, A2 => n1703, Z => n34728);
   U13333 : NAND2_X2 port map( A1 => n37031, A2 => n2883, ZN => n3528);
   U13347 : NOR2_X1 port map( A1 => n11658, A2 => n11582, ZN => n11659);
   U13348 : XOR2_X1 port map( A1 => n2594, A2 => n26395, Z => n36719);
   U13351 : XOR2_X1 port map( A1 => n39078, A2 => n7439, Z => n26395);
   U13384 : OAI21_X2 port map( A1 => n34747, A2 => n34746, B => n24843, ZN => 
                           n3629);
   U13387 : AOI21_X1 port map( A1 => n16803, A2 => n29890, B => n10848, ZN => 
                           n17527);
   U13388 : INV_X2 port map( I => n6720, ZN => n10848);
   U13389 : XOR2_X1 port map( A1 => n10987, A2 => n30733, Z => n6457);
   U13407 : NAND3_X1 port map( A1 => n36789, A2 => n36790, A3 => n16377, ZN => 
                           n36267);
   U13409 : XOR2_X1 port map( A1 => n9979, A2 => n7185, Z => n31773);
   U13411 : XOR2_X1 port map( A1 => n11372, A2 => n29141, Z => n562);
   U13418 : NAND2_X2 port map( A1 => n24089, A2 => n34750, ZN => n24879);
   U13422 : OAI21_X2 port map( A1 => n34751, A2 => n19349, B => n7480, ZN => 
                           n18364);
   U13429 : XOR2_X1 port map( A1 => n2096, A2 => n30489, Z => n2094);
   U13434 : XOR2_X1 port map( A1 => n38201, A2 => n19862, Z => n30519);
   U13448 : BUF_X4 port map( I => n27575, Z => n28290);
   U13456 : XOR2_X1 port map( A1 => n26288, A2 => n26287, Z => n34752);
   U13482 : NOR3_X1 port map( A1 => n35253, A2 => n18402, A3 => n24382, ZN => 
                           n34758);
   U13488 : XNOR2_X1 port map( A1 => n15219, A2 => n27574, ZN => n27677);
   U13495 : XOR2_X1 port map( A1 => n34760, A2 => n34056, Z => n33347);
   U13497 : XOR2_X1 port map( A1 => n27643, A2 => n27497, Z => n34760);
   U13504 : AND2_X1 port map( A1 => n27341, A2 => n27338, Z => n4668);
   U13518 : AOI22_X2 port map( A1 => n27909, A2 => n28298, B1 => n28268, B2 => 
                           n28301, ZN => n28790);
   U13522 : OAI22_X2 port map( A1 => n27907, A2 => n28753, B1 => n16303, B2 => 
                           n27908, ZN => n28268);
   U13523 : XOR2_X1 port map( A1 => n20571, A2 => n19809, Z => n25694);
   U13525 : XOR2_X1 port map( A1 => n27769, A2 => n27798, Z => n2758);
   U13531 : AOI22_X2 port map( A1 => n35417, A2 => n35694, B1 => n37056, B2 => 
                           n28004, ZN => n34762);
   U13539 : INV_X4 port map( I => n11867, ZN => n5130);
   U13542 : XOR2_X1 port map( A1 => n248, A2 => n15270, Z => n28867);
   U13545 : NAND2_X2 port map( A1 => n10148, A2 => n34763, ZN => n33813);
   U13548 : INV_X2 port map( I => n34764, ZN => n31669);
   U13566 : XOR2_X1 port map( A1 => n3649, A2 => n34766, Z => n9033);
   U13569 : OAI21_X1 port map( A1 => n9032, A2 => n12846, B => n9031, ZN => 
                           n34766);
   U13575 : XOR2_X1 port map( A1 => n26548, A2 => n26541, Z => n34878);
   U13586 : AOI22_X2 port map( A1 => n34767, A2 => n20423, B1 => n26973, B2 => 
                           n16000, ZN => n15999);
   U13612 : XOR2_X1 port map( A1 => n8364, A2 => n27781, Z => n27718);
   U13638 : OR3_X1 port map( A1 => n17410, A2 => n988, A3 => n13081, Z => 
                           n27976);
   U13640 : NAND2_X1 port map( A1 => n29396, A2 => n19157, ZN => n29398);
   U13652 : OAI21_X2 port map( A1 => n20651, A2 => n34772, B => n23197, ZN => 
                           n13982);
   U13664 : XOR2_X1 port map( A1 => n28876, A2 => n35633, Z => n34773);
   U13669 : OAI22_X2 port map( A1 => n8347, A2 => n29700, B1 => n8346, B2 => 
                           n8345, ZN => n18042);
   U13671 : XOR2_X1 port map( A1 => n35637, A2 => n7714, Z => n35636);
   U13673 : OAI21_X2 port map( A1 => n10038, A2 => n5641, B => n10906, ZN => 
                           n34774);
   U13680 : XOR2_X1 port map( A1 => n27804, A2 => n27802, Z => n15994);
   U13681 : XOR2_X1 port map( A1 => n1466, A2 => n36384, Z => n27804);
   U13697 : NAND2_X1 port map( A1 => n31647, A2 => n36424, ZN => n8820);
   U13698 : XOR2_X1 port map( A1 => n34778, A2 => n16562, Z => Ciphertext(187))
                           ;
   U13726 : AOI21_X2 port map( A1 => n37065, A2 => n24120, B => n5854, ZN => 
                           n24753);
   U13727 : XOR2_X1 port map( A1 => n34780, A2 => n28973, Z => n28975);
   U13728 : XOR2_X1 port map( A1 => n28972, A2 => n39220, Z => n34780);
   U13735 : OAI21_X2 port map( A1 => n34105, A2 => n33125, B => n33705, ZN => 
                           n24672);
   U13740 : XOR2_X1 port map( A1 => n10854, A2 => n10855, Z => n853);
   U13741 : XOR2_X1 port map( A1 => n28977, A2 => n29125, Z => n16359);
   U13767 : AOI21_X2 port map( A1 => n28314, A2 => n31045, B => n4926, ZN => 
                           n28972);
   U13774 : XOR2_X1 port map( A1 => n22405, A2 => n7432, Z => n6474);
   U13787 : NAND2_X1 port map( A1 => n34357, A2 => n39194, ZN => n32068);
   U13795 : NOR2_X2 port map( A1 => n21725, A2 => n4913, ZN => n36281);
   U13800 : INV_X2 port map( I => n20605, ZN => n1564);
   U13815 : AOI22_X2 port map( A1 => n23038, A2 => n23540, B1 => n6301, B2 => 
                           n18746, ZN => n23686);
   U13830 : XOR2_X1 port map( A1 => n32776, A2 => n24052, Z => n18683);
   U13833 : NAND2_X1 port map( A1 => n34842, A2 => n27081, ZN => n34841);
   U13866 : XOR2_X1 port map( A1 => n10540, A2 => n34785, Z => n31978);
   U13870 : XOR2_X1 port map( A1 => n10538, A2 => n10539, Z => n34785);
   U13881 : NAND2_X2 port map( A1 => n36425, A2 => n37775, ZN => n15268);
   U13882 : INV_X2 port map( I => n9218, ZN => n259);
   U13908 : XOR2_X1 port map( A1 => n6719, A2 => n5542, Z => n34787);
   U13922 : OR2_X1 port map( A1 => n7387, A2 => n38724, Z => n34924);
   U13924 : XOR2_X1 port map( A1 => n16138, A2 => n23900, Z => n18857);
   U13927 : OAI22_X2 port map( A1 => n23508, A2 => n13829, B1 => n13832, B2 => 
                           n13831, ZN => n16138);
   U13931 : XOR2_X1 port map( A1 => n35987, A2 => n34999, Z => n11230);
   U13934 : XOR2_X1 port map( A1 => n34789, A2 => n35112, Z => n34999);
   U13938 : NAND2_X1 port map( A1 => n14428, A2 => n21270, ZN => n19704);
   U13957 : NAND3_X2 port map( A1 => n27873, A2 => n27872, A3 => n27871, ZN => 
                           n13601);
   U13973 : XOR2_X1 port map( A1 => n22742, A2 => n8312, Z => n22551);
   U13979 : OAI21_X1 port map( A1 => n5977, A2 => n29701, B => n20982, ZN => 
                           n34793);
   U13981 : AOI21_X2 port map( A1 => n13780, A2 => n35182, B => n11164, ZN => 
                           n5757);
   U13984 : OAI21_X1 port map( A1 => n29758, A2 => n19348, B => n34795, ZN => 
                           n29759);
   U13992 : OAI21_X1 port map( A1 => n34182, A2 => n29753, B => n29756, ZN => 
                           n34795);
   U14052 : AOI22_X2 port map( A1 => n3935, A2 => n37103, B1 => n3961, B2 => 
                           n1494, ZN => n34799);
   U14077 : XOR2_X1 port map( A1 => n31314, A2 => n10579, Z => n34800);
   U14080 : AOI21_X2 port map( A1 => n15024, A2 => n12653, B => n89, ZN => 
                           n34801);
   U14081 : XOR2_X1 port map( A1 => n34802, A2 => n32773, Z => n35896);
   U14093 : XNOR2_X1 port map( A1 => n37593, A2 => n26599, ZN => n26419);
   U14098 : AOI21_X2 port map( A1 => n17144, A2 => n26975, B => n17143, ZN => 
                           n27325);
   U14103 : NAND2_X2 port map( A1 => n2946, A2 => n35499, ZN => n36555);
   U14118 : XOR2_X1 port map( A1 => n19428, A2 => n21095, Z => n34809);
   U14119 : NAND2_X1 port map( A1 => n9169, A2 => n28004, ZN => n27893);
   U14121 : NAND2_X2 port map( A1 => n35666, A2 => n3307, ZN => n15467);
   U14143 : NAND2_X2 port map( A1 => n2341, A2 => n19422, ZN => n24663);
   U14144 : NAND2_X2 port map( A1 => n20229, A2 => n20227, ZN => n19422);
   U14162 : XOR2_X1 port map( A1 => n39536, A2 => n29838, Z => n29839);
   U14180 : NAND2_X2 port map( A1 => n5439, A2 => n5438, ZN => n5089);
   U14182 : NOR2_X1 port map( A1 => n2965, A2 => n32168, ZN => n36682);
   U14183 : XOR2_X1 port map( A1 => n33868, A2 => n34814, Z => n36063);
   U14184 : XOR2_X1 port map( A1 => n3317, A2 => n34815, Z => n34814);
   U14189 : INV_X1 port map( I => n1612, ZN => n34815);
   U14195 : NAND2_X2 port map( A1 => n14916, A2 => n23329, ZN => n23783);
   U14199 : XOR2_X1 port map( A1 => n25039, A2 => n25213, Z => n13920);
   U14200 : NAND2_X2 port map( A1 => n26056, A2 => n26089, ZN => n25882);
   U14223 : XOR2_X1 port map( A1 => n33735, A2 => n6154, Z => n2594);
   U14224 : INV_X2 port map( I => n36579, ZN => n33735);
   U14238 : NAND2_X2 port map( A1 => n927, A2 => n26090, ZN => n13502);
   U14244 : AOI21_X2 port map( A1 => n31345, A2 => n22969, B => n13157, ZN => 
                           n13370);
   U14251 : XOR2_X1 port map( A1 => n4269, A2 => n4271, Z => n10071);
   U14258 : XOR2_X1 port map( A1 => n8909, A2 => n34825, Z => n3297);
   U14261 : XOR2_X1 port map( A1 => n3299, A2 => n9106, Z => n34825);
   U14263 : NAND3_X2 port map( A1 => n32586, A2 => n34826, A3 => n2418, ZN => 
                           n11752);
   U14270 : NOR2_X2 port map( A1 => n12329, A2 => n37166, ZN => n14729);
   U14272 : INV_X2 port map( I => n34828, ZN => n14080);
   U14280 : NAND2_X2 port map( A1 => n1577, A2 => n8966, ZN => n13221);
   U14285 : XOR2_X1 port map( A1 => n22529, A2 => n22594, Z => n22771);
   U14286 : NOR2_X2 port map( A1 => n6199, A2 => n33594, ZN => n22529);
   U14289 : OAI21_X2 port map( A1 => n34830, A2 => n26822, B => n14798, ZN => 
                           n34969);
   U14303 : OR2_X1 port map( A1 => n14377, A2 => n26761, Z => n26758);
   U14304 : AND2_X1 port map( A1 => n39112, A2 => n28224, Z => n7326);
   U14308 : INV_X2 port map( I => n26224, ZN => n17048);
   U14309 : NAND2_X2 port map( A1 => n25112, A2 => n18864, ZN => n26224);
   U14310 : OAI21_X1 port map( A1 => n24607, A2 => n12846, B => n29285, ZN => 
                           n9031);
   U14313 : NOR2_X1 port map( A1 => n17451, A2 => n37553, ZN => n36488);
   U14327 : NAND2_X2 port map( A1 => n11631, A2 => n11630, ZN => n24745);
   U14333 : XOR2_X1 port map( A1 => n6384, A2 => n8303, Z => n28842);
   U14337 : NAND2_X2 port map( A1 => n26678, A2 => n34837, ZN => n27436);
   U14339 : NAND3_X1 port map( A1 => n26823, A2 => n20021, A3 => n37643, ZN => 
                           n34837);
   U14342 : NAND2_X2 port map( A1 => n34838, A2 => n18350, ZN => n14808);
   U14343 : OAI21_X2 port map( A1 => n17390, A2 => n27973, B => n28156, ZN => 
                           n34871);
   U14348 : NOR2_X2 port map( A1 => n21239, A2 => n28290, ZN => n27973);
   U14349 : NOR2_X1 port map( A1 => n34841, A2 => n34840, ZN => n10336);
   U14352 : NOR2_X1 port map( A1 => n27164, A2 => n35750, ZN => n34840);
   U14363 : NAND2_X1 port map( A1 => n25849, A2 => n34350, ZN => n25851);
   U14368 : NAND2_X2 port map( A1 => n35327, A2 => n25376, ZN => n25849);
   U14371 : INV_X2 port map( I => n3863, ZN => n36745);
   U14375 : INV_X2 port map( I => n20646, ZN => n22365);
   U14377 : NAND4_X2 port map( A1 => n14912, A2 => n16654, A3 => n16653, A4 => 
                           n34997, ZN => n20646);
   U14382 : NAND3_X1 port map( A1 => n19666, A2 => n39261, A3 => n34924, ZN => 
                           n32487);
   U14395 : XOR2_X1 port map( A1 => n38269, A2 => n34848, Z => n744);
   U14398 : INV_X1 port map( I => n19925, ZN => n34848);
   U14401 : OAI21_X2 port map( A1 => n19215, A2 => n34402, B => n19214, ZN => 
                           n25659);
   U14402 : XOR2_X1 port map( A1 => n3090, A2 => n35350, Z => n36617);
   U14411 : XOR2_X1 port map( A1 => n16284, A2 => n34849, Z => n17084);
   U14412 : XOR2_X1 port map( A1 => n23936, A2 => n35752, Z => n34849);
   U14417 : XOR2_X1 port map( A1 => n19577, A2 => n34850, Z => n20207);
   U14418 : XOR2_X1 port map( A1 => n23793, A2 => n34851, Z => n34850);
   U14431 : XOR2_X1 port map( A1 => n33693, A2 => n34854, Z => n8628);
   U14434 : XOR2_X1 port map( A1 => n8629, A2 => n22560, Z => n34854);
   U14435 : NAND2_X2 port map( A1 => n31325, A2 => n22826, ZN => n34959);
   U14440 : NAND3_X1 port map( A1 => n33565, A2 => n35187, A3 => n30106, ZN => 
                           n34855);
   U14456 : XOR2_X1 port map( A1 => n5586, A2 => n2543, Z => n36884);
   U14457 : NAND2_X2 port map( A1 => n4682, A2 => n12952, ZN => n22880);
   U14507 : NOR2_X2 port map( A1 => n20761, A2 => n15441, ZN => n30800);
   U14510 : NAND2_X2 port map( A1 => n38666, A2 => n18673, ZN => n34863);
   U14514 : NAND2_X2 port map( A1 => n580, A2 => n1202, ZN => n34866);
   U14530 : INV_X1 port map( I => n21735, ZN => n34867);
   U14531 : NAND2_X1 port map( A1 => n34867, A2 => n293, ZN => n20762);
   U14532 : XOR2_X1 port map( A1 => n34869, A2 => n6739, Z => n11948);
   U14533 : XOR2_X1 port map( A1 => n35711, A2 => n26172, Z => n34869);
   U14534 : XOR2_X1 port map( A1 => n22595, A2 => n22594, Z => n11190);
   U14535 : NOR2_X2 port map( A1 => n13296, A2 => n22087, ZN => n22595);
   U14541 : AOI22_X2 port map( A1 => n34870, A2 => n11128, B1 => n8008, B2 => 
                           n1417, ZN => n29819);
   U14543 : NAND3_X1 port map( A1 => n21949, A2 => n21945, A3 => n21784, ZN => 
                           n35623);
   U14569 : NAND2_X1 port map( A1 => n36134, A2 => n36132, ZN => n34877);
   U14572 : XOR2_X1 port map( A1 => n26297, A2 => n34024, Z => n36257);
   U14573 : NOR2_X1 port map( A1 => n36296, A2 => n19886, ZN => n3627);
   U14574 : INV_X4 port map( I => n24557, ZN => n19886);
   U14578 : AOI21_X2 port map( A1 => n36725, A2 => n16644, B => n808, ZN => 
                           n24557);
   U14580 : XOR2_X1 port map( A1 => n21034, A2 => n26545, Z => n13914);
   U14586 : XOR2_X1 port map( A1 => n26455, A2 => n35627, Z => n21034);
   U14588 : XOR2_X1 port map( A1 => n10668, A2 => n34878, Z => n3976);
   U14602 : AOI21_X2 port map( A1 => n29866, A2 => n31545, B => n34882, ZN => 
                           n29883);
   U14604 : NOR2_X1 port map( A1 => n15521, A2 => n16059, ZN => n34882);
   U14616 : OAI21_X2 port map( A1 => n32233, A2 => n32232, B => n34885, ZN => 
                           n26448);
   U14622 : NAND3_X2 port map( A1 => n3434, A2 => n38168, A3 => n32243, ZN => 
                           n34885);
   U14625 : NAND2_X2 port map( A1 => n12650, A2 => n17541, ZN => n16054);
   U14628 : NAND2_X2 port map( A1 => n34886, A2 => n10972, ZN => n25820);
   U14630 : AND2_X1 port map( A1 => n23582, A2 => n23580, Z => n22806);
   U14632 : NAND2_X2 port map( A1 => n8460, A2 => n4698, ZN => n23582);
   U14633 : NOR2_X1 port map( A1 => n5541, A2 => n9740, ZN => n12557);
   U14634 : INV_X2 port map( I => n5518, ZN => n5541);
   U14640 : NAND2_X1 port map( A1 => n3916, A2 => n39676, ZN => n34939);
   U14642 : XOR2_X1 port map( A1 => n9221, A2 => n9219, Z => n14306);
   U14662 : NAND2_X2 port map( A1 => n3076, A2 => n24877, ZN => n24749);
   U14676 : NAND2_X2 port map( A1 => n34890, A2 => n34889, ZN => n6847);
   U14677 : NAND2_X2 port map( A1 => n34891, A2 => n8087, ZN => n36791);
   U14701 : NAND2_X1 port map( A1 => n11306, A2 => n13801, ZN => n34897);
   U14724 : XOR2_X1 port map( A1 => n10253, A2 => n34900, Z => n36264);
   U14725 : XOR2_X1 port map( A1 => n23774, A2 => n23976, Z => n10253);
   U14728 : NAND2_X2 port map( A1 => n7882, A2 => n24246, ZN => n34906);
   U14739 : XOR2_X1 port map( A1 => n25256, A2 => n25116, Z => n34901);
   U14748 : OAI21_X2 port map( A1 => n33365, A2 => n25743, B => n38899, ZN => 
                           n14253);
   U14762 : XOR2_X1 port map( A1 => n23884, A2 => n23774, Z => n23696);
   U14772 : NAND2_X1 port map( A1 => n30066, A2 => n30078, ZN => n3947);
   U14782 : INV_X2 port map( I => n15697, ZN => n36731);
   U14789 : XOR2_X1 port map( A1 => n35998, A2 => n19760, Z => n8908);
   U14796 : XOR2_X1 port map( A1 => n19772, A2 => n8074, Z => n26713);
   U14798 : AOI22_X2 port map( A1 => n1872, A2 => n15163, B1 => n36553, B2 => 
                           n22944, ZN => n10472);
   U14806 : OAI21_X2 port map( A1 => n32795, A2 => n6689, B => n34909, ZN => 
                           n9184);
   U14807 : NAND3_X1 port map( A1 => n27737, A2 => n27346, A3 => n27345, ZN => 
                           n34909);
   U14812 : OAI22_X2 port map( A1 => n6483, A2 => n33354, B1 => n34080, B2 => 
                           n18238, ZN => n24585);
   U14815 : INV_X2 port map( I => n7317, ZN => n33871);
   U14829 : INV_X2 port map( I => n14212, ZN => n25764);
   U14839 : XOR2_X1 port map( A1 => n10195, A2 => n34912, Z => n25631);
   U14841 : XOR2_X1 port map( A1 => n25264, A2 => n25265, Z => n34912);
   U14846 : BUF_X2 port map( I => n26625, Z => n26219);
   U14859 : NAND2_X1 port map( A1 => n30636, A2 => n32769, ZN => n36313);
   U14861 : AND2_X1 port map( A1 => n23907, A2 => n24244, Z => n9384);
   U14865 : NOR2_X2 port map( A1 => n4973, A2 => n34906, ZN => n3793);
   U14874 : XOR2_X1 port map( A1 => n25270, A2 => n9624, Z => n20416);
   U14876 : INV_X2 port map( I => n26807, ZN => n34913);
   U14881 : BUF_X2 port map( I => n33964, Z => n34914);
   U14884 : XOR2_X1 port map( A1 => n26517, A2 => n26602, Z => n26257);
   U14885 : NOR2_X2 port map( A1 => n6400, A2 => n6401, ZN => n26517);
   U14896 : OAI21_X2 port map( A1 => n26937, A2 => n32745, B => n34918, ZN => 
                           n26940);
   U14898 : NAND2_X1 port map( A1 => n10896, A2 => n17198, ZN => n18120);
   U14908 : OAI21_X2 port map( A1 => n6129, A2 => n1680, B => n5232, ZN => 
                           n5231);
   U14910 : NOR2_X2 port map( A1 => n6128, A2 => n22295, ZN => n6129);
   U14914 : OAI21_X2 port map( A1 => n21941, A2 => n4084, B => n36519, ZN => 
                           n36518);
   U14916 : NOR2_X2 port map( A1 => n34923, A2 => n34922, ZN => n21941);
   U14927 : NOR2_X2 port map( A1 => n34926, A2 => n34925, ZN => n17882);
   U14932 : NOR2_X2 port map( A1 => n17970, A2 => n33091, ZN => n34926);
   U14942 : AOI22_X2 port map( A1 => n20593, A2 => n15523, B1 => n15522, B2 => 
                           n17763, ZN => n1812);
   U14952 : XOR2_X1 port map( A1 => n35741, A2 => n12871, Z => n36717);
   U14953 : XOR2_X1 port map( A1 => n22004, A2 => n22003, Z => n22005);
   U14957 : XOR2_X1 port map( A1 => n29255, A2 => n6536, Z => n4461);
   U14960 : NAND2_X1 port map( A1 => n13579, A2 => n13578, ZN => n35483);
   U14979 : NAND3_X2 port map( A1 => n26979, A2 => n11864, A3 => n12290, ZN => 
                           n34930);
   U14983 : NOR3_X2 port map( A1 => n34932, A2 => n34931, A3 => n3480, ZN => 
                           n35399);
   U14995 : XOR2_X1 port map( A1 => n22615, A2 => n8552, Z => n20668);
   U14996 : NOR2_X2 port map( A1 => n9486, A2 => n9484, ZN => n8552);
   U15002 : XOR2_X1 port map( A1 => n3454, A2 => n23429, Z => n36500);
   U15005 : AND2_X1 port map( A1 => n5337, A2 => n12952, Z => n5834);
   U15006 : NAND2_X2 port map( A1 => n6576, A2 => n5077, ZN => n22359);
   U15014 : OAI21_X2 port map( A1 => n30272, A2 => n36368, B => n37335, ZN => 
                           n109);
   U15016 : NOR2_X1 port map( A1 => n39405, A2 => n9197, ZN => n34934);
   U15017 : NAND2_X1 port map( A1 => n33541, A2 => n35137, ZN => n34935);
   U15025 : NOR2_X2 port map( A1 => n1962, A2 => n20673, ZN => n2559);
   U15026 : BUF_X4 port map( I => n3927, Z => n1823);
   U15030 : NAND2_X1 port map( A1 => n24460, A2 => n19466, ZN => n34938);
   U15032 : OR2_X1 port map( A1 => n29755, A2 => n29754, Z => n29735);
   U15034 : NOR2_X2 port map( A1 => n23518, A2 => n23517, ZN => n18475);
   U15046 : AOI21_X1 port map( A1 => n12230, A2 => n4239, B => n13778, ZN => 
                           n35979);
   U15049 : NAND2_X2 port map( A1 => n25400, A2 => n36678, ZN => n34940);
   U15051 : XOR2_X1 port map( A1 => n2582, A2 => n13883, Z => n33112);
   U15052 : XOR2_X1 port map( A1 => n34332, A2 => n27828, Z => n2582);
   U15059 : AOI22_X2 port map( A1 => n937, A2 => n30306, B1 => n17411, B2 => 
                           n12077, ZN => n22333);
   U15063 : XOR2_X1 port map( A1 => n12551, A2 => n31355, Z => n15844);
   U15088 : XOR2_X1 port map( A1 => n27823, A2 => n34945, Z => n754);
   U15092 : INV_X1 port map( I => n19820, ZN => n34945);
   U15109 : OAI21_X2 port map( A1 => n21170, A2 => n21169, B => n17697, ZN => 
                           n27823);
   U15112 : XOR2_X1 port map( A1 => n23755, A2 => n23728, Z => n24013);
   U15116 : NAND2_X2 port map( A1 => n23633, A2 => n23632, ZN => n23728);
   U15143 : INV_X2 port map( I => n36500, ZN => n18116);
   U15145 : OAI21_X2 port map( A1 => n37163, A2 => n12435, B => n12793, ZN => 
                           n34953);
   U15161 : XOR2_X1 port map( A1 => n22370, A2 => n22372, Z => n34955);
   U15167 : INV_X1 port map( I => n17964, ZN => n35073);
   U15172 : INV_X2 port map( I => n34956, ZN => n10004);
   U15188 : NOR2_X2 port map( A1 => n17041, A2 => n21800, ZN => n22622);
   U15190 : INV_X1 port map( I => n18500, ZN => n4748);
   U15192 : NAND2_X1 port map( A1 => n34957, A2 => n18500, ZN => n26930);
   U15193 : XOR2_X1 port map( A1 => n4853, A2 => n26555, Z => n18500);
   U15200 : INV_X2 port map( I => n8966, ZN => n1579);
   U15209 : NAND2_X2 port map( A1 => n34964, A2 => n35057, ZN => n30174);
   U15210 : NAND2_X2 port map( A1 => n31065, A2 => n30196, ZN => n34964);
   U15219 : NOR2_X1 port map( A1 => n16180, A2 => n35187, ZN => n16277);
   U15226 : XOR2_X1 port map( A1 => n21085, A2 => n34966, Z => n26885);
   U15230 : NAND2_X2 port map( A1 => n15082, A2 => n15079, ZN => n10143);
   U15232 : XOR2_X1 port map( A1 => n26376, A2 => n26490, Z => n20656);
   U15238 : OR2_X1 port map( A1 => n35693, A2 => n24735, Z => n10115);
   U15244 : NAND2_X1 port map( A1 => n34217, A2 => n35003, ZN => n34967);
   U15245 : NOR2_X1 port map( A1 => n9963, A2 => n14379, ZN => n14630);
   U15262 : NAND2_X2 port map( A1 => n34972, A2 => n12345, ZN => n13564);
   U15264 : XOR2_X1 port map( A1 => n16797, A2 => n23848, Z => n16795);
   U15289 : INV_X2 port map( I => n29535, ZN => n32317);
   U15300 : XOR2_X1 port map( A1 => n22439, A2 => n31566, Z => n35457);
   U15311 : NOR2_X1 port map( A1 => n7804, A2 => n12630, ZN => n34979);
   U15326 : NAND2_X2 port map( A1 => n13785, A2 => n31379, ZN => n22710);
   U15332 : NAND2_X2 port map( A1 => n2900, A2 => n2899, ZN => n18305);
   U15342 : XOR2_X1 port map( A1 => n25238, A2 => n25298, Z => n25028);
   U15350 : NOR2_X2 port map( A1 => n36110, A2 => n33629, ZN => n36109);
   U15354 : OAI21_X2 port map( A1 => n35028, A2 => n1489, B => n37955, ZN => 
                           n34982);
   U15355 : INV_X4 port map( I => n12168, ZN => n12237);
   U15358 : NOR2_X2 port map( A1 => n11885, A2 => n15605, ZN => n34983);
   U15364 : NOR2_X2 port map( A1 => n12497, A2 => n12498, ZN => n34984);
   U15366 : NAND3_X1 port map( A1 => n1174, A2 => n31569, A3 => n29927, ZN => 
                           n29916);
   U15368 : OAI22_X2 port map( A1 => n34985, A2 => n8587, B1 => n37955, B2 => 
                           n15371, ZN => n17795);
   U15381 : NOR2_X2 port map( A1 => n9805, A2 => n7624, ZN => n24819);
   U15383 : AOI21_X2 port map( A1 => n37144, A2 => n1475, B => n34990, ZN => 
                           n34989);
   U15389 : XOR2_X1 port map( A1 => n4315, A2 => n34993, Z => n4392);
   U15393 : XOR2_X1 port map( A1 => n4313, A2 => n29129, Z => n34993);
   U15395 : AND2_X1 port map( A1 => n28659, A2 => n8366, Z => n6043);
   U15409 : NAND2_X2 port map( A1 => n26075, A2 => n7660, ZN => n26077);
   U15412 : NOR2_X2 port map( A1 => n7874, A2 => n7877, ZN => n7660);
   U15418 : NAND2_X1 port map( A1 => n11497, A2 => n32419, ZN => n11495);
   U15425 : BUF_X2 port map( I => n8972, Z => n33083);
   U15431 : NOR2_X2 port map( A1 => n35470, A2 => n789, ZN => n5323);
   U15440 : OAI22_X2 port map( A1 => n3359, A2 => n20456, B1 => n30644, B2 => 
                           n3356, ZN => n35646);
   U15447 : XOR2_X1 port map( A1 => n18557, A2 => n18556, Z => n21150);
   U15449 : NAND2_X2 port map( A1 => n6078, A2 => n2451, ZN => n6077);
   U15452 : NAND3_X1 port map( A1 => n21844, A2 => n6198, A3 => n18219, ZN => 
                           n34997);
   U15456 : XOR2_X1 port map( A1 => n34999, A2 => n11967, Z => n34998);
   U15468 : NAND2_X1 port map( A1 => n31799, A2 => n1435, ZN => n3844);
   U15482 : NAND3_X2 port map( A1 => n9204, A2 => n20792, A3 => n9203, ZN => 
                           n4353);
   U15487 : NAND2_X2 port map( A1 => n36094, A2 => n3813, ZN => n21068);
   U15498 : AOI21_X2 port map( A1 => n29150, A2 => n4858, B => n29899, ZN => 
                           n19539);
   U15499 : NAND3_X1 port map( A1 => n34007, A2 => n32146, A3 => n974, ZN => 
                           n4857);
   U15503 : INV_X2 port map( I => n36496, ZN => n1472);
   U15512 : XOR2_X1 port map( A1 => n18796, A2 => n33131, Z => n26795);
   U15518 : NOR2_X2 port map( A1 => n3010, A2 => n3011, ZN => n36967);
   U15533 : XOR2_X1 port map( A1 => n27592, A2 => n35334, Z => n27593);
   U15538 : NOR2_X2 port map( A1 => n35791, A2 => n35792, ZN => n35006);
   U15560 : XOR2_X1 port map( A1 => n5965, A2 => n35010, Z => n302);
   U15562 : XOR2_X1 port map( A1 => n9490, A2 => n33388, Z => n35010);
   U15563 : AND2_X1 port map( A1 => n39564, A2 => n5960, Z => n10565);
   U15577 : AOI21_X2 port map( A1 => n34129, A2 => n23480, B => n35013, ZN => 
                           n35012);
   U15588 : NAND2_X2 port map( A1 => n1045, A2 => n16104, ZN => n35016);
   U15590 : NAND2_X1 port map( A1 => n35655, A2 => n20530, ZN => n36598);
   U15598 : XOR2_X1 port map( A1 => n6526, A2 => n6525, Z => n35017);
   U15602 : NAND2_X1 port map( A1 => n1400, A2 => n482, ZN => n28823);
   U15606 : NAND2_X2 port map( A1 => n19630, A2 => n33344, ZN => n16749);
   U15613 : INV_X2 port map( I => n35021, ZN => n20212);
   U15614 : XOR2_X1 port map( A1 => n20210, A2 => n26009, Z => n35021);
   U15625 : INV_X2 port map( I => n33707, ZN => n35023);
   U15627 : OR2_X1 port map( A1 => n28598, A2 => n35023, Z => n28601);
   U15630 : NAND2_X2 port map( A1 => n35025, A2 => n35336, ZN => n15165);
   U15631 : NOR2_X2 port map( A1 => n15169, A2 => n15168, ZN => n35025);
   U15633 : OR2_X1 port map( A1 => n10220, A2 => n35462, Z => n36872);
   U15638 : XNOR2_X1 port map( A1 => n4348, A2 => n19758, ZN => n36494);
   U15640 : AOI22_X2 port map( A1 => n35026, A2 => n14373, B1 => n19403, B2 => 
                           n19768, ZN => n32292);
   U15646 : NAND2_X2 port map( A1 => n19768, A2 => n19262, ZN => n21813);
   U15650 : XOR2_X1 port map( A1 => n10185, A2 => n10183, Z => n35027);
   U15654 : INV_X2 port map( I => n28516, ZN => n9674);
   U15657 : OAI21_X2 port map( A1 => n24391, A2 => n9931, B => n9840, ZN => 
                           n24761);
   U15663 : XOR2_X1 port map( A1 => n22572, A2 => n22595, Z => n22717);
   U15665 : NOR2_X2 port map( A1 => n21829, A2 => n21828, ZN => n22572);
   U15670 : XOR2_X1 port map( A1 => n37957, A2 => n29934, Z => n23744);
   U15689 : OAI21_X2 port map( A1 => n34041, A2 => n28691, B => n33353, ZN => 
                           n2566);
   U15690 : XOR2_X1 port map( A1 => n28845, A2 => n28957, Z => n13630);
   U15697 : XOR2_X1 port map( A1 => n16776, A2 => n9977, Z => n16775);
   U15700 : XOR2_X1 port map( A1 => n8566, A2 => n34053, Z => n24009);
   U15701 : XOR2_X1 port map( A1 => n23762, A2 => n30321, Z => n8566);
   U15706 : XOR2_X1 port map( A1 => n35029, A2 => n19527, Z => Ciphertext(125))
                           ;
   U15716 : NAND2_X1 port map( A1 => n15174, A2 => n29542, ZN => n7436);
   U15717 : NAND2_X1 port map( A1 => n1497, A2 => n15996, ZN => n26670);
   U15720 : NAND2_X1 port map( A1 => n32558, A2 => n14229, ZN => n25651);
   U15740 : OAI21_X2 port map( A1 => n35031, A2 => n12987, B => n7282, ZN => 
                           n7632);
   U15743 : NAND2_X1 port map( A1 => n12986, A2 => n1002, ZN => n35031);
   U15744 : NAND2_X2 port map( A1 => n36664, A2 => n36891, ZN => n24416);
   U15752 : INV_X2 port map( I => n35032, ZN => n30494);
   U15753 : XOR2_X1 port map( A1 => n11117, A2 => n11114, Z => n35032);
   U15755 : XOR2_X1 port map( A1 => n35033, A2 => n27815, Z => n30806);
   U15756 : OAI21_X2 port map( A1 => n29899, A2 => n29898, B => n29949, ZN => 
                           n36843);
   U15761 : OAI22_X2 port map( A1 => n9078, A2 => n22493, B1 => n8692, B2 => 
                           n6303, ZN => n32089);
   U15769 : NAND2_X2 port map( A1 => n36301, A2 => n24517, ZN => n25215);
   U15778 : BUF_X4 port map( I => n28036, Z => n36979);
   U15788 : OAI22_X2 port map( A1 => n35733, A2 => n27996, B1 => n28002, B2 => 
                           n28001, ZN => n3900);
   U15790 : NAND2_X1 port map( A1 => n15232, A2 => n35034, ZN => n4730);
   U15794 : NAND3_X1 port map( A1 => n32317, A2 => n29534, A3 => n18384, ZN => 
                           n35034);
   U15795 : OR2_X1 port map( A1 => n29927, A2 => n29929, Z => n7457);
   U15796 : AOI21_X2 port map( A1 => n8666, A2 => n14600, B => n31356, ZN => 
                           n29927);
   U15802 : XOR2_X1 port map( A1 => n27605, A2 => n35035, Z => n10256);
   U15804 : XOR2_X1 port map( A1 => n557, A2 => n32160, Z => n35035);
   U15820 : NAND2_X1 port map( A1 => n27304, A2 => n31955, ZN => n35749);
   U15825 : BUF_X2 port map( I => n23532, Z => n35039);
   U15828 : BUF_X2 port map( I => n1145, Z => n35040);
   U15830 : NOR3_X1 port map( A1 => n916, A2 => n14423, A3 => n19873, ZN => 
                           n12377);
   U15841 : OAI21_X2 port map( A1 => n7691, A2 => n15512, B => n36112, ZN => 
                           n16968);
   U15855 : NAND2_X2 port map( A1 => n21804, A2 => n36735, ZN => n35042);
   U15874 : XOR2_X1 port map( A1 => n7786, A2 => n7785, Z => n18574);
   U15877 : NAND2_X1 port map( A1 => n36003, A2 => n232, ZN => n35670);
   U15879 : NAND2_X2 port map( A1 => n8332, A2 => n8331, ZN => n35051);
   U15883 : OR2_X1 port map( A1 => n10803, A2 => n29220, Z => n12978);
   U15888 : NOR2_X2 port map( A1 => n25361, A2 => n10686, ZN => n25248);
   U15893 : XOR2_X1 port map( A1 => n33372, A2 => n31720, Z => n17597);
   U15901 : XOR2_X1 port map( A1 => n7530, A2 => n17195, Z => n17987);
   U15906 : OAI21_X2 port map( A1 => n12815, A2 => n12813, B => n12812, ZN => 
                           n17195);
   U15907 : OAI21_X2 port map( A1 => n19409, A2 => n28746, B => n19408, ZN => 
                           n35222);
   U15908 : NAND2_X2 port map( A1 => n34244, A2 => n2147, ZN => n18202);
   U15920 : OAI21_X2 port map( A1 => n35863, A2 => n35045, B => n1316, ZN => 
                           n2796);
   U15921 : NOR2_X1 port map( A1 => n9975, A2 => n20590, ZN => n35045);
   U15927 : AOI22_X2 port map( A1 => n35046, A2 => n35944, B1 => n9882, B2 => 
                           n1934, ZN => n35821);
   U15928 : INV_X2 port map( I => n35047, ZN => n22723);
   U15929 : XOR2_X1 port map( A1 => n22599, A2 => n19819, Z => n35047);
   U15943 : INV_X2 port map( I => n35137, ZN => n35049);
   U15945 : XOR2_X1 port map( A1 => n26598, A2 => n26325, Z => n35656);
   U15949 : XOR2_X1 port map( A1 => n27690, A2 => n33866, Z => n33498);
   U15952 : AND2_X1 port map( A1 => n34717, A2 => n6445, Z => n3515);
   U15972 : INV_X2 port map( I => n22263, ZN => n35526);
   U15975 : NAND3_X1 port map( A1 => n35055, A2 => n1595, A3 => n35054, ZN => 
                           n20250);
   U15980 : NAND2_X1 port map( A1 => n5985, A2 => n1276, ZN => n35054);
   U15984 : INV_X1 port map( I => n20068, ZN => n35055);
   U15994 : NAND2_X2 port map( A1 => n19630, A2 => n24635, ZN => n11711);
   U15997 : NAND2_X2 port map( A1 => n35056, A2 => n11577, ZN => n11710);
   U16000 : AND2_X1 port map( A1 => n28199, A2 => n18061, Z => n35733);
   U16001 : NOR3_X2 port map( A1 => n26014, A2 => n26013, A3 => n33474, ZN => 
                           n20852);
   U16012 : XOR2_X1 port map( A1 => n11899, A2 => n25311, Z => n6233);
   U16013 : XOR2_X1 port map( A1 => n25186, A2 => n19156, Z => n25311);
   U16029 : NOR2_X1 port map( A1 => n27894, A2 => n36253, ZN => n35061);
   U16031 : AOI22_X2 port map( A1 => n14398, A2 => n36663, B1 => n36076, B2 => 
                           n14489, ZN => n6809);
   U16035 : NAND2_X2 port map( A1 => n27180, A2 => n33773, ZN => n31459);
   U16036 : OAI21_X2 port map( A1 => n10699, A2 => n8569, B => n10697, ZN => 
                           n23550);
   U16040 : NOR2_X2 port map( A1 => n24647, A2 => n18569, ZN => n24935);
   U16044 : XOR2_X1 port map( A1 => n35064, A2 => n18432, Z => Ciphertext(127))
                           ;
   U16045 : OAI22_X1 port map( A1 => n29914, A2 => n29931, B1 => n29913, B2 => 
                           n19097, ZN => n35064);
   U16058 : XOR2_X1 port map( A1 => n21087, A2 => n27844, Z => n20140);
   U16061 : XOR2_X1 port map( A1 => n27460, A2 => n1214, Z => n27844);
   U16064 : OAI22_X2 port map( A1 => n2300, A2 => n21845, B1 => n21349, B2 => 
                           n21667, ZN => n37041);
   U16066 : NAND2_X2 port map( A1 => n19517, A2 => n31222, ZN => n2300);
   U16083 : XOR2_X1 port map( A1 => n9028, A2 => n6475, Z => n23080);
   U16085 : XOR2_X1 port map( A1 => n6474, A2 => n6473, Z => n6475);
   U16090 : OR2_X1 port map( A1 => n9649, A2 => n10679, Z => n29954);
   U16102 : NAND2_X2 port map( A1 => n1688, A2 => n22222, ZN => n22224);
   U16103 : NAND2_X2 port map( A1 => n37105, A2 => n3510, ZN => n25052);
   U16106 : XOR2_X1 port map( A1 => n16254, A2 => n13254, Z => n35070);
   U16108 : INV_X2 port map( I => n35072, ZN => n31278);
   U16109 : XOR2_X1 port map( A1 => n3167, A2 => n3166, Z => n35072);
   U16112 : INV_X1 port map( I => n114, ZN => n15337);
   U16118 : NAND2_X1 port map( A1 => n35073, A2 => n114, ZN => n15761);
   U16119 : XOR2_X1 port map( A1 => Plaintext(90), A2 => Key(90), Z => n114);
   U16122 : NOR2_X1 port map( A1 => n32971, A2 => n34458, ZN => n35281);
   U16124 : NAND2_X1 port map( A1 => n38973, A2 => n35281, ZN => n35280);
   U16140 : NAND4_X2 port map( A1 => n18563, A2 => n10969, A3 => n17688, A4 => 
                           n18564, ZN => n20987);
   U16150 : XOR2_X1 port map( A1 => n5866, A2 => n23396, Z => n35076);
   U16151 : INV_X2 port map( I => n35077, ZN => n4048);
   U16154 : XOR2_X1 port map( A1 => n35079, A2 => n35078, Z => n32856);
   U16156 : XOR2_X1 port map( A1 => n11192, A2 => n22606, Z => n35079);
   U16166 : OAI22_X1 port map( A1 => n36976, A2 => n36977, B1 => n10428, B2 => 
                           n14421, ZN => n29217);
   U16167 : INV_X2 port map( I => n35080, ZN => n783);
   U16173 : NAND2_X2 port map( A1 => n31959, A2 => n18311, ZN => n27399);
   U16175 : INV_X1 port map( I => n4761, ZN => n35394);
   U16178 : XOR2_X1 port map( A1 => n22604, A2 => n1161, Z => n35081);
   U16179 : NOR2_X2 port map( A1 => n35082, A2 => n12545, ZN => n29253);
   U16192 : XOR2_X1 port map( A1 => n8533, A2 => n8530, Z => n31976);
   U16193 : XOR2_X1 port map( A1 => n35084, A2 => n35511, Z => n35842);
   U16194 : XOR2_X1 port map( A1 => n25224, A2 => n16674, Z => n35084);
   U16195 : XOR2_X1 port map( A1 => n4461, A2 => n35085, Z => n33023);
   U16196 : XOR2_X1 port map( A1 => n14171, A2 => n19126, Z => n35085);
   U16198 : NAND2_X2 port map( A1 => n601, A2 => n27507, ZN => n36639);
   U16207 : NAND2_X1 port map( A1 => n9682, A2 => n17645, ZN => n13756);
   U16220 : NOR2_X1 port map( A1 => n36304, A2 => n9954, ZN => n6005);
   U16224 : OR2_X2 port map( A1 => n20830, A2 => n20726, Z => n13261);
   U16227 : XOR2_X1 port map( A1 => n1859, A2 => n14218, Z => n35908);
   U16234 : XOR2_X1 port map( A1 => n35087, A2 => n34022, Z => n13352);
   U16236 : XOR2_X1 port map( A1 => n13354, A2 => n22653, Z => n35087);
   U16247 : OR2_X1 port map( A1 => n24558, A2 => n35088, Z => n10774);
   U16249 : XOR2_X1 port map( A1 => n25032, A2 => n5026, Z => n3187);
   U16250 : XOR2_X1 port map( A1 => n25197, A2 => n25149, Z => n5026);
   U16254 : AOI22_X2 port map( A1 => n4713, A2 => n1145, B1 => n4682, B2 => 
                           n15045, ZN => n22969);
   U16261 : NOR2_X2 port map( A1 => n7429, A2 => n5424, ZN => n20621);
   U16266 : NAND2_X2 port map( A1 => n35092, A2 => n18702, ZN => n6263);
   U16268 : NAND2_X2 port map( A1 => n35093, A2 => n11893, ZN => n33100);
   U16274 : OAI21_X2 port map( A1 => n28126, A2 => n27482, B => n11895, ZN => 
                           n35093);
   U16277 : XOR2_X1 port map( A1 => n3887, A2 => n3890, Z => n21159);
   U16288 : AOI22_X1 port map( A1 => n5821, A2 => n9422, B1 => n33168, B2 => 
                           n1339, ZN => n7105);
   U16289 : NOR2_X2 port map( A1 => n37041, A2 => n8073, ZN => n33168);
   U16292 : NAND2_X2 port map( A1 => n30174, A2 => n10101, ZN => n20342);
   U16295 : NAND2_X2 port map( A1 => n35096, A2 => n4799, ZN => n30093);
   U16303 : XOR2_X1 port map( A1 => n29819, A2 => n28817, Z => n29245);
   U16316 : NOR2_X2 port map( A1 => n22128, A2 => n4424, ZN => n18566);
   U16332 : XOR2_X1 port map( A1 => n12575, A2 => n35097, Z => n4866);
   U16334 : XOR2_X1 port map( A1 => n12574, A2 => n32306, Z => n35097);
   U16345 : AOI22_X2 port map( A1 => n31781, A2 => n42, B1 => n8369, B2 => 
                           n1444, ZN => n8366);
   U16346 : XOR2_X1 port map( A1 => n23725, A2 => n1993, Z => n33559);
   U16351 : AOI21_X1 port map( A1 => n38155, A2 => n6287, B => n13379, ZN => 
                           n10272);
   U16372 : OAI22_X1 port map( A1 => n29735, A2 => n29728, B1 => n38143, B2 => 
                           n29750, ZN => n29729);
   U16388 : NOR2_X2 port map( A1 => n36071, A2 => n18786, ZN => n2626);
   U16414 : NOR2_X1 port map( A1 => n2035, A2 => n39296, ZN => n27486);
   U16419 : XOR2_X1 port map( A1 => n36867, A2 => n22644, Z => n16254);
   U16428 : OAI21_X2 port map( A1 => n2060, A2 => n28356, B => n11129, ZN => 
                           n28817);
   U16429 : BUF_X4 port map( I => n26177, Z => n26700);
   U16430 : AOI21_X2 port map( A1 => n1514, A2 => n9175, B => n35102, ZN => 
                           n3519);
   U16431 : INV_X2 port map( I => n26114, ZN => n35102);
   U16441 : XOR2_X1 port map( A1 => n27730, A2 => n27525, Z => n12507);
   U16443 : XOR2_X1 port map( A1 => n29128, A2 => n29126, Z => n21077);
   U16451 : XOR2_X1 port map( A1 => n26523, A2 => n2195, Z => n35105);
   U16455 : NAND2_X1 port map( A1 => n14739, A2 => n37088, ZN => n14742);
   U16460 : NAND3_X2 port map( A1 => n23069, A2 => n6000, A3 => n11366, ZN => 
                           n31594);
   U16466 : XOR2_X1 port map( A1 => n26565, A2 => n29476, Z => n26198);
   U16468 : NAND2_X2 port map( A1 => n33423, A2 => n21198, ZN => n26565);
   U16472 : NAND2_X2 port map( A1 => n20168, A2 => n16581, ZN => n25242);
   U16474 : NAND2_X2 port map( A1 => n24751, A2 => n24750, ZN => n20168);
   U16477 : NAND2_X2 port map( A1 => n37099, A2 => n29491, ZN => n20209);
   U16480 : NAND2_X2 port map( A1 => n35108, A2 => n24199, ZN => n24719);
   U16481 : NAND3_X2 port map( A1 => n37065, A2 => n32491, A3 => n32492, ZN => 
                           n35108);
   U16490 : XOR2_X1 port map( A1 => n19014, A2 => n14610, Z => n31849);
   U16491 : INV_X4 port map( I => n32885, ZN => n1323);
   U16492 : NAND2_X2 port map( A1 => n5063, A2 => n5768, ZN => n24704);
   U16496 : XOR2_X1 port map( A1 => n28840, A2 => n29146, Z => n36545);
   U16501 : OR2_X1 port map( A1 => n9520, A2 => n23907, Z => n10342);
   U16511 : OAI21_X2 port map( A1 => n33725, A2 => n879, B => n37623, ZN => 
                           n6264);
   U16529 : BUF_X4 port map( I => n15933, Z => n12771);
   U16533 : INV_X1 port map( I => n25851, ZN => n36896);
   U16534 : XNOR2_X1 port map( A1 => n9757, A2 => n15401, ZN => n140);
   U16540 : XOR2_X1 port map( A1 => n23777, A2 => n34054, Z => n32610);
   U16545 : BUF_X2 port map( I => n6893, Z => n35112);
   U16547 : NAND3_X2 port map( A1 => n30584, A2 => n7227, A3 => n35113, ZN => 
                           n32404);
   U16560 : INV_X2 port map( I => n1218, ZN => n35114);
   U16570 : NOR2_X2 port map( A1 => n22100, A2 => n9736, ZN => n22176);
   U16584 : NAND3_X1 port map( A1 => n1477, A2 => n997, A3 => n8537, ZN => 
                           n27158);
   U16605 : XOR2_X1 port map( A1 => n25249, A2 => n25299, Z => n11519);
   U16606 : AND2_X1 port map( A1 => n24425, A2 => n14371, Z => n5254);
   U16612 : NAND2_X2 port map( A1 => n14371, A2 => n10073, ZN => n24425);
   U16621 : XOR2_X1 port map( A1 => n34092, A2 => n35120, Z => n36104);
   U16634 : XOR2_X1 port map( A1 => n25156, A2 => n5829, Z => n35120);
   U16635 : INV_X4 port map( I => n18028, ZN => n12927);
   U16636 : OAI21_X2 port map( A1 => n17098, A2 => n17099, B => n35121, ZN => 
                           n11020);
   U16638 : AOI22_X2 port map( A1 => n14830, A2 => n26978, B1 => n14831, B2 => 
                           n33301, ZN => n35121);
   U16644 : NAND2_X1 port map( A1 => n8042, A2 => n10008, ZN => n35122);
   U16653 : NOR2_X1 port map( A1 => n978, A2 => n33100, ZN => n30917);
   U16655 : NOR3_X1 port map( A1 => n35979, A2 => n12377, A3 => n22388, ZN => 
                           n36349);
   U16657 : AOI21_X2 port map( A1 => n2028, A2 => n35822, B => n35194, ZN => 
                           n35193);
   U16660 : NAND2_X2 port map( A1 => n12669, A2 => n8228, ZN => n33437);
   U16673 : NOR2_X2 port map( A1 => n21318, A2 => n19748, ZN => n35124);
   U16695 : XOR2_X1 port map( A1 => n36497, A2 => n2119, Z => n36231);
   U16717 : NAND2_X1 port map( A1 => n9211, A2 => n9213, ZN => n36322);
   U16724 : AOI22_X2 port map( A1 => n22950, A2 => n39752, B1 => n22951, B2 => 
                           n23020, ZN => n22952);
   U16729 : NOR2_X1 port map( A1 => n21609, A2 => n21610, ZN => n36297);
   U16730 : NOR2_X2 port map( A1 => n31437, A2 => n34031, ZN => n35686);
   U16734 : XOR2_X1 port map( A1 => n13917, A2 => n25211, Z => n25039);
   U16740 : AOI21_X1 port map( A1 => n22366, A2 => n22227, B => n20623, ZN => 
                           n21104);
   U16748 : NAND2_X2 port map( A1 => n20643, A2 => n20646, ZN => n22227);
   U16789 : INV_X2 port map( I => n38669, ZN => n36777);
   U16792 : XOR2_X1 port map( A1 => n22462, A2 => n6325, Z => n7931);
   U16793 : XOR2_X1 port map( A1 => n22582, A2 => n18778, Z => n22462);
   U16800 : INV_X1 port map( I => n479, ZN => n27433);
   U16803 : NOR3_X1 port map( A1 => n29433, A2 => n14414, A3 => n18502, ZN => 
                           n29436);
   U16809 : NAND2_X2 port map( A1 => n28569, A2 => n33995, ZN => n28448);
   U16813 : INV_X2 port map( I => n22586, ZN => n1668);
   U16835 : NOR2_X1 port map( A1 => n1313, A2 => n8942, ZN => n10867);
   U16841 : INV_X2 port map( I => n5732, ZN => n8942);
   U16843 : OR2_X1 port map( A1 => n21445, A2 => n21669, Z => n31292);
   U16858 : BUF_X4 port map( I => n19979, Z => n36082);
   U16868 : NAND3_X1 port map( A1 => n30071, A2 => n30076, A3 => n4377, ZN => 
                           n30073);
   U16874 : OAI22_X1 port map( A1 => n22840, A2 => n13042, B1 => n23106, B2 => 
                           n23104, ZN => n22841);
   U16882 : XOR2_X1 port map( A1 => n22391, A2 => n22656, Z => n22457);
   U16887 : XOR2_X1 port map( A1 => n18300, A2 => n8951, Z => n15648);
   U16892 : XOR2_X1 port map( A1 => n17775, A2 => n35139, Z => n33676);
   U16894 : XOR2_X1 port map( A1 => n9979, A2 => n35140, Z => n35139);
   U16902 : NAND2_X1 port map( A1 => n29547, A2 => n35141, ZN => n21069);
   U16907 : INV_X2 port map( I => n19097, ZN => n29932);
   U16908 : XOR2_X1 port map( A1 => n11927, A2 => n11925, Z => n15738);
   U16917 : INV_X2 port map( I => n35143, ZN => n30853);
   U16921 : XOR2_X1 port map( A1 => n29077, A2 => n20622, Z => n29381);
   U16929 : NAND3_X2 port map( A1 => n35144, A2 => n5294, A3 => n5295, ZN => 
                           n36894);
   U16940 : NAND2_X1 port map( A1 => n14127, A2 => n3693, ZN => n35547);
   U16942 : OAI21_X2 port map( A1 => n9292, A2 => n9293, B => n25630, ZN => 
                           n35145);
   U16946 : AOI21_X2 port map( A1 => n35146, A2 => n5509, B => n14642, ZN => 
                           n5705);
   U16953 : NAND2_X2 port map( A1 => n584, A2 => n33860, ZN => n16281);
   U16958 : OAI21_X2 port map( A1 => n17077, A2 => n28311, B => n15211, ZN => 
                           n8911);
   U16970 : XOR2_X1 port map( A1 => n18942, A2 => n35147, Z => n35868);
   U16971 : XOR2_X1 port map( A1 => n35760, A2 => n35148, Z => n35147);
   U16977 : INV_X2 port map( I => n35149, ZN => n21137);
   U16978 : XNOR2_X1 port map( A1 => n18578, A2 => n18580, ZN => n35149);
   U16981 : AOI22_X2 port map( A1 => n19146, A2 => n23321, B1 => n16047, B2 => 
                           n961, ZN => n18485);
   U16983 : XOR2_X1 port map( A1 => n7766, A2 => n28989, Z => n20819);
   U16984 : XOR2_X1 port map( A1 => n12741, A2 => n8939, Z => n28989);
   U16986 : AND2_X1 port map( A1 => n19667, A2 => n34370, Z => n31913);
   U16993 : AOI21_X1 port map( A1 => n33416, A2 => n29735, B => n29733, ZN => 
                           n29736);
   U17003 : NAND2_X2 port map( A1 => n29486, A2 => n14417, ZN => n29444);
   U17019 : NAND2_X2 port map( A1 => n11952, A2 => n35155, ZN => n18289);
   U17031 : AOI21_X1 port map( A1 => n37050, A2 => n955, B => n32105, ZN => 
                           n35156);
   U17036 : XNOR2_X1 port map( A1 => n29073, A2 => n18430, ZN => n9994);
   U17041 : XNOR2_X1 port map( A1 => n15595, A2 => n26397, ZN => n36468);
   U17045 : NAND2_X1 port map( A1 => n25883, A2 => n8006, ZN => n35159);
   U17059 : XOR2_X1 port map( A1 => n208, A2 => n23777, Z => n5510);
   U17061 : BUF_X2 port map( I => n25427, Z => n35160);
   U17063 : XOR2_X1 port map( A1 => n27617, A2 => n27594, Z => n35708);
   U17065 : NAND3_X2 port map( A1 => n26846, A2 => n26844, A3 => n26845, ZN => 
                           n27594);
   U17066 : INV_X2 port map( I => n35161, ZN => n8293);
   U17072 : XOR2_X1 port map( A1 => n35162, A2 => n35389, Z => n32049);
   U17073 : XOR2_X1 port map( A1 => n17349, A2 => n38174, Z => n35162);
   U17076 : XOR2_X1 port map( A1 => n3550, A2 => n3548, Z => n9393);
   U17080 : XOR2_X1 port map( A1 => n21030, A2 => n5116, Z => n35163);
   U17083 : XOR2_X1 port map( A1 => n7582, A2 => n34052, Z => n32432);
   U17105 : OAI21_X2 port map( A1 => n39829, A2 => n35165, B => n28789, ZN => 
                           n30131);
   U17112 : NOR2_X1 port map( A1 => n28788, A2 => n38196, ZN => n35165);
   U17118 : XOR2_X1 port map( A1 => n8958, A2 => n35421, Z => n9470);
   U17121 : XOR2_X1 port map( A1 => n29086, A2 => n35168, Z => n31867);
   U17123 : XOR2_X1 port map( A1 => n8939, A2 => n35169, Z => n35168);
   U17125 : INV_X1 port map( I => n29476, ZN => n35169);
   U17126 : XOR2_X1 port map( A1 => n36869, A2 => n6328, Z => n36932);
   U17131 : AOI21_X1 port map( A1 => n12189, A2 => n6648, B => n35287, ZN => 
                           n13721);
   U17144 : OAI22_X2 port map( A1 => n17475, A2 => n39537, B1 => n20154, B2 => 
                           n35170, ZN => n17474);
   U17147 : XOR2_X1 port map( A1 => n25210, A2 => n25174, Z => n5315);
   U17157 : AOI21_X2 port map( A1 => n9997, A2 => n6337, B => n24600, ZN => 
                           n24128);
   U17158 : NOR3_X2 port map( A1 => n11710, A2 => n3120, A3 => n15332, ZN => 
                           n3124);
   U17159 : INV_X4 port map( I => n29862, ZN => n29956);
   U17164 : OR2_X1 port map( A1 => n35217, A2 => n37060, Z => n19088);
   U17165 : INV_X2 port map( I => n27571, ZN => n35417);
   U17168 : INV_X2 port map( I => n28961, ZN => n29761);
   U17173 : NOR2_X2 port map( A1 => n4322, A2 => n36546, ZN => n25743);
   U17176 : NAND2_X2 port map( A1 => n30260, A2 => n30257, ZN => n30250);
   U17181 : OR2_X2 port map( A1 => n11428, A2 => n39827, Z => n11125);
   U17188 : INV_X2 port map( I => n482, ZN => n30165);
   U17189 : NAND2_X1 port map( A1 => n24235, A2 => n30311, ZN => n8160);
   U17201 : NAND2_X2 port map( A1 => n18873, A2 => n9105, ZN => n20964);
   U17204 : NAND2_X2 port map( A1 => n36859, A2 => n33316, ZN => n13010);
   U17207 : NOR2_X1 port map( A1 => n31587, A2 => n12931, ZN => n35171);
   U17210 : INV_X1 port map( I => n25699, ZN => n1110);
   U17233 : NOR2_X1 port map( A1 => n38164, A2 => n8287, ZN => n20922);
   U17236 : OAI22_X1 port map( A1 => n981, A2 => n1207, B1 => n5469, B2 => 
                           n28290, ZN => n30872);
   U17242 : AOI22_X1 port map( A1 => n29605, A2 => n29604, B1 => n29625, B2 => 
                           n29611, ZN => n30657);
   U17245 : NAND2_X1 port map( A1 => n18306, A2 => n36382, ZN => n29625);
   U17247 : NAND3_X1 port map( A1 => n76, A2 => n17532, A3 => n2877, ZN => 
                           n2666);
   U17252 : NOR2_X2 port map( A1 => n36029, A2 => n10393, ZN => n35173);
   U17263 : OR2_X1 port map( A1 => n13442, A2 => n17262, Z => n19173);
   U17283 : CLKBUF_X12 port map( I => n20512, Z => n31022);
   U17285 : NAND2_X1 port map( A1 => n31022, A2 => n6640, ZN => n2050);
   U17291 : NAND2_X1 port map( A1 => n9141, A2 => n28717, ZN => n11009);
   U17295 : INV_X1 port map( I => n20454, ZN => n20659);
   U17301 : NOR2_X1 port map( A1 => n28490, A2 => n18960, ZN => n12544);
   U17304 : NAND3_X1 port map( A1 => n28490, A2 => n18960, A3 => n4950, ZN => 
                           n28452);
   U17307 : NOR2_X1 port map( A1 => n32781, A2 => n18626, ZN => n18625);
   U17320 : AOI22_X1 port map( A1 => n29688, A2 => n5067, B1 => n29685, B2 => 
                           n29686, ZN => n31914);
   U17321 : INV_X1 port map( I => n18837, ZN => n36767);
   U17323 : INV_X2 port map( I => n23307, ZN => n22493);
   U17324 : NAND3_X1 port map( A1 => n29392, A2 => n29393, A3 => n29391, ZN => 
                           n35676);
   U17338 : NAND2_X1 port map( A1 => n29232, A2 => n35185, ZN => n36232);
   U17339 : NOR2_X1 port map( A1 => n5955, A2 => n7834, ZN => n5954);
   U17351 : OAI21_X1 port map( A1 => n10763, A2 => n13752, B => n11453, ZN => 
                           n35811);
   U17355 : OR2_X1 port map( A1 => n28585, A2 => n28584, Z => n35179);
   U17364 : NAND2_X1 port map( A1 => n30035, A2 => n8039, ZN => n18783);
   U17367 : OAI21_X1 port map( A1 => n20102, A2 => n37021, B => n30059, ZN => 
                           n36268);
   U17381 : AOI22_X1 port map( A1 => n20922, A2 => n17192, B1 => n30129, B2 => 
                           n38164, ZN => n20921);
   U17392 : NOR2_X1 port map( A1 => n36964, A2 => n10708, ZN => n24036);
   U17393 : AOI21_X2 port map( A1 => n10711, A2 => n9011, B => n36965, ZN => 
                           n36964);
   U17397 : BUF_X2 port map( I => n26651, Z => n4138);
   U17400 : NAND2_X1 port map( A1 => n33203, A2 => n30986, ZN => n31764);
   U17401 : INV_X2 port map( I => n29699, ZN => n1182);
   U17405 : NAND2_X1 port map( A1 => n38163, A2 => n20274, ZN => n29007);
   U17407 : NAND2_X1 port map( A1 => n1193, A2 => n28311, ZN => n15211);
   U17417 : NOR2_X1 port map( A1 => n28749, A2 => n28746, ZN => n33106);
   U17418 : NAND2_X1 port map( A1 => n4024, A2 => n28746, ZN => n4023);
   U17438 : NAND2_X1 port map( A1 => n9200, A2 => n38227, ZN => n7797);
   U17446 : NOR2_X1 port map( A1 => n28823, A2 => n30160, ZN => n35183);
   U17448 : AND2_X1 port map( A1 => n29979, A2 => n18896, Z => n33422);
   U17456 : AOI22_X1 port map( A1 => n1442, A2 => n14263, B1 => n1072, B2 => 
                           n28105, ZN => n13249);
   U17475 : INV_X1 port map( I => n27249, ZN => n19918);
   U17479 : AOI22_X1 port map( A1 => n27027, A2 => n13213, B1 => n13212, B2 => 
                           n27247, ZN => n13211);
   U17482 : AOI21_X1 port map( A1 => n8651, A2 => n26961, B => n8556, ZN => 
                           n7607);
   U17488 : INV_X1 port map( I => n29137, ZN => n36668);
   U17500 : AND2_X2 port map( A1 => n9173, A2 => n35673, Z => n35186);
   U17503 : NOR2_X1 port map( A1 => n5825, A2 => n1379, ZN => n36677);
   U17506 : NAND2_X1 port map( A1 => n33963, A2 => n6938, ZN => n30222);
   U17514 : NOR2_X1 port map( A1 => n29310, A2 => n12876, ZN => n12878);
   U17546 : NAND2_X1 port map( A1 => n23159, A2 => n22935, ZN => n18865);
   U17561 : AND2_X1 port map( A1 => n18042, A2 => n29684, Z => n18041);
   U17567 : NOR2_X1 port map( A1 => n29747, A2 => n29740, ZN => n29728);
   U17568 : NAND2_X1 port map( A1 => n16889, A2 => n14858, ZN => n36051);
   U17574 : NOR2_X1 port map( A1 => n20184, A2 => n28143, ZN => n20185);
   U17582 : NAND2_X1 port map( A1 => n28375, A2 => n29635, ZN => n36125);
   U17583 : INV_X1 port map( I => n30141, ZN => n30136);
   U17586 : NOR2_X1 port map( A1 => n28131, A2 => n28229, ZN => n35819);
   U17588 : INV_X1 port map( I => n19891, ZN => n35659);
   U17591 : NAND2_X1 port map( A1 => n8592, A2 => n30047, ZN => n8591);
   U17609 : XNOR2_X1 port map( A1 => n26537, A2 => n26488, ZN => n36077);
   U17611 : INV_X2 port map( I => n10803, ZN => n32209);
   U17613 : INV_X2 port map( I => n18240, ZN => n10803);
   U17619 : NAND2_X2 port map( A1 => n53, A2 => n9739, ZN => n35188);
   U17625 : NOR2_X1 port map( A1 => n28224, A2 => n2868, ZN => n35820);
   U17626 : OR2_X2 port map( A1 => n33262, A2 => n33261, Z => n35189);
   U17631 : OR2_X2 port map( A1 => n33262, A2 => n33261, Z => n35190);
   U17633 : INV_X1 port map( I => n17220, ZN => n36260);
   U17639 : NOR2_X1 port map( A1 => n3003, A2 => n22228, ZN => n22089);
   U17641 : AOI22_X1 port map( A1 => n10868, A2 => n29579, B1 => n10869, B2 => 
                           n29580, ZN => n29619);
   U17644 : INV_X1 port map( I => n29815, ZN => n13574);
   U17655 : INV_X2 port map( I => n4377, ZN => n30078);
   U17678 : NAND2_X1 port map( A1 => n15703, A2 => n26090, ZN => n10511);
   U17696 : INV_X2 port map( I => n25601, ZN => n1254);
   U17698 : INV_X1 port map( I => n26651, ZN => n31254);
   U17708 : NAND2_X1 port map( A1 => n11866, A2 => n35622, ZN => n32142);
   U17712 : NAND2_X2 port map( A1 => n8138, A2 => n32506, ZN => n35196);
   U17717 : NOR2_X1 port map( A1 => n9242, A2 => n35469, ZN => n7839);
   U17720 : NAND3_X1 port map( A1 => n7535, A2 => n7534, A3 => n1302, ZN => 
                           n12269);
   U17732 : OAI21_X1 port map( A1 => n31107, A2 => n11283, B => n7690, ZN => 
                           n35862);
   U17749 : INV_X1 port map( I => n26246, ZN => n10776);
   U17750 : XNOR2_X1 port map( A1 => n28830, A2 => n35320, ZN => n28545);
   U17759 : INV_X2 port map( I => n20156, ZN => n14278);
   U17760 : NAND2_X1 port map( A1 => n4192, A2 => n32046, ZN => n2429);
   U17770 : AND2_X1 port map( A1 => n30173, A2 => n30172, Z => n35254);
   U17778 : INV_X1 port map( I => n1403, ZN => n36269);
   U17780 : NAND2_X1 port map( A1 => n28720, A2 => n28722, ZN => n4980);
   U17784 : NAND3_X1 port map( A1 => n38073, A2 => n7044, A3 => n34011, ZN => 
                           n18460);
   U17786 : OAI21_X1 port map( A1 => n38073, A2 => n37983, B => n32882, ZN => 
                           n17862);
   U17787 : NAND2_X1 port map( A1 => n38073, A2 => n34011, ZN => n17857);
   U17788 : NAND2_X1 port map( A1 => n31328, A2 => n24784, ZN => n24506);
   U17792 : NOR2_X1 port map( A1 => n24784, A2 => n24874, ZN => n24643);
   U17794 : NAND2_X1 port map( A1 => n24784, A2 => n31519, ZN => n31023);
   U17803 : NAND3_X1 port map( A1 => n30822, A2 => n16676, A3 => n20342, ZN => 
                           n11264);
   U17808 : NAND3_X1 port map( A1 => n11264, A2 => n11263, A3 => n30168, ZN => 
                           n30971);
   U17809 : AND3_X1 port map( A1 => n27338, A2 => n27053, A3 => n27341, Z => 
                           n14692);
   U17810 : NOR2_X1 port map( A1 => n20578, A2 => n14601, ZN => n17466);
   U17845 : NAND2_X1 port map( A1 => n28559, A2 => n15792, ZN => n28561);
   U17850 : XNOR2_X1 port map( A1 => n31215, A2 => n14802, ZN => n35197);
   U17851 : AOI21_X1 port map( A1 => n11421, A2 => n34484, B => n35988, ZN => 
                           n35198);
   U17854 : NOR2_X1 port map( A1 => n27441, A2 => n27440, ZN => n160);
   U17865 : INV_X1 port map( I => n28130, ZN => n28228);
   U17867 : NAND2_X1 port map( A1 => n30780, A2 => n36266, ZN => n35199);
   U17869 : NAND2_X1 port map( A1 => n1068, A2 => n28677, ZN => n28675);
   U17877 : OAI21_X2 port map( A1 => n18464, A2 => n14504, B => n18463, ZN => 
                           n35200);
   U17880 : INV_X1 port map( I => n33946, ZN => n32291);
   U17898 : NOR2_X1 port map( A1 => n910, A2 => n2678, ZN => n33032);
   U17904 : NOR2_X1 port map( A1 => n1100, A2 => n34265, ZN => n14650);
   U17911 : NOR2_X1 port map( A1 => n25688, A2 => n25587, ZN => n36412);
   U17913 : NAND2_X1 port map( A1 => n4603, A2 => n25587, ZN => n36592);
   U17919 : CLKBUF_X12 port map( I => n27903, Z => n19743);
   U17924 : NAND2_X1 port map( A1 => n33254, A2 => n27284, ZN => n35905);
   U17925 : OR2_X2 port map( A1 => n7500, A2 => n8128, Z => n16234);
   U17926 : OAI21_X2 port map( A1 => n24968, A2 => n24967, B => n19574, ZN => 
                           n35202);
   U17931 : OAI21_X1 port map( A1 => n29762, A2 => n19568, B => n29764, ZN => 
                           n29637);
   U17939 : CLKBUF_X4 port map( I => n29044, Z => n30964);
   U17940 : INV_X1 port map( I => n3827, ZN => n14412);
   U17965 : OAI21_X1 port map( A1 => n31022, A2 => n20531, B => n200, ZN => 
                           n31001);
   U17970 : NAND2_X1 port map( A1 => n14931, A2 => n89, ZN => n35583);
   U17986 : NAND2_X1 port map( A1 => n12288, A2 => n24158, ZN => n12287);
   U17998 : NAND2_X1 port map( A1 => n25978, A2 => n26031, ZN => n16477);
   U18008 : NAND2_X2 port map( A1 => n3248, A2 => n3250, ZN => n35208);
   U18012 : AOI21_X1 port map( A1 => n2629, A2 => n8393, B => n1742, ZN => 
                           n26275);
   U18016 : INV_X1 port map( I => n28591, ZN => n28674);
   U18017 : XNOR2_X1 port map( A1 => n33962, A2 => n16787, ZN => n35210);
   U18018 : AOI21_X1 port map( A1 => n30055, A2 => n34179, B => n9918, ZN => 
                           n10671);
   U18022 : BUF_X2 port map( I => n30055, Z => n19909);
   U18023 : OAI21_X1 port map( A1 => n12450, A2 => n29486, B => n33425, ZN => 
                           n10259);
   U18029 : NAND2_X1 port map( A1 => n34006, A2 => n29642, ZN => n36100);
   U18037 : OAI21_X1 port map( A1 => n27349, A2 => n27347, B => n35767, ZN => 
                           n35766);
   U18039 : OAI22_X1 port map( A1 => n30017, A2 => n30024, B1 => n30015, B2 => 
                           n15643, ZN => n30013);
   U18043 : AOI22_X2 port map( A1 => n36092, A2 => n34128, B1 => n22060, B2 => 
                           n8618, ZN => n35211);
   U18060 : XOR2_X1 port map( A1 => n16689, A2 => n16687, Z => n35213);
   U18062 : NAND2_X1 port map( A1 => n8235, A2 => n8234, ZN => n35214);
   U18067 : AOI21_X1 port map( A1 => n18406, A2 => n25993, B => n37613, ZN => 
                           n16247);
   U18068 : OAI21_X1 port map( A1 => n23819, A2 => n24116, B => n38224, ZN => 
                           n14255);
   U18069 : AOI21_X2 port map( A1 => n1830, A2 => n23340, B => n1829, ZN => 
                           n35215);
   U18078 : AOI21_X1 port map( A1 => n1830, A2 => n23340, B => n1829, ZN => 
                           n3503);
   U18082 : NAND3_X1 port map( A1 => n17224, A2 => n19559, A3 => n21246, ZN => 
                           n20221);
   U18090 : NAND3_X1 port map( A1 => n9591, A2 => n1174, A3 => n19097, ZN => 
                           n21282);
   U18094 : NOR2_X1 port map( A1 => n20510, A2 => n30128, ZN => n35624);
   U18095 : INV_X2 port map( I => n26089, ZN => n949);
   U18096 : XOR2_X1 port map( A1 => n589, A2 => n14835, Z => n35217);
   U18099 : OR3_X2 port map( A1 => n33919, A2 => n20039, A3 => n8430, Z => 
                           n10969);
   U18109 : INV_X1 port map( I => n20039, ZN => n24787);
   U18110 : NAND2_X1 port map( A1 => n21031, A2 => n37048, ZN => n25479);
   U18115 : AOI21_X1 port map( A1 => n33474, A2 => n1098, B => n26123, ZN => 
                           n26017);
   U18127 : INV_X1 port map( I => n16371, ZN => n29263);
   U18134 : BUF_X2 port map( I => n16371, Z => n16123);
   U18146 : OR2_X2 port map( A1 => n17597, A2 => n16371, Z => n19162);
   U18147 : INV_X1 port map( I => n10371, ZN => n3932);
   U18149 : AOI21_X1 port map( A1 => n20538, A2 => n12301, B => n30176, ZN => 
                           n11263);
   U18151 : NAND2_X1 port map( A1 => n1481, A2 => n36840, ZN => n30588);
   U18153 : INV_X1 port map( I => n27700, ZN => n36566);
   U18163 : NOR2_X1 port map( A1 => n39316, A2 => n33316, ZN => n2085);
   U18167 : NAND2_X1 port map( A1 => n33316, A2 => n35331, ZN => n12212);
   U18181 : NAND2_X1 port map( A1 => n31772, A2 => n13761, ZN => n10685);
   U18183 : INV_X1 port map( I => n24700, ZN => n35219);
   U18184 : AOI21_X2 port map( A1 => n24531, A2 => n8389, B => n8388, ZN => 
                           n35220);
   U18189 : OAI22_X1 port map( A1 => n36677, A2 => n36676, B1 => n17975, B2 => 
                           n17773, ZN => n17974);
   U18196 : OR2_X1 port map( A1 => n14800, A2 => n14801, Z => n35221);
   U18204 : AND2_X2 port map( A1 => n35928, A2 => n18378, Z => n35224);
   U18210 : NOR2_X1 port map( A1 => n378, A2 => n33293, ZN => n14854);
   U18211 : NOR2_X1 port map( A1 => n19448, A2 => n21277, ZN => n20669);
   U18212 : NAND2_X1 port map( A1 => n1823, A2 => n28460, ZN => n32769);
   U18218 : XOR2_X1 port map( A1 => n8403, A2 => n8404, Z => n35225);
   U18224 : NAND2_X1 port map( A1 => n35344, A2 => n10143, ZN => n11776);
   U18225 : NAND2_X2 port map( A1 => n19329, A2 => n8210, ZN => n35229);
   U18234 : NAND2_X1 port map( A1 => n10702, A2 => n19544, ZN => n10703);
   U18236 : OAI21_X1 port map( A1 => n5453, A2 => n2799, B => n4914, ZN => 
                           n5452);
   U18237 : AOI21_X1 port map( A1 => n9161, A2 => n17353, B => n4914, ZN => 
                           n5354);
   U18239 : NAND3_X1 port map( A1 => n4914, A2 => n2799, A3 => n728, ZN => 
                           n13465);
   U18240 : NAND3_X1 port map( A1 => n954, A2 => n4914, A3 => n10104, ZN => 
                           n2958);
   U18253 : INV_X1 port map( I => n19436, ZN => n26879);
   U18255 : CLKBUF_X4 port map( I => n5351, Z => n5239);
   U18264 : INV_X1 port map( I => n23602, ZN => n35230);
   U18271 : AND2_X2 port map( A1 => n34160, A2 => n12836, Z => n2966);
   U18274 : CLKBUF_X2 port map( I => n15332, Z => n10013);
   U18295 : AND2_X2 port map( A1 => n11296, A2 => n13880, Z => n28633);
   U18314 : CLKBUF_X4 port map( I => n39489, Z => n31383);
   U18317 : NAND2_X1 port map( A1 => n25867, A2 => n26019, ZN => n25868);
   U18323 : NAND3_X1 port map( A1 => n856, A2 => n26672, A3 => n17217, ZN => 
                           n11227);
   U18328 : AOI22_X1 port map( A1 => n35274, A2 => n20357, B1 => n19778, B2 => 
                           n3833, ZN => n35231);
   U18344 : NAND2_X2 port map( A1 => n23210, A2 => n23209, ZN => n7014);
   U18347 : NOR2_X1 port map( A1 => n24309, A2 => n24446, ZN => n8681);
   U18349 : INV_X2 port map( I => n24309, ZN => n24086);
   U18358 : NOR2_X1 port map( A1 => n29739, A2 => n29756, ZN => n29752);
   U18374 : INV_X1 port map( I => n21669, ZN => n21446);
   U18384 : INV_X2 port map( I => n23929, ZN => n35235);
   U18387 : AOI21_X1 port map( A1 => n7770, A2 => n7769, B => n38674, ZN => 
                           n30854);
   U18390 : NOR2_X1 port map( A1 => n19065, A2 => n29481, ZN => n16877);
   U18391 : INV_X2 port map( I => n9945, ZN => n23819);
   U18405 : AOI21_X1 port map( A1 => n28137, A2 => n33960, B => n19667, ZN => 
                           n10266);
   U18412 : XOR2_X1 port map( A1 => n1259, A2 => n11698, Z => n35237);
   U18423 : INV_X1 port map( I => n8407, ZN => n19590);
   U18430 : NOR3_X1 port map( A1 => n25661, A2 => n25660, A3 => n25379, ZN => 
                           n25499);
   U18440 : AOI21_X1 port map( A1 => n9277, A2 => n7693, B => n17087, ZN => 
                           n11121);
   U18441 : NAND2_X1 port map( A1 => n10116, A2 => n7693, ZN => n5390);
   U18442 : CLKBUF_X2 port map( I => n7693, Z => n35373);
   U18447 : INV_X1 port map( I => n27213, ZN => n31710);
   U18455 : NOR2_X1 port map( A1 => n19580, A2 => n3213, ZN => n33558);
   U18456 : CLKBUF_X4 port map( I => n25546, Z => n19701);
   U18467 : NOR2_X1 port map( A1 => n4232, A2 => n7023, ZN => n36247);
   U18468 : NOR2_X1 port map( A1 => n17469, A2 => n31527, ZN => n36421);
   U18473 : NAND2_X1 port map( A1 => n861, A2 => n19712, ZN => n36261);
   U18476 : NOR2_X1 port map( A1 => n36716, A2 => n5063, ZN => n31893);
   U18478 : INV_X1 port map( I => n27357, ZN => n13754);
   U18484 : NOR2_X1 port map( A1 => n29534, A2 => n29531, ZN => n15233);
   U18489 : XNOR2_X1 port map( A1 => n35601, A2 => n32890, ZN => n35244);
   U18493 : AND2_X2 port map( A1 => n16445, A2 => n15933, Z => n10690);
   U18497 : INV_X1 port map( I => n29616, ZN => n36548);
   U18510 : XNOR2_X1 port map( A1 => n22736, A2 => n4346, ZN => n35247);
   U18514 : NAND2_X1 port map( A1 => n29858, A2 => n29859, ZN => n29847);
   U18521 : NAND2_X1 port map( A1 => n28312, A2 => n5418, ZN => n35479);
   U18527 : OAI22_X1 port map( A1 => n29881, A2 => n17286, B1 => n29880, B2 => 
                           n29883, ZN => n10845);
   U18531 : OR2_X1 port map( A1 => n17198, A2 => n31596, Z => n35572);
   U18533 : OAI21_X1 port map( A1 => n18384, A2 => n29535, B => n29532, ZN => 
                           n29490);
   U18538 : NOR2_X1 port map( A1 => n22316, A2 => n3863, ZN => n37011);
   U18551 : OAI21_X1 port map( A1 => n19497, A2 => n20672, B => n29683, ZN => 
                           n29685);
   U18557 : XNOR2_X1 port map( A1 => n25146, A2 => n1895, ZN => n25330);
   U18562 : NOR2_X1 port map( A1 => n25539, A2 => n25540, ZN => n25541);
   U18578 : AOI21_X1 port map( A1 => n30786, A2 => n28311, B => n30785, ZN => 
                           n18931);
   U18581 : AOI21_X1 port map( A1 => n841, A2 => n14460, B => n18164, ZN => 
                           n32867);
   U18588 : INV_X1 port map( I => n20536, ZN => n36372);
   U18595 : INV_X1 port map( I => n22639, ZN => n3203);
   U18600 : INV_X1 port map( I => n18920, ZN => n24407);
   U18615 : NAND3_X1 port map( A1 => n20578, A2 => n17237, A3 => n26841, ZN => 
                           n26612);
   U18622 : NAND3_X1 port map( A1 => n31161, A2 => n18148, A3 => n35813, ZN => 
                           n17688);
   U18623 : NAND3_X2 port map( A1 => n13165, A2 => n25796, A3 => n13164, ZN => 
                           n35251);
   U18624 : XOR2_X1 port map( A1 => n21084, A2 => n30956, Z => n35252);
   U18632 : NAND3_X1 port map( A1 => n13165, A2 => n25796, A3 => n13164, ZN => 
                           n26495);
   U18637 : INV_X1 port map( I => n4671, ZN => n13233);
   U18639 : NOR2_X1 port map( A1 => n28655, A2 => n3664, ZN => n28445);
   U18647 : INV_X1 port map( I => n7464, ZN => n1915);
   U18649 : INV_X1 port map( I => n3687, ZN => n30828);
   U18650 : NOR2_X1 port map( A1 => n32259, A2 => n3687, ZN => n11687);
   U18658 : OAI21_X1 port map( A1 => n22265, A2 => n22266, B => n3687, ZN => 
                           n22070);
   U18660 : OAI21_X1 port map( A1 => n12023, A2 => n3687, B => n17307, ZN => 
                           n21263);
   U18666 : XOR2_X1 port map( A1 => n5849, A2 => n5851, Z => n35256);
   U18676 : AND2_X2 port map( A1 => n13156, A2 => n14757, Z => n35258);
   U18699 : NAND2_X1 port map( A1 => n29616, A2 => n29623, ZN => n29622);
   U18709 : NAND2_X1 port map( A1 => n29623, A2 => n35273, ZN => n36382);
   U18712 : NOR2_X1 port map( A1 => n29623, A2 => n29616, ZN => n9046);
   U18713 : INV_X1 port map( I => n31547, ZN => n31898);
   U18724 : INV_X2 port map( I => n1226, ZN => n994);
   U18733 : NOR2_X1 port map( A1 => n22222, A2 => n1688, ZN => n17018);
   U18739 : NAND2_X1 port map( A1 => n30872, A2 => n877, ZN => n6978);
   U18746 : INV_X1 port map( I => n10582, ZN => n9389);
   U18752 : NAND3_X1 port map( A1 => n33591, A2 => n5093, A3 => n16108, ZN => 
                           n28718);
   U18755 : AND2_X2 port map( A1 => n33546, A2 => n15667, Z => n35265);
   U18769 : OAI21_X1 port map( A1 => n25812, A2 => n25813, B => n35671, ZN => 
                           n20451);
   U18772 : INV_X1 port map( I => n9267, ZN => n9295);
   U18776 : OAI22_X2 port map( A1 => n27559, A2 => n34360, B1 => n2381, B2 => 
                           n2380, ZN => n35266);
   U18779 : OAI22_X1 port map( A1 => n27559, A2 => n34360, B1 => n2381, B2 => 
                           n2380, ZN => n27851);
   U18784 : AOI22_X1 port map( A1 => n24701, A2 => n35219, B1 => n33986, B2 => 
                           n13049, ZN => n35267);
   U18793 : AOI22_X1 port map( A1 => n24701, A2 => n35219, B1 => n33986, B2 => 
                           n13049, ZN => n35268);
   U18795 : AOI22_X1 port map( A1 => n24701, A2 => n35219, B1 => n33986, B2 => 
                           n13049, ZN => n25240);
   U18799 : OAI21_X2 port map( A1 => n11486, A2 => n14667, B => n26196, ZN => 
                           n35270);
   U18805 : XNOR2_X1 port map( A1 => n1886, A2 => n1883, ZN => n35271);
   U18808 : NAND2_X1 port map( A1 => n26134, A2 => n9916, ZN => n17003);
   U18809 : NAND2_X1 port map( A1 => n5311, A2 => n2947, ZN => n32861);
   U18826 : NOR2_X1 port map( A1 => n1478, A2 => n6686, ZN => n37039);
   U18833 : AOI22_X2 port map( A1 => n10868, A2 => n29579, B1 => n10869, B2 => 
                           n29580, ZN => n35273);
   U18852 : NAND2_X1 port map( A1 => n32691, A2 => n25798, ZN => n36048);
   U18853 : NAND2_X1 port map( A1 => n25797, A2 => n32691, ZN => n26006);
   U18854 : NAND2_X1 port map( A1 => n31899, A2 => n29568, ZN => n17365);
   U18860 : NAND2_X1 port map( A1 => n23625, A2 => n23430, ZN => n36393);
   U18862 : INV_X1 port map( I => n22854, ZN => n22928);
   U18881 : XOR2_X1 port map( A1 => n36939, A2 => n29817, Z => n11653);
   U18885 : XOR2_X1 port map( A1 => n27663, A2 => n27785, Z => n3320);
   U18888 : XOR2_X1 port map( A1 => n7917, A2 => n11937, Z => n11938);
   U18895 : AOI22_X2 port map( A1 => n7820, A2 => n31787, B1 => n7819, B2 => 
                           n4634, ZN => n7917);
   U18898 : OAI21_X1 port map( A1 => n29618, A2 => n35405, B => n31540, ZN => 
                           n29601);
   U18919 : NAND2_X1 port map( A1 => n27357, A2 => n7632, ZN => n27021);
   U18936 : NOR2_X2 port map( A1 => n10977, A2 => n10976, ZN => n31821);
   U18937 : XOR2_X1 port map( A1 => n10662, A2 => n36002, Z => n2572);
   U18958 : AOI22_X2 port map( A1 => n33663, A2 => n3390, B1 => n32012, B2 => 
                           n3389, ZN => n36866);
   U18973 : NAND2_X2 port map( A1 => n14548, A2 => n35280, ZN => n11321);
   U18977 : XOR2_X1 port map( A1 => n3387, A2 => n20718, Z => n3386);
   U18982 : NAND2_X1 port map( A1 => n1226, A2 => n995, ZN => n8453);
   U18986 : NOR2_X2 port map( A1 => n32444, A2 => n35573, ZN => n1226);
   U18996 : NOR2_X2 port map( A1 => n15465, A2 => n15464, ZN => n27178);
   U19002 : XOR2_X1 port map( A1 => n17703, A2 => n8602, Z => n2615);
   U19013 : XOR2_X1 port map( A1 => n6477, A2 => n16216, Z => n8247);
   U19029 : XOR2_X1 port map( A1 => n22733, A2 => n22734, Z => n35286);
   U19060 : NAND2_X2 port map( A1 => n24585, A2 => n24582, ZN => n5063);
   U19062 : NAND2_X2 port map( A1 => n35294, A2 => n35293, ZN => n31355);
   U19065 : NAND2_X2 port map( A1 => n36705, A2 => n7186, ZN => n33765);
   U19066 : XOR2_X1 port map( A1 => n35255, A2 => n31524, Z => n19067);
   U19075 : NOR2_X2 port map( A1 => n32866, A2 => n5535, ZN => n7464);
   U19079 : NAND2_X1 port map( A1 => n20830, A2 => n29481, ZN => n18290);
   U19091 : NAND2_X2 port map( A1 => n17929, A2 => n17928, ZN => n13029);
   U19099 : NAND3_X1 port map( A1 => n1755, A2 => n36207, A3 => n33861, ZN => 
                           n35330);
   U19106 : INV_X2 port map( I => n2722, ZN => n27583);
   U19110 : AOI22_X2 port map( A1 => n8686, A2 => n7596, B1 => n15142, B2 => 
                           n9646, ZN => n2722);
   U19119 : INV_X2 port map( I => n35300, ZN => n800);
   U19151 : OR2_X2 port map( A1 => n21933, A2 => n36062, Z => n21932);
   U19152 : BUF_X2 port map( I => n27792, Z => n35303);
   U19156 : OAI21_X2 port map( A1 => n16282, A2 => n16283, B => n16281, ZN => 
                           n32886);
   U19159 : NAND2_X2 port map( A1 => n22814, A2 => n22815, ZN => n35534);
   U19160 : AOI21_X2 port map( A1 => n4349, A2 => n4350, B => n31714, ZN => 
                           n24495);
   U19166 : XOR2_X1 port map( A1 => n11236, A2 => n27204, Z => n9196);
   U19180 : XOR2_X1 port map( A1 => n18833, A2 => n21163, Z => n33152);
   U19181 : XNOR2_X1 port map( A1 => n26571, A2 => n12221, ZN => n12903);
   U19189 : MUX2_X1 port map( I0 => n12396, I1 => n39001, S => n23517, Z => 
                           n17788);
   U19202 : XOR2_X1 port map( A1 => n18857, A2 => n24024, Z => n17000);
   U19205 : AOI21_X2 port map( A1 => n28202, A2 => n28203, B => n35309, ZN => 
                           n28680);
   U19213 : OAI21_X2 port map( A1 => n4107, A2 => n14750, B => n35310, ZN => 
                           n23358);
   U19214 : XOR2_X1 port map( A1 => n22735, A2 => n22663, Z => n3800);
   U19222 : XOR2_X1 port map( A1 => n2233, A2 => n19094, Z => n22735);
   U19244 : AOI21_X2 port map( A1 => n6381, A2 => n21787, B => n35315, ZN => 
                           n31960);
   U19245 : AND2_X1 port map( A1 => n21659, A2 => n21660, Z => n35315);
   U19270 : AOI21_X2 port map( A1 => n11187, A2 => n23477, B => n35322, ZN => 
                           n11183);
   U19283 : XOR2_X1 port map( A1 => n16191, A2 => n35323, Z => n30607);
   U19290 : XOR2_X1 port map( A1 => n16190, A2 => n34139, Z => n35323);
   U19301 : NAND2_X2 port map( A1 => n8106, A2 => n8107, ZN => n35900);
   U19303 : XOR2_X1 port map( A1 => n28870, A2 => n35324, Z => n35857);
   U19313 : AOI22_X2 port map( A1 => n35326, A2 => n16206, B1 => n4871, B2 => 
                           n28548, ZN => n15780);
   U19314 : OAI21_X2 port map( A1 => n14631, A2 => n25373, B => n25327, ZN => 
                           n35327);
   U19348 : NAND2_X2 port map( A1 => n17739, A2 => n11388, ZN => n8627);
   U19352 : XOR2_X1 port map( A1 => n25184, A2 => n25176, Z => n25310);
   U19353 : NAND2_X2 port map( A1 => n17904, A2 => n24813, ZN => n25184);
   U19354 : XOR2_X1 port map( A1 => n20065, A2 => n215, Z => n35543);
   U19356 : NOR2_X1 port map( A1 => n27590, A2 => n27591, ZN => n35334);
   U19357 : INV_X4 port map( I => n11678, ZN => n35377);
   U19358 : AOI22_X2 port map( A1 => n35335, A2 => n20815, B1 => n7052, B2 => 
                           n591, ZN => n35448);
   U19359 : NOR2_X2 port map( A1 => n6696, A2 => n2366, ZN => n35335);
   U19361 : XOR2_X1 port map( A1 => n2623, A2 => n2622, Z => n25488);
   U19362 : XOR2_X1 port map( A1 => n26211, A2 => n19900, Z => n26836);
   U19363 : AOI22_X1 port map( A1 => n11446, A2 => n11448, B1 => n32079, B2 => 
                           n32508, ZN => n35340);
   U19364 : XOR2_X1 port map( A1 => n29124, A2 => n28874, Z => n28916);
   U19370 : NAND3_X1 port map( A1 => n14519, A2 => n20605, A3 => n33012, ZN => 
                           n35336);
   U19376 : AOI22_X2 port map( A1 => n7908, A2 => n11803, B1 => n36328, B2 => 
                           n11429, ZN => n7907);
   U19392 : XOR2_X1 port map( A1 => n8922, A2 => n8923, Z => n11780);
   U19396 : XOR2_X1 port map( A1 => n24933, A2 => n34564, Z => n24974);
   U19399 : NAND2_X1 port map( A1 => n35500, A2 => n17132, ZN => n8931);
   U19410 : XOR2_X1 port map( A1 => n25262, A2 => n30519, Z => n12749);
   U19423 : XOR2_X1 port map( A1 => n35340, A2 => n30130, Z => Ciphertext(167))
                           ;
   U19426 : INV_X2 port map( I => n33252, ZN => n35627);
   U19438 : OAI21_X1 port map( A1 => n29956, A2 => n29863, B => n10679, ZN => 
                           n35342);
   U19439 : XOR2_X1 port map( A1 => n35343, A2 => n31815, Z => n22942);
   U19441 : XOR2_X1 port map( A1 => n11887, A2 => n34132, Z => n36971);
   U19443 : NAND2_X2 port map( A1 => n27198, A2 => n4353, ZN => n27397);
   U19444 : INV_X2 port map( I => n26039, ZN => n25830);
   U19445 : NAND2_X2 port map( A1 => n35371, A2 => n2248, ZN => n26039);
   U19453 : XOR2_X1 port map( A1 => n5917, A2 => n9948, Z => n32026);
   U19457 : NOR2_X2 port map( A1 => n1129, A2 => n24360, ZN => n11361);
   U19467 : AOI21_X2 port map( A1 => n30355, A2 => n5935, B => n35345, ZN => 
                           n31959);
   U19475 : XOR2_X1 port map( A1 => n12762, A2 => n12760, Z => n14287);
   U19486 : NAND2_X2 port map( A1 => n71, A2 => n70, ZN => n30574);
   U19500 : INV_X2 port map( I => n16260, ZN => n29412);
   U19504 : NAND2_X2 port map( A1 => n12067, A2 => n35348, ZN => n24877);
   U19506 : NAND2_X2 port map( A1 => n17095, A2 => n31014, ZN => n27402);
   U19512 : XOR2_X1 port map( A1 => n13724, A2 => n21323, Z => n13794);
   U19513 : NAND2_X2 port map( A1 => n35353, A2 => n38168, ZN => n32999);
   U19523 : XOR2_X1 port map( A1 => n5918, A2 => n5920, Z => n8250);
   U19526 : NAND2_X1 port map( A1 => n35813, A2 => n8430, ZN => n8426);
   U19529 : NAND2_X2 port map( A1 => n35355, A2 => n23500, ZN => n17937);
   U19533 : NAND2_X2 port map( A1 => n11323, A2 => n11322, ZN => n19759);
   U19537 : XOR2_X1 port map( A1 => n29127, A2 => n29050, Z => n29292);
   U19555 : NOR2_X1 port map( A1 => n11296, A2 => n975, ZN => n2823);
   U19559 : NAND2_X2 port map( A1 => n6978, A2 => n6980, ZN => n13880);
   U19579 : INV_X4 port map( I => n27349, ZN => n993);
   U19584 : NAND2_X2 port map( A1 => n583, A2 => n21008, ZN => n27349);
   U19595 : XOR2_X1 port map( A1 => Plaintext(8), A2 => Key(8), Z => n35359);
   U19597 : XOR2_X1 port map( A1 => n14110, A2 => n14109, Z => n23189);
   U19600 : AOI22_X2 port map( A1 => n29458, A2 => n19065, B1 => n29454, B2 => 
                           n29455, ZN => n12479);
   U19606 : NAND2_X2 port map( A1 => n12426, A2 => n12175, ZN => n35376);
   U19614 : NAND2_X1 port map( A1 => n14477, A2 => n33840, ZN => n23547);
   U19615 : NAND2_X2 port map( A1 => n12508, A2 => n36001, ZN => n14477);
   U19618 : NOR2_X1 port map( A1 => n31673, A2 => n35450, ZN => n14509);
   U19624 : AOI22_X1 port map( A1 => n30028, A2 => n30027, B1 => n33311, B2 => 
                           n30031, ZN => n18313);
   U19630 : AND2_X1 port map( A1 => n3092, A2 => n27484, Z => n20528);
   U19637 : AOI22_X2 port map( A1 => n6472, A2 => n35696, B1 => n8494, B2 => 
                           n18810, ZN => n35362);
   U19650 : XOR2_X1 port map( A1 => n4209, A2 => n35363, Z => n36390);
   U19651 : XOR2_X1 port map( A1 => n2126, A2 => n12437, Z => n35363);
   U19656 : XOR2_X1 port map( A1 => n27478, A2 => n27850, Z => n27606);
   U19657 : NAND2_X2 port map( A1 => n11040, A2 => n11037, ZN => n27850);
   U19663 : XOR2_X1 port map( A1 => n27495, A2 => n27833, Z => n27646);
   U19664 : XNOR2_X1 port map( A1 => n39161, A2 => n23996, ZN => n6291);
   U19682 : NOR3_X1 port map( A1 => n25498, A2 => n15036, A3 => n14401, ZN => 
                           n25382);
   U19695 : XOR2_X1 port map( A1 => n36971, A2 => n6880, Z => n31078);
   U19697 : NOR2_X1 port map( A1 => n28742, A2 => n17583, ZN => n35370);
   U19702 : OAI21_X2 port map( A1 => n35931, A2 => n33669, B => n35374, ZN => 
                           n33283);
   U19723 : NAND2_X2 port map( A1 => n8656, A2 => n6694, ZN => n8532);
   U19734 : XOR2_X1 port map( A1 => n13001, A2 => n5284, Z => n411);
   U19735 : AOI21_X2 port map( A1 => n14588, A2 => n30434, B => n27231, ZN => 
                           n18641);
   U19737 : OAI22_X2 port map( A1 => n27898, A2 => n28594, B1 => n7905, B2 => 
                           n31088, ZN => n16357);
   U19750 : AOI21_X2 port map( A1 => n14410, A2 => n1024, B => n31574, ZN => 
                           n2461);
   U19752 : NAND2_X2 port map( A1 => n35467, A2 => n8737, ZN => n8683);
   U19762 : AOI21_X2 port map( A1 => n17744, A2 => n36210, B => n35386, ZN => 
                           n17742);
   U19763 : NOR3_X2 port map( A1 => n14901, A2 => n23552, A3 => n34012, ZN => 
                           n35386);
   U19764 : NAND2_X2 port map( A1 => n35387, A2 => n6087, ZN => n8668);
   U19766 : OAI21_X2 port map( A1 => n22956, A2 => n22958, B => n22955, ZN => 
                           n35387);
   U19769 : XOR2_X1 port map( A1 => n27834, A2 => n30104, Z => n35389);
   U19772 : AND2_X1 port map( A1 => n24866, A2 => n36385, Z => n24499);
   U19773 : NAND2_X2 port map( A1 => n24324, A2 => n24323, ZN => n24866);
   U19774 : XOR2_X1 port map( A1 => n6164, A2 => n35390, Z => n11);
   U19778 : XOR2_X1 port map( A1 => n14098, A2 => n3140, Z => n35390);
   U19781 : OAI21_X2 port map( A1 => n5306, A2 => n19480, B => n35391, ZN => 
                           n30210);
   U19784 : NAND3_X1 port map( A1 => n17104, A2 => n35180, A3 => n17103, ZN => 
                           n35392);
   U19787 : OAI21_X2 port map( A1 => n10468, A2 => n34723, B => n1580, ZN => 
                           n9528);
   U19789 : AOI22_X2 port map( A1 => n35394, A2 => n38303, B1 => n31270, B2 => 
                           n5, ZN => n5613);
   U19810 : NAND2_X2 port map( A1 => n18224, A2 => n18223, ZN => n28560);
   U19813 : AND2_X1 port map( A1 => n29880, A2 => n10294, Z => n31968);
   U19818 : INV_X2 port map( I => n35395, ZN => n20359);
   U19832 : AOI21_X2 port map( A1 => n13010, A2 => n9350, B => n39316, ZN => 
                           n9349);
   U19837 : OAI21_X2 port map( A1 => n14474, A2 => n17018, B => n196, ZN => 
                           n35400);
   U19840 : NAND2_X2 port map( A1 => n33485, A2 => n35401, ZN => n35992);
   U19842 : INV_X1 port map( I => n35402, ZN => n1785);
   U19846 : AOI21_X1 port map( A1 => n6274, A2 => n6491, B => n6273, ZN => 
                           n35402);
   U19852 : INV_X1 port map( I => n9360, ZN => n35841);
   U19854 : OR2_X1 port map( A1 => n33948, A2 => n31250, Z => n19964);
   U19870 : OR2_X1 port map( A1 => n29622, A2 => n35405, Z => n17176);
   U19897 : XOR2_X1 port map( A1 => n23887, A2 => n23713, Z => n6277);
   U19905 : INV_X2 port map( I => n35407, ZN => n8556);
   U19908 : XNOR2_X1 port map( A1 => n8557, A2 => n26373, ZN => n35407);
   U19934 : NAND2_X1 port map( A1 => n11838, A2 => n38579, ZN => n35414);
   U19936 : NAND2_X1 port map( A1 => n7220, A2 => n7219, ZN => n35415);
   U19940 : XNOR2_X1 port map( A1 => n1669, A2 => n11541, ZN => n35642);
   U19942 : XOR2_X1 port map( A1 => n6572, A2 => n31791, Z => n7787);
   U19945 : NAND2_X2 port map( A1 => n1865, A2 => n1864, ZN => n22620);
   U19956 : XOR2_X1 port map( A1 => n6460, A2 => n24150, Z => n31348);
   U19960 : NAND2_X1 port map( A1 => n15301, A2 => n1403, ZN => n36403);
   U19963 : XOR2_X1 port map( A1 => n18886, A2 => n28933, Z => n431);
   U19965 : NAND2_X2 port map( A1 => n32186, A2 => n16576, ZN => n27571);
   U19970 : NAND2_X2 port map( A1 => n1351, A2 => n17938, ZN => n21497);
   U19974 : NAND3_X1 port map( A1 => n31184, A2 => n30368, A3 => n24406, ZN => 
                           n30850);
   U19979 : AOI22_X2 port map( A1 => n37257, A2 => n28246, B1 => n37451, B2 => 
                           n19003, ZN => n35420);
   U19980 : XOR2_X1 port map( A1 => n8957, A2 => n27569, Z => n35421);
   U19981 : NAND3_X2 port map( A1 => n1763, A2 => n23167, A3 => n22975, ZN => 
                           n20564);
   U19984 : NAND3_X2 port map( A1 => n1906, A2 => n35735, A3 => n30635, ZN => 
                           n35422);
   U19986 : AOI22_X2 port map( A1 => n35424, A2 => n19132, B1 => n35423, B2 => 
                           n1221, ZN => n27785);
   U19993 : XOR2_X1 port map( A1 => n24025, A2 => n19904, Z => n11180);
   U19995 : NAND2_X2 port map( A1 => n35600, A2 => n321, ZN => n24025);
   U19998 : XOR2_X1 port map( A1 => n11828, A2 => n16439, Z => n35425);
   U20013 : NAND2_X1 port map( A1 => n22928, A2 => n22994, ZN => n22555);
   U20014 : NAND2_X1 port map( A1 => n20616, A2 => n170, ZN => n29993);
   U20016 : XOR2_X1 port map( A1 => n9043, A2 => n18279, Z => n33010);
   U20020 : NAND3_X2 port map( A1 => n3275, A2 => n3276, A3 => n3274, ZN => 
                           n9043);
   U20027 : BUF_X4 port map( I => n8267, Z => n35921);
   U20044 : AOI21_X1 port map( A1 => n18783, A2 => n18782, B => n30037, ZN => 
                           n36848);
   U20048 : NOR2_X1 port map( A1 => n4964, A2 => n35427, ZN => n32696);
   U20059 : OAI21_X2 port map( A1 => n7212, A2 => n22496, B => n36660, ZN => 
                           n35920);
   U20084 : NAND2_X2 port map( A1 => n12993, A2 => n12991, ZN => n11067);
   U20088 : AND2_X1 port map( A1 => n33980, A2 => n12187, Z => n19003);
   U20103 : XOR2_X1 port map( A1 => n35435, A2 => n14046, Z => n35769);
   U20110 : NAND2_X2 port map( A1 => n6252, A2 => n29558, ZN => n29543);
   U20112 : NAND2_X2 port map( A1 => n6253, A2 => n14850, ZN => n29558);
   U20131 : XOR2_X1 port map( A1 => n18106, A2 => n26605, Z => n36915);
   U20133 : XOR2_X1 port map( A1 => n8833, A2 => n17757, Z => n26605);
   U20137 : XOR2_X1 port map( A1 => n35746, A2 => n35747, Z => n4256);
   U20141 : NAND2_X2 port map( A1 => n35437, A2 => n14995, ZN => n21864);
   U20160 : INV_X4 port map( I => n23350, ZN => n36027);
   U20170 : XOR2_X1 port map( A1 => n27837, A2 => n3207, Z => n35438);
   U20171 : AOI21_X2 port map( A1 => n16750, A2 => n16749, B => n35439, ZN => 
                           n7728);
   U20185 : OAI22_X2 port map( A1 => n20414, A2 => n3120, B1 => n24849, B2 => 
                           n33344, ZN => n35439);
   U20187 : NAND3_X2 port map( A1 => n27124, A2 => n27125, A3 => n27129, ZN => 
                           n16736);
   U20189 : NOR2_X1 port map( A1 => n35679, A2 => n25770, ZN => n30568);
   U20203 : NAND2_X1 port map( A1 => n38395, A2 => n17864, ZN => n64);
   U20205 : NOR2_X2 port map( A1 => n10295, A2 => n35441, ZN => n23634);
   U20209 : INV_X2 port map( I => n29005, ZN => n4095);
   U20211 : XOR2_X1 port map( A1 => n3938, A2 => n34183, Z => n29005);
   U20216 : AOI22_X2 port map( A1 => n12891, A2 => n12890, B1 => n36609, B2 => 
                           n34172, ZN => n12889);
   U20225 : XOR2_X1 port map( A1 => n12857, A2 => n7673, Z => n35836);
   U20229 : XOR2_X1 port map( A1 => n35446, A2 => n22438, Z => n35445);
   U20231 : XOR2_X1 port map( A1 => n29253, A2 => n9930, Z => n16553);
   U20232 : NAND4_X2 port map( A1 => n22820, A2 => n7683, A3 => n18856, A4 => 
                           n31748, ZN => n18204);
   U20235 : NAND3_X2 port map( A1 => n17971, A2 => n24778, A3 => n24777, ZN => 
                           n16627);
   U20241 : NAND2_X2 port map( A1 => n16700, A2 => n31638, ZN => n31287);
   U20250 : INV_X2 port map( I => n35450, ZN => n30279);
   U20251 : XNOR2_X1 port map( A1 => n20516, A2 => n20716, ZN => n35450);
   U20273 : NAND3_X2 port map( A1 => n36785, A2 => n16098, A3 => n23338, ZN => 
                           n23658);
   U20274 : INV_X1 port map( I => n32630, ZN => n35569);
   U20277 : NOR2_X2 port map( A1 => n35452, A2 => n7859, ZN => n31862);
   U20281 : NOR2_X2 port map( A1 => n20404, A2 => n33788, ZN => n5955);
   U20284 : NAND2_X2 port map( A1 => n35454, A2 => n25810, ZN => n26437);
   U20285 : NAND2_X2 port map( A1 => n3153, A2 => n3857, ZN => n30076);
   U20286 : AOI21_X2 port map( A1 => n22015, A2 => n20034, B => n22165, ZN => 
                           n35734);
   U20299 : INV_X2 port map( I => n35455, ZN => n14418);
   U20301 : XOR2_X1 port map( A1 => Plaintext(138), A2 => Key(138), Z => n35455
                           );
   U20307 : XOR2_X1 port map( A1 => n35457, A2 => n22667, Z => n10963);
   U20333 : INV_X2 port map( I => n35462, ZN => n24155);
   U20336 : NOR2_X2 port map( A1 => n12064, A2 => n19142, ZN => n35462);
   U20337 : INV_X2 port map( I => n15047, ZN => n17197);
   U20342 : NAND2_X1 port map( A1 => n36623, A2 => n28729, ZN => n15296);
   U20343 : XOR2_X1 port map( A1 => n35463, A2 => n26480, Z => n30551);
   U20346 : NAND2_X2 port map( A1 => n9087, A2 => n9086, ZN => n26480);
   U20347 : INV_X2 port map( I => n27532, ZN => n35464);
   U20348 : NAND2_X1 port map( A1 => n20724, A2 => n29410, ZN => n35677);
   U20365 : XOR2_X1 port map( A1 => n19064, A2 => n25007, Z => n10717);
   U20367 : XOR2_X1 port map( A1 => n12430, A2 => n3395, Z => n35468);
   U20370 : INV_X2 port map( I => n31971, ZN => n35469);
   U20375 : OAI22_X2 port map( A1 => n3714, A2 => n32351, B1 => n2928, B2 => 
                           n3715, ZN => n35470);
   U20376 : XOR2_X1 port map( A1 => n3330, A2 => n35471, Z => n36334);
   U20378 : XOR2_X1 port map( A1 => n35472, A2 => n25033, Z => n8713);
   U20380 : XOR2_X1 port map( A1 => n24997, A2 => n25290, Z => n25033);
   U20387 : XOR2_X1 port map( A1 => n7337, A2 => n35532, Z => n10380);
   U20390 : XOR2_X1 port map( A1 => n22766, A2 => n22624, Z => n7337);
   U20391 : NOR2_X1 port map( A1 => n35474, A2 => n22253, ZN => n17409);
   U20393 : NAND2_X1 port map( A1 => n12930, A2 => n10242, ZN => n35474);
   U20396 : INV_X2 port map( I => n35476, ZN => n2752);
   U20398 : XOR2_X1 port map( A1 => n2754, A2 => n2753, Z => n35476);
   U20410 : XOR2_X1 port map( A1 => n38191, A2 => n12480, Z => n35480);
   U20411 : XOR2_X1 port map( A1 => n24026, A2 => n5238, Z => n35481);
   U20414 : NAND3_X2 port map( A1 => n35483, A2 => n39813, A3 => n13580, ZN => 
                           n10638);
   U20426 : XNOR2_X1 port map( A1 => n17727, A2 => n22562, ZN => n22733);
   U20429 : NAND2_X2 port map( A1 => n6723, A2 => n6721, ZN => n22562);
   U20436 : XNOR2_X1 port map( A1 => n26455, A2 => n29785, ZN => n36511);
   U20450 : NOR2_X2 port map( A1 => n4147, A2 => n17887, ZN => n4148);
   U20457 : INV_X2 port map( I => n31474, ZN => n35705);
   U20460 : XOR2_X1 port map( A1 => n4131, A2 => n36264, Z => n31474);
   U20461 : XOR2_X1 port map( A1 => n39161, A2 => n19629, Z => n23924);
   U20467 : AOI21_X2 port map( A1 => n24506, A2 => n9212, B => n36017, ZN => 
                           n18393);
   U20479 : NAND2_X1 port map( A1 => n14396, A2 => n19586, ZN => n15080);
   U20480 : NOR2_X2 port map( A1 => n31037, A2 => n35487, ZN => n23969);
   U20481 : OAI22_X2 port map( A1 => n23621, A2 => n33496, B1 => n23284, B2 => 
                           n23452, ZN => n35487);
   U20487 : XOR2_X1 port map( A1 => n35490, A2 => n2743, Z => n2742);
   U20488 : XOR2_X1 port map( A1 => n33806, A2 => n22382, Z => n35490);
   U20489 : OAI22_X2 port map( A1 => n13306, A2 => n13304, B1 => n32616, B2 => 
                           n30274, ZN => n23963);
   U20490 : NAND2_X2 port map( A1 => n28345, A2 => n28347, ZN => n28717);
   U20505 : XOR2_X1 port map( A1 => n36863, A2 => n35494, Z => n33553);
   U20506 : XOR2_X1 port map( A1 => n27763, A2 => n27762, Z => n35494);
   U20513 : XOR2_X1 port map( A1 => n32200, A2 => n29247, Z => n12853);
   U20516 : OR2_X1 port map( A1 => n11728, A2 => n18246, Z => n35495);
   U20517 : NAND2_X2 port map( A1 => n28140, A2 => n28139, ZN => n35496);
   U20518 : XOR2_X1 port map( A1 => n26521, A2 => n35498, Z => n11740);
   U20519 : XOR2_X1 port map( A1 => n31941, A2 => n26407, Z => n35498);
   U20521 : AND2_X1 port map( A1 => n28586, A2 => n11030, Z => n36031);
   U20523 : XOR2_X1 port map( A1 => n18635, A2 => n5203, Z => n31933);
   U20525 : XOR2_X1 port map( A1 => n22784, A2 => n1710, Z => n12516);
   U20526 : XOR2_X1 port map( A1 => n14388, A2 => n16553, Z => n16552);
   U20529 : NAND2_X1 port map( A1 => n10171, A2 => n27304, ZN => n35906);
   U20543 : INV_X2 port map( I => n32854, ZN => n35506);
   U20546 : INV_X1 port map( I => n16203, ZN => n35508);
   U20551 : NOR2_X1 port map( A1 => n11030, A2 => n36076, ZN => n36032);
   U20552 : OR2_X1 port map( A1 => n8527, A2 => n38591, Z => n26443);
   U20564 : XOR2_X1 port map( A1 => n25293, A2 => n35511, Z => n35510);
   U20567 : NAND2_X1 port map( A1 => n33086, A2 => n22264, ZN => n35513);
   U20591 : NAND3_X1 port map( A1 => n15215, A2 => n9594, A3 => n16114, ZN => 
                           n35763);
   U20598 : AOI21_X1 port map( A1 => n29389, A2 => n29497, B => n36275, ZN => 
                           n35517);
   U20599 : NAND2_X2 port map( A1 => n6954, A2 => n6953, ZN => n7552);
   U20614 : NOR2_X1 port map( A1 => n24795, A2 => n16238, ZN => n35520);
   U20615 : XOR2_X1 port map( A1 => n11207, A2 => n29306, Z => n35728);
   U20626 : NOR2_X2 port map( A1 => n20102, A2 => n30059, ZN => n6496);
   U20631 : NAND2_X1 port map( A1 => n39676, A2 => n26109, ZN => n25790);
   U20639 : XOR2_X1 port map( A1 => n8371, A2 => n36828, Z => n4898);
   U20668 : AOI21_X2 port map( A1 => n14355, A2 => n26833, B => n7527, ZN => 
                           n26772);
   U20670 : NAND2_X1 port map( A1 => n39155, A2 => n18708, ZN => n9507);
   U20678 : NAND2_X2 port map( A1 => n35689, A2 => n1642, ZN => n23392);
   U20695 : XOR2_X1 port map( A1 => n21207, A2 => n7380, Z => n25552);
   U20704 : NAND2_X2 port map( A1 => n22119, A2 => n22116, ZN => n3687);
   U20705 : AOI22_X2 port map( A1 => n2164, A2 => n31198, B1 => n31257, B2 => 
                           n35968, ZN => n25303);
   U20726 : NOR2_X1 port map( A1 => n13555, A2 => n11449, ZN => n6170);
   U20729 : NAND2_X1 port map( A1 => n19204, A2 => n14636, ZN => n35535);
   U20730 : BUF_X2 port map( I => n23250, Z => n35536);
   U20735 : OAI21_X2 port map( A1 => n10452, A2 => n31958, B => n35541, ZN => 
                           n17849);
   U20737 : XOR2_X1 port map( A1 => n27538, A2 => n34094, Z => n35542);
   U20738 : INV_X1 port map( I => n35233, ZN => n12248);
   U20748 : NOR2_X2 port map( A1 => n22396, A2 => n22397, ZN => n22408);
   U20766 : XOR2_X1 port map( A1 => n22517, A2 => n4123, Z => n22382);
   U20772 : XOR2_X1 port map( A1 => n35544, A2 => n27784, Z => n33522);
   U20786 : XOR2_X1 port map( A1 => n5153, A2 => n29145, Z => n1740);
   U20787 : NAND2_X2 port map( A1 => n28752, A2 => n28751, ZN => n29145);
   U20791 : AND2_X1 port map( A1 => n35550, A2 => n33538, Z => n17787);
   U20794 : NAND2_X1 port map( A1 => n23517, A2 => n19671, ZN => n35550);
   U20801 : NAND3_X2 port map( A1 => n31168, A2 => n16435, A3 => n35553, ZN => 
                           n22728);
   U20802 : AOI22_X1 port map( A1 => n10651, A2 => n9876, B1 => n22341, B2 => 
                           n15350, ZN => n35553);
   U20803 : XOR2_X1 port map( A1 => n8909, A2 => n774, Z => n35554);
   U20818 : NAND2_X2 port map( A1 => n17819, A2 => n17820, ZN => n21802);
   U20821 : XOR2_X1 port map( A1 => n4442, A2 => n35556, Z => n10455);
   U20822 : XOR2_X1 port map( A1 => n22609, A2 => n20350, Z => n35556);
   U20828 : NAND2_X2 port map( A1 => n28460, A2 => n28378, ZN => n31390);
   U20842 : NAND2_X2 port map( A1 => n10, A2 => n14066, ZN => n33840);
   U20858 : NOR2_X1 port map( A1 => n21914, A2 => n938, ZN => n21915);
   U20863 : XOR2_X1 port map( A1 => n19194, A2 => n10413, Z => n10427);
   U20887 : NAND2_X1 port map( A1 => n16832, A2 => n10733, ZN => n36852);
   U20889 : NAND2_X2 port map( A1 => n35563, A2 => n27938, ZN => n16108);
   U20890 : NAND2_X1 port map( A1 => n33613, A2 => n33611, ZN => n35563);
   U20918 : NAND2_X2 port map( A1 => n23355, A2 => n37523, ZN => n23248);
   U20925 : XOR2_X1 port map( A1 => n35566, A2 => n34062, Z => n36454);
   U20930 : XOR2_X1 port map( A1 => n6034, A2 => n5055, Z => n35566);
   U20931 : XOR2_X1 port map( A1 => n8183, A2 => n35267, Z => n24702);
   U20941 : NOR2_X2 port map( A1 => n33032, A2 => n7258, ZN => n35568);
   U20946 : NOR2_X2 port map( A1 => n21420, A2 => n21419, ZN => n36371);
   U20953 : AOI21_X1 port map( A1 => n29645, A2 => n35572, B => n37879, ZN => 
                           n17383);
   U20958 : NAND2_X2 port map( A1 => n22000, A2 => n20298, ZN => n17189);
   U20962 : NAND2_X2 port map( A1 => n17882, A2 => n15652, ZN => n22484);
   U20982 : XOR2_X1 port map( A1 => n2387, A2 => n2388, Z => n31403);
   U20983 : NOR2_X1 port map( A1 => n7445, A2 => n36321, ZN => n20029);
   U20989 : NAND2_X2 port map( A1 => n35948, A2 => n16184, ZN => n36321);
   U21018 : NAND2_X2 port map( A1 => n24662, A2 => n35578, ZN => n35577);
   U21028 : NOR2_X1 port map( A1 => n18383, A2 => n14456, ZN => n19242);
   U21034 : XOR2_X1 port map( A1 => n3709, A2 => n5255, Z => n33057);
   U21042 : XOR2_X1 port map( A1 => n5652, A2 => n15960, Z => n18886);
   U21045 : NAND2_X2 port map( A1 => n6809, A2 => n30748, ZN => n5652);
   U21061 : NAND2_X2 port map( A1 => n6712, A2 => n35584, ZN => n23433);
   U21065 : AOI21_X2 port map( A1 => n22996, A2 => n35586, B => n35585, ZN => 
                           n35584);
   U21076 : NOR2_X2 port map( A1 => n23163, A2 => n35586, ZN => n35585);
   U21079 : INV_X2 port map( I => n23164, ZN => n35586);
   U21086 : INV_X2 port map( I => n23530, ZN => n23528);
   U21088 : NAND4_X2 port map( A1 => n33832, A2 => n20741, A3 => n20744, A4 => 
                           n5464, ZN => n23530);
   U21090 : XOR2_X1 port map( A1 => n12853, A2 => n3297, Z => n12055);
   U21100 : OR2_X1 port map( A1 => n37230, A2 => n33788, Z => n24483);
   U21121 : NOR2_X2 port map( A1 => n8190, A2 => n23374, ZN => n35594);
   U21124 : OAI21_X1 port map( A1 => n16880, A2 => n5061, B => n36425, ZN => 
                           n9715);
   U21126 : NOR2_X2 port map( A1 => n12511, A2 => n12512, ZN => n16880);
   U21134 : XOR2_X1 port map( A1 => n35595, A2 => n18255, Z => n30455);
   U21144 : XOR2_X1 port map( A1 => n37042, A2 => n35596, Z => n35595);
   U21153 : INV_X2 port map( I => n22527, ZN => n35596);
   U21160 : NAND2_X2 port map( A1 => n12394, A2 => n7866, ZN => n25691);
   U21161 : NAND2_X2 port map( A1 => n35598, A2 => n5292, ZN => n14890);
   U21164 : NAND2_X2 port map( A1 => n25568, A2 => n25692, ZN => n35598);
   U21166 : XOR2_X1 port map( A1 => n35599, A2 => n26369, Z => n19810);
   U21167 : XOR2_X1 port map( A1 => n26432, A2 => n16169, Z => n35599);
   U21169 : OR2_X2 port map( A1 => n17464, A2 => n5975, Z => n23072);
   U21175 : BUF_X4 port map( I => n7520, Z => n35960);
   U21178 : AOI22_X2 port map( A1 => n36137, A2 => n38244, B1 => n37209, B2 => 
                           n19686, ZN => n35600);
   U21181 : XOR2_X1 port map( A1 => n35601, A2 => n32890, Z => n33788);
   U21198 : XOR2_X1 port map( A1 => n11794, A2 => n5005, Z => n36000);
   U21201 : NAND3_X2 port map( A1 => n19670, A2 => n24965, A3 => n16819, ZN => 
                           n30520);
   U21221 : XOR2_X1 port map( A1 => n5463, A2 => n22667, Z => n9137);
   U21234 : NAND2_X2 port map( A1 => n12816, A2 => n22965, ZN => n23496);
   U21241 : BUF_X2 port map( I => n27852, Z => n35610);
   U21245 : XOR2_X1 port map( A1 => n9449, A2 => n9448, Z => n35614);
   U21248 : NOR2_X1 port map( A1 => n38839, A2 => n17790, ZN => n8201);
   U21250 : OAI21_X2 port map( A1 => n14326, A2 => n2760, B => n35616, ZN => 
                           n2281);
   U21257 : NOR2_X2 port map( A1 => n8927, A2 => n35619, ZN => n33493);
   U21262 : NOR3_X2 port map( A1 => n1125, A2 => n9371, A3 => n35890, ZN => 
                           n35619);
   U21267 : XOR2_X1 port map( A1 => n8469, A2 => n8471, Z => n29149);
   U21268 : NAND2_X2 port map( A1 => n21786, A2 => n35623, ZN => n22294);
   U21275 : XOR2_X1 port map( A1 => n27500, A2 => n26916, Z => n35626);
   U21288 : XOR2_X1 port map( A1 => n26593, A2 => n36383, Z => n15674);
   U21289 : XOR2_X1 port map( A1 => n26340, A2 => n6757, Z => n26593);
   U21291 : OAI22_X1 port map( A1 => n29414, A2 => n29413, B1 => n29415, B2 => 
                           n29416, ZN => n29417);
   U21298 : XOR2_X1 port map( A1 => n25237, A2 => n11964, Z => n15011);
   U21302 : NAND2_X1 port map( A1 => n19588, A2 => n14561, ZN => n3039);
   U21318 : XOR2_X1 port map( A1 => n24019, A2 => n35630, Z => n16321);
   U21325 : XOR2_X1 port map( A1 => n24020, A2 => n23890, Z => n35630);
   U21326 : XOR2_X1 port map( A1 => n35631, A2 => n24022, Z => n13504);
   U21338 : XOR2_X1 port map( A1 => n24023, A2 => n20317, Z => n35631);
   U21340 : NOR3_X2 port map( A1 => n12927, A2 => n14769, A3 => n1354, ZN => 
                           n3480);
   U21354 : XOR2_X1 port map( A1 => n35636, A2 => n848, Z => n36283);
   U21365 : XOR2_X1 port map( A1 => n24011, A2 => n30150, Z => n35640);
   U21400 : INV_X1 port map( I => n32103, ZN => n17403);
   U21401 : XOR2_X1 port map( A1 => n35642, A2 => n22279, Z => n32103);
   U21420 : NAND3_X2 port map( A1 => n585, A2 => n32507, A3 => n609, ZN => 
                           n35647);
   U21455 : OAI22_X2 port map( A1 => n22333, A2 => n20308, B1 => n20961, B2 => 
                           n937, ZN => n12267);
   U21458 : OR2_X1 port map( A1 => n33786, A2 => n35932, Z => n8416);
   U21466 : NAND3_X2 port map( A1 => n38653, A2 => n34190, A3 => n13485, ZN => 
                           n13406);
   U21480 : OAI21_X1 port map( A1 => n30042, A2 => n30043, B => n5348, ZN => 
                           n35653);
   U21483 : NAND2_X1 port map( A1 => n27213, A2 => n16043, ZN => n17152);
   U21485 : NOR2_X2 port map( A1 => n8627, A2 => n11387, ZN => n27213);
   U21491 : NAND2_X2 port map( A1 => n36672, A2 => n16570, ZN => n24417);
   U21492 : OAI22_X1 port map( A1 => n35744, A2 => n13391, B1 => n1240, B2 => 
                           n26093, ZN => n35655);
   U21493 : NAND3_X2 port map( A1 => n13695, A2 => n13697, A3 => n13696, ZN => 
                           n18875);
   U21496 : NOR2_X1 port map( A1 => n29946, A2 => n29996, ZN => n6600);
   U21497 : INV_X2 port map( I => n29994, ZN => n29946);
   U21501 : XOR2_X1 port map( A1 => n5129, A2 => n10829, Z => n29994);
   U21511 : XOR2_X1 port map( A1 => n343, A2 => n35656, Z => n33695);
   U21514 : NAND3_X1 port map( A1 => n1403, A2 => n37368, A3 => n39828, ZN => 
                           n32762);
   U21518 : NOR2_X2 port map( A1 => n36387, A2 => n20850, ZN => n20849);
   U21523 : INV_X2 port map( I => n5348, ZN => n29997);
   U21543 : XOR2_X1 port map( A1 => n10722, A2 => n38813, Z => n3317);
   U21545 : AND2_X1 port map( A1 => n36833, A2 => n27357, Z => n21170);
   U21555 : XOR2_X1 port map( A1 => n4440, A2 => n22530, Z => n13514);
   U21563 : XOR2_X1 port map( A1 => n12015, A2 => n3239, Z => n22530);
   U21580 : XOR2_X1 port map( A1 => n14346, A2 => n26163, Z => n26401);
   U21583 : NAND2_X2 port map( A1 => n8721, A2 => n8719, ZN => n32366);
   U21589 : AND2_X1 port map( A1 => n35667, A2 => n38282, Z => n20651);
   U21597 : NOR2_X1 port map( A1 => n21365, A2 => n21364, ZN => n35668);
   U21605 : XOR2_X1 port map( A1 => n5553, A2 => n34144, Z => n16558);
   U21610 : XOR2_X1 port map( A1 => n26498, A2 => n4875, Z => n5553);
   U21611 : OAI21_X1 port map( A1 => n10120, A2 => n21839, B => n7278, ZN => 
                           n3868);
   U21619 : OAI21_X2 port map( A1 => n32415, A2 => n14520, B => n20525, ZN => 
                           n35673);
   U21632 : NAND3_X2 port map( A1 => n35675, A2 => n11672, A3 => n8343, ZN => 
                           n22604);
   U21640 : XOR2_X1 port map( A1 => n19640, A2 => n19639, Z => n20524);
   U21653 : XOR2_X1 port map( A1 => n35676, A2 => n29394, Z => Ciphertext(36));
   U21656 : XOR2_X1 port map( A1 => n33509, A2 => n29165, Z => n29816);
   U21658 : NAND2_X2 port map( A1 => n18191, A2 => n28122, ZN => n29165);
   U21659 : NAND2_X1 port map( A1 => n31997, A2 => n35677, ZN => n32462);
   U21670 : XOR2_X1 port map( A1 => n36384, A2 => n900, Z => n35678);
   U21681 : XOR2_X1 port map( A1 => n23886, A2 => n23808, Z => n24060);
   U21683 : NAND2_X2 port map( A1 => n17443, A2 => n17442, ZN => n23886);
   U21689 : INV_X4 port map( I => n35686, ZN => n6977);
   U21692 : NAND3_X2 port map( A1 => n5408, A2 => n36271, A3 => n33581, ZN => 
                           n6014);
   U21717 : INV_X2 port map( I => n35687, ZN => n23165);
   U21737 : NAND2_X2 port map( A1 => n13631, A2 => n21926, ZN => n18595);
   U21738 : XOR2_X1 port map( A1 => n26253, A2 => n26252, Z => n26348);
   U21742 : NAND2_X2 port map( A1 => n11625, A2 => n11623, ZN => n26252);
   U21745 : AOI22_X2 port map( A1 => n12680, A2 => n36716, B1 => n5063, B2 => 
                           n12681, ZN => n35688);
   U21746 : XOR2_X1 port map( A1 => n38021, A2 => n1620, Z => n12026);
   U21749 : INV_X2 port map( I => n37092, ZN => n35689);
   U21759 : OAI22_X1 port map( A1 => n14662, A2 => n33712, B1 => n18238, B2 => 
                           n1606, ZN => n23909);
   U21793 : INV_X2 port map( I => n35693, ZN => n24855);
   U21799 : NAND2_X2 port map( A1 => n15549, A2 => n15550, ZN => n35895);
   U21806 : NAND2_X2 port map( A1 => n28038, A2 => n28039, ZN => n28484);
   U21811 : NAND2_X2 port map( A1 => n13618, A2 => n13621, ZN => n16067);
   U21812 : AOI21_X2 port map( A1 => n35699, A2 => n19856, B => n20832, ZN => 
                           n20831);
   U21820 : NAND2_X2 port map( A1 => n22856, A2 => n19945, ZN => n17917);
   U21823 : XOR2_X1 port map( A1 => n13235, A2 => n22466, Z => n2200);
   U21832 : NAND2_X2 port map( A1 => n4703, A2 => n13629, ZN => n16897);
   U21836 : XOR2_X1 port map( A1 => n18991, A2 => n8183, Z => n24972);
   U21843 : NAND2_X1 port map( A1 => n12119, A2 => n12118, ZN => n33180);
   U21844 : NOR2_X1 port map( A1 => n22222, A2 => n22221, ZN => n15499);
   U21853 : XOR2_X1 port map( A1 => n4201, A2 => n1077, Z => n10396);
   U21860 : INV_X1 port map( I => n29017, ZN => n35702);
   U21879 : NOR2_X2 port map( A1 => n22223, A2 => n22221, ZN => n22135);
   U21881 : NOR2_X2 port map( A1 => n21686, A2 => n21685, ZN => n22223);
   U21882 : XOR2_X1 port map( A1 => n19096, A2 => n11950, Z => n10215);
   U21885 : OAI21_X2 port map( A1 => n30422, A2 => n31698, B => n15208, ZN => 
                           n19096);
   U21891 : XOR2_X1 port map( A1 => n26263, A2 => n35704, Z => n10854);
   U21894 : XOR2_X1 port map( A1 => n26223, A2 => n343, Z => n35704);
   U21895 : AOI21_X1 port map( A1 => n4621, A2 => n9913, B => n1396, ZN => 
                           n6321);
   U21896 : XOR2_X1 port map( A1 => n1929, A2 => n794, Z => n16459);
   U21899 : OR2_X1 port map( A1 => n35732, A2 => n9178, Z => n10795);
   U21900 : XOR2_X1 port map( A1 => n35706, A2 => n3422, Z => n3973);
   U21901 : XOR2_X1 port map( A1 => n31627, A2 => n36999, Z => n35706);
   U21905 : XOR2_X1 port map( A1 => n16378, A2 => n16380, Z => n16388);
   U21907 : INV_X4 port map( I => n32829, ZN => n21248);
   U21921 : INV_X2 port map( I => n35708, ZN => n21036);
   U21924 : NOR2_X1 port map( A1 => n29477, A2 => n7303, ZN => n2449);
   U21931 : XOR2_X1 port map( A1 => n35852, A2 => n27659, Z => n36136);
   U21936 : OR2_X1 port map( A1 => n17607, A2 => n2616, Z => n24798);
   U21943 : XOR2_X1 port map( A1 => n22566, A2 => n35824, Z => n18359);
   U21945 : NAND2_X2 port map( A1 => n9127, A2 => n9126, ZN => n22566);
   U21959 : XOR2_X1 port map( A1 => n15935, A2 => n32610, Z => n15933);
   U21970 : NAND2_X2 port map( A1 => n495, A2 => n1487, ZN => n16520);
   U21972 : NAND2_X2 port map( A1 => n35718, A2 => n16517, ZN => n27607);
   U21978 : XOR2_X1 port map( A1 => n4441, A2 => n22517, Z => n4440);
   U21981 : NAND2_X2 port map( A1 => n1839, A2 => n1837, ZN => n22517);
   U21995 : OAI22_X2 port map( A1 => n1265, A2 => n35893, B1 => n24737, B2 => 
                           n5871, ZN => n24736);
   U21999 : NAND2_X2 port map( A1 => n7845, A2 => n32699, ZN => n25080);
   U22003 : NOR2_X2 port map( A1 => n35723, A2 => n18979, ZN => n36425);
   U22006 : INV_X1 port map( I => n25488, ZN => n220);
   U22011 : INV_X2 port map( I => n35724, ZN => n217);
   U22013 : AOI21_X2 port map( A1 => n1399, A2 => n30220, B => n30159, ZN => 
                           n10568);
   U22014 : XOR2_X1 port map( A1 => n35726, A2 => n15331, Z => n19938);
   U22015 : XOR2_X1 port map( A1 => n411, A2 => n19014, Z => n35726);
   U22042 : NAND2_X1 port map( A1 => n17364, A2 => n29567, ZN => n35731);
   U22050 : NAND2_X2 port map( A1 => n106, A2 => n4138, ZN => n35732);
   U22054 : NAND3_X1 port map( A1 => n35911, A2 => n32575, A3 => n2191, ZN => 
                           n21188);
   U22055 : INV_X2 port map( I => n14213, ZN => n15936);
   U22057 : NOR2_X2 port map( A1 => n16841, A2 => n24416, ZN => n14213);
   U22058 : XOR2_X1 port map( A1 => n27833, A2 => n27731, Z => n17043);
   U22060 : XOR2_X1 port map( A1 => n25194, A2 => n25275, Z => n25103);
   U22061 : NAND2_X2 port map( A1 => n9999, A2 => n4608, ZN => n25275);
   U22066 : AOI21_X2 port map( A1 => n22018, A2 => n22017, B => n35734, ZN => 
                           n22430);
   U22077 : OAI21_X2 port map( A1 => n2190, A2 => n14945, B => n33186, ZN => 
                           n35780);
   U22099 : XOR2_X1 port map( A1 => n28865, A2 => n29252, Z => n28979);
   U22103 : NOR2_X2 port map( A1 => n6046, A2 => n35737, ZN => n36700);
   U22118 : XOR2_X1 port map( A1 => n25286, A2 => n34137, Z => n35741);
   U22123 : XOR2_X1 port map( A1 => n35743, A2 => n6927, Z => n16339);
   U22126 : XOR2_X1 port map( A1 => n27714, A2 => n27805, Z => n35743);
   U22127 : INV_X4 port map( I => n17499, ZN => n1340);
   U22129 : XOR2_X1 port map( A1 => n22458, A2 => n9115, Z => n8172);
   U22130 : XOR2_X1 port map( A1 => n22443, A2 => n8026, Z => n22458);
   U22132 : NOR2_X1 port map( A1 => n15209, A2 => n35179, ZN => n17364);
   U22135 : BUF_X2 port map( I => n33258, Z => n35744);
   U22147 : OAI21_X2 port map( A1 => n16373, A2 => n12533, B => n16372, ZN => 
                           n18407);
   U22151 : XOR2_X1 port map( A1 => n38514, A2 => n36765, Z => n35747);
   U22159 : INV_X1 port map( I => n35748, ZN => n25408);
   U22181 : XOR2_X1 port map( A1 => n27546, A2 => n19808, Z => n5252);
   U22187 : XOR2_X1 port map( A1 => n476, A2 => n5116, Z => n35752);
   U22194 : XOR2_X1 port map( A1 => n32839, A2 => n34151, Z => n36858);
   U22199 : NOR2_X1 port map( A1 => n35756, A2 => n35755, ZN => n30878);
   U22207 : INV_X2 port map( I => n13519, ZN => n35755);
   U22209 : NAND2_X1 port map( A1 => n1335, A2 => n22307, ZN => n35756);
   U22210 : INV_X2 port map( I => n35757, ZN => n15248);
   U22216 : XOR2_X1 port map( A1 => n35758, A2 => n26171, Z => n26689);
   U22219 : XOR2_X1 port map( A1 => n26173, A2 => n36270, Z => n35758);
   U22235 : XOR2_X1 port map( A1 => n1323, A2 => n35211, Z => n35760);
   U22244 : INV_X2 port map( I => n35228, ZN => n27364);
   U22252 : NOR2_X1 port map( A1 => n859, A2 => n26936, ZN => n11339);
   U22255 : OAI21_X2 port map( A1 => n9951, A2 => n4833, B => n306, ZN => 
                           n28417);
   U22257 : NOR2_X2 port map( A1 => n5908, A2 => n35333, ZN => n25920);
   U22262 : NAND2_X1 port map( A1 => n35764, A2 => n35259, ZN => n6246);
   U22264 : XOR2_X1 port map( A1 => n9408, A2 => n9409, Z => n740);
   U22271 : XOR2_X1 port map( A1 => n35765, A2 => n34038, Z => n63);
   U22272 : XOR2_X1 port map( A1 => n29094, A2 => n31811, Z => n35765);
   U22273 : XNOR2_X1 port map( A1 => n18813, A2 => n11722, ZN => n36127);
   U22275 : XOR2_X1 port map( A1 => n2269, A2 => n29122, Z => n11722);
   U22280 : NOR2_X2 port map( A1 => n31453, A2 => n18590, ZN => n18241);
   U22290 : INV_X2 port map( I => n35769, ZN => n730);
   U22326 : OAI22_X2 port map( A1 => n11610, A2 => n5224, B1 => n5223, B2 => 
                           n20038, ZN => n20707);
   U22346 : NAND2_X1 port map( A1 => n28266, A2 => n38996, ZN => n36059);
   U22352 : NAND2_X2 port map( A1 => n10254, A2 => n28124, ZN => n27963);
   U22357 : AND2_X1 port map( A1 => n14075, A2 => n31899, Z => n14073);
   U22360 : NOR2_X2 port map( A1 => n6850, A2 => n5599, ZN => n35779);
   U22367 : XOR2_X1 port map( A1 => n25037, A2 => n9695, Z => n24838);
   U22380 : XOR2_X1 port map( A1 => n27809, A2 => n27529, Z => n27530);
   U22382 : NAND2_X2 port map( A1 => n11581, A2 => n35786, ZN => n17179);
   U22385 : NAND2_X2 port map( A1 => n17673, A2 => n36587, ZN => n19608);
   U22388 : NAND2_X2 port map( A1 => n31580, A2 => n12825, ZN => n25478);
   U22402 : OAI22_X2 port map( A1 => n15215, A2 => n34583, B1 => n20924, B2 => 
                           n541, ZN => n5597);
   U22403 : INV_X2 port map( I => n15261, ZN => n541);
   U22408 : NAND2_X2 port map( A1 => n33535, A2 => n14669, ZN => n35855);
   U22417 : XOR2_X1 port map( A1 => n7659, A2 => n19839, Z => n6363);
   U22420 : NOR2_X2 port map( A1 => n8503, A2 => n8504, ZN => n7659);
   U22430 : NOR2_X1 port map( A1 => n38202, A2 => n36838, ZN => n15695);
   U22433 : NOR2_X1 port map( A1 => n17194, A2 => n13371, ZN => n9366);
   U22445 : OAI21_X2 port map( A1 => n6503, A2 => n26471, B => n35794, ZN => 
                           n7757);
   U22449 : XOR2_X1 port map( A1 => n33498, A2 => n31020, Z => n1825);
   U22456 : OAI21_X2 port map( A1 => n23376, A2 => n23377, B => n23375, ZN => 
                           n33452);
   U22460 : NAND2_X2 port map( A1 => n36866, A2 => n21212, ZN => n16771);
   U22465 : NOR2_X2 port map( A1 => n35795, A2 => n8257, ZN => n27523);
   U22485 : XOR2_X1 port map( A1 => n35796, A2 => n26374, Z => n12012);
   U22499 : NAND2_X2 port map( A1 => n6332, A2 => n29644, ZN => n10868);
   U22504 : NAND2_X2 port map( A1 => n29443, A2 => n10870, ZN => n6332);
   U22533 : AOI21_X2 port map( A1 => n21306, A2 => n25771, B => n21305, ZN => 
                           n10965);
   U22534 : AND2_X1 port map( A1 => n9833, A2 => n25758, Z => n16890);
   U22536 : XOR2_X1 port map( A1 => n25215, A2 => n30973, Z => n36259);
   U22549 : NAND2_X2 port map( A1 => n3192, A2 => n36832, ZN => n28729);
   U22551 : NAND2_X2 port map( A1 => n14754, A2 => n21988, ZN => n22476);
   U22553 : NOR2_X1 port map( A1 => n3293, A2 => n21894, ZN => n21515);
   U22560 : NAND2_X2 port map( A1 => n35803, A2 => n13548, ZN => n17087);
   U22576 : XOR2_X1 port map( A1 => n26387, A2 => n26388, Z => n26474);
   U22590 : XNOR2_X1 port map( A1 => n5730, A2 => n25246, ZN => n36339);
   U22605 : XOR2_X1 port map( A1 => n35810, A2 => n22672, Z => n36291);
   U22607 : XOR2_X1 port map( A1 => n22582, A2 => n36290, Z => n22672);
   U22625 : OAI21_X2 port map( A1 => n13825, A2 => n13824, B => n28682, ZN => 
                           n13823);
   U22628 : INV_X2 port map( I => n35816, ZN => n37043);
   U22633 : XOR2_X1 port map( A1 => n30898, A2 => n784, Z => n35816);
   U22640 : AOI22_X2 port map( A1 => n35818, A2 => n34015, B1 => n8574, B2 => 
                           n21969, ZN => n2193);
   U22643 : OAI21_X2 port map( A1 => n21586, A2 => n119, B => n21584, ZN => 
                           n9876);
   U22659 : NAND2_X2 port map( A1 => n21128, A2 => n36876, ZN => n23900);
   U22660 : XOR2_X1 port map( A1 => n33470, A2 => n990, Z => n31138);
   U22667 : XOR2_X1 port map( A1 => n22592, A2 => n22514, Z => n20609);
   U22670 : NAND2_X1 port map( A1 => n22317, A2 => n36745, ZN => n7093);
   U22678 : AOI21_X2 port map( A1 => n28370, A2 => n28580, B => n16038, ZN => 
                           n35823);
   U22684 : OR2_X1 port map( A1 => n19477, A2 => n8798, Z => n35825);
   U22692 : NAND2_X2 port map( A1 => n35833, A2 => n36464, ZN => n22282);
   U22703 : NAND3_X2 port map( A1 => n33340, A2 => n33369, A3 => n12022, ZN => 
                           n35826);
   U22716 : BUF_X2 port map( I => n35867, Z => n35832);
   U22718 : XOR2_X1 port map( A1 => n17890, A2 => n19758, Z => n7763);
   U22729 : XOR2_X1 port map( A1 => n35834, A2 => n10863, Z => n11048);
   U22732 : INV_X2 port map( I => n35835, ZN => n12101);
   U22734 : OAI22_X1 port map( A1 => n13133, A2 => n13151, B1 => n35224, B2 => 
                           n14193, ZN => n31350);
   U22739 : XOR2_X1 port map( A1 => n35836, A2 => n12858, Z => n12856);
   U22741 : XOR2_X1 port map( A1 => n7250, A2 => n7247, Z => n8199);
   U22751 : NAND2_X1 port map( A1 => n307, A2 => n35837, ZN => n19784);
   U22753 : AOI22_X1 port map( A1 => n12369, A2 => n18873, B1 => n7303, B2 => 
                           n12148, ZN => n35837);
   U22754 : XOR2_X1 port map( A1 => n23948, A2 => n23949, Z => n17790);
   U22763 : XOR2_X1 port map( A1 => n7582, A2 => n34020, Z => n36756);
   U22779 : OAI22_X2 port map( A1 => n35841, A2 => n35840, B1 => n9362, B2 => 
                           n24290, ZN => n24707);
   U22783 : AOI21_X2 port map( A1 => n37118, A2 => n6668, B => n35843, ZN => 
                           n6875);
   U22784 : NOR3_X1 port map( A1 => n5772, A2 => n35228, A3 => n34001, ZN => 
                           n35843);
   U22785 : NAND2_X2 port map( A1 => n35844, A2 => n1437, ZN => n11006);
   U22791 : NOR2_X1 port map( A1 => n27895, A2 => n1445, ZN => n5470);
   U22793 : INV_X2 port map( I => n17755, ZN => n27895);
   U22823 : INV_X1 port map( I => n35847, ZN => n35846);
   U22824 : NAND2_X1 port map( A1 => n39488, A2 => n28238, ZN => n35847);
   U22825 : XOR2_X1 port map( A1 => n22528, A2 => n35848, Z => n494);
   U22827 : NAND2_X2 port map( A1 => n21831, A2 => n21832, ZN => n22528);
   U22833 : OAI21_X2 port map( A1 => n36607, A2 => n35849, B => n30163, ZN => 
                           n30173);
   U22847 : XOR2_X1 port map( A1 => n21036, A2 => n35853, Z => n35852);
   U22850 : OR2_X1 port map( A1 => n15218, A2 => n6581, Z => n6827);
   U22854 : AOI21_X2 port map( A1 => n3798, A2 => n3799, B => n33519, ZN => 
                           n35867);
   U22855 : XOR2_X1 port map( A1 => n35856, A2 => n24942, Z => n8277);
   U22856 : XOR2_X1 port map( A1 => n25284, A2 => n19683, Z => n35856);
   U22859 : XOR2_X1 port map( A1 => n35857, A2 => n2031, Z => n20866);
   U22861 : INV_X2 port map( I => n9900, ZN => n3602);
   U22862 : XOR2_X1 port map( A1 => n32959, A2 => n437, Z => n9900);
   U22864 : XOR2_X1 port map( A1 => n20485, A2 => n15471, Z => n20484);
   U22865 : BUF_X2 port map( I => n29699, Z => n35858);
   U22873 : NAND3_X2 port map( A1 => n16195, A2 => n18460, A3 => n24748, ZN => 
                           n25182);
   U22874 : XOR2_X1 port map( A1 => n11312, A2 => n11309, Z => n35859);
   U22876 : OAI22_X2 port map( A1 => n3618, A2 => n1990, B1 => n18699, B2 => 
                           n20266, ZN => n35860);
   U22894 : NOR2_X2 port map( A1 => n1028, A2 => n18110, ZN => n30421);
   U22897 : NAND2_X2 port map( A1 => n16473, A2 => n17338, ZN => n29034);
   U22914 : XOR2_X1 port map( A1 => n2284, A2 => n13551, Z => n12732);
   U22921 : CLKBUF_X4 port map( I => n21938, Z => n35883);
   U22932 : XOR2_X1 port map( A1 => n11999, A2 => n11998, Z => n861);
   U22935 : XOR2_X1 port map( A1 => n10971, A2 => n10970, Z => n7923);
   U22948 : NAND2_X1 port map( A1 => n2449, A2 => n18873, ZN => n2448);
   U22953 : NAND3_X2 port map( A1 => n9256, A2 => n10773, A3 => n19560, ZN => 
                           n25149);
   U22962 : OR2_X1 port map( A1 => n7303, A2 => n34534, Z => n29480);
   U22968 : XOR2_X1 port map( A1 => n22503, A2 => n21999, Z => n22002);
   U22982 : NAND3_X2 port map( A1 => n20751, A2 => n20750, A3 => n21612, ZN => 
                           n19373);
   U22991 : NOR2_X1 port map( A1 => n13927, A2 => n17378, ZN => n27995);
   U22993 : XOR2_X1 port map( A1 => n31777, A2 => n18060, Z => n13927);
   U22996 : INV_X2 port map( I => n35868, ZN => n20449);
   U23004 : NAND2_X2 port map( A1 => n27988, A2 => n27987, ZN => n28661);
   U23008 : OR2_X1 port map( A1 => n12049, A2 => n36117, Z => n32945);
   U23023 : XOR2_X1 port map( A1 => n12231, A2 => n28987, Z => n12215);
   U23024 : XOR2_X1 port map( A1 => n35871, A2 => n2159, Z => n5966);
   U23026 : XOR2_X1 port map( A1 => n35908, A2 => n8540, Z => n14217);
   U23040 : XOR2_X1 port map( A1 => n8654, A2 => n35874, Z => n4315);
   U23043 : XOR2_X1 port map( A1 => n28851, A2 => n31524, Z => n35874);
   U23051 : OAI22_X2 port map( A1 => n16288, A2 => n14769, B1 => n16287, B2 => 
                           n12927, ZN => n36214);
   U23069 : NAND2_X2 port map( A1 => n26067, A2 => n26066, ZN => n7602);
   U23075 : NAND3_X2 port map( A1 => n15614, A2 => n17219, A3 => n15613, ZN => 
                           n17440);
   U23077 : NAND2_X2 port map( A1 => n1048, A2 => n22184, ZN => n17793);
   U23078 : NAND2_X2 port map( A1 => n23522, A2 => n2273, ZN => n23525);
   U23087 : XOR2_X1 port map( A1 => n22723, A2 => n35879, Z => n35878);
   U23095 : NOR2_X2 port map( A1 => n11646, A2 => n9481, ZN => n35882);
   U23098 : AND2_X1 port map( A1 => n4880, A2 => n34786, Z => n30944);
   U23103 : NAND2_X2 port map( A1 => n17499, A2 => n22307, ZN => n36069);
   U23104 : XOR2_X1 port map( A1 => n22787, A2 => n22672, Z => n17277);
   U23106 : OR2_X1 port map( A1 => n730, A2 => n8069, Z => n8771);
   U23112 : NAND2_X2 port map( A1 => n23065, A2 => n23064, ZN => n23250);
   U23117 : NAND2_X2 port map( A1 => n6213, A2 => n4760, ZN => n23399);
   U23118 : NAND2_X2 port map( A1 => n35886, A2 => n15001, ZN => n25163);
   U23119 : BUF_X2 port map( I => n1254, Z => n35887);
   U23131 : XNOR2_X1 port map( A1 => n22622, A2 => n29223, ZN => n36605);
   U23140 : XOR2_X1 port map( A1 => n35889, A2 => n38226, Z => n184);
   U23146 : AOI22_X2 port map( A1 => n11878, A2 => n33489, B1 => n12169, B2 => 
                           n22367, ZN => n13704);
   U23159 : OR2_X1 port map( A1 => n20077, A2 => n15290, Z => n22783);
   U23160 : NAND2_X2 port map( A1 => n17132, A2 => n12327, ZN => n27398);
   U23163 : NAND2_X2 port map( A1 => n7010, A2 => n22730, ZN => n23637);
   U23190 : XOR2_X1 port map( A1 => n35996, A2 => n35894, Z => n14672);
   U23191 : XNOR2_X1 port map( A1 => n18807, A2 => n18279, ZN => n35970);
   U23197 : NAND2_X1 port map( A1 => n8495, A2 => n16039, ZN => n15115);
   U23199 : XOR2_X1 port map( A1 => n11901, A2 => Key(169), Z => n16039);
   U23200 : NAND2_X2 port map( A1 => n32796, A2 => n13042, ZN => n22838);
   U23220 : INV_X2 port map( I => n35896, ZN => n17594);
   U23223 : OR2_X1 port map( A1 => n7742, A2 => n26249, Z => n2226);
   U23228 : AND2_X1 port map( A1 => n30284, A2 => n14962, Z => n36929);
   U23241 : BUF_X2 port map( I => n27283, Z => n35904);
   U23248 : AOI21_X2 port map( A1 => n27107, A2 => n28052, B => n27962, ZN => 
                           n36029);
   U23250 : NAND2_X1 port map( A1 => n15224, A2 => n36791, ZN => n28733);
   U23275 : AND2_X1 port map( A1 => n30153, A2 => n20525, Z => n8717);
   U23278 : XOR2_X1 port map( A1 => n14425, A2 => n35909, Z => n5002);
   U23279 : XOR2_X1 port map( A1 => n15625, A2 => n29003, Z => n35909);
   U23280 : XOR2_X1 port map( A1 => n19047, A2 => n35910, Z => n30221);
   U23296 : XOR2_X1 port map( A1 => n17159, A2 => n28985, Z => n35910);
   U23297 : XOR2_X1 port map( A1 => n38171, A2 => n1553, Z => n25141);
   U23300 : INV_X2 port map( I => n38629, ZN => n35911);
   U23305 : NAND2_X2 port map( A1 => n14910, A2 => n14908, ZN => n20643);
   U23308 : NAND2_X1 port map( A1 => n17538, A2 => n17617, ZN => n17616);
   U23332 : XOR2_X1 port map( A1 => n26393, A2 => n26466, Z => n13244);
   U23348 : AOI21_X2 port map( A1 => n33849, A2 => n4686, B => n31678, ZN => 
                           n27045);
   U23354 : XOR2_X1 port map( A1 => n25268, A2 => n25162, Z => n10407);
   U23355 : XOR2_X1 port map( A1 => n13917, A2 => n25096, Z => n25162);
   U23361 : INV_X2 port map( I => n31107, ZN => n3662);
   U23365 : NAND2_X1 port map( A1 => n5988, A2 => n31107, ZN => n28235);
   U23389 : INV_X2 port map( I => n11970, ZN => n32017);
   U23404 : AOI21_X2 port map( A1 => n8328, A2 => n18150, B => n8325, ZN => 
                           n28398);
   U23428 : XOR2_X1 port map( A1 => n35923, A2 => n17759, Z => n26906);
   U23435 : NAND2_X2 port map( A1 => n1039, A2 => n30574, ZN => n23039);
   U23436 : OAI21_X2 port map( A1 => n33240, A2 => n2192, B => n35924, ZN => 
                           n14896);
   U23440 : NAND2_X2 port map( A1 => n2518, A2 => n576, ZN => n27637);
   U23459 : AOI22_X2 port map( A1 => n20827, A2 => n15031, B1 => n33285, B2 => 
                           n18005, ZN => n35926);
   U23479 : NAND3_X2 port map( A1 => n7483, A2 => n28154, A3 => n17818, ZN => 
                           n11296);
   U23490 : NAND2_X2 port map( A1 => n35928, A2 => n18378, ZN => n496);
   U23493 : OAI21_X2 port map( A1 => n18379, A2 => n18380, B => n27571, ZN => 
                           n35928);
   U23495 : NOR2_X1 port map( A1 => n5537, A2 => n26852, ZN => n19207);
   U23500 : NOR2_X1 port map( A1 => n5537, A2 => n20660, ZN => n11674);
   U23519 : XOR2_X1 port map( A1 => n25242, A2 => n25229, Z => n25313);
   U23549 : NAND3_X2 port map( A1 => n32182, A2 => n9663, A3 => n18150, ZN => 
                           n9575);
   U23566 : NAND2_X2 port map( A1 => n16235, A2 => n16488, ZN => n23939);
   U23567 : XOR2_X1 port map( A1 => n35941, A2 => n20486, Z => n15471);
   U23569 : XOR2_X1 port map( A1 => n37701, A2 => n35942, Z => n35941);
   U23577 : INV_X2 port map( I => n11937, ZN => n35942);
   U23591 : OAI21_X1 port map( A1 => n20623, A2 => n7357, B => n35943, ZN => 
                           n20148);
   U23600 : BUF_X2 port map( I => n26039, Z => n35944);
   U23623 : XOR2_X1 port map( A1 => n25841, A2 => n30469, Z => n857);
   U23624 : NOR2_X1 port map( A1 => n11678, A2 => n23391, ZN => n4859);
   U23627 : NAND2_X2 port map( A1 => n21634, A2 => n21633, ZN => n36397);
   U23659 : XOR2_X1 port map( A1 => n13550, A2 => n36390, Z => n36150);
   U23676 : XOR2_X1 port map( A1 => n20846, A2 => n20772, Z => n6049);
   U23697 : NAND2_X2 port map( A1 => n25659, A2 => n25658, ZN => n32095);
   U23698 : OAI22_X2 port map( A1 => n22314, A2 => n15004, B1 => n18675, B2 => 
                           n18674, ZN => n18087);
   U23699 : XOR2_X1 port map( A1 => n2042, A2 => n35957, Z => n36357);
   U23729 : INV_X2 port map( I => n2880, ZN => n15388);
   U23739 : XOR2_X1 port map( A1 => n3023, A2 => n3022, Z => n2880);
   U23741 : NAND2_X2 port map( A1 => n8070, A2 => n2148, ZN => n35962);
   U23745 : XOR2_X1 port map( A1 => n35964, A2 => n28630, Z => n28631);
   U23748 : XOR2_X1 port map( A1 => n29052, A2 => n19825, Z => n35964);
   U23762 : NOR3_X1 port map( A1 => n35966, A2 => n35965, A3 => n1406, ZN => 
                           n21196);
   U23763 : NOR2_X1 port map( A1 => n29310, A2 => n29384, ZN => n35965);
   U23770 : XOR2_X1 port map( A1 => n32135, A2 => n34345, Z => n22747);
   U23781 : NAND2_X2 port map( A1 => n37098, A2 => n19179, ZN => n26760);
   U23786 : NOR2_X1 port map( A1 => n14235, A2 => n35915, ZN => n10839);
   U23790 : NAND2_X2 port map( A1 => n13641, A2 => n13640, ZN => n14235);
   U23798 : XOR2_X1 port map( A1 => n35970, A2 => n23649, Z => n35969);
   U23803 : NOR2_X2 port map( A1 => n23942, A2 => n23941, ZN => n11081);
   U23805 : XOR2_X1 port map( A1 => n5629, A2 => n35971, Z => n734);
   U23808 : XOR2_X1 port map( A1 => n36128, A2 => n25025, Z => n35971);
   U23814 : AOI21_X2 port map( A1 => n35976, A2 => n35975, B => n7191, ZN => 
                           n18240);
   U23817 : NAND2_X1 port map( A1 => n7193, A2 => n7194, ZN => n35976);
   U23818 : BUF_X2 port map( I => n21111, Z => n35977);
   U23833 : NAND3_X1 port map( A1 => n27411, A2 => n27311, A3 => n997, ZN => 
                           n35978);
   U23854 : XOR2_X1 port map( A1 => n4646, A2 => n35983, Z => n12431);
   U23859 : XOR2_X1 port map( A1 => n37129, A2 => n35984, Z => n35983);
   U23861 : INV_X1 port map( I => n30122, ZN => n35984);
   U23879 : NAND2_X2 port map( A1 => n7805, A2 => n7808, ZN => n8402);
   U23925 : XOR2_X1 port map( A1 => n35993, A2 => n33357, Z => n384);
   U23927 : XOR2_X1 port map( A1 => n26545, A2 => n744, Z => n35993);
   U23930 : NOR2_X2 port map( A1 => n20670, A2 => n22153, ZN => n20335);
   U23931 : INV_X2 port map( I => n37643, ZN => n16686);
   U23933 : NAND2_X2 port map( A1 => n15502, A2 => n11671, ZN => n30881);
   U23935 : INV_X1 port map( I => n36815, ZN => n30436);
   U23938 : AND2_X1 port map( A1 => n36815, A2 => n36658, Z => n19215);
   U23950 : XOR2_X1 port map( A1 => n11215, A2 => n19991, Z => n9221);
   U23955 : NAND2_X2 port map( A1 => n22062, A2 => n32886, ZN => n32885);
   U23986 : NOR2_X2 port map( A1 => n9803, A2 => n10775, ZN => n26001);
   U23987 : XOR2_X1 port map( A1 => n26450, A2 => n26451, Z => n6681);
   U23996 : OR2_X1 port map( A1 => n28389, A2 => n18960, Z => n11911);
   U23999 : AOI22_X2 port map( A1 => n22083, A2 => n23114, B1 => n23115, B2 => 
                           n8569, ZN => n36001);
   U24015 : NOR2_X2 port map( A1 => n36004, A2 => n8265, ZN => n32002);
   U24020 : NOR2_X1 port map( A1 => n2969, A2 => n36801, ZN => n2967);
   U24029 : XOR2_X1 port map( A1 => n26448, A2 => n37380, Z => n659);
   U24040 : NAND2_X2 port map( A1 => n20551, A2 => n12568, ZN => n22645);
   U24041 : XOR2_X1 port map( A1 => n36013, A2 => n19937, Z => Ciphertext(164))
                           ;
   U24055 : NOR3_X1 port map( A1 => n21248, A2 => n27508, A3 => n31287, ZN => 
                           n27187);
   U24060 : INV_X4 port map( I => n36532, ZN => n15677);
   U24062 : NAND2_X2 port map( A1 => n5454, A2 => n5452, ZN => n36532);
   U24067 : XOR2_X1 port map( A1 => n19096, A2 => n2318, Z => n2317);
   U24074 : OAI21_X2 port map( A1 => n36020, A2 => n20105, B => n911, ZN => 
                           n18349);
   U24119 : INV_X2 port map( I => n36024, ZN => n11060);
   U24120 : XOR2_X1 port map( A1 => n11061, A2 => n11062, Z => n36024);
   U24124 : XOR2_X1 port map( A1 => n22543, A2 => n18751, Z => n1947);
   U24140 : NOR2_X1 port map( A1 => n17931, A2 => n23354, ZN => n36026);
   U24145 : NAND3_X1 port map( A1 => n31192, A2 => n2888, A3 => n3575, ZN => 
                           n2889);
   U24149 : NOR2_X1 port map( A1 => n36794, A2 => n24896, ZN => n25584);
   U24158 : XOR2_X1 port map( A1 => n36030, A2 => n36205, Z => n14481);
   U24159 : XOR2_X1 port map( A1 => n25265, A2 => n14672, Z => n36030);
   U24172 : INV_X2 port map( I => n25283, ZN => n30318);
   U24177 : NAND2_X2 port map( A1 => n24546, A2 => n4694, ZN => n25283);
   U24180 : NAND2_X1 port map( A1 => n24146, A2 => n1602, ZN => n8501);
   U24206 : NAND3_X2 port map( A1 => n29767, A2 => n31059, A3 => n31517, ZN => 
                           n29792);
   U24208 : NAND2_X2 port map( A1 => n20028, A2 => n24439, ZN => n36075);
   U24211 : XOR2_X1 port map( A1 => n11753, A2 => n29528, Z => n11207);
   U24213 : XOR2_X1 port map( A1 => n36034, A2 => n5103, Z => n14411);
   U24215 : OAI21_X2 port map( A1 => n33380, A2 => n20870, B => n36036, ZN => 
                           n27781);
   U24223 : NAND2_X1 port map( A1 => n21461, A2 => n21868, ZN => n3564);
   U24229 : XOR2_X1 port map( A1 => n2068, A2 => n2067, Z => n2066);
   U24238 : XOR2_X1 port map( A1 => n22592, A2 => n36038, Z => n22596);
   U24260 : NAND2_X2 port map( A1 => n32337, A2 => n11683, ZN => n15871);
   U24274 : XOR2_X1 port map( A1 => n32646, A2 => n36040, Z => n2352);
   U24277 : NAND2_X1 port map( A1 => n28807, A2 => n19759, ZN => n28289);
   U24280 : XOR2_X1 port map( A1 => n27598, A2 => n32686, Z => n36041);
   U24282 : NAND2_X2 port map( A1 => n5777, A2 => n5776, ZN => n9824);
   U24301 : INV_X2 port map( I => n36044, ZN => n1589);
   U24304 : XNOR2_X1 port map( A1 => n36646, A2 => n2398, ZN => n36044);
   U24309 : NOR2_X2 port map( A1 => n36046, A2 => n4775, ZN => n9999);
   U24313 : XOR2_X1 port map( A1 => n33645, A2 => n29649, Z => n17798);
   U24325 : NOR2_X1 port map( A1 => n38609, A2 => n12235, ZN => n18752);
   U24335 : XOR2_X1 port map( A1 => n26208, A2 => n659, Z => n12412);
   U24364 : OAI21_X1 port map( A1 => n38156, A2 => n16889, B => n36051, ZN => 
                           n9559);
   U24367 : OAI21_X1 port map( A1 => n1208, A2 => n39235, B => n17770, ZN => 
                           n9684);
   U24374 : NAND2_X2 port map( A1 => n36053, A2 => n25339, ZN => n26063);
   U24385 : OAI21_X1 port map( A1 => n566, A2 => n33968, B => n29719, ZN => 
                           n16630);
   U24389 : NAND2_X2 port map( A1 => n7251, A2 => n36935, ZN => n28525);
   U24398 : XOR2_X1 port map( A1 => n3110, A2 => n25182, Z => n25312);
   U24411 : NOR2_X2 port map( A1 => n21709, A2 => n36055, ZN => n22092);
   U24413 : AOI21_X1 port map( A1 => n21706, A2 => n21707, B => n2045, ZN => 
                           n36055);
   U24416 : NOR2_X1 port map( A1 => n5709, A2 => n11622, ZN => n30377);
   U24429 : XOR2_X1 port map( A1 => n2935, A2 => n22453, Z => n36057);
   U24434 : OR2_X1 port map( A1 => n29756, A2 => n29754, Z => n33607);
   U24443 : XOR2_X1 port map( A1 => Plaintext(145), A2 => Key(145), Z => n36062
                           );
   U24445 : NAND2_X2 port map( A1 => n15868, A2 => n17869, ZN => n17335);
   U24449 : INV_X2 port map( I => n36063, ZN => n7240);
   U24450 : INV_X2 port map( I => n36064, ZN => n32775);
   U24466 : XOR2_X1 port map( A1 => n26279, A2 => n19808, Z => n13931);
   U24467 : BUF_X2 port map( I => n23899, Z => n36065);
   U24470 : XOR2_X1 port map( A1 => n36066, A2 => n6764, Z => n24285);
   U24483 : XOR2_X1 port map( A1 => n22597, A2 => n33177, Z => n12863);
   U24486 : XOR2_X1 port map( A1 => n36068, A2 => n24016, Z => n3454);
   U24492 : XOR2_X1 port map( A1 => n23667, A2 => n11739, Z => n24016);
   U24499 : AOI21_X1 port map( A1 => n36069, A2 => n1335, B => n17989, ZN => 
                           n4126);
   U24509 : XOR2_X1 port map( A1 => n22574, A2 => n6047, Z => n30661);
   U24552 : AOI21_X2 port map( A1 => n4384, A2 => n1547, B => n36133, ZN => 
                           n36071);
   U24557 : OAI21_X2 port map( A1 => n4456, A2 => n27946, B => n36072, ZN => 
                           n28651);
   U24564 : XOR2_X1 port map( A1 => n36074, A2 => n873, Z => n9373);
   U24566 : XOR2_X1 port map( A1 => n27605, A2 => n32021, Z => n36074);
   U24584 : BUF_X2 port map( I => n10907, Z => n36076);
   U24586 : XOR2_X1 port map( A1 => n36077, A2 => n6963, Z => n26177);
   U24587 : XOR2_X1 port map( A1 => n26554, A2 => n26245, Z => n26488);
   U24591 : NAND2_X2 port map( A1 => n4431, A2 => n4430, ZN => n26245);
   U24599 : XOR2_X1 port map( A1 => n26161, A2 => n29269, Z => n9932);
   U24618 : NAND2_X2 port map( A1 => n3013, A2 => n25799, ZN => n3434);
   U24619 : XOR2_X1 port map( A1 => n23997, A2 => n36079, Z => n19960);
   U24624 : OAI22_X2 port map( A1 => n36080, A2 => n1220, B1 => n2998, B2 => 
                           n10946, ZN => n12341);
   U24625 : XOR2_X1 port map( A1 => n36970, A2 => n36081, Z => n33479);
   U24627 : XOR2_X1 port map( A1 => n17363, A2 => n8780, Z => n36081);
   U24634 : XOR2_X1 port map( A1 => n15592, A2 => n19797, Z => n1886);
   U24635 : XOR2_X1 port map( A1 => n22670, A2 => n36290, Z => n20412);
   U24640 : NAND2_X2 port map( A1 => n21263, A2 => n21260, ZN => n36290);
   U24646 : INV_X2 port map( I => n6947, ZN => n22326);
   U24656 : OAI22_X2 port map( A1 => n439, A2 => n440, B1 => n13557, B2 => 
                           n13556, ZN => n6947);
   U24657 : INV_X4 port map( I => n7221, ZN => n8082);
   U24663 : NAND2_X2 port map( A1 => n6243, A2 => n6244, ZN => n7221);
   U24669 : XOR2_X1 port map( A1 => n23804, A2 => n6289, Z => n36087);
   U24700 : NAND2_X2 port map( A1 => n22059, A2 => n22100, ZN => n36092);
   U24708 : NAND2_X2 port map( A1 => n12542, A2 => n28492, ZN => n29252);
   U24720 : AOI22_X2 port map( A1 => n9726, A2 => n6775, B1 => n1475, B2 => 
                           n27130, ZN => n27632);
   U24729 : NAND2_X1 port map( A1 => n2339, A2 => n8155, ZN => n36097);
   U24737 : NAND2_X1 port map( A1 => n19285, A2 => n4748, ZN => n36098);
   U24741 : NAND2_X1 port map( A1 => n36099, A2 => n2678, ZN => n33517);
   U24752 : INV_X2 port map( I => n36104, ZN => n30317);
   U24764 : XOR2_X1 port map( A1 => n26279, A2 => n26404, Z => n15530);
   U24766 : NAND2_X2 port map( A1 => n15870, A2 => n15869, ZN => n26404);
   U24775 : NOR2_X2 port map( A1 => n6421, A2 => n6684, ZN => n3309);
   U24778 : INV_X2 port map( I => n23310, ZN => n6421);
   U24786 : NAND2_X2 port map( A1 => n36444, A2 => n2088, ZN => n7693);
   U24802 : NAND3_X2 port map( A1 => n2587, A2 => n2586, A3 => n14597, ZN => 
                           n15346);
   U24803 : NAND2_X2 port map( A1 => n36109, A2 => n36108, ZN => n17732);
   U24806 : INV_X1 port map( I => n36775, ZN => n36108);
   U24810 : XOR2_X1 port map( A1 => n9762, A2 => n36111, Z => n10655);
   U24811 : XOR2_X1 port map( A1 => n16082, A2 => n34161, Z => n36111);
   U24824 : INV_X2 port map( I => n36113, ZN => n2597);
   U24833 : XOR2_X1 port map( A1 => n27837, A2 => n13878, Z => n36114);
   U24835 : OAI22_X2 port map( A1 => n33206, A2 => n33394, B1 => n37083, B2 => 
                           n30196, ZN => n32925);
   U24847 : INV_X2 port map( I => n36117, ZN => n37060);
   U24848 : XOR2_X1 port map( A1 => n6852, A2 => n6855, Z => n36117);
   U24859 : XOR2_X1 port map( A1 => n38514, A2 => n18004, Z => n5119);
   U24871 : XOR2_X1 port map( A1 => n9390, A2 => n36119, Z => n6593);
   U24872 : XOR2_X1 port map( A1 => n31872, A2 => n7990, Z => n36119);
   U24874 : AOI21_X2 port map( A1 => n27232, A2 => n945, B => n36120, ZN => 
                           n20823);
   U24882 : XOR2_X1 port map( A1 => n36123, A2 => n29017, Z => Ciphertext(173))
                           ;
   U24890 : AOI22_X1 port map( A1 => n29015, A2 => n30131, B1 => n29016, B2 => 
                           n3896, ZN => n36123);
   U24892 : XOR2_X1 port map( A1 => n27842, A2 => n7549, Z => n21087);
   U24900 : NAND3_X2 port map( A1 => n20434, A2 => n36126, A3 => n36125, ZN => 
                           n20437);
   U24912 : XOR2_X1 port map( A1 => n5750, A2 => n27855, Z => n10782);
   U24926 : AND2_X2 port map( A1 => n5899, A2 => n5966, Z => n4915);
   U24932 : XOR2_X1 port map( A1 => n13076, A2 => n18395, Z => n36128);
   U24944 : OAI22_X2 port map( A1 => n8968, A2 => n24866, B1 => n7970, B2 => 
                           n8314, ZN => n7967);
   U24947 : OAI21_X1 port map( A1 => n33976, A2 => n36135, B => n25328, ZN => 
                           n36134);
   U24948 : INV_X2 port map( I => n36136, ZN => n4803);
   U24955 : NAND2_X2 port map( A1 => n7781, A2 => n8248, ZN => n16216);
   U24961 : NOR2_X2 port map( A1 => n5734, A2 => n36139, ZN => n4497);
   U24964 : XOR2_X1 port map( A1 => n30913, A2 => n26499, Z => n13673);
   U24972 : OAI21_X2 port map( A1 => n5392, A2 => n5391, B => n36140, ZN => 
                           n5777);
   U24973 : INV_X2 port map( I => n36141, ZN => n36140);
   U24981 : OAI21_X2 port map( A1 => n19587, A2 => n5132, B => n1155, ZN => 
                           n36141);
   U24984 : OAI21_X1 port map( A1 => n18910, A2 => n12543, B => n36144, ZN => 
                           n13028);
   U25004 : NOR3_X1 port map( A1 => n1427, A2 => n28611, A3 => n8787, ZN => 
                           n5927);
   U25008 : XOR2_X1 port map( A1 => n6751, A2 => n6753, Z => n28127);
   U25009 : BUF_X2 port map( I => n9616, Z => n36151);
   U25014 : NAND2_X2 port map( A1 => n20464, A2 => n20463, ZN => n25345);
   U25016 : OAI21_X1 port map( A1 => n19557, A2 => n27337, B => n36152, ZN => 
                           n27135);
   U25043 : XOR2_X1 port map( A1 => n15844, A2 => n34162, Z => n32842);
   U25054 : NAND2_X2 port map( A1 => n29491, A2 => n1179, ZN => n12428);
   U25061 : OR2_X1 port map( A1 => n17072, A2 => n13699, Z => n32962);
   U25062 : NOR2_X2 port map( A1 => n33668, A2 => n16124, ZN => n17072);
   U25068 : NAND2_X2 port map( A1 => n28433, A2 => n39423, ZN => n28460);
   U25083 : OAI21_X2 port map( A1 => n36164, A2 => n26799, B => n10203, ZN => 
                           n7973);
   U25094 : OAI21_X2 port map( A1 => n14409, A2 => n14439, B => n22804, ZN => 
                           n12960);
   U25107 : INV_X2 port map( I => n36160, ZN => n37045);
   U25108 : XOR2_X1 port map( A1 => n5937, A2 => n5936, Z => n36160);
   U25115 : OAI21_X2 port map( A1 => n36816, A2 => n13460, B => n1113, ZN => 
                           n13320);
   U25116 : NAND2_X2 port map( A1 => n5896, A2 => n24492, ZN => n24763);
   U25118 : NAND3_X2 port map( A1 => n36163, A2 => n25070, A3 => n25067, ZN => 
                           n31242);
   U25121 : XOR2_X1 port map( A1 => n8972, A2 => n30126, Z => n25809);
   U25134 : NAND2_X1 port map( A1 => n36524, A2 => n11150, ZN => n30381);
   U25140 : XOR2_X1 port map( A1 => n36168, A2 => n34239, Z => Ciphertext(88));
   U25147 : INV_X2 port map( I => n18032, ZN => n25965);
   U25157 : NAND2_X2 port map( A1 => n30988, A2 => n36612, ZN => n18032);
   U25168 : NAND2_X2 port map( A1 => n36170, A2 => n29173, ZN => n13559);
   U25178 : AND2_X2 port map( A1 => n30597, A2 => n36931, Z => n26727);
   U25183 : INV_X1 port map( I => n29206, ZN => n36171);
   U25189 : NAND2_X2 port map( A1 => n1782, A2 => n1785, ZN => n4302);
   U25207 : NAND3_X1 port map( A1 => n29922, A2 => n31570, A3 => n3860, ZN => 
                           n8583);
   U25230 : NOR2_X2 port map( A1 => n15644, A2 => n36172, ZN => n33512);
   U25233 : INV_X2 port map( I => n36173, ZN => n833);
   U25234 : XOR2_X1 port map( A1 => n15938, A2 => n15937, Z => n36173);
   U25257 : AOI21_X2 port map( A1 => n26834, A2 => n26835, B => n38852, ZN => 
                           n36175);
   U25277 : BUF_X4 port map( I => n23354, Z => n36564);
   U25285 : NOR2_X1 port map( A1 => n22171, A2 => n36176, ZN => n1840);
   U25302 : XOR2_X1 port map( A1 => n13235, A2 => n22638, Z => n4560);
   U25304 : XOR2_X1 port map( A1 => n19725, A2 => n24982, Z => n25245);
   U25307 : NAND2_X2 port map( A1 => n11906, A2 => n24823, ZN => n24982);
   U25308 : NAND2_X2 port map( A1 => n9824, A2 => n4179, ZN => n33581);
   U25314 : NAND2_X1 port map( A1 => n36180, A2 => n24819, ZN => n8648);
   U25321 : XOR2_X1 port map( A1 => n23740, A2 => n36181, Z => n6156);
   U25323 : XOR2_X1 port map( A1 => n6227, A2 => n20317, Z => n36181);
   U25324 : NAND2_X1 port map( A1 => n2487, A2 => n36182, ZN => n2485);
   U25330 : BUF_X2 port map( I => n32205, Z => n36183);
   U25331 : NAND2_X1 port map( A1 => n17691, A2 => n17692, ZN => n36184);
   U25346 : XOR2_X1 port map( A1 => n24436, A2 => n21174, Z => n36205);
   U25349 : INV_X2 port map( I => n19979, ZN => n5896);
   U25350 : INV_X2 port map( I => n24492, ZN => n36186);
   U25384 : NAND2_X2 port map( A1 => n16964, A2 => n385, ZN => n18910);
   U25387 : NAND2_X2 port map( A1 => n28290, A2 => n877, ZN => n27896);
   U25394 : XOR2_X1 port map( A1 => n22736, A2 => n22737, Z => n36190);
   U25405 : NAND2_X2 port map( A1 => n33844, A2 => n36193, ZN => n29437);
   U25413 : NAND2_X2 port map( A1 => n36194, A2 => n25508, ZN => n20851);
   U25415 : OAI21_X2 port map( A1 => n10850, A2 => n38825, B => n33327, ZN => 
                           n36194);
   U25417 : OAI21_X1 port map( A1 => n28750, A2 => n28745, B => n33283, ZN => 
                           n28523);
   U25451 : AOI21_X2 port map( A1 => n22945, A2 => n19488, B => n17083, ZN => 
                           n23390);
   U25454 : XOR2_X1 port map( A1 => n36195, A2 => n1765, Z => n13587);
   U25474 : NAND2_X2 port map( A1 => n12466, A2 => n3097, ZN => n36588);
   U25475 : NAND2_X1 port map( A1 => n36199, A2 => n1598, ZN => n23816);
   U25481 : OAI21_X1 port map( A1 => n24294, A2 => n8824, B => n33939, ZN => 
                           n36199);
   U25490 : AOI22_X1 port map( A1 => n36201, A2 => n626, B1 => n10342, B2 => 
                           n11673, ZN => n31437);
   U25514 : OAI21_X1 port map( A1 => n1606, A2 => n18329, B => n3398, ZN => 
                           n36201);
   U25523 : INV_X2 port map( I => n37014, ZN => n1135);
   U25531 : XOR2_X1 port map( A1 => n36204, A2 => n15932, Z => n30839);
   U25542 : XOR2_X1 port map( A1 => n386, A2 => n19774, Z => n36204);
   U25547 : XOR2_X1 port map( A1 => n16021, A2 => n23790, Z => n36206);
   U25548 : XNOR2_X1 port map( A1 => n4278, A2 => n4277, ZN => n36698);
   U25554 : NAND2_X2 port map( A1 => n11006, A2 => n11005, ZN => n19631);
   U25558 : NAND2_X2 port map( A1 => n25261, A2 => n37052, ZN => n25725);
   U25560 : XOR2_X1 port map( A1 => n1463, A2 => n12999, Z => n36211);
   U25565 : NOR2_X2 port map( A1 => n34121, A2 => n11108, ZN => n36212);
   U25566 : XOR2_X1 port map( A1 => n22490, A2 => n13478, Z => n13477);
   U25568 : NOR2_X1 port map( A1 => n35260, A2 => n9815, ZN => n37049);
   U25571 : NAND2_X1 port map( A1 => n31199, A2 => n23380, ZN => n14974);
   U25572 : NAND2_X2 port map( A1 => n454, A2 => n10670, ZN => n30097);
   U25583 : NAND2_X2 port map( A1 => n30350, A2 => n36936, ZN => n5028);
   U25588 : XOR2_X1 port map( A1 => n25173, A2 => n24921, Z => n11061);
   U25596 : OR2_X1 port map( A1 => n36471, A2 => n35901, Z => n31625);
   U25619 : INV_X2 port map( I => n17353, ZN => n36216);
   U25636 : BUF_X2 port map( I => n14231, Z => n36218);
   U25649 : XNOR2_X1 port map( A1 => n28896, A2 => n32608, ZN => n32465);
   U25676 : XOR2_X1 port map( A1 => n8904, A2 => n35970, Z => n18404);
   U25688 : INV_X2 port map( I => n14015, ZN => n6908);
   U25690 : NAND3_X2 port map( A1 => n30715, A2 => n12565, A3 => n12566, ZN => 
                           n14015);
   U25691 : NAND2_X2 port map( A1 => n17107, A2 => n2114, ZN => n27767);
   U25701 : XOR2_X1 port map( A1 => n8605, A2 => n25040, Z => n17623);
   U25704 : XOR2_X1 port map( A1 => n28796, A2 => n28795, Z => n19224);
   U25707 : XOR2_X1 port map( A1 => n26513, A2 => n844, Z => n5177);
   U25709 : INV_X2 port map( I => n14751, ZN => n24963);
   U25717 : NOR2_X2 port map( A1 => n32347, A2 => n32348, ZN => n32205);
   U25731 : OR3_X2 port map( A1 => n32775, A2 => n25487, A3 => n10938, Z => 
                           n14656);
   U25732 : OR2_X1 port map( A1 => n15865, A2 => n8193, Z => n12564);
   U25745 : XOR2_X1 port map( A1 => n26207, A2 => n1507, Z => n26393);
   U25760 : BUF_X4 port map( I => n30504, Z => n36340);
   U25766 : NOR2_X2 port map( A1 => n21319, A2 => n9846, ZN => n36229);
   U25768 : XOR2_X1 port map( A1 => n36231, A2 => n2120, Z => n2117);
   U25771 : XOR2_X1 port map( A1 => n39209, A2 => n6561, Z => n36233);
   U25775 : XOR2_X1 port map( A1 => n29095, A2 => n29145, Z => n29255);
   U25782 : XOR2_X1 port map( A1 => n7337, A2 => n22714, Z => n22719);
   U25786 : NAND2_X2 port map( A1 => n28091, A2 => n36236, ZN => n28463);
   U25794 : XOR2_X1 port map( A1 => n7055, A2 => n36238, Z => n33315);
   U25799 : INV_X1 port map( I => n22715, ZN => n36238);
   U25800 : NAND2_X2 port map( A1 => n22090, A2 => n7490, ZN => n22715);
   U25806 : NOR2_X1 port map( A1 => n14704, A2 => n30280, ZN => n11760);
   U25814 : NAND2_X2 port map( A1 => n16034, A2 => n20019, ZN => n36320);
   U25840 : XOR2_X1 port map( A1 => n36240, A2 => n36239, Z => n15386);
   U25844 : XOR2_X1 port map( A1 => n8586, A2 => n11050, Z => n36240);
   U25850 : XOR2_X1 port map( A1 => n22710, A2 => n22464, Z => n22667);
   U25855 : XOR2_X1 port map( A1 => n37957, A2 => n23710, Z => n23662);
   U25858 : XOR2_X1 port map( A1 => n31410, A2 => n30756, Z => n31305);
   U25860 : NAND2_X2 port map( A1 => n8305, A2 => n34150, ZN => n260);
   U25864 : BUF_X2 port map( I => n9422, Z => n36245);
   U25865 : NAND2_X1 port map( A1 => n32695, A2 => n20133, ZN => n36250);
   U25870 : INV_X2 port map( I => n36253, ZN => n37057);
   U25875 : INV_X2 port map( I => n38165, ZN => n36254);
   U25883 : INV_X2 port map( I => n36257, ZN => n26763);
   U25884 : XOR2_X1 port map( A1 => n32734, A2 => n36258, Z => n2895);
   U25889 : XOR2_X1 port map( A1 => n25103, A2 => n36259, Z => n36258);
   U25896 : BUF_X4 port map( I => n34603, Z => n36263);
   U25897 : NAND3_X2 port map( A1 => n23069, A2 => n6000, A3 => n11366, ZN => 
                           n19005);
   U25901 : XOR2_X1 port map( A1 => n5721, A2 => n5722, Z => n252);
   U25948 : INV_X2 port map( I => n8182, ZN => n15164);
   U25951 : XOR2_X1 port map( A1 => n27697, A2 => n36260, Z => n8182);
   U25952 : XOR2_X1 port map( A1 => n19717, A2 => n36265, Z => n10239);
   U25957 : NAND2_X2 port map( A1 => n22381, A2 => n22380, ZN => n19717);
   U25959 : NAND2_X2 port map( A1 => n30780, A2 => n36266, ZN => n28677);
   U25965 : NAND2_X1 port map( A1 => n1086, A2 => n27589, ZN => n12263);
   U25980 : NAND2_X2 port map( A1 => n3264, A2 => n9609, ZN => n11937);
   U25990 : XOR2_X1 port map( A1 => n25141, A2 => n15779, Z => n21207);
   U26016 : XOR2_X1 port map( A1 => n26169, A2 => n9776, Z => n36270);
   U26025 : INV_X2 port map( I => n28514, ZN => n1881);
   U26034 : NAND2_X2 port map( A1 => n32759, A2 => n1882, ZN => n28514);
   U26035 : OAI21_X2 port map( A1 => n26, A2 => n12793, B => n37011, ZN => 
                           n36271);
   U26053 : NAND2_X2 port map( A1 => n27192, A2 => n31421, ZN => n19355);
   U26056 : AOI22_X2 port map( A1 => n36273, A2 => n15319, B1 => n32297, B2 => 
                           n14558, ZN => n13624);
   U26078 : INV_X4 port map( I => n17424, ZN => n36275);
   U26085 : XOR2_X1 port map( A1 => n3488, A2 => n11722, Z => n16647);
   U26102 : OAI21_X2 port map( A1 => n33926, A2 => n23328, B => n36279, ZN => 
                           n18279);
   U26106 : NAND2_X1 port map( A1 => n1763, A2 => n531, ZN => n16954);
   U26112 : NAND3_X1 port map( A1 => n12564, A2 => n19426, A3 => n38839, ZN => 
                           n11521);
   U26117 : INV_X2 port map( I => n36283, ZN => n8413);
   U26118 : XOR2_X1 port map( A1 => n2594, A2 => n33653, Z => n36284);
   U26120 : AOI22_X2 port map( A1 => n8686, A2 => n26179, B1 => n924, B2 => 
                           n5746, ZN => n5745);
   U26127 : XOR2_X1 port map( A1 => n36286, A2 => n20874, Z => n23074);
   U26132 : XOR2_X1 port map( A1 => n30444, A2 => n22387, Z => n36286);
   U26143 : NAND2_X2 port map( A1 => n37103, A2 => n1092, ZN => n26817);
   U26152 : OR2_X2 port map( A1 => n19250, A2 => n36655, Z => n36523);
   U26155 : XOR2_X1 port map( A1 => n36289, A2 => n27732, Z => n10002);
   U26159 : XOR2_X1 port map( A1 => n7651, A2 => n7549, Z => n36289);
   U26176 : AOI22_X1 port map( A1 => n12450, A2 => n38420, B1 => n1404, B2 => 
                           n31667, ZN => n2410);
   U26177 : XOR2_X1 port map( A1 => n36291, A2 => n20502, Z => n4633);
   U26185 : NAND2_X1 port map( A1 => n17261, A2 => n187, ZN => n36446);
   U26199 : BUF_X2 port map( I => n33440, Z => n36293);
   U26212 : XOR2_X1 port map( A1 => n8554, A2 => n8553, Z => n9775);
   U26220 : NAND2_X2 port map( A1 => n10650, A2 => n10649, ZN => n17074);
   U26229 : OAI22_X2 port map( A1 => n18028, A2 => n20476, B1 => n32164, B2 => 
                           n14450, ZN => n17923);
   U26236 : XOR2_X1 port map( A1 => n26208, A2 => n32386, Z => n26211);
   U26237 : NOR2_X2 port map( A1 => n36297, A2 => n21614, ZN => n9736);
   U26238 : INV_X2 port map( I => n15113, ZN => n32759);
   U26243 : NAND2_X2 port map( A1 => n13458, A2 => n13455, ZN => n15113);
   U26244 : XOR2_X1 port map( A1 => n1794, A2 => n1792, Z => n20026);
   U26246 : NAND3_X2 port map( A1 => n20999, A2 => n22284, A3 => n21000, ZN => 
                           n22464);
   U26248 : XOR2_X1 port map( A1 => n33179, A2 => n23732, Z => n18922);
   U26255 : INV_X2 port map( I => n12633, ZN => n1122);
   U26256 : NAND2_X2 port map( A1 => n16446, A2 => n16450, ZN => n12633);
   U26277 : XOR2_X1 port map( A1 => n17137, A2 => n17136, Z => n17984);
   U26278 : NAND3_X2 port map( A1 => n14444, A2 => n31820, A3 => n14656, ZN => 
                           n18176);
   U26288 : XOR2_X1 port map( A1 => n22466, A2 => n18189, Z => n10107);
   U26298 : NAND2_X2 port map( A1 => n36300, A2 => n18426, ZN => n26582);
   U26299 : NAND2_X2 port map( A1 => n23242, A2 => n21130, ZN => n36876);
   U26301 : XOR2_X1 port map( A1 => n25312, A2 => n25074, Z => n15937);
   U26304 : XOR2_X1 port map( A1 => n37038, A2 => n24935, Z => n25074);
   U26316 : XOR2_X1 port map( A1 => n13634, A2 => n15625, Z => n21259);
   U26320 : NAND2_X2 port map( A1 => n14593, A2 => n12817, ZN => n15625);
   U26323 : NAND3_X2 port map( A1 => n10795, A2 => n10796, A3 => n21255, ZN => 
                           n27252);
   U26326 : XOR2_X1 port map( A1 => n7256, A2 => n4009, Z => n882);
   U26327 : OAI22_X2 port map( A1 => n14129, A2 => n36263, B1 => n6514, B2 => 
                           n23594, ZN => n11098);
   U26339 : NOR2_X2 port map( A1 => n37237, A2 => n611, ZN => n36302);
   U26359 : XOR2_X1 port map( A1 => n17344, A2 => n1971, Z => n36305);
   U26389 : NAND2_X2 port map( A1 => n30728, A2 => n4916, ZN => n4377);
   U26390 : OAI21_X2 port map( A1 => n8392, A2 => n930, B => n36308, ZN => 
                           n18631);
   U26391 : NAND3_X2 port map( A1 => n7258, A2 => n2534, A3 => n9959, ZN => 
                           n36308);
   U26395 : NOR2_X1 port map( A1 => n36310, A2 => n36309, ZN => n20187);
   U26396 : NOR2_X1 port map( A1 => n19813, A2 => n6448, ZN => n36310);
   U26397 : XOR2_X1 port map( A1 => n25141, A2 => n20409, Z => n15265);
   U26412 : XOR2_X1 port map( A1 => n22604, A2 => n6893, Z => n22755);
   U26416 : XOR2_X1 port map( A1 => n10112, A2 => n36311, Z => n10111);
   U26418 : XOR2_X1 port map( A1 => n26468, A2 => n34157, Z => n36311);
   U26428 : OAI21_X1 port map( A1 => n36490, A2 => n13998, B => n21555, ZN => 
                           n7414);
   U26447 : INV_X1 port map( I => n5750, ZN => n36317);
   U26452 : XOR2_X1 port map( A1 => n26370, A2 => n26486, Z => n12114);
   U26461 : OAI22_X1 port map( A1 => n34156, A2 => n9529, B1 => n26063, B2 => 
                           n19793, ZN => n9086);
   U26473 : NAND2_X2 port map( A1 => n36322, A2 => n9209, ZN => n19670);
   U26479 : OAI22_X1 port map( A1 => n17985, A2 => n20671, B1 => n17422, B2 => 
                           n11910, ZN => n17420);
   U26489 : XOR2_X1 port map( A1 => n3956, A2 => n36326, Z => n3134);
   U26493 : XOR2_X1 port map( A1 => n26529, A2 => n745, Z => n36326);
   U26498 : XOR2_X1 port map( A1 => n12818, A2 => n36327, Z => n3663);
   U26506 : XOR2_X1 port map( A1 => n22772, A2 => n37042, Z => n36327);
   U26507 : NOR2_X1 port map( A1 => n14011, A2 => n35232, ZN => n43);
   U26513 : XOR2_X1 port map( A1 => n26279, A2 => n32003, Z => n25735);
   U26533 : XOR2_X1 port map( A1 => n15222, A2 => n27816, Z => n36329);
   U26539 : OR2_X1 port map( A1 => n19203, A2 => n27383, Z => n33370);
   U26553 : NAND2_X2 port map( A1 => n2657, A2 => n25532, ZN => n11292);
   U26569 : NAND2_X2 port map( A1 => n9175, A2 => n5356, ZN => n26083);
   U26580 : OR2_X1 port map( A1 => n28152, A2 => n32186, Z => n36712);
   U26601 : XOR2_X1 port map( A1 => n36334, A2 => n3331, Z => n36447);
   U26606 : XOR2_X1 port map( A1 => n36335, A2 => n11553, Z => n17292);
   U26607 : XOR2_X1 port map( A1 => n14385, A2 => n25155, Z => n36335);
   U26616 : NOR2_X2 port map( A1 => n36337, A2 => n36336, ZN => n12567);
   U26620 : INV_X2 port map( I => n36338, ZN => n11512);
   U26669 : NAND2_X2 port map( A1 => n17810, A2 => n19070, ZN => n36341);
   U26681 : OAI22_X1 port map( A1 => n21678, A2 => n36455, B1 => n21825, B2 => 
                           n21861, ZN => n21679);
   U26682 : OAI22_X2 port map( A1 => n36346, A2 => n14549, B1 => n18712, B2 => 
                           n18710, ZN => n18711);
   U26694 : XOR2_X1 port map( A1 => n36349, A2 => n1169, Z => n17812);
   U26696 : OAI21_X1 port map( A1 => n39830, A2 => n21023, B => n35252, ZN => 
                           n18107);
   U26697 : BUF_X2 port map( I => n21858, Z => n36351);
   U26707 : OR2_X1 port map( A1 => n14139, A2 => n22262, Z => n21990);
   U26714 : OR2_X1 port map( A1 => n33644, A2 => n7512, Z => n36352);
   U26722 : NOR2_X2 port map( A1 => n36606, A2 => n36353, ZN => n33140);
   U26724 : INV_X1 port map( I => n36354, ZN => n21919);
   U26727 : AOI21_X2 port map( A1 => n21921, A2 => n36354, B => n8468, ZN => 
                           n15441);
   U26728 : NAND2_X1 port map( A1 => n670, A2 => n293, ZN => n36354);
   U26746 : NAND2_X2 port map( A1 => n423, A2 => n422, ZN => n36471);
   U26749 : INV_X2 port map( I => n36357, ZN => n12246);
   U26756 : OAI21_X2 port map( A1 => n1351, A2 => n36887, B => n21656, ZN => 
                           n36358);
   U26760 : XOR2_X1 port map( A1 => n36360, A2 => n37129, Z => n27643);
   U26769 : XOR2_X1 port map( A1 => n27523, A2 => n27852, Z => n36360);
   U26773 : INV_X2 port map( I => n22215, ZN => n6576);
   U26775 : OAI22_X2 port map( A1 => n15274, A2 => n15292, B1 => n11172, B2 => 
                           n21629, ZN => n22215);
   U26781 : XOR2_X1 port map( A1 => n37101, A2 => n36364, Z => n36363);
   U26789 : INV_X1 port map( I => n29983, ZN => n36364);
   U26796 : XOR2_X1 port map( A1 => n4039, A2 => n26500, Z => n36366);
   U26811 : XNOR2_X1 port map( A1 => n23904, A2 => n23681, ZN => n36646);
   U26816 : INV_X2 port map( I => n11354, ZN => n36369);
   U26818 : AOI22_X1 port map( A1 => n18483, A2 => n30112, B1 => n32933, B2 => 
                           n30102, ZN => n30105);
   U26826 : OAI22_X2 port map( A1 => n28611, A2 => n35173, B1 => n1434, B2 => 
                           n28496, ZN => n28539);
   U26827 : NAND2_X2 port map( A1 => n33620, A2 => n15570, ZN => n28356);
   U26831 : OR2_X1 port map( A1 => n34019, A2 => n21001, Z => n20999);
   U26834 : XOR2_X1 port map( A1 => n36372, A2 => n36373, Z => n33008);
   U26846 : NAND2_X1 port map( A1 => n35895, A2 => n27320, ZN => n18669);
   U26858 : XOR2_X1 port map( A1 => n36377, A2 => n29162, Z => n11384);
   U26860 : XOR2_X1 port map( A1 => n9131, A2 => n1411, Z => n36377);
   U26861 : NOR2_X2 port map( A1 => n1603, A2 => n15320, ZN => n32297);
   U26864 : XOR2_X1 port map( A1 => n31563, A2 => n34135, Z => n12830);
   U26880 : XOR2_X1 port map( A1 => n24006, A2 => n24007, Z => n36379);
   U26888 : XOR2_X1 port map( A1 => n25155, A2 => n24922, Z => n14214);
   U26890 : NAND2_X2 port map( A1 => n685, A2 => n10652, ZN => n15350);
   U26897 : XOR2_X1 port map( A1 => n13504, A2 => n36388, Z => n13503);
   U26898 : XOR2_X1 port map( A1 => n8113, A2 => n8982, Z => n36388);
   U26903 : XOR2_X1 port map( A1 => n11372, A2 => n23898, Z => n36389);
   U26904 : OR2_X1 port map( A1 => n25808, A2 => n33997, Z => n3806);
   U26928 : INV_X2 port map( I => n20573, ZN => n36392);
   U26932 : XOR2_X1 port map( A1 => n17039, A2 => n6433, Z => n28946);
   U26937 : AOI21_X2 port map( A1 => n28799, A2 => n28798, B => n28670, ZN => 
                           n17039);
   U26947 : INV_X2 port map( I => n19675, ZN => n28669);
   U26948 : OAI22_X2 port map( A1 => n15204, A2 => n31832, B1 => n15014, B2 => 
                           n17477, ZN => n19675);
   U26953 : INV_X2 port map( I => n36396, ZN => n37061);
   U26968 : NOR2_X2 port map( A1 => n1119, A2 => n7810, ZN => n548);
   U26995 : XOR2_X1 port map( A1 => n7744, A2 => n30122, Z => n9777);
   U26998 : NOR2_X2 port map( A1 => n38302, A2 => n6849, ZN => n6850);
   U26999 : XOR2_X1 port map( A1 => n36400, A2 => n30682, Z => Ciphertext(130))
                           ;
   U27010 : NOR2_X1 port map( A1 => n31726, A2 => n31727, ZN => n36400);
   U27013 : XOR2_X1 port map( A1 => n11667, A2 => n38218, Z => n25595);
   U27016 : XOR2_X1 port map( A1 => n28984, A2 => n31398, Z => n31377);
   U27017 : XOR2_X1 port map( A1 => n10237, A2 => n36406, Z => n10247);
   U27027 : NAND2_X2 port map( A1 => n36408, A2 => n2635, ZN => n25284);
   U27047 : AOI21_X1 port map( A1 => n31231, A2 => n13986, B => n15189, ZN => 
                           n36410);
   U27049 : OAI21_X2 port map( A1 => n36412, A2 => n36411, B => n19813, ZN => 
                           n20186);
   U27080 : NOR3_X1 port map( A1 => n36415, A2 => n36413, A3 => n5152, ZN => 
                           n5151);
   U27083 : NOR2_X1 port map( A1 => n36671, A2 => n36414, ZN => n36413);
   U27093 : AND2_X1 port map( A1 => n36671, A2 => n31015, Z => n36415);
   U27097 : NAND2_X2 port map( A1 => n36416, A2 => n15017, ZN => n12243);
   U27099 : NAND3_X1 port map( A1 => n34019, A2 => n13980, A3 => n21001, ZN => 
                           n36416);
   U27100 : XOR2_X1 port map( A1 => n24838, A2 => n36418, Z => n7377);
   U27103 : XOR2_X1 port map( A1 => n34142, A2 => n24836, Z => n36418);
   U27108 : OR2_X1 port map( A1 => n11726, A2 => n8413, Z => n3255);
   U27112 : XOR2_X1 port map( A1 => n23782, A2 => n599, Z => n3167);
   U27116 : XOR2_X1 port map( A1 => n31563, A2 => n34032, Z => n36423);
   U27126 : NAND2_X1 port map( A1 => n16366, A2 => n18920, ZN => n30368);
   U27132 : AOI21_X2 port map( A1 => n4226, A2 => n4225, B => n34123, ZN => 
                           n4224);
   U27143 : OAI21_X2 port map( A1 => n14065, A2 => n3449, B => n20004, ZN => 
                           n33001);
   U27154 : INV_X2 port map( I => n36435, ZN => n12066);
   U27157 : NAND2_X2 port map( A1 => n16237, A2 => n997, ZN => n27011);
   U27176 : NOR2_X2 port map( A1 => n9835, A2 => n23477, ZN => n12008);
   U27187 : OAI21_X2 port map( A1 => n36441, A2 => n20752, B => n21939, ZN => 
                           n20751);
   U27194 : OAI21_X2 port map( A1 => n36621, A2 => n36622, B => n24357, ZN => 
                           n33224);
   U27200 : XOR2_X1 port map( A1 => n12997, A2 => n9808, Z => n13413);
   U27206 : NAND2_X2 port map( A1 => n36446, A2 => n4372, ZN => n5084);
   U27209 : INV_X2 port map( I => n36447, ZN => n32623);
   U27217 : BUF_X2 port map( I => n32024, Z => n36448);
   U27218 : NOR2_X1 port map( A1 => n36450, A2 => n3509, ZN => n36449);
   U27220 : INV_X1 port map( I => n16569, ZN => n36451);
   U27224 : INV_X1 port map( I => n36452, ZN => n28172);
   U27227 : NAND2_X1 port map( A1 => n19467, A2 => n32474, ZN => n36452);
   U27234 : NAND2_X2 port map( A1 => n4, A2 => n3, ZN => n1487);
   U27241 : INV_X2 port map( I => n36454, ZN => n7160);
   U27247 : INV_X1 port map( I => n21858, ZN => n36455);
   U27249 : XOR2_X1 port map( A1 => Plaintext(46), A2 => Key(46), Z => n21858);
   U27262 : XOR2_X1 port map( A1 => n13673, A2 => n13674, Z => n36456);
   U27269 : XOR2_X1 port map( A1 => n3530, A2 => n3529, Z => n20482);
   U27276 : NAND2_X1 port map( A1 => n37776, A2 => n28458, ZN => n28383);
   U27286 : BUF_X2 port map( I => n23873, Z => n36461);
   U27290 : XOR2_X1 port map( A1 => n29294, A2 => n5991, Z => n36939);
   U27301 : AOI21_X1 port map( A1 => n27311, A2 => n16243, B => n27412, ZN => 
                           n33261);
   U27303 : XOR2_X1 port map( A1 => n8782, A2 => n9038, Z => n8781);
   U27306 : OAI21_X2 port map( A1 => n21940, A2 => n21941, B => n21939, ZN => 
                           n36464);
   U27339 : XOR2_X1 port map( A1 => n22704, A2 => n22702, Z => n36869);
   U27344 : XOR2_X1 port map( A1 => n22464, A2 => n19931, Z => n22702);
   U27349 : XOR2_X1 port map( A1 => n7762, A2 => n5517, Z => n5709);
   U27357 : INV_X1 port map( I => n4123, ZN => n22483);
   U27365 : NAND2_X2 port map( A1 => n4121, A2 => n4122, ZN => n4123);
   U27371 : XOR2_X1 port map( A1 => n36468, A2 => n14302, Z => n14060);
   U27372 : AOI22_X2 port map( A1 => n12079, A2 => n2186, B1 => n22030, B2 => 
                           n11508, ZN => n11507);
   U27374 : NOR2_X2 port map( A1 => n5075, A2 => n37217, ZN => n12079);
   U27398 : XOR2_X1 port map( A1 => n22543, A2 => n6711, Z => n6710);
   U27399 : XOR2_X1 port map( A1 => n23933, A2 => n23883, Z => n23835);
   U27410 : NOR2_X2 port map( A1 => n16758, A2 => n16757, ZN => n23933);
   U27423 : NOR2_X2 port map( A1 => n27053, A2 => n27337, ZN => n27344);
   U27425 : INV_X2 port map( I => n36470, ZN => n19426);
   U27426 : XNOR2_X1 port map( A1 => n16942, A2 => n20767, ZN => n36470);
   U27433 : XOR2_X1 port map( A1 => n18359, A2 => n22603, Z => n17284);
   U27441 : NAND2_X1 port map( A1 => n3869, A2 => n24477, ZN => n16159);
   U27447 : OAI21_X2 port map( A1 => n20565, A2 => n25526, B => n1539, ZN => 
                           n36472);
   U27456 : OR2_X1 port map( A1 => n20735, A2 => n21145, Z => n36474);
   U27462 : NAND2_X2 port map( A1 => n36476, A2 => n13698, ZN => n27392);
   U27485 : OAI21_X2 port map( A1 => n34040, A2 => n24514, B => n31797, ZN => 
                           n25104);
   U27499 : XOR2_X1 port map( A1 => n26290, A2 => n26379, Z => n26242);
   U27524 : AND2_X1 port map( A1 => n18157, A2 => n33550, Z => n33141);
   U27537 : BUF_X2 port map( I => n24411, Z => n36485);
   U27553 : AOI21_X2 port map( A1 => n36885, A2 => n32930, B => n32024, ZN => 
                           n17093);
   U27561 : INV_X2 port map( I => n39820, ZN => n36486);
   U27562 : NOR2_X2 port map( A1 => n36488, A2 => n36487, ZN => n18838);
   U27581 : NAND2_X2 port map( A1 => n18605, A2 => n30585, ZN => n16835);
   U27584 : XNOR2_X1 port map( A1 => n14902, A2 => n22787, ZN => n16802);
   U27590 : XOR2_X1 port map( A1 => n22671, A2 => n16798, Z => n14902);
   U27602 : OAI22_X2 port map( A1 => n34067, A2 => n36490, B1 => n19483, B2 => 
                           n10144, ZN => n11173);
   U27603 : INV_X2 port map( I => n13959, ZN => n36490);
   U27610 : XOR2_X1 port map( A1 => n36491, A2 => n19879, Z => Ciphertext(63));
   U27615 : NAND3_X2 port map( A1 => n7437, A2 => n7436, A3 => n7435, ZN => 
                           n36491);
   U27622 : XOR2_X1 port map( A1 => n2662, A2 => n36493, Z => n33947);
   U27636 : XOR2_X1 port map( A1 => n24981, A2 => n36494, Z => n36493);
   U27652 : OAI22_X2 port map( A1 => n20496, A2 => n20495, B1 => n28460, B2 => 
                           n28378, ZN => n20492);
   U27665 : XOR2_X1 port map( A1 => n28041, A2 => n36498, Z => n19920);
   U27666 : XOR2_X1 port map( A1 => n28040, A2 => n18159, Z => n36498);
   U27673 : NAND2_X2 port map( A1 => n3004, A2 => n36499, ZN => n2349);
   U27679 : INV_X4 port map( I => n3455, ZN => n16200);
   U27681 : NAND2_X2 port map( A1 => n3175, A2 => n30813, ZN => n3455);
   U27682 : NAND2_X2 port map( A1 => n18718, A2 => n19504, ZN => n36840);
   U27687 : NAND2_X2 port map( A1 => n8990, A2 => n36501, ZN => n8798);
   U27696 : NAND2_X2 port map( A1 => n36502, A2 => n24856, ZN => n18536);
   U27703 : OAI21_X2 port map( A1 => n20690, A2 => n20689, B => n24853, ZN => 
                           n36502);
   U27726 : OR2_X1 port map( A1 => n28205, A2 => n118, Z => n14361);
   U27732 : XOR2_X1 port map( A1 => n26181, A2 => n34165, Z => n26368);
   U27742 : NOR3_X1 port map( A1 => n10436, A2 => n8452, A3 => n23159, ZN => 
                           n36506);
   U27753 : NOR2_X1 port map( A1 => n16786, A2 => n14254, ZN => n7194);
   U27754 : XOR2_X1 port map( A1 => n33962, A2 => n16787, Z => n16786);
   U27760 : NAND3_X2 port map( A1 => n33675, A2 => n8914, A3 => n8913, ZN => 
                           n29052);
   U27767 : XOR2_X1 port map( A1 => n32766, A2 => n26542, Z => n36508);
   U27776 : XOR2_X1 port map( A1 => n26415, A2 => n36511, Z => n36510);
   U27791 : XOR2_X1 port map( A1 => n36758, A2 => n36513, Z => n746);
   U27813 : INV_X2 port map( I => n36514, ZN => n30186);
   U27827 : XOR2_X1 port map( A1 => n7944, A2 => n36516, Z => n36515);
   U27830 : INV_X2 port map( I => n3448, ZN => n36516);
   U27835 : NAND2_X2 port map( A1 => n25354, A2 => n25353, ZN => n36922);
   U27844 : NAND2_X2 port map( A1 => n35232, A2 => n31612, ZN => n23636);
   U27858 : OAI21_X2 port map( A1 => n18742, A2 => n15437, B => n36518, ZN => 
                           n9616);
   U27862 : XOR2_X1 port map( A1 => n19862, A2 => n1553, Z => n2184);
   U27868 : INV_X4 port map( I => n36523, ZN => n5101);
   U27880 : NAND2_X1 port map( A1 => n17710, A2 => n24145, ZN => n14051);
   U27899 : INV_X2 port map( I => n28117, ZN => n3159);
   U27905 : NOR2_X1 port map( A1 => n36532, A2 => n1827, ZN => n8156);
   U27921 : XOR2_X1 port map( A1 => n21098, A2 => n20082, Z => n14319);
   U27934 : NOR2_X1 port map( A1 => n34279, A2 => n31433, ZN => n30486);
   U27937 : OAI21_X2 port map( A1 => n26353, A2 => n18606, B => n14824, ZN => 
                           n31433);
   U27943 : INV_X2 port map( I => n29113, ZN => n5153);
   U27944 : NAND2_X2 port map( A1 => n5154, A2 => n1741, ZN => n29113);
   U27945 : XOR2_X1 port map( A1 => n36537, A2 => n12179, Z => n14401);
   U27954 : AND2_X1 port map( A1 => n6592, A2 => n18545, Z => n25676);
   U27974 : XOR2_X1 port map( A1 => n23959, A2 => n36541, Z => n36540);
   U27976 : INV_X2 port map( I => n23487, ZN => n21247);
   U27977 : NAND2_X2 port map( A1 => n22983, A2 => n22984, ZN => n23487);
   U28002 : NAND2_X1 port map( A1 => n5207, A2 => n5206, ZN => n5205);
   U28012 : INV_X2 port map( I => n36543, ZN => n668);
   U28013 : XOR2_X1 port map( A1 => Plaintext(180), A2 => Key(180), Z => n36543
                           );
   U28024 : XOR2_X1 port map( A1 => n6513, A2 => n6511, Z => n18707);
   U28035 : INV_X1 port map( I => n26828, ZN => n32892);
   U28036 : NAND2_X1 port map( A1 => n15386, A2 => n32623, ZN => n26828);
   U28044 : NOR2_X1 port map( A1 => n29384, A2 => n31279, ZN => n36550);
   U28048 : NAND2_X2 port map( A1 => n21246, A2 => n36551, ZN => n23600);
   U28049 : INV_X2 port map( I => n22973, ZN => n36554);
   U28064 : NAND2_X1 port map( A1 => n21052, A2 => n35809, ZN => n30728);
   U28069 : NAND2_X1 port map( A1 => n23034, A2 => n23035, ZN => n23037);
   U28078 : NOR2_X1 port map( A1 => n28048, A2 => n34410, ZN => n36558);
   U28081 : INV_X1 port map( I => n4975, ZN => n36559);
   U28085 : NOR2_X1 port map( A1 => n30015, A2 => n30037, ZN => n30031);
   U28113 : XOR2_X1 port map( A1 => n23980, A2 => n32174, Z => n21267);
   U28116 : NAND2_X2 port map( A1 => n8138, A2 => n32506, ZN => n23980);
   U28121 : OAI21_X2 port map( A1 => n2574, A2 => n36568, B => n2679, ZN => 
                           n5031);
   U28157 : INV_X4 port map( I => n23426, ZN => n2798);
   U28195 : XOR2_X1 port map( A1 => n27756, A2 => n9184, Z => n10818);
   U28196 : NOR2_X1 port map( A1 => n29683, A2 => n31538, ZN => n18794);
   U28235 : AND2_X1 port map( A1 => n36571, A2 => n33440, Z => n10889);
   U28248 : XOR2_X1 port map( A1 => n23852, A2 => n36572, Z => n16245);
   U28249 : XOR2_X1 port map( A1 => n13978, A2 => n6561, Z => n36572);
   U28252 : XOR2_X1 port map( A1 => n36576, A2 => n24990, Z => n25546);
   U28255 : XOR2_X1 port map( A1 => n9389, A2 => n729, Z => n36576);
   U28267 : NAND2_X2 port map( A1 => n36577, A2 => n17441, ZN => n23888);
   U28295 : OAI21_X2 port map( A1 => n6514, A2 => n36263, B => n19232, ZN => 
                           n23416);
   U28304 : XOR2_X1 port map( A1 => n26454, A2 => n26433, Z => n11072);
   U28311 : NAND2_X2 port map( A1 => n14988, A2 => n14990, ZN => n27448);
   U28324 : NOR3_X1 port map( A1 => n11226, A2 => n36480, A3 => n38377, ZN => 
                           n3402);
   U28338 : NAND2_X1 port map( A1 => n13226, A2 => n1143, ZN => n22369);
   U28345 : NAND2_X1 port map( A1 => n6543, A2 => n25860, ZN => n36581);
   U28365 : NAND2_X2 port map( A1 => n1587, A2 => n24398, ZN => n9583);
   U28366 : NAND2_X2 port map( A1 => n9783, A2 => n33574, ZN => n10079);
   U28373 : INV_X1 port map( I => n998, ZN => n27189);
   U28384 : NOR2_X2 port map( A1 => n36584, A2 => n24163, ZN => n7770);
   U28420 : NAND2_X1 port map( A1 => n17677, A2 => n38656, ZN => n36587);
   U28429 : OR2_X1 port map( A1 => n7291, A2 => n9875, Z => n36679);
   U28457 : NAND2_X2 port map( A1 => n20604, A2 => n36589, ZN => n21272);
   U28480 : NOR2_X2 port map( A1 => n29779, A2 => n29776, ZN => n36590);
   U28506 : AOI21_X2 port map( A1 => n36593, A2 => n36592, B => n35611, ZN => 
                           n18565);
   U28513 : NAND2_X2 port map( A1 => n36594, A2 => n3083, ZN => n11922);
   U28521 : NOR2_X2 port map( A1 => n12324, A2 => n12325, ZN => n20353);
   U28546 : OAI21_X2 port map( A1 => n21564, A2 => n19397, B => n11433, ZN => 
                           n22113);
   U28547 : NOR2_X2 port map( A1 => n30835, A2 => n9190, ZN => n16236);
   U28548 : NAND2_X2 port map( A1 => n36598, A2 => n14762, ZN => n18273);
   U28553 : OR2_X1 port map( A1 => n12235, A2 => n8205, Z => n16666);
   U28557 : XOR2_X1 port map( A1 => n32219, A2 => n14978, Z => n15037);
   U28558 : OAI21_X1 port map( A1 => n4192, A2 => n32566, B => n38187, ZN => 
                           n2502);
   U28559 : AOI21_X2 port map( A1 => n2428, A2 => n3088, B => n32940, ZN => 
                           n27845);
   U28562 : NOR2_X2 port map( A1 => n33412, A2 => n24821, ZN => n6770);
   U28589 : NAND2_X1 port map( A1 => n29699, A2 => n29195, ZN => n29633);
   U28605 : INV_X2 port map( I => n36601, ZN => n858);
   U28611 : XOR2_X1 port map( A1 => n15818, A2 => n15821, Z => n36601);
   U28614 : NOR2_X1 port map( A1 => n36981, A2 => n27240, ZN => n17354);
   U28618 : XOR2_X1 port map( A1 => n36603, A2 => n36602, Z => n31272);
   U28644 : NOR2_X1 port map( A1 => n28330, A2 => n17583, ZN => n28738);
   U28662 : XOR2_X1 port map( A1 => n14294, A2 => n36604, Z => n550);
   U28663 : XOR2_X1 port map( A1 => n9937, A2 => n36605, Z => n36604);
   U28669 : NOR3_X1 port map( A1 => n14600, A2 => n14158, A3 => n29815, ZN => 
                           n17912);
   U28670 : AOI21_X2 port map( A1 => n21558, A2 => n21559, B => n21920, ZN => 
                           n36606);
   U28673 : XOR2_X1 port map( A1 => n36608, A2 => n8547, Z => n8546);
   U28674 : XOR2_X1 port map( A1 => n17812, A2 => n22444, Z => n36608);
   U28703 : XOR2_X1 port map( A1 => n31563, A2 => n3576, Z => n3579);
   U28737 : NOR2_X2 port map( A1 => n2759, A2 => n21672, ZN => n31480);
   U28755 : NAND2_X1 port map( A1 => n14877, A2 => n19724, ZN => n14876);
   U28759 : AOI21_X2 port map( A1 => n36611, A2 => n20515, B => n3602, ZN => 
                           n10775);
   U28767 : NAND2_X2 port map( A1 => n7802, A2 => n19495, ZN => n36611);
   U28775 : NAND2_X1 port map( A1 => n29632, A2 => n29701, ZN => n29197);
   U28778 : XOR2_X1 port map( A1 => n36613, A2 => n33309, Z => n21126);
   U28789 : XOR2_X1 port map( A1 => n36223, A2 => n10673, Z => n36613);
   U28810 : XOR2_X1 port map( A1 => n32448, A2 => n11923, Z => n11015);
   U28832 : AND3_X1 port map( A1 => n16240, A2 => n31362, A3 => n33514, Z => 
                           n7888);
   U28837 : NAND3_X2 port map( A1 => n36615, A2 => n10676, A3 => n35777, ZN => 
                           n9955);
   U28854 : OAI21_X1 port map( A1 => n32651, A2 => n24565, B => n36618, ZN => 
                           n20301);
   U28876 : NAND2_X2 port map( A1 => n17687, A2 => n18986, ZN => n27466);
   U28877 : INV_X2 port map( I => n36620, ZN => n10047);
   U28880 : XOR2_X1 port map( A1 => n16563, A2 => n16560, Z => n36620);
   U28890 : XOR2_X1 port map( A1 => n5836, A2 => n3233, Z => n3232);
   U28892 : NOR2_X2 port map( A1 => n11173, A2 => n11174, ZN => n11327);
   U28918 : NOR2_X1 port map( A1 => n32099, A2 => n19499, ZN => n7261);
   U28921 : NAND2_X2 port map( A1 => n7263, A2 => n10791, ZN => n9053);
   U28934 : XOR2_X1 port map( A1 => n27840, A2 => n18650, Z => n13791);
   U29008 : NAND2_X2 port map( A1 => n19539, A2 => n19540, ZN => n30096);
   U29018 : AOI21_X2 port map( A1 => n18328, A2 => n30526, B => n1606, ZN => 
                           n36626);
   U29024 : XOR2_X1 port map( A1 => n36627, A2 => n27881, Z => n29483);
   U29026 : XOR2_X1 port map( A1 => n13381, A2 => n27880, Z => n36627);
   U29029 : OAI21_X2 port map( A1 => n10564, A2 => n10565, B => n32009, ZN => 
                           n31048);
   U29031 : XOR2_X1 port map( A1 => n38560, A2 => n30865, Z => n16431);
   U29033 : OAI21_X1 port map( A1 => n31859, A2 => n1331, B => n31860, ZN => 
                           n18729);
   U29041 : XOR2_X1 port map( A1 => n31261, A2 => n19881, Z => n32001);
   U29051 : XOR2_X1 port map( A1 => n4612, A2 => n23717, Z => n23722);
   U29056 : XOR2_X1 port map( A1 => n25286, A2 => n25081, Z => n5816);
   U29063 : XOR2_X1 port map( A1 => n11321, A2 => n25014, Z => n25081);
   U29072 : INV_X1 port map( I => n25355, ZN => n25449);
   U29073 : XOR2_X1 port map( A1 => n17108, A2 => n36799, Z => n25355);
   U29074 : NAND2_X2 port map( A1 => n36629, A2 => n12075, ZN => n27697);
   U29077 : NOR2_X2 port map( A1 => n12073, A2 => n12072, ZN => n36629);
   U29081 : OAI21_X2 port map( A1 => n36443, A2 => n32609, B => n36631, ZN => 
                           n9735);
   U29086 : NAND2_X2 port map( A1 => n36632, A2 => n32609, ZN => n36631);
   U29122 : XOR2_X1 port map( A1 => n36637, A2 => n8401, Z => n8301);
   U29143 : XOR2_X1 port map( A1 => n9712, A2 => n32203, Z => n17198);
   U29148 : INV_X2 port map( I => n2430, ZN => n22899);
   U29152 : XOR2_X1 port map( A1 => n2200, A2 => n2198, Z => n2430);
   U29171 : NAND2_X1 port map( A1 => n5966, A2 => n17405, ZN => n28045);
   U29180 : XOR2_X1 port map( A1 => n25809, A2 => n16294, Z => n36644);
   U29203 : XOR2_X1 port map( A1 => n12515, A2 => n16278, Z => n36645);
   U29204 : XOR2_X1 port map( A1 => n737, A2 => n26401, Z => n6963);
   U29209 : NAND2_X1 port map( A1 => n5174, A2 => n11616, ZN => n36957);
   U29214 : BUF_X2 port map( I => n4342, Z => n36649);
   U29219 : OR2_X1 port map( A1 => n13998, A2 => n18959, Z => n13956);
   U29220 : OAI21_X1 port map( A1 => n34066, A2 => n21645, B => n36651, ZN => 
                           n21648);
   U29223 : NAND2_X1 port map( A1 => n21642, A2 => n21645, ZN => n36651);
   U29226 : NAND2_X2 port map( A1 => n16732, A2 => n16731, ZN => n32024);
   U29228 : NAND2_X1 port map( A1 => n22822, A2 => n7387, ZN => n36654);
   U29240 : XOR2_X1 port map( A1 => n10399, A2 => n1457, Z => n36656);
   U29246 : NAND2_X2 port map( A1 => n2736, A2 => n2737, ZN => n4108);
   U29247 : XOR2_X1 port map( A1 => n5802, A2 => n12139, Z => n13205);
   U29259 : AOI22_X2 port map( A1 => n13009, A2 => n11044, B1 => n8792, B2 => 
                           n196, ZN => n13008);
   U29276 : NAND2_X2 port map( A1 => n32832, A2 => n8362, ZN => n17454);
   U29286 : OAI21_X2 port map( A1 => n7216, A2 => n1339, B => n36661, ZN => 
                           n36660);
   U29287 : XOR2_X1 port map( A1 => n13977, A2 => n19344, Z => n19343);
   U29295 : XOR2_X1 port map( A1 => n25263, A2 => n18432, Z => n17593);
   U29297 : BUF_X2 port map( I => n7063, Z => n36663);
   U29298 : XOR2_X1 port map( A1 => n31823, A2 => n26480, Z => n26182);
   U29306 : XOR2_X1 port map( A1 => n36727, A2 => n16753, Z => n33182);
   U29312 : NAND2_X2 port map( A1 => n32292, A2 => n18825, ZN => n22240);
   U29333 : INV_X2 port map( I => n26128, ZN => n36666);
   U29371 : XOR2_X1 port map( A1 => n4875, A2 => n6523, Z => n5534);
   U29377 : NAND2_X1 port map( A1 => n36674, A2 => n8691, ZN => n20074);
   U29386 : OAI21_X2 port map( A1 => n29988, A2 => n30051, B => n10943, ZN => 
                           n30038);
   U29392 : OAI22_X2 port map( A1 => n15936, A2 => n36673, B1 => n7267, B2 => 
                           n24799, ZN => n14781);
   U29400 : NAND2_X2 port map( A1 => n22828, A2 => n20907, ZN => n5258);
   U29445 : XOR2_X1 port map( A1 => n38816, A2 => n31218, Z => n36687);
   U29470 : XOR2_X1 port map( A1 => n6661, A2 => n30101, Z => n28986);
   U29483 : NAND2_X1 port map( A1 => n29207, A2 => n11973, ZN => n9807);
   U29494 : NOR2_X1 port map( A1 => n19610, A2 => n36691, ZN => n19482);
   U29498 : NOR2_X1 port map( A1 => n21141, A2 => n19893, ZN => n36691);
   U29516 : XOR2_X1 port map( A1 => n20554, A2 => n36692, Z => n30562);
   U29517 : XOR2_X1 port map( A1 => n25016, A2 => n25324, Z => n36692);
   U29518 : XOR2_X1 port map( A1 => n23725, A2 => n17563, Z => n10941);
   U29520 : NAND3_X1 port map( A1 => n15043, A2 => n15044, A3 => n29410, ZN => 
                           n7733);
   U29528 : AND2_X1 port map( A1 => n31287, A2 => n27424, Z => n30475);
   U29529 : NAND2_X1 port map( A1 => n33201, A2 => n33202, ZN => n33200);
   U29541 : NAND2_X2 port map( A1 => n22805, A2 => n36696, ZN => n14856);
   U29552 : OAI22_X2 port map( A1 => n12960, A2 => n32740, B1 => n22892, B2 => 
                           n33925, ZN => n36696);
   U29553 : OAI22_X1 port map( A1 => n3039, A2 => n5569, B1 => n38601, B2 => 
                           n3040, ZN => n16197);
   U29554 : XOR2_X1 port map( A1 => n4279, A2 => n36698, Z => n31920);
   U29557 : NOR2_X1 port map( A1 => n31271, A2 => n8193, ZN => n5);
   U29561 : NOR2_X2 port map( A1 => n29591, A2 => n28550, ZN => n2296);
   U29585 : XOR2_X1 port map( A1 => n29835, A2 => n36702, Z => n12763);
   U29587 : XOR2_X1 port map( A1 => n12765, A2 => n28819, Z => n36702);
   U29588 : AOI21_X2 port map( A1 => n9816, A2 => n13375, B => n12417, ZN => 
                           n12416);
   U29594 : NOR2_X2 port map( A1 => n39671, A2 => n20740, ZN => n27232);
   U29607 : NOR2_X1 port map( A1 => n16154, A2 => n37671, ZN => n36703);
   U29615 : XOR2_X1 port map( A1 => n3521, A2 => n5185, Z => n12973);
   U29619 : INV_X2 port map( I => n18994, ZN => n1245);
   U29635 : NAND2_X1 port map( A1 => n1046, A2 => n23140, ZN => n21047);
   U29667 : AOI22_X2 port map( A1 => n20411, A2 => n3120, B1 => n11710, B2 => 
                           n24847, ZN => n24731);
   U29671 : OR2_X1 port map( A1 => n21339, A2 => n21687, Z => n4750);
   U29682 : AOI21_X2 port map( A1 => n9721, A2 => n36712, B => n33902, ZN => 
                           n30837);
   U29716 : OAI22_X2 port map( A1 => n1071, A2 => n20157, B1 => n28118, B2 => 
                           n19667, ZN => n28140);
   U29717 : XOR2_X1 port map( A1 => n22754, A2 => n18001, Z => n5571);
   U29737 : INV_X2 port map( I => n36717, ZN => n37051);
   U29745 : XOR2_X1 port map( A1 => n36718, A2 => n13928, Z => n17022);
   U29749 : XOR2_X1 port map( A1 => n31790, A2 => n26408, Z => n36718);
   U29753 : XOR2_X1 port map( A1 => n3553, A2 => n36719, Z => n5078);
   U29760 : XOR2_X1 port map( A1 => n35065, A2 => n13193, Z => n2739);
   U29779 : NOR2_X2 port map( A1 => n15466, A2 => n12044, ZN => n21929);
   U29797 : NAND2_X2 port map( A1 => n32577, A2 => n26717, ZN => n21101);
   U29799 : XOR2_X1 port map( A1 => n22678, A2 => n36723, Z => n23131);
   U29801 : XOR2_X1 port map( A1 => n11985, A2 => n11984, Z => n36723);
   U29802 : NAND2_X1 port map( A1 => n22313, A2 => n36151, ZN => n22314);
   U29804 : NOR2_X2 port map( A1 => n18636, A2 => n32753, ZN => n36726);
   U29806 : XOR2_X1 port map( A1 => n10982, A2 => n10984, Z => n27882);
   U29816 : XOR2_X1 port map( A1 => n1658, A2 => n4819, Z => n36727);
   U29820 : NOR2_X2 port map( A1 => n22254, A2 => n32675, ZN => n22126);
   U29826 : XOR2_X1 port map( A1 => n10484, A2 => n10486, Z => n19746);
   U29833 : OAI21_X1 port map( A1 => n1787, A2 => n1095, B => n14380, ZN => 
                           n26954);
   U29849 : NAND2_X2 port map( A1 => n13096, A2 => n26958, ZN => n19529);
   U29852 : OAI21_X2 port map( A1 => n12461, A2 => n12460, B => n36729, ZN => 
                           n25301);
   U29861 : XOR2_X1 port map( A1 => n24974, A2 => n36730, Z => n31410);
   U29863 : XOR2_X1 port map( A1 => n26376, A2 => n26289, Z => n8844);
   U29882 : XOR2_X1 port map( A1 => n19384, A2 => n26582, Z => n26286);
   U29888 : XOR2_X1 port map( A1 => n36734, A2 => n25311, Z => n15034);
   U29891 : XOR2_X1 port map( A1 => n25031, A2 => n6066, Z => n36734);
   U29899 : XOR2_X1 port map( A1 => Plaintext(55), A2 => Key(55), Z => n7703);
   U29900 : INV_X2 port map( I => n13359, ZN => n36735);
   U29918 : NAND2_X1 port map( A1 => n36738, A2 => n30217, ZN => n36737);
   U29941 : NAND3_X1 port map( A1 => n14869, A2 => n30211, A3 => n33437, ZN => 
                           n31987);
   U29945 : NOR2_X1 port map( A1 => n1068, A2 => n28591, ZN => n4992);
   U29948 : OAI22_X2 port map( A1 => n36944, A2 => n28176, B1 => n28265, B2 => 
                           n28175, ZN => n28591);
   U29958 : OR2_X1 port map( A1 => n26090, A2 => n35828, Z => n25363);
   U29961 : NAND2_X1 port map( A1 => n28267, A2 => n37079, ZN => n31766);
   U29963 : NAND2_X2 port map( A1 => n36741, A2 => n37279, ZN => n2950);
   U29966 : NAND2_X2 port map( A1 => n23340, A2 => n23341, ZN => n36741);
   U29973 : NAND3_X2 port map( A1 => n13282, A2 => n13281, A3 => n13280, ZN => 
                           n6130);
   U29979 : NAND2_X1 port map( A1 => n18412, A2 => n35977, ZN => n8467);
   U29983 : AND2_X1 port map( A1 => n38848, A2 => n33996, Z => n18459);
   U29992 : NAND2_X1 port map( A1 => n36745, A2 => n22317, ZN => n36902);
   U29994 : NOR2_X1 port map( A1 => n31766, A2 => n31765, ZN => n36944);
   U29998 : OAI21_X2 port map( A1 => n9735, A2 => n38746, B => n9734, ZN => 
                           n22657);
   U29999 : XOR2_X1 port map( A1 => n35221, A2 => n22775, Z => n22689);
   U30000 : NOR2_X2 port map( A1 => n14800, A2 => n14801, ZN => n11644);
   U30008 : AOI22_X1 port map( A1 => n15230, A2 => n23042, B1 => n38329, B2 => 
                           n4714, ZN => n11914);
   U30020 : INV_X2 port map( I => n24038, ZN => n36748);
   U30024 : XOR2_X1 port map( A1 => n36894, A2 => n19801, Z => n16857);
   U30025 : XOR2_X1 port map( A1 => n29245, A2 => n11127, Z => n19727);
   U30026 : AOI21_X2 port map( A1 => n21631, A2 => n36519, B => n36751, ZN => 
                           n21634);
   U30031 : OR2_X1 port map( A1 => n10631, A2 => n20238, Z => n36753);
   U30032 : XOR2_X1 port map( A1 => n3823, A2 => n4118, Z => n36992);
   U30033 : XNOR2_X1 port map( A1 => n29300, A2 => n15617, ZN => n28836);
   U30036 : NAND2_X2 port map( A1 => n15514, A2 => n19726, ZN => n29300);
   U30040 : OAI22_X2 port map( A1 => n11213, A2 => n15237, B1 => n12090, B2 => 
                           n13186, ZN => n31132);
   U30057 : XOR2_X1 port map( A1 => n3616, A2 => n12664, Z => n36759);
   U30062 : NAND2_X2 port map( A1 => n7614, A2 => n36857, ZN => n20159);
   U30063 : NAND2_X2 port map( A1 => n33893, A2 => n5363, ZN => n27452);
   U30069 : INV_X2 port map( I => n9917, ZN => n28749);
   U30076 : NOR2_X2 port map( A1 => n31934, A2 => n36761, ZN => n17687);
   U30083 : BUF_X2 port map( I => n6205, Z => n36764);
   U30094 : XOR2_X1 port map( A1 => Plaintext(29), A2 => Key(29), Z => n36772);
   U30102 : INV_X2 port map( I => n36772, ZN => n21445);
   U30124 : NAND2_X1 port map( A1 => n33765, A2 => n31664, ZN => n36774);
   U30125 : NAND2_X2 port map( A1 => n28700, A2 => n36777, ZN => n36776);
   U30128 : NAND2_X2 port map( A1 => n21956, A2 => n21957, ZN => n22580);
   U30133 : NAND2_X2 port map( A1 => n21486, A2 => n36779, ZN => n22085);
   U30136 : AOI21_X2 port map( A1 => n21120, A2 => n36782, B => n21119, ZN => 
                           n23473);
   U30140 : NAND2_X1 port map( A1 => n13373, A2 => n36783, ZN => n36782);
   U30151 : XOR2_X1 port map( A1 => n30842, A2 => n9420, Z => n18433);
   U30157 : XOR2_X1 port map( A1 => n16492, A2 => n25269, Z => n25161);
   U30160 : NAND3_X2 port map( A1 => n16747, A2 => n2503, A3 => n16746, ZN => 
                           n16492);
   U30177 : INV_X2 port map( I => n9339, ZN => n10698);
   U30180 : NAND2_X1 port map( A1 => n23152, A2 => n2572, ZN => n9339);
   U30206 : XOR2_X1 port map( A1 => n10039, A2 => n10248, Z => n25581);
   U30208 : XOR2_X1 port map( A1 => n24892, A2 => n24891, Z => n36799);
   U30209 : XOR2_X1 port map( A1 => n23736, A2 => n10771, Z => n8016);
   U30216 : NOR3_X1 port map( A1 => n14704, A2 => n4986, A3 => n12771, ZN => 
                           n36800);
   U30217 : XOR2_X1 port map( A1 => n19009, A2 => n11458, Z => n11459);
   U30221 : XOR2_X1 port map( A1 => n12588, A2 => n26285, Z => n36803);
   U30222 : XOR2_X1 port map( A1 => n479, A2 => n27648, Z => n36804);
   U30230 : AOI21_X2 port map( A1 => n25878, A2 => n25879, B => n25877, ZN => 
                           n6989);
   U30232 : NAND2_X2 port map( A1 => n12889, A2 => n12888, ZN => n28886);
   U30233 : OAI21_X2 port map( A1 => n1521, A2 => n11036, B => n36807, ZN => 
                           n26403);
   U30239 : AOI21_X2 port map( A1 => n37116, A2 => n1521, B => n11032, ZN => 
                           n36807);
   U30244 : AOI21_X1 port map( A1 => n24228, A2 => n24328, B => n1607, ZN => 
                           n15496);
   U30250 : XOR2_X1 port map( A1 => n36808, A2 => n1358, Z => Ciphertext(107));
   U30257 : XOR2_X1 port map( A1 => n27673, A2 => n36809, Z => n31043);
   U30259 : OAI21_X2 port map( A1 => n18924, A2 => n13289, B => n12240, ZN => 
                           n27843);
   U30260 : NAND3_X2 port map( A1 => n25405, A2 => n25406, A3 => n25404, ZN => 
                           n3413);
   U30261 : AOI22_X1 port map( A1 => n30185, A2 => n31846, B1 => n39122, B2 => 
                           n30182, ZN => n4780);
   U30270 : XOR2_X1 port map( A1 => n29246, A2 => n36837, Z => n16787);
   U30272 : NAND2_X2 port map( A1 => n33833, A2 => n13818, ZN => n29246);
   U30278 : XOR2_X1 port map( A1 => n36812, A2 => n19200, Z => n15463);
   U30288 : INV_X2 port map( I => n30597, ZN => n3449);
   U30297 : XOR2_X1 port map( A1 => n38269, A2 => n38502, Z => n26415);
   U30303 : NAND2_X2 port map( A1 => n38874, A2 => n2716, ZN => n36817);
   U30305 : NAND3_X2 port map( A1 => n24511, A2 => n30414, A3 => n31986, ZN => 
                           n24869);
   U30306 : XOR2_X1 port map( A1 => n36822, A2 => n17406, Z => n17405);
   U30309 : NAND2_X1 port map( A1 => n30058, A2 => n37253, ZN => n36824);
   U30323 : NAND2_X1 port map( A1 => n37014, A2 => n36829, ZN => n37010);
   U30330 : XOR2_X1 port map( A1 => n36830, A2 => n16225, Z => n16704);
   U30337 : XOR2_X1 port map( A1 => n28979, A2 => n2914, Z => n36830);
   U30338 : INV_X2 port map( I => n36831, ZN => n30443);
   U30340 : XOR2_X1 port map( A1 => n28983, A2 => n17880, Z => n29026);
   U30343 : NAND2_X2 port map( A1 => n15295, A2 => n7030, ZN => n17880);
   U30347 : NAND2_X2 port map( A1 => n15360, A2 => n3313, ZN => n36833);
   U30350 : XOR2_X1 port map( A1 => n31339, A2 => n39136, Z => n12818);
   U30352 : NOR2_X2 port map( A1 => n22376, A2 => n22375, ZN => n31339);
   U30364 : AOI21_X2 port map( A1 => n10618, A2 => n36835, B => n888, ZN => 
                           n3221);
   U30372 : XOR2_X1 port map( A1 => n29289, A2 => n29081, Z => n36837);
   U30374 : BUF_X2 port map( I => n4472, Z => n36839);
   U30376 : XOR2_X1 port map( A1 => n21267, A2 => n23784, Z => n182);
   U30377 : XOR2_X1 port map( A1 => n22542, A2 => n22656, Z => n6709);
   U30378 : NAND2_X2 port map( A1 => n36843, A2 => n8419, ZN => n18081);
   U30379 : NOR2_X1 port map( A1 => n6657, A2 => n32486, ZN => n12131);
   U30380 : OAI22_X2 port map( A1 => n11848, A2 => n33263, B1 => n8481, B2 => 
                           n834, ZN => n25819);
   U30392 : XOR2_X1 port map( A1 => n22771, A2 => n22393, Z => n18914);
   U30400 : XOR2_X1 port map( A1 => n36847, A2 => n13426, Z => n13425);
   U30403 : XOR2_X1 port map( A1 => n26258, A2 => n26257, Z => n15453);
   U30407 : XOR2_X1 port map( A1 => n35231, A2 => n19749, Z => n16458);
   U30421 : XOR2_X1 port map( A1 => n32309, A2 => n7481, Z => n36851);
   U30427 : OAI21_X2 port map( A1 => n26640, A2 => n26918, B => n36853, ZN => 
                           n5554);
   U30428 : NAND2_X1 port map( A1 => n11700, A2 => n13786, ZN => n13363);
   U30438 : NAND2_X2 port map( A1 => n12379, A2 => n12378, ZN => n12989);
   U30442 : OR2_X1 port map( A1 => n25991, A2 => n25760, Z => n33328);
   U30446 : INV_X2 port map( I => n36856, ZN => n31557);
   U30450 : XOR2_X1 port map( A1 => n4334, A2 => n4332, Z => n36856);
   U30457 : XOR2_X1 port map( A1 => n2739, A2 => n2738, Z => n9022);
   U30458 : NAND2_X1 port map( A1 => n550, A2 => n18415, ZN => n6499);
   U30459 : NOR3_X1 port map( A1 => n23042, A2 => n39096, A3 => n33431, ZN => 
                           n14882);
   U30462 : XOR2_X1 port map( A1 => n18051, A2 => n6523, Z => n26500);
   U30463 : NAND2_X2 port map( A1 => n5705, A2 => n16063, ZN => n31015);
   U30465 : NAND2_X2 port map( A1 => n21732, A2 => n11124, ZN => n17126);
   U30466 : NAND2_X2 port map( A1 => n33148, A2 => n21730, ZN => n21732);
   U30467 : OAI22_X2 port map( A1 => n20813, A2 => n1512, B1 => n10015, B2 => 
                           n26215, ZN => n26038);
   U30468 : OAI22_X2 port map( A1 => n12826, A2 => n17183, B1 => n31843, B2 => 
                           n31842, ZN => n26215);
   U30474 : XOR2_X1 port map( A1 => n27730, A2 => n9164, Z => n36861);
   U30487 : XOR2_X1 port map( A1 => n25080, A2 => n25196, Z => n25286);
   U30495 : XOR2_X1 port map( A1 => n33027, A2 => n26338, Z => n26450);
   U30497 : AOI21_X2 port map( A1 => n26053, A2 => n926, B => n34153, ZN => 
                           n2751);
   U30498 : INV_X2 port map( I => n36868, ZN => n13686);
   U30499 : XOR2_X1 port map( A1 => n10485, A2 => n25289, Z => n10484);
   U30512 : INV_X4 port map( I => n36871, ZN => n23531);
   U30513 : OAI22_X2 port map( A1 => n23206, A2 => n36422, B1 => n23207, B2 => 
                           n14994, ZN => n36871);
   U30515 : XOR2_X1 port map( A1 => n26358, A2 => n32386, Z => n33385);
   U30522 : INV_X1 port map( I => n21617, ZN => n37033);
   U30540 : AOI22_X1 port map( A1 => n122, A2 => n36910, B1 => n29218, B2 => 
                           n12691, ZN => n33350);
   U30549 : NAND2_X2 port map( A1 => n5258, A2 => n23523, ZN => n23526);
   U30552 : XOR2_X1 port map( A1 => n36880, A2 => n15398, Z => n32154);
   U30558 : INV_X1 port map( I => n13374, ZN => n1469);
   U30559 : XNOR2_X1 port map( A1 => n13374, A2 => n27787, ZN => n27748);
   U30563 : NAND2_X2 port map( A1 => n18586, A2 => n15979, ZN => n27358);
   U30565 : XOR2_X1 port map( A1 => n5587, A2 => n36884, Z => n29769);
   U30566 : XOR2_X1 port map( A1 => n22758, A2 => n9205, Z => n3529);
   U30580 : XOR2_X1 port map( A1 => n10317, A2 => n10546, Z => n10316);
   U30581 : INV_X4 port map( I => n36889, ZN => n9231);
   U30586 : INV_X2 port map( I => n36890, ZN => n30484);
   U30587 : XOR2_X1 port map( A1 => n4967, A2 => n5743, Z => n36890);
   U30600 : OAI21_X2 port map( A1 => n24326, A2 => n13884, B => n24390, ZN => 
                           n36891);
   U30601 : OR2_X2 port map( A1 => n21395, A2 => n21394, Z => n17869);
   U30602 : OR2_X1 port map( A1 => n25540, A2 => n30317, Z => n16825);
   U30603 : NOR2_X2 port map( A1 => n17800, A2 => n11614, ZN => n36892);
   U30604 : NAND2_X1 port map( A1 => n253, A2 => n30494, ZN => n16884);
   U30609 : XOR2_X1 port map( A1 => n17461, A2 => n36899, Z => n22854);
   U30610 : XOR2_X1 port map( A1 => n10939, A2 => n2234, Z => n36899);
   U30612 : AOI22_X2 port map( A1 => n23090, A2 => n19488, B1 => n15163, B2 => 
                           n23091, ZN => n32025);
   U30615 : XOR2_X1 port map( A1 => n8068, A2 => n8065, Z => n8539);
   U30619 : OR2_X1 port map( A1 => n24536, A2 => n33946, Z => n25680);
   U30620 : XOR2_X1 port map( A1 => n38905, A2 => n23914, Z => n30502);
   U30623 : NAND3_X1 port map( A1 => n37010, A2 => n39133, A3 => n15941, ZN => 
                           n6521);
   U30627 : INV_X2 port map( I => n36909, ZN => n18959);
   U30628 : XOR2_X1 port map( A1 => Plaintext(175), A2 => Key(175), Z => n36909
                           );
   U30629 : INV_X2 port map( I => n33581, ZN => n12435);
   U30635 : XOR2_X1 port map( A1 => n37855, A2 => n10131, Z => n36916);
   U30636 : NOR2_X1 port map( A1 => n32696, A2 => n3605, ZN => n32695);
   U30640 : XOR2_X1 port map( A1 => n36919, A2 => n19799, Z => Ciphertext(86));
   U30641 : OR2_X1 port map( A1 => n26058, A2 => n38416, Z => n14573);
   U30642 : OAI21_X2 port map( A1 => n34065, A2 => n12353, B => n36923, ZN => 
                           n21300);
   U30643 : NAND2_X2 port map( A1 => n9394, A2 => n5414, ZN => n36924);
   U30645 : INV_X2 port map( I => n28790, ZN => n7288);
   U30646 : XOR2_X1 port map( A1 => n6795, A2 => n36925, Z => n6796);
   U30647 : XOR2_X1 port map( A1 => n38816, A2 => n6847, Z => n36925);
   U30648 : NAND3_X1 port map( A1 => n30931, A2 => n18960, A3 => n28653, ZN => 
                           n4523);
   U30649 : XOR2_X1 port map( A1 => n22772, A2 => n11315, Z => n11314);
   U30650 : XOR2_X1 port map( A1 => n25313, A2 => n25312, Z => n4273);
   U30651 : AOI22_X2 port map( A1 => n7897, A2 => n36926, B1 => n8519, B2 => 
                           n7896, ZN => n7895);
   U30652 : NAND2_X2 port map( A1 => n1328, A2 => n22287, ZN => n36926);
   U30655 : NOR2_X2 port map( A1 => n36930, A2 => n17544, ZN => n11568);
   U30657 : INV_X2 port map( I => n36932, ZN => n6327);
   U30661 : XOR2_X1 port map( A1 => n8400, A2 => n6360, Z => n11451);
   U30662 : NAND2_X2 port map( A1 => n3352, A2 => n2771, ZN => n23069);
   U30664 : OAI21_X2 port map( A1 => n36938, A2 => n31277, B => n15251, ZN => 
                           n27424);
   U30666 : OAI22_X2 port map( A1 => n34077, A2 => n7440, B1 => n2439, B2 => 
                           n1031, ZN => n23942);
   U30669 : NAND2_X1 port map( A1 => n33894, A2 => n33609, ZN => n23341);
   U30671 : AOI21_X2 port map( A1 => n14203, A2 => n14205, B => n24185, ZN => 
                           n17351);
   U30672 : NAND2_X2 port map( A1 => n6303, A2 => n23484, ZN => n23306);
   U30674 : NOR2_X1 port map( A1 => n9751, A2 => n19746, ZN => n36940);
   U30675 : NOR2_X2 port map( A1 => n26727, A2 => n13588, ZN => n26774);
   U30676 : OAI21_X2 port map( A1 => n14966, A2 => n1489, B => n36942, ZN => 
                           n14949);
   U30678 : INV_X1 port map( I => n28848, ZN => n1178);
   U30682 : NOR2_X1 port map( A1 => n4318, A2 => n22225, ZN => n36946);
   U30685 : OAI22_X1 port map( A1 => n21837, A2 => n8736, B1 => n690, B2 => 
                           n21435, ZN => n14909);
   U30689 : NAND2_X1 port map( A1 => n28562, A2 => n28563, ZN => n28564);
   U30690 : NAND2_X2 port map( A1 => n10640, A2 => n13484, ZN => n6384);
   U30693 : XOR2_X1 port map( A1 => n36959, A2 => n10748, Z => n15883);
   U30695 : XOR2_X1 port map( A1 => n29056, A2 => n29028, Z => n12039);
   U30696 : NOR2_X2 port map( A1 => n21370, A2 => n21369, ZN => n31573);
   U30697 : XOR2_X1 port map( A1 => n26473, A2 => n26472, Z => n36961);
   U30698 : NOR2_X2 port map( A1 => n4849, A2 => n344, ZN => n20289);
   U30699 : XOR2_X1 port map( A1 => n36962, A2 => n12228, Z => n33144);
   U30703 : AND2_X1 port map( A1 => n20660, A2 => n14453, Z => n15668);
   U30704 : XOR2_X1 port map( A1 => n27809, A2 => n10983, Z => n10982);
   U30709 : OAI21_X2 port map( A1 => n3012, A2 => n7075, B => n36967, ZN => 
                           n7901);
   U30710 : XOR2_X1 port map( A1 => n31581, A2 => n23660, Z => n8512);
   U30713 : OAI22_X1 port map( A1 => n6851, A2 => n29421, B1 => n20018, B2 => 
                           n32946, ZN => n36968);
   U30715 : XOR2_X1 port map( A1 => n12411, A2 => n26145, Z => n5737);
   U30718 : XNOR2_X1 port map( A1 => n27855, A2 => n27607, ZN => n27732);
   U30719 : NAND2_X2 port map( A1 => n15772, A2 => n27453, ZN => n27855);
   U30720 : NOR2_X1 port map( A1 => n4116, A2 => n7935, ZN => n21723);
   U30723 : NAND2_X2 port map( A1 => n8595, A2 => n36974, ZN => n3313);
   U30724 : NOR3_X1 port map( A1 => n37378, A2 => n17791, A3 => n36798, ZN => 
                           n15831);
   U30727 : NAND2_X2 port map( A1 => n27068, A2 => n15120, ZN => n27864);
   U30730 : XOR2_X1 port map( A1 => n33132, A2 => n35900, Z => n36980);
   U30734 : NAND2_X2 port map( A1 => n36985, A2 => n18098, ZN => n2);
   U30735 : NAND2_X2 port map( A1 => n15015, A2 => n31194, ZN => n36985);
   U30736 : NAND2_X2 port map( A1 => n29270, A2 => n29271, ZN => n19085);
   U30738 : NAND2_X1 port map( A1 => n36216, A2 => n10104, ZN => n13467);
   U30744 : XOR2_X1 port map( A1 => n26393, A2 => n20212, Z => n12622);
   U30745 : AOI22_X2 port map( A1 => n29461, A2 => n29389, B1 => n17426, B2 => 
                           n19151, ZN => n29402);
   U30748 : XOR2_X1 port map( A1 => n17653, A2 => n31112, Z => n24836);
   U30749 : INV_X2 port map( I => n24928, ZN => n31112);
   U30750 : AOI22_X2 port map( A1 => n24834, A2 => n1271, B1 => n24866, B2 => 
                           n13220, ZN => n24928);
   U30751 : OAI21_X1 port map( A1 => n3792, A2 => n3793, B => n24733, ZN => 
                           n4063);
   U30755 : NAND2_X2 port map( A1 => n33929, A2 => n21424, ZN => n4179);
   U30757 : OAI21_X2 port map( A1 => n2668, A2 => n2671, B => n9341, ZN => 
                           n22443);
   U30758 : NAND3_X2 port map( A1 => n32196, A2 => n1529, A3 => n35333, ZN => 
                           n26218);
   U30760 : NAND3_X1 port map( A1 => n29673, A2 => n19497, A3 => n20672, ZN => 
                           n18944);
   U30762 : NAND2_X1 port map( A1 => n16838, A2 => n1387, ZN => n18431);
   U30766 : BUF_X2 port map( I => n22943, Z => n36996);
   U30767 : NOR2_X1 port map( A1 => n36998, A2 => n36997, ZN => n16837);
   U30768 : INV_X1 port map( I => n8399, ZN => n36998);
   U30769 : XOR2_X1 port map( A1 => n33308, A2 => n31791, Z => n36999);
   U30773 : NOR2_X1 port map( A1 => n459, A2 => n1483, ZN => n37002);
   U30774 : INV_X2 port map( I => n37003, ZN => n6106);
   U30775 : XOR2_X1 port map( A1 => n6109, A2 => n6107, Z => n37003);
   U30777 : NAND2_X1 port map( A1 => n2981, A2 => n2983, ZN => n37006);
   U30778 : OR2_X2 port map( A1 => n20897, A2 => n19167, Z => n23121);
   U30779 : NAND2_X2 port map( A1 => n37007, A2 => n25967, ZN => n26516);
   U30780 : NOR2_X1 port map( A1 => n25964, A2 => n25962, ZN => n37008);
   U30782 : NAND2_X2 port map( A1 => n528, A2 => n530, ZN => n9611);
   U30783 : AOI22_X2 port map( A1 => n27287, A2 => n27218, B1 => n31146, B2 => 
                           n30486, ZN => n27564);
   U30784 : OAI21_X2 port map( A1 => n34359, A2 => n1470, B => n6013, ZN => 
                           n27287);
   U30787 : NOR2_X1 port map( A1 => n1297, A2 => n23468, ZN => n37012);
   U30788 : INV_X2 port map( I => n37013, ZN => n20616);
   U30789 : XNOR2_X1 port map( A1 => n4140, A2 => n4141, ZN => n37013);
   U30791 : NAND2_X2 port map( A1 => n24571, A2 => n37017, ZN => n13200);
   U30792 : AND2_X1 port map( A1 => n3389, A2 => n37018, Z => n5535);
   U30793 : XOR2_X1 port map( A1 => n16833, A2 => n37019, Z => n331);
   U30794 : XOR2_X1 port map( A1 => n8704, A2 => n23980, Z => n37019);
   U30795 : INV_X2 port map( I => n37020, ZN => n37056);
   U30796 : XOR2_X1 port map( A1 => n2757, A2 => n2758, Z => n37020);
   U30798 : XOR2_X1 port map( A1 => n30966, A2 => n14043, Z => n14045);
   U30804 : AOI21_X2 port map( A1 => n37026, A2 => n14082, B => n7097, ZN => 
                           n26086);
   U30805 : OR2_X1 port map( A1 => n14257, A2 => n25642, Z => n37026);
   U30808 : INV_X2 port map( I => n20616, ZN => n32894);
   U30809 : NAND2_X2 port map( A1 => n37027, A2 => n9313, ZN => n9290);
   U30810 : OAI21_X2 port map( A1 => n30369, A2 => n10236, B => n18603, ZN => 
                           n37027);
   U30815 : NAND3_X2 port map( A1 => n13858, A2 => n13859, A3 => n13855, ZN => 
                           n37030);
   U30816 : OR3_X1 port map( A1 => n38159, A2 => n17751, A3 => n8944, Z => 
                           n9745);
   U30824 : NAND3_X2 port map( A1 => n14994, A2 => n14409, A3 => n31300, ZN => 
                           n31918);
   U30825 : NAND2_X2 port map( A1 => n20831, A2 => n21552, ZN => n22349);
   U30830 : XOR2_X1 port map( A1 => n37034, A2 => n12918, Z => n9973);
   U30833 : NAND2_X2 port map( A1 => n37036, A2 => n18822, ZN => n18819);
   U30834 : OAI22_X2 port map( A1 => n32740, A2 => n14994, B1 => n13946, B2 => 
                           n14439, ZN => n37036);
   U30838 : XOR2_X1 port map( A1 => n10837, A2 => n37038, Z => n37037);
   U30840 : XOR2_X1 port map( A1 => n5317, A2 => n5318, Z => n12829);
   U30842 : OAI21_X2 port map( A1 => n32837, A2 => n30288, B => n27182, ZN => 
                           n27746);
   U30843 : XOR2_X1 port map( A1 => n11059, A2 => n10593, Z => n10592);
   U30845 : NOR2_X1 port map( A1 => n37039, A2 => n7175, ZN => n19563);
   U30846 : BUF_X2 port map( I => n27417, Z => n37040);
   U30847 : BUF_X2 port map( I => n7560, Z => n37042);
   U30848 : XOR2_X1 port map( A1 => n22517, A2 => n37660, Z => n1868);
   U30849 : INV_X2 port map( I => n35469, ZN => n274);
   U30850 : INV_X2 port map( I => n32191, ZN => n1082);
   U30853 : INV_X2 port map( I => n32838, ZN => n10659);
   U30854 : INV_X2 port map( I => n24316, ZN => n24467);
   U30855 : XOR2_X1 port map( A1 => n2107, A2 => n2104, Z => n37047);
   U30857 : OAI21_X2 port map( A1 => n13340, A2 => n32019, B => n17453, ZN => 
                           n31579);
   U30858 : OAI22_X2 port map( A1 => n2746, A2 => n37202, B1 => n16541, B2 => 
                           n2745, ZN => n31543);
   U30859 : XOR2_X1 port map( A1 => n12830, A2 => n12833, Z => n37048);
   U30863 : INV_X2 port map( I => n13877, ZN => n12999);
   U30867 : INV_X1 port map( I => n29210, ZN => n17121);
   U30868 : OAI21_X2 port map( A1 => n15141, A2 => n15139, B => n15138, ZN => 
                           n29802);
   U241 : NAND2_X2 port map( A1 => n2, A2 => n5543, ZN => n6317);
   U5878 : INV_X2 port map( I => n8253, ZN => n8385);
   U1627 : INV_X2 port map( I => n8173, ZN => n32619);
   U7284 : INV_X2 port map( I => n668, ZN => n21910);
   U4261 : NAND2_X2 port map( A1 => n17118, A2 => n22177, ZN => n22137);
   U59 : INV_X2 port map( I => n10118, ZN => n1052);
   U20202 : NAND2_X2 port map( A1 => n27266, A2 => n35990, ZN => n20403);
   U1704 : OAI21_X2 port map( A1 => n959, A2 => n33712, B => n18238, ZN => 
                           n33354);
   U5464 : NAND2_X2 port map( A1 => n16579, A2 => n1843, ZN => n1842);
   U2347 : NAND2_X2 port map( A1 => n38629, A2 => n1419, ZN => n28682);
   U6509 : INV_X2 port map( I => n22359, ZN => n36337);
   U10258 : INV_X2 port map( I => n18429, ZN => n4318);
   U23027 : INV_X2 port map( I => n20995, ZN => n17047);
   U967 : BUF_X4 port map( I => n18983, Z => n12159);
   U17487 : OAI22_X2 port map( A1 => n2842, A2 => n2841, B1 => n1671, B2 => 
                           n22182, ZN => n1745);
   U5236 : INV_X2 port map( I => n22897, ZN => n1654);
   U12157 : NAND2_X2 port map( A1 => n7724, A2 => n26134, ZN => n3244);
   U5990 : NAND2_X2 port map( A1 => n35779, A2 => n19053, ZN => n12067);
   U7621 : INV_X2 port map( I => n30131, ZN => n30144);
   U2525 : NAND2_X2 port map( A1 => n36960, A2 => n35780, ZN => n17813);
   U6787 : INV_X2 port map( I => n6291, ZN => n5802);
   U6080 : BUF_X4 port map( I => n24140, Z => n2439);
   U1379 : INV_X4 port map( I => n25867, ZN => n5886);
   U2394 : NAND2_X2 port map( A1 => n14130, A2 => n34013, ZN => n22959);
   U17116 : INV_X2 port map( I => n24515, ZN => n1270);
   U22586 : INV_X2 port map( I => n10679, ZN => n29960);
   U10169 : OAI21_X2 port map( A1 => n1778, A2 => n14028, B => n14038, ZN => 
                           n1777);
   U1092 : INV_X2 port map( I => n37593, ZN => n34513);
   U6911 : INV_X4 port map( I => n14472, ZN => n8070);
   U4968 : INV_X2 port map( I => n36913, ZN => n7088);
   U5911 : INV_X2 port map( I => n26796, ZN => n26734);
   U28603 : NAND3_X2 port map( A1 => n978, A2 => n13508, A3 => n33100, ZN => 
                           n12604);
   U2367 : OAI21_X2 port map( A1 => n14130, A2 => n34013, B => n17691, ZN => 
                           n34715);
   U8654 : NAND2_X2 port map( A1 => n20579, A2 => n20581, ZN => n21980);
   U1610 : NOR2_X2 port map( A1 => n12460, A2 => n31712, ZN => n31711);
   U3407 : AOI21_X2 port map( A1 => n27883, A2 => n28255, B => n27885, ZN => 
                           n10151);
   U20427 : INV_X2 port map( I => n7674, ZN => n20372);
   U3791 : BUF_X4 port map( I => n6106, Z => n32105);
   U17987 : NAND2_X2 port map( A1 => n22402, A2 => n22183, ZN => n22398);
   U28416 : NAND2_X2 port map( A1 => n35429, A2 => n1047, ZN => n22183);
   U6937 : INV_X2 port map( I => n20614, ZN => n18831);
   U16853 : INV_X4 port map( I => n1276, ZN => n24336);
   U326 : INV_X2 port map( I => n28250, ZN => n13457);
   U861 : NAND2_X2 port map( A1 => n20094, A2 => n26831, ZN => n36507);
   U4971 : NOR2_X2 port map( A1 => n13502, A2 => n19889, ZN => n13501);
   U23874 : INV_X2 port map( I => n35901, ZN => n15664);
   U2138 : INV_X2 port map( I => n23967, ZN => n34451);
   U7170 : INV_X4 port map( I => n22935, ZN => n1042);
   U4267 : BUF_X2 port map( I => n13989, Z => n33516);
   U15517 : INV_X2 port map( I => n7810, ZN => n8127);
   U2172 : NAND2_X2 port map( A1 => n25337, A2 => n20052, ZN => n25550);
   U18960 : INV_X2 port map( I => n6550, ZN => n28159);
   U1338 : INV_X2 port map( I => n2047, ZN => n1143);
   U17145 : INV_X2 port map( I => n29672, ZN => n20672);
   U3603 : NAND2_X2 port map( A1 => n1072, A2 => n34008, ZN => n28108);
   U1687 : NOR2_X2 port map( A1 => n3451, A2 => n25359, ZN => n31900);
   U7601 : OAI21_X2 port map( A1 => n29990, A2 => n3986, B => n621, ZN => n4011
                           );
   U1206 : NAND2_X2 port map( A1 => n19889, A2 => n11003, ZN => n4852);
   U7206 : NAND2_X2 port map( A1 => n26761, A2 => n26809, ZN => n26653);
   U22538 : OAI21_X2 port map( A1 => n19261, A2 => n22137, B => n35802, ZN => 
                           n5874);
   U589 : INV_X4 port map( I => n14408, ZN => n1493);
   U3542 : INV_X2 port map( I => n23404, ZN => n3366);
   U6276 : BUF_X2 port map( I => n13704, Z => n35505);
   U302 : INV_X2 port map( I => n16108, ZN => n15112);
   U359 : NAND2_X2 port map( A1 => n28281, A2 => n37754, ZN => n11280);
   U20032 : INV_X2 port map( I => n32010, ZN => n33937);
   U28095 : INV_X2 port map( I => n27745, ZN => n27535);
   U7386 : NAND2_X2 port map( A1 => n9217, A2 => n13495, ZN => n6409);
   U5213 : BUF_X4 port map( I => n2319, Z => n35062);
   U18781 : INV_X2 port map( I => n5960, ZN => n9147);
   U729 : NAND2_X2 port map( A1 => n26870, A2 => n7973, ZN => n27007);
   U18464 : OAI21_X2 port map( A1 => n12146, A2 => n10008, B => n33104, ZN => 
                           n31759);
   U141 : INV_X2 port map( I => n34179, ZN => n30052);
   U653 : INV_X2 port map( I => n4815, ZN => n21149);
   U29506 : NAND2_X2 port map( A1 => n7635, A2 => n28023, ZN => n27918);
   U5757 : INV_X4 port map( I => n11003, ZN => n927);
   U3026 : INV_X2 port map( I => n17529, ZN => n1671);
   U30812 : INV_X4 port map( I => n31994, ZN => n37028);
   U3834 : INV_X2 port map( I => n34526, ZN => n24708);
   U5877 : INV_X2 port map( I => n16627, ZN => n35722);
   U18045 : AOI22_X2 port map( A1 => n17309, A2 => n32385, B1 => n11980, B2 => 
                           n38694, ZN => n35212);
   U3923 : INV_X2 port map( I => n24317, ZN => n17546);
   U13744 : INV_X2 port map( I => n692, ZN => n25999);
   U11009 : NOR2_X1 port map( A1 => n32497, A2 => n35720, ZN => n18218);
   U5270 : INV_X2 port map( I => n24285, ZN => n24119);
   U6679 : INV_X4 port map( I => n22682, ZN => n22856);
   U1384 : BUF_X4 port map( I => n18987, Z => n596);
   U9089 : NOR2_X2 port map( A1 => n33669, A2 => n39132, ZN => n2614);
   U2391 : NOR2_X2 port map( A1 => n1045, A2 => n20173, ZN => n35863);
   U5605 : BUF_X4 port map( I => n12667, Z => n6131);
   U4655 : INV_X2 port map( I => n9165, ZN => n10681);
   U5742 : NAND2_X2 port map( A1 => n27011, A2 => n31875, ZN => n10357);
   U28849 : NAND2_X1 port map( A1 => n4239, A2 => n22390, ZN => n36616);
   U22096 : INV_X2 port map( I => n9958, ZN => n12302);
   U2254 : INV_X4 port map( I => n11033, ZN => n930);
   U3343 : INV_X4 port map( I => n217, ZN => n5702);
   U7714 : BUF_X2 port map( I => n3014, Z => n33841);
   U22616 : NOR2_X2 port map( A1 => n32542, A2 => n20732, ZN => n8925);
   U2242 : NOR2_X2 port map( A1 => n217, A2 => n7160, ZN => n22932);
   U19626 : INV_X2 port map( I => n7133, ZN => n26244);
   U2369 : INV_X2 port map( I => n25337, ZN => n25460);
   U10213 : NOR2_X1 port map( A1 => n16432, A2 => n34382, ZN => n6104);
   U6587 : OAI21_X2 port map( A1 => n38555, A2 => n31383, B => n21995, ZN => 
                           n20089);
   U1721 : NOR2_X2 port map( A1 => n31698, A2 => n18148, ZN => n20038);
   U1080 : NOR2_X2 port map( A1 => n26056, A2 => n9743, ZN => n15703);
   U17473 : OAI22_X2 port map( A1 => n39576, A2 => n16468, B1 => n1057, B2 => 
                           n30051, ZN => n7166);
   U3191 : NAND2_X2 port map( A1 => n9363, A2 => n24707, ZN => n34192);
   U12702 : NOR2_X2 port map( A1 => n33986, A2 => n34526, ZN => n9363);
   U12056 : NAND2_X2 port map( A1 => n9326, A2 => n19241, ZN => n1849);
   U5051 : NOR2_X2 port map( A1 => n37072, A2 => n39454, ZN => n9326);
   U652 : INV_X2 port map( I => n8402, ZN => n8302);
   U28451 : INV_X4 port map( I => n34562, ZN => n33369);
   U12405 : NOR2_X2 port map( A1 => n6894, A2 => n560, ZN => n21136);
   U650 : INV_X2 port map( I => n27825, ZN => n1463);
   U238 : NAND2_X2 port map( A1 => n10587, A2 => n9648, ZN => n33724);
   U5564 : OAI21_X2 port map( A1 => n20134, A2 => n20612, B => n34417, ZN => 
                           n16643);
   U4895 : NAND2_X2 port map( A1 => n19546, A2 => n32138, ZN => n12751);
   U17390 : INV_X2 port map( I => n5921, ZN => n17708);
   U5702 : NOR2_X2 port map( A1 => n39085, A2 => n1027, ZN => n11199);
   U2048 : INV_X2 port map( I => n690, ZN => n1158);
   U4150 : BUF_X4 port map( I => n8742, Z => n557);
   U17960 : AOI22_X2 port map( A1 => n21449, A2 => n1342, B1 => n32817, B2 => 
                           n22173, ZN => n21453);
   U2310 : NOR2_X2 port map( A1 => n12946, A2 => n20696, ZN => n31123);
   U3897 : OR2_X1 port map( A1 => n10896, A2 => n31596, Z => n10870);
   U16641 : NAND2_X2 port map( A1 => n28238, A2 => n1453, ZN => n4150);
   U17288 : INV_X2 port map( I => n16054, ZN => n3395);
   U8624 : NAND2_X2 port map( A1 => n9242, A2 => n31971, ZN => n2604);
   U1120 : NOR2_X2 port map( A1 => n32157, A2 => n32156, ZN => n34883);
   U18281 : NAND2_X2 port map( A1 => n18062, A2 => n25801, ZN => n25903);
   U17589 : INV_X2 port map( I => n30894, ZN => n89);
   U17232 : NAND2_X2 port map( A1 => n29986, A2 => n16468, ZN => n6602);
   U6855 : NAND2_X2 port map( A1 => n24337, A2 => n14558, ZN => n7811);
   U600 : INV_X2 port map( I => n27730, ZN => n27833);
   U17064 : AND2_X2 port map( A1 => n889, A2 => n13492, Z => n14642);
   U3387 : BUF_X2 port map( I => n17425, Z => n15089);
   U3233 : INV_X2 port map( I => n19260, ZN => n29525);
   U2112 : INV_X2 port map( I => n36272, ZN => n14558);
   U464 : AOI21_X2 port map( A1 => n35846, A2 => n16851, B => n4152, ZN => 
                           n12466);
   U19587 : NOR2_X2 port map( A1 => n1650, A2 => n9472, ZN => n5215);
   U3424 : NAND2_X2 port map( A1 => n6161, A2 => n32617, ZN => n6732);
   U5846 : INV_X4 port map( I => n25498, ZN => n25379);
   U18651 : AOI21_X2 port map( A1 => n21996, A2 => n3687, B => n22071, ZN => 
                           n16028);
   U7232 : INV_X4 port map( I => n11149, ZN => n22267);
   U1888 : INV_X4 port map( I => n6944, ZN => n24723);
   U26225 : INV_X2 port map( I => n32080, ZN => n20572);
   U1256 : NAND2_X2 port map( A1 => n37151, A2 => n26008, ZN => n20049);
   U9258 : OAI21_X2 port map( A1 => n3224, A2 => n11130, B => n33858, ZN => 
                           n3095);
   U5583 : INV_X4 port map( I => n29598, ZN => n1404);
   U7182 : INV_X2 port map( I => n57, ZN => n14304);
   U5821 : INV_X4 port map( I => n32617, ZN => n21762);
   U13678 : NAND2_X2 port map( A1 => n17635, A2 => n22107, ZN => n17634);
   U4236 : AOI21_X2 port map( A1 => n15715, A2 => n33061, B => n38527, ZN => 
                           n15713);
   U13781 : INV_X2 port map( I => n7768, ZN => n8621);
   U8954 : INV_X4 port map( I => n33384, ZN => n30694);
   U4001 : AND2_X1 port map( A1 => n11562, A2 => n26269, Z => n854);
   U24461 : OAI21_X2 port map( A1 => n18734, A2 => n4664, B => n32419, ZN => 
                           n16809);
   U6750 : NOR2_X2 port map( A1 => n23528, A2 => n36539, ZN => n23529);
   U4277 : INV_X2 port map( I => n24337, ZN => n8174);
   U608 : INV_X2 port map( I => n28219, ZN => n36860);
   U11367 : INV_X2 port map( I => n28141, ZN => n28142);
   U4175 : INV_X2 port map( I => n14463, ZN => n10477);
   U1717 : INV_X2 port map( I => n25194, ZN => n2318);
   U3806 : INV_X2 port map( I => n3313, ZN => n992);
   U9200 : INV_X1 port map( I => n1472, ZN => n3088);
   U18104 : AOI21_X2 port map( A1 => n31680, A2 => n16480, B => n16479, ZN => 
                           n6110);
   U10313 : AOI22_X1 port map( A1 => n21756, A2 => n11916, B1 => n11917, B2 => 
                           n11918, ZN => n10324);
   U9128 : INV_X2 port map( I => n28153, ZN => n1203);
   U177 : INV_X2 port map( I => n29642, ZN => n35571);
   U12780 : INV_X1 port map( I => n16502, ZN => n1581);
   U2120 : INV_X4 port map( I => n1589, ZN => n2396);
   U3264 : NAND2_X2 port map( A1 => n29981, A2 => n29968, ZN => n29971);
   U6363 : INV_X2 port map( I => n20408, ZN => n5907);
   U4208 : BUF_X4 port map( I => n28807, Z => n33577);
   U1099 : INV_X2 port map( I => n801, ZN => n24267);
   U6925 : AOI22_X2 port map( A1 => n24084, A2 => n24853, B1 => n24855, B2 => 
                           n32064, ZN => n24085);
   U5747 : INV_X2 port map( I => n23464, ZN => n23238);
   U17203 : NAND2_X2 port map( A1 => n35960, A2 => n24637, ZN => n20414);
   U13900 : OAI22_X2 port map( A1 => n21605, A2 => n16128, B1 => n21944, B2 => 
                           n19133, ZN => n11302);
   U2363 : AOI22_X2 port map( A1 => n22863, A2 => n1650, B1 => n1651, B2 => 
                           n6385, ZN => n4160);
   U79 : INV_X2 port map( I => n31428, ZN => n3693);
   U857 : AOI21_X2 port map( A1 => n17785, A2 => n11513, B => n35877, ZN => 
                           n36520);
   U1736 : OAI21_X2 port map( A1 => n11271, A2 => n37106, B => n11082, ZN => 
                           n13494);
   U14416 : NOR2_X2 port map( A1 => n37137, A2 => n20625, ZN => n31465);
   U14439 : NOR2_X2 port map( A1 => n948, A2 => n26660, ZN => n31264);
   U3419 : INV_X4 port map( I => n35377, ZN => n21130);
   U11532 : INV_X2 port map( I => n30959, ZN => n28168);
   U6368 : INV_X2 port map( I => n8765, ZN => n962);
   U2518 : INV_X2 port map( I => n22335, ZN => n36632);
   U27619 : INV_X2 port map( I => n19458, ZN => n29998);
   U21142 : NOR2_X2 port map( A1 => n8818, A2 => n18261, ZN => n28111);
   U9685 : NAND2_X2 port map( A1 => n9584, A2 => n34620, ZN => n9580);
   U5741 : BUF_X4 port map( I => n5126, Z => n31827);
   U1604 : OAI21_X2 port map( A1 => n4625, A2 => n2149, B => n34636, ZN => 
                           n7695);
   U3466 : INV_X4 port map( I => n1275, ZN => n9101);
   U10220 : OAI22_X1 port map( A1 => n22889, A2 => n19469, B1 => n5656, B2 => 
                           n23125, ZN => n34713);
   U676 : INV_X2 port map( I => n27595, ZN => n31163);
   U1432 : NAND2_X2 port map( A1 => n1048, A2 => n22108, ZN => n22107);
   U203 : INV_X2 port map( I => n20006, ZN => n11721);
   U1615 : NOR2_X2 port map( A1 => n25327, A2 => n37237, ZN => n18786);
   U18361 : NAND2_X2 port map( A1 => n32902, A2 => n28377, ZN => n9111);
   U6087 : CLKBUF_X4 port map( I => n23992, Z => n24443);
   U15189 : INV_X2 port map( I => n13193, ZN => n24018);
   U5798 : INV_X2 port map( I => n22122, ZN => n22266);
   U6996 : AOI21_X2 port map( A1 => n2057, A2 => n7210, B => n20989, ZN => 
                           n20988);
   U2922 : AOI22_X2 port map( A1 => n38851, A2 => n19538, B1 => n1314, B2 => 
                           n14725, ZN => n33706);
   U1628 : NAND2_X2 port map( A1 => n37238, A2 => n5798, ZN => n34636);
   U7856 : INV_X4 port map( I => n2532, ZN => n21751);
   U13217 : INV_X2 port map( I => n23365, ZN => n1953);
   U11385 : INV_X2 port map( I => n35895, ZN => n32961);
   U20655 : INV_X2 port map( I => n32151, ZN => n3969);
   U8715 : INV_X4 port map( I => n18205, ZN => n21788);
   U4466 : NOR2_X2 port map( A1 => n27326, A2 => n39216, ZN => n8763);
   U4911 : INV_X4 port map( I => n12443, ZN => n28103);
   U4215 : NAND2_X2 port map( A1 => n7552, A2 => n39681, ZN => n11126);
   U3875 : OR2_X1 port map( A1 => n31558, A2 => n7584, Z => n23161);
   U3133 : INV_X2 port map( I => n20372, ZN => n23082);
   U13650 : OAI21_X2 port map( A1 => n37189, A2 => n14823, B => n9715, ZN => 
                           n14822);
   U13530 : NOR2_X2 port map( A1 => n35586, A2 => n19870, ZN => n4099);
   U27421 : OAI21_X2 port map( A1 => n1625, A2 => n6217, B => n23528, ZN => 
                           n23283);
   U877 : INV_X4 port map( I => n21254, ZN => n954);
   U2106 : OAI21_X2 port map( A1 => n4993, A2 => n19837, B => n18163, ZN => 
                           n33487);
   U7027 : NAND2_X2 port map( A1 => n955, A2 => n15541, ZN => n25452);
   U15586 : INV_X2 port map( I => n24427, ZN => n19070);
   U7035 : OAI21_X2 port map( A1 => n32085, A2 => n560, B => n17353, ZN => 
                           n5355);
   U1055 : AND2_X2 port map( A1 => n36283, A2 => n12682, Z => n26955);
   U3812 : INV_X2 port map( I => n20087, ZN => n344);
   U6938 : INV_X2 port map( I => n6106, ZN => n14708);
   U2233 : NAND2_X2 port map( A1 => n35545, A2 => n39316, ZN => n9011);
   U6128 : INV_X2 port map( I => n3779, ZN => n4152);
   U2968 : OAI22_X2 port map( A1 => n6181, A2 => n1390, B1 => n29662, B2 => 
                           n39689, ZN => n29665);
   U2523 : OAI21_X2 port map( A1 => n5945, A2 => n1989, B => n5944, ZN => n4328
                           );
   U6300 : INV_X2 port map( I => n22038, ZN => n34216);
   U344 : INV_X2 port map( I => n28717, ZN => n35491);
   U25211 : INV_X2 port map( I => n25557, ZN => n17281);
   U7051 : OAI21_X2 port map( A1 => n38531, A2 => n31310, B => n1524, ZN => 
                           n35956);
   U51 : NOR2_X2 port map( A1 => n3818, A2 => n30076, ZN => n30066);
   U29543 : AOI22_X2 port map( A1 => n6534, A2 => n36911, B1 => n39632, B2 => 
                           n7542, ZN => n3920);
   U3384 : NOR2_X2 port map( A1 => n20498, A2 => n17730, ZN => n29717);
   U1696 : NOR2_X2 port map( A1 => n9781, A2 => n18077, ZN => n35748);
   U3414 : INV_X2 port map( I => n34120, ZN => n17477);
   U319 : AOI22_X2 port map( A1 => n18910, A2 => n6932, B1 => n28651, B2 => 
                           n11120, ZN => n28389);
   U5475 : NAND2_X2 port map( A1 => n22038, A2 => n21802, ZN => n22076);
   U4805 : NAND2_X2 port map( A1 => n13114, A2 => n1284, ZN => n13113);
   U4580 : NAND2_X2 port map( A1 => n39401, A2 => n23426, ZN => n31787);
   U1473 : NOR2_X2 port map( A1 => n1346, A2 => n11703, ZN => n35);
   U5994 : INV_X2 port map( I => n4862, ZN => n21143);
   U7569 : INV_X2 port map( I => n29761, ZN => n30747);
   U5472 : INV_X2 port map( I => n28339, ZN => n34007);
   U7356 : NAND2_X2 port map( A1 => n1227, A2 => n3313, ZN => n11140);
   U428 : INV_X2 port map( I => n19631, ZN => n32338);
   U430 : NAND2_X2 port map( A1 => n13601, A2 => n28728, ZN => n15752);
   U5724 : INV_X4 port map( I => n13555, ZN => n7086);
   U7444 : BUF_X4 port map( I => n28033, Z => n37);
   U2953 : NAND2_X2 port map( A1 => n5430, A2 => n28272, ZN => n31027);
   U19589 : NOR2_X2 port map( A1 => n32926, A2 => n33593, ZN => n27245);
   U2441 : INV_X2 port map( I => n13352, ZN => n23124);
   U5809 : INV_X2 port map( I => n11703, ZN => n9288);
   U3944 : AOI21_X2 port map( A1 => n25690, A2 => n14481, B => n19963, ZN => 
                           n25687);
   U4159 : NAND2_X2 port map( A1 => n38610, A2 => n29040, ZN => n15733);
   U4253 : AOI21_X2 port map( A1 => n2927, A2 => n39266, B => n12699, ZN => 
                           n12698);
   U626 : NOR2_X2 port map( A1 => n1070, A2 => n1448, ZN => n4375);
   U3680 : BUF_X2 port map( I => n29456, Z => n19065);
   U19672 : NAND3_X1 port map( A1 => n1893, A2 => n1894, A3 => n17521, ZN => 
                           n445);
   U1312 : NAND2_X2 port map( A1 => n30443, A2 => n11658, ZN => n23100);
   U10327 : OAI21_X2 port map( A1 => n21810, A2 => n13472, B => n2166, ZN => 
                           n21566);
   U2404 : AOI21_X2 port map( A1 => n22303, A2 => n22076, B => n33886, ZN => 
                           n14363);
   U4953 : INV_X2 port map( I => n14601, ZN => n34004);
   U1139 : INV_X2 port map( I => n15679, ZN => n20317);
   U30862 : NAND2_X2 port map( A1 => n26863, A2 => n1230, ZN => n37055);
   U6872 : INV_X2 port map( I => n5897, ZN => n6273);
   U14903 : INV_X2 port map( I => n20416, ZN => n25716);
   U791 : NOR2_X2 port map( A1 => n27213, A2 => n16043, ZN => n27214);
   U1909 : NAND2_X2 port map( A1 => n24784, A2 => n32898, ZN => n24875);
   U5315 : NAND2_X2 port map( A1 => n37227, A2 => n17709, ZN => n19028);
   U16552 : NAND2_X2 port map( A1 => n3694, A2 => n15996, ZN => n15822);
   U14240 : NOR2_X1 port map( A1 => n34821, A2 => n15735, ZN => n18715);
   U2027 : AND2_X2 port map( A1 => n8151, A2 => n11643, Z => n22870);
   U4819 : OR2_X2 port map( A1 => n35252, A2 => n20087, Z => n29581);
   U2614 : NOR2_X2 port map( A1 => n21412, A2 => n21475, ZN => n21564);
   U7815 : INV_X2 port map( I => n35287, ZN => n27410);
   U13447 : AND2_X2 port map( A1 => n32855, A2 => n21767, Z => n21766);
   U15198 : AOI22_X2 port map( A1 => n27990, A2 => n28103, B1 => n27991, B2 => 
                           n2740, ZN => n27993);
   U4152 : NAND2_X2 port map( A1 => n28394, A2 => n28395, ZN => n33574);
   U8429 : NOR2_X2 port map( A1 => n14088, A2 => n30659, ZN => n9140);
   U1334 : INV_X4 port map( I => n21132, ZN => n3803);
   U24379 : INV_X2 port map( I => n22796, ZN => n18750);
   U22261 : INV_X2 port map( I => n10111, ZN => n14394);
   U1269 : AOI21_X2 port map( A1 => n26081, A2 => n13869, B => n10724, ZN => 
                           n30659);
   U20968 : NAND2_X2 port map( A1 => n7494, A2 => n7612, ZN => n27037);
   U9845 : NAND2_X2 port map( A1 => n23331, A2 => n23636, ZN => n3264);
   U6085 : INV_X4 port map( I => n17240, ZN => n971);
   U4590 : INV_X2 port map( I => n24802, ZN => n34354);
   U9574 : INV_X2 port map( I => n14045, ZN => n1252);
   U21057 : INV_X1 port map( I => n8517, ZN => n21839);
   U2348 : NAND2_X2 port map( A1 => n12696, A2 => n10299, ZN => n35441);
   U18313 : OAI22_X2 port map( A1 => n3930, A2 => n11364, B1 => n31383, B2 => 
                           n22328, ZN => n8503);
   U10176 : NOR2_X2 port map( A1 => n13163, A2 => n22326, ZN => n8504);
   U30215 : INV_X4 port map( I => n18619, ZN => n24395);
   U1826 : NOR2_X2 port map( A1 => n4225, A2 => n1566, ZN => n18063);
   U19371 : AOI21_X2 port map( A1 => n7535, A2 => n6969, B => n5487, ZN => 
                           n23244);
   U16955 : INV_X2 port map( I => n28159, ZN => n19541);
   U3078 : INV_X4 port map( I => n15153, ZN => n5669);
   U8410 : NOR2_X2 port map( A1 => n31234, A2 => n34307, ZN => n19119);
   U555 : NAND2_X2 port map( A1 => n37056, A2 => n28153, ZN => n28420);
   U3431 : NAND2_X2 port map( A1 => n2639, A2 => n8476, ZN => n28369);
   U4825 : NOR2_X1 port map( A1 => n4126, A2 => n30878, ZN => n30877);
   U178 : INV_X2 port map( I => n5977, ZN => n29632);
   U595 : INV_X2 port map( I => n17934, ZN => n26660);
   U18103 : NAND2_X2 port map( A1 => n20039, A2 => n35813, ZN => n24872);
   U325 : INV_X2 port map( I => n32682, ZN => n34861);
   U8003 : INV_X4 port map( I => n9242, ZN => n28278);
   U2329 : NAND3_X2 port map( A1 => n35208, A2 => n13823, A3 => n37248, ZN => 
                           n13818);
   U6054 : CLKBUF_X2 port map( I => Key(64), Z => n19583);
   U27621 : NAND2_X1 port map( A1 => n9444, A2 => n28504, ZN => n28507);
   U17464 : NAND2_X2 port map( A1 => n6602, A2 => n39576, ZN => n454);
   U30129 : OAI21_X2 port map( A1 => n15568, A2 => n15569, B => n28229, ZN => 
                           n33620);
   U5501 : AOI21_X2 port map( A1 => n35694, A2 => n16576, B => n1203, ZN => 
                           n10466);
   U24952 : INV_X2 port map( I => n4120, ZN => n32902);
   U6367 : BUF_X2 port map( I => n22796, Z => n23128);
   U16980 : INV_X1 port map( I => n38228, ZN => n27576);
   U17212 : OAI21_X2 port map( A1 => n6160, A2 => n31275, B => n31785, ZN => 
                           n31554);
   U1389 : INV_X2 port map( I => n36666, ZN => n34745);
   U17370 : INV_X2 port map( I => n35151, ZN => n26112);
   U9383 : NAND2_X1 port map( A1 => n17213, A2 => n25939, ZN => n13525);
   U37 : NOR2_X2 port map( A1 => n18384, A2 => n29534, ZN => n29519);
   U3236 : AOI22_X2 port map( A1 => n26775, A2 => n26866, B1 => n20004, B2 => 
                           n26774, ZN => n30617);
   U4350 : BUF_X4 port map( I => n14401, Z => n1109);
   U14216 : INV_X2 port map( I => n19559, ZN => n23602);
   U3710 : OAI21_X2 port map( A1 => n20396, A2 => n21310, B => n1126, ZN => 
                           n24135);
   U5504 : OR2_X2 port map( A1 => n16382, A2 => n13062, Z => n14271);
   U17520 : NAND2_X2 port map( A1 => n29341, A2 => n29336, ZN => n29333);
   U4290 : INV_X4 port map( I => n34717, ZN => n1217);
   U30362 : INV_X2 port map( I => n19515, ZN => n33782);
   U171 : INV_X2 port map( I => n15270, ZN => n15271);
   U1565 : NAND2_X2 port map( A1 => n13516, A2 => n19886, ZN => n12161);
   U1025 : NOR2_X2 port map( A1 => n26920, A2 => n26922, ZN => n35629);
   U9803 : INV_X2 port map( I => n9458, ZN => n1275);
   U25808 : NAND2_X2 port map( A1 => n9514, A2 => n759, ZN => n15334);
   U2943 : NAND2_X2 port map( A1 => n19728, A2 => n8527, ZN => n2158);
   U25872 : INV_X2 port map( I => n39528, ZN => n15448);
   U2578 : INV_X4 port map( I => n22294, ZN => n22246);
   U5807 : NAND2_X2 port map( A1 => n14083, A2 => n25642, ZN => n34465);
   U25074 : NOR2_X2 port map( A1 => n16140, A2 => n35290, ZN => n15890);
   U3851 : INV_X4 port map( I => n22899, ZN => n22849);
   U25188 : NAND2_X1 port map( A1 => n14657, A2 => n24775, ZN => n17971);
   U598 : INV_X4 port map( I => n15594, ZN => n26354);
   U16592 : OAI21_X2 port map( A1 => n36095, A2 => n22915, B => n19293, ZN => 
                           n4102);
   U2296 : NOR2_X2 port map( A1 => n35377, A2 => n31944, ZN => n2633);
   U17752 : BUF_X4 port map( I => n20156, Z => n7251);
   U11629 : NAND2_X2 port map( A1 => n26790, A2 => n4781, ZN => n12352);
   U9121 : OAI21_X2 port map( A1 => n13366, A2 => n14480, B => n17447, ZN => 
                           n11408);
   U17830 : NAND2_X2 port map( A1 => n8735, A2 => n16366, ZN => n35782);
   U1516 : NAND2_X1 port map( A1 => n7696, A2 => n21868, ZN => n12332);
   U221 : NOR2_X2 port map( A1 => n35173, A2 => n28356, ZN => n28535);
   U2463 : INV_X2 port map( I => n35859, ZN => n11307);
   U26558 : AOI21_X2 port map( A1 => n13339, A2 => n15272, B => n20782, ZN => 
                           n33135);
   U2429 : INV_X2 port map( I => n23085, ZN => n20230);
   U2414 : INV_X2 port map( I => n29792, ZN => n29782);
   U6027 : INV_X2 port map( I => n22197, ZN => n1687);
   U17715 : AOI21_X2 port map( A1 => n28649, A2 => n29494, B => n29420, ZN => 
                           n18725);
   U25963 : OAI21_X2 port map( A1 => n5653, A2 => n5210, B => n24909, ZN => 
                           n5209);
   U1381 : INV_X2 port map( I => n11308, ZN => n11315);
   U26557 : NOR2_X2 port map( A1 => n14079, A2 => n17034, ZN => n26662);
   U7539 : OAI21_X2 port map( A1 => n8658, A2 => n8657, B => n1066, ZN => n8656
                           );
   U3591 : OAI22_X2 port map( A1 => n24136, A2 => n24086, B1 => n24309, B2 => 
                           n7730, ZN => n11630);
   U13880 : NAND2_X2 port map( A1 => n9539, A2 => n21854, ZN => n6270);
   U10197 : OAI21_X2 port map( A1 => n9546, A2 => n38246, B => n7916, ZN => 
                           n19011);
   U10892 : BUF_X2 port map( I => n16009, Z => n4849);
   U5955 : INV_X2 port map( I => n524, ZN => n35088);
   U28586 : AOI21_X2 port map( A1 => n23010, A2 => n23009, B => n23308, ZN => 
                           n23016);
   U165 : NAND2_X2 port map( A1 => n35571, A2 => n19962, ZN => n7373);
   U1910 : NAND2_X2 port map( A1 => n17087, A2 => n24623, ZN => n35693);
   U4585 : NAND2_X2 port map( A1 => n10143, A2 => n39401, ZN => n31164);
   U13563 : INV_X4 port map( I => n17692, ZN => n14130);
   U627 : OAI21_X2 port map( A1 => n944, A2 => n1475, B => n19662, ZN => n31498
                           );
   U2212 : OAI21_X2 port map( A1 => n13489, A2 => n12236, B => n37289, ZN => 
                           n13488);
   U4763 : AOI21_X2 port map( A1 => n38283, A2 => n19645, B => n19469, ZN => 
                           n15627);
   U1070 : INV_X4 port map( I => n1607, ZN => n24330);
   U10308 : OAI22_X2 port map( A1 => n21635, A2 => n32138, B1 => n12754, B2 => 
                           n21944, ZN => n11303);
   U1445 : INV_X2 port map( I => n21802, ZN => n22073);
   U17386 : NAND3_X2 port map( A1 => n13294, A2 => n8262, A3 => n5101, ZN => 
                           n27242);
   U6392 : NOR2_X2 port map( A1 => n20034, A2 => n39284, ZN => n9485);
   U15413 : NAND2_X2 port map( A1 => n24076, A2 => n23911, ZN => n7114);
   U10141 : INV_X2 port map( I => n33510, ZN => n36517);
   U18633 : BUF_X4 port map( I => n11562, Z => n948);
   U761 : INV_X2 port map( I => n16736, ZN => n944);
   U16132 : OAI21_X2 port map( A1 => n36461, A2 => n30775, B => n6583, ZN => 
                           n24056);
   U2488 : AOI21_X2 port map( A1 => n22359, A2 => n22358, B => n31939, ZN => 
                           n14801);
   U13069 : INV_X2 port map( I => n19188, ZN => n8884);
   U16788 : AOI21_X2 port map( A1 => n7404, A2 => n36922, B => n34402, ZN => 
                           n14722);
   U13846 : OAI21_X2 port map( A1 => n19553, A2 => n39672, B => n19552, ZN => 
                           n21686);
   U6399 : INV_X2 port map( I => n22041, ZN => n17530);
   U18840 : AND2_X1 port map( A1 => n16039, A2 => n15370, Z => n11900);
   U2586 : NOR2_X2 port map( A1 => n31480, A2 => n6102, ZN => n6099);
   U26196 : INV_X2 port map( I => n14481, ZN => n19813);
   U27605 : INV_X2 port map( I => n10231, ZN => n26645);
   U7712 : INV_X4 port map( I => n33957, ZN => n12784);
   U6160 : INV_X2 port map( I => n35191, ZN => n1634);
   U5901 : NAND2_X2 port map( A1 => n28698, A2 => n28696, ZN => n28366);
   U16229 : BUF_X4 port map( I => n33736, Z => n31504);
   U12420 : NOR2_X2 port map( A1 => n23389, A2 => n38408, ZN => n20450);
   U24220 : BUF_X2 port map( I => n15463, Z => n32815);
   U2294 : CLKBUF_X4 port map( I => n39401, Z => n36885);
   U9933 : INV_X2 port map( I => n18866, ZN => n23404);
   U282 : NAND3_X2 port map( A1 => n28213, A2 => n28212, A3 => n16869, ZN => 
                           n28352);
   U6782 : INV_X2 port map( I => n10370, ZN => n5699);
   U14110 : INV_X2 port map( I => n13966, ZN => n31198);
   U31 : INV_X2 port map( I => n11067, ZN => n13804);
   U675 : NAND2_X2 port map( A1 => n17994, A2 => n25954, ZN => n9589);
   U7443 : NOR2_X2 port map( A1 => n1446, A2 => n8368, ZN => n14585);
   U11624 : OAI21_X2 port map( A1 => n27391, A2 => n27035, B => n27200, ZN => 
                           n27036);
   U1420 : NAND3_X2 port map( A1 => n25697, A2 => n25698, A3 => n32654, ZN => 
                           n32615);
   U6608 : NAND2_X2 port map( A1 => n5616, A2 => n5618, ZN => n34259);
   U18277 : NAND2_X2 port map( A1 => n2340, A2 => n15136, ZN => n31723);
   U14576 : INV_X4 port map( I => n2153, ZN => n22262);
   U26313 : INV_X2 port map( I => n22247, ZN => n16140);
   U8237 : BUF_X4 port map( I => n3441, Z => n2747);
   U1469 : AOI21_X2 port map( A1 => n10044, A2 => n21693, B => n8971, ZN => 
                           n21494);
   U6672 : NAND2_X2 port map( A1 => n22129, A2 => n8245, ZN => n16463);
   U1137 : OAI21_X2 port map( A1 => n25764, A2 => n10724, B => n25989, ZN => 
                           n4801);
   U7164 : INV_X2 port map( I => n15290, ZN => n6647);
   U19558 : INV_X2 port map( I => n13880, ZN => n975);
   U17979 : NAND2_X2 port map( A1 => n16115, A2 => n33845, ZN => n18673);
   U1647 : NOR2_X2 port map( A1 => n34689, A2 => n32131, ZN => n18438);
   U17873 : AOI22_X2 port map( A1 => n31326, A2 => n29990, B1 => n30045, B2 => 
                           n4011, ZN => n35234);
   U3278 : NAND3_X2 port map( A1 => n98, A2 => n9346, A3 => n23413, ZN => 
                           n36927);
   U21040 : INV_X2 port map( I => n36075, ZN => n10199);
   U151 : NAND2_X2 port map( A1 => n37100, A2 => n14422, ZN => n29449);
   U3626 : AOI22_X2 port map( A1 => n14249, A2 => n33086, B1 => n14250, B2 => 
                           n14139, ZN => n14248);
   U18355 : INV_X2 port map( I => n36623, ZN => n17714);
   U3241 : OAI21_X2 port map( A1 => n32802, A2 => n39537, B => n17343, ZN => 
                           n20959);
   U13554 : NAND2_X2 port map( A1 => n23166, A2 => n22973, ZN => n23088);
   U5042 : INV_X4 port map( I => n5541, ZN => n12533);
   U19815 : INV_X4 port map( I => n20931, ZN => n29990);
   U2248 : NOR2_X2 port map( A1 => n23480, A2 => n9078, ZN => n35013);
   U18419 : NAND2_X2 port map( A1 => n3633, A2 => n11923, ZN => n36594);
   U28460 : NAND2_X2 port map( A1 => n20638, A2 => n20408, ZN => n5464);
   U7517 : AOI21_X2 port map( A1 => n28608, A2 => n11390, B => n34737, ZN => 
                           n6095);
   U7151 : OAI21_X2 port map( A1 => n19944, A2 => n23171, B => n23172, ZN => 
                           n18331);
   U2609 : INV_X2 port map( I => n17923, ZN => n16288);
   U16342 : INV_X2 port map( I => n26112, ZN => n33753);
   U2676 : OAI21_X2 port map( A1 => n17433, A2 => n33226, B => n38878, ZN => 
                           n17435);
   U2789 : NOR2_X2 port map( A1 => n10931, A2 => n37355, ZN => n32641);
   U3467 : INV_X2 port map( I => n14704, ZN => n11265);
   U833 : INV_X4 port map( I => n12327, ZN => n11910);
   U1023 : INV_X4 port map( I => n19886, ZN => n1027);
   U15338 : NOR3_X2 port map( A1 => n365, A2 => n33871, A3 => n13971, ZN => 
                           n25759);
   U3448 : BUF_X2 port map( I => n7696, Z => n19549);
   U832 : INV_X2 port map( I => n7676, ZN => n35184);
   U25604 : NAND3_X1 port map( A1 => n36217, A2 => n4976, A3 => n36216, ZN => 
                           n11252);
   U1655 : INV_X4 port map( I => n4914, ZN => n35449);
   U1162 : OAI21_X2 port map( A1 => n33464, A2 => n33465, B => n25345, ZN => 
                           n26067);
   U5159 : INV_X2 port map( I => n5044, ZN => n23572);
   U18267 : NAND2_X2 port map( A1 => n4013, A2 => n18988, ZN => n31114);
   U894 : INV_X2 port map( I => n5271, ZN => n25154);
   U18275 : NAND2_X2 port map( A1 => n18348, A2 => n37259, ZN => n18347);
   U5713 : NAND2_X2 port map( A1 => n37732, A2 => n20339, ZN => n16881);
   U3037 : NAND2_X2 port map( A1 => n9310, A2 => n32870, ZN => n27270);
   U18602 : INV_X2 port map( I => n26063, ZN => n25742);
   U1135 : OAI21_X2 port map( A1 => n14793, A2 => n1106, B => n3356, ZN => 
                           n36574);
   U3732 : INV_X2 port map( I => n25943, ZN => n6302);
   U17046 : OAI21_X2 port map( A1 => n10055, A2 => n12629, B => n34010, ZN => 
                           n12601);
   U3020 : NAND2_X2 port map( A1 => n30210, A2 => n30213, ZN => n30212);
   U351 : INV_X2 port map( I => n37079, ZN => n17032);
   U4773 : AND2_X1 port map( A1 => n11044, A2 => n22222, Z => n14474);
   U1512 : NAND2_X2 port map( A1 => n18028, A2 => n20476, ZN => n18954);
   U8844 : INV_X4 port map( I => n33514, ZN => n13971);
   U17449 : NAND2_X2 port map( A1 => n9265, A2 => n35290, ZN => n164);
   U5070 : BUF_X2 port map( I => n23083, Z => n19865);
   U1855 : OAI21_X2 port map( A1 => n10840, A2 => n1301, B => n32401, ZN => 
                           n10842);
   U467 : NAND2_X2 port map( A1 => n1074, A2 => n28180, ZN => n27946);
   U235 : OAI21_X2 port map( A1 => n35369, A2 => n35370, B => n31269, ZN => 
                           n34395);
   U379 : INV_X2 port map( I => n10883, ZN => n33424);
   U2931 : NOR2_X2 port map( A1 => n19728, A2 => n8527, ZN => n8587);
   U5903 : NAND2_X2 port map( A1 => n24558, A2 => n24757, ZN => n31257);
   U12427 : INV_X4 port map( I => n25468, ZN => n25409);
   U10149 : NAND3_X2 port map( A1 => n12091, A2 => n937, A3 => n22252, ZN => 
                           n22000);
   U1713 : INV_X2 port map( I => n24938, ZN => n25031);
   U9464 : NAND2_X2 port map( A1 => n14025, A2 => n1115, ZN => n11954);
   U2764 : INV_X4 port map( I => n33933, ZN => n20872);
   U5800 : AOI22_X2 port map( A1 => n35157, A2 => n35156, B1 => n25592, B2 => 
                           n32105, ZN => n19401);
   U15187 : OAI21_X2 port map( A1 => n33094, A2 => n37936, B => n33093, ZN => 
                           n28960);
   U245 : INV_X2 port map( I => n28673, ZN => n1068);
   U5648 : NOR2_X2 port map( A1 => n26972, A2 => n5935, ZN => n16000);
   U2928 : NOR2_X2 port map( A1 => n30197, A2 => n30198, ZN => n30199);
   U858 : NOR2_X2 port map( A1 => n20052, A2 => n31809, ZN => n8980);
   U6404 : NOR2_X2 port map( A1 => n21879, A2 => n21878, ZN => n22041);
   U4271 : NOR2_X2 port map( A1 => n23550, A2 => n38614, ZN => n23347);
   U143 : AND2_X2 port map( A1 => n10422, A2 => n36426, Z => n17444);
   U22681 : NAND2_X2 port map( A1 => n4699, A2 => n3669, ZN => n10321);
   U12074 : OAI22_X2 port map( A1 => n25903, A2 => n33474, B1 => n26016, B2 => 
                           n38825, ZN => n12458);
   U7041 : INV_X4 port map( I => n20517, ZN => n1032);
   U2355 : NOR2_X2 port map( A1 => n6005, A2 => n36230, ZN => n32943);
   U2214 : NAND2_X2 port map( A1 => n17816, A2 => n39371, ZN => n32207);
   U30050 : NAND2_X1 port map( A1 => n8580, A2 => n8579, ZN => n7971);
   U217 : INV_X2 port map( I => n28791, ZN => n248);
   U7056 : NAND2_X2 port map( A1 => n25820, A2 => n36798, ZN => n25931);
   U14845 : INV_X2 port map( I => n37954, ZN => n24228);
   U2500 : NAND2_X2 port map( A1 => n5876, A2 => n22236, ZN => n35802);
   U3497 : NOR2_X2 port map( A1 => n13038, A2 => n23349, ZN => n16443);
   U276 : NOR2_X2 port map( A1 => n14232, A2 => n28012, ZN => n11876);
   U3373 : INV_X2 port map( I => n18545, ZN => n1546);
   U5707 : INV_X1 port map( I => n37355, ZN => n1578);
   U6876 : INV_X4 port map( I => n26086, ZN => n25874);
   U7479 : INV_X2 port map( I => n1448, ZN => n986);
   U1970 : INV_X2 port map( I => n9583, ZN => n9579);
   U11548 : INV_X4 port map( I => n9893, ZN => n955);
   U8376 : NAND2_X2 port map( A1 => n23537, A2 => n23539, ZN => n23225);
   U7258 : INV_X2 port map( I => n8413, ZN => n8103);
   U3909 : INV_X2 port map( I => n38194, ZN => n14064);
   U12366 : INV_X2 port map( I => n13988, ZN => n9541);
   U18050 : AOI22_X2 port map( A1 => n36092, A2 => n34128, B1 => n22060, B2 => 
                           n8618, ZN => n22784);
   U3868 : NOR2_X2 port map( A1 => n7387, A2 => n38724, ZN => n36137);
   U9750 : OAI21_X2 port map( A1 => n18141, A2 => n13710, B => n1601, ZN => 
                           n13709);
   U13820 : AND2_X2 port map( A1 => n15697, A2 => n4342, Z => n8618);
   U7045 : INV_X2 port map( I => n24095, ZN => n24477);
   U2142 : INV_X2 port map( I => n23697, ZN => n23779);
   U26305 : INV_X2 port map( I => n17605, ZN => n22762);
   U666 : NOR2_X2 port map( A1 => n16904, A2 => n16903, ZN => n21265);
   U27173 : OAI21_X2 port map( A1 => n28226, A2 => n35659, B => n19921, ZN => 
                           n20226);
   U2178 : AOI21_X2 port map( A1 => n13691, A2 => n23645, B => n35312, ZN => 
                           n35285);
   U20709 : INV_X4 port map( I => n39678, ZN => n8014);
   U9861 : NAND2_X2 port map( A1 => n23462, A2 => n18090, ZN => n18155);
   U21571 : NOR2_X1 port map( A1 => n1275, A2 => n1131, ZN => n9459);
   U7796 : OAI21_X2 port map( A1 => n3515, A2 => n3514, B => n27072, ZN => 
                           n4492);
   U6867 : NAND2_X2 port map( A1 => n7198, A2 => n24795, ZN => n9614);
   U465 : AOI22_X2 port map( A1 => n8880, A2 => n28194, B1 => n9897, B2 => 
                           n37251, ZN => n3846);
   U6314 : NOR2_X2 port map( A1 => n14392, A2 => n24300, ZN => n13112);
   U21139 : AOI21_X2 port map( A1 => n23452, A2 => n10480, B => n8668, ZN => 
                           n16713);
   U14727 : NOR2_X2 port map( A1 => n34399, A2 => n11003, ZN => n31299);
   U4925 : NAND2_X2 port map( A1 => n8971, A2 => n21804, ZN => n4298);
   U12575 : NAND2_X2 port map( A1 => n24736, A2 => n37687, ZN => n2850);
   U2684 : NAND3_X2 port map( A1 => n19123, A2 => n19124, A3 => n19125, ZN => 
                           n36072);
   U16810 : NAND2_X2 port map( A1 => n32974, A2 => n25874, ZN => n26088);
   U2570 : INV_X2 port map( I => n31573, ZN => n36960);
   U5030 : INV_X2 port map( I => n35244, ZN => n1288);
   U6950 : NAND2_X2 port map( A1 => n14999, A2 => n13966, ZN => n24757);
   U3557 : AOI21_X2 port map( A1 => n25840, A2 => n11807, B => n8233, ZN => 
                           n8234);
   U450 : AOI22_X2 port map( A1 => n37136, A2 => n28283, B1 => n13993, B2 => 
                           n16544, ZN => n28170);
   U14100 : NAND2_X1 port map( A1 => n34805, A2 => n29587, ZN => n34804);
   U27288 : INV_X2 port map( I => n22349, ZN => n1332);
   U30631 : BUF_X4 port map( I => n21912, Z => n36912);
   U3571 : OAI22_X2 port map( A1 => n14495, A2 => n15651, B1 => n16171, B2 => 
                           n30238, ZN => n5632);
   U2491 : BUF_X2 port map( I => n32932, Z => n31607);
   U16049 : OAI21_X1 port map( A1 => n980, A2 => n28690, B => n2639, ZN => 
                           n31461);
   U6695 : INV_X2 port map( I => n9845, ZN => n14451);
   U13752 : NOR2_X2 port map( A1 => n14251, A2 => n22259, ZN => n17001);
   U8351 : INV_X4 port map( I => n15461, ZN => n1128);
   U4436 : INV_X4 port map( I => n31679, ZN => n1265);
   U13118 : NAND3_X2 port map( A1 => n17959, A2 => n17958, A3 => n38055, ZN => 
                           n16031);
   U9114 : NOR2_X2 port map( A1 => n18277, A2 => n18276, ZN => n7034);
   U17676 : AND2_X1 port map( A1 => n31917, A2 => n26090, Z => n5682);
   U8835 : INV_X2 port map( I => n3257, ZN => n27624);
   U1392 : INV_X2 port map( I => n260, ZN => n16073);
   U10933 : BUF_X2 port map( I => n29296, Z => n4816);
   U4450 : OR2_X1 port map( A1 => n36827, A2 => n7023, Z => n28606);
   U571 : NOR2_X2 port map( A1 => n12260, A2 => n876, ZN => n13984);
   U4244 : NAND2_X1 port map( A1 => n5034, A2 => n9503, ZN => n31640);
   U1790 : NAND3_X2 port map( A1 => n13896, A2 => n30412, A3 => n27259, ZN => 
                           n5374);
   U7096 : NOR2_X2 port map( A1 => n603, A2 => n25797, ZN => n25855);
   U18732 : NAND3_X2 port map( A1 => n30470, A2 => n25519, A3 => n20924, ZN => 
                           n5902);
   U454 : OAI22_X2 port map( A1 => n33481, A2 => n28152, B1 => n16412, B2 => 
                           n8960, ZN => n28402);
   U1649 : NAND2_X2 port map( A1 => n31509, A2 => n5541, ZN => n25416);
   U16912 : INV_X4 port map( I => n9733, ZN => n32671);
   U22334 : INV_X4 port map( I => n28771, ZN => n35777);
   U190 : INV_X4 port map( I => n28768, ZN => n28771);
   U213 : NAND2_X2 port map( A1 => n11488, A2 => n11490, ZN => n28529);
   U668 : NAND2_X2 port map( A1 => n10946, A2 => n36865, ZN => n1835);
   U994 : INV_X4 port map( I => n17993, ZN => n32745);
   U60 : OAI21_X2 port map( A1 => n16988, A2 => n6863, B => n39392, ZN => 
                           n29273);
   U6141 : INV_X2 port map( I => n27777, ZN => n1460);
   U1085 : NAND2_X2 port map( A1 => n14378, A2 => n17709, ZN => n14123);
   U15923 : NAND2_X2 port map( A1 => n30290, A2 => n27282, ZN => n26264);
   U39 : INV_X2 port map( I => n29568, ZN => n29567);
   U6211 : INV_X2 port map( I => n23214, ZN => n17568);
   U6165 : NAND2_X2 port map( A1 => n36035, A2 => n35536, ZN => n31475);
   U4426 : OR2_X1 port map( A1 => n19658, A2 => n33937, Z => n24225);
   U25352 : NOR2_X2 port map( A1 => n20585, A2 => n21328, ZN => n22306);
   U936 : INV_X2 port map( I => n26743, ZN => n35877);
   U7482 : INV_X2 port map( I => n31279, ZN => n1406);
   U6045 : INV_X2 port map( I => n21577, ZN => n21593);
   U1695 : INV_X2 port map( I => n37050, ZN => n17246);
   U7050 : NAND2_X2 port map( A1 => n39301, A2 => n8212, ZN => n8211);
   U8924 : NAND2_X2 port map( A1 => n25604, A2 => n9029, ZN => n34261);
   U7617 : INV_X2 port map( I => n29517, ZN => n33427);
   U929 : OAI21_X2 port map( A1 => n19886, A2 => n36296, B => n12159, ZN => 
                           n11198);
   U4755 : BUF_X2 port map( I => n12396, Z => n33538);
   U10452 : BUF_X2 port map( I => Key(6), Z => n29649);
   U7502 : INV_X4 port map( I => n28396, ZN => n32791);
   U4845 : INV_X2 port map( I => n1154, ZN => n31649);
   U9957 : NOR2_X2 port map( A1 => n10297, A2 => n10296, ZN => n10295);
   U8476 : OAI21_X2 port map( A1 => n8707, A2 => n1313, B => n23142, ZN => 
                           n10297);
   U25462 : INV_X1 port map( I => n36196, ZN => n6898);
   U30103 : OAI22_X2 port map( A1 => n25991, A2 => n11807, B1 => n18289, B2 => 
                           n9883, ZN => n4854);
   U1949 : INV_X2 port map( I => n23619, ZN => n20835);
   U2353 : NAND2_X2 port map( A1 => n34185, A2 => n34184, ZN => n22907);
   U12977 : NOR2_X2 port map( A1 => n32683, A2 => n37107, ZN => n4244);
   U3798 : NAND2_X2 port map( A1 => n22055, A2 => n22132, ZN => n22056);
   U4186 : AND2_X1 port map( A1 => n25782, A2 => n8407, Z => n13119);
   U826 : AOI21_X2 port map( A1 => n25562, A2 => n25637, B => n25436, ZN => 
                           n25439);
   U9703 : NOR2_X2 port map( A1 => n9634, A2 => n13809, ZN => n21211);
   U17990 : BUF_X2 port map( I => n27211, Z => n36203);
   U30119 : INV_X2 port map( I => n28109, ZN => n33612);
   U4628 : NAND2_X2 port map( A1 => n3013, A2 => n38168, ZN => n9962);
   U9353 : INV_X4 port map( I => n19332, ZN => n1235);
   U11454 : INV_X4 port map( I => n27478, ZN => n27815);
   U13732 : NAND2_X2 port map( A1 => n22107, A2 => n7613, ZN => n17898);
   U13611 : INV_X2 port map( I => n22573, ZN => n13768);
   U14090 : BUF_X4 port map( I => n3713, Z => n32260);
   U11321 : NAND2_X2 port map( A1 => n15389, A2 => n42, ZN => n27936);
   U5951 : INV_X2 port map( I => n24794, ZN => n1563);
   U166 : NOR2_X2 port map( A1 => n1175, A2 => n35210, ZN => n34619);
   U6772 : INV_X2 port map( I => n5323, ZN => n23831);
   U14696 : OAI21_X2 port map( A1 => n20395, A2 => n12286, B => n24156, ZN => 
                           n34895);
   U13555 : INV_X2 port map( I => n23189, ZN => n1647);
   U23637 : NAND2_X2 port map( A1 => n935, A2 => n35684, ZN => n8869);
   U808 : OAI21_X2 port map( A1 => n36262, A2 => n33026, B => n33025, ZN => 
                           n26153);
   U438 : INV_X2 port map( I => n27506, ZN => n601);
   U17190 : OAI21_X2 port map( A1 => n35897, A2 => n21248, B => n30544, ZN => 
                           n27506);
   U4167 : INV_X2 port map( I => n24308, ZN => n24446);
   U7300 : INV_X2 port map( I => n1217, ZN => n34943);
   U23074 : NOR2_X2 port map( A1 => n1094, A2 => n1786, ZN => n26957);
   U3411 : OAI21_X2 port map( A1 => n13053, A2 => n27955, B => n17477, ZN => 
                           n385);
   U1698 : NOR2_X2 port map( A1 => n25725, A2 => n38661, ZN => n36686);
   U5411 : OAI21_X2 port map( A1 => n14712, A2 => n14713, B => n28627, ZN => 
                           n36255);
   U8929 : NOR2_X2 port map( A1 => n13714, A2 => n20896, ZN => n27955);
   U9604 : AOI22_X2 port map( A1 => n34666, A2 => n1121, B1 => n24782, B2 => 
                           n24658, ZN => n4694);
   U9478 : NAND2_X2 port map( A1 => n4217, A2 => n4216, ZN => n4215);
   U1164 : AOI21_X2 port map( A1 => n10290, A2 => n35109, B => n20769, ZN => 
                           n20768);
   U2385 : NAND2_X2 port map( A1 => n18365, A2 => n17578, ZN => n7012);
   U695 : OAI21_X2 port map( A1 => n37191, A2 => n3998, B => n3996, ZN => 
                           n35037);
   U7833 : INV_X4 port map( I => n35919, ZN => n1081);
   U604 : INV_X4 port map( I => n26695, ZN => n1495);
   U4602 : NAND2_X2 port map( A1 => n24693, A2 => n24721, ZN => n30862);
   U18359 : INV_X4 port map( I => n30161, ZN => n33277);
   U5689 : INV_X4 port map( I => n25434, ZN => n25674);
   U3970 : INV_X2 port map( I => n6686, ZN => n27416);
   U960 : OAI21_X2 port map( A1 => n14921, A2 => n14922, B => n1490, ZN => 
                           n12684);
   U7912 : BUF_X2 port map( I => n20394, Z => n17076);
   U24130 : NAND2_X2 port map( A1 => n25622, A2 => n33785, ZN => n2417);
   U16 : INV_X2 port map( I => n19297, ZN => n29658);
   U1205 : NOR2_X2 port map( A1 => n39061, A2 => n39160, ZN => n4455);
   U4058 : OAI22_X2 port map( A1 => n11009, A2 => n31321, B1 => n28716, B2 => 
                           n33591, ZN => n16503);
   U25465 : AOI21_X1 port map( A1 => n26606, A2 => n13219, B => n26986, ZN => 
                           n36196);
   U24725 : INV_X2 port map( I => n15004, ZN => n16935);
   U5876 : INV_X2 port map( I => n4192, ZN => n991);
   U12916 : OAI21_X2 port map( A1 => n24142, A2 => n18302, B => n14123, ZN => 
                           n14780);
   U1567 : OAI21_X1 port map( A1 => n18218, A2 => n34156, B => n18217, ZN => 
                           n25655);
   U22515 : NAND2_X2 port map( A1 => n32526, A2 => n15324, ZN => n16055);
   U3436 : NAND2_X2 port map( A1 => n1783, A2 => n24700, ZN => n1782);
   U12045 : NOR2_X2 port map( A1 => n25781, A2 => n25774, ZN => n15870);
   U2323 : INV_X4 port map( I => n21068, ZN => n23518);
   U1231 : NAND3_X2 port map( A1 => n25409, A2 => n14635, A3 => n25467, ZN => 
                           n25339);
   U14496 : AOI21_X2 port map( A1 => n24426, A2 => n3142, B => n8041, ZN => 
                           n2089);
   U4515 : NAND2_X2 port map( A1 => n33392, A2 => n19507, ZN => n12517);
   U13240 : NAND2_X2 port map( A1 => n23362, A2 => n23480, ZN => n15681);
   U1905 : AOI22_X2 port map( A1 => n8916, A2 => n20863, B1 => n20864, B2 => 
                           n38302, ZN => n11577);
   U16866 : BUF_X4 port map( I => n24745, Z => n35137);
   U10799 : INV_X2 port map( I => n17978, ZN => n30858);
   U5928 : INV_X2 port map( I => n17458, ZN => n1243);
   U7235 : INV_X2 port map( I => n11327, ZN => n22360);
   U7082 : INV_X2 port map( I => n17269, ZN => n9227);
   U2078 : NAND2_X2 port map( A1 => n253, A2 => n24443, ZN => n24310);
   U18655 : AOI22_X2 port map( A1 => n22072, A2 => n3687, B1 => n22071, B2 => 
                           n33623, ZN => n22380);
   U13831 : AOI22_X2 port map( A1 => n17264, A2 => n18417, B1 => n14542, B2 => 
                           n21712, ZN => n12024);
   U17461 : INV_X4 port map( I => n19410, ZN => n20157);
   U6740 : INV_X2 port map( I => n6176, ZN => n20972);
   U968 : NOR2_X2 port map( A1 => n36262, A2 => n36261, ZN => n7859);
   U1858 : INV_X2 port map( I => n24707, ZN => n24700);
   U12911 : AOI22_X2 port map( A1 => n1274, A2 => n232, B1 => n1123, B2 => 
                           n24116, ZN => n11133);
   U5343 : NOR2_X2 port map( A1 => n1602, A2 => n23819, ZN => n8690);
   U1585 : INV_X2 port map( I => n12836, ZN => n26876);
   U8683 : NAND2_X2 port map( A1 => n21727, A2 => n18293, ZN => n11172);
   U20951 : INV_X4 port map( I => n1029, ZN => n35578);
   U9958 : AOI21_X2 port map( A1 => n11301, A2 => n33361, B => n11299, ZN => 
                           n18034);
   U10200 : NOR2_X2 port map( A1 => n1675, A2 => n18656, ZN => n17156);
   U13890 : OAI21_X1 port map( A1 => n21715, A2 => n21714, B => n21713, ZN => 
                           n21716);
   U813 : NAND2_X2 port map( A1 => n26148, A2 => n36262, ZN => n33025);
   U706 : NAND2_X2 port map( A1 => n5297, A2 => n1217, ZN => n35144);
   U4544 : BUF_X2 port map( I => n10665, Z => n33785);
   U678 : NOR2_X2 port map( A1 => n15245, A2 => n35604, ZN => n35603);
   U22843 : NOR2_X2 port map( A1 => n17691, A2 => n17692, ZN => n11159);
   U30570 : NOR2_X2 port map( A1 => n12814, A2 => n22270, ZN => n5147);
   U17894 : BUF_X4 port map( I => n26893, Z => n33396);
   U8952 : NAND3_X2 port map( A1 => n35392, A2 => n29520, A3 => n29521, ZN => 
                           n29523);
   U2374 : NAND2_X2 port map( A1 => n8707, A2 => n35591, ZN => n8706);
   U16487 : AOI21_X2 port map( A1 => n14229, A2 => n13712, B => n1019, ZN => 
                           n14224);
   U9520 : NAND2_X2 port map( A1 => n25665, A2 => n4001, ZN => n20442);
   U118 : NAND2_X2 port map( A1 => n19896, A2 => n17295, ZN => n17294);
   U1631 : INV_X2 port map( I => n20153, ZN => n25327);
   U19123 : AOI21_X2 port map( A1 => n6375, A2 => n6374, B => n28287, ZN => 
                           n6587);
   U6749 : INV_X2 port map( I => n20418, ZN => n12638);
   U502 : OAI21_X2 port map( A1 => n20941, A2 => n18013, B => n14152, ZN => 
                           n34965);
   U1880 : NOR2_X2 port map( A1 => n2553, A2 => n23456, ZN => n18763);
   U26905 : INV_X4 port map( I => n14501, ZN => n21656);
   U4572 : AOI21_X2 port map( A1 => n35023, A2 => n37081, B => n38529, ZN => 
                           n16255);
   U946 : INV_X4 port map( I => n5935, ZN => n3694);
   U8047 : INV_X2 port map( I => n29794, ZN => n16682);
   U911 : NAND2_X2 port map( A1 => n26840, A2 => n32345, ZN => n18095);
   U11048 : BUF_X4 port map( I => n19771, Z => n7486);
   U19876 : NAND3_X2 port map( A1 => n14437, A2 => n16060, A3 => n36850, ZN => 
                           n31980);
   U2923 : NAND2_X1 port map( A1 => n35787, A2 => n14664, ZN => n16075);
   U9029 : INV_X2 port map( I => n8944, ZN => n1433);
   U6630 : NAND2_X2 port map( A1 => n20372, A2 => n34419, ZN => n22843);
   U6459 : INV_X2 port map( I => n21982, ZN => n1686);
   U1154 : AOI21_X2 port map( A1 => n26107, A2 => n25825, B => n16200, ZN => 
                           n15551);
   U5905 : NOR2_X2 port map( A1 => n18541, A2 => n16908, ZN => n24716);
   U30576 : INV_X2 port map( I => n39067, ZN => n24464);
   U8360 : INV_X2 port map( I => n23590, ZN => n23874);
   U3855 : INV_X4 port map( I => n23053, ZN => n1043);
   U8427 : NAND2_X2 port map( A1 => n31644, A2 => n32260, ZN => n3714);
   U7546 : BUF_X2 port map( I => n29042, Z => n31782);
   U17525 : INV_X2 port map( I => n16539, ZN => n31891);
   U15894 : NOR2_X1 port map( A1 => n936, A2 => n14089, ZN => n2272);
   U947 : OAI21_X2 port map( A1 => n2929, A2 => n20578, B => n38238, ZN => 
                           n17416);
   U4700 : OR2_X1 port map( A1 => n17594, A2 => n37085, Z => n25615);
   U2621 : NAND2_X2 port map( A1 => n5075, A2 => n9252, ZN => n29);
   U2129 : INV_X4 port map( I => n23819, ZN => n1123);
   U28774 : NAND2_X2 port map( A1 => n33648, A2 => n18031, ZN => n36612);
   U6157 : INV_X2 port map( I => n21808, ZN => n1345);
   U6869 : NOR2_X2 port map( A1 => n19484, A2 => n38884, ZN => n24518);
   U24437 : NAND2_X2 port map( A1 => n16729, A2 => n7379, ZN => n16728);
   U6213 : AOI22_X2 port map( A1 => n37073, A2 => n11858, B1 => n25888, B2 => 
                           n928, ZN => n12941);
   U2284 : NAND2_X2 port map( A1 => n36263, A2 => n17887, ZN => n36131);
   U7531 : AOI21_X2 port map( A1 => n33229, A2 => n28478, B => n2191, ZN => 
                           n16036);
   U2859 : AOI21_X2 port map( A1 => n18999, A2 => n5821, B => n31649, ZN => 
                           n31953);
   U17703 : NAND2_X1 port map( A1 => n21220, A2 => n20885, ZN => n4901);
   U1356 : NAND2_X2 port map( A1 => n34898, A2 => n26075, ZN => n26079);
   U1707 : INV_X2 port map( I => n25392, ZN => n25587);
   U8256 : INV_X4 port map( I => n32091, ZN => n19484);
   U4265 : INV_X4 port map( I => n17118, ZN => n22236);
   U5715 : NAND2_X2 port map( A1 => n20545, A2 => n38899, ZN => n36458);
   U2447 : AOI22_X2 port map( A1 => n20590, A2 => n20344, B1 => n22793, B2 => 
                           n20174, ZN => n34664);
   U8480 : NOR2_X2 port map( A1 => n23121, A2 => n19440, ZN => n30663);
   U1407 : INV_X2 port map( I => n31809, ZN => n1537);
   U12649 : INV_X2 port map( I => n24770, ZN => n12460);
   U6643 : INV_X2 port map( I => n20638, ZN => n14524);
   U413 : INV_X4 port map( I => n36320, ZN => n2191);
   U2366 : AOI21_X2 port map( A1 => n36234, A2 => n27149, B => n27235, ZN => 
                           n5997);
   U8553 : INV_X2 port map( I => n17021, ZN => n22921);
   U11612 : NAND2_X2 port map( A1 => n5082, A2 => n37076, ZN => n5297);
   U704 : NAND2_X2 port map( A1 => n31150, A2 => n31298, ZN => n34579);
   U288 : AOI21_X2 port map( A1 => n33436, A2 => n1194, B => n1431, ZN => 
                           n19688);
   U1361 : INV_X4 port map( I => n35059, ZN => n20813);
   U9851 : NAND2_X1 port map( A1 => n9862, A2 => n23555, ZN => n15325);
   U2736 : NAND2_X2 port map( A1 => n27149, A2 => n27436, ZN => n15983);
   U14432 : OAI21_X2 port map( A1 => n11042, A2 => n11041, B => n2035, ZN => 
                           n11040);
   U338 : INV_X2 port map( I => n28570, ZN => n37018);
   U19003 : OAI21_X2 port map( A1 => n18617, A2 => n34121, B => n34245, ZN => 
                           n6463);
   U20220 : NOR2_X2 port map( A1 => n11547, A2 => n1532, ZN => n7513);
   U2058 : INV_X2 port map( I => n30000, ZN => n21167);
   U10718 : OAI22_X2 port map( A1 => n6862, A2 => n11056, B1 => n29421, B2 => 
                           n13153, ZN => n6866);
   U2493 : NOR2_X2 port map( A1 => n36085, A2 => n36084, ZN => n4111);
   U262 : NAND2_X2 port map( A1 => n12543, A2 => n28651, ZN => n36144);
   U3128 : NOR2_X2 port map( A1 => n19865, A2 => n20372, ZN => n10470);
   U845 : AOI21_X2 port map( A1 => n39117, A2 => n14079, B => n1008, ZN => 
                           n12405);
   U23083 : OAI21_X2 port map( A1 => n365, A2 => n34154, B => n2942, ZN => 
                           n2941);
   U12117 : NOR2_X2 port map( A1 => n39824, A2 => n11616, ZN => n31018);
   U399 : INV_X2 port map( I => n32002, ZN => n36775);
   U6627 : INV_X2 port map( I => n13686, ZN => n925);
   U22234 : INV_X2 port map( I => n21721, ZN => n21645);
   U24714 : AOI21_X2 port map( A1 => n21573, A2 => n15839, B => n20580, ZN => 
                           n20579);
   U13703 : NOR2_X2 port map( A1 => n18129, A2 => n1148, ZN => n7868);
   U9921 : OAI21_X2 port map( A1 => n17556, A2 => n23569, B => n23543, ZN => 
                           n23546);
   U17034 : INV_X2 port map( I => n25602, ZN => n35157);
   U4232 : NAND2_X2 port map( A1 => n1029, A2 => n9825, ZN => n24752);
   U19849 : OAI22_X2 port map( A1 => n31975, A2 => n17266, B1 => n21745, B2 => 
                           n19542, ZN => n19906);
   U19188 : NAND2_X2 port map( A1 => n1148, A2 => n584, ZN => n6450);
   U11103 : INV_X4 port map( I => n865, ZN => n6615);
   U6579 : NAND2_X2 port map( A1 => n22133, A2 => n22132, ZN => n4121);
   U154 : NAND2_X2 port map( A1 => n36924, A2 => n12353, ZN => n36923);
   U5748 : INV_X2 port map( I => n14477, ZN => n1136);
   U1063 : INV_X2 port map( I => n36858, ZN => n865);
   U6959 : INV_X4 port map( I => n17658, ZN => n1118);
   U8298 : NAND2_X1 port map( A1 => n30651, A2 => n2889, ZN => n4460);
   U1156 : INV_X4 port map( I => n18142, ZN => n31133);
   U2555 : NAND2_X2 port map( A1 => n33571, A2 => n35290, ZN => n22141);
   U14770 : OAI21_X2 port map( A1 => n4367, A2 => n30175, B => n39122, ZN => 
                           n34903);
   U15651 : NAND2_X2 port map( A1 => n39501, A2 => n17658, ZN => n24161);
   U1479 : OAI21_X2 port map( A1 => n14666, A2 => n9602, B => n1249, ZN => 
                           n35492);
   U30066 : NAND2_X2 port map( A1 => n1432, A2 => n4232, ZN => n28605);
   U20475 : NAND2_X1 port map( A1 => n16868, A2 => n12192, ZN => n18019);
   U28376 : NOR3_X2 port map( A1 => n39284, A2 => n32039, A3 => n196, ZN => 
                           n21965);
   U6028 : OAI21_X2 port map( A1 => n18752, A2 => n30378, B => n16081, ZN => 
                           n36725);
   U10271 : NOR2_X2 port map( A1 => n34025, A2 => n34393, ZN => n34392);
   U11881 : NOR2_X2 port map( A1 => n26982, A2 => n26979, ZN => n4982);
   U2182 : NOR3_X2 port map( A1 => n32858, A2 => n1297, A3 => n6969, ZN => 
                           n18680);
   U1200 : NAND3_X2 port map( A1 => n17003, A2 => n26133, A3 => n25936, ZN => 
                           n21306);
   U11593 : NAND2_X2 port map( A1 => n37201, A2 => n27284, ZN => n9493);
   U13792 : AND3_X1 port map( A1 => n22315, A2 => n15004, A3 => n22277, Z => 
                           n14508);
   U24678 : INV_X2 port map( I => n35832, ZN => n20692);
   U12796 : NOR2_X1 port map( A1 => n19453, A2 => n12040, ZN => n33468);
   U9714 : NOR2_X2 port map( A1 => n5714, A2 => n20653, ZN => n5713);
   U22491 : OAI21_X2 port map( A1 => n23060, A2 => n36724, B => n19535, ZN => 
                           n22705);
   U5216 : BUF_X4 port map( I => n23592, Z => n4147);
   U2161 : INV_X2 port map( I => n23976, ZN => n1616);
   U9243 : AOI21_X2 port map( A1 => n26667, A2 => n17237, B => n1002, ZN => 
                           n14280);
   U442 : AOI21_X2 port map( A1 => n6714, A2 => n879, B => n38365, ZN => n6713)
                           ;
   U17069 : INV_X4 port map( I => n33453, ZN => n6217);
   U19489 : NOR2_X2 port map( A1 => n6770, A2 => n37210, ZN => n14168);
   U6947 : OR2_X2 port map( A1 => n1118, A2 => n24226, Z => n24964);
   U9365 : INV_X2 port map( I => n26463, ZN => n1238);
   U747 : INV_X2 port map( I => n27404, ZN => n1079);
   U24476 : NAND2_X1 port map( A1 => n2726, A2 => n17319, ZN => n2725);
   U1552 : OAI21_X2 port map( A1 => n13949, A2 => n13948, B => n26986, ZN => 
                           n13947);
   U6723 : INV_X4 port map( I => n34962, ZN => n1642);
   U6488 : OAI21_X2 port map( A1 => n22265, A2 => n19515, B => n22267, ZN => 
                           n33781);
   U1906 : BUF_X4 port map( I => n22234, Z => n19261);
   U6331 : NOR2_X1 port map( A1 => n23529, A2 => n18236, ZN => n8928);
   U13093 : NOR2_X1 port map( A1 => n36248, A2 => n36247, ZN => n36246);
   U2530 : OAI21_X2 port map( A1 => n1327, A2 => n11329, B => n22287, ZN => 
                           n34822);
   U1539 : INV_X1 port map( I => n21722, ZN => n21640);
   U15423 : OAI21_X2 port map( A1 => n10473, A2 => n32782, B => n25748, ZN => 
                           n26478);
   U7851 : OAI21_X2 port map( A1 => n3417, A2 => n1500, B => n33689, ZN => 
                           n2238);
   U1781 : BUF_X4 port map( I => n7923, Z => n2576);
   U3927 : INV_X1 port map( I => n25490, ZN => n25517);
   U13238 : AOI22_X2 port map( A1 => n23556, A2 => n31234, B1 => n16443, B2 => 
                           n32616, ZN => n23558);
   U8589 : AOI21_X2 port map( A1 => n916, A2 => n22349, B => n2910, ZN => n7814
                           );
   U11772 : OAI21_X2 port map( A1 => n10678, A2 => n10187, B => n26354, ZN => 
                           n10186);
   U12438 : OAI21_X2 port map( A1 => n9526, A2 => n18837, B => n38685, ZN => 
                           n12599);
   U7247 : BUF_X4 port map( I => n22113, Z => n1049);
   U13230 : NOR2_X1 port map( A1 => n596, A2 => n3926, ZN => n32721);
   U2420 : NAND2_X2 port map( A1 => n10345, A2 => n21402, ZN => n14846);
   U8518 : INV_X4 port map( I => n33745, ZN => n11328);
   U17009 : AOI21_X2 port map( A1 => n683, A2 => n123, B => n35153, ZN => 
                           n10128);
   U17565 : NAND2_X1 port map( A1 => n9278, A2 => n17456, ZN => n5015);
   U4658 : OR3_X1 port map( A1 => n15414, A2 => n20128, A3 => n14064, Z => 
                           n13664);
   U7848 : NAND2_X2 port map( A1 => n13156, A2 => n14757, ZN => n27390);
   U532 : OAI21_X2 port map( A1 => n1494, A2 => n20211, B => n13757, ZN => 
                           n20636);
   U14844 : INV_X4 port map( I => n2395, ZN => n12733);
   U5615 : OAI21_X2 port map( A1 => n4776, A2 => n25897, B => n37582, ZN => 
                           n6397);
   U4467 : INV_X4 port map( I => n1302, ZN => n17167);
   U27294 : INV_X4 port map( I => n18585, ZN => n19262);
   U5845 : CLKBUF_X4 port map( I => n25157, Z => n25754);
   U7360 : NOR2_X2 port map( A1 => n13266, A2 => n1079, ZN => n36080);
   U17528 : NOR2_X2 port map( A1 => n12955, A2 => n10569, ZN => n12954);
   U8412 : OAI21_X2 port map( A1 => n23588, A2 => n19686, B => n37757, ZN => 
                           n8046);
   U9898 : NOR2_X2 port map( A1 => n23620, A2 => n33080, ZN => n9587);
   U6873 : BUF_X2 port map( I => n13779, Z => n31385);
   U24081 : INV_X2 port map( I => n13635, ZN => n17691);
   U247 : NAND2_X2 port map( A1 => n35479, A2 => n35478, ZN => n30786);
   U2312 : CLKBUF_X4 port map( I => n18525, Z => n20525);
   U25847 : INV_X4 port map( I => n1257, ZN => n25467);
   U167 : NOR2_X2 port map( A1 => n14437, A2 => n29937, ZN => n12275);
   U2213 : INV_X4 port map( I => n1109, ZN => n25661);
   U21661 : INV_X2 port map( I => n9539, ZN => n11598);
   U17981 : NAND2_X2 port map( A1 => n24244, A2 => n11673, ZN => n30526);
   U14842 : INV_X4 port map( I => n2393, ZN => n24327);
   U10361 : NAND2_X2 port map( A1 => n36728, A2 => n35116, ZN => n21945);
   U24378 : NAND2_X2 port map( A1 => n18524, A2 => n4664, ZN => n17232);
   U24896 : OAI22_X2 port map( A1 => n18734, A2 => n19637, B1 => n25386, B2 => 
                           n4048, ZN => n18524);
   U30001 : NOR2_X2 port map( A1 => n13491, A2 => n37671, ZN => n3234);
   U10331 : BUF_X4 port map( I => n35828, Z => n34399);
   U22940 : INV_X4 port map( I => n8042, ZN => n33104);
   U4657 : OAI22_X2 port map( A1 => n10160, A2 => n37525, B1 => n35901, B2 => 
                           n10161, ZN => n10159);
   U7969 : OAI21_X2 port map( A1 => n17179, A2 => n10807, B => n17178, ZN => 
                           n25441);
   U5721 : AOI21_X2 port map( A1 => n26805, A2 => n26804, B => n13713, ZN => 
                           n20245);
   U5393 : BUF_X4 port map( I => n28550, Z => n29596);
   U10376 : OAI21_X2 port map( A1 => n21751, A2 => n17102, B => n21889, ZN => 
                           n5979);
   U17679 : OAI21_X2 port map( A1 => n38100, A2 => n15555, B => n7024, ZN => 
                           n35191);
   U1265 : OAI21_X2 port map( A1 => n20105, A2 => n31131, B => n32722, ZN => 
                           n31634);
   U13030 : INV_X2 port map( I => n39815, ZN => n8581);
   U16389 : NOR2_X2 port map( A1 => n28051, A2 => n19750, ZN => n10516);
   U24736 : INV_X2 port map( I => n35116, ZN => n20242);
   U6633 : INV_X4 port map( I => n28238, ZN => n2740);
   U21976 : OAI21_X1 port map( A1 => n15967, A2 => n13411, B => n22258, ZN => 
                           n22767);
   U6032 : NAND2_X2 port map( A1 => n7608, A2 => n5305, ZN => n22197);
   U9334 : NOR2_X2 port map( A1 => n39117, A2 => n1008, ZN => n12173);
   U20405 : NAND2_X2 port map( A1 => n14085, A2 => n37075, ZN => n14084);
   U5172 : INV_X2 port map( I => n15423, ZN => n23380);
   U7407 : AOI21_X2 port map( A1 => n32961, A2 => n27391, B => n13699, ZN => 
                           n14797);
   U835 : NAND3_X2 port map( A1 => n33333, A2 => n4007, A3 => n26933, ZN => 
                           n26644);
   U13686 : NOR2_X2 port map( A1 => n5932, A2 => n34776, ZN => n17221);
   U11810 : NAND2_X2 port map( A1 => n20562, A2 => n26610, ZN => n7855);
   U16642 : NAND2_X1 port map( A1 => n17811, A2 => n35122, ZN => n24380);
   U12311 : INV_X2 port map( I => n25470, ZN => n2962);
   U7028 : NAND2_X2 port map( A1 => n1257, A2 => n10004, ZN => n25470);
   U13024 : BUF_X2 port map( I => n18269, Z => n10008);
   U24401 : NOR2_X1 port map( A1 => n15206, A2 => n15205, ZN => n15223);
   U3969 : NOR2_X2 port map( A1 => n32488, A2 => n36634, ZN => n10374);
   U3952 : BUF_X4 port map( I => n16174, Z => n2771);
   U18553 : NOR2_X2 port map( A1 => n5707, A2 => n5706, ZN => n28713);
   U25670 : INV_X1 port map( I => n17197, ZN => n28192);
   U18765 : NOR2_X2 port map( A1 => n32944, A2 => n12056, ZN => n31810);
   U3548 : CLKBUF_X4 port map( I => n3903, Z => n32012);
   U3312 : CLKBUF_X4 port map( I => n21567, Z => n3293);
   U30070 : INV_X4 port map( I => n37107, ZN => n33580);
   U12637 : NOR2_X2 port map( A1 => n10606, A2 => n10605, ZN => n31060);
   U886 : INV_X2 port map( I => n7377, ZN => n24896);
   U1270 : NAND3_X2 port map( A1 => n7026, A2 => n7025, A3 => n6366, ZN => 
                           n6860);
   U18192 : AOI21_X2 port map( A1 => n1404, A2 => n29486, B => n31667, ZN => 
                           n33425);
   U11967 : BUF_X2 port map( I => n26512, Z => n26934);
   U1349 : INV_X2 port map( I => n16678, ZN => n23011);
   U11965 : BUF_X2 port map( I => n26779, Z => n5537);
   U3713 : OAI22_X2 port map( A1 => n27300, A2 => n36989, B1 => n27171, B2 => 
                           n27170, ZN => n27172);
   U8197 : INV_X4 port map( I => n9526, ZN => n1115);
   U25231 : BUF_X2 port map( I => n17915, Z => n32924);
   U2388 : INV_X2 port map( I => n18204, ZN => n1630);
   U7272 : NAND2_X1 port map( A1 => n9614, A2 => n36321, ZN => n9612);
   U12025 : NOR2_X2 port map( A1 => n4794, A2 => n6062, ZN => n8135);
   U4681 : OR3_X1 port map( A1 => n33333, A2 => n26932, A3 => n37235, Z => 
                           n32072);
   U2996 : NAND2_X2 port map( A1 => n6366, A2 => n8245, ZN => n8594);
   U161 : NAND2_X2 port map( A1 => n14178, A2 => n14179, ZN => n8726);
   U17632 : INV_X4 port map( I => n19544, ZN => n31603);
   U976 : NAND2_X2 port map( A1 => n30348, A2 => n38238, ZN => n17739);
   U7986 : NAND3_X2 port map( A1 => n26076, A2 => n11807, A3 => n26077, ZN => 
                           n7171);
   U3363 : BUF_X4 port map( I => n17810, Z => n33101);
   U21858 : INV_X2 port map( I => n37498, ZN => n25316);
   U1140 : AOI21_X2 port map( A1 => n25996, A2 => n25995, B => n37211, ZN => 
                           n36949);
   U1225 : BUF_X2 port map( I => n2349, Z => n586);
   U618 : INV_X2 port map( I => n37104, ZN => n7195);
   U919 : OAI21_X2 port map( A1 => n26805, A2 => n13713, B => n1091, ZN => 
                           n31447);
   U15833 : INV_X4 port map( I => n34813, ZN => n916);
   U5644 : INV_X2 port map( I => n4458, ZN => n13713);
   U1614 : NAND2_X2 port map( A1 => n6696, A2 => n591, ZN => n14443);
   U4909 : BUF_X4 port map( I => n13973, Z => n1890);
   U18222 : INV_X2 port map( I => n10143, ZN => n35313);
   U2761 : AOI21_X2 port map( A1 => n15084, A2 => n33745, B => n35564, ZN => 
                           n15082);
   U2448 : NAND2_X2 port map( A1 => n18244, A2 => n23101, ZN => n35528);
   U883 : NOR2_X2 port map( A1 => n4748, A2 => n18870, ZN => n2339);
   U2023 : INV_X2 port map( I => n27385, ZN => n19132);
   U796 : NOR2_X2 port map( A1 => n31710, A2 => n31708, ZN => n34776);
   U12396 : NOR2_X1 port map( A1 => n7583, A2 => n35271, ZN => n1873);
   U7234 : NOR2_X2 port map( A1 => n26794, A2 => n925, ZN => n12172);
   U6161 : BUF_X4 port map( I => n3092, Z => n2035);
   U3982 : NOR2_X1 port map( A1 => n20363, A2 => n20362, ZN => n14351);
   U6503 : INV_X2 port map( I => n17127, ZN => n18867);
   U17097 : NAND2_X2 port map( A1 => n17693, A2 => n16271, ZN => n17711);
   U26779 : INV_X4 port map( I => n36361, ZN => n14501);
   U1575 : NAND2_X2 port map( A1 => n24612, A2 => n6977, ZN => n32367);
   U1258 : NOR2_X1 port map( A1 => n32510, A2 => n26134, ZN => n6749);
   U5423 : AOI21_X2 port map( A1 => n30740, A2 => n28480, B => n3532, ZN => 
                           n34266);
   U4817 : BUF_X2 port map( I => n8365, Z => n591);
   U9387 : OAI22_X2 port map( A1 => n1242, A2 => n5883, B1 => n1523, B2 => 
                           n5882, ZN => n5881);
   U9279 : NAND2_X2 port map( A1 => n16267, A2 => n22352, ZN => n3972);
   U9999 : OAI22_X2 port map( A1 => n18072, A2 => n22799, B1 => n22800, B2 => 
                           n23209, ZN => n22801);
   U7267 : INV_X2 port map( I => n21912, ZN => n1155);
   U18123 : INV_X2 port map( I => n5131, ZN => n19587);
   U18540 : AOI22_X2 port map( A1 => n39365, A2 => n37880, B1 => n37981, B2 => 
                           n28302, ZN => n28304);
   U10893 : INV_X1 port map( I => n29900, ZN => n6204);
   U6353 : INV_X1 port map( I => n21687, ZN => n6234);
   U554 : INV_X2 port map( I => n26802, ZN => n26804);
   U23858 : NAND2_X1 port map( A1 => n32743, A2 => n39595, ZN => n33302);
   U12245 : NOR2_X2 port map( A1 => n12096, A2 => n12097, ZN => n31028);
   U9095 : NOR2_X2 port map( A1 => n30952, A2 => n30951, ZN => n18891);
   U17524 : INV_X2 port map( I => n31584, ZN => n31585);
   U11503 : AOI21_X1 port map( A1 => n36969, A2 => n27214, B => n2922, ZN => 
                           n8645);
   U7446 : NOR2_X2 port map( A1 => n1200, A2 => n4457, ZN => n32585);
   U10975 : NOR2_X1 port map( A1 => n14787, A2 => n14773, ZN => n31717);
   U12131 : NAND2_X2 port map( A1 => n491, A2 => n18420, ZN => n31795);
   U6656 : NAND2_X2 port map( A1 => n8197, A2 => n1831, ZN => n7025);
   U10316 : AOI21_X2 port map( A1 => n21909, A2 => n21462, B => n668, ZN => 
                           n7526);
   U16553 : BUF_X2 port map( I => n38901, Z => n15996);
   U1100 : INV_X2 port map( I => n8193, ZN => n20537);
   U8671 : AOI21_X2 port map( A1 => n6349, A2 => n6350, B => n21561, ZN => 
                           n6348);
   U9244 : OAI21_X1 port map( A1 => n30942, A2 => n1493, B => n4651, ZN => 
                           n11306);
   U724 : INV_X2 port map( I => n13712, ZN => n14228);
   U27468 : NOR2_X2 port map( A1 => n35839, A2 => n19084, ZN => n21943);
   U18100 : INV_X2 port map( I => n24419, ZN => n16917);
   U28291 : INV_X2 port map( I => n21602, ZN => n21662);
   U4607 : NAND2_X2 port map( A1 => n5662, A2 => n38566, ZN => n36615);
   U26165 : NOR2_X2 port map( A1 => n21987, A2 => n22342, ZN => n22345);
   U3256 : NOR2_X2 port map( A1 => n24694, A2 => n24590, ZN => n24576);
   U17051 : INV_X1 port map( I => n9828, ZN => n35175);
   U13887 : NAND2_X2 port map( A1 => n21580, A2 => n1847, ZN => n10652);
   U7129 : AOI21_X2 port map( A1 => n25979, A2 => n34265, B => n37175, ZN => 
                           n25984);
   U17137 : OR2_X1 port map( A1 => n33561, A2 => n17022, Z => n20666);
   U20873 : CLKBUF_X4 port map( I => n19713, Z => n35560);
   U12626 : OR3_X2 port map( A1 => n19586, A2 => n31093, A3 => n33745, Z => 
                           n22820);
   U9570 : BUF_X4 port map( I => n13410, Z => n9526);
   U10499 : NAND2_X1 port map( A1 => n37228, A2 => n13817, ZN => n20969);
   U3291 : INV_X4 port map( I => n5089, ZN => n30851);
   U27549 : INV_X2 port map( I => n19298, ZN => n26932);
   U4697 : INV_X4 port map( I => n22307, ZN => n4200);
   U13183 : OAI22_X2 port map( A1 => n20278, A2 => n37014, B1 => n20620, B2 => 
                           n22987, ZN => n7041);
   U4932 : NOR2_X2 port map( A1 => n19549, A2 => n16305, ZN => n21336);
   U797 : NAND2_X2 port map( A1 => n27347, A2 => n19477, ZN => n8165);
   U25461 : INV_X1 port map( I => n25412, ZN => n17020);
   U27706 : INV_X2 port map( I => n21869, ZN => n21570);
   U12063 : NAND3_X2 port map( A1 => n34116, A2 => n1781, A3 => n1777, ZN => 
                           n22742);
   U17311 : INV_X2 port map( I => n197, ZN => n35176);
   U4992 : INV_X2 port map( I => n4210, ZN => n15513);
   U12867 : NAND2_X2 port map( A1 => n18256, A2 => n15143, ZN => n16744);
   U24787 : NAND2_X2 port map( A1 => n19697, A2 => n12392, ZN => n19530);
   U6048 : INV_X2 port map( I => n20778, ZN => n14499);
   U2173 : OAI21_X2 port map( A1 => n9669, A2 => n9670, B => n20588, ZN => 
                           n17819);
   U1527 : INV_X2 port map( I => n21484, ZN => n9670);
   U12501 : INV_X2 port map( I => n20333, ZN => n16673);
   U4309 : INV_X2 port map( I => n24817, ZN => n24828);
   U15603 : NOR2_X2 port map( A1 => n35019, A2 => n22030, ZN => n35818);
   U2948 : NAND2_X2 port map( A1 => n8734, A2 => n28725, ZN => n8733);
   U5573 : OAI21_X2 port map( A1 => n30696, A2 => n30695, B => n26004, ZN => 
                           n16118);
   U1474 : INV_X2 port map( I => n19543, ZN => n6504);
   U242 : AOI21_X2 port map( A1 => n37018, A2 => n28448, B => n979, ZN => 
                           n13806);
   U5543 : NAND2_X1 port map( A1 => n33887, A2 => n34037, ZN => n10949);
   U18695 : NOR2_X2 port map( A1 => n15155, A2 => n32114, ZN => n32113);
   U829 : NAND3_X2 port map( A1 => n10567, A2 => n10098, A3 => n17047, ZN => 
                           n18605);
   U30485 : NAND2_X2 port map( A1 => n6615, A2 => n16834, ZN => n10098);
   U5298 : OAI21_X2 port map( A1 => n21661, A2 => n21946, B => n32664, ZN => 
                           n15805);
   U22541 : NAND2_X1 port map( A1 => n28770, A2 => n28769, ZN => n10596);
   U7487 : AOI22_X2 port map( A1 => n32324, A2 => n2876, B1 => n32705, B2 => 
                           n39132, ZN => n2873);
   U17811 : OR2_X1 port map( A1 => n3827, A2 => n3826, Z => n3825);
   U426 : NAND2_X2 port map( A1 => n17735, A2 => n33765, ZN => n14737);
   U2642 : CLKBUF_X4 port map( I => n7062, Z => n35071);
   U20317 : INV_X2 port map( I => n26512, ZN => n26937);
   U825 : NAND2_X2 port map( A1 => n26774, A2 => n3919, ZN => n3918);
   U18052 : INV_X1 port map( I => n11297, ZN => n17535);
   U1014 : BUF_X4 port map( I => n26485, Z => n33194);
   U29427 : NAND2_X2 port map( A1 => n30629, A2 => n17458, ZN => n25889);
   U7957 : INV_X1 port map( I => n25261, ZN => n3568);
   U2773 : NAND2_X2 port map( A1 => n28544, A2 => n13372, ZN => n34870);
   U24516 : NOR2_X2 port map( A1 => n15314, A2 => n32849, ZN => n8595);
   U7722 : INV_X2 port map( I => n28205, ZN => n1438);
   U2189 : NOR2_X2 port map( A1 => n39666, A2 => n12144, ZN => n33226);
   U16786 : INV_X2 port map( I => n6548, ZN => n11375);
   U6281 : INV_X2 port map( I => n2186, ZN => n35019);
   U11781 : INV_X4 port map( I => n27184, ZN => n30986);
   U9382 : AOI21_X2 port map( A1 => n26083, A2 => n4163, B => n3277, ZN => 
                           n9174);
   U18471 : INV_X2 port map( I => n37094, ZN => n17117);
   U811 : NAND3_X2 port map( A1 => n30851, A2 => n35904, A3 => n27081, ZN => 
                           n30556);
   U2287 : CLKBUF_X4 port map( I => n23523, Z => n30835);
   U23582 : OR2_X2 port map( A1 => n10379, A2 => n37043, Z => n10378);
   U8168 : CLKBUF_X4 port map( I => n38197, Z => n10055);
   U13618 : BUF_X4 port map( I => n22573, Z => n9874);
   U9497 : NOR2_X2 port map( A1 => n13218, A2 => n19367, ZN => n13197);
   U23019 : NAND2_X2 port map( A1 => n11484, A2 => n12446, ZN => n15287);
   U3003 : INV_X4 port map( I => n23108, ZN => n1142);
   U10229 : INV_X2 port map( I => n20397, ZN => n19778);
   U27068 : BUF_X4 port map( I => n23108, Z => n33196);
   U14277 : NAND2_X2 port map( A1 => n19028, A2 => n1597, ZN => n13026);
   U22577 : INV_X2 port map( I => n10655, ZN => n17237);
   U23963 : INV_X2 port map( I => n13417, ZN => n20018);
   U1592 : INV_X4 port map( I => n24694, ZN => n9656);
   U4652 : BUF_X2 port map( I => n30447, Z => n545);
   U1739 : NAND3_X2 port map( A1 => n7847, A2 => n18509, A3 => n37389, ZN => 
                           n13629);
   U22895 : NOR2_X2 port map( A1 => n37033, A2 => n37032, ZN => n14813);
   U3135 : OAI21_X2 port map( A1 => n12983, A2 => n3101, B => n1116, ZN => 
                           n17173);
   U2767 : NAND2_X2 port map( A1 => n31283, A2 => n5570, ZN => n29188);
   U11952 : BUF_X2 port map( I => n26919, Z => n13392);
   U1087 : INV_X2 port map( I => n6130, ZN => n26573);
   U6374 : INV_X2 port map( I => n2147, ZN => n28750);
   U6761 : INV_X2 port map( I => n9518, ZN => n9154);
   U8315 : NAND2_X2 port map( A1 => n34216, A2 => n38687, ZN => n22303);
   U1688 : OAI21_X2 port map( A1 => n38702, A2 => n15049, B => n17163, ZN => 
                           n33187);
   U2229 : NAND2_X2 port map( A1 => n23039, A2 => n17995, ZN => n15799);
   U924 : NAND2_X2 port map( A1 => n26810, A2 => n14377, ZN => n26812);
   U16861 : NOR2_X2 port map( A1 => n35135, A2 => n30384, ZN => n33755);
   U16864 : NAND2_X2 port map( A1 => n4321, A2 => n18744, ZN => n35135);
   U8716 : NOR2_X2 port map( A1 => n14499, A2 => n21521, ZN => n21412);
   U17723 : NAND2_X2 port map( A1 => n2878, A2 => n11283, ZN => n2874);
   U287 : NOR2_X2 port map( A1 => n17532, A2 => n32705, ZN => n2878);
   U13281 : INV_X2 port map( I => n23039, ZN => n11797);
   U9 : INV_X2 port map( I => n20437, ZN => n29570);
   U5489 : INV_X2 port map( I => n25509, ZN => n33834);
   U27814 : INV_X4 port map( I => n15102, ZN => n16460);
   U4483 : INV_X1 port map( I => n20566, ZN => n5384);
   U19771 : OAI21_X2 port map( A1 => n27278, A2 => n9875, B => n38305, ZN => 
                           n7694);
   U1531 : INV_X2 port map( I => n21857, ZN => n21860);
   U12137 : NAND2_X2 port map( A1 => n1012, A2 => n6506, ZN => n8236);
   U23407 : NAND2_X2 port map( A1 => n18188, A2 => n19410, ZN => n28119);
   U11905 : NAND2_X2 port map( A1 => n5997, A2 => n5998, ZN => n34836);
   U9841 : NAND3_X2 port map( A1 => n18155, A2 => n23459, A3 => n35808, ZN => 
                           n23241);
   U5687 : BUF_X4 port map( I => n25720, Z => n18519);
   U18131 : AOI21_X1 port map( A1 => n5145, A2 => n29813, B => n5144, ZN => 
                           n5143);
   U15731 : NOR2_X2 port map( A1 => n33270, A2 => n831, ZN => n4952);
   U622 : OAI21_X2 port map( A1 => n31000, A2 => n11088, B => n35114, ZN => 
                           n11087);
   U10036 : AOI22_X2 port map( A1 => n19054, A2 => n33969, B1 => n38752, B2 => 
                           n1653, ZN => n18748);
   U1566 : OR2_X2 port map( A1 => n15159, A2 => n30844, Z => n12705);
   U12252 : NAND2_X1 port map( A1 => n12780, A2 => n12779, ZN => n12778);
   U7202 : INV_X4 port map( I => n10440, ZN => n30795);
   U18567 : INV_X2 port map( I => n19473, ZN => n24309);
   U24402 : NOR2_X2 port map( A1 => n277, A2 => n24168, ZN => n24182);
   U14366 : INV_X4 port map( I => n2416, ZN => n25622);
   U199 : INV_X1 port map( I => n11348, ZN => n35870);
   U24756 : OAI21_X2 port map( A1 => n18408, A2 => n1676, B => n17869, ZN => 
                           n17557);
   U2671 : NOR2_X2 port map( A1 => n10441, A2 => n10442, ZN => n35038);
   U22419 : INV_X2 port map( I => n39096, ZN => n22937);
   U17684 : OAI21_X2 port map( A1 => n38100, A2 => n15555, B => n7024, ZN => 
                           n35192);
   U3356 : INV_X2 port map( I => n12856, ZN => n17810);
   U8687 : OAI21_X2 port map( A1 => n21551, A2 => n21763, B => n33771, ZN => 
                           n6670);
   U17635 : BUF_X4 port map( I => n21608, Z => n12144);
   U1925 : AOI21_X2 port map( A1 => n34046, A2 => n33513, B => n35086, ZN => 
                           n5330);
   U12417 : NAND2_X2 port map( A1 => n19767, A2 => n32722, ZN => n4454);
   U2823 : BUF_X4 port map( I => n33417, Z => n32131);
   U17634 : INV_X2 port map( I => n21608, ZN => n17233);
   U4245 : NOR2_X2 port map( A1 => n12144, A2 => n21779, ZN => n21535);
   U11213 : NOR2_X2 port map( A1 => n17615, A2 => n32352, ZN => n17085);
   U9411 : AOI21_X2 port map( A1 => n12457, A2 => n25751, B => n1522, ZN => 
                           n12456);
   U4919 : NAND3_X2 port map( A1 => n21788, A2 => n32456, A3 => n21787, ZN => 
                           n16951);
   U11913 : NOR2_X2 port map( A1 => n7978, A2 => n26703, ZN => n13644);
   U8907 : INV_X2 port map( I => n29777, ZN => n1402);
   U13724 : NAND2_X1 port map( A1 => n1838, A2 => n554, ZN => n1837);
   U10418 : BUF_X2 port map( I => n15354, Z => n11274);
   U2257 : OAI21_X2 port map( A1 => n21208, A2 => n37012, B => n17167, ZN => 
                           n12268);
   U9858 : AOI21_X2 port map( A1 => n23462, A2 => n1140, B => n5083, ZN => 
                           n23299);
   U1377 : OR2_X2 port map( A1 => n25351, A2 => n18121, Z => n19264);
   U15862 : INV_X4 port map( I => n1606, ZN => n9547);
   U3705 : INV_X2 port map( I => n33997, ZN => n1107);
   U4444 : AOI21_X2 port map( A1 => n14810, A2 => n26110, B => n33753, ZN => 
                           n33752);
   U4243 : BUF_X2 port map( I => n21857, Z => n455);
   U5548 : INV_X2 port map( I => n26018, ZN => n1239);
   U1911 : INV_X2 port map( I => n24732, ZN => n24839);
   U17362 : INV_X2 port map( I => n20208, ZN => n35180);
   U15281 : OAI21_X2 port map( A1 => n2812, A2 => n38748, B => n36210, ZN => 
                           n2813);
   U27275 : OAI21_X2 port map( A1 => n21588, A2 => n19397, B => n17792, ZN => 
                           n18560);
   U10447 : BUF_X2 port map( I => Key(143), Z => n29647);
   U3165 : BUF_X2 port map( I => n21270, Z => n32720);
   U4868 : BUF_X4 port map( I => n5988, Z => n36854);
   U20147 : NAND2_X2 port map( A1 => n32041, A2 => n32040, ZN => n23065);
   U13343 : INV_X2 port map( I => n4847, ZN => n33893);
   U6306 : INV_X4 port map( I => n19915, ZN => n1127);
   U17411 : NAND2_X2 port map( A1 => n22342, A2 => n17074, ZN => n21966);
   U6507 : INV_X2 port map( I => n17074, ZN => n22171);
   U6718 : AOI21_X2 port map( A1 => n22803, A2 => n5657, B => n8461, ZN => 
                           n8460);
   U20454 : INV_X4 port map( I => n16200, ZN => n10807);
   U15541 : INV_X4 port map( I => n585, ZN => n5572);
   U2249 : AOI22_X2 port map( A1 => n18606, A2 => n26740, B1 => n6615, B2 => 
                           n18706, ZN => n30585);
   U2754 : NOR3_X2 port map( A1 => n1417, A2 => n209, A3 => n1192, ZN => n5156)
                           ;
   U8956 : NOR2_X2 port map( A1 => n27653, A2 => n11412, ZN => n14237);
   U5954 : NAND2_X2 port map( A1 => n978, A2 => n13508, ZN => n32004);
   U4693 : AOI21_X2 port map( A1 => n37737, A2 => n24746, B => n32882, ZN => 
                           n2549);
   U7489 : BUF_X2 port map( I => n8944, Z => n36796);
   U4614 : AOI22_X2 port map( A1 => n9352, A2 => n38566, B1 => n9353, B2 => 
                           n10618, ZN => n33686);
   U2533 : BUF_X4 port map( I => n19712, Z => n31157);
   U30561 : INV_X2 port map( I => n8556, ZN => n2292);
   U2712 : NOR2_X2 port map( A1 => n12702, A2 => n12703, ZN => n56);
   U19298 : INV_X2 port map( I => n6591, ZN => n19589);
   U4899 : INV_X4 port map( I => n14378, ZN => n1597);
   U1065 : BUF_X4 port map( I => n18500, Z => n17194);
   U7256 : NOR2_X1 port map( A1 => n17617, A2 => n5405, ZN => n36307);
   U395 : INV_X2 port map( I => n36791, ZN => n13133);
   U1267 : NAND2_X2 port map( A1 => n26119, A2 => n7423, ZN => n35401);
   U13658 : NOR2_X2 port map( A1 => n11012, A2 => n21965, ZN => n9343);
   U9987 : NAND2_X2 port map( A1 => n22959, A2 => n11157, ZN => n11156);
   U9197 : NAND2_X1 port map( A1 => n18730, A2 => n1331, ZN => n31860);
   U10552 : OAI22_X1 port map( A1 => n25363, A2 => n424, B1 => n9568, B2 => 
                           n26090, ZN => n34413);
   U12706 : CLKBUF_X8 port map( I => n2634, Z => n2340);
   U25964 : OAI21_X2 port map( A1 => n12477, A2 => n13081, B => n37057, ZN => 
                           n36266);
   U12801 : OAI21_X2 port map( A1 => n28590, A2 => n3598, B => n14701, ZN => 
                           n35961);
   U8847 : NAND2_X2 port map( A1 => n31583, A2 => n37061, ZN => n20371);
   U3650 : NAND3_X2 port map( A1 => n32712, A2 => n27146, A3 => n27354, ZN => 
                           n36492);
   U30348 : NOR2_X1 port map( A1 => n9056, A2 => n154, ZN => n36834);
   U13033 : OR3_X2 port map( A1 => n18342, A2 => n12951, A3 => n11795, Z => 
                           n7279);
   U1794 : BUF_X2 port map( I => n30454, Z => n33240);
   U2217 : AOI22_X2 port map( A1 => n23253, A2 => n23610, B1 => n9639, B2 => 
                           n1132, ZN => n33702);
   U18766 : NOR2_X1 port map( A1 => n32619, A2 => n32618, ZN => n3761);
   U8616 : NAND2_X1 port map( A1 => n23548, A2 => n23472, ZN => n2688);
   U1112 : NOR2_X2 port map( A1 => n6104, A2 => n6103, ZN => n6154);
   U8261 : OAI21_X1 port map( A1 => n4531, A2 => n32703, B => n32702, ZN => 
                           n10640);
   U19812 : NAND2_X2 port map( A1 => n15121, A2 => n1101, ZN => n7135);
   U179 : INV_X2 port map( I => n36595, ZN => n3633);
   U128 : INV_X4 port map( I => n37100, ZN => n29446);
   U2343 : NOR3_X2 port map( A1 => n14396, A2 => n19538, A3 => n31093, ZN => 
                           n35564);
   U3860 : BUF_X2 port map( I => n29307, Z => n29498);
   U689 : OR2_X2 port map( A1 => n27108, A2 => n6686, Z => n30434);
   U13020 : OR2_X2 port map( A1 => n10733, A2 => n14290, Z => n15775);
   U1290 : NAND2_X2 port map( A1 => n32436, A2 => n260, ZN => n31964);
   U21579 : NAND2_X2 port map( A1 => n35665, A2 => n34087, ZN => n32436);
   U23324 : INV_X4 port map( I => n12066, ZN => n12065);
   U26021 : NAND2_X1 port map( A1 => n33054, A2 => n33052, ZN => n33051);
   U6860 : INV_X2 port map( I => n17915, ZN => n1528);
   U28144 : NAND2_X2 port map( A1 => n19238, A2 => n17112, ZN => n21511);
   U7081 : INV_X2 port map( I => n32377, ZN => n23579);
   U908 : INV_X2 port map( I => n10987, ZN => n3426);
   U27577 : INV_X2 port map( I => n16835, ZN => n19334);
   U1664 : NAND2_X2 port map( A1 => n32831, A2 => n24878, ZN => n8125);
   U12267 : OAI21_X2 port map( A1 => n25687, A2 => n25686, B => n25685, ZN => 
                           n20008);
   U7494 : NOR2_X2 port map( A1 => n11412, A2 => n11164, ZN => n11163);
   U20357 : NOR2_X1 port map( A1 => n32950, A2 => n6534, ZN => n35466);
   U3496 : CLKBUF_X4 port map( I => n9847, Z => n2018);
   U17621 : INV_X1 port map( I => n38199, ZN => n26754);
   U3984 : BUF_X4 port map( I => n33987, Z => n33986);
   U9688 : OAI21_X2 port map( A1 => n19027, A2 => n13026, B => n19026, ZN => 
                           n23754);
   U5631 : NAND2_X2 port map( A1 => n26696, A2 => n923, ZN => n4583);
   U21152 : NOR2_X2 port map( A1 => n17040, A2 => n7730, ZN => n8682);
   U1128 : NAND2_X2 port map( A1 => n20088, A2 => n26021, ZN => n33423);
   U3975 : NAND2_X2 port map( A1 => n34969, A2 => n8537, ZN => n13364);
   U1347 : NOR2_X2 port map( A1 => n37238, A2 => n5798, ZN => n13034);
   U2416 : INV_X2 port map( I => n12909, ZN => n14461);
   U3919 : NAND2_X1 port map( A1 => n27114, A2 => n33088, ZN => n32757);
   U1313 : NAND2_X2 port map( A1 => n8006, A2 => n17008, ZN => n7941);
   U9327 : INV_X2 port map( I => n1091, ZN => n10890);
   U7490 : INV_X2 port map( I => n15187, ZN => n18667);
   U2709 : CLKBUF_X4 port map( I => n22854, Z => n22993);
   U7310 : BUF_X2 port map( I => Key(51), Z => n29223);
   U5332 : INV_X1 port map( I => n37916, ZN => n1279);
   U313 : OAI21_X2 port map( A1 => n20188, A2 => n33842, B => n21239, ZN => 
                           n14330);
   U4042 : OAI21_X2 port map( A1 => n1112, A2 => n7866, B => n33950, ZN => 
                           n11332);
   U8188 : INV_X4 port map( I => n25692, ZN => n1112);
   U5006 : NAND2_X2 port map( A1 => n21806, A2 => n36735, ZN => n21274);
   U11830 : AOI21_X2 port map( A1 => n3125, A2 => n35960, B => n3124, ZN => 
                           n35022);
   U2610 : NOR2_X2 port map( A1 => n123, A2 => n19545, ZN => n9041);
   U3623 : NAND2_X2 port map( A1 => n22080, A2 => n38337, ZN => n4337);
   U10888 : INV_X2 port map( I => n11573, ZN => n30220);
   U13567 : INV_X2 port map( I => n20077, ZN => n1653);
   U7002 : NAND3_X1 port map( A1 => n24269, A2 => n24444, A3 => n24311, ZN => 
                           n11104);
   U272 : AOI21_X2 port map( A1 => n27996, A2 => n16461, B => n27995, ZN => 
                           n28002);
   U4425 : NOR2_X2 port map( A1 => n2078, A2 => n3541, ZN => n2077);
   U8187 : INV_X1 port map( I => n37604, ZN => n32634);
   U22313 : NAND2_X2 port map( A1 => n17501, A2 => n32747, ZN => n10224);
   U4090 : AND3_X1 port map( A1 => n24812, A2 => n24565, A3 => n19294, Z => 
                           n14532);
   U840 : INV_X4 port map( I => n25487, ZN => n1535);
   U2320 : INV_X2 port map( I => n23296, ZN => n35808);
   U5454 : AOI21_X1 port map( A1 => n15372, A2 => n28220, B => n11650, ZN => 
                           n11649);
   U14028 : CLKBUF_X2 port map( I => Key(44), Z => n30090);
   U14385 : INV_X2 port map( I => n2000, ZN => n13758);
   U12324 : NOR2_X2 port map( A1 => n8222, A2 => n7866, ZN => n8221);
   U25311 : NAND2_X2 port map( A1 => n28361, A2 => n28362, ZN => n18836);
   U8719 : NOR2_X2 port map( A1 => n14499, A2 => n8597, ZN => n8599);
   U6769 : INV_X4 port map( I => n14488, ZN => n26823);
   U16404 : NAND2_X1 port map( A1 => n35447, A2 => n20306, ZN => n36972);
   U1918 : NOR2_X2 port map( A1 => n17120, A2 => n9996, ZN => n12669);
   U6267 : AOI21_X2 port map( A1 => n1267, A2 => n2341, B => n1576, ZN => n6636
                           );
   U11337 : OAI21_X2 port map( A1 => n15313, A2 => n28720, B => n37311, ZN => 
                           n15312);
   U4439 : NOR2_X2 port map( A1 => n25586, A2 => n10062, ZN => n32157);
   U12668 : INV_X2 port map( I => n18110, ZN => n16211);
   U16802 : NAND2_X2 port map( A1 => n4345, A2 => n9201, ZN => n3998);
   U3892 : NAND2_X2 port map( A1 => n16922, A2 => n16921, ZN => n16920);
   U9048 : AOI22_X2 port map( A1 => n19139, A2 => n1446, B1 => n20577, B2 => 
                           n28111, ZN => n18309);
   U13295 : INV_X2 port map( I => n23347, ZN => n10048);
   U8382 : CLKBUF_X4 port map( I => n10162, Z => n36422);
   U2872 : CLKBUF_X4 port map( I => n28704, Z => n18281);
   U2457 : BUF_X2 port map( I => n22887, Z => n31300);
   U6118 : BUF_X4 port map( I => n9878, Z => n2937);
   U4395 : NOR2_X2 port map( A1 => n19777, A2 => n5698, ZN => n17841);
   U5785 : INV_X2 port map( I => n18246, ZN => n19564);
   U20025 : AOI22_X2 port map( A1 => n16105, A2 => n16104, B1 => n1316, B2 => 
                           n20173, ZN => n7366);
   U4360 : NOR2_X2 port map( A1 => n7320, A2 => n26304, ZN => n31274);
   U15070 : NAND2_X2 port map( A1 => n6446, A2 => n27070, ZN => n34944);
   U11969 : INV_X1 port map( I => n26358, ZN => n4591);
   U7592 : CLKBUF_X2 port map( I => n14422, Z => n357);
   U8865 : NOR2_X2 port map( A1 => n9394, A2 => n5669, ZN => n30190);
   U6442 : INV_X2 port map( I => n3443, ZN => n9316);
   U2967 : NAND3_X1 port map( A1 => n4919, A2 => n16985, A3 => n20480, ZN => 
                           n32188);
   U9530 : INV_X2 port map( I => n12394, ZN => n1536);
   U12314 : NAND2_X2 port map( A1 => n25444, A2 => n38338, ZN => n9503);
   U9962 : NAND2_X2 port map( A1 => n2049, A2 => n1989, ZN => n5944);
   U13802 : INV_X2 port map( I => n17869, ZN => n17207);
   U16333 : INV_X2 port map( I => n5080, ZN => n25328);
   U6419 : INV_X2 port map( I => n21923, ZN => n1689);
   U5402 : NOR2_X2 port map( A1 => n37852, A2 => n8954, ZN => n8968);
   U28226 : BUF_X4 port map( I => n16760, Z => n33359);
   U2625 : NOR2_X2 port map( A1 => n4759, A2 => n21888, ZN => n21601);
   U2505 : NAND2_X2 port map( A1 => n22342, A2 => n22341, ZN => n10487);
   U2009 : NOR3_X2 port map( A1 => n17127, A2 => n1989, A3 => n37791, ZN => 
                           n33034);
   U7099 : NOR2_X2 port map( A1 => n26135, A2 => n31626, ZN => n15449);
   U5287 : NAND2_X2 port map( A1 => n15240, A2 => n1608, ZN => n20083);
   U565 : INV_X2 port map( I => n33960, ZN => n32977);
   U1185 : OR2_X2 port map( A1 => n34609, A2 => n4553, Z => n25916);
   U1936 : INV_X4 port map( I => n1140, ZN => n32061);
   U11230 : AOI22_X2 port map( A1 => n28759, A2 => n18701, B1 => n1416, B2 => 
                           n30917, ZN => n28761);
   U21369 : OAI21_X1 port map( A1 => n29741, A2 => n29754, B => n29737, ZN => 
                           n29726);
   U18388 : INV_X2 port map( I => n17567, ZN => n17784);
   U6545 : INV_X4 port map( I => n11329, ZN => n8520);
   U20121 : NAND2_X2 port map( A1 => n7062, A2 => n32456, ZN => n21794);
   U3701 : OAI21_X2 port map( A1 => n923, A2 => n37102, B => n26695, ZN => 
                           n16707);
   U12116 : NOR2_X2 port map( A1 => n25758, A2 => n33514, ZN => n2498);
   U17498 : INV_X2 port map( I => n27786, ZN => n18733);
   U7434 : NOR2_X2 port map( A1 => n36197, A2 => n28278, ZN => n7840);
   U27642 : BUF_X4 port map( I => n18342, Z => n33289);
   U7461 : NAND2_X2 port map( A1 => n18461, A2 => n38262, ZN => n18457);
   U24181 : NAND2_X2 port map( A1 => n19043, A2 => n17714, ZN => n13890);
   U15745 : INV_X1 port map( I => n14130, ZN => n23178);
   U30764 : INV_X1 port map( I => n36995, ZN => n30338);
   U6813 : AOI21_X2 port map( A1 => n9892, A2 => n931, B => n7460, ZN => n24968
                           );
   U12532 : NAND3_X1 port map( A1 => n18264, A2 => n24413, A3 => n18263, ZN => 
                           n24415);
   U1208 : NOR2_X2 port map( A1 => n32044, A2 => n2957, ZN => n2955);
   U8260 : NAND2_X2 port map( A1 => n1028, A2 => n24782, ZN => n13415);
   U16321 : INV_X2 port map( I => n9385, ZN => n14211);
   U1072 : INV_X2 port map( I => n18238, ZN => n1591);
   U13291 : OAI21_X2 port map( A1 => n8459, A2 => n8458, B => n19469, ZN => 
                           n4698);
   U28818 : AOI21_X2 port map( A1 => n34906, A2 => n24732, B => n4973, ZN => 
                           n24254);
   U11861 : BUF_X2 port map( I => n27141, Z => n9593);
   U1975 : NOR2_X2 port map( A1 => n5942, A2 => n5943, ZN => n5946);
   U12443 : NAND2_X2 port map( A1 => n25467, A2 => n38210, ZN => n14679);
   U8096 : NAND2_X1 port map( A1 => n17038, A2 => n17020, ZN => n17037);
   U16531 : OAI21_X2 port map( A1 => n1689, A2 => n9316, B => n37612, ZN => 
                           n4057);
   U7438 : NAND2_X2 port map( A1 => n28214, A2 => n11512, ZN => n18020);
   U22803 : NAND2_X2 port map( A1 => n8385, A2 => n11083, ZN => n13178);
   U17154 : AOI21_X2 port map( A1 => n7767, A2 => n17212, B => n834, ZN => 
                           n25772);
   U4221 : NAND3_X2 port map( A1 => n36638, A2 => n33247, A3 => n3683, ZN => 
                           n31343);
   U8352 : INV_X2 port map( I => n14491, ZN => n24453);
   U2174 : NOR2_X2 port map( A1 => n37190, A2 => n34981, ZN => n4538);
   U24744 : NOR2_X2 port map( A1 => n33709, A2 => n15879, ZN => n7625);
   U8959 : OAI21_X2 port map( A1 => n33424, A2 => n18035, B => n11030, ZN => 
                           n4926);
   U495 : NAND2_X1 port map( A1 => n27981, A2 => n28047, ZN => n36914);
   U27151 : INV_X1 port map( I => n36755, ZN => n36433);
   U27903 : INV_X2 port map( I => n20958, ZN => n23076);
   U3087 : NOR2_X1 port map( A1 => n18884, A2 => n8480, ZN => n16642);
   U4737 : INV_X2 port map( I => n23198, ZN => n1044);
   U12043 : OR2_X1 port map( A1 => n19137, A2 => n16510, Z => n10148);
   U11727 : NOR2_X2 port map( A1 => n4927, A2 => n34569, ZN => n32206);
   U21872 : AOI22_X2 port map( A1 => n18822, A2 => n22892, B1 => n13946, B2 => 
                           n22804, ZN => n32397);
   U13287 : NOR2_X2 port map( A1 => n30386, A2 => n3761, ZN => n36729);
   U6369 : NAND2_X2 port map( A1 => n19375, A2 => n34923, ZN => n21778);
   U5621 : NAND2_X2 port map( A1 => n34658, A2 => n26316, ZN => n31253);
   U12843 : NOR2_X2 port map( A1 => n6914, A2 => n6170, ZN => n6913);
   U347 : INV_X4 port map( I => n20860, ZN => n7872);
   U10032 : NOR2_X2 port map( A1 => n31005, A2 => n20872, ZN => n16892);
   U17394 : INV_X1 port map( I => n26905, ZN => n15485);
   U19238 : AOI21_X2 port map( A1 => n23174, A2 => n3803, B => n20840, ZN => 
                           n11157);
   U11937 : AOI21_X1 port map( A1 => n38548, A2 => n14212, B => n25951, ZN => 
                           n12869);
   U7198 : INV_X1 port map( I => n735, ZN => n26470);
   U4473 : BUF_X2 port map( I => n18062, Z => n31719);
   U1738 : INV_X2 port map( I => n37395, ZN => n34746);
   U7826 : NAND2_X2 port map( A1 => n7612, A2 => n5035, ZN => n5366);
   U15781 : INV_X1 port map( I => n33995, ZN => n31513);
   U26689 : NAND2_X2 port map( A1 => n5366, A2 => n5367, ZN => n5361);
   U14613 : NOR2_X2 port map( A1 => n9587, A2 => n9588, ZN => n34884);
   U18928 : AOI21_X1 port map( A1 => n2681, A2 => n38248, B => n31836, ZN => 
                           n2684);
   U6010 : AOI21_X2 port map( A1 => n17793, A2 => n22108, B => n1684, ZN => 
                           n12155);
   U24726 : INV_X2 port map( I => n22272, ZN => n15029);
   U23396 : NAND2_X2 port map( A1 => n17167, A2 => n12191, ZN => n23334);
   U22203 : OAI21_X2 port map( A1 => n14392, A2 => n24184, B => n35690, ZN => 
                           n10046);
   U2221 : NAND3_X2 port map( A1 => n23494, A2 => n33638, A3 => n36630, ZN => 
                           n23500);
   U575 : INV_X2 port map( I => n38002, ZN => n26840);
   U2063 : NAND2_X2 port map( A1 => n37216, A2 => n36227, ZN => n31168);
   U1261 : INV_X4 port map( I => n23399, ZN => n961);
   U9189 : NAND3_X1 port map( A1 => n28042, A2 => n28043, A3 => n1073, ZN => 
                           n36832);
   U1310 : NOR2_X1 port map( A1 => n832, A2 => n14778, ZN => n30945);
   U11875 : NAND2_X2 port map( A1 => n6909, A2 => n35537, ZN => n12566);
   U29184 : NOR3_X2 port map( A1 => n26240, A2 => n26239, A3 => n26238, ZN => 
                           n26439);
   U6654 : NAND2_X2 port map( A1 => n18948, A2 => n15925, ZN => n18696);
   U29248 : OAI21_X2 port map( A1 => n33689, A2 => n37585, B => n26444, ZN => 
                           n26445);
   U2930 : AOI21_X2 port map( A1 => n14382, A2 => n19728, B => n1500, ZN => 
                           n26444);
   U6647 : NOR2_X2 port map( A1 => n16638, A2 => n22993, ZN => n34643);
   U2116 : OR2_X2 port map( A1 => n30280, A2 => n31278, Z => n15018);
   U506 : OAI21_X2 port map( A1 => n7934, A2 => n8498, B => n28045, ZN => 
                           n27988);
   U21197 : NOR2_X2 port map( A1 => n27507, A2 => n35265, ZN => n35604);
   U11492 : NAND2_X2 port map( A1 => n8092, A2 => n8093, ZN => n34525);
   U29054 : OAI22_X2 port map( A1 => n33428, A2 => n33427, B1 => n29536, B2 => 
                           n29519, ZN => n29510);
   U24877 : NAND3_X2 port map( A1 => n24118, A2 => n24372, A3 => n38609, ZN => 
                           n14895);
   U5915 : INV_X2 port map( I => n26541, ZN => n16169);
   U18303 : BUF_X4 port map( I => n38669, Z => n31088);
   U17576 : INV_X2 port map( I => n4841, ZN => n28238);
   U9581 : NOR2_X2 port map( A1 => n35000, A2 => n33640, ZN => n2328);
   U8854 : NOR2_X2 port map( A1 => n17374, A2 => n19120, ZN => n13388);
   U20065 : NOR2_X2 port map( A1 => n5415, A2 => n8112, ZN => n33281);
   U6554 : AOI21_X2 port map( A1 => n12353, A2 => n5669, B => n30155, ZN => 
                           n8112);
   U15056 : OAI21_X2 port map( A1 => n32802, A2 => n37097, B => n2608, ZN => 
                           n2607);
   U13252 : NAND2_X2 port map( A1 => n14739, A2 => n8146, ZN => n8145);
   U2413 : INV_X2 port map( I => n30304, ZN => n8093);
   U12285 : AOI21_X1 port map( A1 => n33826, A2 => n19237, B => n19236, ZN => 
                           n17868);
   U2201 : NAND2_X2 port map( A1 => n3497, A2 => n15787, ZN => n36394);
   U8423 : OAI21_X2 port map( A1 => n23624, A2 => n35938, B => n3498, ZN => 
                           n3497);
   U3992 : OAI22_X2 port map( A1 => n10906, A2 => n36663, B1 => n18871, B2 => 
                           n10883, ZN => n28314);
   U3396 : AOI22_X2 port map( A1 => n14484, A2 => n19366, B1 => n28148, B2 => 
                           n18392, ZN => n30608);
   U8398 : NOR2_X2 port map( A1 => n1298, A2 => n32351, ZN => n5790);
   U16680 : AOI22_X2 port map( A1 => n12544, A2 => n12543, B1 => n36145, B2 => 
                           n18961, ZN => n12542);
   U20222 : BUF_X4 port map( I => n30504, Z => n35443);
   U13147 : AOI22_X2 port map( A1 => n8390, A2 => n32858, B1 => n23421, B2 => 
                           n1302, ZN => n7482);
   U17287 : BUF_X2 port map( I => n36397, Z => n35754);
   U4688 : OAI21_X1 port map( A1 => n24626, A2 => n24627, B => n9847, ZN => 
                           n13747);
   U28297 : INV_X2 port map( I => n9736, ZN => n22334);
   U15163 : INV_X2 port map( I => n7324, ZN => n31353);
   U26622 : NAND2_X2 port map( A1 => n26964, A2 => n26963, ZN => n17602);
   U1073 : NAND3_X2 port map( A1 => n30665, A2 => n35537, A3 => n1231, ZN => 
                           n26963);
   U27859 : INV_X4 port map( I => n21939, ZN => n36519);
   U4458 : NAND2_X1 port map( A1 => n27011, A2 => n16263, ZN => n8196);
   U12784 : OAI21_X2 port map( A1 => n6175, A2 => n10690, B => n9844, ZN => 
                           n16406);
   U26478 : NAND2_X2 port map( A1 => n5351, A2 => n36325, ZN => n7325);
   U1344 : INV_X1 port map( I => n23102, ZN => n23103);
   U17540 : INV_X2 port map( I => n29555, ZN => n29541);
   U6705 : OAI22_X2 port map( A1 => n22809, A2 => n36554, B1 => n531, B2 => 
                           n23169, ZN => n22812);
   U23409 : NOR2_X2 port map( A1 => n16081, A2 => n24373, ZN => n24191);
   U671 : NAND2_X2 port map( A1 => n26084, A2 => n26114, ZN => n4372);
   U3287 : INV_X4 port map( I => n14729, ZN => n1577);
   U29245 : INV_X2 port map( I => n26439, ZN => n26440);
   U1801 : BUF_X4 port map( I => n39816, Z => n250);
   U30574 : INV_X1 port map( I => n23654, ZN => n238);
   U7060 : INV_X2 port map( I => n23599, ZN => n23601);
   U5864 : INV_X2 port map( I => n20896, ZN => n941);
   U2590 : AOI22_X2 port map( A1 => n8434, A2 => n21834, B1 => n8436, B2 => 
                           n21436, ZN => n34220);
   U25457 : INV_X2 port map( I => n25716, ZN => n25562);
   U2977 : NAND2_X2 port map( A1 => n23308, A2 => n38704, ZN => n23311);
   U5697 : AOI21_X2 port map( A1 => n24708, A2 => n24529, B => n33986, ZN => 
                           n8389);
   U12187 : NOR2_X2 port map( A1 => n26079, A2 => n15283, ZN => n7170);
   U19536 : AOI21_X2 port map( A1 => n30702, A2 => n28133, B => n2870, ZN => 
                           n3070);
   U5437 : NAND2_X1 port map( A1 => n4874, A2 => n13837, ZN => n6556);
   U10037 : OR2_X1 port map( A1 => n1484, A2 => n32870, Z => n16480);
   U9587 : INV_X2 port map( I => n24944, ZN => n13259);
   U1339 : INV_X4 port map( I => n34014, ZN => n9050);
   U105 : INV_X4 port map( I => n8805, ZN => n3986);
   U19058 : NOR2_X1 port map( A1 => n20915, A2 => n14692, ZN => n20914);
   U860 : NOR2_X1 port map( A1 => n20815, A2 => n35271, ZN => n219);
   U12684 : BUF_X4 port map( I => n8805, Z => n34652);
   U14559 : NOR2_X1 port map( A1 => n4459, A2 => n2140, ZN => n10903);
   U19714 : NOR2_X2 port map( A1 => n32543, A2 => n28486, ZN => n8657);
   U1916 : NAND2_X2 port map( A1 => n31945, A2 => n30506, ZN => n32598);
   U866 : NOR2_X2 port map( A1 => n13427, A2 => n4686, ZN => n27044);
   U1558 : BUF_X2 port map( I => n24819, Z => n31714);
   U541 : AOI22_X2 port map( A1 => n13984, A2 => n27969, B1 => n12257, B2 => 
                           n13983, ZN => n14277);
   U27587 : NAND3_X2 port map( A1 => n24906, A2 => n32802, A3 => n24905, ZN => 
                           n24907);
   U4035 : INV_X2 port map( I => n18302, ZN => n20058);
   U4111 : NAND2_X2 port map( A1 => n21117, A2 => n38448, ZN => n2128);
   U1726 : INV_X2 port map( I => n20774, ZN => n1209);
   U183 : NAND2_X2 port map( A1 => n6163, A2 => n8805, ZN => n29992);
   U18027 : BUF_X2 port map( I => Key(99), Z => n30094);
   U17379 : CLKBUF_X4 port map( I => n14462, Z => n12443);
   U4082 : CLKBUF_X4 port map( I => n9383, Z => n1606);
   U1064 : INV_X2 port map( I => n39648, ZN => n7658);
   U17193 : INV_X2 port map( I => n33316, ZN => n36965);
   U6800 : INV_X2 port map( I => n9214, ZN => n26901);
   U780 : NOR2_X2 port map( A1 => n27273, A2 => n27274, ZN => n8382);
   U10909 : INV_X1 port map( I => n7766, ZN => n28947);
   U6603 : BUF_X2 port map( I => n15871, Z => n35532);
   U11801 : NOR2_X1 port map( A1 => n7393, A2 => n7392, ZN => n14966);
   U23787 : NOR2_X2 port map( A1 => n10806, A2 => n39571, ZN => n32727);
   U17347 : NAND2_X2 port map( A1 => n33116, A2 => n8272, ZN => n35529);
   U226 : OAI21_X2 port map( A1 => n18096, A2 => n37295, B => n5662, ZN => 
                           n19726);
   U10110 : INV_X2 port map( I => n23140, ZN => n22949);
   U2766 : AOI21_X2 port map( A1 => n25365, A2 => n25623, B => n1532, ZN => 
                           n3012);
   U7106 : INV_X2 port map( I => n25856, ZN => n26008);
   U20992 : NAND2_X1 port map( A1 => n32215, A2 => n15411, ZN => n11222);
   U6973 : NOR2_X2 port map( A1 => n24824, A2 => n24819, ZN => n24629);
   U26800 : OAI21_X2 port map( A1 => n32425, A2 => n38292, B => n38042, ZN => 
                           n23328);
   U15239 : NAND3_X2 port map( A1 => n16520, A2 => n27406, A3 => n2947, ZN => 
                           n16516);
   U13676 : INV_X2 port map( I => n22352, ZN => n4993);
   U29724 : OAI21_X2 port map( A1 => n24509, A2 => n14213, B => n24799, ZN => 
                           n7396);
   U24157 : OAI21_X2 port map( A1 => n1038, A2 => n32424, B => n1635, ZN => 
                           n15702);
   U28768 : INV_X2 port map( I => n25797, ZN => n25912);
   U4633 : OR3_X1 port map( A1 => n38168, A2 => n35855, A3 => n14375, Z => 
                           n13282);
   U28682 : NAND3_X2 port map( A1 => n34494, A2 => n37279, A3 => n17927, ZN => 
                           n23627);
   U6053 : INV_X2 port map( I => n24257, ZN => n36342);
   U9069 : NOR2_X2 port map( A1 => n30431, A2 => n30714, ZN => n11026);
   U4789 : NOR2_X2 port map( A1 => n20968, A2 => n20967, ZN => n20966);
   U3773 : INV_X2 port map( I => n32601, ZN => n23477);
   U1481 : OAI21_X1 port map( A1 => n18593, A2 => n18592, B => n21431, ZN => 
                           n18591);
   U14791 : NAND2_X1 port map( A1 => n26945, A2 => n34908, ZN => n35613);
   U80 : NAND3_X2 port map( A1 => n481, A2 => n29776, A3 => n34914, ZN => n9063
                           );
   U10253 : NAND3_X2 port map( A1 => n8869, A2 => n8491, A3 => n18865, ZN => 
                           n30815);
   U2098 : NOR3_X2 port map( A1 => n6849, A2 => n20537, A3 => n24469, ZN => 
                           n34366);
   U20236 : OAI21_X1 port map( A1 => n20305, A2 => n28064, B => n21239, ZN => 
                           n35447);
   U2177 : OAI21_X2 port map( A1 => n34996, A2 => n7333, B => n38292, ZN => 
                           n14012);
   U21960 : NAND3_X1 port map( A1 => n37210, A2 => n24387, A3 => n31714, ZN => 
                           n4938);
   U21714 : NOR2_X2 port map( A1 => n32359, A2 => n972, ZN => n6649);
   U14587 : OAI21_X2 port map( A1 => n22843, A2 => n19865, B => n2163, ZN => 
                           n22456);
   U6014 : AOI22_X2 port map( A1 => n28425, A2 => n39724, B1 => n9935, B2 => 
                           n10906, ZN => n30748);
   U7830 : INV_X2 port map( I => n27399, ZN => n1473);
   U3516 : BUF_X2 port map( I => n22802, Z => n272);
   U6318 : INV_X2 port map( I => n12612, ZN => n24116);
   U21797 : NOR2_X1 port map( A1 => n24822, A2 => n13214, ZN => n24823);
   U5709 : NAND2_X1 port map( A1 => n25854, A2 => n36048, ZN => n15919);
   U5016 : NOR2_X2 port map( A1 => n1686, A2 => n3644, ZN => n21421);
   U9890 : NOR2_X2 port map( A1 => n10174, A2 => n13150, ZN => n15624);
   U5467 : INV_X2 port map( I => n7324, ZN => n1197);
   U18205 : NAND2_X2 port map( A1 => n28418, A2 => n9169, ZN => n18378);
   U1466 : NOR2_X2 port map( A1 => n11851, A2 => n543, ZN => n6671);
   U24299 : NAND2_X2 port map( A1 => n17577, A2 => n14196, ZN => n17576);
   U13758 : OAI21_X2 port map( A1 => n2458, A2 => n18408, B => n16511, ZN => 
                           n17577);
   U14811 : NOR2_X2 port map( A1 => n35782, A2 => n24406, ZN => n35781);
   U22230 : INV_X4 port map( I => n6684, ZN => n19869);
   U1921 : NAND2_X1 port map( A1 => n31267, A2 => n36157, ZN => n34438);
   U6240 : INV_X4 port map( I => n16043, ZN => n15276);
   U871 : NOR2_X1 port map( A1 => n14989, A2 => n3402, ZN => n14988);
   U8387 : NAND3_X1 port map( A1 => n3048, A2 => n15123, A3 => n9924, ZN => 
                           n15324);
   U1037 : NAND2_X2 port map( A1 => n24118, A2 => n24372, ZN => n24430);
   U5143 : INV_X4 port map( I => n22709, ZN => n1650);
   U30763 : NAND2_X2 port map( A1 => n31574, A2 => n39389, ZN => n13537);
   U3625 : INV_X2 port map( I => n293, ZN => n21917);
   U15421 : NOR2_X2 port map( A1 => n2439, A2 => n2975, ZN => n2974);
   U7204 : NOR2_X2 port map( A1 => n22287, A2 => n22197, ZN => n22134);
   U8827 : NAND2_X1 port map( A1 => n9046, A2 => n35405, ZN => n9045);
   U2245 : NAND2_X2 port map( A1 => n8964, A2 => n35536, ZN => n8138);
   U2512 : AOI22_X2 port map( A1 => n23215, A2 => n23413, B1 => n23412, B2 => 
                           n6421, ZN => n18381);
   U7610 : NAND3_X1 port map( A1 => n30136, A2 => n34177, A3 => n18588, ZN => 
                           n31258);
   U13474 : NAND3_X2 port map( A1 => n23068, A2 => n3906, A3 => n37984, ZN => 
                           n11366);
   U1192 : OAI22_X2 port map( A1 => n25916, A2 => n34265, B1 => n26034, B2 => 
                           n37300, ZN => n12708);
   U24789 : OAI21_X2 port map( A1 => n22962, A2 => n39303, B => n22816, ZN => 
                           n19528);
   U29311 : NAND2_X2 port map( A1 => n26777, A2 => n32256, ZN => n26778);
   U8390 : NOR2_X2 port map( A1 => n32858, A2 => n5487, ZN => n21208);
   U12561 : OAI22_X2 port map( A1 => n7938, A2 => n31055, B1 => n30345, B2 => 
                           n33864, ZN => n3348);
   U3652 : AOI21_X2 port map( A1 => n13150, A2 => n32377, B => n1626, ZN => 
                           n10613);
   U15442 : INV_X2 port map( I => n23226, ZN => n31332);
   U3132 : OAI21_X2 port map( A1 => n32425, A2 => n6637, B => n6639, ZN => 
                           n6994);
   U6726 : AOI21_X2 port map( A1 => n6638, A2 => n6637, B => n30881, ZN => 
                           n6639);
   U253 : NAND2_X2 port map( A1 => n36814, A2 => n27907, ZN => n12312);
   U2134 : NAND2_X2 port map( A1 => n22150, A2 => n33678, ZN => n16511);
   U17799 : INV_X2 port map( I => n33937, ZN => n18455);
   U4824 : INV_X2 port map( I => n22465, ZN => n30322);
   U6218 : INV_X4 port map( I => n25962, ZN => n25803);
   U2340 : NAND2_X1 port map( A1 => n27374, A2 => n27373, ZN => n27375);
   U23915 : INV_X1 port map( I => n11636, ZN => n1095);
   U2805 : INV_X1 port map( I => n29087, ZN => n6675);
   U8640 : NAND3_X1 port map( A1 => n3333, A2 => n39507, A3 => n13065, ZN => 
                           n3332);
   U2049 : INV_X2 port map( I => n22528, ZN => n22454);
   U23222 : INV_X2 port map( I => n26249, ZN => n36801);
   U17959 : AOI21_X2 port map( A1 => n10857, A2 => n38275, B => n32075, ZN => 
                           n10856);
   U23093 : INV_X1 port map( I => n686, ZN => n35881);
   U10687 : OAI21_X2 port map( A1 => n8717, A2 => n8716, B => n29183, ZN => 
                           n20219);
   U7123 : NAND2_X2 port map( A1 => n22803, A2 => n37883, ZN => n4439);
   U12807 : NOR2_X2 port map( A1 => n24293, A2 => n24295, ZN => n13809);
   U3725 : OAI21_X2 port map( A1 => n25401, A2 => n37926, B => n16234, ZN => 
                           n24937);
   U18040 : INV_X2 port map( I => n22263, ZN => n19471);
   U21490 : NAND2_X1 port map( A1 => n841, A2 => n25495, ZN => n19311);
   U16658 : NAND2_X2 port map( A1 => n38483, A2 => n26970, ZN => n4171);
   U5655 : BUF_X4 port map( I => n37054, Z => n1786);
   U8583 : NOR2_X2 port map( A1 => n37217, A2 => n2186, ZN => n11508);
   U3883 : NOR2_X1 port map( A1 => n27420, A2 => n31287, ZN => n13793);
   U13722 : NAND2_X2 port map( A1 => n10433, A2 => n35019, ZN => n4122);
   U13184 : NOR3_X2 port map( A1 => n5380, A2 => n34014, A3 => n22958, ZN => 
                           n34716);
   U21107 : INV_X2 port map( I => n14383, ZN => n14382);
   U10184 : NAND2_X2 port map( A1 => n22132, A2 => n37217, ZN => n22029);
   U26315 : NAND2_X1 port map( A1 => n16146, A2 => n34720, ZN => n16147);
   U6563 : NAND2_X2 port map( A1 => n14037, A2 => n14038, ZN => n14036);
   U3351 : OAI21_X2 port map( A1 => n29760, A2 => n29764, B => n29762, ZN => 
                           n17540);
   U1232 : INV_X2 port map( I => n25702, ZN => n16072);
   U4185 : NAND2_X2 port map( A1 => n38408, A2 => n1627, ZN => n8146);
   U12242 : NOR2_X1 port map( A1 => n8689, A2 => n25723, ZN => n7239);
   U7052 : NAND2_X2 port map( A1 => n20450, A2 => n1627, ZN => n5839);
   U9237 : BUF_X4 port map( I => n14015, Z => n2761);
   U3942 : OR2_X2 port map( A1 => n14481, A2 => n19963, Z => n25685);
   U26215 : AOI21_X2 port map( A1 => n24472, A2 => n19818, B => n33085, ZN => 
                           n20378);
   U11896 : NAND2_X1 port map( A1 => n18946, A2 => n6606, ZN => n8019);
   U27342 : AOI21_X2 port map( A1 => n20150, A2 => n18743, B => n38079, ZN => 
                           n20149);
   U15367 : NAND2_X2 port map( A1 => n31390, A2 => n31389, ZN => n28435);
   U1287 : NAND2_X2 port map( A1 => n1044, A2 => n38282, ZN => n5658);
   U3646 : NOR2_X2 port map( A1 => n2451, A2 => n33396, ZN => n6313);
   U27520 : AND2_X1 port map( A1 => n14583, A2 => n11227, Z => n36483);
   U3353 : NAND2_X2 port map( A1 => n17105, A2 => n29764, ZN => n28962);
   U5792 : OAI21_X2 port map( A1 => n27319, A2 => n2304, B => n1081, ZN => 
                           n2303);
   U3039 : INV_X4 port map( I => n17105, ZN => n29762);
   U1403 : NOR2_X2 port map( A1 => n22115, A2 => n22114, ZN => n22375);
   U12854 : OAI21_X2 port map( A1 => n32590, A2 => n1312, B => n31081, ZN => 
                           n31080);
   U8286 : NOR2_X1 port map( A1 => n7085, A2 => n7084, ZN => n7083);
   U11571 : AOI21_X2 port map( A1 => n27295, A2 => n39531, B => n35485, ZN => 
                           n27296);
   U10518 : NAND2_X1 port map( A1 => n12321, A2 => n15840, ZN => n12320);
   U2246 : NOR2_X2 port map( A1 => n36430, A2 => n36431, ZN => n36429);
   U30203 : NAND2_X2 port map( A1 => n2127, A2 => n2128, ZN => n36795);
   U2076 : NOR2_X1 port map( A1 => n7504, A2 => n20109, ZN => n20108);
   U3381 : OAI21_X2 port map( A1 => n11095, A2 => n11468, B => n38055, ZN => 
                           n2933);
   U17348 : NAND2_X2 port map( A1 => n33116, A2 => n8272, ZN => n35255);
   U28550 : NAND3_X2 port map( A1 => n23213, A2 => n14561, A3 => n4472, ZN => 
                           n23510);
   U23721 : NAND2_X1 port map( A1 => n35959, A2 => n35958, ZN => n32394);
   U7280 : INV_X1 port map( I => n686, ZN => n1352);
   U6923 : INV_X4 port map( I => n13300, ZN => n19507);
   U6154 : NAND2_X2 port map( A1 => n32740, A2 => n36422, ZN => n30326);
   U7470 : BUF_X4 port map( I => n20453, Z => n1399);
   U16080 : NOR2_X2 port map( A1 => n24333, A2 => n14581, ZN => n31484);
   U333 : NAND2_X2 port map( A1 => n28221, A2 => n18841, ZN => n19852);
   U11741 : NAND2_X2 port map( A1 => n14135, A2 => n33689, ZN => n14134);
   U15969 : NOR2_X1 port map( A1 => n32808, A2 => n18274, ZN => n19907);
   U2346 : NOR2_X2 port map( A1 => n37984, A2 => n23143, ZN => n23156);
   U15653 : NOR2_X2 port map( A1 => n1118, A2 => n38794, ZN => n12407);
   U696 : OAI21_X1 port map( A1 => n35768, A2 => n35767, B => n35766, ZN => 
                           n27052);
   U23016 : NAND2_X1 port map( A1 => n3430, A2 => n19765, ZN => n10209);
   U4293 : INV_X2 port map( I => n14450, ZN => n21498);
   U8128 : NOR2_X2 port map( A1 => n25583, A2 => n1253, ZN => n17815);
   U4935 : OAI22_X1 port map( A1 => n7302, A2 => n7303, B1 => n29464, B2 => 
                           n9105, ZN => n616);
   U11900 : OAI21_X2 port map( A1 => n27226, A2 => n35427, B => n11256, ZN => 
                           n27228);
   U11091 : NAND2_X2 port map( A1 => n28705, A2 => n31088, ZN => n8272);
   U1994 : NOR3_X2 port map( A1 => n18867, A2 => n35442, A3 => n1989, ZN => 
                           n5943);
   U12436 : INV_X2 port map( I => n25625, ZN => n1532);
   U17686 : NAND2_X2 port map( A1 => n15803, A2 => n15802, ZN => n15801);
   U8358 : INV_X2 port map( I => n6402, ZN => n1131);
   U23194 : INV_X2 port map( I => n16039, ZN => n20277);
   U25228 : NAND3_X2 port map( A1 => n8674, A2 => n8673, A3 => n20872, ZN => 
                           n33138);
   U12360 : NAND3_X2 port map( A1 => n24943, A2 => n1112, A3 => n1531, ZN => 
                           n12391);
   U2104 : NAND2_X2 port map( A1 => n15175, A2 => n16635, ZN => n17943);
   U23638 : NAND2_X1 port map( A1 => n16982, A2 => n24214, ZN => n35948);
   U23102 : NAND2_X2 port map( A1 => n7861, A2 => n36262, ZN => n32607);
   U1985 : NAND2_X1 port map( A1 => n18402, A2 => n24383, ZN => n35985);
   U30527 : INV_X2 port map( I => n33895, ZN => n20423);
   U10822 : NAND2_X2 port map( A1 => n15424, A2 => n29776, ZN => n5923);
   U20997 : NAND2_X1 port map( A1 => n18534, A2 => n33726, ZN => n32215);
   U21785 : NAND2_X2 port map( A1 => n28475, A2 => n31088, ZN => n9673);
   U24674 : NOR2_X1 port map( A1 => n4800, A2 => n36188, ZN => n13480);
   U15371 : INV_X2 port map( I => n34987, ZN => n20407);
   U13393 : NOR3_X1 port map( A1 => n18506, A2 => n17578, A3 => n18462, ZN => 
                           n18505);
   U17057 : NAND3_X2 port map( A1 => n26645, A2 => n26751, A3 => n26754, ZN => 
                           n26352);
   U232 : NAND3_X2 port map( A1 => n31347, A2 => n2469, A3 => n1195, ZN => 
                           n6370);
   U816 : INV_X1 port map( I => n25481, ZN => n1534);
   U28387 : NOR2_X2 port map( A1 => n1152, A2 => n22092, ZN => n22091);
   U9110 : INV_X2 port map( I => n10255, ZN => n19750);
   U6598 : OAI21_X2 port map( A1 => n22093, A2 => n22094, B => n35060, ZN => 
                           n22095);
   U10599 : NAND3_X1 port map( A1 => n16126, A2 => n31662, A3 => n31661, ZN => 
                           n34416);
   U3320 : NAND2_X2 port map( A1 => n8131, A2 => n28807, ZN => n2469);
   U8333 : INV_X4 port map( I => n24266, ZN => n1601);
   U13275 : NOR2_X2 port map( A1 => n7939, A2 => n38119, ZN => n7938);
   U29242 : NAND2_X2 port map( A1 => n34892, A2 => n1089, ZN => n26422);
   U2637 : AOI21_X2 port map( A1 => n36912, A2 => n6604, B => n5392, ZN => 
                           n35699);
   U17385 : NAND2_X1 port map( A1 => n15719, A2 => n36649, ZN => n4745);
   U7417 : NAND2_X2 port map( A1 => n11574, A2 => n1177, ZN => n10408);
   U3936 : AND2_X1 port map( A1 => n14450, A2 => n19313, Z => n32410);
   U11545 : NAND2_X1 port map( A1 => n16919, A2 => n1000, ZN => n27024);
   U21539 : INV_X1 port map( I => n32310, ZN => n33450);
   U10216 : NOR2_X1 port map( A1 => n3435, A2 => n1687, ZN => n4902);
   U7858 : INV_X4 port map( I => n27306, ZN => n1086);
   U8078 : NOR2_X1 port map( A1 => n5664, A2 => n33662, ZN => n33908);
   U12076 : INV_X2 port map( I => n26021, ZN => n10474);
   U13773 : NAND2_X2 port map( A1 => n31940, A2 => n35754, ZN => n22212);
   U1427 : AOI22_X2 port map( A1 => n2246, A2 => n36083, B1 => n2247, B2 => 
                           n517, ZN => n35371);
   U605 : INV_X2 port map( I => n26974, ZN => n1497);
   U7329 : INV_X4 port map( I => n1746, ZN => n2840);
   U6912 : BUF_X2 port map( I => n25106, Z => n25448);
   U10096 : NAND2_X1 port map( A1 => n35440, A2 => n4647, ZN => n36053);
   U10003 : NAND2_X2 port map( A1 => n22886, A2 => n20638, ZN => n18365);
   U7896 : AOI21_X2 port map( A1 => n1231, A2 => n35537, B => n8651, ZN => 
                           n12694);
   U12282 : INV_X2 port map( I => n11332, ZN => n11331);
   U329 : NAND2_X2 port map( A1 => n36414, A2 => n36671, ZN => n35478);
   U20217 : NAND2_X1 port map( A1 => n32063, A2 => n32062, ZN => n24624);
   U4288 : NAND2_X2 port map( A1 => n13542, A2 => n935, ZN => n465);
   U29360 : BUF_X4 port map( I => n31132, Z => n36673);
   U130 : INV_X1 port map( I => n19783, ZN => n30232);
   U2751 : BUF_X4 port map( I => n36791, Z => n209);
   U28975 : INV_X2 port map( I => n25469, ZN => n25609);
   U16916 : NOR2_X1 port map( A1 => n5682, A2 => n4677, ZN => n5679);
   U13025 : INV_X4 port map( I => n19990, ZN => n21310);
   U770 : NOR2_X1 port map( A1 => n34660, A2 => n37241, ZN => n35768);
   U2335 : NOR2_X2 port map( A1 => n33737, A2 => n36506, ZN => n35361);
   U954 : AOI22_X2 port map( A1 => n26994, A2 => n1229, B1 => n26996, B2 => 
                           n19364, ZN => n34257);
   U15884 : OAI21_X1 port map( A1 => n7418, A2 => n27180, B => n31459, ZN => 
                           n27004);
   U7415 : AOI21_X2 port map( A1 => n29420, A2 => n505, B => n12262, ZN => 
                           n12261);
   U95 : NOR3_X2 port map( A1 => n505, A2 => n9993, A3 => n29494, ZN => n12262)
                           ;
   U3064 : BUF_X2 port map( I => n18866, Z => n9190);
   U19330 : NOR2_X1 port map( A1 => n18628, A2 => n1073, ZN => n36060);
   U1114 : INV_X2 port map( I => n39055, ZN => n13446);
   U11169 : INV_X2 port map( I => n24661, ZN => n1028);
   U6885 : OAI21_X2 port map( A1 => n16779, A2 => n9922, B => n7949, ZN => 
                           n32250);
   U13344 : NOR2_X2 port map( A1 => n11583, A2 => n4963, ZN => n12254);
   U10343 : NAND2_X2 port map( A1 => n21413, A2 => n19543, ZN => n11433);
   U8037 : BUF_X4 port map( I => n20406, Z => n1755);
   U24051 : NOR2_X2 port map( A1 => n19488, A2 => n1763, ZN => n23091);
   U10593 : INV_X1 port map( I => n12369, ZN => n7302);
   U2979 : OAI21_X2 port map( A1 => n35830, A2 => n12543, B => n34702, ZN => 
                           n18259);
   U8776 : BUF_X4 port map( I => Key(102), Z => n30170);
   U24360 : NAND2_X1 port map( A1 => n372, A2 => n20921, ZN => n32884);
   U5368 : NAND2_X2 port map( A1 => n35330, A2 => n35329, ZN => n139);
   U18416 : NOR2_X2 port map( A1 => n31994, A2 => n34265, ZN => n25981);
   U6379 : NAND3_X1 port map( A1 => n17998, A2 => n1049, A3 => n21117, ZN => 
                           n10744);
   U5974 : BUF_X4 port map( I => n24276, Z => n14378);
   U14792 : INV_X2 port map( I => n26019, ZN => n31310);
   U22277 : AOI21_X2 port map( A1 => n38673, A2 => n10154, B => n22114, ZN => 
                           n11439);
   U5355 : NAND2_X2 port map( A1 => n33855, A2 => n9799, ZN => n34688);
   U3274 : AND2_X2 port map( A1 => n15461, A2 => n7240, Z => n24472);
   U7615 : NAND2_X2 port map( A1 => n28069, A2 => n5020, ZN => n10826);
   U7016 : OAI21_X2 port map( A1 => n24314, A2 => n33077, B => n5572, ZN => 
                           n1877);
   U1115 : INV_X2 port map( I => n16590, ZN => n20791);
   U20266 : NOR2_X1 port map( A1 => n28270, A2 => n1198, ZN => n12497);
   U21317 : NOR2_X1 port map( A1 => n34063, A2 => n35629, ZN => n36853);
   U18431 : INV_X4 port map( I => n5558, ZN => n5935);
   U17458 : INV_X4 port map( I => n11092, ZN => n20924);
   U1095 : INV_X1 port map( I => n18790, ZN => n24372);
   U9707 : NAND3_X2 port map( A1 => n17592, A2 => n24242, A3 => n1593, ZN => 
                           n17591);
   U6770 : NAND2_X1 port map( A1 => n30507, A2 => n16079, ZN => n16078);
   U3112 : OAI21_X2 port map( A1 => n17900, A2 => n30851, B => n30556, ZN => 
                           n16953);
   U9591 : INV_X4 port map( I => n24925, ZN => n1259);
   U20051 : OAI21_X2 port map( A1 => n16841, A2 => n37355, B => n17350, ZN => 
                           n24509);
   U5516 : NOR2_X1 port map( A1 => n7840, A2 => n7839, ZN => n35523);
   U26685 : BUF_X2 port map( I => n10054, Z => n33151);
   U6820 : NOR2_X1 port map( A1 => n4821, A2 => n24395, ZN => n12803);
   U18877 : OAI22_X2 port map( A1 => n36244, A2 => n7978, B1 => n26702, B2 => 
                           n30795, ZN => n26707);
   U2072 : NAND2_X2 port map( A1 => n2192, A2 => n36500, ZN => n4183);
   U22999 : INV_X4 port map( I => n3644, ZN => n22114);
   U4408 : INV_X2 port map( I => n18722, ZN => n21478);
   U1107 : INV_X2 port map( I => n13584, ZN => n10747);
   U23700 : NAND2_X2 port map( A1 => n17294, A2 => n17296, ZN => n32714);
   U25012 : AOI21_X2 port map( A1 => n29481, A2 => n29454, B => n29426, ZN => 
                           n17296);
   U5125 : BUF_X2 port map( I => n8646, Z => n33412);
   U20574 : AOI21_X1 port map( A1 => n3067, A2 => n3066, B => n3065, ZN => 
                           n32132);
   U12665 : NAND2_X2 port map( A1 => n12517, A2 => n37421, ZN => n9826);
   U13734 : NAND2_X1 port map( A1 => n28507, A2 => n34794, ZN => n34781);
   U12873 : NAND2_X1 port map( A1 => n12803, A2 => n24397, ZN => n12802);
   U23107 : OAI21_X2 port map( A1 => n28342, A2 => n28401, B => n28341, ZN => 
                           n11665);
   U4651 : NAND2_X1 port map( A1 => n18384, A2 => n29531, ZN => n17103);
   U13533 : INV_X4 port map( I => n6885, ZN => n17286);
   U9129 : INV_X2 port map( I => n31494, ZN => n1204);
   U3879 : BUF_X4 port map( I => n3213, Z => n362);
   U12858 : OAI21_X2 port map( A1 => n7730, A2 => n19745, B => n13707, ZN => 
                           n13706);
   U6352 : NAND2_X2 port map( A1 => n5907, A2 => n20638, ZN => n20637);
   U5784 : NAND2_X1 port map( A1 => n32266, A2 => n31359, ZN => n35440);
   U28397 : OAI21_X1 port map( A1 => n25469, A2 => n32556, B => n19968, ZN => 
                           n32266);
   U13453 : OAI21_X2 port map( A1 => n22512, A2 => n23213, B => n1312, ZN => 
                           n2253);
   U2102 : OAI21_X2 port map( A1 => n8682, A2 => n8681, B => n24448, ZN => 
                           n11631);
   U13149 : INV_X1 port map( I => n26497, ZN => n34712);
   U2790 : AOI22_X2 port map( A1 => n29482, A2 => n19896, B1 => n29378, B2 => 
                           n31521, ZN => n6734);
   U7994 : INV_X1 port map( I => n27969, ZN => n28233);
   U4692 : NOR2_X2 port map( A1 => n5392, A2 => n37351, ZN => n5451);
   U24613 : OAI21_X2 port map( A1 => n7284, A2 => n1255, B => n1256, ZN => 
                           n16411);
   U7412 : BUF_X2 port map( I => n11083, Z => n34360);
   U4694 : OAI22_X2 port map( A1 => n27207, A2 => n27325, B1 => n27326, B2 => 
                           n1473, ZN => n556);
   U5415 : INV_X4 port map( I => n19499, ZN => n6337);
   U5352 : NAND2_X2 port map( A1 => n30746, A2 => n30745, ZN => n36947);
   U5523 : CLKBUF_X4 port map( I => n28174, Z => n3989);
   U20441 : CLKBUF_X4 port map( I => n24195, Z => n6515);
   U21584 : NAND3_X2 port map( A1 => n24710, A2 => n6491, A3 => n33986, ZN => 
                           n9364);
   U5637 : BUF_X2 port map( I => n13770, Z => n36424);
   U14370 : OR2_X2 port map( A1 => n32986, A2 => n31254, Z => n18575);
   U1 : NAND3_X1 port map( A1 => n32452, A2 => n18795, A3 => n20862, ZN => 
                           n36919);
   U9583 : INV_X2 port map( I => n19572, ZN => n19941);
   U4603 : NOR3_X2 port map( A1 => n11271, A2 => n11081, A3 => n9218, ZN => 
                           n9474);
   U11324 : NAND2_X2 port map( A1 => n8351, A2 => n11407, ZN => n8350);
   U2576 : BUF_X2 port map( I => n28157, Z => n28269);
   U17629 : NAND2_X2 port map( A1 => n13593, A2 => n18187, ZN => n19305);
   U25549 : INV_X1 port map( I => n19631, ZN => n976);
   U7159 : INV_X2 port map( I => n962, ZN => n1313);
   U8105 : AOI22_X2 port map( A1 => n2799, A2 => n954, B1 => n728, B2 => n21254
                           , ZN => n4132);
   U7176 : INV_X2 port map( I => n23162, ZN => n22996);
   U4910 : BUF_X4 port map( I => n17650, Z => n9776);
   U1924 : OAI22_X2 port map( A1 => n15828, A2 => n24433, B1 => n1608, B2 => 
                           n30897, ZN => n15826);
   U29080 : INV_X2 port map( I => n36263, ZN => n36630);
   U9286 : NAND2_X2 port map( A1 => n26996, A2 => n17655, ZN => n20562);
   U2974 : NOR3_X2 port map( A1 => n19412, A2 => n19411, A3 => n29656, ZN => 
                           n18243);
   U1900 : INV_X4 port map( I => n3708, ZN => n23521);
   U7092 : BUF_X2 port map( I => n25798, Z => n34961);
   U612 : INV_X1 port map( I => n875, ZN => n11337);
   U6652 : INV_X2 port map( I => n19823, ZN => n23070);
   U4129 : OAI21_X2 port map( A1 => n13111, A2 => n19364, B => n26692, ZN => 
                           n17826);
   U2241 : NAND2_X2 port map( A1 => n23413, A2 => n5591, ZN => n34635);
   U9127 : BUF_X2 port map( I => n27481, Z => n28123);
   U5330 : BUF_X2 port map( I => n24369, Z => n19942);
   U1175 : INV_X2 port map( I => n25820, ZN => n1511);
   U11215 : NOR2_X1 port map( A1 => n3055, A2 => n3056, ZN => n36709);
   U1053 : INV_X1 port map( I => n24296, ZN => n1598);
   U2034 : NAND2_X2 port map( A1 => n20783, A2 => n1142, ZN => n15272);
   U5245 : NAND2_X1 port map( A1 => n15940, A2 => n17470, ZN => n21128);
   U4974 : INV_X4 port map( I => n22132, ZN => n22030);
   U21390 : INV_X4 port map( I => n11653, ZN => n19544);
   U3088 : BUF_X2 port map( I => n12673, Z => n30995);
   U7265 : BUF_X2 port map( I => n26665, Z => n12290);
   U8761 : CLKBUF_X2 port map( I => Key(139), Z => n19839);
   U20443 : NOR2_X2 port map( A1 => n12705, A2 => n38685, ZN => n12702);
   U29406 : NAND2_X2 port map( A1 => n22302, A2 => n22303, ZN => n22305);
   U7335 : AOI21_X2 port map( A1 => n26980, A2 => n26687, B => n12290, ZN => 
                           n12590);
   U8224 : NOR2_X2 port map( A1 => n2697, A2 => n1996, ZN => n1995);
   U12115 : AOI21_X2 port map( A1 => n13168, A2 => n9605, B => n32109, ZN => 
                           n11764);
   U14296 : OAI21_X2 port map( A1 => n27956, A2 => n16325, B => n34832, ZN => 
                           n11208);
   U1234 : NAND2_X1 port map( A1 => n31432, A2 => n17952, ZN => n35353);
   U13138 : NAND2_X2 port map( A1 => n3383, A2 => n23117, ZN => n3382);
   U16707 : BUF_X2 port map( I => n19467, Z => n28048);
   U25124 : NAND2_X1 port map( A1 => n23271, A2 => n23355, ZN => n18197);
   U2065 : BUF_X4 port map( I => n7536, Z => n123);
   U26094 : NAND2_X1 port map( A1 => n28479, A2 => n1419, ZN => n21190);
   U11778 : AOI21_X1 port map( A1 => n21171, A2 => n26219, B => n16298, ZN => 
                           n5560);
   U11596 : OAI21_X1 port map( A1 => n20709, A2 => n7499, B => n20708, ZN => 
                           n8208);
   U7905 : NOR2_X2 port map( A1 => n21099, A2 => n26970, ZN => n3541);
   U8936 : NAND2_X2 port map( A1 => n1416, A2 => n2022, ZN => n8849);
   U6984 : INV_X4 port map( I => n9276, ZN => n10116);
   U5027 : INV_X2 port map( I => n22711, ZN => n1322);
   U1393 : BUF_X4 port map( I => n25718, Z => n19400);
   U18172 : NOR2_X2 port map( A1 => n38609, A2 => n31697, ZN => n13);
   U6688 : BUF_X4 port map( I => n18229, Z => n12392);
   U7731 : INV_X2 port map( I => n1445, ZN => n1207);
   U25190 : NAND2_X1 port map( A1 => n33109, A2 => n14839, ZN => n12105);
   U17941 : OAI22_X1 port map( A1 => n23309, A2 => n39626, B1 => n23607, B2 => 
                           n23311, ZN => n5592);
   U9789 : AOI22_X2 port map( A1 => n863, A2 => n1093, B1 => n36477, B2 => 
                           n34163, ZN => n34335);
   U4442 : INV_X2 port map( I => n19465, ZN => n10902);
   U2137 : BUF_X4 port map( I => n27249, Z => n7676);
   U28428 : NAND2_X1 port map( A1 => n33370, A2 => n33369, ZN => n7806);
   U17638 : NOR2_X2 port map( A1 => n38914, A2 => n25849, ZN => n2424);
   U4949 : NAND3_X1 port map( A1 => n4750, A2 => n7367, A3 => n21808, ZN => 
                           n7999);
   U12040 : NOR2_X2 port map( A1 => n11858, A2 => n26068, ZN => n2541);
   U25423 : BUF_X2 port map( I => n22674, Z => n18072);
   U8009 : BUF_X2 port map( I => n3158, Z => n3032);
   U2959 : CLKBUF_X4 port map( I => n13545, Z => n611);
   U10467 : CLKBUF_X2 port map( I => Key(80), Z => n29282);
   U4333 : BUF_X2 port map( I => n20591, Z => n20173);
   U8395 : INV_X1 port map( I => n10174, ZN => n1626);
   U12653 : NAND2_X1 port map( A1 => n34646, A2 => n34645, ZN => n25972);
   U13547 : NAND3_X1 port map( A1 => n10146, A2 => n10147, A3 => n971, ZN => 
                           n34763);
   U5793 : INV_X4 port map( I => n7357, ZN => n18429);
   U315 : NAND2_X2 port map( A1 => n7325, A2 => n8056, ZN => n7946);
   U6658 : NOR2_X1 port map( A1 => n10353, A2 => n36090, ZN => n10354);
   U19807 : INV_X4 port map( I => n28560, ZN => n28654);
   U5780 : OAI21_X2 port map( A1 => n22301, A2 => n22075, B => n22076, ZN => 
                           n20356);
   U4449 : NAND2_X1 port map( A1 => n24917, A2 => n18876, ZN => n33209);
   U12201 : NAND2_X1 port map( A1 => n17037, A2 => n39821, ZN => n36693);
   U2539 : NAND3_X1 port map( A1 => n13723, A2 => n13441, A3 => n18997, ZN => 
                           n2555);
   U5363 : NOR2_X1 port map( A1 => n29425, A2 => n20830, ZN => n35296);
   U10323 : OR2_X1 port map( A1 => n34483, A2 => n34597, Z => n34613);
   U1105 : INV_X2 port map( I => n12235, ZN => n24118);
   U14436 : NAND2_X1 port map( A1 => n34855, A2 => n31430, ZN => n18554);
   U312 : AOI21_X1 port map( A1 => n36742, A2 => n35804, B => n32800, ZN => 
                           n6371);
   U10105 : INV_X4 port map( I => n37589, ZN => n23213);
   U6924 : NOR2_X2 port map( A1 => n9703, A2 => n24853, ZN => n14934);
   U22350 : OAI22_X2 port map( A1 => n10116, A2 => n17087, B1 => n9277, B2 => 
                           n32064, ZN => n9703);
   U5629 : NAND2_X1 port map( A1 => n5070, A2 => n33708, ZN => n14201);
   U11229 : NAND3_X1 port map( A1 => n27986, A2 => n38874, A3 => n20053, ZN => 
                           n27987);
   U5496 : AOI21_X2 port map( A1 => n13826, A2 => n11806, B => n1117, ZN => 
                           n32365);
   U18278 : NAND2_X1 port map( A1 => n18346, A2 => n13653, ZN => n9280);
   U4568 : INV_X2 port map( I => n9861, ZN => n31139);
   U13757 : NOR2_X1 port map( A1 => n14777, A2 => n22245, ZN => n20731);
   U3473 : NOR2_X2 port map( A1 => n24698, A2 => n37097, ZN => n1909);
   U11832 : NAND2_X1 port map( A1 => n31238, A2 => n31237, ZN => n31236);
   U5969 : INV_X2 port map( I => n24408, ZN => n24406);
   U30367 : INV_X2 port map( I => n14234, ZN => n23115);
   U12136 : INV_X2 port map( I => n25889, ZN => n7293);
   U12184 : NAND2_X2 port map( A1 => n26079, A2 => n1012, ZN => n18876);
   U30742 : BUF_X4 port map( I => n5831, Z => n36989);
   U21912 : NAND2_X1 port map( A1 => n30393, A2 => n21533, ZN => n16930);
   U7792 : NAND3_X2 port map( A1 => n27072, A2 => n34943, A3 => n39338, ZN => 
                           n5294);
   U23072 : INV_X2 port map( I => n12141, ZN => n14933);
   U1045 : INV_X2 port map( I => n20936, ZN => n35764);
   U3434 : BUF_X4 port map( I => n29897, Z => n30059);
   U27300 : INV_X2 port map( I => n33244, ZN => n33935);
   U5591 : INV_X1 port map( I => n16520, ZN => n27310);
   U4781 : AOI21_X1 port map( A1 => n3637, A2 => n12527, B => n33647, ZN => 
                           n31036);
   U9968 : INV_X2 port map( I => n6355, ZN => n27412);
   U7402 : AOI21_X2 port map( A1 => n29378, A2 => n31521, B => n16877, ZN => 
                           n16876);
   U21016 : INV_X1 port map( I => n23202, ZN => n35576);
   U17427 : INV_X2 port map( I => n13414, ZN => n1036);
   U11732 : NAND2_X1 port map( A1 => n11222, A2 => n11220, ZN => n11225);
   U1424 : INV_X2 port map( I => n20351, ZN => n1329);
   U8178 : NAND2_X2 port map( A1 => n32223, A2 => n32221, ZN => n24365);
   U13405 : NAND2_X2 port map( A1 => n3683, A2 => n22902, ZN => n14331);
   U5278 : BUF_X4 port map( I => n35614, Z => n34014);
   U4671 : OR2_X2 port map( A1 => n24483, A2 => n32360, Z => n30373);
   U24465 : NAND2_X1 port map( A1 => n25708, A2 => n33218, ZN => n18215);
   U1579 : NAND2_X2 port map( A1 => n39258, A2 => n1909, ZN => n3399);
   U7845 : NAND3_X2 port map( A1 => n4583, A2 => n946, A3 => n4582, ZN => n4581
                           );
   U8368 : AOI21_X2 port map( A1 => n20036, A2 => n23559, B => n23560, ZN => 
                           n20035);
   U3546 : NAND2_X2 port map( A1 => n23430, A2 => n34494, ZN => n20036);
   U3524 : NOR2_X2 port map( A1 => n26980, A2 => n26687, ZN => n14830);
   U9322 : INV_X2 port map( I => n26655, ZN => n13645);
   U200 : OAI22_X2 port map( A1 => n9692, A2 => n7063, B1 => n18035, B2 => 
                           n39724, ZN => n14091);
   U21510 : OR2_X2 port map( A1 => n35748, A2 => n25606, Z => n25608);
   U1285 : NAND2_X2 port map( A1 => n7941, A2 => n31523, ZN => n35499);
   U12537 : OAI21_X1 port map( A1 => n2704, A2 => n2703, B => n33195, ZN => 
                           n2701);
   U30108 : BUF_X2 port map( I => n15922, Z => n33603);
   U4782 : INV_X1 port map( I => n12527, ZN => n1430);
   U909 : NAND2_X2 port map( A1 => n34538, A2 => n37585, ZN => n9535);
   U21060 : INV_X4 port map( I => n8526, ZN => n19728);
   U5801 : NOR2_X1 port map( A1 => n9926, A2 => n27187, ZN => n27192);
   U5949 : BUF_X4 port map( I => n28660, Z => n33436);
   U1174 : NAND3_X2 port map( A1 => n8860, A2 => n8858, A3 => n34482, ZN => 
                           n34481);
   U10226 : NOR2_X2 port map( A1 => n34085, A2 => n25435, ZN => n11442);
   U6978 : INV_X4 port map( I => n19507, ZN => n20696);
   U2040 : NOR2_X1 port map( A1 => n8979, A2 => n8978, ZN => n8977);
   U657 : NAND2_X2 port map( A1 => n2518, A2 => n576, ZN => n35218);
   U8287 : OAI21_X1 port map( A1 => n12975, A2 => n24433, B => n10023, ZN => 
                           n13072);
   U7495 : INV_X2 port map( I => n6317, ZN => n5542);
   U3998 : INV_X4 port map( I => n28669, ZN => n14209);
   U10148 : NAND2_X2 port map( A1 => n36008, A2 => n36007, ZN => n25845);
   U12251 : AOI21_X2 port map( A1 => n11268, A2 => n953, B => n11944, ZN => 
                           n16737);
   U1524 : OAI21_X2 port map( A1 => n2288, A2 => n33480, B => n30941, ZN => 
                           n171);
   U26698 : INV_X4 port map( I => n18077, ZN => n25468);
   U9815 : NAND2_X2 port map( A1 => n33804, A2 => n33805, ZN => n34342);
   U26201 : NOR3_X2 port map( A1 => n17346, A2 => n26564, A3 => n17194, ZN => 
                           n15879);
   U10247 : NOR2_X1 port map( A1 => n6822, A2 => n24527, ZN => n15168);
   U21967 : NAND3_X1 port map( A1 => n32485, A2 => n21224, A3 => n36844, ZN => 
                           n32411);
   U27278 : INV_X2 port map( I => n33242, ZN => n728);
   U1056 : OAI21_X1 port map( A1 => n33539, A2 => n1239, B => n7415, ZN => 
                           n20802);
   U26367 : INV_X1 port map( I => n26643, ZN => n36306);
   U1679 : NOR2_X2 port map( A1 => n33532, A2 => n33530, ZN => n33529);
   U12423 : INV_X1 port map( I => n25483, ZN => n6248);
   U11821 : OAI21_X1 port map( A1 => n14427, A2 => n21091, B => n18469, ZN => 
                           n17144);
   U24050 : AOI21_X2 port map( A1 => n23169, A2 => n1763, B => n22810, ZN => 
                           n22811);
   U7008 : OAI21_X1 port map( A1 => n25614, A2 => n25613, B => n25612, ZN => 
                           n25618);
   U11560 : NAND2_X1 port map( A1 => n26622, A2 => n1500, ZN => n34538);
   U6073 : NOR2_X2 port map( A1 => n21236, A2 => n9048, ZN => n9047);
   U24577 : OR2_X2 port map( A1 => n6163, A2 => n7140, Z => n7141);
   U8953 : NAND4_X2 port map( A1 => n29847, A2 => n5108, A3 => n5107, A4 => 
                           n34267, ZN => n34552);
   U1355 : INV_X4 port map( I => n9854, ZN => n23160);
   U2468 : INV_X2 port map( I => n12393, ZN => n34789);
   U14922 : INV_X4 port map( I => n35883, ZN => n34923);
   U4815 : INV_X2 port map( I => n20321, ZN => n26841);
   U13190 : NAND2_X1 port map( A1 => n23249, A2 => n6637, ZN => n11528);
   U2008 : CLKBUF_X2 port map( I => n22993, Z => n32084);
   U10473 : BUF_X2 port map( I => Key(11), Z => n29849);
   U4871 : BUF_X2 port map( I => n34122, Z => n33899);
   U14314 : INV_X2 port map( I => n9266, ZN => n17447);
   U6468 : BUF_X2 port map( I => Key(49), Z => n17428);
   U10482 : BUF_X2 port map( I => Key(21), Z => n19755);
   U14049 : BUF_X2 port map( I => Key(148), Z => n19534);
   U10445 : BUF_X2 port map( I => Key(12), Z => n19722);
   U7313 : BUF_X2 port map( I => Key(126), Z => n19815);
   U14053 : BUF_X2 port map( I => Key(86), Z => n19879);
   U10448 : CLKBUF_X2 port map( I => Key(155), Z => n30122);
   U28501 : INV_X1 port map( I => Key(3), ZN => n29528);
   U8760 : BUF_X2 port map( I => Key(22), Z => n19730);
   U6466 : BUF_X2 port map( I => Key(187), Z => n19761);
   U20774 : INV_X1 port map( I => n29887, ZN => n32174);
   U10437 : CLKBUF_X4 port map( I => n21790, Z => n18205);
   U8863 : INV_X1 port map( I => n28821, ZN => n30682);
   U10411 : INV_X2 port map( I => n8936, ZN => n21833);
   U25516 : INV_X1 port map( I => n19763, ZN => n14820);
   U26977 : INV_X1 port map( I => n29463, ZN => n33184);
   U8722 : INV_X2 port map( I => n34122, ZN => n21923);
   U30573 : CLKBUF_X2 port map( I => n32370, Z => n36887);
   U27790 : INV_X1 port map( I => n30016, ZN => n33311);
   U7296 : CLKBUF_X4 port map( I => n11576, Z => n10120);
   U14006 : CLKBUF_X2 port map( I => n21752, Z => n19416);
   U4969 : BUF_X2 port map( I => n21496, Z => n16128);
   U14007 : INV_X1 port map( I => n29141, ZN => n18700);
   U26650 : CLKBUF_X2 port map( I => n695, Z => n33148);
   U1518 : INV_X2 port map( I => n17209, ZN => n21894);
   U4879 : CLKBUF_X2 port map( I => n12670, Z => n33885);
   U14002 : CLKBUF_X2 port map( I => n21841, Z => n18152);
   U25500 : INV_X1 port map( I => n29337, ZN => n20479);
   U6436 : CLKBUF_X2 port map( I => n20810, Z => n10044);
   U8662 : INV_X2 port map( I => n34247, ZN => n20923);
   U23225 : INV_X2 port map( I => n21761, ZN => n11851);
   U7866 : INV_X2 port map( I => n17799, ZN => n18028);
   U27618 : CLKBUF_X2 port map( I => n21840, Z => n33285);
   U27516 : INV_X1 port map( I => n21789, ZN => n21527);
   U23244 : OR2_X1 port map( A1 => n11900, A2 => n18293, Z => n15274);
   U22005 : NAND2_X1 port map( A1 => n21728, A2 => n36721, ZN => n35723);
   U17056 : NAND2_X1 port map( A1 => n21867, A2 => n15359, ZN => n12333);
   U13825 : AOI21_X1 port map( A1 => n21059, A2 => n21058, B => n7640, ZN => 
                           n21057);
   U20143 : OAI21_X1 port map( A1 => n17866, A2 => n21859, B => n36351, ZN => 
                           n35437);
   U7728 : BUF_X2 port map( I => n8040, Z => n3676);
   U3304 : CLKBUF_X4 port map( I => n22354, Z => n9685);
   U16900 : NAND2_X1 port map( A1 => n4424, A2 => n20679, ZN => n5796);
   U21260 : CLKBUF_X2 port map( I => n22122, Z => n32259);
   U4045 : BUF_X2 port map( I => n2696, Z => n32434);
   U5791 : CLKBUF_X4 port map( I => n11327, Z => n11171);
   U15527 : INV_X2 port map( I => n22292, ZN => n33713);
   U27270 : CLKBUF_X2 port map( I => n8882, Z => n36457);
   U30132 : BUF_X2 port map( I => n19773, Z => n33623);
   U1426 : INV_X2 port map( I => n22281, ZN => n19486);
   U25788 : CLKBUF_X4 port map( I => n19655, Z => n36237);
   U6495 : AOI21_X1 port map( A1 => n1686, A2 => n13191, B => n38375, ZN => 
                           n11234);
   U6021 : INV_X1 port map( I => n22045, ZN => n10924);
   U17744 : INV_X1 port map( I => n12964, ZN => n20773);
   U10144 : NOR2_X1 port map( A1 => n22199, A2 => n8518, ZN => n14270);
   U14112 : CLKBUF_X4 port map( I => n1326, Z => n34808);
   U28422 : NAND2_X1 port map( A1 => n22353, A2 => n21288, ZN => n22208);
   U17545 : NAND2_X1 port map( A1 => n22009, A2 => n22214, ZN => n21105);
   U28413 : OAI21_X1 port map( A1 => n22204, A2 => n19837, B => n22207, ZN => 
                           n22163);
   U2531 : CLKBUF_X4 port map( I => n22334, Z => n36443);
   U24186 : OAI21_X1 port map( A1 => n15294, A2 => n13910, B => n22156, ZN => 
                           n13909);
   U20007 : NAND2_X1 port map( A1 => n12433, A2 => n7093, ZN => n36436);
   U6564 : NOR2_X1 port map( A1 => n8701, A2 => n22172, ZN => n33228);
   U27606 : NAND2_X1 port map( A1 => n22144, A2 => n33438, ZN => n19430);
   U27748 : INV_X1 port map( I => n21298, ZN => n20239);
   U25088 : AOI21_X1 port map( A1 => n21337, A2 => n14024, B => n33359, ZN => 
                           n19216);
   U2208 : NAND2_X1 port map( A1 => n21335, A2 => n21334, ZN => n21338);
   U13690 : NAND2_X1 port map( A1 => n11142, A2 => n1149, ZN => n11141);
   U4162 : INV_X1 port map( I => n34345, ZN => n36778);
   U2938 : CLKBUF_X4 port map( I => n6014, Z => n5284);
   U24425 : INV_X1 port map( I => n16798, ZN => n22174);
   U20955 : NAND2_X1 port map( A1 => n22026, A2 => n22027, ZN => n4630);
   U8053 : BUF_X2 port map( I => n3528, Z => n34188);
   U6266 : CLKBUF_X2 port map( I => n33227, Z => n36362);
   U13602 : BUF_X1 port map( I => n22773, Z => n19848);
   U15263 : NAND2_X1 port map( A1 => n33072, A2 => n33780, ZN => n34972);
   U20866 : CLKBUF_X2 port map( I => n15346, Z => n35559);
   U25494 : INV_X2 port map( I => n22430, ZN => n21215);
   U6258 : INV_X1 port map( I => n7560, ZN => n34691);
   U11465 : CLKBUF_X2 port map( I => n22711, Z => n30950);
   U6239 : CLKBUF_X2 port map( I => n23140, Z => n36763);
   U23928 : CLKBUF_X2 port map( I => n5337, Z => n35994);
   U10088 : CLKBUF_X4 port map( I => n23152, Z => n8569);
   U4008 : CLKBUF_X1 port map( I => n12631, Z => n31183);
   U6231 : CLKBUF_X2 port map( I => n13668, Z => n34419);
   U2006 : BUF_X2 port map( I => n22709, Z => n383);
   U2462 : INV_X2 port map( I => n8539, ZN => n33925);
   U2458 : CLKBUF_X2 port map( I => n407, Z => n32515);
   U6224 : BUF_X2 port map( I => n23164, Z => n36095);
   U6235 : CLKBUF_X4 port map( I => n22946, Z => n34013);
   U13568 : CLKBUF_X4 port map( I => n23102, Z => n18244);
   U8550 : INV_X2 port map( I => n14442, ZN => n1147);
   U1368 : INV_X2 port map( I => n7160, ZN => n16678);
   U6655 : BUF_X2 port map( I => n21291, Z => n11582);
   U4784 : BUF_X2 port map( I => n39811, Z => n33082);
   U6617 : INV_X1 port map( I => n12029, ZN => n35667);
   U23236 : INV_X1 port map( I => n32636, ZN => n23052);
   U1359 : INV_X1 port map( I => n22864, ZN => n22994);
   U13469 : NAND2_X1 port map( A1 => n9255, A2 => n23123, ZN => n3046);
   U6226 : INV_X1 port map( I => n11913, ZN => n35851);
   U2432 : INV_X2 port map( I => n23020, ZN => n23138);
   U14767 : INV_X2 port map( I => n22833, ZN => n1141);
   U10563 : NAND2_X1 port map( A1 => n32084, A2 => n15239, ZN => n15238);
   U1326 : INV_X2 port map( I => n781, ZN => n1045);
   U8481 : NOR2_X1 port map( A1 => n17124, A2 => n35442, ZN => n5810);
   U25339 : NAND2_X1 port map( A1 => n23177, A2 => n23174, ZN => n36185);
   U4031 : OR2_X1 port map( A1 => n23066, A2 => n22994, Z => n14747);
   U27440 : NAND2_X1 port map( A1 => n19013, A2 => n14390, ZN => n22918);
   U5264 : NOR2_X1 port map( A1 => n33763, A2 => n19697, ZN => n36043);
   U2349 : NOR2_X1 port map( A1 => n14879, A2 => n30394, ZN => n35347);
   U19635 : NAND2_X1 port map( A1 => n22997, A2 => n35586, ZN => n9330);
   U6192 : NAND2_X1 port map( A1 => n3811, A2 => n10828, ZN => n36094);
   U19030 : INV_X1 port map( I => n13719, ZN => n23184);
   U19691 : INV_X1 port map( I => n19528, ZN => n7010);
   U6182 : NAND2_X1 port map( A1 => n36043, A2 => n18386, ZN => n35092);
   U23540 : OAI21_X1 port map( A1 => n23020, A2 => n36763, B => n35939, ZN => 
                           n4690);
   U22717 : NAND2_X1 port map( A1 => n22280, A2 => n22833, ZN => n32552);
   U28599 : OAI21_X1 port map( A1 => n23063, A2 => n23062, B => n23061, ZN => 
                           n23064);
   U3226 : OAI21_X1 port map( A1 => n37062, A2 => n22999, B => n23000, ZN => 
                           n8058);
   U3391 : CLKBUF_X4 port map( I => n38704, Z => n5591);
   U13332 : BUF_X2 port map( I => n23464, Z => n5083);
   U13475 : INV_X1 port map( I => n17968, ZN => n23185);
   U5231 : CLKBUF_X4 port map( I => n33453, Z => n31685);
   U2302 : CLKBUF_X2 port map( I => n12028, Z => n35525);
   U7100 : CLKBUF_X4 port map( I => n11669, Z => n6637);
   U14384 : INV_X2 port map( I => n4644, ZN => n35545);
   U9956 : CLKBUF_X2 port map( I => n31908, Z => n34357);
   U14940 : INV_X2 port map( I => n15953, ZN => n23539);
   U23171 : BUF_X4 port map( I => n23631, Z => n32616);
   U2215 : CLKBUF_X4 port map( I => n23251, Z => n23493);
   U7097 : INV_X2 port map( I => n16013, ZN => n16774);
   U4270 : BUF_X2 port map( I => n38614, Z => n36210);
   U13178 : NAND2_X1 port map( A1 => n3174, A2 => n20322, ZN => n3031);
   U13341 : CLKBUF_X2 port map( I => n23530, Z => n18086);
   U28117 : BUF_X2 port map( I => n13038, Z => n33349);
   U18884 : INV_X2 port map( I => n9395, ZN => n23452);
   U23135 : INV_X1 port map( I => n23622, ZN => n23621);
   U20806 : CLKBUF_X4 port map( I => n9395, Z => n33080);
   U9936 : INV_X2 port map( I => n15122, ZN => n17960);
   U13330 : INV_X1 port map( I => n23586, ZN => n13897);
   U6127 : INV_X1 port map( I => n19389, ZN => n35344);
   U9971 : INV_X1 port map( I => n38881, ZN => n1307);
   U13288 : NOR2_X1 port map( A1 => n13897, A2 => n39261, ZN => n7629);
   U7868 : INV_X1 port map( I => n31164, ZN => n23469);
   U1915 : NAND2_X1 port map( A1 => n30789, A2 => n23321, ZN => n30788);
   U1940 : NAND2_X1 port map( A1 => n7387, A2 => n19686, ZN => n23324);
   U3447 : NAND2_X1 port map( A1 => n23216, A2 => n23606, ZN => n18382);
   U13206 : INV_X1 port map( I => n23397, ZN => n20066);
   U24028 : CLKBUF_X4 port map( I => n9968, Z => n36011);
   U13191 : INV_X1 port map( I => n7224, ZN => n11097);
   U2153 : INV_X1 port map( I => n9347, ZN => n35279);
   U27764 : NAND2_X1 port map( A1 => n19923, A2 => n19922, ZN => n23633);
   U13198 : NAND2_X1 port map( A1 => n16863, A2 => n15842, ZN => n7487);
   U16327 : INV_X1 port map( I => n37957, ZN => n2512);
   U25120 : INV_X1 port map( I => n20509, ZN => n24059);
   U5277 : INV_X1 port map( I => n23777, ZN => n12857);
   U2159 : NOR2_X1 port map( A1 => n1616, A2 => n10110, ZN => n10109);
   U13065 : INV_X1 port map( I => n23663, ZN => n7360);
   U13075 : INV_X1 port map( I => n14220, ZN => n23716);
   U1808 : INV_X1 port map( I => n18602, ZN => n24203);
   U2371 : INV_X1 port map( I => n19949, ZN => n20457);
   U3544 : CLKBUF_X2 port map( I => n19949, Z => n277);
   U9823 : CLKBUF_X2 port map( I => n14471, Z => n10152);
   U9819 : CLKBUF_X2 port map( I => n24095, Z => n23694);
   U3822 : BUF_X2 port map( I => n8250, Z => n30311);
   U3316 : CLKBUF_X2 port map( I => n19295, Z => n10073);
   U4702 : CLKBUF_X2 port map( I => n16816, Z => n32069);
   U9808 : INV_X2 port map( I => n23827, ZN => n1276);
   U24838 : NOR2_X1 port map( A1 => n24133, A2 => n19864, ZN => n18277);
   U9820 : BUF_X2 port map( I => n16179, Z => n9066);
   U5302 : INV_X1 port map( I => n24271, ZN => n1124);
   U1763 : INV_X2 port map( I => n9371, ZN => n33513);
   U1797 : CLKBUF_X4 port map( I => n15754, Z => n3869);
   U27662 : CLKBUF_X4 port map( I => n24420, Z => n19584);
   U1132 : CLKBUF_X4 port map( I => n18790, Z => n16081);
   U13745 : BUF_X1 port map( I => n94, Z => n34783);
   U2028 : INV_X2 port map( I => n15385, ZN => n19382);
   U5967 : INV_X1 port map( I => n24370, ZN => n12580);
   U8582 : INV_X2 port map( I => n24381, ZN => n24214);
   U19754 : CLKBUF_X1 port map( I => n24169, Z => n35384);
   U28796 : INV_X1 port map( I => n24412, ZN => n24112);
   U5319 : BUF_X2 port map( I => n24427, Z => n3142);
   U12971 : INV_X2 port map( I => n800, ZN => n18466);
   U9786 : NOR2_X1 port map( A1 => n24168, A2 => n24169, ZN => n4821);
   U14752 : INV_X1 port map( I => n32250, ZN => n3190);
   U1982 : NAND2_X1 port map( A1 => n23845, A2 => n34620, ZN => n17584);
   U22797 : INV_X2 port map( I => n3142, ZN => n32937);
   U28804 : NAND2_X1 port map( A1 => n24137, A2 => n17040, ZN => n24138);
   U12861 : NOR2_X1 port map( A1 => n24398, A2 => n12801, ZN => n12800);
   U25570 : NOR2_X1 port map( A1 => n24081, A2 => n1126, ZN => n24082);
   U12938 : AOI21_X1 port map( A1 => n1034, A2 => n305, B => n4286, ZN => n5014
                           );
   U26853 : BUF_X2 port map( I => n19499, Z => n36376);
   U12602 : NAND2_X1 port map( A1 => n34637, A2 => n4051, ZN => n4050);
   U5337 : NOR2_X1 port map( A1 => n10783, A2 => n31003, ZN => n10777);
   U6932 : INV_X2 port map( I => n24903, ZN => n20155);
   U18783 : INV_X2 port map( I => n24799, ZN => n24655);
   U5074 : CLKBUF_X4 port map( I => n14283, Z => n19);
   U12728 : INV_X2 port map( I => n17087, ZN => n19868);
   U1945 : CLKBUF_X4 port map( I => n9385, Z => n4973);
   U3976 : CLKBUF_X4 port map( I => n32831, Z => n30843);
   U30856 : CLKBUF_X4 port map( I => n7810, Z => n3076);
   U23317 : INV_X2 port map( I => n24668, ZN => n24750);
   U1675 : NOR2_X1 port map( A1 => n24735, A2 => n24814, ZN => n33818);
   U3785 : CLKBUF_X4 port map( I => n12686, Z => n8314);
   U12648 : INV_X1 port map( I => n36955, ZN => n3122);
   U6909 : INV_X2 port map( I => n6357, ZN => n24686);
   U17781 : BUF_X2 port map( I => n24877, Z => n33705);
   U19777 : INV_X1 port map( I => n24566, ZN => n3624);
   U27110 : CLKBUF_X4 port map( I => n24883, Z => n18114);
   U6968 : NAND2_X1 port map( A1 => n14338, A2 => n24762, ZN => n12632);
   U27670 : NAND2_X1 port map( A1 => n24840, A2 => n24843, ZN => n19597);
   U22944 : INV_X2 port map( I => n24250, ZN => n24733);
   U17383 : INV_X1 port map( I => n24763, ZN => n6023);
   U9666 : NAND2_X1 port map( A1 => n31722, A2 => n1582, ZN => n16669);
   U24858 : NAND2_X1 port map( A1 => n4601, A2 => n20926, ZN => n20925);
   U3490 : NAND2_X1 port map( A1 => n15688, A2 => n2018, ZN => n14782);
   U1785 : NAND2_X1 port map( A1 => n17495, A2 => n34947, ZN => n36672);
   U12550 : NAND2_X1 port map( A1 => n10115, A2 => n4688, ZN => n7321);
   U21908 : AOI22_X1 port map( A1 => n32400, A2 => n13901, B1 => n38973, B2 => 
                           n13903, ZN => n12817);
   U26868 : OAI21_X1 port map( A1 => n34115, A2 => n9277, B => n14936, ZN => 
                           n14935);
   U11218 : NOR2_X1 port map( A1 => n1119, A2 => n30915, ZN => n31144);
   U1573 : NAND2_X1 port map( A1 => n13746, A2 => n24832, ZN => n30930);
   U29350 : NAND2_X1 port map( A1 => n25052, A2 => n1273, ZN => n36669);
   U12539 : NAND2_X1 port map( A1 => n18844, A2 => n6336, ZN => n24580);
   U5931 : NAND2_X1 port map( A1 => n2076, A2 => n2075, ZN => n36295);
   U20341 : OAI21_X1 port map( A1 => n15849, A2 => n24648, B => n15848, ZN => 
                           n32087);
   U27669 : NAND2_X1 port map( A1 => n19597, A2 => n24841, ZN => n19596);
   U2216 : NAND2_X1 port map( A1 => n31520, A2 => n31891, ZN => n33043);
   U9600 : CLKBUF_X4 port map( I => n8542, Z => n30761);
   U1709 : INV_X1 port map( I => n25016, ZN => n34653);
   U5853 : INV_X1 port map( I => n39600, ZN => n34856);
   U9596 : CLKBUF_X4 port map( I => n7328, Z => n5208);
   U11907 : CLKBUF_X2 port map( I => n25569, Z => n31004);
   U12482 : CLKBUF_X4 port map( I => n25309, Z => n25469);
   U4547 : CLKBUF_X4 port map( I => n10584, Z => n31780);
   U4527 : BUF_X2 port map( I => n835, Z => n32580);
   U2640 : BUF_X2 port map( I => n25421, Z => n12309);
   U12477 : CLKBUF_X2 port map( I => n25598, Z => n9815);
   U6252 : CLKBUF_X2 port map( I => n5709, Z => n5519);
   U8181 : CLKBUF_X4 port map( I => n13018, Z => n12500);
   U9569 : BUF_X2 port map( I => n25694, Z => n19767);
   U17341 : CLKBUF_X4 port map( I => n25613, Z => n18031);
   U17603 : INV_X1 port map( I => n25158, ZN => n13811);
   U9571 : CLKBUF_X4 port map( I => n25552, Z => n12825);
   U4353 : CLKBUF_X2 port map( I => n16203, Z => n3985);
   U8183 : CLKBUF_X4 port map( I => n25722, Z => n19367);
   U4522 : CLKBUF_X2 port map( I => n252, Z => n32868);
   U1665 : CLKBUF_X2 port map( I => n33948, Z => n19548);
   U3375 : NOR2_X1 port map( A1 => n18545, A2 => n19589, ZN => n14257);
   U5325 : CLKBUF_X2 port map( I => n25355, Z => n25583);
   U30302 : CLKBUF_X2 port map( I => n34576, Z => n36816);
   U9535 : CLKBUF_X4 port map( I => n730, Z => n7986);
   U7460 : NAND2_X1 port map( A1 => n15541, A2 => n1552, ZN => n25349);
   U1676 : NOR2_X1 port map( A1 => n35508, A2 => n36162, ZN => n36142);
   U15988 : AOI21_X1 port map( A1 => n18545, A2 => n19589, B => n25502, ZN => 
                           n15254);
   U23740 : CLKBUF_X4 port map( I => n25696, Z => n32722);
   U26410 : INV_X2 port map( I => n7075, ZN => n33115);
   U5039 : CLKBUF_X1 port map( I => n31010, Z => n35696);
   U10742 : CLKBUF_X2 port map( I => n14805, Z => n34436);
   U15948 : NOR2_X1 port map( A1 => n31619, A2 => n33115, ZN => n7924);
   U5480 : NAND2_X1 port map( A1 => n17815, A2 => n36792, ZN => n4216);
   U819 : NOR2_X1 port map( A1 => n4469, A2 => n1545, ZN => n4465);
   U9448 : NAND2_X1 port map( A1 => n10788, A2 => n1534, ZN => n10787);
   U12333 : NOR2_X1 port map( A1 => n6748, A2 => n25666, ZN => n25667);
   U12320 : NAND2_X1 port map( A1 => n12462, A2 => n12463, ZN => n12996);
   U29082 : AOI22_X1 port map( A1 => n25633, A2 => n25728, B1 => n16168, B2 => 
                           n18294, ZN => n25634);
   U29061 : OAI21_X1 port map( A1 => n1022, A2 => n14413, B => n36019, ZN => 
                           n25515);
   U27461 : NAND2_X1 port map( A1 => n36475, A2 => n36793, ZN => n20626);
   U9467 : OAI21_X1 port map( A1 => n25528, A2 => n517, B => n25333, ZN => 
                           n1992);
   U19228 : NOR2_X1 port map( A1 => n25478, A2 => n8980, ZN => n8979);
   U11749 : INV_X1 port map( I => n34572, ZN => n34571);
   U17665 : NAND2_X1 port map( A1 => n15404, A2 => n14679, ZN => n4888);
   U27104 : NAND2_X1 port map( A1 => n33204, A2 => n30381, ZN => n15445);
   U18322 : AOI21_X1 port map( A1 => n30633, A2 => n32279, B => n19398, ZN => 
                           n32278);
   U12241 : OAI21_X1 port map( A1 => n17868, A2 => n19235, B => n19234, ZN => 
                           n25573);
   U3364 : NAND2_X1 port map( A1 => n11549, A2 => n25621, ZN => n10041);
   U14629 : NAND2_X1 port map( A1 => n4756, A2 => n4754, ZN => n34886);
   U12294 : NAND2_X1 port map( A1 => n6173, A2 => n6172, ZN => n6171);
   U7920 : INV_X2 port map( I => n26106, ZN => n1017);
   U4994 : BUF_X1 port map( I => n37393, Z => n34417);
   U12206 : INV_X2 port map( I => n37393, ZN => n11848);
   U3679 : CLKBUF_X4 port map( I => n26115, Z => n30302);
   U725 : INV_X2 port map( I => n33293, ZN => n1106);
   U4050 : NAND2_X1 port map( A1 => n26093, A2 => n26329, ZN => n15003);
   U2706 : CLKBUF_X4 port map( I => n33909, Z => n31205);
   U16974 : INV_X2 port map( I => n26124, ZN => n5098);
   U18849 : INV_X2 port map( I => n32691, ZN => n26003);
   U4302 : CLKBUF_X4 port map( I => n7901, Z => n3013);
   U7103 : BUF_X2 port map( I => n33644, Z => n31263);
   U6848 : CLKBUF_X4 port map( I => n18032, Z => n16407);
   U4470 : CLKBUF_X4 port map( I => n34609, Z => n30883);
   U775 : INV_X2 port map( I => n37730, ZN => n1524);
   U3090 : CLKBUF_X4 port map( I => n18994, Z => n7767);
   U3259 : INV_X2 port map( I => n17400, ZN => n1011);
   U1923 : CLKBUF_X4 port map( I => n26070, Z => n11858);
   U27612 : AOI21_X1 port map( A1 => n39729, A2 => n33237, B => n35744, ZN => 
                           n19439);
   U12096 : AOI21_X1 port map( A1 => n949, A2 => n18003, B => n18002, ZN => 
                           n11010);
   U26145 : NOR2_X1 port map( A1 => n25459, A2 => n33348, ZN => n18314);
   U12122 : OAI21_X1 port map( A1 => n931, A2 => n7460, B => n13067, ZN => 
                           n13066);
   U1255 : NAND2_X1 port map( A1 => n34647, A2 => n39676, ZN => n34646);
   U29110 : NAND2_X1 port map( A1 => n25959, A2 => n25793, ZN => n25794);
   U23049 : OAI21_X1 port map( A1 => n25957, A2 => n11552, B => n11551, ZN => 
                           n18745);
   U8004 : AOI21_X1 port map( A1 => n12569, A2 => n26012, B => n39661, ZN => 
                           n4401);
   U6826 : INV_X1 port map( I => n26072, ZN => n11859);
   U5698 : NAND2_X1 port map( A1 => n36766, A2 => n26214, ZN => n25833);
   U4355 : NOR2_X1 port map( A1 => n195, A2 => n30436, ZN => n36300);
   U11799 : INV_X1 port map( I => n8858, ZN => n9378);
   U9039 : NAND2_X1 port map( A1 => n25857, A2 => n26072, ZN => n34275);
   U672 : AOI21_X1 port map( A1 => n10889, A2 => n7110, B => n7111, ZN => n9983
                           );
   U3345 : NAND2_X1 port map( A1 => n12105, A2 => n34685, ZN => n10016);
   U7119 : NAND2_X1 port map( A1 => n25651, A2 => n39015, ZN => n3914);
   U1893 : OAI21_X1 port map( A1 => n11859, A2 => n26071, B => n15796, ZN => 
                           n17187);
   U6577 : INV_X1 port map( I => n26565, ZN => n1507);
   U1138 : CLKBUF_X4 port map( I => n14393, Z => n37024);
   U7101 : INV_X1 port map( I => n9174, ZN => n10269);
   U12021 : NAND2_X1 port map( A1 => n34595, A2 => n36293, ZN => n9077);
   U4427 : CLKBUF_X2 port map( I => n18490, Z => n31941);
   U11997 : BUF_X2 port map( I => n26565, Z => n19289);
   U8798 : CLKBUF_X4 port map( I => n2055, Z => n33812);
   U4430 : CLKBUF_X4 port map( I => n14346, Z => n33308);
   U5682 : CLKBUF_X1 port map( I => n17455, Z => n36765);
   U8831 : INV_X2 port map( I => n26234, ZN => n7603);
   U4424 : CLKBUF_X4 port map( I => n26559, Z => n32464);
   U15549 : CLKBUF_X2 port map( I => n20613, Z => n19700);
   U17950 : CLKBUF_X2 port map( I => n3827, Z => n36480);
   U4390 : CLKBUF_X2 port map( I => n36355, Z => n31502);
   U5662 : CLKBUF_X4 port map( I => n26809, Z => n14377);
   U11963 : CLKBUF_X2 port map( I => n26796, Z => n7725);
   U2698 : CLKBUF_X2 port map( I => n14440, Z => n7516);
   U11075 : CLKBUF_X2 port map( I => n14488, Z => n34484);
   U21952 : OR2_X1 port map( A1 => n35197, A2 => n19442, Z => n14659);
   U27962 : CLKBUF_X2 port map( I => n384, Z => n33333);
   U9357 : CLKBUF_X2 port map( I => n14080, Z => n14079);
   U21256 : CLKBUF_X4 port map( I => n8413, Z => n32256);
   U3996 : CLKBUF_X2 port map( I => n26885, Z => n7305);
   U7181 : CLKBUF_X4 port map( I => n14962, Z => n34892);
   U21017 : INV_X2 port map( I => n8479, ZN => n10187);
   U11834 : NAND2_X1 port map( A1 => n18575, A2 => n106, ZN => n20790);
   U15099 : INV_X1 port map( I => n11224, ZN => n11226);
   U3939 : BUF_X2 port map( I => n17252, Z => n33301);
   U11892 : INV_X1 port map( I => n26652, ZN => n26738);
   U27513 : NAND2_X1 port map( A1 => n26798, A2 => n26797, ZN => n19210);
   U11803 : NAND2_X1 port map( A1 => n16049, A2 => n26721, ZN => n27124);
   U530 : INV_X2 port map( I => n26751, ZN => n26898);
   U3933 : NOR2_X1 port map( A1 => n26987, A2 => n26986, ZN => n5480);
   U9315 : NAND2_X1 port map( A1 => n26907, A2 => n26926, ZN => n26912);
   U11524 : NAND2_X1 port map( A1 => n26912, A2 => n9166, ZN => n30958);
   U15275 : OAI21_X1 port map( A1 => n11616, A2 => n26751, B => n26738, ZN => 
                           n34974);
   U12023 : NOR2_X1 port map( A1 => n15594, A2 => n20797, ZN => n9015);
   U19272 : NAND2_X1 port map( A1 => n17514, A2 => n6555, ZN => n6554);
   U16934 : OAI21_X1 port map( A1 => n4459, A2 => n12549, B => n33952, ZN => 
                           n4580);
   U30395 : NOR2_X1 port map( A1 => n26843, A2 => n1002, ZN => n36846);
   U11867 : NAND2_X1 port map( A1 => n26911, A2 => n26910, ZN => n12659);
   U14290 : NAND2_X1 port map( A1 => n16939, A2 => n14659, ZN => n34830);
   U5625 : NAND2_X1 port map( A1 => n31226, A2 => n31225, ZN => n36938);
   U11811 : OR2_X1 port map( A1 => n26898, A2 => n15317, Z => n5172);
   U7328 : NAND2_X1 port map( A1 => n26352, A2 => n34843, ZN => n5590);
   U3050 : OAI21_X1 port map( A1 => n17279, A2 => n17278, B => n1236, ZN => 
                           n15550);
   U25286 : NAND2_X1 port map( A1 => n9619, A2 => n17786, ZN => n36521);
   U523 : NAND2_X1 port map( A1 => n4689, A2 => n9075, ZN => n26733);
   U14128 : INV_X2 port map( I => n1788, ZN => n8137);
   U5627 : INV_X1 port map( I => n26760, ZN => n11517);
   U12726 : NOR2_X1 port map( A1 => n9015, A2 => n9014, ZN => n36501);
   U11789 : INV_X1 port map( I => n14280, ZN => n3136);
   U11747 : CLKBUF_X2 port map( I => n5831, Z => n3513);
   U11774 : NAND2_X1 port map( A1 => n26138, A2 => n11522, ZN => n15685);
   U15140 : CLKBUF_X2 port map( I => n27358, Z => n34952);
   U5767 : CLKBUF_X4 port map( I => n21272, Z => n2760);
   U13593 : CLKBUF_X2 port map( I => n19135, Z => n34769);
   U5888 : CLKBUF_X2 port map( I => n27399, Z => n18228);
   U7361 : CLKBUF_X1 port map( I => n27131, Z => n7620);
   U755 : INV_X2 port map( I => n33662, ZN => n14261);
   U4915 : BUF_X2 port map( I => n9267, Z => n31672);
   U7391 : CLKBUF_X4 port map( I => n9037, Z => n2522);
   U8573 : INV_X2 port map( I => n27288, ZN => n1470);
   U7819 : NAND2_X1 port map( A1 => n19334, A2 => n18195, ZN => n9488);
   U23329 : INV_X2 port map( I => n17166, ZN => n12074);
   U7821 : CLKBUF_X4 port map( I => n27275, Z => n10677);
   U5745 : CLKBUF_X4 port map( I => n27435, Z => n17754);
   U18229 : OAI21_X1 port map( A1 => n18232, A2 => n19619, B => n27271, ZN => 
                           n19329);
   U11644 : AOI21_X1 port map( A1 => n27273, A2 => n20244, B => n38900, ZN => 
                           n20243);
   U406 : NOR2_X1 port map( A1 => n11854, A2 => n11853, ZN => n11855);
   U18566 : NAND2_X1 port map( A1 => n34520, A2 => n33803, ZN => n7403);
   U25327 : NOR2_X1 port map( A1 => n2208, A2 => n32557, ZN => n33376);
   U13598 : NAND2_X1 port map( A1 => n34770, A2 => n27388, ZN => n36036);
   U7414 : NOR2_X1 port map( A1 => n17354, A2 => n7894, ZN => n18861);
   U11582 : NAND2_X1 port map( A1 => n16360, A2 => n27273, ZN => n14057);
   U12138 : CLKBUF_X1 port map( I => n27738, Z => n31020);
   U23651 : INV_X1 port map( I => n27528, ZN => n35986);
   U3906 : CLKBUF_X2 port map( I => n14456, Z => n32783);
   U30258 : INV_X1 port map( I => n27843, ZN => n36809);
   U7704 : CLKBUF_X4 port map( I => n18688, Z => n1454);
   U30386 : CLKBUF_X2 port map( I => n28117, Z => n36844);
   U559 : CLKBUF_X4 port map( I => n20531, Z => n7635);
   U371 : INV_X1 port map( I => n21159, ZN => n19417);
   U7725 : CLKBUF_X2 port map( I => n9775, Z => n7591);
   U5403 : CLKBUF_X4 port map( I => n28093, Z => n28214);
   U17906 : CLKBUF_X2 port map( I => n17533, Z => n32324);
   U3318 : CLKBUF_X4 port map( I => n28125, Z => n10254);
   U7719 : INV_X2 port map( I => n19435, ZN => n1071);
   U7720 : CLKBUF_X4 port map( I => n28186, Z => n15357);
   U2421 : CLKBUF_X2 port map( I => n8148, Z => n288);
   U22708 : CLKBUF_X2 port map( I => n6990, Z => n35827);
   U19801 : CLKBUF_X2 port map( I => n33955, Z => n31966);
   U17964 : OR2_X1 port map( A1 => n20531, A2 => n6640, Z => n14618);
   U4098 : CLKBUF_X4 port map( I => n28188, Z => n9969);
   U4266 : INV_X1 port map( I => n27989, ZN => n33020);
   U4132 : OR3_X1 port map( A1 => n9688, A2 => n17314, A3 => n32352, Z => 
                           n27994);
   U299 : NAND2_X1 port map( A1 => n13714, A2 => n1212, ZN => n13663);
   U22782 : AOI21_X1 port map( A1 => n15597, A2 => n20896, B => n18603, ZN => 
                           n11055);
   U11340 : INV_X1 port map( I => n28108, ZN => n6789);
   U3358 : INV_X2 port map( I => n36838, ZN => n28194);
   U9047 : OAI21_X1 port map( A1 => n35607, A2 => n19280, B => n13251, ZN => 
                           n13250);
   U7670 : OAI21_X1 port map( A1 => n35607, A2 => n1205, B => n11147, ZN => 
                           n6790);
   U5490 : AOI21_X1 port map( A1 => n20993, A2 => n28045, B => n4915, ZN => 
                           n32869);
   U5483 : INV_X1 port map( I => n28420, ZN => n18380);
   U14234 : NAND2_X1 port map( A1 => n13250, A2 => n13249, ZN => n5237);
   U11329 : NAND2_X1 port map( A1 => n19324, A2 => n19325, ZN => n5906);
   U11189 : NAND2_X1 port map( A1 => n35657, A2 => n19946, ZN => n4724);
   U21877 : NAND2_X1 port map( A1 => n27891, A2 => n34447, ZN => n14736);
   U3675 : CLKBUF_X4 port map( I => n28578, Z => n34667);
   U3619 : CLKBUF_X4 port map( I => n9290, Z => n5662);
   U3899 : BUF_X2 port map( I => n28595, Z => n16295);
   U4421 : BUF_X2 port map( I => n1882, Z => n31321);
   U30153 : CLKBUF_X2 port map( I => n20445, Z => n36788);
   U11179 : NAND2_X1 port map( A1 => n12487, A2 => n12486, ZN => n7745);
   U3900 : CLKBUF_X4 port map( I => n6932, Z => n30931);
   U9019 : BUF_X2 port map( I => n9575, Z => n7555);
   U7505 : CLKBUF_X4 port map( I => n28396, Z => n36814);
   U260 : INV_X2 port map( I => n28433, ZN => n28458);
   U29584 : OAI22_X1 port map( A1 => n7454, A2 => n36788, B1 => n28354, B2 => 
                           n28353, ZN => n28355);
   U18088 : NAND2_X1 port map( A1 => n28533, A2 => n8743, ZN => n28504);
   U3999 : CLKBUF_X4 port map( I => n13880, Z => n33843);
   U9757 : INV_X2 port map( I => n8743, ZN => n17800);
   U5477 : INV_X2 port map( I => n28356, ZN => n28611);
   U28689 : CLKBUF_X4 port map( I => n28494, Z => n36609);
   U7526 : INV_X2 port map( I => n17800, ZN => n5890);
   U14818 : NAND2_X1 port map( A1 => n1430, A2 => n28726, ZN => n12610);
   U11167 : CLKBUF_X4 port map( I => n28696, Z => n9648);
   U18299 : NAND2_X1 port map( A1 => n12610, A2 => n32178, ZN => n12607);
   U5420 : NAND2_X1 port map( A1 => n10361, A2 => n36567, ZN => n31404);
   U20539 : NAND2_X1 port map( A1 => n21188, A2 => n21190, ZN => n18103);
   U19562 : NAND2_X1 port map( A1 => n28366, A2 => n37081, ZN => n16343);
   U10992 : NAND2_X1 port map( A1 => n13060, A2 => n17045, ZN => n7647);
   U10947 : OAI21_X1 port map( A1 => n4025, A2 => n28746, B => n4023, ZN => 
                           n28752);
   U3271 : NAND2_X1 port map( A1 => n35030, A2 => n15964, ZN => n4878);
   U19561 : NOR2_X1 port map( A1 => n17322, A2 => n37081, ZN => n17321);
   U229 : NAND2_X1 port map( A1 => n7478, A2 => n34305, ZN => n2900);
   U205 : AOI22_X1 port map( A1 => n9598, A2 => n17320, B1 => n17321, B2 => 
                           n10587, ZN => n17338);
   U16698 : INV_X2 port map( I => n7710, ZN => n29832);
   U6574 : BUF_X2 port map( I => n29249, Z => n18242);
   U4121 : INV_X1 port map( I => n28869, ZN => n31841);
   U6808 : OAI21_X1 port map( A1 => n16656, A2 => n16655, B => n5645, ZN => 
                           n33375);
   U4298 : CLKBUF_X4 port map( I => n18305, Z => n467);
   U17403 : CLKBUF_X2 port map( I => n29903, Z => n18222);
   U8046 : BUF_X2 port map( I => n11415, Z => n482);
   U18373 : CLKBUF_X1 port map( I => n38186, Z => n33404);
   U2781 : CLKBUF_X2 port map( I => n15853, Z => n105);
   U1671 : CLKBUF_X4 port map( I => n28899, Z => n29491);
   U19034 : OAI21_X1 port map( A1 => n30229, A2 => n19765, B => n10590, ZN => 
                           n14281);
   U97 : INV_X2 port map( I => n17238, ZN => n1175);
   U2444 : NAND2_X1 port map( A1 => n8726, A2 => n29286, ZN => n32648);
   U109 : NAND2_X1 port map( A1 => n20405, A2 => n35695, ZN => n35057);
   U4094 : INV_X1 port map( I => n21290, ZN => n32499);
   U7398 : AOI21_X1 port map( A1 => n29629, A2 => n31511, B => n13722, ZN => 
                           n2554);
   U4101 : BUF_X1 port map( I => n30049, Z => n32628);
   U24292 : NOR2_X1 port map( A1 => n30165, A2 => n14184, ZN => n14183);
   U30605 : NAND2_X1 port map( A1 => n36893, A2 => n29389, ZN => n8147);
   U21880 : NAND2_X1 port map( A1 => n29861, A2 => n17779, ZN => n17302);
   U23989 : NAND2_X1 port map( A1 => n32762, A2 => n30001, ZN => n15644);
   U10651 : NAND2_X1 port map( A1 => n29953, A2 => n19196, ZN => n19195);
   U10594 : BUF_X2 port map( I => n29930, Z => n9591);
   U17354 : CLKBUF_X4 port map( I => n19260, Z => n18384);
   U10618 : BUF_X2 port map( I => n29530, Z => n19362);
   U5340 : CLKBUF_X2 port map( I => n30178, Z => n35899);
   U27 : INV_X4 port map( I => n9231, ZN => n30024);
   U29181 : AOI21_X1 port map( A1 => n35175, A2 => n30093, B => n1382, ZN => 
                           n30083);
   U24024 : NAND3_X1 port map( A1 => n9263, A2 => n9264, A3 => n32508, ZN => 
                           n36005);
   U4291 : OR2_X1 port map( A1 => n30180, A2 => n17997, Z => n896);
   U9638 : AOI22_X1 port map( A1 => n29669, A2 => n29668, B1 => n29676, B2 => 
                           n29670, ZN => n34323);
   U4 : NOR2_X1 port map( A1 => n13606, A2 => n29811, ZN => n36365);
   U8792 : CLKBUF_X2 port map( I => Key(112), Z => n19735);
   U6461 : CLKBUF_X2 port map( I => Key(100), Z => n19674);
   U10457 : CLKBUF_X2 port map( I => Key(123), Z => n28821);
   U8754 : CLKBUF_X2 port map( I => Key(114), Z => n19943);
   U8758 : CLKBUF_X2 port map( I => Key(34), Z => n29666);
   U10475 : CLKBUF_X2 port map( I => Key(72), Z => n30104);
   U10483 : CLKBUF_X2 port map( I => Key(115), Z => n19729);
   U8784 : BUF_X2 port map( I => Key(159), Z => n19835);
   U4064 : INV_X1 port map( I => n19786, ZN => n33866);
   U30194 : INV_X1 port map( I => n19943, ZN => n33661);
   U27794 : INV_X1 port map( I => n19883, ZN => n36513);
   U16870 : AOI22_X1 port map( A1 => n21902, A2 => n526, B1 => n35921, B2 => 
                           n7304, ZN => n21904);
   U25073 : NOR2_X1 port map( A1 => n21748, A2 => n21713, ZN => n21649);
   U6313 : CLKBUF_X2 port map( I => n22042, Z => n36428);
   U1444 : INV_X2 port map( I => n22306, ZN => n1335);
   U4848 : BUF_X2 port map( I => n8431, Z => n32817);
   U25402 : OR2_X1 port map( A1 => n22293, A2 => n9265, Z => n14498);
   U29160 : CLKBUF_X2 port map( I => n22348, Z => n36641);
   U2096 : CLKBUF_X4 port map( I => n22549, Z => n7055);
   U1376 : NAND2_X2 port map( A1 => n17339, A2 => n17340, ZN => n22700);
   U21821 : CLKBUF_X4 port map( I => n2126, Z => n36596);
   U4801 : CLKBUF_X2 port map( I => n23214, Z => n32590);
   U23587 : INV_X2 port map( I => n9797, ZN => n23061);
   U6685 : INV_X2 port map( I => n22895, ZN => n20174);
   U8464 : OAI21_X1 port map( A1 => n9770, A2 => n9769, B => n22964, ZN => 
                           n12816);
   U17624 : INV_X2 port map( I => n388, ZN => n1635);
   U2289 : CLKBUF_X4 port map( I => n14235, Z => n35963);
   U6152 : CLKBUF_X2 port map( I => n5357, Z => n35130);
   U6756 : CLKBUF_X4 port map( I => n17508, Z => n15176);
   U27904 : CLKBUF_X1 port map( I => n23337, Z => n36530);
   U1163 : AOI21_X1 port map( A1 => n35664, A2 => n12597, B => n11969, ZN => 
                           n20222);
   U13315 : NOR2_X1 port map( A1 => n16774, A2 => n37431, ZN => n16863);
   U14360 : CLKBUF_X1 port map( I => n3609, Z => n34844);
   U3979 : CLKBUF_X2 port map( I => n18602, Z => n33314);
   U8354 : CLKBUF_X2 port map( I => n8193, Z => n5599);
   U4171 : CLKBUF_X2 port map( I => n14463, Z => n370);
   U17265 : INV_X2 port map( I => n24203, ZN => n7210);
   U4537 : CLKBUF_X1 port map( I => n24202, Z => n18304);
   U5204 : BUF_X2 port map( I => n35134, Z => n35690);
   U9726 : NAND2_X1 port map( A1 => n24294, A2 => n8463, ZN => n9083);
   U2030 : AOI21_X1 port map( A1 => n24214, A2 => n6567, B => n34673, ZN => 
                           n34252);
   U12603 : NOR2_X1 port map( A1 => n4053, A2 => n1031, ZN => n34637);
   U8282 : INV_X1 port map( I => n24737, ZN => n1582);
   U5072 : INV_X2 port map( I => n31986, ZN => n24648);
   U27711 : NAND2_X1 port map( A1 => n39196, A2 => n19565, ZN => n6169);
   U26565 : NAND2_X1 port map( A1 => n24839, A2 => n34906, ZN => n24840);
   U17737 : NAND2_X1 port map( A1 => n6187, A2 => n24806, ZN => n6183);
   U17983 : CLKBUF_X2 port map( I => n31181, Z => n35972);
   U4539 : CLKBUF_X4 port map( I => n15030, Z => n518);
   U4222 : CLKBUF_X4 port map( I => n24924, Z => n449);
   U5866 : CLKBUF_X2 port map( I => n25266, Z => n35953);
   U3920 : BUF_X2 port map( I => n15907, Z => n371);
   U17442 : CLKBUF_X2 port map( I => n20416, Z => n31574);
   U5827 : CLKBUF_X2 port map( I => n20838, Z => n36019);
   U12757 : CLKBUF_X2 port map( I => n25158, Z => n25756);
   U23936 : INV_X1 port map( I => n25727, ZN => n16168);
   U5471 : CLKBUF_X2 port map( I => n17594, Z => n13460);
   U27987 : NAND2_X1 port map( A1 => n15329, A2 => n15172, ZN => n33204);
   U2648 : AOI21_X1 port map( A1 => n32172, A2 => n16677, B => n25449, ZN => 
                           n4620);
   U11751 : AOI21_X1 port map( A1 => n20888, A2 => n19463, B => n25616, ZN => 
                           n34572);
   U9409 : NOR2_X1 port map( A1 => n12768, A2 => n9944, ZN => n34309);
   U12292 : NOR2_X1 port map( A1 => n8123, A2 => n8122, ZN => n8121);
   U754 : INV_X1 port map( I => n9833, ZN => n19121);
   U6868 : BUF_X2 port map( I => n26106, Z => n18162);
   U4489 : BUF_X2 port map( I => n26215, Z => n9868);
   U17021 : INV_X1 port map( I => n15992, ZN => n35155);
   U8039 : INV_X2 port map( I => n14890, ZN => n25928);
   U25607 : BUF_X2 port map( I => n10834, Z => n32979);
   U4475 : BUF_X2 port map( I => n21204, Z => n31340);
   U5540 : BUF_X2 port map( I => n19240, Z => n33474);
   U4977 : CLKBUF_X2 port map( I => n26131, Z => n35109);
   U3950 : BUF_X2 port map( I => n25900, Z => n33327);
   U1342 : NAND2_X1 port map( A1 => n1019, A2 => n35151, ZN => n34647);
   U5442 : OAI21_X1 port map( A1 => n11835, A2 => n11833, B => n19740, ZN => 
                           n12523);
   U11715 : NAND2_X1 port map( A1 => n34573, A2 => n34574, ZN => n34565);
   U21264 : NAND2_X1 port map( A1 => n25110, A2 => n25510, ZN => n18864);
   U1598 : CLKBUF_X2 port map( I => n26968, Z => n13181);
   U10521 : AND2_X1 port map( A1 => n34160, A2 => n26968, Z => n2969);
   U11966 : CLKBUF_X2 port map( I => n20891, Z => n19972);
   U3941 : CLKBUF_X2 port map( I => n866, Z => n31701);
   U7229 : BUF_X2 port map( I => n20704, Z => n9178);
   U11951 : CLKBUF_X2 port map( I => n26630, Z => n26811);
   U4398 : CLKBUF_X2 port map( I => n11224, Z => n33726);
   U2564 : NAND2_X1 port map( A1 => n26860, A2 => n12682, ZN => n11652);
   U21897 : INV_X1 port map( I => n35732, ZN => n30347);
   U20632 : NOR2_X1 port map( A1 => n26812, A2 => n33849, ZN => n12795);
   U2735 : BUF_X2 port map( I => n27436, Z => n30671);
   U11707 : CLKBUF_X2 port map( I => n27252, Z => n9756);
   U5599 : BUF_X2 port map( I => n35051, Z => n34689);
   U760 : CLKBUF_X4 port map( I => n8537, Z => n31875);
   U720 : AND2_X2 port map( A1 => n8798, A2 => n27349, Z => n27351);
   U23578 : CLKBUF_X2 port map( I => n27253, Z => n32697);
   U4342 : CLKBUF_X2 port map( I => n30358, Z => n31683);
   U3610 : INV_X1 port map( I => n27492, ZN => n4885);
   U5401 : BUF_X2 port map( I => n36838, Z => n19657);
   U5474 : CLKBUF_X4 port map( I => n28651, Z => n35830);
   U11115 : CLKBUF_X2 port map( I => n28596, Z => n9598);
   U4852 : CLKBUF_X2 port map( I => n33100, Z => n34915);
   U17300 : CLKBUF_X2 port map( I => n5028, Z => n32595);
   U17206 : BUF_X2 port map( I => n12168, Z => n33647);
   U23047 : NAND2_X1 port map( A1 => n10618, A2 => n32286, ZN => n35875);
   U25962 : BUF_X2 port map( I => n29052, Z => n33041);
   U6102 : CLKBUF_X2 port map( I => n29120, Z => n29286);
   U24059 : BUF_X2 port map( I => n21299, Z => n32777);
   U19231 : NAND2_X1 port map( A1 => n8445, A2 => n6496, ZN => n30001);
   U2847 : BUF_X2 port map( I => n18896, Z => n13705);
   U16847 : CLKBUF_X4 port map( I => n17347, Z => n6252);
   U6505 : INV_X2 port map( I => n13559, ZN => n1382);
   U8839 : INV_X1 port map( I => n3896, ZN => n3897);
   U5675 : BUF_X4 port map( I => n7959, Z => n36244);
   U6382 : BUF_X4 port map( I => n21387, Z => n18417);
   U9503 : NAND2_X1 port map( A1 => n32053, A2 => n7915, ZN => n30808);
   U405 : NAND2_X2 port map( A1 => n30370, A2 => n28118, ZN => n20410);
   U11968 : BUF_X2 port map( I => n26770, Z => n19442);
   U27212 : OAI21_X2 port map( A1 => n19660, A2 => n19659, B => n23070, ZN => 
                           n19360);
   U4311 : NAND2_X1 port map( A1 => n19596, A2 => n19595, ZN => n14826);
   U2885 : OR2_X1 port map( A1 => n37079, A2 => n8604, Z => n27989);
   U27188 : NOR2_X2 port map( A1 => n34923, A2 => n19350, ZN => n36441);
   U5038 : OAI21_X2 port map( A1 => n24685, A2 => n12460, B => n7930, ZN => 
                           n8107);
   U30500 : NAND2_X2 port map( A1 => n33284, A2 => n15876, ZN => n29401);
   U1215 : NOR2_X2 port map( A1 => n30936, A2 => n25467, ZN => n33270);
   U25361 : INV_X4 port map( I => n12049, ZN => n32946);
   U2149 : BUF_X4 port map( I => n23963, Z => n30612);
   U12851 : NOR2_X2 port map( A1 => n24336, A2 => n24332, ZN => n24333);
   U6777 : BUF_X4 port map( I => n855, Z => n12373);
   U5280 : INV_X4 port map( I => n12953, ZN => n1603);
   U6425 : INV_X4 port map( I => n21692, ZN => n1355);
   U8062 : NOR2_X2 port map( A1 => n1018, A2 => n31626, ZN => n1852);
   U3978 : BUF_X2 port map( I => n205, Z => n33379);
   U15539 : BUF_X4 port map( I => n4322, Z => n32974);
   U13480 : NAND2_X1 port map( A1 => n16955, A2 => n16954, ZN => n22945);
   U13923 : NOR2_X2 port map( A1 => n14577, A2 => n21932, ZN => n18025);
   U12758 : NOR2_X2 port map( A1 => n10691, A2 => n10690, ZN => n10689);
   U20527 : NAND3_X2 port map( A1 => n13738, A2 => n13739, A3 => n29286, ZN => 
                           n35502);
   U19520 : OAI21_X2 port map( A1 => n23596, A2 => n36720, B => n23595, ZN => 
                           n14993);
   U4154 : OR2_X1 port map( A1 => n2572, A2 => n18433, Z => n32636);
   U21069 : INV_X4 port map( I => n36214, ZN => n14196);
   U17660 : NAND2_X2 port map( A1 => n4948, A2 => n17465, ZN => n12415);
   U17271 : NOR2_X2 port map( A1 => n7631, A2 => n8757, ZN => n6519);
   U18926 : NAND2_X2 port map( A1 => n9700, A2 => n9698, ZN => n31835);
   U360 : NAND2_X2 port map( A1 => n36478, A2 => n28537, ZN => n4228);
   U7154 : INV_X2 port map( I => n26009, ZN => n26158);
   U4112 : BUF_X2 port map( I => n30154, Z => n33081);
   U14850 : NAND2_X2 port map( A1 => n7941, A2 => n31318, ZN => n31654);
   U3491 : NOR2_X2 port map( A1 => n26140, A2 => n11485, ZN => n11484);
   U18774 : NAND2_X2 port map( A1 => n24770, A2 => n5957, ZN => n24351);
   U12968 : INV_X4 port map( I => n921, ZN => n9508);
   U12925 : NOR2_X1 port map( A1 => n10695, A2 => n1283, ZN => n10694);
   U2140 : INV_X2 port map( I => n8113, ZN => n1993);
   U2951 : INV_X2 port map( I => n29166, ZN => n36928);
   U800 : BUF_X4 port map( I => n39583, Z => n33088);
   U2615 : NAND2_X2 port map( A1 => n19075, A2 => n21778, ZN => n36346);
   U11756 : NOR2_X2 port map( A1 => n16401, A2 => n12177, ZN => n8332);
   U5781 : INV_X2 port map( I => n22075, ZN => n22039);
   U27543 : NAND3_X2 port map( A1 => n1299, A2 => n33538, A3 => n19283, ZN => 
                           n23266);
   U144 : NOR2_X2 port map( A1 => n29286, A2 => n1062, ZN => n11409);
   U11724 : AND2_X2 port map( A1 => n27583, A2 => n27304, Z => n8696);
   U13414 : OAI21_X1 port map( A1 => n23050, A2 => n9854, B => n4566, ZN => 
                           n4565);
   U12781 : NAND2_X2 port map( A1 => n24135, A2 => n24464, ZN => n7033);
   U29924 : NOR2_X2 port map( A1 => n4182, A2 => n33531, ZN => n33530);
   U18667 : BUF_X4 port map( I => n26553, Z => n31791);
   U16476 : OAI21_X2 port map( A1 => n11709, A2 => n11708, B => n11707, ZN => 
                           n17415);
   U22564 : NOR2_X1 port map( A1 => n13547, A2 => n24029, ZN => n35803);
   U2686 : BUF_X4 port map( I => n17220, Z => n36384);
   U3695 : NAND2_X2 port map( A1 => n26802, A2 => n26747, ZN => n4458);
   U19982 : INV_X4 port map( I => n35422, ZN => n15102);
   U14442 : INV_X4 port map( I => n27275, ZN => n4434);
   U16578 : BUF_X4 port map( I => n24104, Z => n24328);
   U2858 : NAND2_X2 port map( A1 => n29483, A2 => n29643, ZN => n29443);
   U14919 : INV_X1 port map( I => n21776, ZN => n34922);
   U22578 : INV_X1 port map( I => n10656, ZN => n21868);
   U2288 : INV_X1 port map( I => n7062, ZN => n2990);
   U5009 : INV_X1 port map( I => n12670, ZN => n21895);
   U22214 : INV_X1 port map( I => n18027, ZN => n14769);
   U3520 : BUF_X2 port map( I => n7304, Z => n275);
   U10419 : INV_X2 port map( I => n19262, ZN => n1350);
   U5816 : NOR2_X1 port map( A1 => n35883, A2 => n21465, ZN => n4084);
   U22693 : INV_X2 port map( I => n13998, ZN => n19483);
   U2199 : INV_X1 port map( I => n21713, ZN => n30731);
   U23516 : INV_X2 port map( I => n15359, ZN => n16305);
   U19590 : INV_X2 port map( I => n35359, ZN => n5392);
   U1538 : INV_X1 port map( I => n13996, ZN => n13959);
   U24311 : INV_X1 port map( I => n14245, ZN => n14373);
   U15320 : INV_X1 port map( I => n31381, ZN => n17242);
   U7304 : INV_X1 port map( I => n20810, ZN => n21492);
   U10426 : INV_X1 port map( I => n694, ZN => n1353);
   U28217 : NAND2_X1 port map( A1 => n19822, A2 => n1372, ZN => n21393);
   U30656 : AOI21_X1 port map( A1 => n17847, A2 => n21839, B => n452, ZN => 
                           n36930);
   U25067 : NOR2_X1 port map( A1 => n21893, A2 => n21568, ZN => n21569);
   U8658 : NAND2_X1 port map( A1 => n19036, A2 => n21702, ZN => n9425);
   U1477 : NOR2_X1 port map( A1 => n19479, A2 => n21775, ZN => n18742);
   U4639 : NOR2_X1 port map( A1 => n21762, A2 => n9642, ZN => n538);
   U13955 : NOR2_X1 port map( A1 => n21894, A2 => n21893, ZN => n21896);
   U8686 : INV_X2 port map( I => n21840, ZN => n15031);
   U6427 : INV_X2 port map( I => n19434, ZN => n21592);
   U10338 : INV_X1 port map( I => n19483, ZN => n6654);
   U4917 : BUF_X2 port map( I => n21517, Z => n587);
   U30029 : NOR2_X1 port map( A1 => n19375, A2 => n8700, ZN => n36751);
   U7855 : INV_X2 port map( I => n21751, ZN => n15910);
   U4933 : NAND2_X1 port map( A1 => n21897, A2 => n17242, ZN => n21838);
   U6413 : NAND2_X1 port map( A1 => n21507, A2 => n9670, ZN => n21591);
   U19081 : NAND2_X1 port map( A1 => n19016, A2 => n21432, ZN => n21825);
   U2655 : NOR2_X1 port map( A1 => n21684, A2 => n19262, ZN => n19403);
   U1525 : INV_X1 port map( I => n9316, ZN => n21724);
   U8690 : NAND2_X1 port map( A1 => n21429, A2 => n14373, ZN => n13805);
   U1520 : INV_X1 port map( I => n21823, ZN => n21861);
   U20008 : NAND2_X1 port map( A1 => n37111, A2 => n32123, ZN => n10345);
   U27635 : INV_X1 port map( I => n21655, ZN => n21779);
   U1495 : INV_X2 port map( I => n10120, ZN => n1159);
   U21870 : NOR2_X1 port map( A1 => n19768, A2 => n21682, ZN => n21812);
   U28187 : INV_X1 port map( I => n21835, ZN => n21837);
   U4918 : INV_X1 port map( I => n21849, ZN => n21667);
   U2814 : NOR2_X1 port map( A1 => n21659, A2 => n21660, ZN => n13257);
   U28206 : OAI21_X1 port map( A1 => n21660, A2 => n21767, B => n21788, ZN => 
                           n21384);
   U19315 : NAND2_X1 port map( A1 => n6604, A2 => n33154, ZN => n21718);
   U6433 : INV_X1 port map( I => n21767, ZN => n21528);
   U18302 : INV_X2 port map( I => n5392, ZN => n21914);
   U5140 : AND2_X1 port map( A1 => n21492, A2 => n21805, Z => n683);
   U17280 : NAND2_X1 port map( A1 => n20266, A2 => n21478, ZN => n14946);
   U24732 : NOR2_X1 port map( A1 => n19434, A2 => n19238, ZN => n20587);
   U13950 : NAND2_X1 port map( A1 => n21787, A2 => n21528, ZN => n4829);
   U3245 : AOI21_X1 port map( A1 => n14783, A2 => n20277, B => n15466, ZN => 
                           n14811);
   U29319 : NAND2_X1 port map( A1 => n6198, A2 => n31604, ZN => n21448);
   U16014 : NAND2_X1 port map( A1 => n2533, A2 => n21751, ZN => n15928);
   U13925 : INV_X1 port map( I => n21850, ZN => n21423);
   U19078 : INV_X1 port map( I => n21825, ZN => n17866);
   U10283 : NAND3_X1 port map( A1 => n15115, A2 => n21727, A3 => n917, ZN => 
                           n14848);
   U17891 : NAND2_X1 port map( A1 => n8441, A2 => n21899, ZN => n8440);
   U8691 : NAND2_X1 port map( A1 => n21817, A2 => n2155, ZN => n2154);
   U28145 : NAND2_X1 port map( A1 => n21327, A2 => n21511, ZN => n21328);
   U13853 : AOI21_X1 port map( A1 => n20762, A2 => n19756, B => n35977, ZN => 
                           n20761);
   U6412 : NAND2_X1 port map( A1 => n19470, A2 => n6241, ZN => n21483);
   U6411 : INV_X1 port map( I => n21924, ZN => n21469);
   U7301 : INV_X1 port map( I => n20923, ZN => n21636);
   U3721 : INV_X2 port map( I => n21339, ZN => n1156);
   U22705 : OAI21_X1 port map( A1 => n10915, A2 => n10918, B => n21804, ZN => 
                           n10914);
   U17011 : NOR3_X1 port map( A1 => n19545, A2 => n21806, A3 => n21410, ZN => 
                           n35153);
   U28971 : INV_X1 port map( I => n1847, ZN => n33413);
   U6037 : AOI21_X1 port map( A1 => n4373, A2 => n19133, B => n16130, ZN => 
                           n16129);
   U10298 : NOR2_X1 port map( A1 => n11378, A2 => n21414, ZN => n21415);
   U26061 : NAND2_X1 port map( A1 => n17966, A2 => n39627, ZN => n15802);
   U4649 : CLKBUF_X2 port map( I => n32617, Z => n543);
   U28312 : NOR2_X1 port map( A1 => n21433, A2 => n18174, ZN => n36578);
   U4662 : NAND2_X1 port map( A1 => n15761, A2 => n13855, ZN => n17763);
   U27980 : NAND2_X1 port map( A1 => n21775, A2 => n19479, ZN => n21612);
   U28302 : NOR2_X1 port map( A1 => n21942, A2 => n21770, ZN => n21637);
   U28746 : NAND2_X1 port map( A1 => n19517, A2 => n21445, ZN => n2759);
   U1475 : INV_X1 port map( I => n21810, ZN => n1346);
   U2193 : NAND2_X1 port map( A1 => n18174, A2 => n36351, ZN => n30874);
   U17279 : NOR2_X1 port map( A1 => n21478, A2 => n19388, ZN => n533);
   U1465 : INV_X1 port map( I => n9616, ZN => n14928);
   U10299 : OAI22_X1 port map( A1 => n5047, A2 => n6234, B1 => n21854, B2 => 
                           n1156, ZN => n21855);
   U10907 : AOI21_X1 port map( A1 => n30874, A2 => n455, B => n33053, ZN => 
                           n21419);
   U2620 : OAI21_X1 port map( A1 => n12927, A2 => n21498, B => n32164, ZN => 
                           n15125);
   U17562 : NAND3_X1 port map( A1 => n35071, A2 => n21789, A3 => n4829, ZN => 
                           n21529);
   U24512 : NAND2_X1 port map( A1 => n21779, A2 => n21656, ZN => n17161);
   U24526 : NAND2_X1 port map( A1 => n39426, A2 => n5132, ZN => n19856);
   U3063 : NAND2_X1 port map( A1 => n21644, A2 => n19647, ZN => n7954);
   U16182 : OAI21_X1 port map( A1 => n37155, A2 => n21515, B => n3670, ZN => 
                           n21516);
   U28165 : NOR2_X1 port map( A1 => n18174, A2 => n19609, ZN => n21342);
   U18894 : NOR2_X1 port map( A1 => n14868, A2 => n19392, ZN => n6102);
   U10326 : AOI21_X1 port map( A1 => n21582, A2 => n19699, B => n21581, ZN => 
                           n21586);
   U10320 : NAND2_X1 port map( A1 => n5505, A2 => n5391, ZN => n5504);
   U10286 : AOI21_X1 port map( A1 => n10127, A2 => n8971, B => n10125, ZN => 
                           n10126);
   U2606 : AOI21_X1 port map( A1 => n21448, A2 => n31292, B => n21672, ZN => 
                           n35737);
   U1486 : NAND2_X1 port map( A1 => n9041, A2 => n21492, ZN => n4296);
   U21448 : NOR2_X1 port map( A1 => n12927, A2 => n35651, ZN => n21797);
   U28277 : AOI21_X1 port map( A1 => n32544, A2 => n21509, B => n33852, ZN => 
                           n21510);
   U10304 : NAND2_X1 port map( A1 => n12852, A2 => n15369, ZN => n2481);
   U5141 : AND2_X1 port map( A1 => n16165, A2 => n1766, Z => n685);
   U16180 : NAND2_X1 port map( A1 => n21583, A2 => n3670, ZN => n21584);
   U3881 : AOI21_X1 port map( A1 => n17112, A2 => n38480, B => n21592, ZN => 
                           n21597);
   U26124 : NOR2_X1 port map( A1 => n21497, A2 => n21656, ZN => n17482);
   U7251 : NOR2_X1 port map( A1 => n21836, A2 => n1158, ZN => n15952);
   U18740 : INV_X2 port map( I => n36425, ZN => n1680);
   U28278 : NAND2_X1 port map( A1 => n21511, A2 => n21510, ZN => n21512);
   U1478 : NOR2_X1 port map( A1 => n4373, A2 => n2645, ZN => n2644);
   U13936 : OAI21_X1 port map( A1 => n21457, A2 => n21456, B => n19337, ZN => 
                           n13789);
   U19124 : INV_X1 port map( I => n6381, ZN => n21501);
   U23732 : NAND2_X1 port map( A1 => n21648, A2 => n21647, ZN => n22008);
   U20711 : INV_X1 port map( I => n10820, ZN => n22221);
   U5806 : INV_X1 port map( I => n22047, ZN => n22108);
   U17771 : NOR2_X1 port map( A1 => n8493, A2 => n22155, ZN => n4935);
   U8603 : INV_X1 port map( I => n31202, ZN => n7046);
   U4647 : INV_X2 port map( I => n22100, ZN => n20391);
   U21068 : NOR2_X1 port map( A1 => n33678, A2 => n14196, ZN => n4765);
   U6540 : NAND2_X1 port map( A1 => n22362, A2 => n36397, ZN => n22358);
   U13754 : INV_X1 port map( I => n2840, ZN => n14038);
   U9374 : INV_X2 port map( I => n5061, ZN => n1149);
   U27208 : INV_X2 port map( I => n14423, ZN => n12230);
   U30354 : INV_X1 port map( I => n38375, ZN => n10930);
   U6292 : BUF_X2 port map( I => n22243, Z => n35429);
   U7219 : NAND2_X1 port map( A1 => n22040, A2 => n2839, ZN => n22181);
   U6020 : INV_X1 port map( I => n16880, ZN => n11091);
   U13816 : INV_X1 port map( I => n22277, ZN => n22313);
   U10205 : NAND2_X1 port map( A1 => n1680, A2 => n16880, ZN => n7578);
   U8628 : INV_X2 port map( I => n19737, ZN => n22229);
   U26324 : INV_X1 port map( I => n22130, ZN => n22189);
   U10270 : INV_X1 port map( I => n17861, ZN => n17897);
   U8631 : INV_X1 port map( I => n22177, ZN => n20943);
   U13736 : NOR2_X1 port map( A1 => n11044, A2 => n196, ZN => n8948);
   U3402 : INV_X2 port map( I => n21864, ZN => n1047);
   U4961 : BUF_X2 port map( I => n8493, Z => n396);
   U4957 : NAND2_X1 port map( A1 => n19471, A2 => n33738, ZN => n22079);
   U26617 : NOR2_X1 port map( A1 => n22358, A2 => n5077, ZN => n36336);
   U7224 : INV_X1 port map( I => n22353, ZN => n1678);
   U6533 : NOR2_X1 port map( A1 => n1328, A2 => n22196, ZN => n20758);
   U15455 : OAI21_X1 port map( A1 => n31407, A2 => n19655, B => n17359, ZN => 
                           n22026);
   U26109 : NAND3_X1 port map( A1 => n8749, A2 => n21864, A3 => n8439, ZN => 
                           n36680);
   U1429 : INV_X1 port map( I => n2257, ZN => n6297);
   U29244 : CLKBUF_X2 port map( I => n21864, Z => n33438);
   U6435 : INV_X2 port map( I => n39075, ZN => n5232);
   U2118 : INV_X1 port map( I => n22296, ZN => n13626);
   U2566 : INV_X1 port map( I => n34379, ZN => n34407);
   U26262 : BUF_X2 port map( I => n474, Z => n33091);
   U3025 : NAND2_X1 port map( A1 => n2840, A2 => n17530, ZN => n17529);
   U8606 : NAND2_X1 port map( A1 => n22267, A2 => n22122, ZN => n17308);
   U8588 : NOR2_X1 port map( A1 => n22190, A2 => n5819, ZN => n21002);
   U22300 : BUF_X2 port map( I => n22306, Z => n32478);
   U3768 : BUF_X2 port map( I => n22332, Z => n30306);
   U16390 : INV_X2 port map( I => n22322, ZN => n11276);
   U18729 : INV_X1 port map( I => n22222, ZN => n22017);
   U1428 : INV_X1 port map( I => n22295, ZN => n22248);
   U5778 : NAND2_X1 port map( A1 => n4388, A2 => n22038, ZN => n3266);
   U5796 : INV_X1 port map( I => n133, ZN => n1684);
   U17680 : NOR2_X1 port map( A1 => n22151, A2 => n35771, ZN => n15175);
   U9113 : INV_X1 port map( I => n22310, ZN => n34282);
   U4443 : INV_X1 port map( I => n22058, ZN => n20234);
   U2619 : NAND2_X1 port map( A1 => n10154, A2 => n10930, ZN => n2127);
   U6530 : NOR2_X1 port map( A1 => n19471, A2 => n33086, ZN => n35014);
   U2549 : INV_X1 port map( I => n22080, ZN => n35514);
   U25635 : NAND2_X1 port map( A1 => n22176, A2 => n20234, ZN => n4746);
   U13707 : NAND2_X1 port map( A1 => n4932, A2 => n17793, ZN => n8348);
   U21476 : NAND2_X1 port map( A1 => n17897, A2 => n20996, ZN => n35652);
   U13710 : NAND2_X1 port map( A1 => n16888, A2 => n22238, ZN => n21826);
   U19515 : NOR2_X1 port map( A1 => n32313, A2 => n35526, ZN => n6807);
   U17507 : OAI21_X1 port map( A1 => n39075, A2 => n6128, B => n1680, ZN => 
                           n14823);
   U19291 : NOR2_X1 port map( A1 => n35618, A2 => n22364, ZN => n22157);
   U4108 : OAI21_X1 port map( A1 => n22313, A2 => n15493, B => n14925, ZN => 
                           n14924);
   U8587 : OAI22_X1 port map( A1 => n1684, A2 => n21972, B1 => n21971, B2 => 
                           n1048, ZN => n17027);
   U16812 : NAND3_X1 port map( A1 => n8520, A2 => n22197, A3 => n22196, ZN => 
                           n22198);
   U10203 : NOR2_X1 port map( A1 => n39075, A2 => n16880, ZN => n18271);
   U8594 : NAND2_X1 port map( A1 => n22323, A2 => n22324, ZN => n1866);
   U15126 : INV_X1 port map( I => n7355, ZN => n14181);
   U26683 : OAI21_X1 port map( A1 => n19253, A2 => n15499, B => n11044, ZN => 
                           n9342);
   U13716 : AOI21_X1 port map( A1 => n7294, A2 => n16936, B => n16935, ZN => 
                           n16934);
   U10245 : NOR2_X1 port map( A1 => n35429, A2 => n1047, ZN => n2434);
   U20719 : NOR2_X1 port map( A1 => n22143, A2 => n8679, ZN => n8029);
   U25089 : NOR2_X1 port map( A1 => n22236, A2 => n33860, ZN => n16227);
   U29791 : NAND3_X1 port map( A1 => n3266, A2 => n22073, A3 => n3269, ZN => 
                           n3265);
   U16722 : NOR2_X1 port map( A1 => n12230, A2 => n4240, ZN => n22172);
   U13133 : NOR2_X1 port map( A1 => n14035, A2 => n14034, ZN => n22043);
   U7203 : NAND2_X1 port map( A1 => n8949, A2 => n22224, ZN => n8745);
   U6589 : INV_X2 port map( I => n36006, ZN => n1344);
   U24769 : NOR2_X1 port map( A1 => n22017, A2 => n32039, ZN => n18803);
   U4775 : NAND2_X1 port map( A1 => n32408, A2 => n22222, ZN => n22015);
   U24264 : NAND2_X1 port map( A1 => n6127, A2 => n1149, ZN => n18928);
   U16829 : NOR2_X1 port map( A1 => n22101, A2 => n22335, ZN => n22103);
   U13811 : NOR2_X1 port map( A1 => n1342, A2 => n20679, ZN => n22173);
   U4032 : INV_X1 port map( I => n22194, ZN => n30996);
   U1419 : INV_X1 port map( I => n20643, ZN => n22225);
   U2509 : NAND2_X1 port map( A1 => n36649, A2 => n36731, ZN => n502);
   U18038 : NOR2_X1 port map( A1 => n22261, A2 => n19471, ZN => n19975);
   U24424 : INV_X1 port map( I => n22059, ZN => n15347);
   U6556 : BUF_X2 port map( I => n22058, Z => n32609);
   U6504 : NAND2_X1 port map( A1 => n1047, A2 => n37089, ZN => n8751);
   U20876 : OAI22_X1 port map( A1 => n22006, A2 => n8275, B1 => n22007, B2 => 
                           n22225, ZN => n21103);
   U5002 : AOI21_X1 port map( A1 => n22065, A2 => n22066, B => n39151, ZN => 
                           n4479);
   U5000 : NOR2_X1 port map( A1 => n22034, A2 => n18854, ZN => n22037);
   U10175 : AOI21_X1 port map( A1 => n11276, A2 => n33091, B => n31092, ZN => 
                           n17537);
   U17071 : OAI21_X1 port map( A1 => n12814, A2 => n36683, B => n22154, ZN => 
                           n12813);
   U16674 : OAI21_X1 port map( A1 => n35755, A2 => n33359, B => n32478, ZN => 
                           n4198);
   U24545 : NOR3_X1 port map( A1 => n22328, A2 => n36303, A3 => n38555, ZN => 
                           n22329);
   U27009 : OAI21_X1 port map( A1 => n11276, A2 => n18253, B => n22324, ZN => 
                           n17782);
   U4406 : NAND2_X1 port map( A1 => n13632, A2 => n22146, ZN => n7911);
   U6381 : NOR2_X1 port map( A1 => n14269, A2 => n22134, ZN => n9391);
   U2083 : OAI21_X1 port map( A1 => n22236, A2 => n19261, B => n33859, ZN => 
                           n20386);
   U10191 : AOI21_X1 port map( A1 => n8751, A2 => n8749, B => n35429, ZN => 
                           n8750);
   U1443 : INV_X1 port map( I => n22254, ZN => n20308);
   U3515 : OAI21_X1 port map( A1 => n8687, A2 => n33438, B => n19430, ZN => 
                           n13614);
   U2081 : OAI21_X1 port map( A1 => n1048, A2 => n32640, B => n20254, ZN => 
                           n33655);
   U25383 : OAI21_X1 port map( A1 => n6724, A2 => n12255, B => n22281, ZN => 
                           n6723);
   U13695 : NAND2_X1 port map( A1 => n15029, A2 => n31649, ZN => n19654);
   U19954 : NOR2_X1 port map( A1 => n584, A2 => n19261, ZN => n15837);
   U8072 : NAND2_X1 port map( A1 => n35754, A2 => n22360, ZN => n34189);
   U28839 : NAND2_X1 port map( A1 => n36616, A2 => n916, ZN => n2883);
   U23468 : NOR2_X1 port map( A1 => n18928, A2 => n22248, ZN => n12325);
   U19836 : OAI21_X1 port map( A1 => n18803, A2 => n18804, B => n35400, ZN => 
                           n19819);
   U1394 : NAND2_X1 port map( A1 => n18429, A2 => n22227, ZN => n22367);
   U5586 : INV_X1 port map( I => n19815, ZN => n31771);
   U30434 : NAND2_X1 port map( A1 => n15852, A2 => n22272, ZN => n22499);
   U30329 : INV_X1 port map( I => n22740, ZN => n33756);
   U26083 : NAND2_X1 port map( A1 => n15837, A2 => n20351, ZN => n15836);
   U10180 : OAI21_X1 port map( A1 => n18999, A2 => n36661, B => n7131, ZN => 
                           n7132);
   U4022 : NAND2_X1 port map( A1 => n17782, A2 => n32803, ZN => n21832);
   U13606 : INV_X1 port map( I => n22651, ZN => n7530);
   U6373 : NOR3_X1 port map( A1 => n3109, A2 => n9485, A3 => n8947, ZN => n3106
                           );
   U8071 : AOI21_X1 port map( A1 => n34189, A2 => n34246, B => n22361, ZN => 
                           n14800);
   U28502 : INV_X1 port map( I => n29528, ZN => n27739);
   U16661 : INV_X1 port map( I => n22648, ZN => n20608);
   U13614 : INV_X1 port map( I => n22542, ZN => n13236);
   U2292 : BUF_X2 port map( I => n3610, Z => n2585);
   U6437 : INV_X1 port map( I => n30085, ZN => n1713);
   U8738 : INV_X1 port map( I => n19407, ZN => n1375);
   U1380 : INV_X1 port map( I => n29325, ZN => n1718);
   U2054 : INV_X2 port map( I => n12195, ZN => n22670);
   U6441 : INV_X1 port map( I => Key(97), ZN => n1697);
   U13639 : INV_X1 port map( I => n17756, ZN => n1664);
   U8557 : INV_X1 port map( I => n22371, ZN => n22732);
   U5823 : INV_X1 port map( I => n19835, ZN => n965);
   U8745 : INV_X1 port map( I => n19940, ZN => n1369);
   U16168 : INV_X1 port map( I => n12818, ZN => n22482);
   U14160 : INV_X1 port map( I => n1805, ZN => n7584);
   U1365 : INV_X1 port map( I => n23074, ZN => n20873);
   U8537 : INV_X1 port map( I => n7584, ZN => n1320);
   U18789 : INV_X2 port map( I => n5976, ZN => n14390);
   U26964 : INV_X2 port map( I => n906, ZN => n23077);
   U26497 : INV_X1 port map( I => n16593, ZN => n23164);
   U2401 : INV_X1 port map( I => n15289, ZN => n19307);
   U26695 : INV_X1 port map( I => n33152, ZN => n14560);
   U30835 : AND2_X1 port map( A1 => n407, A2 => n10162, Z => n22892);
   U3735 : BUF_X4 port map( I => n19680, Z => n6366);
   U27875 : NAND2_X1 port map( A1 => n23188, A2 => n23190, ZN => n20364);
   U5046 : NAND3_X1 port map( A1 => n23078, A2 => n23077, A3 => n33933, ZN => 
                           n23079);
   U24561 : NAND2_X1 port map( A1 => n33925, A2 => n22892, ZN => n20264);
   U25859 : NAND2_X1 port map( A1 => n33817, A2 => n22935, ZN => n17205);
   U2822 : INV_X1 port map( I => n7518, ZN => n12630);
   U4281 : INV_X1 port map( I => n18220, ZN => n7960);
   U13496 : INV_X1 port map( I => n20782, ZN => n13336);
   U6626 : CLKBUF_X2 port map( I => n2047, Z => n35442);
   U10056 : INV_X2 port map( I => n23060, ZN => n14765);
   U23680 : NOR2_X1 port map( A1 => n301, A2 => n12729, ZN => n33544);
   U1305 : NAND2_X1 port map( A1 => n7266, A2 => n14442, ZN => n22979);
   U5997 : INV_X2 port map( I => n10436, ZN => n935);
   U4007 : BUF_X2 port map( I => n22798, Z => n3273);
   U1367 : INV_X2 port map( I => n20267, ZN => n936);
   U6629 : INV_X1 port map( I => n36554, ZN => n34467);
   U5020 : INV_X2 port map( I => n640, ZN => n23013);
   U13328 : INV_X2 port map( I => n33925, ZN => n32740);
   U10061 : INV_X2 port map( I => n3452, ZN => n22919);
   U7167 : INV_X1 port map( I => n22368, ZN => n20439);
   U10094 : INV_X1 port map( I => n20407, ZN => n18071);
   U29917 : CLKBUF_X2 port map( I => n10334, Z => n36736);
   U1323 : INV_X2 port map( I => n23149, ZN => n9699);
   U7171 : INV_X1 port map( I => n23165, ZN => n22975);
   U3183 : INV_X2 port map( I => n22795, ZN => n5380);
   U28543 : INV_X1 port map( I => n23129, ZN => n22958);
   U8554 : INV_X1 port map( I => n12631, ZN => n23095);
   U8497 : INV_X1 port map( I => n39527, ZN => n1318);
   U7175 : INV_X1 port map( I => n550, ZN => n22859);
   U23017 : INV_X1 port map( I => n11481, ZN => n20840);
   U27279 : AND2_X1 port map( A1 => n217, A2 => n32981, Z => n23012);
   U1325 : INV_X1 port map( I => n19697, ZN => n23110);
   U7169 : INV_X1 port map( I => n16174, ZN => n3906);
   U2995 : INV_X2 port map( I => n8245, ZN => n1831);
   U5085 : NOR2_X1 port map( A1 => n32815, A2 => n22915, ZN => n22997);
   U2433 : NOR2_X1 port map( A1 => n23169, A2 => n23167, ZN => n17498);
   U15618 : NOR3_X1 port map( A1 => n9797, A2 => n23058, A3 => n23060, ZN => 
                           n284);
   U16549 : NOR2_X1 port map( A1 => n22804, A2 => n301, ZN => n14880);
   U20148 : NAND2_X1 port map( A1 => n14765, A2 => n23058, ZN => n32040);
   U21147 : OAI21_X1 port map( A1 => n20872, A2 => n23077, B => n23182, ZN => 
                           n8676);
   U10065 : INV_X1 port map( I => n23047, ZN => n8720);
   U6616 : NOR2_X1 port map( A1 => n2350, A2 => n22900, ZN => n15199);
   U27432 : NAND2_X1 port map( A1 => n19082, A2 => n17131, ZN => n20373);
   U3302 : NOR2_X1 port map( A1 => n2771, A2 => n8942, ZN => n10296);
   U16752 : NOR2_X1 port map( A1 => n35684, A2 => n17205, ZN => n35791);
   U16335 : NAND2_X1 port map( A1 => n14130, A2 => n3803, ZN => n15741);
   U13503 : INV_X1 port map( I => n9080, ZN => n11160);
   U6661 : INV_X1 port map( I => n37922, ZN => n22926);
   U13485 : NAND2_X1 port map( A1 => n20590, A2 => n1316, ZN => n15678);
   U13521 : NAND2_X1 port map( A1 => n1315, A2 => n15290, ZN => n5309);
   U28578 : NOR2_X1 port map( A1 => n19697, A2 => n20782, ZN => n22982);
   U13463 : INV_X1 port map( I => n14804, ZN => n15041);
   U1297 : INV_X1 port map( I => n15388, ZN => n5569);
   U27230 : BUF_X2 port map( I => n18415, Z => n36453);
   U7150 : NOR2_X1 port map( A1 => n7960, A2 => n19293, ZN => n18572);
   U2297 : INV_X2 port map( I => n22920, ZN => n18518);
   U7177 : BUF_X2 port map( I => n19167, Z => n19134);
   U16736 : INV_X2 port map( I => n33431, ZN => n22833);
   U1330 : INV_X1 port map( I => n17691, ZN => n23177);
   U7160 : INV_X1 port map( I => n33935, ZN => n19614);
   U29294 : CLKBUF_X2 port map( I => n23101, Z => n36662);
   U10100 : NOR2_X1 port map( A1 => n23095, A2 => n6466, ZN => n22985);
   U5770 : INV_X1 port map( I => n19840, ZN => n19440);
   U7136 : NAND2_X1 port map( A1 => n1313, A2 => n5581, ZN => n8705);
   U18429 : NOR2_X1 port map( A1 => n4713, A2 => n15045, ZN => n5555);
   U10109 : INV_X1 port map( I => n39155, ZN => n1319);
   U2406 : OR2_X1 port map( A1 => n4472, A2 => n2880, Z => n9155);
   U5531 : INV_X1 port map( I => n14395, ZN => n14725);
   U5019 : INV_X1 port map( I => n9472, ZN => n1651);
   U5054 : INV_X1 port map( I => n39811, ZN => n23098);
   U2024 : NAND2_X1 port map( A1 => n33972, A2 => n217, ZN => n5038);
   U10073 : NAND2_X1 port map( A1 => n1652, A2 => n17226, ZN => n10299);
   U13520 : NOR2_X1 port map( A1 => n1316, A2 => n22895, ZN => n16105);
   U21527 : AOI21_X1 port map( A1 => n19134, A2 => n19351, B => n32228, ZN => 
                           n9255);
   U17651 : NAND3_X1 port map( A1 => n23028, A2 => n20077, A3 => n15290, ZN => 
                           n17009);
   U18735 : AOI22_X1 port map( A1 => n17578, A2 => n23211, B1 => n23209, B2 => 
                           n5907, ZN => n18065);
   U14555 : AOI21_X1 port map( A1 => n23020, A2 => n22949, B => n37108, ZN => 
                           n35880);
   U2854 : NAND3_X1 port map( A1 => n5380, A2 => n19621, A3 => n59, ZN => n3628
                           );
   U24269 : AOI22_X1 port map( A1 => n18572, A2 => n22915, B1 => n32815, B2 => 
                           n22870, ZN => n8013);
   U1990 : NAND2_X1 port map( A1 => n35040, A2 => n22880, ZN => n30599);
   U8488 : NOR2_X1 port map( A1 => n1648, A2 => n1316, ZN => n2795);
   U15062 : NAND3_X1 port map( A1 => n6366, A2 => n19614, A3 => n1831, ZN => 
                           n18660);
   U16505 : OAI22_X1 port map( A1 => n36736, A2 => n8730, B1 => n4714, B2 => 
                           n1144, ZN => n22280);
   U3647 : NOR2_X1 port map( A1 => n36453, A2 => n10074, ZN => n5413);
   U2557 : NOR3_X1 port map( A1 => n34014, A2 => n19621, A3 => n34457, ZN => 
                           n11240);
   U7135 : AOI21_X1 port map( A1 => n37589, A2 => n36839, B => n38601, ZN => 
                           n13275);
   U3858 : NAND3_X1 port map( A1 => n1146, A2 => n23053, A3 => n14556, ZN => 
                           n13077);
   U15310 : NOR2_X1 port map( A1 => n34979, A2 => n22985, ZN => n10876);
   U30740 : NOR2_X1 port map( A1 => n2771, A2 => n15911, ZN => n2772);
   U6356 : NOR2_X1 port map( A1 => n15330, A2 => n23098, ZN => n7590);
   U28443 : NOR3_X1 port map( A1 => n13734, A2 => n18244, A3 => n19788, ZN => 
                           n22397);
   U10101 : NAND2_X1 port map( A1 => n23138, A2 => n34368, ZN => n12618);
   U22906 : OAI22_X1 port map( A1 => n18518, A2 => n9725, B1 => n22682, B2 => 
                           n22920, ZN => n11301);
   U13514 : OAI21_X1 port map( A1 => n1824, A2 => n13734, B => n36662, ZN => 
                           n23081);
   U26175 : AOI22_X1 port map( A1 => n33075, A2 => n33074, B1 => n1824, B2 => 
                           n18244, ZN => n3145);
   U2762 : NAND3_X1 port map( A1 => n14396, A2 => n19586, A3 => n33745, ZN => 
                           n31748);
   U15585 : NAND2_X1 port map( A1 => n35016, A2 => n35918, ZN => n4611);
   U13298 : OAI21_X1 port map( A1 => n34727, A2 => n34726, B => n39356, ZN => 
                           n7722);
   U20637 : NAND2_X1 port map( A1 => n6466, A2 => n6366, ZN => n7902);
   U2000 : NOR2_X1 port map( A1 => n1044, A2 => n19469, ZN => n32873);
   U8504 : NOR2_X1 port map( A1 => n13650, A2 => n39811, ZN => n2658);
   U22032 : NAND3_X1 port map( A1 => n23045, A2 => n15330, A3 => n13650, ZN => 
                           n36903);
   U24034 : NAND3_X1 port map( A1 => n18867, A2 => n19181, A3 => n1989, ZN => 
                           n32918);
   U13371 : NAND2_X1 port map( A1 => n15041, A2 => n32270, ZN => n3535);
   U28570 : NOR2_X1 port map( A1 => n22949, A2 => n1046, ZN => n22951);
   U13534 : NOR2_X1 port map( A1 => n19966, A2 => n16104, ZN => n2794);
   U5754 : NAND3_X1 port map( A1 => n20637, A2 => n18072, A3 => n22886, ZN => 
                           n18066);
   U4366 : NOR2_X1 port map( A1 => n5702, A2 => n39350, ZN => n6901);
   U24734 : NOR2_X1 port map( A1 => n6646, A2 => n20077, ZN => n19944);
   U28446 : INV_X1 port map( I => n22838, ZN => n22396);
   U5089 : INV_X1 port map( I => n16967, ZN => n23031);
   U2395 : NOR2_X1 port map( A1 => n23209, A2 => n23135, ZN => n35806);
   U24549 : NOR2_X1 port map( A1 => n15289, A2 => n23028, ZN => n23171);
   U30324 : INV_X2 port map( I => n2553, ZN => n36829);
   U26757 : NAND2_X1 port map( A1 => n19083, A2 => n20373, ZN => n23145);
   U5165 : NAND2_X1 port map( A1 => n22923, A2 => n5838, ZN => n5837);
   U13426 : OAI21_X1 port map( A1 => n13311, A2 => n23028, B => n6646, ZN => 
                           n18330);
   U1276 : OAI22_X1 port map( A1 => n23197, A2 => n31049, B1 => n23199, B2 => 
                           n23198, ZN => n15589);
   U13483 : AOI22_X1 port map( A1 => n17226, A2 => n23142, B1 => n5581, B2 => 
                           n8508, ZN => n8507);
   U8460 : NAND2_X1 port map( A1 => n23012, A2 => n23011, ZN => n6903);
   U6701 : OAI22_X1 port map( A1 => n1045, A2 => n22884, B1 => n20590, B2 => 
                           n4340, ZN => n4704);
   U2356 : AOI22_X1 port map( A1 => n2795, A2 => n22895, B1 => n2794, B2 => 
                           n20173, ZN => n31657);
   U13461 : NAND2_X1 port map( A1 => n23155, A2 => n37674, ZN => n9700);
   U1282 : NOR2_X1 port map( A1 => n23123, A2 => n22876, ZN => n22878);
   U6692 : NAND2_X1 port map( A1 => n5582, A2 => n1652, ZN => n36527);
   U18811 : NAND3_X1 port map( A1 => n8706, A2 => n8705, A3 => n1652, ZN => 
                           n6000);
   U21412 : OAI21_X1 port map( A1 => n35851, A2 => n9322, B => n1141, ZN => 
                           n35644);
   U15119 : OAI21_X1 port map( A1 => n23031, A2 => n22954, B => n18750, ZN => 
                           n6087);
   U16650 : OAI21_X1 port map( A1 => n5413, A2 => n4162, B => n383, ZN => n4161
                           );
   U17375 : NAND2_X1 port map( A1 => n4143, A2 => n9080, ZN => n7639);
   U24441 : INV_X1 port map( I => n22937, ZN => n23096);
   U13524 : INV_X1 port map( I => n23156, ZN => n3561);
   U6349 : NAND2_X1 port map( A1 => n16617, A2 => n7130, ZN => n23432);
   U6348 : OAI21_X1 port map( A1 => n10698, A2 => n23114, B => n1043, ZN => 
                           n10697);
   U1268 : NOR2_X1 port map( A1 => n15740, A2 => n15742, ZN => n6088);
   U7140 : NAND2_X1 port map( A1 => n9339, A2 => n9699, ZN => n9698);
   U13465 : NOR2_X1 port map( A1 => n23187, A2 => n14724, ZN => n4936);
   U5752 : OAI21_X1 port map( A1 => n18072, A2 => n18065, B => n18066, ZN => 
                           n23464);
   U6690 : OR2_X1 port map( A1 => n9155, A2 => n17568, Z => n23511);
   U6336 : INV_X1 port map( I => n17931, ZN => n12093);
   U1237 : INV_X1 port map( I => n35534, ZN => n1306);
   U2508 : CLKBUF_X2 port map( I => n23352, Z => n32158);
   U5247 : BUF_X2 port map( I => n23587, Z => n19686);
   U2293 : BUF_X2 port map( I => n4644, Z => n36859);
   U1264 : NAND2_X1 port map( A1 => n8569, A2 => n23151, ZN => n23158);
   U8435 : INV_X1 port map( I => n23303, ZN => n23488);
   U5744 : INV_X1 port map( I => n7712, ZN => n12083);
   U1955 : INV_X1 port map( I => n23349, ZN => n13305);
   U11695 : INV_X1 port map( I => n17508, ZN => n34558);
   U5169 : INV_X1 port map( I => n23613, ZN => n14739);
   U8475 : INV_X2 port map( I => n23237, ZN => n1140);
   U5261 : INV_X1 port map( I => n31908, ZN => n1290);
   U6722 : INV_X2 port map( I => n35915, ZN => n4207);
   U2332 : NOR2_X1 port map( A1 => n16013, A2 => n23390, ZN => n23622);
   U9901 : NAND2_X1 port map( A1 => n14011, A2 => n23637, ZN => n7009);
   U4255 : INV_X1 port map( I => n7577, ZN => n32425);
   U1239 : INV_X1 port map( I => n23461, ZN => n23370);
   U6732 : INV_X1 port map( I => n35664, ZN => n1632);
   U12178 : INV_X2 port map( I => n4147, ZN => n36130);
   U1914 : NOR2_X1 port map( A1 => n10839, A2 => n35545, ZN => n32401);
   U17322 : INV_X1 port map( I => n22493, ZN => n4542);
   U8330 : INV_X1 port map( I => n18682, ZN => n1297);
   U8407 : INV_X1 port map( I => n23535, ZN => n23537);
   U9963 : INV_X2 port map( I => n36539, ZN => n1300);
   U1954 : INV_X1 port map( I => n10480, ZN => n52);
   U13218 : INV_X2 port map( I => n7379, ZN => n23645);
   U6727 : NAND2_X1 port map( A1 => n23325, A2 => n35534, ZN => n23586);
   U2602 : NOR2_X1 port map( A1 => n23639, A2 => n7712, ZN => n10633);
   U3361 : NAND2_X1 port map( A1 => n34506, A2 => n23548, ZN => n13752);
   U9954 : INV_X1 port map( I => n18425, ZN => n1295);
   U8453 : INV_X2 port map( I => n12028, ZN => n1310);
   U5022 : INV_X1 port map( I => n23532, ZN => n1625);
   U1242 : INV_X1 port map( I => n23473, ZN => n1139);
   U7197 : INV_X2 port map( I => n8668, ZN => n33496);
   U4922 : INV_X2 port map( I => n36810, ZN => n23401);
   U18705 : INV_X1 port map( I => n23478, ZN => n23483);
   U2319 : INV_X1 port map( I => n6159, ZN => n35367);
   U7835 : AND2_X1 port map( A1 => n23423, A2 => n17094, Z => n34121);
   U19428 : AND2_X1 port map( A1 => n39194, A2 => n7225, Z => n20031);
   U17353 : INV_X1 port map( I => n33840, ZN => n960);
   U25144 : OAI22_X1 port map( A1 => n23483, A2 => n9078, B1 => n23361, B2 => 
                           n6176, ZN => n23363);
   U25639 : NAND2_X1 port map( A1 => n23526, A2 => n23404, ZN => n36219);
   U10227 : INV_X2 port map( I => n36564, ZN => n23270);
   U13169 : INV_X1 port map( I => n23227, ZN => n23277);
   U8433 : NOR2_X1 port map( A1 => n23325, A2 => n19481, ZN => n23264);
   U9896 : NOR2_X1 port map( A1 => n23306, A2 => n23483, ZN => n8784);
   U28637 : NOR2_X1 port map( A1 => n18284, A2 => n35808, ZN => n23298);
   U13299 : NAND2_X1 port map( A1 => n23347, A2 => n14845, ZN => n5253);
   U8619 : NAND2_X1 port map( A1 => n7335, A2 => n3496, ZN => n23343);
   U6771 : AOI22_X1 port map( A1 => n7598, A2 => n4600, B1 => n32226, B2 => 
                           n23425, ZN => n18370);
   U20764 : NAND2_X1 port map( A1 => n23302, A2 => n37774, ZN => n32407);
   U13273 : NAND2_X1 port map( A1 => n23533, A2 => n23534, ZN => n16369);
   U7078 : NAND2_X1 port map( A1 => n15642, A2 => n35377, ZN => n2632);
   U6345 : CLKBUF_X2 port map( I => n23461, Z => n18090);
   U24169 : NAND2_X1 port map( A1 => n5591, A2 => n32246, ZN => n23010);
   U21138 : NOR2_X1 port map( A1 => n23453, A2 => n605, ZN => n9588);
   U1210 : INV_X1 port map( I => n23358, ZN => n8965);
   U15352 : NOR2_X1 port map( A1 => n23306, A2 => n8692, ZN => n34981);
   U6138 : NAND2_X1 port map( A1 => n36027, A2 => n36026, ZN => n23275);
   U6728 : NOR2_X1 port map( A1 => n32425, A2 => n6638, ZN => n22989);
   U18763 : NAND2_X1 port map( A1 => n1644, A2 => n37923, ZN => n23286);
   U13266 : INV_X1 port map( I => n23534, ZN => n16086);
   U13246 : INV_X1 port map( I => n23620, ZN => n13603);
   U9879 : NAND2_X1 port map( A1 => n8239, A2 => n10763, ZN => n10207);
   U18870 : BUF_X2 port map( I => n23567, Z => n31829);
   U2316 : NOR2_X1 port map( A1 => n23251, A2 => n5357, ZN => n36888);
   U4740 : INV_X1 port map( I => n23572, ZN => n33721);
   U5237 : INV_X2 port map( I => n2798, ZN => n31661);
   U15472 : NOR2_X1 port map( A1 => n31787, A2 => n35313, ZN => n35312);
   U7091 : INV_X2 port map( I => n23577, ZN => n1134);
   U2290 : BUF_X2 port map( I => n36442, Z => n9835);
   U11244 : INV_X1 port map( I => n23441, ZN => n11095);
   U1209 : INV_X2 port map( I => n23531, ZN => n18236);
   U24170 : NOR2_X1 port map( A1 => n1631, A2 => n5591, ZN => n23215);
   U9869 : NAND2_X1 port map( A1 => n36564, A2 => n23350, ZN => n30974);
   U5180 : NAND2_X1 port map( A1 => n23572, A2 => n1134, ZN => n33719);
   U8369 : AOI21_X1 port map( A1 => n35039, A2 => n39812, B => n4396, ZN => 
                           n4251);
   U6763 : AOI21_X1 port map( A1 => n23444, A2 => n4207, B => n36859, ZN => 
                           n23447);
   U8372 : NAND3_X1 port map( A1 => n23599, A2 => n23489, A3 => n12597, ZN => 
                           n7825);
   U30624 : AOI22_X1 port map( A1 => n8680, A2 => n36885, B1 => n18391, B2 => 
                           n33287, ZN => n36945);
   U13193 : OAI21_X1 port map( A1 => n22989, A2 => n23256, B => n1293, ZN => 
                           n17441);
   U22903 : NAND3_X1 port map( A1 => n23553, A2 => n14623, A3 => n18236, ZN => 
                           n35864);
   U9855 : NOR2_X1 port map( A1 => n23397, A2 => n23264, ZN => n7630);
   U5255 : NOR3_X1 port map( A1 => n30440, A2 => n35001, A3 => n18763, ZN => 
                           n7042);
   U2258 : INV_X1 port map( I => n23526, ZN => n36878);
   U28271 : OAI21_X1 port map( A1 => n2853, A2 => n6637, B => n6638, ZN => 
                           n36577);
   U24384 : OAI21_X1 port map( A1 => n23493, A2 => n23315, B => n19358, ZN => 
                           n23418);
   U20402 : NOR2_X1 port map( A1 => n9192, A2 => n7426, ZN => n35477);
   U5217 : INV_X1 port map( I => n23476, ZN => n12009);
   U15286 : OAI21_X1 port map( A1 => n20991, A2 => n20992, B => n16182, ZN => 
                           n31376);
   U1228 : INV_X1 port map( I => n23400, ZN => n19146);
   U1193 : OAI21_X1 port map( A1 => n16086, A2 => n23533, B => n5184, ZN => 
                           n5183);
   U19184 : NAND2_X1 port map( A1 => n39012, A2 => n6217, ZN => n18237);
   U1835 : AOI21_X1 port map( A1 => n23286, A2 => n31091, B => n33080, ZN => 
                           n31037);
   U19736 : OAI21_X1 port map( A1 => n31949, A2 => n16456, B => n36564, ZN => 
                           n15604);
   U25123 : INV_X1 port map( I => n23581, ZN => n21297);
   U6764 : NAND2_X1 port map( A1 => n23275, A2 => n23274, ZN => n9889);
   U2665 : NAND2_X1 port map( A1 => n5371, A2 => n16370, ZN => n31074);
   U25848 : NAND2_X1 port map( A1 => n12642, A2 => n12641, ZN => n36241);
   U9918 : INV_X1 port map( I => n23560, ZN => n17927);
   U15823 : NAND2_X1 port map( A1 => n23525, A2 => n3365, ZN => n3364);
   U13234 : NAND2_X1 port map( A1 => n12638, A2 => n1304, ZN => n23262);
   U5021 : NAND2_X1 port map( A1 => n31829, A2 => n32260, ZN => n4417);
   U1179 : INV_X1 port map( I => n23554, ZN => n6286);
   U2151 : INV_X1 port map( I => n24012, ZN => n23659);
   U25150 : OAI21_X1 port map( A1 => n18762, A2 => n39133, B => n18763, ZN => 
                           n16056);
   U8377 : OAI22_X1 port map( A1 => n23365, A2 => n3715, B1 => n32260, B2 => 
                           n2921, ZN => n2920);
   U25152 : AOI21_X1 port map( A1 => n23278, A2 => n31332, B => n23277, ZN => 
                           n15562);
   U28591 : NAND2_X1 port map( A1 => n39214, A2 => n30524, ZN => n23038);
   U13215 : NAND3_X1 port map( A1 => n18237, A2 => n18235, A3 => n18086, ZN => 
                           n23224);
   U3861 : NAND2_X1 port map( A1 => n37279, A2 => n23560, ZN => n8238);
   U26540 : OAI21_X1 port map( A1 => n37923, A2 => n23452, B => n16713, ZN => 
                           n16712);
   U28594 : NAND3_X1 port map( A1 => n23040, A2 => n34386, A3 => n18090, ZN => 
                           n23041);
   U13095 : NAND2_X1 port map( A1 => n30364, A2 => n5999, ZN => n7149);
   U2255 : NAND2_X1 port map( A1 => n37005, A2 => n23458, ZN => n23239);
   U26162 : AOI22_X1 port map( A1 => n23640, A2 => n32226, B1 => n1310, B2 => 
                           n43, ZN => n3275);
   U5212 : INV_X1 port map( I => n2319, ZN => n34315);
   U20242 : NAND2_X1 port map( A1 => n18680, A2 => n23468, ZN => n12413);
   U13179 : NAND2_X1 port map( A1 => n23579, A2 => n15624, ZN => n23329);
   U13194 : NAND2_X1 port map( A1 => n7425, A2 => n7427, ZN => n3795);
   U5978 : NOR2_X1 port map( A1 => n23054, A2 => n23048, ZN => n23597);
   U6776 : BUF_X2 port map( I => n9611, Z => n36895);
   U1155 : INV_X1 port map( I => n23873, ZN => n2390);
   U13089 : INV_X1 port map( I => n23695, ZN => n14345);
   U7811 : INV_X1 port map( I => n23900, ZN => n1620);
   U14958 : AOI22_X1 port map( A1 => n18918, A2 => n18917, B1 => n16047, B2 => 
                           n23403, ZN => n23712);
   U1145 : INV_X1 port map( I => n23667, ZN => n1617);
   U2141 : INV_X1 port map( I => n18301, ZN => n34498);
   U28056 : INV_X1 port map( I => n23655, ZN => n24005);
   U1144 : INV_X1 port map( I => n17925, ZN => n23930);
   U13088 : INV_X1 port map( I => n16055, ZN => n23661);
   U1829 : INV_X1 port map( I => n23778, ZN => n31227);
   U3007 : INV_X1 port map( I => n9979, ZN => n12174);
   U9003 : INV_X1 port map( I => n34269, ZN => n15532);
   U6324 : INV_X1 port map( I => n23671, ZN => n24024);
   U6786 : INV_X1 port map( I => n24015, ZN => n3571);
   U1131 : BUF_X2 port map( I => n24463, Z => n19864);
   U27146 : INV_X2 port map( I => n18178, ZN => n18402);
   U28803 : NAND2_X1 port map( A1 => n17076, A2 => n19864, ZN => n24134);
   U6822 : BUF_X2 port map( I => n4243, Z => n33061);
   U12973 : NOR2_X1 port map( A1 => n9371, A2 => n17911, ZN => n9370);
   U13052 : BUF_X2 port map( I => n24164, Z => n24346);
   U1077 : INV_X1 port map( I => n1609, ZN => n24478);
   U1791 : INV_X1 port map( I => n24196, ZN => n31452);
   U6805 : NAND2_X1 port map( A1 => n12733, A2 => n24327, ZN => n24329);
   U22682 : CLKBUF_X2 port map( I => n9520, Z => n33712);
   U5033 : INV_X1 port map( I => n24169, ZN => n24398);
   U7039 : NAND2_X1 port map( A1 => n24087, A2 => n802, ZN => n24223);
   U12996 : BUF_X2 port map( I => n24404, Z => n12360);
   U3377 : BUF_X2 port map( I => n24287, Z => n232);
   U5300 : INV_X2 port map( I => n6515, ZN => n24282);
   U2206 : BUF_X2 port map( I => n31403, Z => n8735);
   U15201 : INV_X2 port map( I => n2741, ZN => n14392);
   U6536 : INV_X1 port map( I => n16832, ZN => n1285);
   U9829 : INV_X1 port map( I => n13144, ZN => n1283);
   U7941 : INV_X2 port map( I => n18402, ZN => n17066);
   U15863 : INV_X1 port map( I => n15892, ZN => n18238);
   U7897 : INV_X1 port map( I => n7240, ZN => n16377);
   U8342 : INV_X1 port map( I => n17709, ZN => n24143);
   U23367 : INV_X1 port map( I => n12138, ZN => n19880);
   U8348 : INV_X1 port map( I => n37230, ZN => n1282);
   U13043 : NAND2_X1 port map( A1 => n2192, A2 => n24366, ZN => n4182);
   U1767 : INV_X2 port map( I => n38886, ZN => n2336);
   U18971 : INV_X1 port map( I => n6226, ZN => n21043);
   U7014 : INV_X1 port map( I => n24360, ZN => n24458);
   U15853 : INV_X2 port map( I => n1129, ZN => n1031);
   U24247 : NOR2_X1 port map( A1 => n1131, A2 => n1275, ZN => n17163);
   U6830 : NOR2_X1 port map( A1 => n37134, A2 => n3226, ZN => n3228);
   U3711 : NAND3_X1 port map( A1 => n21310, A2 => n24461, A3 => n19864, ZN => 
                           n24305);
   U8296 : NOR2_X1 port map( A1 => n1595, A2 => n5985, ZN => n4359);
   U8320 : NAND2_X1 port map( A1 => n37045, A2 => n39815, ZN => n24400);
   U1770 : NAND3_X1 port map( A1 => n24390, A2 => n9963, A3 => n13584, ZN => 
                           n30580);
   U4312 : NAND2_X1 port map( A1 => n13884, A2 => n10747, ZN => n12481);
   U4155 : INV_X1 port map( I => n807, ZN => n17040);
   U19458 : INV_X1 port map( I => n39699, ZN => n1035);
   U9811 : INV_X1 port map( I => n33599, ZN => n24283);
   U5972 : INV_X2 port map( I => n19426, ZN => n20863);
   U4679 : NOR2_X1 port map( A1 => n9370, A2 => n24282, ZN => n32322);
   U2094 : INV_X1 port map( I => n13412, ZN => n14004);
   U4699 : BUF_X2 port map( I => n24241, Z => n32360);
   U8149 : INV_X1 port map( I => n39415, ZN => n34210);
   U5732 : INV_X1 port map( I => n9066, ZN => n1599);
   U6288 : AOI21_X1 port map( A1 => n1586, A2 => n17709, B => n36757, ZN => 
                           n6215);
   U12797 : INV_X1 port map( I => n24466, ZN => n12288);
   U12875 : NAND2_X1 port map( A1 => n24312, A2 => n24313, ZN => n12329);
   U5193 : CLKBUF_X2 port map( I => n1609, Z => n36740);
   U9825 : BUF_X2 port map( I => n18721, Z => n12146);
   U1044 : NOR2_X1 port map( A1 => n914, A2 => n14558, ZN => n24338);
   U9788 : INV_X1 port map( I => n16366, ZN => n1594);
   U19565 : INV_X1 port map( I => n18721, ZN => n24258);
   U20142 : INV_X1 port map( I => n24279, ZN => n32891);
   U1086 : NAND2_X1 port map( A1 => n1032, A2 => n13555, ZN => n7082);
   U18848 : NOR2_X1 port map( A1 => n1129, A2 => n24140, ZN => n24141);
   U26437 : NOR2_X1 port map( A1 => n12733, A2 => n2396, ZN => n24166);
   U8347 : INV_X1 port map( I => n24287, ZN => n1602);
   U8353 : INV_X1 port map( I => n35134, ZN => n1284);
   U17515 : OR2_X1 port map( A1 => n10073, A2 => n5211, Z => n17456);
   U6312 : INV_X1 port map( I => n24116, ZN => n1274);
   U2082 : INV_X1 port map( I => n16459, ZN => n33077);
   U18559 : INV_X1 port map( I => n18342, ZN => n20027);
   U5973 : INV_X1 port map( I => n33939, ZN => n24295);
   U20627 : INV_X1 port map( I => n17871, ZN => n7883);
   U9738 : AOI21_X1 port map( A1 => n1033, A2 => n24346, B => n34330, ZN => 
                           n23702);
   U3716 : NOR2_X1 port map( A1 => n24134, A2 => n21310, ZN => n18276);
   U2021 : NAND2_X1 port map( A1 => n5953, A2 => n24346, ZN => n35916);
   U5733 : NAND2_X1 port map( A1 => n34547, A2 => n9066, ZN => n24293);
   U2689 : AOI22_X1 port map( A1 => n24231, A2 => n15385, B1 => n1595, B2 => 
                           n24335, ZN => n4360);
   U5147 : OAI21_X1 port map( A1 => n38302, A2 => n24469, B => n5599, ZN => 
                           n35504);
   U7023 : NOR3_X1 port map( A1 => n1609, A2 => n3869, A3 => n94, ZN => n15755)
                           ;
   U26670 : NOR2_X1 port map( A1 => n23702, A2 => n23704, ZN => n36343);
   U1753 : NOR2_X1 port map( A1 => n24412, A2 => n24411, ZN => n4308);
   U19628 : INV_X1 port map( I => n36852, ZN => n13167);
   U12998 : NOR2_X1 port map( A1 => n18116, A2 => n2192, ZN => n3620);
   U1061 : OAI21_X1 port map( A1 => n23820, A2 => n14704, B => n15018, ZN => 
                           n9846);
   U6847 : NOR2_X1 port map( A1 => n8735, A2 => n18920, ZN => n15872);
   U1036 : NOR2_X1 port map( A1 => n19426, A2 => n8193, ZN => n13350);
   U1066 : NAND2_X1 port map( A1 => n17711, A2 => n14378, ZN => n19026);
   U9787 : NOR2_X1 port map( A1 => n35314, A2 => n33061, ZN => n14899);
   U6286 : OAI21_X1 port map( A1 => n24136, A2 => n24267, B => n19745, ZN => 
                           n24139);
   U15329 : NOR2_X1 port map( A1 => n24233, A2 => n23694, ZN => n15206);
   U3712 : NOR2_X1 port map( A1 => n19864, A2 => n21310, ZN => n12286);
   U25044 : OAI21_X1 port map( A1 => n2336, A2 => n7440, B => n2439, ZN => 
                           n36154);
   U1742 : INV_X1 port map( I => n4475, ZN => n9909);
   U21215 : OAI21_X1 port map( A1 => n11169, A2 => n19864, B => n19466, ZN => 
                           n32247);
   U21728 : OAI21_X1 port map( A1 => n24166, A2 => n24327, B => n1607, ZN => 
                           n24167);
   U1048 : NAND3_X1 port map( A1 => n12367, A2 => n19007, A3 => n7082, ZN => 
                           n7081);
   U10659 : OAI21_X1 port map( A1 => n24214, A2 => n18402, B => n7210, ZN => 
                           n7209);
   U12887 : NAND2_X1 port map( A1 => n23844, A2 => n24395, ZN => n18101);
   U9816 : NOR2_X1 port map( A1 => n12771, A2 => n9844, ZN => n10695);
   U28844 : NAND2_X1 port map( A1 => n19415, A2 => n18455, ZN => n24429);
   U2041 : NAND3_X1 port map( A1 => n15145, A2 => n15146, A3 => n24330, ZN => 
                           n36209);
   U9752 : NOR2_X1 port map( A1 => n13708, A2 => n1601, ZN => n13707);
   U15930 : AOI22_X1 port map( A1 => n11132, A2 => n24119, B1 => n14684, B2 => 
                           n23819, ZN => n11131);
   U9760 : NAND2_X1 port map( A1 => n24114, A2 => n12771, ZN => n7344);
   U23110 : NAND2_X1 port map( A1 => n11673, A2 => n24245, ZN => n21081);
   U7902 : INV_X1 port map( I => n24140, ZN => n24459);
   U4617 : BUF_X2 port map( I => n16445, Z => n14705);
   U3392 : NOR2_X1 port map( A1 => n1593, A2 => n35244, ZN => n24165);
   U7017 : INV_X1 port map( I => n1128, ZN => n1588);
   U9804 : INV_X1 port map( I => n19857, ZN => n1604);
   U7746 : AND2_X1 port map( A1 => n32518, A2 => n9520, Z => n34080);
   U2969 : AOI21_X1 port map( A1 => n13446, A2 => n1032, B => n13444, ZN => 
                           n13445);
   U6062 : AND2_X1 port map( A1 => n18721, A2 => n18269, Z => n34044);
   U9692 : NOR2_X1 port map( A1 => n11317, A2 => n34074, ZN => n9805);
   U5719 : OAI22_X1 port map( A1 => n24293, A2 => n326, B1 => n1599, B2 => 
                           n24295, ZN => n8840);
   U24077 : NAND2_X1 port map( A1 => n24353, A2 => n24233, ZN => n13625);
   U19593 : AOI21_X1 port map( A1 => n37134, A2 => n24298, B => n17081, ZN => 
                           n13308);
   U6857 : AOI22_X1 port map( A1 => n24149, A2 => n12248, B1 => n20839, B2 => 
                           n24207, ZN => n7179);
   U6293 : OAI21_X1 port map( A1 => n18698, A2 => n18697, B => n24274, ZN => 
                           n19537);
   U17821 : NAND3_X1 port map( A1 => n37651, A2 => n24407, A3 => n39504, ZN => 
                           n20583);
   U30294 : NAND2_X1 port map( A1 => n33727, A2 => n12360, ZN => n17299);
   U9705 : AOI21_X1 port map( A1 => n10220, A2 => n9101, B => n15049, ZN => 
                           n9888);
   U1969 : OAI21_X1 port map( A1 => n2348, A2 => n39478, B => n36561, ZN => 
                           n16069);
   U1928 : OAI21_X1 port map( A1 => n35873, A2 => n35872, B => n18348, ZN => 
                           n30914);
   U6865 : OAI21_X1 port map( A1 => n16829, A2 => n14630, B => n36378, ZN => 
                           n6953);
   U18916 : NAND2_X1 port map( A1 => n39478, A2 => n9963, ZN => n24391);
   U6850 : AOI21_X1 port map( A1 => n19382, A2 => n1127, B => n24102, ZN => 
                           n30652);
   U1986 : NAND2_X1 port map( A1 => n13386, A2 => n36852, ZN => n9840);
   U28822 : NAND2_X1 port map( A1 => n807, A2 => n1601, ZN => n24265);
   U22345 : NOR2_X1 port map( A1 => n24402, A2 => n32484, ZN => n13741);
   U6829 : INV_X1 port map( I => n24129, ZN => n3949);
   U23985 : AOI21_X1 port map( A1 => n19426, A2 => n38302, B => n20537, ZN => 
                           n13481);
   U12943 : NOR2_X1 port map( A1 => n11758, A2 => n24173, ZN => n9842);
   U12852 : OAI22_X1 port map( A1 => n19381, A2 => n24176, B1 => n24336, B2 => 
                           n18295, ZN => n6956);
   U21430 : NAND2_X1 port map( A1 => n31270, A2 => n37803, ZN => n19052);
   U22627 : NOR2_X1 port map( A1 => n35815, A2 => n35814, ZN => n1949);
   U12963 : NOR2_X1 port map( A1 => n585, A2 => n32507, ZN => n34690);
   U19100 : NAND2_X1 port map( A1 => n7083, A2 => n7081, ZN => n6357);
   U14702 : NOR2_X1 port map( A1 => n17509, A2 => n24459, ZN => n34899);
   U21103 : AOI21_X1 port map( A1 => n24401, A2 => n8581, B => n39703, ZN => 
                           n24301);
   U12903 : NOR2_X1 port map( A1 => n19682, A2 => n36378, ZN => n9931);
   U26358 : INV_X1 port map( I => n33108, ZN => n23765);
   U1759 : OAI21_X1 port map( A1 => n24441, A2 => n20903, B => n19584, ZN => 
                           n33616);
   U20590 : OAI22_X1 port map( A1 => n7800, A2 => n24346, B1 => n39156, B2 => 
                           n24348, ZN => n12050);
   U19505 : NAND2_X1 port map( A1 => n13481, A2 => n19052, ZN => n35348);
   U10751 : OAI21_X1 port map( A1 => n34899, A2 => n35854, B => n19895, ZN => 
                           n34437);
   U1672 : INV_X1 port map( I => n24746, ZN => n16196);
   U3973 : CLKBUF_X2 port map( I => n24864, Z => n32093);
   U1643 : CLKBUF_X2 port map( I => n24661, Z => n16210);
   U1669 : CLKBUF_X2 port map( I => n3760, Z => n3487);
   U13510 : OAI21_X1 port map( A1 => n13351, A2 => n13350, B => n5613, ZN => 
                           n31519);
   U23619 : INV_X2 port map( I => n24634, ZN => n12672);
   U5704 : INV_X2 port map( I => n17986, ZN => n24630);
   U6890 : INV_X2 port map( I => n15281, ZN => n934);
   U4249 : INV_X2 port map( I => n9197, ZN => n457);
   U1844 : NAND2_X1 port map( A1 => n12672, A2 => n36634, ZN => n36690);
   U4048 : INV_X1 port map( I => n19713, ZN => n24876);
   U20221 : INV_X2 port map( I => n10116, ZN => n32064);
   U1886 : INV_X2 port map( I => n11081, ZN => n13495);
   U14275 : INV_X1 port map( I => n13221, ZN => n24833);
   U8250 : INV_X1 port map( I => n24589, ZN => n1263);
   U21709 : BUF_X2 port map( I => n17986, Z => n33012);
   U8144 : NAND2_X1 port map( A1 => n37389, A2 => n24589, ZN => n34199);
   U25924 : NAND2_X1 port map( A1 => n24226, A2 => n2747, ZN => n25018);
   U1815 : CLKBUF_X2 port map( I => n24683, Z => n33392);
   U15871 : NOR2_X1 port map( A1 => n15332, A2 => n24847, ZN => n36955);
   U1673 : INV_X1 port map( I => n16238, ZN => n7198);
   U1897 : INV_X1 port map( I => n1265, ZN => n34198);
   U6994 : INV_X2 port map( I => n5056, ZN => n24692);
   U12679 : NAND2_X1 port map( A1 => n9581, A2 => n9580, ZN => n9578);
   U5952 : INV_X1 port map( I => n17101, ZN => n1267);
   U993 : INV_X1 port map( I => n24814, ZN => n24853);
   U1629 : INV_X1 port map( I => n24686, ZN => n31712);
   U8247 : INV_X1 port map( I => n7770, ZN => n36716);
   U17043 : INV_X1 port map( I => n20326, ZN => n24826);
   U1834 : NAND2_X1 port map( A1 => n37983, A2 => n24746, ZN => n2906);
   U9623 : NAND2_X1 port map( A1 => n24572, A2 => n24832, ZN => n4188);
   U15182 : NOR2_X1 port map( A1 => n13045, A2 => n5897, ZN => n6492);
   U15510 : NAND2_X1 port map( A1 => n13966, A2 => n24864, ZN => n21018);
   U27302 : INV_X2 port map( I => n24883, ZN => n18845);
   U27540 : NOR2_X1 port map( A1 => n16990, A2 => n24737, ZN => n19278);
   U21937 : NOR2_X1 port map( A1 => n24828, A2 => n11081, ZN => n32403);
   U1583 : NOR3_X1 port map( A1 => n1271, A2 => n933, A3 => n7286, ZN => n32504
                           );
   U5413 : NAND3_X1 port map( A1 => n16097, A2 => n32045, A3 => n37411, ZN => 
                           n9209);
   U30055 : NAND2_X1 port map( A1 => n24699, A2 => n37097, ZN => n2608);
   U21025 : NAND2_X1 port map( A1 => n24663, A2 => n1029, ZN => n35579);
   U17431 : NOR2_X1 port map( A1 => n19484, A2 => n36376, ZN => n443);
   U6878 : INV_X2 port map( I => n2340, ZN => n15137);
   U5944 : NAND2_X1 port map( A1 => n36988, A2 => n36340, ZN => n15427);
   U28903 : INV_X1 port map( I => n37067, ZN => n24743);
   U28878 : NOR2_X1 port map( A1 => n11271, A2 => n24630, ZN => n24569);
   U3492 : NAND3_X1 port map( A1 => n31625, A2 => n23705, A3 => n2018, ZN => 
                           n20975);
   U21043 : NAND2_X1 port map( A1 => n30282, A2 => n24691, ZN => n32223);
   U977 : INV_X2 port map( I => n24877, ZN => n1119);
   U6883 : BUF_X2 port map( I => n24545, Z => n34666);
   U25713 : INV_X1 port map( I => n15136, ZN => n20930);
   U8142 : NOR2_X1 port map( A1 => n34199, A2 => n34198, ZN => n34197);
   U1650 : BUF_X4 port map( I => n33919, Z => n31161);
   U23783 : BUF_X2 port map( I => n24863, Z => n35968);
   U5375 : BUF_X2 port map( I => n7506, Z => n33317);
   U6282 : INV_X2 port map( I => n6977, ZN => n9212);
   U1806 : INV_X1 port map( I => n36321, ZN => n35521);
   U17710 : CLKBUF_X2 port map( I => n8966, Z => n30554);
   U14264 : INV_X1 port map( I => n24698, ZN => n24900);
   U6908 : NAND3_X1 port map( A1 => n24824, A2 => n24821, A3 => n24819, ZN => 
                           n4351);
   U6893 : INV_X1 port map( I => n30534, ZN => n36920);
   U7690 : AND2_X1 port map( A1 => n24250, A2 => n9385, Z => n34055);
   U5037 : INV_X1 port map( I => n9825, ZN => n4601);
   U15985 : NOR2_X1 port map( A1 => n3510, A2 => n24912, ZN => n5210);
   U5372 : OAI21_X1 port map( A1 => n24789, A2 => n24788, B => n20039, ZN => 
                           n24510);
   U9654 : NAND2_X1 port map( A1 => n957, A2 => n1026, ZN => n13581);
   U3005 : AOI21_X1 port map( A1 => n36988, A2 => n19901, B => n37477, ZN => 
                           n24651);
   U12577 : INV_X1 port map( I => n12643, ZN => n1560);
   U1824 : AOI22_X1 port map( A1 => n17496, A2 => n24799, B1 => n19679, B2 => 
                           n37355, ZN => n34947);
   U9669 : NOR2_X1 port map( A1 => n31698, A2 => n31161, ZN => n4909);
   U22559 : NAND3_X1 port map( A1 => n6822, A2 => n5431, A3 => n24828, ZN => 
                           n24571);
   U10989 : AOI21_X1 port map( A1 => n2904, A2 => n30699, B => n37983, ZN => 
                           n2903);
   U3218 : NAND2_X1 port map( A1 => n1030, A2 => n35952, ZN => n24558);
   U3142 : NAND2_X1 port map( A1 => n14241, A2 => n36340, ZN => n33666);
   U12306 : OAI21_X1 port map( A1 => n14523, A2 => n18504, B => n1263, ZN => 
                           n11907);
   U12620 : NAND2_X1 port map( A1 => n457, A2 => n9198, ZN => n11751);
   U24018 : NOR2_X1 port map( A1 => n24659, A2 => n19, ZN => n36046);
   U1756 : NAND2_X1 port map( A1 => n16815, A2 => n34906, ZN => n34747);
   U2626 : NAND2_X1 port map( A1 => n6838, A2 => n4323, ZN => n6574);
   U9617 : AOI21_X1 port map( A1 => n6337, A2 => n19484, B => n9997, ZN => 
                           n10793);
   U24239 : AOI21_X1 port map( A1 => n2340, A2 => n24664, B => n1029, ZN => 
                           n20927);
   U1811 : NAND2_X1 port map( A1 => n35579, A2 => n35577, ZN => n24666);
   U5916 : NAND2_X1 port map( A1 => n24177, A2 => n19, ZN => n35697);
   U2729 : NAND2_X1 port map( A1 => n3122, A2 => n24593, ZN => n62);
   U14779 : AOI21_X1 port map( A1 => n32403, A2 => n6822, B => n9474, ZN => 
                           n34905);
   U12660 : NAND2_X1 port map( A1 => n24569, A2 => n37106, ZN => n13202);
   U1734 : INV_X1 port map( I => n31161, ZN => n5224);
   U8273 : NOR2_X1 port map( A1 => n35968, A2 => n32093, ZN => n4226);
   U4203 : OAI21_X1 port map( A1 => n2731, A2 => n934, B => n38794, ZN => n2746
                           );
   U9595 : NOR2_X1 port map( A1 => n24965, A2 => n38631, ZN => n9177);
   U6261 : INV_X1 port map( I => n9021, ZN => n11642);
   U7928 : AND2_X1 port map( A1 => n36321, A2 => n16238, Z => n34138);
   U23260 : NOR2_X1 port map( A1 => n19679, A2 => n31213, ZN => n11943);
   U19939 : AOI21_X1 port map( A1 => n934, A2 => n15282, B => n12409, ZN => 
                           n12408);
   U15787 : AOI21_X1 port map( A1 => n24752, A2 => n1576, B => n24664, ZN => 
                           n5245);
   U28773 : OAI21_X1 port map( A1 => n17658, A2 => n18115, B => n2731, ZN => 
                           n11769);
   U8229 : AOI21_X1 port map( A1 => n24639, A2 => n34906, B => n14211, ZN => 
                           n2505);
   U1837 : AOI22_X1 port map( A1 => n3487, A2 => n11846, B1 => n9921, B2 => 
                           n5957, ZN => n12461);
   U3585 : NAND3_X1 port map( A1 => n14241, A2 => n19901, A3 => n38848, ZN => 
                           n15846);
   U25192 : NAND3_X1 port map( A1 => n9656, A2 => n958, A3 => n24692, ZN => 
                           n24210);
   U30027 : OAI22_X1 port map( A1 => n24728, A2 => n25048, B1 => n12672, B2 => 
                           n25053, ZN => n14827);
   U12583 : NAND2_X1 port map( A1 => n24629, A2 => n24821, ZN => n24389);
   U1535 : AOI21_X1 port map( A1 => n6957, A2 => n24696, B => n957, ZN => 
                           n12503);
   U1962 : AOI22_X1 port map( A1 => n24644, A2 => n6977, B1 => n32045, B2 => 
                           n24643, ZN => n9683);
   U14889 : OAI22_X1 port map( A1 => n5653, A2 => n24909, B1 => n25053, B2 => 
                           n37105, ZN => n13030);
   U5424 : NAND2_X1 port map( A1 => n16841, A2 => n24799, ZN => n32643);
   U12556 : NAND2_X1 port map( A1 => n37210, A2 => n24629, ZN => n14165);
   U15132 : NOR2_X1 port map( A1 => n34138, A2 => n1563, ZN => n13340);
   U3672 : NAND2_X1 port map( A1 => n24736, A2 => n7846, ZN => n7845);
   U25652 : AOI21_X1 port map( A1 => n20158, A2 => n38285, B => n33317, ZN => 
                           n17343);
   U4581 : NAND2_X1 port map( A1 => n8317, A2 => n8318, ZN => n8316);
   U12590 : NAND2_X1 port map( A1 => n24709, A2 => n13050, ZN => n13049);
   U950 : AOI21_X1 port map( A1 => n24556, A2 => n19886, B => n14532, ZN => 
                           n15586);
   U1775 : NAND2_X1 port map( A1 => n6023, A2 => n24691, ZN => n36918);
   U12991 : AOI21_X1 port map( A1 => n6707, A2 => n19484, B => n6706, ZN => 
                           n4840);
   U28881 : NAND2_X1 port map( A1 => n24579, A2 => n24578, ZN => n24885);
   U1784 : NAND2_X1 port map( A1 => n36280, A2 => n7831, ZN => n10467);
   U2547 : AOI21_X1 port map( A1 => n14523, A2 => n37687, B => n13628, ZN => 
                           n4703);
   U9609 : NOR2_X1 port map( A1 => n11943, A2 => n36673, ZN => n3879);
   U22571 : OAI22_X1 port map( A1 => n2340, A2 => n35578, B1 => n38523, B2 => 
                           n2341, ZN => n20438);
   U24255 : INV_X1 port map( I => n33271, ZN => n33197);
   U12517 : INV_X1 port map( I => n24991, ZN => n5845);
   U3635 : INV_X1 port map( I => n12534, ZN => n10837);
   U1768 : NOR3_X1 port map( A1 => n20411, A2 => n24847, A3 => n11710, ZN => 
                           n12388);
   U6941 : NAND2_X1 port map( A1 => n20806, A2 => n19507, ZN => n20697);
   U18491 : OAI22_X1 port map( A1 => n24730, A2 => n39157, B1 => n24731, B2 => 
                           n11712, ZN => n35245);
   U4561 : BUF_X2 port map( I => n19725, Z => n32195);
   U15170 : AOI21_X1 port map( A1 => n24531, A2 => n8389, B => n8388, ZN => 
                           n25229);
   U5693 : AOI21_X1 port map( A1 => n24499, A2 => n38369, B => n12207, ZN => 
                           n12206);
   U5427 : INV_X1 port map( I => n24959, ZN => n25225);
   U21794 : INV_X1 port map( I => n3015, ZN => n11756);
   U896 : INV_X1 port map( I => n24994, ZN => n25083);
   U8202 : INV_X1 port map( I => n25263, ZN => n5308);
   U4579 : INV_X1 port map( I => n2653, ZN => n31628);
   U25184 : INV_X1 port map( I => n25160, ZN => n24676);
   U9836 : INV_X1 port map( I => n16526, ZN => n7352);
   U15344 : NAND2_X1 port map( A1 => n16542, A2 => n9528, ZN => n25238);
   U5691 : INV_X1 port map( I => n15030, ZN => n1558);
   U26312 : NOR2_X1 port map( A1 => n25022, A2 => n25021, ZN => n25165);
   U12586 : INV_X1 port map( I => n24985, ZN => n1561);
   U6945 : INV_X1 port map( I => n24922, ZN => n25192);
   U25179 : INV_X1 port map( I => n4302, ZN => n25076);
   U6943 : INV_X1 port map( I => n25247, ZN => n3647);
   U22530 : INV_X1 port map( I => n24927, ZN => n16674);
   U16155 : NAND2_X1 port map( A1 => n817, A2 => n9181, ZN => n25202);
   U6987 : INV_X1 port map( I => n24931, ZN => n4348);
   U30582 : INV_X1 port map( I => n15907, ZN => n8304);
   U13535 : NOR2_X1 port map( A1 => n5100, A2 => n32989, ZN => n31156);
   U3139 : INV_X2 port map( I => n841, ZN => n1116);
   U9580 : BUF_X2 port map( I => n14751, Z => n5798);
   U5041 : INV_X1 port map( I => n34483, ZN => n9740);
   U10664 : INV_X1 port map( I => n34427, ZN => n319);
   U1683 : INV_X1 port map( I => n25421, ZN => n34576);
   U26453 : INV_X1 port map( I => n18121, ZN => n25574);
   U876 : INV_X1 port map( I => n25581, ZN => n1253);
   U8167 : INV_X1 port map( I => n18831, ZN => n19235);
   U25214 : NAND2_X1 port map( A1 => n25558, A2 => n25557, ZN => n17450);
   U3193 : INV_X1 port map( I => n31557, ZN => n36593);
   U9528 : NOR2_X1 port map( A1 => n33826, A2 => n25721, ZN => n10532);
   U1613 : INV_X2 port map( I => n25540, ZN => n36991);
   U1639 : NAND2_X1 port map( A1 => n12309, A2 => n17594, ZN => n20888);
   U3719 : INV_X1 port map( I => n33130, ZN => n9481);
   U24174 : INV_X1 port map( I => n13873, ZN => n16264);
   U11620 : INV_X2 port map( I => n25606, ZN => n31359);
   U1748 : NAND2_X1 port map( A1 => n8771, A2 => n24963, ZN => n4625);
   U19881 : INV_X1 port map( I => n12162, ZN => n7236);
   U3788 : CLKBUF_X2 port map( I => n8069, Z => n2148);
   U5458 : INV_X1 port map( I => n25647, ZN => n32279);
   U21244 : CLKBUF_X2 port map( I => n733, Z => n35611);
   U4530 : CLKBUF_X2 port map( I => n25543, Z => n517);
   U27493 : INV_X2 port map( I => n19153, ZN => n25577);
   U30851 : INV_X2 port map( I => n36105, ZN => n1249);
   U5522 : NAND2_X1 port map( A1 => n25665, A2 => n25361, ZN => n4469);
   U30171 : INV_X1 port map( I => n19941, ZN => n36792);
   U9562 : INV_X2 port map( I => n24536, ZN => n19398);
   U1387 : INV_X1 port map( I => n25600, ZN => n32101);
   U9568 : INV_X1 port map( I => n14473, ZN => n25401);
   U25594 : AND2_X1 port map( A1 => n11060, A2 => n16186, Z => n16316);
   U12480 : INV_X1 port map( I => n31305, ZN => n1551);
   U5942 : INV_X1 port map( I => n21042, ZN => n25670);
   U9529 : INV_X1 port map( I => n33947, ZN => n7802);
   U10529 : INV_X1 port map( I => n39061, ZN => n1022);
   U5683 : INV_X1 port map( I => n25696, ZN => n911);
   U23534 : AND2_X1 port map( A1 => n36105, A2 => n25619, Z => n25142);
   U28861 : NAND2_X1 port map( A1 => n25682, A2 => n30633, ZN => n24535);
   U5843 : NAND2_X1 port map( A1 => n32580, A2 => n30377, ZN => n16372);
   U1363 : NAND3_X1 port map( A1 => n25399, A2 => n25400, A3 => n25401, ZN => 
                           n32789);
   U15349 : NAND2_X1 port map( A1 => n9526, A2 => n25307, ZN => n13849);
   U6906 : NOR2_X1 port map( A1 => n25487, A2 => n35216, ZN => n7052);
   U12388 : NAND2_X1 port map( A1 => n25603, A2 => n14708, ZN => n5857);
   U7926 : INV_X2 port map( I => n25513, ZN => n13461);
   U9488 : NOR2_X1 port map( A1 => n9893, A2 => n826, ZN => n8739);
   U2037 : INV_X1 port map( I => n25484, ZN => n1547);
   U12402 : NAND2_X1 port map( A1 => n12616, A2 => n826, ZN => n9029);
   U1657 : NAND2_X1 port map( A1 => n7705, A2 => n33946, ZN => n25679);
   U823 : NAND2_X1 port map( A1 => n25545, A2 => n1539, ZN => n13375);
   U27888 : AOI21_X1 port map( A1 => n10674, A2 => n19863, B => n25379, ZN => 
                           n12462);
   U12428 : INV_X1 port map( I => n1252, ZN => n6064);
   U870 : INV_X2 port map( I => n14081, ZN => n25642);
   U18245 : NOR2_X1 port map( A1 => n4914, A2 => n11060, ZN => n13468);
   U12316 : NAND2_X1 port map( A1 => n25435, A2 => n25248, ZN => n11441);
   U6249 : NAND2_X1 port map( A1 => n16246, A2 => n19696, ZN => n25698);
   U1286 : AOI21_X1 port map( A1 => n15443, A2 => n19095, B => n31984, ZN => 
                           n31158);
   U9465 : OAI21_X1 port map( A1 => n5011, A2 => n5010, B => n8014, ZN => n5277
                           );
   U12355 : AOI21_X1 port map( A1 => n20440, A2 => n20442, B => n25361, ZN => 
                           n7339);
   U1275 : NOR2_X1 port map( A1 => n14619, A2 => n10530, ZN => n31159);
   U9517 : AOI21_X1 port map( A1 => n7075, A2 => n30694, B => n37905, ZN => 
                           n7926);
   U17465 : INV_X1 port map( I => n15443, ZN => n15329);
   U29571 : INV_X1 port map( I => n6592, ZN => n20855);
   U1581 : NAND2_X1 port map( A1 => n19400, A2 => n14410, ZN => n36907);
   U4428 : INV_X1 port map( I => n138, ZN => n15406);
   U8112 : NAND2_X1 port map( A1 => n12825, A2 => n19581, ZN => n11278);
   U1632 : OR2_X1 port map( A1 => n16203, A2 => n33949, Z => n4384);
   U18573 : AND2_X1 port map( A1 => n25498, A2 => n25380, Z => n12404);
   U3479 : AND2_X1 port map( A1 => n25695, A2 => n25694, Z => n20105);
   U3254 : AND2_X1 port map( A1 => n31669, A2 => n20838, Z => n25514);
   U814 : INV_X1 port map( I => n34150, ZN => n19296);
   U2146 : INV_X1 port map( I => n541, ZN => n15215);
   U6898 : INV_X1 port map( I => n25660, ZN => n25381);
   U1277 : AOI21_X1 port map( A1 => n12394, A2 => n20648, B => n8014, ZN => 
                           n32255);
   U9451 : NAND2_X1 port map( A1 => n4048, A2 => n4664, ZN => n8907);
   U6899 : OAI21_X1 port map( A1 => n10563, A2 => n9915, B => n9441, ZN => 
                           n9440);
   U1546 : NOR2_X1 port map( A1 => n15406, A2 => n36708, ZN => n36941);
   U1463 : NAND2_X1 port map( A1 => n36907, A2 => n1024, ZN => n21220);
   U19435 : OAI21_X1 port map( A1 => n25637, A2 => n6731, B => n37993, ZN => 
                           n20885);
   U12370 : NAND2_X1 port map( A1 => n952, A2 => n15406, ZN => n8568);
   U6954 : NAND2_X1 port map( A1 => n24937, A2 => n14805, ZN => n31165);
   U10963 : INV_X1 port map( I => n20855, ZN => n34464);
   U9555 : NAND2_X1 port map( A1 => n10882, A2 => n16836, ZN => n11641);
   U17261 : NAND2_X1 port map( A1 => n35449, A2 => n18909, ZN => n36217);
   U1522 : NAND2_X1 port map( A1 => n25625, A2 => n25365, ZN => n34719);
   U4049 : AOI21_X1 port map( A1 => n12382, A2 => n33950, B => n12500, ZN => 
                           n35117);
   U4496 : NAND2_X1 port map( A1 => n31984, A2 => n30705, ZN => n9427);
   U12335 : NAND2_X1 port map( A1 => n1112, A2 => n12500, ZN => n4642);
   U14381 : AOI21_X1 port map( A1 => n36345, A2 => n1984, B => n7924, ZN => 
                           n34846);
   U30037 : OAI21_X1 port map( A1 => n25422, A2 => n18031, B => n12309, ZN => 
                           n36755);
   U9456 : OAI21_X1 port map( A1 => n2416, A2 => n2576, B => n33785, ZN => 
                           n11547);
   U23541 : NOR2_X1 port map( A1 => n12675, A2 => n25754, ZN => n32684);
   U30529 : INV_X1 port map( I => n25566, ZN => n33897);
   U24913 : NOR2_X1 port map( A1 => n25474, A2 => n36486, ZN => n16026);
   U2999 : INV_X1 port map( I => n25577, ZN => n25662);
   U12412 : NAND2_X1 port map( A1 => n13016, A2 => n12500, ZN => n13015);
   U12271 : AOI21_X1 port map( A1 => n20746, A2 => n17613, B => n7802, ZN => 
                           n9803);
   U9495 : NOR2_X1 port map( A1 => n11278, A2 => n20052, ZN => n10719);
   U12415 : NOR2_X1 port map( A1 => n25756, A2 => n38338, ZN => n25627);
   U9772 : NOR2_X1 port map( A1 => n31745, A2 => n10034, ZN => n14794);
   U8944 : NAND2_X1 port map( A1 => n32207, A2 => n4214, ZN => n34264);
   U1254 : NOR2_X1 port map( A1 => n10674, A2 => n25660, ZN => n229);
   U1662 : NAND2_X1 port map( A1 => n35882, A2 => n11647, ZN => n30813);
   U12411 : INV_X1 port map( I => n11363, ZN => n14316);
   U9501 : NOR2_X1 port map( A1 => n15172, A2 => n1108, ZN => n15924);
   U3093 : OAI21_X1 port map( A1 => n36486, A2 => n13461, B => n13744, ZN => 
                           n25476);
   U3286 : NOR2_X1 port map( A1 => n25608, A2 => n25472, ZN => n17013);
   U8154 : INV_X1 port map( I => n25545, ZN => n25480);
   U1217 : NAND2_X1 port map( A1 => n25195, A2 => n32722, ZN => n2496);
   U1471 : NOR2_X1 port map( A1 => n25682, A2 => n25681, ZN => n34393);
   U29092 : NAND3_X1 port map( A1 => n20856, A2 => n25677, A3 => n14081, ZN => 
                           n25678);
   U12336 : NAND2_X1 port map( A1 => n25448, A2 => n39371, ZN => n14486);
   U15458 : OAI21_X1 port map( A1 => n3005, A2 => n591, B => n38245, ZN => 
                           n3004);
   U22205 : OAI21_X1 port map( A1 => n14472, A2 => n32450, B => n32449, ZN => 
                           n15881);
   U776 : NOR2_X1 port map( A1 => n32101, A2 => n3058, ZN => n3057);
   U4627 : INV_X2 port map( I => n25887, ZN => n928);
   U18221 : NAND3_X1 port map( A1 => n31707, A2 => n12675, A3 => n9441, ZN => 
                           n25755);
   U27394 : NOR2_X1 port map( A1 => n33251, A2 => n33250, ZN => n2248);
   U1405 : NAND3_X1 port map( A1 => n34078, A2 => n25562, A3 => n35349, ZN => 
                           n1855);
   U3802 : INV_X2 port map( I => n25345, ZN => n9530);
   U18873 : OAI21_X1 port map( A1 => n10973, A2 => n7987, B => n6065, ZN => 
                           n10972);
   U8103 : NAND2_X1 port map( A1 => n4792, A2 => n4791, ZN => n25775);
   U1401 : AOI21_X1 port map( A1 => n2576, A2 => n25623, B => n34719, ZN => 
                           n11548);
   U16146 : NOR2_X1 port map( A1 => n14613, A2 => n16428, ZN => n36897);
   U7069 : INV_X2 port map( I => n18062, ZN => n26016);
   U12228 : NAND2_X1 port map( A1 => n11734, A2 => n26128, ZN => n1827);
   U16489 : INV_X2 port map( I => n25971, ZN => n1019);
   U6859 : INV_X2 port map( I => n8683, ZN => n1012);
   U17864 : INV_X2 port map( I => n9412, ZN => n18406);
   U1314 : NOR2_X1 port map( A1 => n26016, A2 => n26015, ZN => n10850);
   U12234 : NAND2_X1 port map( A1 => n15991, A2 => n37184, ZN => n11952);
   U3948 : NAND2_X1 port map( A1 => n31375, A2 => n26020, ZN => n31312);
   U1396 : OAI21_X1 port map( A1 => n954, A2 => n4914, B => n17353, ZN => 
                           n36624);
   U7058 : INV_X2 port map( I => n17791, ZN => n26135);
   U7741 : BUF_X2 port map( I => n10223, Z => n30595);
   U1399 : NAND2_X1 port map( A1 => n26019, A2 => n26020, ZN => n26045);
   U8051 : INV_X1 port map( I => n18176, ZN => n19793);
   U764 : INV_X1 port map( I => n25993, ZN => n25957);
   U1371 : BUF_X2 port map( I => n35903, Z => n31994);
   U3803 : INV_X1 port map( I => n38416, ZN => n20456);
   U15898 : INV_X1 port map( I => n33879, ZN => n26185);
   U6823 : INV_X1 port map( I => n25941, ZN => n26061);
   U735 : INV_X2 port map( I => n10015, ZN => n5908);
   U28208 : INV_X2 port map( I => n15085, ZN => n36571);
   U1333 : INV_X1 port map( I => n31362, ZN => n25998);
   U7076 : INV_X2 port map( I => n37613, ZN => n11552);
   U1336 : NAND2_X1 port map( A1 => n18176, A2 => n25345, ZN => n25769);
   U1332 : NOR2_X1 port map( A1 => n596, A2 => n25941, ZN => n35720);
   U7077 : NOR2_X1 port map( A1 => n3356, A2 => n36226, ZN => n34382);
   U17766 : NAND2_X1 port map( A1 => n26045, A2 => n5886, ZN => n20088);
   U22033 : NOR2_X1 port map( A1 => n25822, A2 => n18142, ZN => n15832);
   U722 : INV_X1 port map( I => n25798, ZN => n26004);
   U12194 : CLKBUF_X2 port map( I => n8683, Z => n9883);
   U24604 : NAND2_X1 port map( A1 => n25971, A2 => n18661, ZN => n26110);
   U3068 : CLKBUF_X2 port map( I => n6830, Z => n2888);
   U14591 : NAND2_X1 port map( A1 => n1017, A2 => n17180, ZN => n26042);
   U18601 : NAND2_X1 port map( A1 => n25770, A2 => n26063, ZN => n26060);
   U1978 : INV_X1 port map( I => n26001, ZN => n9379);
   U17783 : INV_X1 port map( I => n26116, ZN => n31624);
   U12195 : INV_X1 port map( I => n7136, ZN => n15121);
   U1186 : INV_X1 port map( I => n18827, ZN => n19259);
   U5562 : INV_X2 port map( I => n39030, ZN => n26005);
   U4250 : INV_X1 port map( I => n17180, ZN => n1518);
   U20294 : INV_X1 port map( I => n10834, ZN => n929);
   U16575 : INV_X2 port map( I => n8375, ZN => n6056);
   U17697 : INV_X1 port map( I => n13717, ZN => n9380);
   U16033 : INV_X1 port map( I => n9413, ZN => n12234);
   U1303 : INV_X1 port map( I => n26329, ZN => n1240);
   U730 : INV_X1 port map( I => n2349, ZN => n926);
   U12210 : AOI21_X1 port map( A1 => n25975, A2 => n17458, B => n6056, ZN => 
                           n25793);
   U1089 : INV_X2 port map( I => n6222, ZN => n33365);
   U1130 : NAND3_X1 port map( A1 => n13869, A2 => n38548, A3 => n10724, ZN => 
                           n2418);
   U29127 : NOR2_X1 port map( A1 => n25876, A2 => n25875, ZN => n25877);
   U8718 : NAND3_X1 port map( A1 => n38548, A2 => n35003, A3 => n14212, ZN => 
                           n30674);
   U25248 : AOI21_X1 port map( A1 => n33263, A2 => n15178, B => n18884, ZN => 
                           n15177);
   U9378 : NAND2_X1 port map( A1 => n14375, A2 => n31263, ZN => n4293);
   U14581 : NOR2_X1 port map( A1 => n8156, A2 => n25738, ZN => n10510);
   U8041 : NOR2_X1 port map( A1 => n6506, A2 => n8683, ZN => n25760);
   U1248 : NOR2_X1 port map( A1 => n32196, A2 => n31340, ZN => n35046);
   U18574 : NOR2_X1 port map( A1 => n25874, A2 => n4322, ZN => n2891);
   U28982 : OAI21_X1 port map( A1 => n25995, A2 => n318, B => n25111, ZN => 
                           n25110);
   U7086 : NAND2_X1 port map( A1 => n11807, A2 => n9883, ZN => n24917);
   U12102 : NAND2_X1 port map( A1 => n10062, A2 => n1102, ZN => n8710);
   U25238 : NAND2_X1 port map( A1 => n25657, A2 => n34402, ZN => n19214);
   U12012 : INV_X1 port map( I => n26083, ZN => n11773);
   U16125 : INV_X1 port map( I => n7961, ZN => n33366);
   U12244 : INV_X1 port map( I => n9694, ZN => n26032);
   U17284 : NOR2_X1 port map( A1 => n30302, A2 => n4163, ZN => n25788);
   U4409 : INV_X1 port map( I => n35855, ZN => n1527);
   U14965 : BUF_X2 port map( I => n26054, Z => n32109);
   U18025 : BUF_X2 port map( I => n1011, Z => n36722);
   U12205 : INV_X1 port map( I => n19259, ZN => n2835);
   U8077 : INV_X1 port map( I => n11734, ZN => n26126);
   U4465 : CLKBUF_X2 port map( I => n6180, Z => n33795);
   U12204 : CLKBUF_X2 port map( I => n26329, Z => n7460);
   U1271 : NAND2_X1 port map( A1 => n26016, A2 => n26015, ZN => n26123);
   U14780 : NAND2_X1 port map( A1 => n1239, A2 => n586, ZN => n25745);
   U4135 : INV_X1 port map( I => n26031, ZN => n1016);
   U8060 : INV_X1 port map( I => n6506, ZN => n15283);
   U12243 : INV_X1 port map( I => n1107, ZN => n12711);
   U10608 : INV_X1 port map( I => n26070, ZN => n15796);
   U6879 : INV_X1 port map( I => n26054, ZN => n1020);
   U5740 : AND2_X1 port map( A1 => n26054, A2 => n2349, Z => n34153);
   U12106 : OAI21_X1 port map( A1 => n25886, A2 => n15796, B => n928, ZN => 
                           n25858);
   U684 : AOI22_X1 port map( A1 => n25862, A2 => n33218, B1 => n38982, B2 => 
                           n25861, ZN => n15946);
   U7109 : BUF_X2 port map( I => n25836, Z => n31954);
   U12162 : AOI22_X1 port map( A1 => n33348, A2 => n26050, B1 => n31311, B2 => 
                           n1523, ZN => n26051);
   U2568 : OAI22_X1 port map( A1 => n32056, A2 => n32690, B1 => n26005, B2 => 
                           n26006, ZN => n25531);
   U24608 : NAND2_X1 port map( A1 => n20813, A2 => n31340, ZN => n26213);
   U6201 : NAND3_X1 port map( A1 => n10724, A2 => n30937, A3 => n12199, ZN => 
                           n12152);
   U8867 : NOR2_X1 port map( A1 => n16200, A2 => n38760, ZN => n19218);
   U12049 : AOI21_X1 port map( A1 => n5326, A2 => n25870, B => n17501, ZN => 
                           n5325);
   U659 : NAND3_X1 port map( A1 => n30900, A2 => n425, A3 => n32052, ZN => 
                           n25406);
   U12145 : NAND2_X1 port map( A1 => n25855, A2 => n26004, ZN => n16612);
   U11034 : AOI21_X1 port map( A1 => n25768, A2 => n4832, B => n1097, ZN => 
                           n21307);
   U14726 : AOI22_X1 port map( A1 => n31299, A2 => n9743, B1 => n927, B2 => 
                           n949, ZN => n19368);
   U1054 : NOR2_X1 port map( A1 => n9568, A2 => n15703, ZN => n31470);
   U7105 : OAI21_X1 port map( A1 => n17502, A2 => n950, B => n10765, ZN => 
                           n26099);
   U19147 : NOR2_X1 port map( A1 => n25771, A2 => n35109, ZN => n6401);
   U23128 : OAI21_X1 port map( A1 => n6578, A2 => n34018, B => n35891, ZN => 
                           n9087);
   U1190 : OAI21_X1 port map( A1 => n34519, A2 => n25996, B => n11834, ZN => 
                           n11625);
   U18417 : NAND3_X1 port map( A1 => n16478, A2 => n16477, A3 => n34265, ZN => 
                           n20507);
   U7934 : OAI21_X1 port map( A1 => n32109, A2 => n25745, B => n30611, ZN => 
                           n25746);
   U7063 : NOR2_X1 port map( A1 => n17951, A2 => n14375, ZN => n26186);
   U17921 : NOR3_X1 port map( A1 => n14564, A2 => n31994, A3 => n19898, ZN => 
                           n12709);
   U8717 : NAND2_X1 port map( A1 => n30425, A2 => n30674, ZN => n30934);
   U9375 : NAND3_X1 port map( A1 => n25922, A2 => n18038, A3 => n25803, ZN => 
                           n13165);
   U5674 : BUF_X2 port map( I => n26113, Z => n1521);
   U29111 : NAND3_X1 port map( A1 => n26030, A2 => n10062, A3 => n25965, ZN => 
                           n25796);
   U26997 : NOR2_X1 port map( A1 => n362, A2 => n25835, ZN => n18376);
   U18290 : NAND2_X1 port map( A1 => n5886, A2 => n38531, ZN => n5882);
   U20853 : OR2_X1 port map( A1 => n14854, A2 => n32185, Z => n3361);
   U6158 : INV_X1 port map( I => n26215, ZN => n1529);
   U6214 : INV_X1 port map( I => n8120, ZN => n26078);
   U12082 : INV_X1 port map( I => n26214, ZN => n26212);
   U23358 : NAND2_X1 port map( A1 => n12721, A2 => n32243, ZN => n13281);
   U30826 : NOR2_X1 port map( A1 => n362, A2 => n18375, ZN => n5283);
   U18642 : OAI21_X1 port map( A1 => n26078, A2 => n26075, B => n11762, ZN => 
                           n12151);
   U7980 : AOI22_X1 port map( A1 => n14685, A2 => n6578, B1 => n6302, B2 => 
                           n26061, ZN => n4430);
   U16375 : NAND2_X1 port map( A1 => n35099, A2 => n25977, ZN => n2574);
   U12120 : NAND2_X1 port map( A1 => n25898, A2 => n36293, ZN => n6396);
   U26613 : OAI21_X1 port map( A1 => n36819, A2 => n1015, B => n36581, ZN => 
                           n25838);
   U1136 : AOI22_X1 port map( A1 => n5283, A2 => n1015, B1 => n14694, B2 => 
                           n362, ZN => n34499);
   U27382 : INV_X1 port map( I => n25919, ZN => n18863);
   U7116 : INV_X1 port map( I => n10225, ZN => n31073);
   U4319 : NAND2_X1 port map( A1 => n25831, A2 => n25921, ZN => n25834);
   U640 : BUF_X2 port map( I => n9858, Z => n343);
   U5666 : OAI21_X1 port map( A1 => n14984, A2 => n25749, B => n14983, ZN => 
                           n26165);
   U21416 : OAI21_X1 port map( A1 => n3361, A2 => n3360, B => n35646, ZN => 
                           n3781);
   U14570 : NAND2_X1 port map( A1 => n9077, A2 => n20116, ZN => n26530);
   U3621 : BUF_X2 port map( I => n11752, Z => n291);
   U6811 : INV_X1 port map( I => n6154, ZN => n16294);
   U17617 : NOR2_X1 port map( A1 => n26078, A2 => n9855, ZN => n2421);
   U1016 : NAND2_X1 port map( A1 => n34148, A2 => n18273, ZN => n7862);
   U26588 : INV_X1 port map( I => n26585, ZN => n36333);
   U12005 : INV_X1 port map( I => n32095, ZN => n9870);
   U1599 : INV_X1 port map( I => n17263, ZN => n8110);
   U7963 : INV_X1 port map( I => n1009, ZN => n11298);
   U2131 : NAND2_X1 port map( A1 => n7603, A2 => n7602, ZN => n7781);
   U14386 : AOI22_X1 port map( A1 => n32747, A2 => n32748, B1 => n26097, B2 => 
                           n39351, ZN => n35239);
   U15111 : BUF_X2 port map( I => n4828, Z => n36958);
   U20345 : INV_X1 port map( I => n34768, ZN => n35463);
   U12001 : INV_X1 port map( I => n26436, ZN => n16830);
   U9360 : NAND2_X1 port map( A1 => n3100, A2 => n1504, ZN => n3099);
   U11976 : INV_X1 port map( I => n32464, ZN => n20843);
   U623 : INV_X1 port map( I => n13062, ZN => n26729);
   U6778 : BUF_X2 port map( I => n26861, Z => n8817);
   U1082 : BUF_X2 port map( I => n19423, Z => n34005);
   U17785 : INV_X2 port map( I => n12682, ZN => n14380);
   U16889 : INV_X2 port map( I => n13605, ZN => n26933);
   U7915 : INV_X1 port map( I => n26861, ZN => n20223);
   U26192 : INV_X1 port map( I => n36292, ZN => n14453);
   U1081 : INV_X1 port map( I => n740, ZN => n33858);
   U11972 : INV_X1 port map( I => n37054, ZN => n1787);
   U5362 : INV_X1 port map( I => n30284, ZN => n20004);
   U962 : BUF_X2 port map( I => n10355, Z => n33689);
   U1034 : INV_X2 port map( I => n167, ZN => n26944);
   U7909 : BUF_X2 port map( I => n11335, Z => n11334);
   U13250 : NAND2_X1 port map( A1 => n19353, A2 => n33561, ZN => n26987);
   U4410 : BUF_X2 port map( I => n13528, Z => n33849);
   U16312 : CLKBUF_X2 port map( I => n19615, Z => n36882);
   U10744 : INV_X2 port map( I => n30853, ZN => n14355);
   U4196 : BUF_X2 port map( I => n6454, Z => n441);
   U5656 : INV_X2 port map( I => n26992, ZN => n26692);
   U987 : INV_X1 port map( I => n39825, ZN => n17655);
   U7958 : INV_X1 port map( I => n9118, ZN => n9117);
   U23229 : INV_X1 port map( I => n17252, ZN => n11864);
   U18917 : INV_X1 port map( I => n26746, ZN => n20120);
   U16503 : INV_X2 port map( I => n36392, ZN => n1002);
   U2899 : INV_X1 port map( I => n18210, ZN => n1008);
   U30829 : INV_X1 port map( I => n17022, ZN => n26986);
   U592 : INV_X1 port map( I => n34005, ZN => n26903);
   U550 : INV_X1 port map( I => n10355, ZN => n1491);
   U585 : INV_X2 port map( I => n8527, ZN => n26857);
   U3924 : NOR3_X1 port map( A1 => n15411, A2 => n17217, A3 => n33726, ZN => 
                           n32849);
   U22931 : INV_X1 port map( I => n34160, ZN => n14455);
   U6754 : INV_X2 port map( I => n17047, ZN => n11679);
   U21409 : NAND2_X1 port map( A1 => n11138, A2 => n14412, ZN => n9062);
   U2279 : NAND2_X1 port map( A1 => n26920, A2 => n38188, ZN => n33063);
   U13588 : NOR2_X1 port map( A1 => n1497, A2 => n15996, ZN => n34767);
   U29322 : NOR2_X1 port map( A1 => n20399, A2 => n26863, ZN => n26864);
   U15288 : NOR2_X1 port map( A1 => n26943, A2 => n15670, ZN => n33548);
   U19191 : INV_X1 port map( I => n6454, ZN => n10479);
   U7937 : INV_X1 port map( I => n35197, ZN => n26825);
   U5641 : INV_X1 port map( I => n13056, ZN => n8816);
   U11863 : NOR2_X1 port map( A1 => n14488, A2 => n36882, ZN => n21192);
   U11807 : INV_X1 port map( I => n26950, ZN => n8815);
   U934 : INV_X1 port map( I => n1003, ZN => n32344);
   U887 : INV_X1 port map( I => n14065, ZN => n31225);
   U24812 : NOR2_X1 port map( A1 => n1092, A2 => n13757, ZN => n3961);
   U6779 : INV_X2 port map( I => n14636, ZN => n26701);
   U11946 : INV_X2 port map( I => n4411, ZN => n4007);
   U7895 : NOR2_X1 port map( A1 => n8814, A2 => n8817, ZN => n26731);
   U907 : INV_X1 port map( I => n26860, ZN => n8415);
   U881 : NAND2_X1 port map( A1 => n33849, A2 => n37098, ZN => n31670);
   U5218 : INV_X1 port map( I => n37103, ZN => n1090);
   U21108 : NAND2_X1 port map( A1 => n10355, A2 => n14383, ZN => n15371);
   U15211 : INV_X1 port map( I => n2752, ZN => n26800);
   U1018 : INV_X2 port map( I => n858, ZN => n1490);
   U24471 : INV_X1 port map( I => n26763, ZN => n26923);
   U9300 : INV_X1 port map( I => n14459, ZN => n1229);
   U25629 : INV_X1 port map( I => n32986, ZN => n849);
   U9341 : INV_X1 port map( I => n26770, ZN => n18903);
   U4546 : AOI21_X1 port map( A1 => n5935, A2 => n858, B => n20423, ZN => 
                           n15998);
   U553 : INV_X1 port map( I => n9618, ZN => n26740);
   U23261 : INV_X1 port map( I => n11948, ZN => n17034);
   U5657 : INV_X1 port map( I => n30859, ZN => n13088);
   U26505 : INV_X1 port map( I => n26795, ZN => n20699);
   U9336 : NAND2_X1 port map( A1 => n3449, A2 => n20399, ZN => n3919);
   U9301 : NOR2_X1 port map( A1 => n31982, A2 => n12682, ZN => n3742);
   U5690 : NAND2_X1 port map( A1 => n11696, A2 => n17515, ZN => n15650);
   U25401 : OAI22_X1 port map( A1 => n31670, A2 => n6891, B1 => n26653, B2 => 
                           n37856, ZN => n36655);
   U952 : NAND3_X1 port map( A1 => n26828, A2 => n11138, A3 => n17260, ZN => 
                           n36974);
   U4018 : NOR3_X1 port map( A1 => n30665, A2 => n26961, A3 => n2292, ZN => 
                           n35403);
   U11850 : OAI21_X1 port map( A1 => n14732, A2 => n2491, B => n13588, ZN => 
                           n12887);
   U7281 : NOR2_X1 port map( A1 => n2226, A2 => n32168, ZN => n4172);
   U11760 : NOR2_X1 port map( A1 => n13427, A2 => n37856, ZN => n7627);
   U6760 : OAI21_X1 port map( A1 => n26720, A2 => n1234, B => n735, ZN => 
                           n13454);
   U16918 : OAI21_X1 port map( A1 => n26996, A2 => n14459, B => n26692, ZN => 
                           n13036);
   U996 : OAI21_X1 port map( A1 => n26951, A2 => n31701, B => n35409, ZN => 
                           n31638);
   U24048 : NOR2_X1 port map( A1 => n8478, A2 => n2752, ZN => n10678);
   U999 : NAND2_X1 port map( A1 => n10314, A2 => n5537, ZN => n36147);
   U19273 : NAND2_X1 port map( A1 => n441, A2 => n26639, ZN => n6555);
   U3006 : NAND2_X1 port map( A1 => n8817, A2 => n26780, ZN => n34426);
   U11964 : NAND2_X1 port map( A1 => n26876, A2 => n14455, ZN => n12328);
   U3054 : NAND2_X1 port map( A1 => n26833, A2 => n26724, ZN => n2882);
   U29193 : NAND2_X1 port map( A1 => n26992, A2 => n19364, ZN => n26284);
   U2985 : INV_X2 port map( I => n862, ZN => n18809);
   U24637 : NAND2_X1 port map( A1 => n33279, A2 => n26970, ZN => n15196);
   U30654 : NOR2_X1 port map( A1 => n36929, A2 => n37055, ZN => n31277);
   U930 : NAND3_X1 port map( A1 => n19939, A2 => n37154, A3 => n11334, ZN => 
                           n32036);
   U7223 : NAND2_X1 port map( A1 => n1490, A2 => n5935, ZN => n15823);
   U19266 : AOI21_X1 port map( A1 => n34061, A2 => n11707, B => n36647, ZN => 
                           n35321);
   U2944 : NOR2_X1 port map( A1 => n26857, A2 => n19728, ZN => n35028);
   U30089 : OAI21_X1 port map( A1 => n34108, A2 => n13487, B => n33396, ZN => 
                           n36769);
   U6691 : AOI21_X1 port map( A1 => n32941, A2 => n26679, B => n36078, ZN => 
                           n30500);
   U17539 : NOR2_X1 port map( A1 => n167, A2 => n26614, ZN => n19206);
   U28379 : NAND2_X1 port map( A1 => n14134, A2 => n12220, ZN => n36582);
   U3357 : NAND2_X1 port map( A1 => n1492, A2 => n2140, ZN => n26976);
   U11884 : NOR2_X1 port map( A1 => n852, A2 => n26979, ZN => n14831);
   U1995 : OAI21_X1 port map( A1 => n1088, A2 => n14636, B => n26700, ZN => 
                           n10441);
   U15302 : INV_X2 port map( I => n38519, ZN => n8154);
   U21532 : NAND2_X1 port map( A1 => n9269, A2 => n19225, ZN => n26834);
   U23033 : OAI21_X1 port map( A1 => n26700, A2 => n14636, B => n36244, ZN => 
                           n32602);
   U30553 : INV_X1 port map( I => n3574, ZN => n26663);
   U7210 : INV_X1 port map( I => n7596, ZN => n26710);
   U6796 : INV_X1 port map( I => n13393, ZN => n1232);
   U17248 : OAI22_X1 port map( A1 => n15650, A2 => n18809, B1 => n10479, B2 => 
                           n11696, ZN => n18776);
   U21427 : NAND3_X1 port map( A1 => n13801, A2 => n14807, A3 => n1493, ZN => 
                           n9098);
   U9292 : OAI21_X1 port map( A1 => n13758, A2 => n26220, B => n1092, ZN => 
                           n7691);
   U20661 : OAI21_X1 port map( A1 => n38852, A2 => n38928, B => n26772, ZN => 
                           n19172);
   U943 : NAND3_X1 port map( A1 => n16686, A2 => n14488, A3 => n36882, ZN => 
                           n26427);
   U24941 : AOI21_X1 port map( A1 => n18587, A2 => n19331, B => n14921, ZN => 
                           n18586);
   U19227 : AOI21_X1 port map( A1 => n39824, A2 => n26899, B => n26898, ZN => 
                           n35311);
   U519 : NOR2_X1 port map( A1 => n17574, A2 => n17573, ZN => n19687);
   U8926 : NAND2_X1 port map( A1 => n17097, A2 => n33301, ZN => n34262);
   U29316 : OAI21_X1 port map( A1 => n1091, A2 => n26802, B => n26801, ZN => 
                           n26806);
   U931 : NAND2_X1 port map( A1 => n26877, A2 => n17655, ZN => n13870);
   U948 : NOR2_X1 port map( A1 => n26909, A2 => n9117, ZN => n26787);
   U9230 : NAND2_X1 port map( A1 => n27141, A2 => n946, ZN => n17916);
   U899 : NAND2_X1 port map( A1 => n26653, A2 => n36424, ZN => n31678);
   U9330 : NOR2_X1 port map( A1 => n8155, A2 => n38519, ZN => n7511);
   U15394 : NOR2_X1 port map( A1 => n30347, A2 => n10202, ZN => n36164);
   U959 : NAND2_X1 port map( A1 => n1494, A2 => n37103, ZN => n26838);
   U22316 : NAND3_X1 port map( A1 => n15341, A2 => n14097, A3 => n39117, ZN => 
                           n35772);
   U11809 : NAND2_X1 port map( A1 => n8652, A2 => n35537, ZN => n2129);
   U10293 : OAI21_X1 port map( A1 => n36146, A2 => n36147, B => n34396, ZN => 
                           n32577);
   U26179 : NAND3_X1 port map( A1 => n16686, A2 => n26826, A3 => n18903, ZN => 
                           n26425);
   U20765 : NOR2_X1 port map( A1 => n33633, A2 => n34034, ZN => n33631);
   U889 : NAND2_X1 port map( A1 => n30665, A2 => n35764, ZN => n27129);
   U26321 : INV_X1 port map( I => n12756, ZN => n33097);
   U7903 : INV_X1 port map( I => n26709, ZN => n18606);
   U11889 : INV_X1 port map( I => n2158, ZN => n3417);
   U9302 : OAI21_X1 port map( A1 => n12373, A2 => n11696, B => n441, ZN => 
                           n6078);
   U9287 : NAND2_X1 port map( A1 => n948, A2 => n26696, ZN => n10340);
   U5898 : OAI21_X1 port map( A1 => n9147, A2 => n4946, B => n36873, ZN => 
                           n12936);
   U9239 : AOI21_X1 port map( A1 => n32633, A2 => n32634, B => n1492, ZN => 
                           n17143);
   U15746 : AOI21_X1 port map( A1 => n3283, A2 => n19449, B => n3282, ZN => 
                           n27283);
   U17875 : NAND2_X1 port map( A1 => n26650, A2 => n18719, ZN => n18718);
   U7269 : NAND2_X1 port map( A1 => n20636, A2 => n1090, ZN => n14757);
   U1762 : NOR2_X1 port map( A1 => n1232, A2 => n3606, ZN => n12714);
   U23458 : OAI21_X1 port map( A1 => n30363, A2 => n32669, B => n13392, ZN => 
                           n20792);
   U7288 : INV_X1 port map( I => n32926, ZN => n2660);
   U862 : OAI22_X1 port map( A1 => n32693, A2 => n34004, B1 => n8465, B2 => 
                           n1002, ZN => n35573);
   U2039 : NAND3_X1 port map( A1 => n26564, A2 => n17194, A3 => n26636, ZN => 
                           n26637);
   U4073 : NAND3_X1 port map( A1 => n26750, A2 => n17194, A3 => n15897, ZN => 
                           n15896);
   U890 : NAND2_X1 port map( A1 => n21182, A2 => n36445, ZN => n21050);
   U29844 : NOR2_X1 port map( A1 => n19529, A2 => n27508, ZN => n27420);
   U750 : INV_X1 port map( I => n27361, ZN => n27282);
   U4680 : INV_X1 port map( I => n17132, ZN => n13333);
   U21544 : INV_X1 port map( I => n36833, ZN => n30290);
   U484 : INV_X2 port map( I => n12485, ZN => n17142);
   U806 : BUF_X2 port map( I => n27361, Z => n32557);
   U19721 : INV_X1 port map( I => n39424, ZN => n35381);
   U17978 : INV_X2 port map( I => n11910, ZN => n20671);
   U4474 : INV_X1 port map( I => n7973, ZN => n1480);
   U24262 : INV_X2 port map( I => n34644, ZN => n27081);
   U3188 : INV_X1 port map( I => n35051, ZN => n11736);
   U793 : INV_X2 port map( I => n15360, ZN => n31298);
   U5880 : INV_X2 port map( I => n35500, ZN => n12326);
   U15027 : INV_X2 port map( I => n39826, ZN => n14327);
   U4153 : CLKBUF_X2 port map( I => n5363, Z => n11765);
   U5700 : INV_X1 port map( I => n3540, ZN => n995);
   U28310 : INV_X2 port map( I => n27448, ZN => n16043);
   U8081 : INV_X2 port map( I => n11729, ZN => n27180);
   U5891 : INV_X2 port map( I => n7632, ZN => n1000);
   U30562 : INV_X1 port map( I => n27358, ZN => n1227);
   U19112 : INV_X1 port map( I => n19135, ZN => n35299);
   U5381 : INV_X1 port map( I => n27365, ZN => n5772);
   U5581 : INV_X2 port map( I => n30358, ZN => n10946);
   U2881 : NAND2_X1 port map( A1 => n27415, A2 => n30434, ZN => n33234);
   U23988 : OAI21_X1 port map( A1 => n27372, A2 => n38578, B => n16042, ZN => 
                           n16041);
   U9157 : NAND3_X1 port map( A1 => n13294, A2 => n6534, A3 => n27240, ZN => 
                           n8263);
   U17558 : NOR2_X1 port map( A1 => n27341, A2 => n7096, ZN => n27342);
   U7782 : NAND2_X1 port map( A1 => n36528, A2 => n4192, ZN => n16849);
   U18665 : NAND2_X1 port map( A1 => n36989, A2 => n27379, ZN => n6446);
   U27384 : INV_X1 port map( I => n20740, ZN => n27147);
   U9706 : BUF_X2 port map( I => n19529, Z => n30768);
   U3576 : INV_X1 port map( I => n8537, ZN => n16263);
   U29390 : NAND2_X1 port map( A1 => n39414, A2 => n27240, ZN => n27238);
   U19794 : INV_X2 port map( I => n27269, ZN => n19662);
   U29382 : NAND2_X1 port map( A1 => n12326, A2 => n38060, ZN => n27206);
   U17192 : NAND2_X1 port map( A1 => n1225, A2 => n7096, ZN => n4037);
   U21123 : NOR3_X1 port map( A1 => n17467, A2 => n20574, A3 => n8627, ZN => 
                           n27092);
   U16275 : NAND2_X1 port map( A1 => n13526, A2 => n20377, ZN => n12375);
   U4654 : NAND2_X1 port map( A1 => n27108, A2 => n6686, ZN => n27181);
   U18865 : INV_X2 port map( I => n993, ZN => n33146);
   U18483 : NAND3_X1 port map( A1 => n1000, A2 => n31298, A3 => n27357, ZN => 
                           n15429);
   U6588 : INV_X1 port map( I => n20133, ZN => n9512);
   U479 : INV_X1 port map( I => n27424, ZN => n3059);
   U16313 : INV_X1 port map( I => n7975, ZN => n27247);
   U7344 : NAND2_X1 port map( A1 => n27275, A2 => n27314, ZN => n6648);
   U788 : INV_X1 port map( I => n18743, ZN => n7706);
   U507 : INV_X1 port map( I => n15616, ZN => n1080);
   U746 : INV_X1 port map( I => n4034, ZN => n1224);
   U18683 : INV_X1 port map( I => n39583, ZN => n1481);
   U18369 : NAND2_X1 port map( A1 => n6191, A2 => n27292, ZN => n27295);
   U728 : NOR2_X1 port map( A1 => n38578, A2 => n19662, ZN => n3470);
   U3486 : NAND2_X1 port map( A1 => n27251, A2 => n35184, ZN => n2377);
   U6143 : AOI21_X1 port map( A1 => n16170, A2 => n19997, B => n1477, ZN => 
                           n8640);
   U9182 : OAI21_X1 port map( A1 => n38630, A2 => n27409, B => n10677, ZN => 
                           n4570);
   U30226 : AOI21_X1 port map( A1 => n27250, A2 => n27007, B => n27027, ZN => 
                           n36806);
   U30081 : NOR3_X1 port map( A1 => n11765, A2 => n15276, A3 => n33893, ZN => 
                           n36761);
   U6155 : NAND3_X1 port map( A1 => n37653, A2 => n13278, A3 => n35485, ZN => 
                           n17500);
   U9191 : NOR2_X1 port map( A1 => n2761, A2 => n39826, ZN => n2580);
   U22453 : NAND2_X1 port map( A1 => n2035, A2 => n27402, ZN => n3978);
   U18444 : NOR2_X1 port map( A1 => n38926, A2 => n2923, ZN => n14634);
   U11604 : INV_X1 port map( I => n27299, ZN => n27377);
   U656 : NAND2_X1 port map( A1 => n27297, A2 => n27225, ZN => n31273);
   U686 : NOR2_X1 port map( A1 => n1475, A2 => n27269, ZN => n34990);
   U5743 : INV_X1 port map( I => n10032, ZN => n17903);
   U663 : INV_X1 port map( I => n27245, ZN => n33619);
   U24248 : NAND2_X1 port map( A1 => n14086, A2 => n8385, ZN => n14085);
   U799 : NAND2_X1 port map( A1 => n27398, A2 => n17142, ZN => n32631);
   U13451 : NAND3_X1 port map( A1 => n31150, A2 => n11140, A3 => n15360, ZN => 
                           n15120);
   U28843 : NAND2_X1 port map( A1 => n13178, A2 => n33403, ZN => n11591);
   U9148 : NOR2_X1 port map( A1 => n12074, A2 => n27090, ZN => n12073);
   U18648 : CLKBUF_X2 port map( I => n27407, Z => n7606);
   U2378 : NAND2_X1 port map( A1 => n31298, A2 => n34952, ZN => n27360);
   U14328 : NAND2_X1 port map( A1 => n16849, A2 => n16847, ZN => n16848);
   U29275 : NOR2_X1 port map( A1 => n37598, A2 => n36203, ZN => n26623);
   U30772 : BUF_X2 port map( I => n495, Z => n37001);
   U11529 : NOR2_X1 port map( A1 => n1220, A2 => n1797, ZN => n1796);
   U687 : NOR2_X1 port map( A1 => n17754, A2 => n945, ZN => n36120);
   U14209 : INV_X1 port map( I => n27408, ZN => n27155);
   U19128 : INV_X1 port map( I => n27347, ZN => n11682);
   U7347 : INV_X1 port map( I => n36989, ZN => n27072);
   U705 : OAI22_X1 port map( A1 => n4037, A2 => n8486, B1 => n27133, B2 => 
                           n1225, ZN => n36467);
   U14448 : NAND2_X1 port map( A1 => n15360, A2 => n27357, ZN => n2207);
   U721 : INV_X1 port map( I => n495, ZN => n27154);
   U9144 : AOI22_X1 port map( A1 => n30429, A2 => n11682, B1 => n993, B2 => 
                           n27348, ZN => n18075);
   U29365 : NAND3_X1 port map( A1 => n1486, A2 => n27196, A3 => n27364, ZN => 
                           n27122);
   U29405 : NAND3_X1 port map( A1 => n27371, A2 => n1475, A3 => n944, ZN => 
                           n27376);
   U2446 : AOI21_X1 port map( A1 => n1472, A2 => n27447, B => n32926, ZN => 
                           n1940);
   U6148 : AOI21_X1 port map( A1 => n8453, A2 => n27403, B => n35258, ZN => 
                           n15464);
   U434 : NAND3_X1 port map( A1 => n1217, A2 => n1224, A3 => n3513, ZN => 
                           n27382);
   U29375 : NAND3_X1 port map( A1 => n18246, A2 => n1085, A3 => n27416, ZN => 
                           n27182);
   U3111 : AOI21_X1 port map( A1 => n30851, A2 => n33254, B => n27081, ZN => 
                           n10337);
   U5773 : AOI22_X1 port map( A1 => n38146, A2 => n27403, B1 => n33803, B2 => 
                           n994, ZN => n32184);
   U24245 : AOI22_X1 port map( A1 => n36865, A2 => n27404, B1 => n27390, B2 => 
                           n13730, ZN => n2998);
   U6703 : OAI21_X1 port map( A1 => n27560, A2 => n1082, B => n10508, ZN => 
                           n27078);
   U16550 : NAND2_X1 port map( A1 => n35115, A2 => n35114, ZN => n35113);
   U1653 : NAND3_X1 port map( A1 => n37198, A2 => n39203, A3 => n27154, ZN => 
                           n27083);
   U21956 : NAND2_X1 port map( A1 => n10359, A2 => n13364, ZN => n10358);
   U11551 : NAND2_X1 port map( A1 => n27329, A2 => n27328, ZN => n21164);
   U628 : AOI21_X1 port map( A1 => n27245, A2 => n4192, B => n2006, ZN => n2114
                           );
   U4898 : NOR2_X1 port map( A1 => n34606, A2 => n4782, ZN => n8933);
   U18422 : NAND2_X1 port map( A1 => n17903, A2 => n27284, ZN => n17902);
   U22390 : NAND2_X1 port map( A1 => n16248, A2 => n4743, ZN => n35790);
   U21642 : NAND2_X1 port map( A1 => n27319, A2 => n37508, ZN => n9491);
   U9174 : OAI21_X1 port map( A1 => n18768, A2 => n2580, B => n27291, ZN => 
                           n18767);
   U1988 : NAND2_X1 port map( A1 => n10066, A2 => n18268, ZN => n19803);
   U25260 : NOR2_X1 port map( A1 => n1217, A2 => n27072, ZN => n19062);
   U11577 : NAND2_X1 port map( A1 => n37162, A2 => n7291, ZN => n20561);
   U14203 : OAI21_X1 port map( A1 => n27155, A2 => n5311, B => n37001, ZN => 
                           n3674);
   U4479 : AOI21_X1 port map( A1 => n27006, A2 => n7973, B => n32976, ZN => 
                           n5769);
   U15066 : NAND2_X1 port map( A1 => n34944, A2 => n34943, ZN => n35293);
   U4307 : NAND2_X1 port map( A1 => n33088, A2 => n31668, ZN => n27258);
   U20969 : NOR2_X1 port map( A1 => n7494, A2 => n39448, ZN => n13895);
   U2810 : NAND2_X1 port map( A1 => n36797, A2 => n19203, ZN => n35423);
   U392 : INV_X1 port map( I => n27852, ZN => n1458);
   U11506 : OAI21_X1 port map( A1 => n27065, A2 => n26273, B => n1221, ZN => 
                           n6027);
   U19471 : NAND3_X1 port map( A1 => n20740, A2 => n36234, A3 => n945, ZN => 
                           n27148);
   U11543 : NAND2_X1 port map( A1 => n7694, A2 => n17058, ZN => n10953);
   U22752 : NAND2_X1 port map( A1 => n37162, A2 => n38305, ZN => n10999);
   U3053 : INV_X1 port map( I => n37881, ZN => n4709);
   U3535 : INV_X1 port map( I => n27834, ZN => n32160);
   U25272 : OAI21_X1 port map( A1 => n14482, A2 => n15986, B => n17754, ZN => 
                           n15985);
   U381 : INV_X1 port map( I => n27554, ZN => n27853);
   U17733 : INV_X1 port map( I => n8894, ZN => n33595);
   U18800 : OAI21_X1 port map( A1 => n11486, A2 => n14667, B => n26196, ZN => 
                           n27794);
   U16663 : BUF_X2 port map( I => n19606, Z => n32931);
   U19263 : BUF_X2 port map( I => n10301, Z => n35318);
   U10104 : INV_X1 port map( I => n27464, ZN => n27669);
   U5835 : INV_X1 port map( I => n27672, ZN => n27849);
   U11447 : INV_X1 port map( I => n27756, ZN => n16972);
   U5810 : INV_X1 port map( I => n27760, ZN => n9162);
   U6697 : INV_X1 port map( I => n14260, ZN => n27676);
   U17329 : NAND2_X1 port map( A1 => n36639, A2 => n35603, ZN => n35178);
   U6696 : INV_X1 port map( I => n27607, ZN => n27460);
   U7750 : INV_X1 port map( I => n17417, ZN => n17418);
   U5829 : INV_X1 port map( I => n27830, ZN => n1456);
   U5524 : BUF_X2 port map( I => n28204, Z => n9514);
   U557 : INV_X2 port map( I => n10817, ZN => n7528);
   U12018 : INV_X1 port map( I => n34594, ZN => n12218);
   U5860 : INV_X1 port map( I => n759, ZN => n1441);
   U3907 : INV_X2 port map( I => n5352, ZN => n1442);
   U13947 : AOI21_X1 port map( A1 => n1212, A2 => n15357, B => n32783, ZN => 
                           n15204);
   U497 : INV_X2 port map( I => n19750, ZN => n1451);
   U24082 : INV_X1 port map( I => n13989, ZN => n15038);
   U343 : INV_X1 port map( I => n8148, ZN => n8149);
   U27296 : INV_X1 port map( I => n36463, ZN => n879);
   U340 : NOR2_X1 port map( A1 => n1202, A2 => n15704, ZN => n10779);
   U19758 : NOR2_X1 port map( A1 => n1209, A2 => n8078, ZN => n11737);
   U2914 : NAND2_X1 port map( A1 => n1439, A2 => n28205, ZN => n16261);
   U4134 : INV_X1 port map( I => n17314, ZN => n28102);
   U21722 : BUF_X2 port map( I => n28237, Z => n32352);
   U6648 : INV_X1 port map( I => n877, ZN => n28156);
   U26373 : INV_X2 port map( I => n28279, ZN => n1076);
   U543 : INV_X1 port map( I => n12673, ZN => n5020);
   U9665 : AND2_X1 port map( A1 => n34166, A2 => n35225, Z => n28064);
   U29356 : INV_X1 port map( I => n27481, ZN => n28050);
   U6650 : INV_X1 port map( I => n7528, ZN => n27980);
   U23243 : INV_X1 port map( I => n32638, ZN => n13081);
   U593 : INV_X1 port map( I => n28133, ZN => n28015);
   U28028 : NOR2_X1 port map( A1 => n33603, A2 => n879, ZN => n20941);
   U6644 : NAND3_X1 port map( A1 => n18673, A2 => n13769, A3 => n15704, ZN => 
                           n7717);
   U584 : NAND2_X1 port map( A1 => n19410, A2 => n19667, ZN => n345);
   U461 : NAND2_X1 port map( A1 => n20053, A2 => n15925, ZN => n27940);
   U514 : NOR2_X1 port map( A1 => n4915, A2 => n2717, ZN => n36818);
   U334 : INV_X1 port map( I => n878, ZN => n28001);
   U515 : INV_X1 port map( I => n12038, ZN => n32728);
   U7467 : AOI21_X1 port map( A1 => n12784, A2 => n28283, B => n16544, ZN => 
                           n30565);
   U2678 : BUF_X2 port map( I => n18261, Z => n42);
   U522 : NOR2_X1 port map( A1 => n983, A2 => n10836, ZN => n10519);
   U572 : CLKBUF_X2 port map( I => n5352, Z => n35607);
   U2333 : BUF_X2 port map( I => n15692, Z => n9897);
   U6677 : NOR2_X1 port map( A1 => n883, A2 => n20860, ZN => n20977);
   U510 : INV_X2 port map( I => n28024, ZN => n33331);
   U17028 : INV_X2 port map( I => n8818, ZN => n28109);
   U20871 : INV_X2 port map( I => n27894, ZN => n28165);
   U2501 : INV_X1 port map( I => n9534, ZN => n11754);
   U15417 : OR2_X1 port map( A1 => n15922, A2 => n28159, Z => n11501);
   U8017 : AND2_X1 port map( A1 => n19891, A2 => n19605, Z => n34170);
   U11342 : AND2_X1 port map( A1 => n20010, A2 => n19995, Z => n15623);
   U549 : INV_X1 port map( I => n37056, ZN => n28151);
   U9111 : INV_X1 port map( I => n28157, ZN => n28012);
   U322 : INV_X1 port map( I => n886, ZN => n1205);
   U7713 : INV_X2 port map( I => n18261, ZN => n1444);
   U6684 : INV_X1 port map( I => n14451, ZN => n28230);
   U15061 : INV_X2 port map( I => n5988, ZN => n7690);
   U18125 : INV_X2 port map( I => n2716, ZN => n1440);
   U3455 : OAI21_X1 port map( A1 => n1070, A2 => n28215, B => n1448, ZN => 
                           n28081);
   U20416 : NAND3_X1 port map( A1 => n8232, A2 => n28229, A3 => n28228, ZN => 
                           n19921);
   U9755 : NAND2_X1 port map( A1 => n3983, A2 => n30773, ZN => n15622);
   U20545 : NAND2_X1 port map( A1 => n3032, A2 => n3159, ZN => n35507);
   U16253 : AOI21_X1 port map( A1 => n11375, A2 => n32080, B => n28159, ZN => 
                           n5671);
   U3665 : NOR2_X1 port map( A1 => n37057, A2 => n988, ZN => n13469);
   U13223 : INV_X1 port map( I => n889, ZN => n7310);
   U27952 : AOI21_X1 port map( A1 => n11754, A2 => n27948, B => n33331, ZN => 
                           n10352);
   U30038 : INV_X1 port map( I => n28043, ZN => n2664);
   U26487 : NAND2_X1 port map( A1 => n18603, A2 => n15357, ZN => n15518);
   U3216 : NOR2_X1 port map( A1 => n11628, A2 => n28272, ZN => n13776);
   U11331 : NAND2_X1 port map( A1 => n18392, A2 => n12260, ZN => n12258);
   U25824 : NAND2_X1 port map( A1 => n36818, A2 => n36817, ZN => n16034);
   U11360 : INV_X2 port map( I => n1074, ZN => n19124);
   U3931 : NAND2_X1 port map( A1 => n19366, A2 => n99, ZN => n28053);
   U27193 : NOR2_X1 port map( A1 => n1207, A2 => n28290, ZN => n28291);
   U7729 : INV_X1 port map( I => n9089, ZN => n21020);
   U9058 : OAI21_X1 port map( A1 => n6050, A2 => n5239, B => n35607, ZN => 
                           n13695);
   U7702 : INV_X1 port map( I => n30484, ZN => n1435);
   U30818 : INV_X1 port map( I => n8604, ZN => n28266);
   U6135 : INV_X1 port map( I => n38579, ZN => n28217);
   U501 : INV_X1 port map( I => n1454, ZN => n1073);
   U14558 : NOR2_X1 port map( A1 => n9969, A2 => n28189, ZN => n28190);
   U482 : NAND2_X1 port map( A1 => n28215, A2 => n987, ZN => n16971);
   U4338 : NOR2_X1 port map( A1 => n38996, A2 => n14562, ZN => n31765);
   U11271 : NOR2_X1 port map( A1 => n28032, A2 => n4347, ZN => n6114);
   U7622 : NAND3_X1 port map( A1 => n9534, A2 => n27948, A3 => n28024, ZN => 
                           n18149);
   U463 : NAND2_X1 port map( A1 => n21239, A2 => n27896, ZN => n31848);
   U6131 : INV_X1 port map( I => n20977, ZN => n28216);
   U9027 : AOI21_X1 port map( A1 => n9702, A2 => n18841, B => n1069, ZN => 
                           n27711);
   U7394 : NOR2_X1 port map( A1 => n15014, A2 => n27955, ZN => n10052);
   U29492 : NAND2_X1 port map( A1 => n1200, A2 => n19124, ZN => n27872);
   U16785 : NOR2_X1 port map( A1 => n1446, A2 => n4306, ZN => n28242);
   U3376 : NAND2_X1 port map( A1 => n14397, A2 => n28181, ZN => n19123);
   U29560 : NAND3_X1 port map( A1 => n28171, A2 => n19601, A3 => n28260, ZN => 
                           n28173);
   U400 : OAI21_X1 port map( A1 => n14562, A2 => n1454, B => n1206, ZN => n3230
                           );
   U6660 : OAI21_X1 port map( A1 => n1202, A2 => n38666, B => n11737, ZN => 
                           n9237);
   U19708 : OAI21_X1 port map( A1 => n31616, A2 => n33292, B => n31607, ZN => 
                           n13455);
   U11206 : NOR2_X1 port map( A1 => n28227, A2 => n19891, ZN => n20225);
   U2376 : NAND2_X1 port map( A1 => n27900, A2 => n11461, ZN => n28203);
   U14904 : NAND2_X1 port map( A1 => n7635, A2 => n31022, ZN => n28085);
   U5895 : NAND2_X1 port map( A1 => n17770, A2 => n7851, ZN => n16994);
   U11170 : NOR2_X1 port map( A1 => n4415, A2 => n3832, ZN => n2667);
   U9036 : OAI21_X1 port map( A1 => n6245, A2 => n7223, B => n38762, ZN => 
                           n6244);
   U29476 : NOR2_X1 port map( A1 => n36689, A2 => n6693, ZN => n6243);
   U24491 : NAND2_X1 port map( A1 => n15572, A2 => n15571, ZN => n15570);
   U26253 : NOR2_X1 port map( A1 => n31607, A2 => n28114, ZN => n15993);
   U2683 : NAND2_X1 port map( A1 => n28274, A2 => n37057, ZN => n33867);
   U339 : INV_X2 port map( I => n37671, ZN => n3235);
   U17395 : AND2_X1 port map( A1 => n11368, A2 => n28286, Z => n31871);
   U18268 : NAND2_X1 port map( A1 => n28661, A2 => n28660, ZN => n6041);
   U296 : NAND3_X1 port map( A1 => n1451, A2 => n27962, A3 => n10254, ZN => 
                           n11893);
   U7668 : AOI21_X1 port map( A1 => n15249, A2 => n42, B => n28111, ZN => 
                           n11518);
   U19497 : OAI22_X1 port map( A1 => n27918, A2 => n200, B1 => n7635, B2 => 
                           n6777, ZN => n20533);
   U6129 : INV_X1 port map( I => n16261, ZN => n7541);
   U5923 : NAND2_X1 port map( A1 => n28284, A2 => n28283, ZN => n11323);
   U29384 : NAND2_X1 port map( A1 => n38579, A2 => n28079, ZN => n28351);
   U18987 : NAND2_X1 port map( A1 => n7555, A2 => n28458, ZN => n31854);
   U28497 : NOR2_X1 port map( A1 => n14615, A2 => n36591, ZN => n16964);
   U353 : OAI21_X1 port map( A1 => n28168, A2 => n20398, B => n30995, ZN => 
                           n11322);
   U1992 : AOI21_X1 port map( A1 => n27920, A2 => n1070, B => n987, ZN => 
                           n27921);
   U22881 : AOI21_X1 port map( A1 => n33669, A2 => n32705, B => n35862, ZN => 
                           n17476);
   U9023 : AOI21_X1 port map( A1 => n28243, A2 => n1444, B => n28242, ZN => 
                           n28244);
   U3197 : NAND2_X1 port map( A1 => n6117, A2 => n8149, ZN => n6116);
   U28075 : OAI21_X1 port map( A1 => n36559, A2 => n36558, B => n3990, ZN => 
                           n28263);
   U17455 : NAND2_X1 port map( A1 => n7719, A2 => n1072, ZN => n7718);
   U29512 : NAND2_X1 port map( A1 => n27935, A2 => n28142, ZN => n28346);
   U3059 : NAND2_X1 port map( A1 => n12227, A2 => n33048, ZN => n28087);
   U17250 : BUF_X2 port map( I => n19675, Z => n16777);
   U4600 : INV_X1 port map( I => n3664, ZN => n28657);
   U10584 : INV_X1 port map( I => n1823, ZN => n31855);
   U328 : OAI21_X1 port map( A1 => n28660, A2 => n1431, B => n6041, ZN => n6040
                           );
   U22893 : INV_X2 port map( I => n1195, ZN => n28812);
   U7492 : NOR2_X1 port map( A1 => n3252, A2 => n28369, ZN => n13820);
   U23003 : INV_X1 port map( I => n28661, ZN => n28553);
   U387 : NAND2_X1 port map( A1 => n2822, A2 => n89, ZN => n36986);
   U29630 : NAND2_X1 port map( A1 => n16778, A2 => n16777, ZN => n12653);
   U14405 : NAND2_X1 port map( A1 => n31597, A2 => n14760, ZN => n15024);
   U17068 : NAND2_X1 port map( A1 => n11005, A2 => n11006, ZN => n31542);
   U1605 : INV_X2 port map( I => n2191, ZN => n1419);
   U424 : INV_X2 port map( I => n37758, ZN => n28554);
   U16637 : CLKBUF_X2 port map( I => n16067, Z => n32543);
   U6124 : INV_X1 port map( I => n8476, ZN => n28690);
   U11158 : OR2_X1 port map( A1 => n496, A2 => n14193, Z => n16398);
   U12547 : INV_X1 port map( I => n20445, ZN => n1434);
   U23536 : INV_X2 port map( I => n28677, ZN => n18883);
   U3620 : INV_X1 port map( I => n9290, ZN => n9329);
   U6611 : INV_X1 port map( I => n28728, ZN => n28323);
   U15324 : INV_X1 port map( I => n3538, ZN => n14987);
   U5123 : INV_X2 port map( I => n6405, ZN => n28378);
   U2443 : NOR2_X1 port map( A1 => n28724, A2 => n37311, ZN => n20736);
   U11085 : INV_X1 port map( I => n15024, ZN => n12715);
   U10699 : NOR2_X1 port map( A1 => n28727, A2 => n15752, ZN => n34433);
   U11001 : NAND2_X1 port map( A1 => n3252, A2 => n38556, ZN => n3250);
   U7577 : NAND2_X1 port map( A1 => n974, A2 => n28339, ZN => n12539);
   U18307 : NAND3_X1 port map( A1 => n36775, A2 => n38669, A3 => n36774, ZN => 
                           n36773);
   U19673 : NAND2_X1 port map( A1 => n32791, A2 => n28753, ZN => n12313);
   U194 : OAI21_X1 port map( A1 => n28697, A2 => n9648, B => n10587, ZN => 
                           n16495);
   U11011 : NOR2_X1 port map( A1 => n14605, A2 => n28654, ZN => n11800);
   U16960 : NOR2_X1 port map( A1 => n2330, A2 => n33436, ZN => n33640);
   U309 : INV_X1 port map( I => n6067, ZN => n33046);
   U420 : INV_X2 port map( I => n33047, ZN => n28639);
   U1817 : INV_X2 port map( I => n11164, ZN => n9444);
   U224 : NAND2_X1 port map( A1 => n14621, A2 => n11697, ZN => n28444);
   U6609 : INV_X2 port map( I => n6892, ZN => n28530);
   U6623 : INV_X1 port map( I => n15224, ZN => n1192);
   U24550 : INV_X1 port map( I => n28434, ZN => n28380);
   U211 : INV_X2 port map( I => n13690, ZN => n18871);
   U23547 : INV_X1 port map( I => n9575, ZN => n20494);
   U5598 : INV_X1 port map( I => n19759, ZN => n28808);
   U6112 : INV_X1 port map( I => n11831, ZN => n1066);
   U7572 : INV_X1 port map( I => n31015, ZN => n28312);
   U16872 : NAND2_X1 port map( A1 => n1194, A2 => n28659, ZN => n28555);
   U7522 : OAI21_X1 port map( A1 => n28732, A2 => n17073, B => n32595, ZN => 
                           n13784);
   U26291 : NAND3_X1 port map( A1 => n15112, A2 => n31321, A3 => n28717, ZN => 
                           n28709);
   U19535 : NAND2_X1 port map( A1 => n35777, A2 => n902, ZN => n18088);
   U11089 : NAND2_X1 port map( A1 => n13061, A2 => n8349, ZN => n13060);
   U9101 : NOR2_X1 port map( A1 => n36892, A2 => n13891, ZN => n31206);
   U2375 : NOR2_X1 port map( A1 => n28765, A2 => n28812, ZN => n13964);
   U27381 : NAND2_X1 port map( A1 => n1426, A2 => n39363, ZN => n18859);
   U27004 : NOR2_X1 port map( A1 => n10618, A2 => n17771, ZN => n18096);
   U17230 : NAND3_X1 port map( A1 => n18281, A2 => n36775, A3 => n37863, ZN => 
                           n8320);
   U16199 : OAI22_X1 port map( A1 => n28554, A2 => n28551, B1 => n28427, B2 => 
                           n1431, ZN => n28428);
   U15567 : INV_X1 port map( I => n36685, ZN => n28415);
   U2583 : INV_X1 port map( I => n18960, ZN => n28450);
   U8947 : NOR2_X1 port map( A1 => n12539, A2 => n11488, ZN => n12538);
   U22568 : INV_X1 port map( I => n32338, ZN => n35804);
   U13367 : INV_X1 port map( I => n39435, ZN => n34737);
   U7519 : NAND2_X1 port map( A1 => n16255, A2 => n16295, ZN => n16256);
   U12528 : AOI21_X1 port map( A1 => n8637, A2 => n12336, B => n34559, ZN => 
                           n34627);
   U5444 : INV_X1 port map( I => n18972, ZN => n36145);
   U8841 : NAND2_X1 port map( A1 => n32376, A2 => n14222, ZN => n16657);
   U7508 : NAND2_X1 port map( A1 => n33100, A2 => n978, ZN => n15457);
   U6575 : NAND2_X1 port map( A1 => n14816, A2 => n14604, ZN => n21145);
   U185 : INV_X2 port map( I => n28530, ZN => n11390);
   U284 : BUF_X2 port map( I => n28638, Z => n4369);
   U305 : NAND2_X1 port map( A1 => n33436, A2 => n1431, ZN => n28439);
   U2817 : NOR2_X1 port map( A1 => n3598, A2 => n18883, ZN => n32952);
   U18767 : AND2_X1 port map( A1 => n28478, A2 => n1414, Z => n28309);
   U5417 : NAND2_X1 port map( A1 => n7486, A2 => n38231, ZN => n34958);
   U30542 : NOR2_X1 port map( A1 => n11438, A2 => n11490, ZN => n33910);
   U17096 : NAND2_X1 port map( A1 => n28494, A2 => n1434, ZN => n12890);
   U7528 : NOR2_X1 port map( A1 => n28530, A2 => n12237, ZN => n10910);
   U19623 : NAND2_X1 port map( A1 => n18972, A2 => n30931, ZN => n28489);
   U23221 : NAND2_X1 port map( A1 => n32703, A2 => n15580, ZN => n14506);
   U3465 : OAI21_X1 port map( A1 => n4969, A2 => n28510, B => n28715, ZN => 
                           n7799);
   U13605 : OAI21_X1 port map( A1 => n888, A2 => n28293, B => n32286, ZN => 
                           n15514);
   U19563 : NAND3_X1 port map( A1 => n10587, A2 => n9598, A3 => n37081, ZN => 
                           n28520);
   U27412 : NAND2_X1 port map( A1 => n34244, A2 => n9917, ZN => n28522);
   U1705 : OAI21_X1 port map( A1 => n28386, A2 => n4950, B => n4949, ZN => 
                           n27958);
   U1812 : NAND2_X1 port map( A1 => n28754, A2 => n28755, ZN => n16922);
   U1700 : OAI21_X1 port map( A1 => n28368, A2 => n18972, B => n28490, ZN => 
                           n9625);
   U11043 : NAND2_X1 port map( A1 => n28293, A2 => n28771, ZN => n11465);
   U2832 : OAI21_X1 port map( A1 => n27457, A2 => n28535, B => n28537, ZN => 
                           n3129);
   U5991 : NAND2_X1 port map( A1 => n28756, A2 => n21027, ZN => n21026);
   U25310 : OAI21_X1 port map( A1 => n37758, A2 => n33436, B => n19688, ZN => 
                           n28558);
   U10926 : NAND2_X1 port map( A1 => n28343, A2 => n34007, ZN => n11664);
   U9282 : AOI21_X1 port map( A1 => n38556, A2 => n28604, B => n34298, ZN => 
                           n35621);
   U258 : AOI21_X1 port map( A1 => n28617, A2 => n3664, B => n28654, ZN => 
                           n28618);
   U11039 : OAI21_X1 port map( A1 => n9638, A2 => n28348, B => n9141, ZN => 
                           n16932);
   U16555 : OAI22_X1 port map( A1 => n5399, A2 => n5396, B1 => n9586, B2 => 
                           n38203, ZN => n5398);
   U7504 : OAI21_X1 port map( A1 => n11438, A2 => n7913, B => n11490, ZN => 
                           n8854);
   U6591 : NOR2_X1 port map( A1 => n20497, A2 => n1823, ZN => n20493);
   U6105 : NAND3_X1 port map( A1 => n12990, A2 => n28453, A3 => n37204, ZN => 
                           n12378);
   U4056 : CLKBUF_X2 port map( I => n11695, Z => n3703);
   U8935 : OR2_X1 port map( A1 => n28529, A2 => n37619, Z => n11491);
   U29616 : NOR2_X1 port map( A1 => n36777, A2 => n28516, ZN => n28518);
   U8940 : AOI22_X1 port map( A1 => n12605, A2 => n28608, B1 => n11390, B2 => 
                           n33647, ZN => n6094);
   U4645 : OAI21_X1 port map( A1 => n8323, A2 => n8322, B => n7555, ZN => n8321
                           );
   U5406 : CLKBUF_X2 port map( I => n7744, Z => n32448);
   U20153 : CLKBUF_X2 port map( I => n29160, Z => n33511);
   U12735 : INV_X1 port map( I => n10079, ZN => n29127);
   U16185 : AOI21_X1 port map( A1 => n28808, A2 => n33577, B => n35083, ZN => 
                           n35082);
   U24689 : INV_X1 port map( I => n28874, ZN => n16310);
   U16688 : INV_X1 port map( I => n9787, ZN => n21007);
   U16761 : BUF_X2 port map( I => n20465, Z => n2392);
   U12189 : BUF_X2 port map( I => n9036, Z => n3665);
   U10970 : INV_X1 port map( I => n10080, ZN => n28927);
   U15141 : INV_X1 port map( I => n14941, ZN => n28977);
   U209 : INV_X1 port map( I => n28827, ZN => n28978);
   U14654 : INV_X2 port map( I => n20686, ZN => n29862);
   U3894 : INV_X2 port map( I => n10896, ZN => n19962);
   U15637 : INV_X1 port map( I => n6163, ZN => n31428);
   U3162 : INV_X2 port map( I => n21270, ZN => n13441);
   U10903 : CLKBUF_X2 port map( I => n29424, Z => n19896);
   U15438 : BUF_X2 port map( I => n28436, Z => n29700);
   U27831 : INV_X2 port map( I => n19424, ZN => n1407);
   U15667 : INV_X1 port map( I => n32251, ZN => n29195);
   U138 : INV_X2 port map( I => n18315, ZN => n29595);
   U30866 : INV_X1 port map( I => n12829, ZN => n31279);
   U189 : INV_X1 port map( I => n20026, ZN => n29310);
   U14084 : INV_X1 port map( I => n18288, ZN => n30195);
   U18048 : INV_X1 port map( I => n14254, ZN => n17238);
   U7442 : NAND2_X1 port map( A1 => n1179, A2 => n18720, ZN => n4655);
   U30865 : INV_X1 port map( I => n18667, ZN => n33928);
   U3505 : INV_X1 port map( I => n29701, ZN => n8941);
   U5081 : INV_X2 port map( I => n30043, ZN => n1056);
   U4102 : OR2_X1 port map( A1 => n30049, A2 => n33256, Z => n4255);
   U19400 : INV_X1 port map( I => n16217, ZN => n29935);
   U8853 : INV_X2 port map( I => n20979, ZN => n30680);
   U4963 : INV_X1 port map( I => n15854, ZN => n29996);
   U30098 : NAND2_X1 port map( A1 => n6019, A2 => n1057, ZN => n29986);
   U6555 : INV_X2 port map( I => n30220, ZN => n1177);
   U18092 : INV_X1 port map( I => n16599, ZN => n20982);
   U8079 : INV_X2 port map( I => n34000, ZN => n29779);
   U180 : OR2_X1 port map( A1 => n33256, A2 => n11896, Z => n30048);
   U1576 : INV_X1 port map( I => n20687, ZN => n29863);
   U127 : INV_X1 port map( I => n11428, ZN => n30162);
   U156 : INV_X1 port map( I => n33967, ZN => n29445);
   U94 : INV_X1 port map( I => n21023, ZN => n17644);
   U10035 : NOR2_X1 port map( A1 => n20525, A2 => n30153, ZN => n30796);
   U23169 : INV_X1 port map( I => n11783, ZN => n30241);
   U74 : INV_X2 port map( I => n29596, ZN => n12450);
   U16855 : NAND2_X1 port map( A1 => n3700, A2 => n3631, ZN => n3698);
   U27617 : NOR2_X1 port map( A1 => n30048, A2 => n32628, ZN => n19454);
   U9831 : INV_X1 port map( I => n34344, ZN => n18007);
   U4808 : NOR2_X1 port map( A1 => n32945, A2 => n13153, ZN => n32944);
   U25496 : INV_X1 port map( I => n29586, ZN => n21264);
   U2753 : NAND2_X1 port map( A1 => n9394, A2 => n15153, ZN => n14495);
   U23797 : NAND2_X1 port map( A1 => n16510, A2 => n971, ZN => n13085);
   U3284 : INV_X1 port map( I => n20982, ZN => n1398);
   U10835 : NOR2_X1 port map( A1 => n30187, A2 => n39280, ZN => n29061);
   U7483 : NAND2_X1 port map( A1 => n29777, A2 => n33964, ZN => n29780);
   U87 : INV_X2 port map( I => n6019, ZN => n29987);
   U8856 : AOI21_X1 port map( A1 => n771, A2 => n29446, B => n1401, ZN => 
                           n16508);
   U2816 : AOI21_X1 port map( A1 => n29378, A2 => n29458, B => n29377, ZN => 
                           n29345);
   U7413 : AOI21_X1 port map( A1 => n5570, A2 => n921, B => n3700, ZN => n9799)
                           ;
   U8875 : INV_X1 port map( I => n1399, ZN => n11574);
   U120 : INV_X1 port map( I => n21285, ZN => n21287);
   U7399 : NOR2_X1 port map( A1 => n28864, A2 => n29587, ZN => n13670);
   U29771 : INV_X1 port map( I => n32906, ZN => n29266);
   U15054 : NOR2_X1 port map( A1 => n29348, A2 => n29286, ZN => n29211);
   U116 : INV_X1 port map( I => n20018, ZN => n11056);
   U4964 : NAND2_X1 port map( A1 => n29946, A2 => n32571, ZN => n19137);
   U5374 : OR2_X1 port map( A1 => n29701, A2 => n16599, Z => n34180);
   U10861 : AND2_X1 port map( A1 => n21023, A2 => n28843, Z => n29634);
   U142 : INV_X1 port map( I => n29941, ZN => n30051);
   U5584 : INV_X1 port map( I => n344, ZN => n16209);
   U5587 : INV_X2 port map( I => n32946, ZN => n907);
   U111 : NOR2_X1 port map( A1 => n1181, A2 => n30160, ZN => n35849);
   U6526 : NOR2_X1 port map( A1 => n2456, A2 => n19992, ZN => n2016);
   U3536 : NOR2_X1 port map( A1 => n29449, A2 => n771, ZN => n29350);
   U7400 : NAND2_X1 port map( A1 => n16074, A2 => n14151, ZN => n2132);
   U7388 : NOR2_X1 port map( A1 => n13670, A2 => n13672, ZN => n13669);
   U2459 : NOR2_X1 port map( A1 => n1404, A2 => n29595, ZN => n2378);
   U29679 : NAND2_X1 port map( A1 => n30159, A2 => n1399, ZN => n33488);
   U10754 : OAI21_X1 port map( A1 => n14755, A2 => n12054, B => n38262, ZN => 
                           n12060);
   U16558 : INV_X1 port map( I => n32894, ZN => n30045);
   U30336 : AOI21_X1 port map( A1 => n29694, A2 => n21037, B => n2559, ZN => 
                           n33760);
   U14473 : NAND2_X1 port map( A1 => n33094, A2 => n34858, ZN => n30396);
   U3084 : NAND2_X1 port map( A1 => n33277, A2 => n1400, ZN => n7908);
   U2418 : OAI21_X1 port map( A1 => n29634, A2 => n29704, B => n16209, ZN => 
                           n17348);
   U93 : NAND2_X1 port map( A1 => n36207, A2 => n1755, ZN => n33393);
   U3540 : NOR2_X1 port map( A1 => n29449, A2 => n1176, ZN => n19791);
   U10808 : OAI21_X1 port map( A1 => n2121, A2 => n18815, B => n19508, ZN => 
                           n3245);
   U27258 : OAI21_X1 port map( A1 => n29843, A2 => n773, B => n18477, ZN => 
                           n29873);
   U67 : NOR2_X1 port map( A1 => n33394, A2 => n33393, ZN => n18590);
   U77 : NOR2_X1 port map( A1 => n34973, A2 => n29378, ZN => n35295);
   U75 : NAND2_X1 port map( A1 => n36023, A2 => n36022, ZN => n4799);
   U18838 : INV_X1 port map( I => n6332, ZN => n10869);
   U16296 : AOI21_X1 port map( A1 => n17842, A2 => n39416, B => n14183, ZN => 
                           n35096);
   U17289 : INV_X1 port map( I => n9828, ZN => n14126);
   U72 : INV_X1 port map( I => n20208, ZN => n29534);
   U26258 : INV_X2 port map( I => n18081, ZN => n1174);
   U4068 : INV_X1 port map( I => n29277, ZN => n1379);
   U46 : INV_X2 port map( I => n9105, ZN => n969);
   U26874 : INV_X1 port map( I => n29659, ZN => n17382);
   U9482 : INV_X1 port map( I => n29930, ZN => n29922);
   U5567 : CLKBUF_X2 port map( I => n29475, Z => n18873);
   U2906 : CLKBUF_X2 port map( I => n30079, Z => n31120);
   U2890 : INV_X1 port map( I => n17469, ZN => n30129);
   U3016 : INV_X1 port map( I => n29979, ZN => n29975);
   U23831 : INV_X1 port map( I => n29208, ZN => n13142);
   U61 : INV_X1 port map( I => n29367, ZN => n16683);
   U6126 : INV_X1 port map( I => n30262, ZN => n1172);
   U49 : NOR2_X1 port map( A1 => n28585, A2 => n28584, ZN => n17262);
   U4040 : INV_X1 port map( I => n29684, ZN => n29675);
   U18806 : NAND2_X1 port map( A1 => n31821, A2 => n10978, ZN => n30134);
   U41 : INV_X1 port map( I => n20078, ZN => n30069);
   U6066 : INV_X1 port map( I => n20307, ZN => n30132);
   U55 : AND2_X1 port map( A1 => n31821, A2 => n10978, Z => n34177);
   U29921 : INV_X1 port map( I => n33437, ZN => n36738);
   U5831 : INV_X1 port map( I => n29929, ZN => n3860);
   U23 : INV_X1 port map( I => n30022, ZN => n30035);
   U17382 : NAND2_X1 port map( A1 => n38164, A2 => n17192, ZN => n33207);
   U2186 : NAND2_X1 port map( A1 => n29478, A2 => n29468, ZN => n29464);
   U7363 : INV_X1 port map( I => n29981, ZN => n29977);
   U30801 : INV_X1 port map( I => n30107, ZN => n30119);
   U14 : INV_X1 port map( I => n13192, ZN => n29811);
   U3836 : INV_X1 port map( I => n15509, ZN => n29209);
   U3577 : NAND2_X1 port map( A1 => n30038, A2 => n9231, ZN => n30014);
   U47 : INV_X2 port map( I => n29859, ZN => n29851);
   U17211 : NOR2_X1 port map( A1 => n1385, A2 => n32508, ZN => n8286);
   U2919 : NAND2_X1 port map( A1 => n29567, A2 => n31899, ZN => n29565);
   U7371 : INV_X1 port map( I => n29530, ZN => n29527);
   U17564 : INV_X1 port map( I => n29740, ZN => n19348);
   U7370 : INV_X1 port map( I => n30093, ZN => n30098);
   U19739 : INV_X1 port map( I => n37096, ZN => n29369);
   U18 : INV_X1 port map( I => n17192, ZN => n17193);
   U20893 : NAND2_X1 port map( A1 => n10813, A2 => n8286, ZN => n9261);
   U2 : NAND3_X1 port map( A1 => n29368, A2 => n13839, A3 => n13804, ZN => 
                           n39677);
   U6 : AOI22_X1 port map( A1 => n19090, A2 => n5530, B1 => n29277, B2 => 
                           n37157, ZN => n17773);
   U7 : AND2_X1 port map( A1 => n4368, A2 => n12198, Z => n4367);
   U8 : NOR2_X1 port map( A1 => n20538, A2 => n4368, ZN => n30171);
   U10 : INV_X1 port map( I => n29336, ZN => n29335);
   U11 : NAND2_X1 port map( A1 => n2792, A2 => n29802, ZN => n29806);
   U15 : NAND2_X1 port map( A1 => n10118, A2 => n30117, ZN => n30106);
   U20 : BUF_X2 port map( I => n3096, Z => n36096);
   U21 : INV_X1 port map( I => n29231, ZN => n1387);
   U22 : INV_X1 port map( I => n29802, ZN => n29813);
   U24 : AND2_X1 port map( A1 => n30097, A2 => n31601, Z => n16471);
   U26 : NAND2_X1 port map( A1 => n35272, A2 => n16260, ZN => n15044);
   U30 : INV_X1 port map( I => n85, ZN => n9913);
   U33 : INV_X1 port map( I => n29678, ZN => n1173);
   U34 : INV_X2 port map( I => n12198, ZN => n20538);
   U36 : INV_X2 port map( I => n20274, ZN => n10813);
   U38 : INV_X1 port map( I => n30213, ZN => n33521);
   U45 : INV_X1 port map( I => n31899, ZN => n1053);
   U48 : NOR2_X1 port map( A1 => n38164, A2 => n1385, ZN => n37724);
   U52 : NAND2_X1 port map( A1 => n29810, A2 => n13192, ZN => n5970);
   U54 : OR2_X1 port map( A1 => n19475, A2 => n20160, Z => n37157);
   U56 : NAND2_X1 port map( A1 => n4072, A2 => n33071, ZN => n33070);
   U57 : INV_X2 port map( I => n8039, ZN => n30034);
   U58 : AOI22_X1 port map( A1 => n29595, A2 => n2296, B1 => n31667, B2 => 
                           n14417, ZN => n36193);
   U62 : NAND2_X1 port map( A1 => n29427, A2 => n29449, ZN => n38805);
   U66 : AOI21_X1 port map( A1 => n30165, A2 => n30046, B => n39416, ZN => 
                           n36023);
   U69 : OAI21_X1 port map( A1 => n7207, A2 => n39322, B => n19162, ZN => 
                           n20160);
   U70 : AND2_X1 port map( A1 => n29942, A2 => n30059, Z => n37177);
   U71 : OAI21_X1 port map( A1 => n29485, A2 => n19962, B => n32197, ZN => 
                           n29489);
   U76 : NAND2_X1 port map( A1 => n37752, A2 => n20673, ZN => n5924);
   U83 : NAND2_X1 port map( A1 => n37376, A2 => n37614, ZN => n37375);
   U84 : NAND2_X1 port map( A1 => n16508, A2 => n32671, ZN => n37797);
   U85 : OAI21_X1 port map( A1 => n38919, A2 => n6938, B => n29202, ZN => 
                           n38773);
   U86 : OAI21_X1 port map( A1 => n20289, A2 => n29635, B => n18107, ZN => 
                           n35762);
   U89 : NAND2_X1 port map( A1 => n2954, A2 => n29459, ZN => n34194);
   U99 : OAI22_X1 port map( A1 => n29457, A2 => n31521, B1 => n13261, B2 => 
                           n29458, ZN => n8924);
   U102 : AOI22_X1 port map( A1 => n29939, A2 => n6019, B1 => n29987, B2 => 
                           n30051, ZN => n34681);
   U103 : AND2_X1 port map( A1 => n5348, A2 => n20080, Z => n29899);
   U107 : INV_X1 port map( I => n773, ZN => n29867);
   U110 : INV_X1 port map( I => n28882, ZN => n8762);
   U113 : NAND2_X1 port map( A1 => n16672, A2 => n1755, ZN => n31065);
   U122 : CLKBUF_X2 port map( I => n29454, Z => n39647);
   U123 : OR2_X1 port map( A1 => n1056, A2 => n4220, Z => n37082);
   U124 : CLKBUF_X4 port map( I => n4879, Z => n37936);
   U125 : OAI21_X1 port map( A1 => n37729, A2 => n37728, B => n37727, ZN => 
                           n29011);
   U129 : NOR2_X1 port map( A1 => n36102, A2 => n30680, ZN => n36101);
   U133 : NAND2_X1 port map( A1 => n11634, A2 => n29263, ZN => n11595);
   U136 : NAND2_X1 port map( A1 => n773, A2 => n4879, ZN => n33093);
   U140 : NAND2_X1 port map( A1 => n36481, A2 => n30160, ZN => n38883);
   U145 : NAND2_X1 port map( A1 => n29781, A2 => n34000, ZN => n10746);
   U146 : INV_X1 port map( I => n15089, ZN => n37858);
   U148 : OAI21_X1 port map( A1 => n37368, A2 => n29942, B => n30059, ZN => 
                           n29171);
   U149 : BUF_X4 port map( I => n29500, Z => n38051);
   U152 : INV_X1 port map( I => n29642, ZN => n37879);
   U155 : BUF_X2 port map( I => n30195, Z => n36225);
   U159 : INV_X1 port map( I => n28843, ZN => n28882);
   U164 : INV_X1 port map( I => n29346, ZN => n38822);
   U168 : CLKBUF_X2 port map( I => n777, Z => n39322);
   U170 : INV_X1 port map( I => n3631, ZN => n38709);
   U172 : NAND2_X1 port map( A1 => n29642, A2 => n29643, ZN => n38129);
   U173 : INV_X1 port map( I => n30156, ZN => n29210);
   U174 : BUF_X2 port map( I => n4671, Z => n31511);
   U175 : INV_X2 port map( I => n30057, ZN => n37021);
   U176 : INV_X1 port map( I => n19428, ZN => n31689);
   U184 : NOR2_X1 port map( A1 => n35823, A2 => n16036, ZN => n38161);
   U186 : NAND2_X1 port map( A1 => n28636, A2 => n10061, ZN => n29025);
   U187 : INV_X1 port map( I => n19571, ZN => n37726);
   U188 : INV_X1 port map( I => n28830, ZN => n1410);
   U192 : NAND2_X1 port map( A1 => n5342, A2 => n8048, ZN => n37637);
   U195 : NOR2_X1 port map( A1 => n38855, A2 => n39473, ZN => n38463);
   U196 : NOR2_X1 port map( A1 => n34173, A2 => n35997, ZN => n37555);
   U197 : NAND2_X1 port map( A1 => n34958, A2 => n39555, ZN => n28331);
   U198 : NAND2_X1 port map( A1 => n39000, A2 => n38997, ZN => n28648);
   U202 : OAI21_X1 port map( A1 => n3018, A2 => n3019, B => n28390, ZN => 
                           n37990);
   U206 : NAND2_X1 port map( A1 => n38399, A2 => n37285, ZN => n31393);
   U207 : NOR2_X1 port map( A1 => n9444, A2 => n11614, ZN => n37558);
   U208 : NAND2_X1 port map( A1 => n28268, A2 => n16691, ZN => n15109);
   U210 : NAND2_X1 port map( A1 => n28439, A2 => n34176, ZN => n37577);
   U214 : NAND2_X1 port map( A1 => n28336, A2 => n32178, ZN => n38062);
   U215 : OAI22_X1 port map( A1 => n28525, A2 => n28735, B1 => n28736, B2 => 
                           n38172, ZN => n38017);
   U216 : AND2_X1 port map( A1 => n18871, A2 => n28686, Z => n18996);
   U218 : OAI21_X1 port map( A1 => n28726, A2 => n12237, B => n38500, ZN => 
                           n3634);
   U220 : AND2_X1 port map( A1 => n9878, A2 => n28620, Z => n28401);
   U223 : NOR2_X1 port map( A1 => n28386, A2 => n28653, ZN => n28368);
   U225 : NOR2_X1 port map( A1 => n2937, A2 => n1189, ZN => n7913);
   U227 : NAND2_X1 port map( A1 => n39664, A2 => n28755, ZN => n21027);
   U228 : NOR2_X1 port map( A1 => n28485, A2 => n28390, ZN => n28178);
   U230 : NAND2_X1 port map( A1 => n36776, A2 => n36773, ZN => n38469);
   U233 : AND2_X1 port map( A1 => n1186, A2 => n14987, Z => n37128);
   U236 : OAI21_X1 port map( A1 => n16307, A2 => n17596, B => n5396, ZN => 
                           n9585);
   U237 : NAND3_X1 port map( A1 => n28721, A2 => n28362, A3 => n28361, ZN => 
                           n38399);
   U250 : BUF_X2 port map( I => n28464, Z => n19827);
   U251 : OAI21_X1 port map( A1 => n37561, A2 => n37560, B => n28724, ZN => 
                           n36585);
   U255 : NOR2_X1 port map( A1 => n15235, A2 => n15737, ZN => n38861);
   U257 : NAND3_X1 port map( A1 => n15709, A2 => n37981, A3 => n28639, ZN => 
                           n35351);
   U263 : AND2_X1 port map( A1 => n16559, A2 => n16067, Z => n34173);
   U266 : INV_X1 port map( I => n28730, ZN => n50);
   U267 : NOR2_X1 port map( A1 => n37080, A2 => n33283, ZN => n32781);
   U271 : NAND2_X1 port map( A1 => n31888, A2 => n28473, ZN => n8094);
   U275 : NAND2_X1 port map( A1 => n28580, A2 => n1196, ZN => n3052);
   U277 : NOR2_X1 port map( A1 => n28485, A2 => n16559, ZN => n3018);
   U278 : NOR2_X1 port map( A1 => n16067, A2 => n28484, ZN => n6629);
   U281 : NOR2_X1 port map( A1 => n28699, A2 => n28698, ZN => n38503);
   U285 : INV_X1 port map( I => n1823, ZN => n37777);
   U286 : OR2_X1 port map( A1 => n38159, A2 => n17751, Z => n28725);
   U290 : NAND2_X1 port map( A1 => n28716, A2 => n1882, ZN => n28515);
   U291 : NAND2_X1 port map( A1 => n31663, A2 => n37758, ZN => n28440);
   U294 : INV_X2 port map( I => n33283, ZN => n28746);
   U297 : OR2_X1 port map( A1 => n38203, A2 => n39227, Z => n8158);
   U303 : OR2_X1 port map( A1 => n28720, A2 => n28723, Z => n14604);
   U304 : INV_X2 port map( I => n5418, ZN => n36414);
   U306 : BUF_X2 port map( I => n28503, Z => n13891);
   U314 : BUF_X2 port map( I => n28676, Z => n9599);
   U316 : NAND2_X1 port map( A1 => n34861, A2 => n7251, ZN => n38065);
   U317 : AND2_X1 port map( A1 => n28686, A2 => n39724, Z => n10038);
   U318 : AND2_X1 port map( A1 => n10883, A2 => n7063, Z => n5641);
   U321 : NAND2_X1 port map( A1 => n8082, A2 => n11831, ZN => n21141);
   U330 : OR2_X1 port map( A1 => n39227, A2 => n37484, Z => n34510);
   U331 : NOR2_X1 port map( A1 => n28700, A2 => n19349, ZN => n33793);
   U332 : NOR2_X1 port map( A1 => n976, A2 => n13170, ZN => n38657);
   U345 : NAND2_X1 port map( A1 => n38231, A2 => n7429, ZN => n28073);
   U348 : NAND3_X1 port map( A1 => n11330, A2 => n12527, A3 => n36588, ZN => 
                           n38500);
   U352 : NAND2_X1 port map( A1 => n28643, A2 => n14448, ZN => n38999);
   U354 : INV_X1 port map( I => n7905, ZN => n36110);
   U365 : INV_X2 port map( I => n36588, ZN => n39435);
   U366 : AND2_X1 port map( A1 => n31027, A2 => n30668, Z => n38231);
   U368 : NOR2_X1 port map( A1 => n35203, A2 => n34559, ZN => n36742);
   U369 : INV_X2 port map( I => n31663, ZN => n1194);
   U370 : BUF_X2 port map( I => n31378, Z => n902);
   U373 : BUF_X1 port map( I => n31663, Z => n39147);
   U374 : INV_X1 port map( I => n28503, ZN => n28533);
   U383 : CLKBUF_X2 port map( I => n33765, Z => n33629);
   U386 : INV_X2 port map( I => n17234, ZN => n32682);
   U390 : INV_X2 port map( I => n34695, ZN => n1196);
   U396 : OAI21_X1 port map( A1 => n15389, A2 => n1444, B => n8368, ZN => 
                           n20584);
   U401 : NAND2_X1 port map( A1 => n11512, A2 => n36643, ZN => n28349);
   U404 : NAND2_X1 port map( A1 => n37785, A2 => n37782, ZN => n27925);
   U411 : BUF_X4 port map( I => n8366, Z => n37758);
   U412 : OAI21_X1 port map( A1 => n39795, A2 => n39794, B => n898, ZN => 
                           n27938);
   U416 : NAND2_X1 port map( A1 => n38490, A2 => n14461, ZN => n28038);
   U417 : NAND3_X1 port map( A1 => n13491, A2 => n37671, A3 => n19525, ZN => 
                           n28144);
   U418 : OAI21_X1 port map( A1 => n30623, A2 => n28028, B => n27948, ZN => 
                           n38288);
   U421 : OAI21_X1 port map( A1 => n12784, A2 => n30995, B => n16544, ZN => 
                           n28284);
   U427 : OAI22_X1 port map( A1 => n36979, A2 => n9969, B1 => n13851, B2 => 
                           n16325, ZN => n38490);
   U432 : NAND3_X1 port map( A1 => n35507, A2 => n21238, A3 => n28249, ZN => 
                           n38923);
   U433 : NOR2_X1 port map( A1 => n37642, A2 => n17057, ZN => n17055);
   U436 : NAND2_X1 port map( A1 => n13409, A2 => n27969, ZN => n35005);
   U437 : NAND3_X1 port map( A1 => n37322, A2 => n28199, A3 => n16461, ZN => 
                           n28202);
   U439 : INV_X1 port map( I => n3990, ZN => n39188);
   U440 : NAND2_X1 port map( A1 => n37784, A2 => n1204, ZN => n37782);
   U443 : NOR2_X1 port map( A1 => n28024, A2 => n14829, ZN => n30623);
   U445 : OR2_X1 port map( A1 => n8207, A2 => n288, Z => n37126);
   U446 : NAND2_X1 port map( A1 => n4347, A2 => n1435, ZN => n38308);
   U453 : OAI22_X1 port map( A1 => n37057, A2 => n988, B1 => n13081, B2 => 
                           n14399, ZN => n8946);
   U456 : NOR3_X1 port map( A1 => n7872, A2 => n1448, A3 => n38579, ZN => 
                           n38868);
   U457 : INV_X1 port map( I => n38419, ZN => n20577);
   U460 : NAND2_X1 port map( A1 => n14562, A2 => n18689, ZN => n27887);
   U468 : NAND2_X1 port map( A1 => n10466, A2 => n10465, ZN => n37334);
   U469 : AOI21_X1 port map( A1 => n37159, A2 => n27896, B => n27973, ZN => 
                           n16706);
   U470 : BUF_X2 port map( I => n27964, Z => n28118);
   U473 : NAND2_X1 port map( A1 => n35061, A2 => n28274, ZN => n32374);
   U474 : NAND2_X1 port map( A1 => n3990, A2 => n3989, ZN => n27981);
   U476 : NAND3_X1 port map( A1 => n28165, A2 => n10642, A3 => n988, ZN => 
                           n37035);
   U477 : NAND3_X1 port map( A1 => n11375, A2 => n11501, A3 => n37078, ZN => 
                           n406);
   U485 : OR2_X1 port map( A1 => n28152, A2 => n16576, Z => n10465);
   U490 : AND2_X1 port map( A1 => n28152, A2 => n16576, Z => n18770);
   U492 : INV_X1 port map( I => n31494, ZN => n37783);
   U498 : OR2_X1 port map( A1 => n9242, A2 => n36197, Z => n2603);
   U503 : NAND2_X1 port map( A1 => n28282, A2 => n33957, ZN => n28067);
   U504 : CLKBUF_X2 port map( I => n18689, Z => n38996);
   U505 : NOR2_X1 port map( A1 => n31942, A2 => n28214, ZN => n34817);
   U508 : NOR2_X1 port map( A1 => n14397, A2 => n36573, ZN => n4767);
   U511 : NAND3_X1 port map( A1 => n37, A2 => n1448, A3 => n38579, ZN => n28325
                           );
   U512 : OAI21_X1 port map( A1 => n38307, A2 => n30995, B => n7528, ZN => 
                           n12809);
   U513 : AOI21_X1 port map( A1 => n37754, A2 => n37753, B => n30773, ZN => 
                           n38327);
   U525 : INV_X1 port map( I => n16576, ZN => n10420);
   U526 : NAND3_X1 port map( A1 => n18777, A2 => n16261, A3 => n34447, ZN => 
                           n12420);
   U535 : NAND2_X1 port map( A1 => n39126, A2 => n39127, ZN => n38678);
   U536 : NAND2_X1 port map( A1 => n28238, A2 => n28236, ZN => n17615);
   U537 : INV_X1 port map( I => n18853, ZN => n39112);
   U544 : BUF_X2 port map( I => n7741, Z => n38579);
   U545 : BUF_X2 port map( I => n33957, Z => n38307);
   U547 : NOR2_X1 port map( A1 => n14397, A2 => n28181, ZN => n39696);
   U548 : INV_X1 port map( I => n11676, ZN => n1436);
   U551 : INV_X1 port map( I => n38453, ZN => n34166);
   U561 : BUF_X2 port map( I => n17405, Z => n2717);
   U562 : INV_X1 port map( I => n2281, ZN => n38620);
   U566 : INV_X1 port map( I => n13877, ZN => n37307);
   U568 : INV_X1 port map( I => n21093, ZN => n38648);
   U569 : INV_X1 port map( I => n31355, ZN => n8364);
   U573 : AOI21_X1 port map( A1 => n27287, A2 => n1080, B => n6010, ZN => 
                           n16162);
   U576 : NAND3_X1 port map( A1 => n10998, A2 => n27059, A3 => n10999, ZN => 
                           n10997);
   U577 : BUF_X2 port map( I => n31767, Z => n37812);
   U579 : NOR2_X1 port map( A1 => n27172, A2 => n19062, ZN => n27549);
   U587 : AND2_X1 port map( A1 => n8253, A2 => n1082, Z => n8252);
   U590 : NAND3_X1 port map( A1 => n37552, A2 => n16514, A3 => n16516, ZN => 
                           n35718);
   U594 : NAND2_X1 port map( A1 => n3672, A2 => n3674, ZN => n38078);
   U596 : OAI22_X1 port map( A1 => n5059, A2 => n27310, B1 => n37001, B2 => 
                           n27155, ZN => n35123);
   U599 : OR2_X1 port map( A1 => n16520, A2 => n27153, Z => n37552);
   U601 : OAI21_X1 port map( A1 => n30871, A2 => n2035, B => n33335, ZN => 
                           n30584);
   U603 : AOI21_X1 port map( A1 => n27250, A2 => n27007, B => n27251, ZN => 
                           n5770);
   U607 : NAND2_X1 port map( A1 => n30582, A2 => n37170, ZN => n17107);
   U609 : NAND2_X1 port map( A1 => n10032, A2 => n35905, ZN => n38047);
   U610 : OAI21_X1 port map( A1 => n37704, A2 => n37703, B => n37040, ZN => 
                           n35914);
   U611 : NAND2_X1 port map( A1 => n36744, A2 => n33619, ZN => n16306);
   U613 : NAND2_X1 port map( A1 => n37512, A2 => n27398, ZN => n27073);
   U614 : INV_X1 port map( I => n35243, ZN => n31584);
   U620 : OAI22_X1 port map( A1 => n14327, A2 => n6908, B1 => n2761, B2 => 
                           n27165, ZN => n14326);
   U621 : NOR2_X1 port map( A1 => n2207, A2 => n32020, ZN => n39236);
   U624 : NAND2_X1 port map( A1 => n5059, A2 => n39206, ZN => n38481);
   U631 : OAI21_X1 port map( A1 => n39632, A2 => n6534, B => n38690, ZN => 
                           n34570);
   U634 : AND2_X1 port map( A1 => n17095, A2 => n3977, Z => n11038);
   U636 : NAND3_X1 port map( A1 => n7588, A2 => n33088, A3 => n18717, ZN => 
                           n10578);
   U639 : INV_X1 port map( I => n26749, ZN => n491);
   U645 : INV_X1 port map( I => n27393, ZN => n31400);
   U646 : NAND2_X1 port map( A1 => n39632, A2 => n6534, ZN => n37854);
   U648 : NAND2_X1 port map( A1 => n37655, A2 => n37652, ZN => n32545);
   U649 : NOR2_X1 port map( A1 => n32555, A2 => n34167, ZN => n39230);
   U655 : NOR2_X1 port map( A1 => n32566, A2 => n38187, ZN => n3531);
   U658 : NAND2_X1 port map( A1 => n12020, A2 => n35826, ZN => n39565);
   U660 : NOR2_X1 port map( A1 => n161, A2 => n160, ZN => n30667);
   U664 : CLKBUF_X2 port map( I => n1226, Z => n34520);
   U665 : OR2_X1 port map( A1 => n32926, A2 => n36496, Z => n37170);
   U667 : INV_X1 port map( I => n37603, ZN => n30732);
   U674 : NAND2_X1 port map( A1 => n27021, A2 => n15360, ZN => n38276);
   U677 : NAND2_X1 port map( A1 => n38489, A2 => n38488, ZN => n6195);
   U679 : NAND2_X1 port map( A1 => n13294, A2 => n36911, ZN => n38565);
   U680 : OR2_X1 port map( A1 => n14881, A2 => n35895, Z => n32960);
   U682 : NAND2_X1 port map( A1 => n14327, A2 => n27389, ZN => n34733);
   U691 : NAND2_X1 port map( A1 => n20133, A2 => n10051, ZN => n37465);
   U693 : NAND2_X1 port map( A1 => n35332, A2 => n27304, ZN => n39283);
   U694 : NOR2_X1 port map( A1 => n27230, A2 => n1085, ZN => n37704);
   U698 : NAND3_X1 port map( A1 => n4782, A2 => n16782, A3 => n33593, ZN => 
                           n36744);
   U700 : OAI21_X1 port map( A1 => n27270, A2 => n27196, B => n27272, ZN => 
                           n38739);
   U701 : OAI21_X1 port map( A1 => n19557, A2 => n7096, B => n1225, ZN => 
                           n39573);
   U707 : NAND2_X1 port map( A1 => n27357, A2 => n27358, ZN => n2208);
   U708 : NAND2_X1 port map( A1 => n5101, A2 => n39414, ZN => n27456);
   U709 : OR2_X1 port map( A1 => n10171, A2 => n2722, Z => n27090);
   U711 : OR2_X1 port map( A1 => n1788, A2 => n7757, Z => n37076);
   U712 : AND2_X1 port map( A1 => n31006, A2 => n7424, Z => n37246);
   U713 : INV_X2 port map( I => n27164, ZN => n20981);
   U714 : OR2_X1 port map( A1 => n27248, A2 => n7975, Z => n35730);
   U716 : BUF_X2 port map( I => n3540, Z => n36865);
   U717 : NAND2_X1 port map( A1 => n27378, A2 => n1788, ZN => n27071);
   U718 : NAND2_X1 port map( A1 => n11083, A2 => n14153, ZN => n14086);
   U727 : OAI22_X1 port map( A1 => n998, A2 => n35265, B1 => n32829, B2 => 
                           n27424, ZN => n9268);
   U731 : AND2_X1 port map( A1 => n19455, A2 => n27197, Z => n14695);
   U733 : INV_X1 port map( I => n31014, ZN => n30758);
   U734 : NAND2_X1 port map( A1 => n36200, A2 => n34969, ZN => n16170);
   U736 : INV_X1 port map( I => n27452, ZN => n5932);
   U737 : INV_X1 port map( I => n36969, ZN => n2923);
   U738 : INV_X1 port map( I => n27095, ZN => n33593);
   U743 : INV_X1 port map( I => n5588, ZN => n39546);
   U748 : INV_X2 port map( I => n9875, ZN => n21144);
   U752 : NAND2_X1 port map( A1 => n27211, A2 => n34977, ZN => n27441);
   U762 : INV_X2 port map( I => n11820, ZN => n10051);
   U765 : INV_X1 port map( I => n27434, ZN => n39150);
   U766 : CLKBUF_X4 port map( I => n32566, Z => n36528);
   U768 : NAND3_X1 port map( A1 => n4782, A2 => n2660, A3 => n36496, ZN => 
                           n38618);
   U769 : NAND2_X1 port map( A1 => n4272, A2 => n6191, ZN => n15641);
   U771 : INV_X2 port map( I => n39050, ZN => n39826);
   U772 : BUF_X2 port map( I => n27446, Z => n4782);
   U773 : OAI21_X1 port map( A1 => n30365, A2 => n32958, B => n36477, ZN => 
                           n36476);
   U774 : BUF_X2 port map( I => n998, Z => n30544);
   U777 : NAND3_X1 port map( A1 => n26892, A2 => n4325, A3 => n33396, ZN => 
                           n4324);
   U778 : NOR3_X1 port map( A1 => n26663, A2 => n32009, A3 => n26662, ZN => 
                           n39754);
   U782 : NOR2_X1 port map( A1 => n38234, A2 => n38233, ZN => n38232);
   U784 : NOR2_X1 port map( A1 => n35403, A2 => n37373, ZN => n37694);
   U787 : NAND2_X1 port map( A1 => n37133, A2 => n38393, ZN => n5264);
   U789 : NOR2_X1 port map( A1 => n9058, A2 => n15352, ZN => n37735);
   U792 : NAND2_X1 port map( A1 => n26755, A2 => n38268, ZN => n32917);
   U798 : NAND2_X1 port map( A1 => n38955, A2 => n6261, ZN => n31406);
   U802 : NAND2_X1 port map( A1 => n38498, A2 => n4489, ZN => n30689);
   U803 : OAI21_X1 port map( A1 => n14458, A2 => n39342, B => n7596, ZN => 
                           n3283);
   U804 : NAND2_X1 port map( A1 => n10736, A2 => n26695, ZN => n32928);
   U805 : OAI21_X1 port map( A1 => n26661, A2 => n19449, B => n16773, ZN => 
                           n3282);
   U807 : AOI21_X1 port map( A1 => n26799, A2 => n39514, B => n18773, ZN => 
                           n9240);
   U809 : NAND2_X1 port map( A1 => n7619, A2 => n1235, ZN => n10567);
   U815 : NAND2_X1 port map( A1 => n4007, A2 => n33352, ZN => n30643);
   U817 : NAND2_X1 port map( A1 => n26618, A2 => n31701, ZN => n20604);
   U818 : AOI21_X1 port map( A1 => n875, A2 => n26937, B => n11334, ZN => 
                           n37549);
   U824 : NAND2_X1 port map( A1 => n26459, A2 => n735, ZN => n9166);
   U828 : NOR2_X1 port map( A1 => n1231, A2 => n30665, ZN => n26624);
   U838 : AND2_X1 port map( A1 => n849, A2 => n9178, Z => n37074);
   U844 : NAND2_X1 port map( A1 => n33063, A2 => n33062, ZN => n37766);
   U847 : NAND2_X1 port map( A1 => n38715, A2 => n16941, ZN => n39222);
   U848 : OAI21_X1 port map( A1 => n11325, A2 => n4970, B => n1093, ZN => 
                           n38498);
   U850 : INV_X1 port map( I => n11334, ZN => n38824);
   U851 : NAND2_X1 port map( A1 => n26944, A2 => n26849, ZN => n38393);
   U853 : INV_X1 port map( I => n26943, ZN => n36146);
   U864 : OAI21_X1 port map( A1 => n278, A2 => n1786, B => n8917, ZN => n37562)
                           ;
   U867 : NOR2_X1 port map( A1 => n26639, A2 => n862, ZN => n37286);
   U872 : INV_X1 port map( I => n37288, ZN => n37287);
   U873 : NAND2_X1 port map( A1 => n17047, A2 => n6615, ZN => n38684);
   U875 : NAND2_X1 port map( A1 => n11248, A2 => n26910, ZN => n38549);
   U878 : OAI21_X1 port map( A1 => n5935, A2 => n19331, B => n15998, ZN => 
                           n39646);
   U879 : NOR3_X1 port map( A1 => n13686, A2 => n5960, A3 => n14080, ZN => 
                           n5963);
   U880 : AOI22_X1 port map( A1 => n21192, A2 => n26826, B1 => n26769, B2 => 
                           n14488, ZN => n39557);
   U882 : NAND2_X1 port map( A1 => n39758, A2 => n26923, ZN => n39508);
   U884 : NOR2_X1 port map( A1 => n13854, A2 => n13088, ZN => n38233);
   U885 : AOI21_X1 port map( A1 => n278, A2 => n1786, B => n8415, ZN => n34601)
                           ;
   U888 : NAND3_X1 port map( A1 => n26991, A2 => n26989, A3 => n26990, ZN => 
                           n5477);
   U891 : NAND3_X1 port map( A1 => n11616, A2 => n38644, A3 => n10231, ZN => 
                           n38268);
   U895 : AND2_X1 port map( A1 => n20321, A2 => n37084, Z => n2929);
   U901 : AND2_X1 port map( A1 => n11636, A2 => n38280, Z => n26777);
   U910 : AND2_X1 port map( A1 => n15037, A2 => n35256, Z => n2491);
   U918 : INV_X1 port map( I => n860, ZN => n37955);
   U926 : NOR2_X1 port map( A1 => n32345, A2 => n20211, ZN => n3935);
   U927 : NOR2_X1 port map( A1 => n33279, A2 => n32168, ZN => n37281);
   U928 : BUF_X2 port map( I => n26704, Z => n7978);
   U932 : NOR2_X1 port map( A1 => n441, A2 => n26639, ZN => n34108);
   U937 : OR2_X1 port map( A1 => n875, A2 => n17993, Z => n37154);
   U941 : NOR2_X1 port map( A1 => n2451, A2 => n26639, ZN => n12236);
   U953 : OR2_X1 port map( A1 => n26932, A2 => n37235, Z => n17617);
   U955 : AOI21_X1 port map( A1 => n862, A2 => n9690, B => n37289, ZN => n37288
                           );
   U956 : INV_X1 port map( I => n33455, ZN => n9081);
   U958 : INV_X1 port map( I => n9801, ZN => n38591);
   U969 : INV_X1 port map( I => n19728, ZN => n38592);
   U971 : INV_X1 port map( I => n859, ZN => n36477);
   U973 : INV_X1 port map( I => n13528, ZN => n37856);
   U974 : INV_X1 port map( I => n26704, ZN => n6190);
   U980 : OR2_X1 port map( A1 => n18390, A2 => n31897, Z => n35622);
   U984 : INV_X1 port map( I => n26988, ZN => n26819);
   U986 : CLKBUF_X2 port map( I => n5274, Z => n33352);
   U988 : OR2_X1 port map( A1 => n20321, A2 => n37084, Z => n26667);
   U989 : NAND2_X1 port map( A1 => n30859, A2 => n26988, ZN => n26606);
   U990 : INV_X1 port map( I => n36355, ZN => n36873);
   U992 : INV_X1 port map( I => n36931, ZN => n30284);
   U997 : INV_X1 port map( I => n39353, ZN => n36355);
   U998 : INV_X1 port map( I => n39207, ZN => n39825);
   U1001 : INV_X1 port map( I => n37588, ZN => n6454);
   U1003 : INV_X1 port map( I => n26511, ZN => n39561);
   U1006 : BUF_X2 port map( I => n32253, Z => n38844);
   U1007 : CLKBUF_X2 port map( I => n31965, Z => n36758);
   U1008 : INV_X1 port map( I => n26420, ZN => n3330);
   U1011 : INV_X1 port map( I => n13853, ZN => n26451);
   U1015 : INV_X1 port map( I => n26356, ZN => n33504);
   U1017 : BUF_X2 port map( I => n10076, Z => n39129);
   U1021 : INV_X2 port map( I => n26517, ZN => n39662);
   U1024 : AOI21_X1 port map( A1 => n26236, A2 => n26237, B => n30883, ZN => 
                           n26240);
   U1030 : NOR2_X1 port map( A1 => n25785, A2 => n30595, ZN => n10457);
   U1033 : AOI21_X1 port map( A1 => n38953, A2 => n10724, B => n13869, ZN => 
                           n11424);
   U1035 : INV_X1 port map( I => n6989, ZN => n39135);
   U1039 : NOR2_X1 port map( A1 => n38437, A2 => n8407, ZN => n13121);
   U1042 : NAND2_X1 port map( A1 => n37745, A2 => n38501, ZN => n32380);
   U1047 : OAI21_X1 port map( A1 => n20235, A2 => n25800, B => n17951, ZN => 
                           n37618);
   U1050 : NOR2_X1 port map( A1 => n34339, A2 => n12910, ZN => n38386);
   U1051 : NOR2_X1 port map( A1 => n16867, A2 => n25965, ZN => n2837);
   U1057 : NAND2_X1 port map( A1 => n16977, A2 => n37996, ZN => n25918);
   U1060 : NAND3_X1 port map( A1 => n1098, A2 => n38409, A3 => n26119, ZN => 
                           n20062);
   U1071 : NAND2_X1 port map( A1 => n3518, A2 => n26084, ZN => n10270);
   U1076 : NAND2_X1 port map( A1 => n32243, A2 => n18354, ZN => n18353);
   U1078 : OAI21_X1 port map( A1 => n14650, A2 => n25978, B => n31496, ZN => 
                           n37365);
   U1079 : NAND3_X1 port map( A1 => n25764, A2 => n13869, A3 => n34217, ZN => 
                           n30571);
   U1088 : AOI22_X1 port map( A1 => n1515, A2 => n7460, B1 => n8005, B2 => 
                           n1240, ZN => n34554);
   U1090 : AOI22_X1 port map( A1 => n25788, A2 => n1514, B1 => n17371, B2 => 
                           n17372, ZN => n13389);
   U1111 : INV_X1 port map( I => n9859, ZN => n25886);
   U1116 : INV_X1 port map( I => n34399, ZN => n37416);
   U1118 : INV_X1 port map( I => n37462, ZN => n34117);
   U1122 : NOR2_X1 port map( A1 => n25836, A2 => n3213, ZN => n25861);
   U1125 : NAND2_X1 port map( A1 => n35151, A2 => n18661, ZN => n26111);
   U1129 : BUF_X2 port map( I => n7512, Z => n32243);
   U1146 : NOR2_X1 port map( A1 => n15832, A2 => n15831, ZN => n39509);
   U1147 : AOI22_X1 port map( A1 => n11552, A2 => n25993, B1 => n25956, B2 => 
                           n9413, ZN => n25510);
   U1148 : INV_X1 port map( I => n31624, ZN => n3518);
   U1149 : CLKBUF_X2 port map( I => n9802, Z => n33218);
   U1151 : NAND2_X1 port map( A1 => n32924, A2 => n38432, ZN => n33764);
   U1158 : AND2_X1 port map( A1 => n26125, A2 => n39454, Z => n4191);
   U1159 : NAND2_X1 port map( A1 => n38437, A2 => n26041, ZN => n34254);
   U1165 : NAND2_X1 port map( A1 => n39030, A2 => n32690, ZN => n25910);
   U1166 : NAND2_X1 port map( A1 => n10223, A2 => n10764, ZN => n7915);
   U1172 : OR2_X1 port map( A1 => n26015, A2 => n25801, Z => n26121);
   U1176 : NOR2_X1 port map( A1 => n26120, A2 => n25903, ZN => n39143);
   U1184 : OAI21_X1 port map( A1 => n25978, A2 => n1100, B => n34265, ZN => 
                           n37930);
   U1191 : OAI22_X1 port map( A1 => n1523, A2 => n25868, B1 => n26021, B2 => 
                           n1524, ZN => n13440);
   U1195 : AND2_X1 port map( A1 => n6904, A2 => n26124, Z => n37072);
   U1196 : BUF_X2 port map( I => n26048, Z => n1523);
   U1197 : INV_X2 port map( I => n35003, ZN => n13869);
   U1212 : INV_X2 port map( I => n3575, ZN => n6222);
   U1214 : NOR3_X1 port map( A1 => n37683, A2 => n1012, A3 => n25992, ZN => 
                           n8233);
   U1216 : BUF_X2 port map( I => n14890, Z => n4163);
   U1219 : CLKBUF_X4 port map( I => n10986, Z => n446);
   U1220 : NAND2_X1 port map( A1 => n25989, A2 => n34217, ZN => n38550);
   U1224 : INV_X1 port map( I => n598, ZN => n1018);
   U1226 : CLKBUF_X4 port map( I => n6904, Z => n4602);
   U1227 : NAND2_X1 port map( A1 => n32196, A2 => n20813, ZN => n38509);
   U1229 : NAND2_X1 port map( A1 => n951, A2 => n13712, ZN => n32558);
   U1236 : INV_X2 port map( I => n26134, ZN => n1105);
   U1238 : NAND2_X1 port map( A1 => n37393, A2 => n17212, ZN => n17211);
   U1241 : INV_X1 port map( I => n34350, ZN => n10404);
   U1243 : NAND2_X1 port map( A1 => n38663, A2 => n39782, ZN => n38185);
   U1247 : NAND2_X1 port map( A1 => n12548, A2 => n25798, ZN => n25856);
   U1249 : BUF_X2 port map( I => n10015, Z => n32196);
   U1251 : CLKBUF_X2 port map( I => n598, Z => n38247);
   U1252 : INV_X2 port map( I => n6830, ZN => n6390);
   U1253 : CLKBUF_X2 port map( I => n25801, Z => n7423);
   U1257 : AOI22_X1 port map( A1 => n25541, A2 => n36486, B1 => n5042, B2 => 
                           n25542, ZN => n39782);
   U1260 : NOR2_X1 port map( A1 => n38675, A2 => n13301, ZN => n37596);
   U1272 : OAI21_X1 port map( A1 => n39390, A2 => n37174, B => n11951, ZN => 
                           n32827);
   U1274 : OAI21_X1 port map( A1 => n33597, A2 => n25364, B => n37905, ZN => 
                           n38662);
   U1279 : NOR2_X1 port map( A1 => n25697, A2 => n37119, ZN => n16230);
   U1283 : OAI21_X1 port map( A1 => n25622, A2 => n25365, B => n33114, ZN => 
                           n7890);
   U1289 : NAND2_X1 port map( A1 => n33268, A2 => n25248, ZN => n9146);
   U1291 : AND2_X1 port map( A1 => n25699, A2 => n31721, Z => n37181);
   U1292 : NOR2_X1 port map( A1 => n39327, A2 => n30317, ZN => n38675);
   U1293 : AND2_X1 port map( A1 => n14401, A2 => n19863, Z => n34099);
   U1295 : OAI21_X1 port map( A1 => n32076, A2 => n2149, B => n1530, ZN => 
                           n39144);
   U1296 : AND2_X1 port map( A1 => n25577, A2 => n1109, Z => n37174);
   U1301 : NOR2_X1 port map( A1 => n37336, A2 => n19767, ZN => n36020);
   U1302 : OAI21_X1 port map( A1 => n25448, A2 => n25583, B => n38782, ZN => 
                           n38004);
   U1316 : AND2_X1 port map( A1 => n15515, A2 => n32026, Z => n25525);
   U1317 : NAND2_X1 port map( A1 => n7926, A2 => n36345, ZN => n39352);
   U1320 : NOR2_X1 port map( A1 => n10158, A2 => n7284, ZN => n16410);
   U1321 : OAI21_X1 port map( A1 => n31721, A2 => n25699, B => n12931, ZN => 
                           n5034);
   U1324 : NOR2_X1 port map( A1 => n25381, A2 => n1109, ZN => n39390);
   U1327 : NOR3_X1 port map( A1 => n15443, A2 => n11150, A3 => n14553, ZN => 
                           n15422);
   U1328 : OAI21_X1 port map( A1 => n19336, A2 => n25248, B => n12896, ZN => 
                           n37647);
   U1337 : OAI21_X1 port map( A1 => n6747, A2 => n20441, B => n38223, ZN => 
                           n9336);
   U1340 : NAND2_X1 port map( A1 => n25682, A2 => n25681, ZN => n19490);
   U1343 : INV_X1 port map( I => n25489, ZN => n38364);
   U1345 : OR2_X1 port map( A1 => n13413, A2 => n11060, Z => n16315);
   U1353 : OR2_X1 port map( A1 => n19941, A2 => n24896, Z => n20296);
   U1354 : BUF_X2 port map( I => n25513, Z => n39327);
   U1358 : NAND2_X1 port map( A1 => n1551, A2 => n371, ZN => n14805);
   U1360 : CLKBUF_X2 port map( I => n25359, Z => n39321);
   U1366 : CLKBUF_X2 port map( I => n25619, Z => n9594);
   U1370 : CLKBUF_X1 port map( I => n24741, Z => n36249);
   U1372 : NOR2_X1 port map( A1 => n10055, A2 => n6300, ZN => n4824);
   U1374 : NOR2_X1 port map( A1 => n33114, A2 => n33384, ZN => n33113);
   U1375 : OAI21_X1 port map( A1 => n25142, A2 => n20924, B => n37844, ZN => 
                           n39568);
   U1397 : NAND2_X1 port map( A1 => n37845, A2 => n38782, ZN => n4217);
   U1400 : NOR2_X1 port map( A1 => n20924, A2 => n11874, ZN => n11873);
   U1404 : NAND2_X1 port map( A1 => n9132, A2 => n37051, ZN => n2462);
   U1410 : NAND2_X1 port map( A1 => n25674, A2 => n25677, ZN => n39700);
   U1415 : NAND3_X1 port map( A1 => n6065, A2 => n32450, A3 => n1252, ZN => 
                           n35710);
   U1416 : AOI21_X1 port map( A1 => n25600, A2 => n33491, B => n25601, ZN => 
                           n37348);
   U1417 : INV_X1 port map( I => n32989, ZN => n19678);
   U1418 : INV_X1 port map( I => n33491, ZN => n34755);
   U1421 : INV_X1 port map( I => n38849, ZN => n18545);
   U1422 : INV_X1 port map( I => n32775, ZN => n20815);
   U1423 : CLKBUF_X2 port map( I => n31669, Z => n39160);
   U1425 : CLKBUF_X2 port map( I => n19941, Z => n39371);
   U1433 : AND2_X1 port map( A1 => n20595, A2 => n19696, Z => n34060);
   U1434 : NAND2_X1 port map( A1 => n12944, A2 => n20924, ZN => n37844);
   U1435 : BUF_X2 port map( I => n32989, Z => n5166);
   U1439 : INV_X1 port map( I => n25619, ZN => n11874);
   U1447 : NOR2_X1 port map( A1 => n25449, A2 => n25582, ZN => n37845);
   U1448 : NOR2_X1 port map( A1 => n1548, A2 => n17774, ZN => n15620);
   U1449 : INV_X1 port map( I => n39778, ZN => n34150);
   U1450 : INV_X1 port map( I => n25072, ZN => n5800);
   U1451 : INV_X1 port map( I => n25254, ZN => n20347);
   U1452 : INV_X1 port map( I => n15930, ZN => n25250);
   U1457 : CLKBUF_X2 port map( I => n25136, Z => n39756);
   U1460 : INV_X1 port map( I => n13935, ZN => n6984);
   U1480 : INV_X1 port map( I => n25237, ZN => n39582);
   U1482 : INV_X2 port map( I => n25259, ZN => n1260);
   U1483 : INV_X1 port map( I => n9701, ZN => n38336);
   U1487 : NAND2_X1 port map( A1 => n38242, A2 => n2505, ZN => n2503);
   U1488 : INV_X1 port map( I => n25079, ZN => n25258);
   U1502 : OAI21_X1 port map( A1 => n33317, A2 => n37115, B => n38521, ZN => 
                           n20665);
   U1509 : NAND2_X1 port map( A1 => n39469, A2 => n33666, ZN => n38083);
   U1511 : CLKBUF_X2 port map( I => n36908, Z => n36228);
   U1513 : CLKBUF_X2 port map( I => n20411, Z => n39157);
   U1514 : NOR2_X1 port map( A1 => n31698, A2 => n39704, ZN => n33449);
   U1521 : AOI21_X1 port map( A1 => n31213, A2 => n37355, B => n24655, ZN => 
                           n24657);
   U1526 : NOR2_X1 port map( A1 => n24789, A2 => n20039, ZN => n37830);
   U1542 : NAND2_X1 port map( A1 => n33317, A2 => n24899, ZN => n38521);
   U1544 : NAND2_X1 port map( A1 => n957, A2 => n31845, ZN => n15585);
   U1547 : AND2_X1 port map( A1 => n2731, A2 => n24674, Z => n37202);
   U1548 : NOR2_X1 port map( A1 => n19886, A2 => n24565, ZN => n39712);
   U1549 : NAND2_X1 port map( A1 => n6791, A2 => n1784, ZN => n1783);
   U1550 : AND2_X1 port map( A1 => n24715, A2 => n39268, Z => n16908);
   U1555 : AOI21_X1 port map( A1 => n24909, A2 => n36634, B => n36752, ZN => 
                           n6229);
   U1562 : NOR2_X1 port map( A1 => n31198, A2 => n3697, ZN => n37684);
   U1564 : NOR2_X1 port map( A1 => n1120, A2 => n36082, ZN => n24765);
   U1568 : NAND2_X1 port map( A1 => n38978, A2 => n8264, ZN => n33401);
   U1570 : NAND2_X1 port map( A1 => n39817, A2 => n5888, ZN => n9071);
   U1574 : INV_X1 port map( I => n34141, ZN => n38293);
   U1580 : NOR2_X1 port map( A1 => n31861, A2 => n38182, ZN => n20944);
   U1582 : NOR3_X1 port map( A1 => n24775, A2 => n24292, A3 => n35801, ZN => 
                           n4578);
   U1586 : NAND2_X1 port map( A1 => n5063, A2 => n37474, ZN => n38286);
   U1591 : NOR2_X1 port map( A1 => n39085, A2 => n37276, ZN => n37275);
   U1597 : NOR2_X1 port map( A1 => n9197, A2 => n9198, ZN => n30384);
   U1600 : NAND2_X1 port map( A1 => n2731, A2 => n15282, ZN => n38795);
   U1606 : OAI21_X1 port map( A1 => n36988, A2 => n24648, B => n37477, ZN => 
                           n24514);
   U1612 : AOI21_X1 port map( A1 => n31385, A2 => n24866, B => n30554, ZN => 
                           n7970);
   U1618 : NOR2_X1 port map( A1 => n16210, A2 => n18110, ZN => n16949);
   U1619 : NOR2_X1 port map( A1 => n24899, A2 => n1268, ZN => n35170);
   U1620 : NOR3_X1 port map( A1 => n9921, A2 => n24685, A3 => n24686, ZN => 
                           n815);
   U1623 : INV_X1 port map( I => n24572, ZN => n16208);
   U1625 : NAND2_X1 port map( A1 => n24529, A2 => n5897, ZN => n13050);
   U1633 : NAND3_X1 port map( A1 => n34662, A2 => n16815, A3 => n37395, ZN => 
                           n38389);
   U1637 : CLKBUF_X2 port map( I => n39098, Z => n38984);
   U1641 : INV_X1 port map( I => n24712, ZN => n24899);
   U1642 : INV_X1 port map( I => n39279, ZN => n30699);
   U1644 : INV_X1 port map( I => n10054, ZN => n14857);
   U1652 : INV_X2 port map( I => n14283, ZN => n1121);
   U1654 : INV_X1 port map( I => n35250, ZN => n16815);
   U1656 : NAND2_X1 port map( A1 => n35443, A2 => n24650, ZN => n24868);
   U1660 : INV_X2 port map( I => n37477, ZN => n14241);
   U1667 : BUF_X2 port map( I => n5634, Z => n37737);
   U1668 : BUF_X2 port map( I => n2616, Z => n31213);
   U1677 : NAND2_X1 port map( A1 => n24811, A2 => n37277, ZN => n37276);
   U1678 : INV_X1 port map( I => n24227, ZN => n38744);
   U1680 : CLKBUF_X2 port map( I => n32637, Z => n39085);
   U1681 : NOR2_X1 port map( A1 => n7871, A2 => n1577, ZN => n37318);
   U1686 : INV_X2 port map( I => n3510, ZN => n36752);
   U1690 : NOR2_X1 port map( A1 => n36716, A2 => n5768, ZN => n6744);
   U1691 : NOR2_X1 port map( A1 => n24875, A2 => n24876, ZN => n36017);
   U1694 : AOI21_X1 port map( A1 => n24829, A2 => n14064, B => n13665, ZN => 
                           n13666);
   U1703 : NOR2_X1 port map( A1 => n24565, A2 => n32637, ZN => n24528);
   U1708 : AOI21_X1 port map( A1 => n24592, A2 => n24847, B => n35960, ZN => 
                           n24593);
   U1710 : NAND2_X1 port map( A1 => n23857, A2 => n31845, ZN => n37537);
   U1714 : NAND2_X1 port map( A1 => n24855, A2 => n35373, ZN => n24856);
   U1716 : INV_X2 port map( I => n39406, ZN => n9198);
   U1718 : NAND2_X1 port map( A1 => n39523, A2 => n36395, ZN => n24897);
   U1720 : NOR2_X1 port map( A1 => n38658, A2 => n24783, ZN => n24177);
   U1724 : NOR2_X1 port map( A1 => n8317, A2 => n31385, ZN => n31483);
   U1725 : OR2_X1 port map( A1 => n5282, A2 => n38749, Z => n32390);
   U1727 : INV_X1 port map( I => n39098, ZN => n18324);
   U1731 : NOR2_X1 port map( A1 => n31796, A2 => n38848, ZN => n39265);
   U1733 : AOI21_X1 port map( A1 => n31845, A2 => n1574, B => n1026, ZN => 
                           n10403);
   U1740 : NAND2_X1 port map( A1 => n7810, A2 => n32831, ZN => n38978);
   U1746 : INV_X1 port map( I => n32651, ZN => n37277);
   U1747 : INV_X1 port map( I => n30845, ZN => n24820);
   U1750 : INV_X1 port map( I => n15414, ZN => n13665);
   U1751 : INV_X1 port map( I => n36908, ZN => n38973);
   U1758 : BUF_X2 port map( I => n14729, Z => n7286);
   U1760 : BUF_X2 port map( I => n24827, Z => n5431);
   U1765 : BUF_X4 port map( I => n24817, Z => n37106);
   U1766 : NAND2_X1 port map( A1 => n19420, A2 => n36385, ZN => n7871);
   U1773 : NOR2_X1 port map( A1 => n1120, A2 => n39098, ZN => n18168);
   U1779 : BUF_X2 port map( I => n18788, Z => n9997);
   U1780 : NAND2_X1 port map( A1 => n24674, A2 => n15281, ZN => n24226);
   U1782 : NAND2_X1 port map( A1 => n24746, A2 => n39279, ZN => n24602);
   U1786 : OAI21_X1 port map( A1 => n12250, A2 => n12277, B => n19915, ZN => 
                           n12249);
   U1789 : BUF_X4 port map( I => n32136, Z => n37097);
   U1799 : NOR2_X1 port map( A1 => n5957, A2 => n3760, ZN => n5495);
   U1800 : OR2_X1 port map( A1 => n1125, A2 => n9371, Z => n37065);
   U1802 : OR2_X1 port map( A1 => n24098, A2 => n24403, Z => n2342);
   U1803 : NOR2_X1 port map( A1 => n39398, A2 => n39397, ZN => n39244);
   U1805 : AOI22_X1 port map( A1 => n37068, A2 => n1128, B1 => n1588, B2 => 
                           n2579, ZN => n38036);
   U1810 : NAND2_X1 port map( A1 => n24140, A2 => n2336, ZN => n31267);
   U1816 : NOR2_X1 port map( A1 => n4308, A2 => n32818, ZN => n37977);
   U1818 : NAND2_X1 port map( A1 => n36740, A2 => n24234, ZN => n38821);
   U1819 : NAND2_X1 port map( A1 => n39381, A2 => n33531, ZN => n39243);
   U1820 : AOI21_X1 port map( A1 => n24395, A2 => n24182, B => n19739, ZN => 
                           n38526);
   U1821 : NOR2_X1 port map( A1 => n250, A2 => n24443, ZN => n24441);
   U1822 : INV_X1 port map( I => n35314, ZN => n39397);
   U1832 : OAI21_X1 port map( A1 => n8987, A2 => n24219, B => n1124, ZN => 
                           n37388);
   U1839 : NOR2_X1 port map( A1 => n5853, A2 => n31464, ZN => n37672);
   U1840 : NOR2_X1 port map( A1 => n9101, A2 => n1131, ZN => n38405);
   U1841 : NAND2_X1 port map( A1 => n34422, A2 => n33531, ZN => n15365);
   U1845 : INV_X1 port map( I => n32683, ZN => n39398);
   U1848 : OR2_X1 port map( A1 => n1130, A2 => n7240, Z => n37068);
   U1849 : INV_X1 port map( I => n35954, ZN => n35958);
   U1850 : OR2_X1 port map( A1 => n1276, A2 => n15385, Z => n19381);
   U1851 : INV_X1 port map( I => n6715, ZN => n38422);
   U1852 : NOR2_X1 port map( A1 => n24401, A2 => n14392, ZN => n24402);
   U1854 : NAND2_X1 port map( A1 => n33104, A2 => n24258, ZN => n24378);
   U1859 : AOI22_X1 port map( A1 => n10220, A2 => n15049, B1 => n1131, B2 => 
                           n19140, ZN => n38446);
   U1862 : NOR2_X1 port map( A1 => n24382, A2 => n24381, ZN => n17067);
   U1863 : OAI22_X1 port map( A1 => n39156, A2 => n35916, B1 => n24345, B2 => 
                           n20404, ZN => n24350);
   U1864 : NOR2_X1 port map( A1 => n11361, A2 => n24141, ZN => n2989);
   U1865 : NAND2_X1 port map( A1 => n24225, A2 => n16081, ZN => n37958);
   U1866 : AOI22_X1 port map( A1 => n24331, A2 => n24327, B1 => n24174, B2 => 
                           n39057, ZN => n36640);
   U1868 : NAND2_X1 port map( A1 => n24484, A2 => n24241, ZN => n24345);
   U1879 : NAND2_X1 port map( A1 => n1131, A2 => n2597, ZN => n4702);
   U1881 : INV_X1 port map( I => n24433, ZN => n15240);
   U1885 : AND2_X1 port map( A1 => n35233, A2 => n15903, Z => n24207);
   U1889 : AND2_X1 port map( A1 => n12759, A2 => n12758, Z => n24231);
   U1890 : INV_X1 port map( I => n24216, ZN => n38527);
   U1891 : NOR2_X1 port map( A1 => n14655, A2 => n15751, ZN => n12926);
   U1892 : NAND2_X1 port map( A1 => n32683, A2 => n33580, ZN => n24261);
   U1894 : CLKBUF_X2 port map( I => n17693, Z => n37377);
   U1896 : INV_X2 port map( I => n2192, ZN => n39373);
   U1907 : NAND2_X1 port map( A1 => n24328, A2 => n1589, ZN => n15146);
   U1917 : NAND3_X1 port map( A1 => n2439, A2 => n24458, A3 => n38431, ZN => 
                           n32881);
   U1930 : NAND2_X1 port map( A1 => n24169, A2 => n20457, ZN => n24397);
   U1931 : NOR2_X1 port map( A1 => n33314, A2 => n20196, ZN => n20989);
   U1932 : OR2_X1 port map( A1 => n20619, A2 => n24470, Z => n24132);
   U1934 : NAND2_X1 port map( A1 => n16449, A2 => n1283, ZN => n23820);
   U1939 : NAND2_X1 port map( A1 => n35450, A2 => n37267, ZN => n24133);
   U1941 : INV_X1 port map( I => n30494, ZN => n1289);
   U1943 : NAND2_X1 port map( A1 => n1129, A2 => n24360, ZN => n24457);
   U1944 : CLKBUF_X1 port map( I => n6226, Z => n34786);
   U1948 : NOR2_X1 port map( A1 => n2395, A2 => n1589, ZN => n38948);
   U1951 : BUF_X2 port map( I => n33599, Z => n39605);
   U1952 : INV_X1 port map( I => n35242, ZN => n39055);
   U1959 : INV_X1 port map( I => n23598, ZN => n36067);
   U1960 : INV_X1 port map( I => n23775, ZN => n38022);
   U1961 : INV_X1 port map( I => n20205, ZN => n39314);
   U1965 : CLKBUF_X4 port map( I => n39161, Z => n38021);
   U1968 : INV_X1 port map( I => n24034, ZN => n37861);
   U1972 : OAI21_X1 port map( A1 => n23600, A2 => n12597, B => n37649, ZN => 
                           n14107);
   U1980 : BUF_X2 port map( I => n23419, Z => n39408);
   U1981 : NAND2_X1 port map( A1 => n3506, A2 => n23561, ZN => n1830);
   U1996 : AOI21_X1 port map( A1 => n37278, A2 => n17927, B => n23625, ZN => 
                           n17926);
   U1998 : OAI21_X1 port map( A1 => n16715, A2 => n23455, B => n605, ZN => 
                           n33155);
   U1999 : INV_X1 port map( I => n23939, ZN => n39412);
   U2003 : INV_X1 port map( I => n23636, ZN => n23640);
   U2005 : INV_X1 port map( I => n23460, ZN => n37005);
   U2011 : NOR2_X1 port map( A1 => n23521, A2 => n2273, ZN => n9672);
   U2019 : INV_X2 port map( I => n23430, ZN => n37279);
   U2020 : NAND2_X1 port map( A1 => n33869, A2 => n38806, ZN => n18538);
   U2022 : NAND2_X1 port map( A1 => n37528, A2 => n30506, ZN => n32596);
   U2026 : NOR2_X1 port map( A1 => n38335, A2 => n38334, ZN => n35398);
   U2029 : NOR2_X1 port map( A1 => n23522, A2 => n2273, ZN => n23405);
   U2031 : NOR2_X1 port map( A1 => n16728, A2 => n2798, ZN => n39281);
   U2033 : OR2_X1 port map( A1 => n23272, A2 => n36564, Z => n15603);
   U2043 : AND2_X1 port map( A1 => n33786, A2 => n10216, Z => n7886);
   U2046 : NAND2_X1 port map( A1 => n23401, A2 => n32471, ZN => n20867);
   U2052 : NOR2_X1 port map( A1 => n39805, A2 => n17768, ZN => n37482);
   U2055 : NAND2_X1 port map( A1 => n39012, A2 => n23283, ZN => n33911);
   U2056 : OAI21_X1 port map( A1 => n37207, A2 => n36448, B => n37802, ZN => 
                           n23648);
   U2059 : NOR2_X1 port map( A1 => n37839, A2 => n16726, ZN => n34942);
   U2061 : NOR2_X1 port map( A1 => n21130, A2 => n38380, ZN => n23393);
   U2062 : NAND2_X1 port map( A1 => n15458, A2 => n1644, ZN => n37320);
   U2067 : NAND2_X1 port map( A1 => n23302, A2 => n12597, ZN => n37649);
   U2070 : NOR2_X1 port map( A1 => n17995, A2 => n39133, ZN => n37976);
   U2074 : INV_X1 port map( I => n23453, ZN => n16715);
   U2075 : AND2_X1 port map( A1 => n35938, A2 => n23430, Z => n37278);
   U2077 : NOR2_X1 port map( A1 => n3174, A2 => n32061, ZN => n32060);
   U2080 : NAND2_X1 port map( A1 => n23116, A2 => n23117, ZN => n23335);
   U2085 : OAI21_X1 port map( A1 => n11097, A2 => n20031, B => n1036, ZN => 
                           n39276);
   U2086 : NOR2_X1 port map( A1 => n1136, A2 => n38248, ZN => n37569);
   U2087 : OAI21_X1 port map( A1 => n4859, A2 => n1642, B => n23392, ZN => 
                           n6052);
   U2090 : AND2_X1 port map( A1 => n23531, A2 => n33453, Z => n39812);
   U2092 : INV_X1 port map( I => n23505, ZN => n39301);
   U2105 : INV_X1 port map( I => n23568, ZN => n1298);
   U2107 : AND2_X1 port map( A1 => n23440, A2 => n9862, Z => n2454);
   U2109 : NOR2_X1 port map( A1 => n23459, A2 => n35808, ZN => n36431);
   U2114 : NOR3_X1 port map( A1 => n31685, A2 => n18086, A3 => n36539, ZN => 
                           n4396);
   U2115 : CLKBUF_X2 port map( I => n4618, Z => n32351);
   U2122 : NOR2_X1 port map( A1 => n7379, A2 => n10143, ZN => n18391);
   U2133 : NAND2_X1 port map( A1 => n5044, A2 => n6159, ZN => n23574);
   U2135 : NAND2_X1 port map( A1 => n23401, A2 => n33703, ZN => n22872);
   U2136 : NOR2_X1 port map( A1 => n39803, A2 => n9772, ZN => n39428);
   U2143 : CLKBUF_X2 port map( I => n23577, Z => n39214);
   U2144 : BUF_X2 port map( I => n3708, Z => n36103);
   U2145 : CLKBUF_X2 port map( I => n23518, Z => n38252);
   U2148 : NOR2_X1 port map( A1 => n23645, A2 => n37839, ZN => n30417);
   U2150 : NOR2_X1 port map( A1 => n23460, A2 => n23458, ZN => n36430);
   U2156 : NAND2_X1 port map( A1 => n23360, A2 => n14974, ZN => n37779);
   U2157 : NAND2_X1 port map( A1 => n22680, A2 => n22681, ZN => n37514);
   U2163 : NAND2_X1 port map( A1 => n23611, A2 => n4525, ZN => n38651);
   U2165 : NAND2_X1 port map( A1 => n1634, A2 => n38614, ZN => n11436);
   U2169 : INV_X2 port map( I => n23580, ZN => n1138);
   U2170 : NAND2_X1 port map( A1 => n23620, A2 => n16774, ZN => n38971);
   U2180 : NOR2_X1 port map( A1 => n1299, A2 => n39001, ZN => n7048);
   U2184 : INV_X1 port map( I => n38792, ZN => n20278);
   U2185 : AND2_X1 port map( A1 => n12966, A2 => n9862, Z => n23282);
   U2187 : NOR2_X1 port map( A1 => n15353, A2 => n8692, ZN => n32111);
   U2192 : NAND2_X1 port map( A1 => n23637, A2 => n12028, ZN => n23247);
   U2195 : BUF_X2 port map( I => n7644, Z => n32930);
   U2196 : AND2_X1 port map( A1 => n8660, A2 => n38704, Z => n23412);
   U2198 : CLKBUF_X2 port map( I => n35331, Z => n39316);
   U2204 : INV_X1 port map( I => n38614, ZN => n23346);
   U2209 : NOR2_X1 port map( A1 => n38441, A2 => n39070, ZN => n23556);
   U2219 : INV_X2 port map( I => n33747, ZN => n23571);
   U2224 : INV_X2 port map( I => n23337, ZN => n31331);
   U2226 : NAND2_X1 port map( A1 => n17931, A2 => n13029, ZN => n23272);
   U2227 : NAND2_X1 port map( A1 => n23456, A2 => n2553, ZN => n15941);
   U2231 : NOR2_X1 port map( A1 => n30574, A2 => n2553, ZN => n38792);
   U2234 : CLKBUF_X2 port map( I => n10216, Z => n8190);
   U2235 : NAND2_X1 port map( A1 => n19559, A2 => n23487, ZN => n36551);
   U2237 : INV_X2 port map( I => n39001, ZN => n7049);
   U2238 : INV_X1 port map( I => n23296, ZN => n37308);
   U2240 : CLKBUF_X2 port map( I => n33840, Z => n39805);
   U2244 : AOI21_X1 port map( A1 => n33082, A2 => n22907, B => n22906, ZN => 
                           n38173);
   U2250 : INV_X2 port map( I => n13733, ZN => n37774);
   U2251 : INV_X2 port map( I => n37088, ZN => n23389);
   U2252 : CLKBUF_X2 port map( I => n30299, Z => n38119);
   U2253 : BUF_X4 port map( I => n20346, Z => n39401);
   U2256 : NOR2_X1 port map( A1 => n35950, A2 => n37063, ZN => n34615);
   U2259 : NAND2_X1 port map( A1 => n19481, A2 => n35534, ZN => n9856);
   U2264 : INV_X1 port map( I => n16094, ZN => n21293);
   U2268 : NAND2_X1 port map( A1 => n23160, A2 => n38074, ZN => n32909);
   U2269 : NAND2_X1 port map( A1 => n22830, A2 => n22831, ZN => n37980);
   U2272 : OAI21_X1 port map( A1 => n23162, A2 => n22871, B => n22915, ZN => 
                           n37548);
   U2273 : OAI22_X1 port map( A1 => n4714, A2 => n36736, B1 => n1144, B2 => 
                           n8730, ZN => n2102);
   U2275 : NOR2_X1 port map( A1 => n35684, A2 => n10436, ZN => n38074);
   U2276 : NOR2_X1 port map( A1 => n18415, A2 => n22859, ZN => n22863);
   U2277 : NAND2_X1 port map( A1 => n11295, A2 => n22802, ZN => n23123);
   U2278 : NOR2_X1 port map( A1 => n37500, A2 => n284, ZN => n37749);
   U2280 : NAND2_X1 port map( A1 => n18147, A2 => n38789, ZN => n36374);
   U2282 : OAI21_X1 port map( A1 => n1146, A2 => n23053, B => n23114, ZN => 
                           n19229);
   U2283 : NOR2_X1 port map( A1 => n6691, A2 => n37629, ZN => n36167);
   U2285 : INV_X1 port map( I => n11476, ZN => n10507);
   U2286 : NAND3_X1 port map( A1 => n15330, A2 => n13650, A3 => n38986, ZN => 
                           n39819);
   U2298 : NAND2_X1 port map( A1 => n9854, A2 => n35684, ZN => n39526);
   U2300 : AOI21_X1 port map( A1 => n22558, A2 => n39518, B => n6674, ZN => 
                           n38559);
   U2303 : NOR2_X1 port map( A1 => n37589, A2 => n23212, ZN => n38492);
   U2306 : NOR2_X1 port map( A1 => n7071, A2 => n1042, ZN => n38541);
   U2311 : NAND2_X1 port map( A1 => n22836, A2 => n23047, ZN => n38800);
   U2313 : CLKBUF_X4 port map( I => n23125, Z => n37883);
   U2314 : NAND2_X1 port map( A1 => n3862, A2 => n23066, ZN => n35310);
   U2315 : AOI21_X1 port map( A1 => n20872, A2 => n23078, B => n23077, ZN => 
                           n15040);
   U2318 : INV_X1 port map( I => n22800, ZN => n23210);
   U2322 : NAND2_X1 port map( A1 => n5515, A2 => n20372, ZN => n12163);
   U2324 : NAND2_X1 port map( A1 => n14765, A2 => n19535, ZN => n39046);
   U2325 : NAND2_X1 port map( A1 => n17128, A2 => n9651, ZN => n17319);
   U2326 : INV_X1 port map( I => n15330, ZN => n11584);
   U2331 : OAI21_X1 port map( A1 => n936, A2 => n10047, B => n14089, ZN => 
                           n34368);
   U2339 : NOR2_X1 port map( A1 => n15163, A2 => n22944, ZN => n17497);
   U2345 : NAND2_X1 port map( A1 => n12729, A2 => n36422, ZN => n14877);
   U2351 : INV_X1 port map( I => n38790, ZN => n38789);
   U2354 : OAI21_X1 port map( A1 => n10047, A2 => n39303, B => n22816, ZN => 
                           n12621);
   U2361 : NOR2_X1 port map( A1 => n23188, A2 => n22979, ZN => n39205);
   U2362 : NAND2_X1 port map( A1 => n7160, A2 => n33972, ZN => n22473);
   U2365 : INV_X1 port map( I => n4573, ZN => n4931);
   U2368 : OR2_X1 port map( A1 => n7518, A2 => n39446, Z => n23047);
   U2370 : INV_X2 port map( I => n783, ZN => n37922);
   U2373 : BUF_X2 port map( I => n37218, Z => n4713);
   U2379 : CLKBUF_X2 port map( I => n15388, Z => n38601);
   U2383 : OAI21_X1 port map( A1 => n23169, A2 => n36554, B => n23167, ZN => 
                           n38790);
   U2386 : NAND2_X1 port map( A1 => n39811, A2 => n19938, ZN => n23099);
   U2389 : INV_X1 port map( I => n780, ZN => n8730);
   U2390 : NAND2_X1 port map( A1 => n13995, A2 => n17127, ZN => n17124);
   U2392 : BUF_X2 port map( I => n14494, Z => n6646);
   U2397 : INV_X1 port map( I => n11307, ZN => n20783);
   U2398 : INV_X1 port map( I => n22678, ZN => n37764);
   U2399 : BUF_X2 port map( I => n22740, Z => n31863);
   U2407 : CLKBUF_X2 port map( I => n19931, Z => n39682);
   U2409 : INV_X1 port map( I => n19814, ZN => n39559);
   U2411 : OAI21_X1 port map( A1 => n35014, A2 => n34090, B => n22125, ZN => 
                           n36849);
   U2419 : NAND2_X1 port map( A1 => n37454, A2 => n37302, ZN => n17536);
   U2425 : NOR2_X1 port map( A1 => n16403, A2 => n8618, ZN => n38747);
   U2430 : NAND2_X1 port map( A1 => n7355, A2 => n1344, ZN => n38479);
   U2436 : NOR2_X1 port map( A1 => n20299, A2 => n1673, ZN => n20298);
   U2437 : OAI21_X1 port map( A1 => n38287, A2 => n2816, B => n36006, ZN => 
                           n6808);
   U2438 : NAND3_X1 port map( A1 => n554, A2 => n22171, A3 => n18766, ZN => 
                           n16435);
   U2439 : NAND3_X1 port map( A1 => n5345, A2 => n18360, A3 => n5894, ZN => 
                           n39111);
   U2449 : NAND2_X1 port map( A1 => n22152, A2 => n17335, ZN => n22153);
   U2450 : AND2_X1 port map( A1 => n21968, A2 => n35780, Z => n8574);
   U2451 : AND2_X1 port map( A1 => n22349, A2 => n34813, Z => n2909);
   U2452 : AOI21_X1 port map( A1 => n21974, A2 => n21975, B => n32640, ZN => 
                           n21976);
   U2454 : NAND2_X1 port map( A1 => n37794, A2 => n37793, ZN => n22062);
   U2461 : OAI21_X1 port map( A1 => n20758, A2 => n20759, B => n37911, ZN => 
                           n38869);
   U2465 : NOR2_X1 port map( A1 => n33713, A2 => n22294, ZN => n39237);
   U2470 : NOR2_X1 port map( A1 => n7768, A2 => n1332, ZN => n38911);
   U2475 : OAI22_X1 port map( A1 => n37838, A2 => n22360, B1 => n11171, B2 => 
                           n31940, ZN => n11379);
   U2477 : NAND2_X1 port map( A1 => n33489, A2 => n22365, ZN => n22006);
   U2479 : NAND2_X1 port map( A1 => n11276, A2 => n22324, ZN => n37454);
   U2480 : NAND2_X1 port map( A1 => n5894, A2 => n5693, ZN => n4874);
   U2482 : AOI21_X1 port map( A1 => n4108, A2 => n6361, B => n22327, ZN => 
                           n34790);
   U2484 : OR2_X1 port map( A1 => n915, A2 => n3863, Z => n38917);
   U2486 : OAI21_X1 port map( A1 => n6485, A2 => n21002, B => n9987, ZN => 
                           n15017);
   U2492 : NAND3_X1 port map( A1 => n39010, A2 => n1337, A3 => n6297, ZN => 
                           n22020);
   U2494 : NOR2_X1 port map( A1 => n1049, A2 => n3907, ZN => n22045);
   U2496 : OR2_X1 port map( A1 => n22277, A2 => n8493, Z => n37199);
   U2497 : BUF_X2 port map( I => n15697, Z => n38830);
   U2498 : NAND2_X1 port map( A1 => n14423, A2 => n32107, ZN => n22390);
   U2503 : INV_X1 port map( I => n9938, ZN => n37838);
   U2507 : NOR2_X1 port map( A1 => n19873, A2 => n22349, ZN => n38007);
   U2513 : NAND3_X1 port map( A1 => n30893, A2 => n14020, A3 => n38448, ZN => 
                           n37709);
   U2514 : BUF_X2 port map( I => n22240, Z => n16888);
   U2520 : NAND2_X1 port map( A1 => n22073, A2 => n38687, ZN => n39377);
   U2526 : INV_X1 port map( I => n584, ZN => n37794);
   U2527 : NOR2_X1 port map( A1 => n22324, A2 => n22322, ZN => n7636);
   U2529 : INV_X2 port map( I => n33086, ZN => n22261);
   U2532 : NOR2_X1 port map( A1 => n22282, A2 => n22281, ZN => n38700);
   U2534 : BUF_X2 port map( I => n11568, Z => n2910);
   U2538 : BUF_X2 port map( I => n7497, Z => n584);
   U2540 : BUF_X2 port map( I => n20397, Z => n33886);
   U2541 : NAND2_X1 port map( A1 => n32313, A2 => n22263, ZN => n39357);
   U2550 : INV_X2 port map( I => n35780, ZN => n2186);
   U2553 : BUF_X2 port map( I => n18929, Z => n6127);
   U2554 : OR2_X1 port map( A1 => n21345, A2 => n21433, Z => n37180);
   U2556 : BUF_X4 port map( I => n22400, Z => n37089);
   U2558 : AOI21_X1 port map( A1 => n39620, A2 => n21713, B => n39619, ZN => 
                           n39618);
   U2561 : NAND2_X1 port map( A1 => n38546, A2 => n39192, ZN => n38545);
   U2567 : NOR2_X1 port map( A1 => n19650, A2 => n21876, ZN => n21455);
   U2569 : INV_X1 port map( I => n38546, ZN => n39620);
   U2571 : NAND2_X1 port map( A1 => n1372, A2 => n21702, ZN => n38340);
   U2573 : OR2_X1 port map( A1 => n18968, A2 => n917, Z => n37142);
   U2577 : AOI21_X1 port map( A1 => n21784, A2 => n21405, B => n21783, ZN => 
                           n38938);
   U2580 : NOR3_X1 port map( A1 => n21869, A2 => n21870, A3 => n15359, ZN => 
                           n684);
   U2584 : NOR2_X1 port map( A1 => n21808, A2 => n39639, ZN => n21690);
   U2585 : NOR2_X1 port map( A1 => n21914, A2 => n1352, ZN => n5505);
   U2589 : OR2_X1 port map( A1 => n37939, A2 => n39411, Z => n21789);
   U2591 : CLKBUF_X2 port map( I => n33154, Z => n39426);
   U2598 : BUF_X2 port map( I => n21848, Z => n19517);
   U2600 : OR2_X1 port map( A1 => n21669, A2 => n21848, Z => n21850);
   U2603 : NAND2_X1 port map( A1 => n21902, A2 => n35921, ZN => n21422);
   U2604 : NOR2_X1 port map( A1 => n21577, A2 => n21594, ZN => n18784);
   U2617 : AND2_X1 port map( A1 => n20476, A2 => n14769, Z => n14577);
   U2618 : NAND2_X1 port map( A1 => n4094, A2 => n19262, ZN => n39368);
   U2628 : NAND2_X1 port map( A1 => n19084, A2 => n21944, ZN => n12752);
   U2630 : NAND3_X1 port map( A1 => n20277, A2 => n21928, A3 => n12044, ZN => 
                           n21728);
   U2631 : INV_X2 port map( I => n1157, ZN => n38546);
   U2633 : CLKBUF_X2 port map( I => n18467, Z => n5132);
   U2638 : AOI21_X2 port map( A1 => n35302, A2 => n31739, B => n23610, ZN => 
                           n31816);
   U2650 : NAND3_X2 port map( A1 => n30680, A2 => n19147, A3 => n19962, ZN => 
                           n32197);
   U2651 : NAND2_X2 port map( A1 => n30881, A2 => n388, ZN => n8362);
   U2654 : NAND2_X2 port map( A1 => n39305, A2 => n27449, ZN => n31708);
   U2656 : NAND2_X2 port map( A1 => n33091, A2 => n11344, ZN => n11277);
   U2658 : INV_X2 port map( I => n25691, ZN => n17271);
   U2663 : AOI22_X2 port map( A1 => n18562, A2 => n5220, B1 => n5219, B2 => 
                           n1221, ZN => n7680);
   U2664 : INV_X2 port map( I => n25351, ZN => n25614);
   U2667 : INV_X4 port map( I => n29241, ZN => n1062);
   U2668 : AND2_X1 port map( A1 => n16933, A2 => n15515, Z => n2246);
   U2670 : BUF_X4 port map( I => n32304, Z => n10702);
   U2677 : AND2_X1 port map( A1 => n15330, A2 => n20570, Z => n37124);
   U2679 : NOR2_X2 port map( A1 => n6443, A2 => n30153, ZN => n14520);
   U2680 : BUF_X4 port map( I => n30249, Z => n19663);
   U2682 : BUF_X4 port map( I => n20987, Z => n39320);
   U2690 : BUF_X2 port map( I => n29166, Z => n39798);
   U2692 : NOR2_X2 port map( A1 => n24526, A2 => n37106, ZN => n15169);
   U2693 : NAND2_X2 port map( A1 => n9265, A2 => n38719, ZN => n38718);
   U2694 : NAND2_X1 port map( A1 => n31652, A2 => n18231, ZN => n39234);
   U2695 : BUF_X2 port map( I => n8116, Z => n124);
   U2697 : BUF_X4 port map( I => n16080, Z => n36678);
   U2699 : BUF_X2 port map( I => n29174, Z => n30160);
   U2700 : NOR2_X2 port map( A1 => n28171, A2 => n28257, ZN => n27885);
   U2702 : INV_X4 port map( I => n25801, ZN => n1098);
   U2710 : OAI21_X2 port map( A1 => n854, A2 => n26697, B => n10736, ZN => 
                           n26698);
   U2714 : NAND2_X2 port map( A1 => n30587, A2 => n37432, ZN => n5459);
   U2715 : NOR2_X2 port map( A1 => n9310, A2 => n32870, ZN => n27368);
   U2716 : BUF_X2 port map( I => n30454, Z => n37319);
   U2717 : NAND3_X2 port map( A1 => n17176, A2 => n37298, A3 => n9957, ZN => 
                           n38697);
   U2718 : INV_X2 port map( I => n15368, ZN => n15421);
   U2719 : NAND2_X1 port map( A1 => n36485, A2 => n12425, ZN => n12424);
   U2725 : BUF_X2 port map( I => n11297, Z => n38491);
   U2728 : BUF_X2 port map( I => n6327, Z => n37629);
   U2731 : AOI21_X2 port map( A1 => n29182, A2 => n3986, B => n32894, ZN => 
                           n4072);
   U2732 : BUF_X4 port map( I => n32854, Z => n34307);
   U2733 : INV_X2 port map( I => n18785, ZN => n3965);
   U2738 : NAND2_X2 port map( A1 => n4525, A2 => n23610, ZN => n4527);
   U2739 : AOI21_X2 port map( A1 => n39159, A2 => n27288, B => n27069, ZN => 
                           n6010);
   U2740 : INV_X4 port map( I => n22324, ZN => n1683);
   U2742 : NOR2_X2 port map( A1 => n14705, A2 => n16449, ZN => n12772);
   U2743 : NAND2_X2 port map( A1 => n39065, A2 => n31433, ZN => n17661);
   U2744 : AOI22_X2 port map( A1 => n21359, A2 => n1158, B1 => n21666, B2 => 
                           n19620, ZN => n21362);
   U2745 : NAND2_X2 port map( A1 => n23056, A2 => n23160, ZN => n8758);
   U2746 : INV_X4 port map( I => n11150, ZN => n952);
   U2747 : INV_X2 port map( I => n33347, ZN => n28049);
   U2748 : OAI22_X2 port map( A1 => n29335, A2 => n29341, B1 => n18601, B2 => 
                           n16889, ZN => n29340);
   U2749 : NAND2_X2 port map( A1 => n37859, A2 => n37858, ZN => n37857);
   U2750 : INV_X2 port map( I => n33956, ZN => n27996);
   U2755 : AOI21_X2 port map( A1 => n9082, A2 => n18749, B => n27318, ZN => 
                           n3849);
   U2756 : BUF_X4 port map( I => n24034, Z => n1614);
   U2759 : BUF_X2 port map( I => n39443, Z => n37614);
   U2765 : INV_X2 port map( I => n197, ZN => n691);
   U2768 : INV_X4 port map( I => n23889, ZN => n17850);
   U2769 : INV_X2 port map( I => n4493, ZN => n39176);
   U2775 : BUF_X4 port map( I => n26031, Z => n37300);
   U2776 : INV_X2 port map( I => n13587, ZN => n22944);
   U2778 : NOR2_X2 port map( A1 => n13471, A2 => n35919, ZN => n16101);
   U2780 : OAI22_X2 port map( A1 => n26103, A2 => n18827, B1 => n1021, B2 => 
                           n17624, ZN => n5327);
   U2782 : BUF_X4 port map( I => n7106, Z => n269);
   U2784 : INV_X2 port map( I => n19318, ZN => n29664);
   U2786 : INV_X4 port map( I => n12478, ZN => n1531);
   U2787 : NOR2_X2 port map( A1 => n24788, A2 => n19255, ZN => n24609);
   U2791 : INV_X2 port map( I => n31433, ZN => n34359);
   U2792 : INV_X2 port map( I => n18433, ZN => n38604);
   U2796 : OR2_X2 port map( A1 => n4899, A2 => n34987, Z => n22886);
   U2797 : INV_X2 port map( I => n27564, ZN => n990);
   U2798 : NAND2_X2 port map( A1 => n4457, A2 => n36573, ZN => n19125);
   U2800 : NAND2_X2 port map( A1 => n12793, A2 => n4179, ZN => n22154);
   U2801 : INV_X2 port map( I => n35705, ZN => n38367);
   U2806 : NOR2_X2 port map( A1 => n36371, A2 => n21982, ZN => n21618);
   U2807 : AOI22_X2 port map( A1 => n22176, A2 => n32609, B1 => n20234, B2 => 
                           n21616, ZN => n2586);
   U2809 : INV_X2 port map( I => n17425, ZN => n19151);
   U2813 : OAI21_X2 port map( A1 => n1515, A2 => n37150, B => n17008, ZN => 
                           n39773);
   U2820 : NOR2_X2 port map( A1 => n24753, A2 => n6756, ZN => n24600);
   U2824 : INV_X1 port map( I => n37023, ZN => n3734);
   U2825 : NAND2_X2 port map( A1 => n13981, A2 => n29367, ZN => n15958);
   U2826 : NAND2_X2 port map( A1 => n11734, A2 => n5126, ZN => n2139);
   U2827 : AOI21_X2 port map( A1 => n23544, A2 => n17017, B => n32351, ZN => 
                           n23545);
   U2829 : NAND3_X2 port map( A1 => n35193, A2 => n4497, A3 => n4493, ZN => 
                           n4494);
   U2830 : INV_X2 port map( I => n2150, ZN => n39386);
   U2834 : INV_X2 port map( I => n21687, ZN => n38439);
   U2835 : NAND2_X2 port map( A1 => n23468, A2 => n3256, ZN => n7535);
   U2836 : BUF_X4 port map( I => n16631, Z => n1448);
   U2838 : NAND2_X2 port map( A1 => n5953, A2 => n1033, ZN => n17592);
   U2839 : NAND2_X2 port map( A1 => n26178, A2 => n26655, ZN => n32482);
   U2842 : INV_X2 port map( I => n22475, ZN => n22570);
   U2844 : NAND2_X1 port map( A1 => n18070, A2 => n15259, ZN => n15483);
   U2845 : NAND2_X1 port map( A1 => n29236, A2 => n29231, ZN => n15259);
   U2846 : OR2_X1 port map( A1 => n28715, A2 => n19844, Z => n28712);
   U2851 : BUF_X2 port map( I => n19844, Z => n33460);
   U2852 : NOR2_X1 port map( A1 => n33384, A2 => n25622, ZN => n33597);
   U2853 : CLKBUF_X4 port map( I => n11657, Z => n33384);
   U2855 : NOR2_X1 port map( A1 => n759, A2 => n28205, ZN => n7851);
   U2862 : NOR2_X1 port map( A1 => n1439, A2 => n28205, ZN => n39702);
   U2864 : INV_X1 port map( I => n30041, ZN => n1405);
   U2866 : NAND2_X1 port map( A1 => n16328, A2 => n30041, ZN => n4220);
   U2867 : CLKBUF_X4 port map( I => n29149, Z => n30041);
   U2871 : NAND2_X1 port map( A1 => n39686, A2 => n39420, ZN => n39567);
   U2873 : NAND2_X1 port map( A1 => n4387, A2 => n3820, ZN => n39420);
   U2875 : INV_X1 port map( I => n24040, ZN => n30321);
   U2876 : NAND2_X1 port map( A1 => n36824, A2 => n29171, ZN => n36170);
   U2878 : NAND2_X1 port map( A1 => n23392, A2 => n15642, ZN => n23242);
   U2880 : INV_X1 port map( I => n23392, ZN => n37528);
   U2883 : INV_X1 port map( I => n21813, ZN => n35026);
   U2884 : OAI22_X1 port map( A1 => n21813, A2 => n21682, B1 => n1350, B2 => 
                           n21684, ZN => n21375);
   U2888 : NOR2_X1 port map( A1 => n30196, A2 => n19693, ZN => n38255);
   U2889 : NOR3_X1 port map( A1 => n18261, A2 => n15248, A3 => n28109, ZN => 
                           n38374);
   U2891 : CLKBUF_X2 port map( I => n22968, Z => n45);
   U2894 : AOI22_X1 port map( A1 => n35250, A2 => n34055, B1 => n12782, B2 => 
                           n14211, ZN => n30960);
   U2901 : NOR2_X1 port map( A1 => n9385, A2 => n35250, ZN => n21049);
   U2904 : NAND2_X1 port map( A1 => n5077, A2 => n22008, ZN => n22214);
   U2908 : NOR2_X1 port map( A1 => n25616, A2 => n25574, ZN => n25420);
   U2909 : NAND2_X1 port map( A1 => n25574, A2 => n38625, ZN => n35419);
   U2911 : INV_X1 port map( I => n27470, ZN => n27761);
   U2912 : INV_X2 port map( I => n14858, ZN => n29338);
   U2915 : INV_X1 port map( I => n29501, ZN => n37374);
   U2916 : OAI21_X1 port map( A1 => n18374, A2 => n18743, B => n10677, ZN => 
                           n12108);
   U2917 : NAND2_X1 port map( A1 => n18374, A2 => n35051, ZN => n20150);
   U2920 : INV_X1 port map( I => n871, ZN => n36223);
   U2924 : AOI22_X1 port map( A1 => n18388, A2 => n33538, B1 => n18475, B2 => 
                           n7049, ZN => n36091);
   U2925 : AOI22_X1 port map( A1 => n1382, A2 => n30096, B1 => n14126, B2 => 
                           n30097, ZN => n30099);
   U2927 : CLKBUF_X2 port map( I => n9267, Z => n37890);
   U2933 : AOI22_X1 port map( A1 => n3470, A2 => n9295, B1 => n3469, B2 => 
                           n16042, ZN => n3468);
   U2939 : NAND2_X1 port map( A1 => n8372, A2 => n19352, ZN => n35424);
   U2950 : CLKBUF_X2 port map( I => n27095, Z => n32046);
   U2952 : NAND2_X1 port map( A1 => n14362, A2 => n3252, ZN => n37809);
   U2954 : NOR2_X1 port map( A1 => n6892, A2 => n12527, ZN => n10908);
   U2955 : NAND2_X1 port map( A1 => n11330, A2 => n6892, ZN => n28726);
   U2956 : INV_X1 port map( I => n13223, ZN => n27065);
   U2960 : NAND2_X1 port map( A1 => n13223, A2 => n34562, ZN => n12020);
   U2961 : BUF_X2 port map( I => n889, Z => n13851);
   U2965 : NAND3_X1 port map( A1 => n28189, A2 => n889, A3 => n16325, ZN => 
                           n13322);
   U2966 : OAI21_X1 port map( A1 => n39202, A2 => n32343, B => n11513, ZN => 
                           n31130);
   U2970 : NOR2_X1 port map( A1 => n26748, A2 => n26800, ZN => n2802);
   U2983 : INV_X1 port map( I => n31538, ZN => n31539);
   U2987 : AOI21_X1 port map( A1 => n28192, A2 => n9897, B => n9553, ZN => 
                           n15691);
   U2988 : NOR2_X1 port map( A1 => n9897, A2 => n17598, ZN => n33598);
   U2989 : INV_X2 port map( I => n20056, ZN => n17598);
   U2990 : NAND2_X1 port map( A1 => n27387, A2 => n2761, ZN => n27289);
   U2991 : NAND2_X1 port map( A1 => n11111, A2 => n4255, ZN => n35787);
   U2992 : NAND2_X1 port map( A1 => n30092, A2 => n30086, ZN => n29175);
   U2997 : INV_X1 port map( I => n30096, ZN => n30092);
   U3000 : NAND2_X1 port map( A1 => n18562, A2 => n19203, ZN => n13223);
   U3004 : INV_X2 port map( I => n27383, ZN => n18562);
   U3008 : AND2_X1 port map( A1 => n2522, A2 => n1891, Z => n37191);
   U3012 : OAI21_X1 port map( A1 => n35903, A2 => n9694, B => n25978, ZN => 
                           n31496);
   U3013 : NOR2_X1 port map( A1 => n1221, A2 => n27385, ZN => n13222);
   U3014 : CLKBUF_X1 port map( I => n15854, Z => n32571);
   U3015 : NAND2_X1 port map( A1 => n28657, A2 => n1197, ZN => n14605);
   U3018 : NOR2_X1 port map( A1 => n1197, A2 => n28560, ZN => n38681);
   U3019 : NAND2_X1 port map( A1 => n37592, A2 => n33383, ZN => n37591);
   U3021 : INV_X1 port map( I => n29067, ZN => n38087);
   U3022 : OR2_X1 port map( A1 => n13587, A2 => n20555, Z => n22974);
   U3024 : NAND2_X1 port map( A1 => n7096, A2 => n27131, ZN => n26889);
   U3031 : NAND2_X1 port map( A1 => n12689, A2 => n2150, ZN => n2152);
   U3032 : NAND2_X1 port map( A1 => n29212, A2 => n13762, ZN => n32267);
   U3034 : INV_X1 port map( I => n2139, ZN => n4868);
   U3036 : AOI21_X1 port map( A1 => n2139, A2 => n34745, B => n1103, ZN => 
                           n36387);
   U3038 : AOI22_X1 port map( A1 => n2760, A2 => n2761, B1 => n34769, B2 => 
                           n20871, ZN => n38873);
   U3040 : NOR2_X1 port map( A1 => n30484, A2 => n1211, ZN => n6733);
   U3041 : NAND2_X1 port map( A1 => n1211, A2 => n30484, ZN => n28032);
   U3042 : AOI21_X1 port map( A1 => n8206, A2 => n1211, B => n31808, ZN => 
                           n30962);
   U3043 : INV_X1 port map( I => n14980, ZN => n19765);
   U3045 : CLKBUF_X2 port map( I => n14980, Z => n9872);
   U3047 : NAND3_X1 port map( A1 => n34733, A2 => n35617, A3 => n2760, ZN => 
                           n35616);
   U3048 : OAI22_X1 port map( A1 => n9541, A2 => n18519, B1 => n18520, B2 => 
                           n19980, ZN => n9540);
   U3049 : NAND2_X1 port map( A1 => n19367, A2 => n18519, ZN => n18520);
   U3051 : NAND2_X1 port map( A1 => n38716, A2 => n18519, ZN => n4792);
   U3052 : NAND3_X1 port map( A1 => n3662, A2 => n36854, A3 => n32324, ZN => 
                           n32752);
   U3055 : NOR2_X1 port map( A1 => n7690, A2 => n3662, ZN => n6058);
   U3056 : NAND2_X1 port map( A1 => n38767, A2 => n4232, ZN => n4005);
   U3060 : NAND2_X1 port map( A1 => n34819, A2 => n28369, ZN => n38767);
   U3062 : INV_X2 port map( I => n2269, ZN => n29131);
   U3066 : AOI21_X1 port map( A1 => n37858, A2 => n37375, B => n37374, ZN => 
                           n30353);
   U3067 : INV_X2 port map( I => n17017, ZN => n1137);
   U3069 : NAND2_X1 port map( A1 => n17017, A2 => n23566, ZN => n23543);
   U3070 : NAND2_X1 port map( A1 => n6040, A2 => n39147, ZN => n6039);
   U3072 : NOR2_X1 port map( A1 => n12218, A2 => n14426, ZN => n5427);
   U3073 : CLKBUF_X1 port map( I => n30038, Z => n35103);
   U3075 : NAND3_X1 port map( A1 => n13006, A2 => n14997, A3 => n39603, ZN => 
                           n38371);
   U3076 : OAI21_X1 port map( A1 => n4882, A2 => n15615, B => n30177, ZN => 
                           n39603);
   U3077 : BUF_X1 port map( I => n35465, Z => n37095);
   U3081 : AOI21_X1 port map( A1 => n30255, A2 => n31529, B => n39234, ZN => 
                           n30256);
   U3082 : CLKBUF_X2 port map( I => n30262, Z => n31529);
   U3086 : AOI22_X1 port map( A1 => n19909, A2 => n29987, B1 => n29989, B2 => 
                           n31629, ZN => n16589);
   U3091 : AOI22_X1 port map( A1 => n907, A2 => n20018, B1 => n10451, B2 => 
                           n8918, ZN => n35541);
   U3095 : OAI22_X1 port map( A1 => n29176, A2 => n29175, B1 => n30099, B2 => 
                           n30087, ZN => n37935);
   U3096 : NAND3_X1 port map( A1 => n34621, A2 => n18431, A3 => n18070, ZN => 
                           n20559);
   U3097 : NAND2_X1 port map( A1 => n29351, A2 => n29385, ZN => n29080);
   U3098 : INV_X1 port map( I => n29384, ZN => n29351);
   U3101 : NAND2_X1 port map( A1 => n16663, A2 => n13605, ZN => n26643);
   U3103 : OAI21_X1 port map( A1 => n26933, A2 => n4411, B => n16663, ZN => 
                           n18946);
   U3104 : BUF_X2 port map( I => n15855, Z => n10587);
   U3106 : INV_X1 port map( I => n15855, ZN => n28699);
   U3110 : CLKBUF_X2 port map( I => n15855, Z => n38529);
   U3113 : NAND2_X1 port map( A1 => n33784, A2 => n30241, ZN => n7749);
   U3114 : NOR2_X1 port map( A1 => n17501, A2 => n26098, ZN => n25872);
   U3117 : INV_X1 port map( I => n26098, ZN => n25447);
   U3120 : OR2_X1 port map( A1 => n26098, A2 => n3874, Z => n25445);
   U3121 : NAND3_X1 port map( A1 => n33815, A2 => n26098, A3 => n31367, ZN => 
                           n32053);
   U3122 : NAND2_X1 port map( A1 => n26098, A2 => n10223, ZN => n39250);
   U3124 : OAI21_X1 port map( A1 => n26903, A2 => n26901, B => n26652, ZN => 
                           n17228);
   U3125 : INV_X1 port map( I => n26901, ZN => n39287);
   U3126 : NAND3_X1 port map( A1 => n34005, A2 => n26754, A3 => n26901, ZN => 
                           n26755);
   U3127 : CLKBUF_X4 port map( I => n29347, Z => n17225);
   U3134 : NOR2_X1 port map( A1 => n2059, A2 => n36788, ZN => n28538);
   U3136 : NOR2_X1 port map( A1 => n2059, A2 => n1434, ZN => n27457);
   U3145 : BUF_X1 port map( I => n8787, Z => n2059);
   U3146 : NOR3_X1 port map( A1 => n24266, A2 => n19745, A3 => n24267, ZN => 
                           n24029);
   U3147 : OR2_X1 port map( A1 => n39277, A2 => n14709, Z => n9020);
   U3148 : NAND2_X1 port map( A1 => n18398, A2 => n37809, ZN => n12046);
   U3149 : NOR2_X1 port map( A1 => n10346, A2 => n29586, ZN => n29629);
   U3154 : NAND2_X1 port map( A1 => n39018, A2 => n29810, ZN => n29799);
   U3156 : NAND2_X1 port map( A1 => n25924, A2 => n26027, ZN => n15377);
   U3157 : AOI22_X1 port map( A1 => n28657, A2 => n38681, B1 => n28442, B2 => 
                           n28559, ZN => n3050);
   U3158 : OAI22_X1 port map( A1 => n29904, A2 => n14600, B1 => n18222, B2 => 
                           n1407, ZN => n31356);
   U3159 : INV_X1 port map( I => n12940, ZN => n37914);
   U3166 : NAND2_X1 port map( A1 => n12940, A2 => n18667, ZN => n11597);
   U3169 : NOR2_X1 port map( A1 => n12940, A2 => n19783, ZN => n17794);
   U3170 : BUF_X2 port map( I => n33368, Z => n38580);
   U3172 : NOR2_X1 port map( A1 => n29630, A2 => n21269, ZN => n10081);
   U3174 : NOR2_X1 port map( A1 => n33784, A2 => n30796, ZN => n31238);
   U3175 : AND2_X1 port map( A1 => n30178, A2 => n12198, Z => n4882);
   U3178 : NAND2_X1 port map( A1 => n38407, A2 => n13757, ZN => n20635);
   U3180 : NAND3_X1 port map( A1 => n13757, A2 => n38407, A3 => n32345, ZN => 
                           n26626);
   U3181 : AOI22_X1 port map( A1 => n8761, A2 => n28882, B1 => n20085, B2 => 
                           n8762, ZN => n38698);
   U3182 : NOR2_X1 port map( A1 => n33482, A2 => n14417, ZN => n2294);
   U3187 : BUF_X1 port map( I => n29591, Z => n33482);
   U3190 : NAND2_X1 port map( A1 => n105, A2 => n29996, ZN => n21290);
   U3192 : NAND3_X1 port map( A1 => n33130, A2 => n841, A3 => n21042, ZN => 
                           n33304);
   U3195 : OAI21_X1 port map( A1 => n841, A2 => n12131, B => n25359, ZN => 
                           n10935);
   U3198 : NOR2_X1 port map( A1 => n5963, A2 => n3573, ZN => n6012);
   U3205 : INV_X2 port map( I => n15189, ZN => n38141);
   U3207 : NAND2_X1 port map( A1 => n29732, A2 => n29755, ZN => n29750);
   U3208 : NAND2_X1 port map( A1 => n4368, A2 => n20342, ZN => n30180);
   U3210 : NAND2_X1 port map( A1 => n39274, A2 => n29459, ZN => n37859);
   U3212 : AND2_X1 port map( A1 => n25867, A2 => n5859, Z => n25747);
   U3217 : NAND2_X1 port map( A1 => n25367, A2 => n25513, ZN => n15788);
   U3222 : NOR3_X1 port map( A1 => n25367, A2 => n25540, A3 => n30317, ZN => 
                           n16428);
   U3223 : INV_X2 port map( I => n25539, ZN => n25367);
   U3227 : AOI21_X1 port map( A1 => n29642, A2 => n30680, B => n37303, ZN => 
                           n29488);
   U3230 : NAND2_X1 port map( A1 => n7373, A2 => n37304, ZN => n37303);
   U3232 : INV_X1 port map( I => n28714, ZN => n17077);
   U3234 : NAND2_X1 port map( A1 => n1425, A2 => n31015, ZN => n28714);
   U3238 : NAND3_X1 port map( A1 => n35731, A2 => n15307, A3 => n15310, ZN => 
                           n17366);
   U3243 : NAND2_X1 port map( A1 => n14158, A2 => n19424, ZN => n29904);
   U3246 : NOR2_X1 port map( A1 => n8677, A2 => n14158, ZN => n10610);
   U3247 : INV_X1 port map( I => n9106, ZN => n34740);
   U3249 : INV_X1 port map( I => n26441, ZN => n38530);
   U3251 : NAND3_X1 port map( A1 => n28051, A2 => n11891, A3 => n28123, ZN => 
                           n17236);
   U3252 : OAI22_X1 port map( A1 => n29787, A2 => n15867, B1 => n29788, B2 => 
                           n29789, ZN => n37781);
   U3257 : NAND2_X1 port map( A1 => n30665, A2 => n34075, ZN => n12565);
   U3262 : CLKBUF_X2 port map( I => n30043, Z => n35809);
   U3265 : NOR2_X1 port map( A1 => n30042, A2 => n16328, ZN => n29898);
   U3267 : INV_X1 port map( I => n36827, ZN => n980);
   U3270 : NOR2_X1 port map( A1 => n8476, A2 => n36827, ZN => n28604);
   U3275 : NAND2_X1 port map( A1 => n8476, A2 => n36827, ZN => n10542);
   U3276 : NAND2_X1 port map( A1 => n27452, A2 => n15276, ZN => n40);
   U3277 : INV_X1 port map( I => n12350, ZN => n30139);
   U3279 : NAND3_X1 port map( A1 => n34180, A2 => n37565, A3 => n35858, ZN => 
                           n8996);
   U3289 : AOI21_X1 port map( A1 => n27822, A2 => n28257, B => n9880, ZN => 
                           n12529);
   U3290 : NAND2_X1 port map( A1 => n33928, A2 => n14940, ZN => n37545);
   U3292 : CLKBUF_X2 port map( I => n30233, Z => n14940);
   U3293 : OAI21_X1 port map( A1 => n36481, A2 => n30046, B => n29185, ZN => 
                           n36328);
   U3296 : BUF_X2 port map( I => n14559, Z => n36481);
   U3297 : OAI21_X1 port map( A1 => n30162, A2 => n29185, B => n36481, ZN => 
                           n28822);
   U3299 : NAND2_X1 port map( A1 => n30034, A2 => n30033, ZN => n30017);
   U3301 : NAND2_X1 port map( A1 => n30033, A2 => n30022, ZN => n30032);
   U3307 : NAND2_X1 port map( A1 => n30033, A2 => n8039, ZN => n30026);
   U3309 : INV_X1 port map( I => n38196, ZN => n37813);
   U3310 : CLKBUF_X2 port map( I => n19050, Z => n38196);
   U3311 : BUF_X2 port map( I => n19226, Z => n26764);
   U3313 : NOR2_X1 port map( A1 => n19349, A2 => n32002, ZN => n30334);
   U3315 : OAI21_X1 port map( A1 => n19497, A2 => n5067, B => n20672, ZN => 
                           n29668);
   U3317 : NAND2_X1 port map( A1 => n36471, A2 => n24802, ZN => n13748);
   U3319 : INV_X1 port map( I => n36471, ZN => n24804);
   U3321 : NAND2_X1 port map( A1 => n26097, A2 => n17700, ZN => n15618);
   U3322 : NOR2_X1 port map( A1 => n39305, A2 => n36969, ZN => n36762);
   U3324 : NOR2_X1 port map( A1 => n27265, A2 => n39305, ZN => n31934);
   U3325 : OAI21_X1 port map( A1 => n29597, A2 => n29595, B => n29596, ZN => 
                           n39006);
   U3327 : NAND2_X1 port map( A1 => n2292, A2 => n26959, ZN => n2100);
   U3328 : INV_X2 port map( I => n26959, ZN => n8651);
   U3329 : CLKBUF_X4 port map( I => n26959, Z => n30665);
   U3333 : AOI21_X1 port map( A1 => n29960, A2 => n29955, B => n29862, ZN => 
                           n17148);
   U3337 : NAND3_X1 port map( A1 => n29960, A2 => n19878, A3 => n29862, ZN => 
                           n29845);
   U3338 : INV_X1 port map( I => n5344, ZN => n37638);
   U3342 : NOR2_X1 port map( A1 => n865, A2 => n17535, ZN => n39202);
   U3344 : OAI22_X1 port map( A1 => n28714, A2 => n28715, B1 => n28712, B2 => 
                           n1193, ZN => n37862);
   U3347 : AOI21_X1 port map( A1 => n31015, A2 => n33460, B => n1193, ZN => 
                           n8216);
   U3349 : OAI22_X1 port map( A1 => n29533, A2 => n35180, B1 => n37605, B2 => 
                           n29536, ZN => n30645);
   U3350 : CLKBUF_X4 port map( I => n17730, Z => n5921);
   U3352 : AND2_X1 port map( A1 => n8293, A2 => n20361, Z => n7962);
   U3354 : OAI21_X1 port map( A1 => n38658, A2 => n34666, B => n30421, ZN => 
                           n24546);
   U3355 : INV_X1 port map( I => n34609, ZN => n1100);
   U3359 : INV_X1 port map( I => n13365, ZN => n7790);
   U3362 : NAND2_X1 port map( A1 => n32791, A2 => n9848, ZN => n17191);
   U3366 : INV_X1 port map( I => n9848, ZN => n27907);
   U3367 : BUF_X2 port map( I => n9848, Z => n39664);
   U3368 : NAND2_X1 port map( A1 => n26687, A2 => n17097, ZN => n11866);
   U3370 : NOR2_X1 port map( A1 => n28723, A2 => n28722, ZN => n15313);
   U3374 : NAND2_X1 port map( A1 => n38145, A2 => n28722, ZN => n28679);
   U3378 : CLKBUF_X2 port map( I => n29696, Z => n29763);
   U3380 : NAND2_X1 port map( A1 => n37349, A2 => n28637, ZN => n38818);
   U3385 : NAND2_X1 port map( A1 => n19115, A2 => n5009, ZN => n37349);
   U3388 : AOI22_X1 port map( A1 => n7048, A2 => n38535, B1 => n2175, B2 => 
                           n37463, ZN => n38025);
   U3389 : INV_X1 port map( I => n28262, ZN => n28257);
   U3393 : CLKBUF_X2 port map( I => n28262, Z => n3990);
   U3394 : BUF_X1 port map( I => n33967, Z => n31095);
   U3395 : CLKBUF_X4 port map( I => n15573, Z => n15447);
   U3400 : NAND2_X1 port map( A1 => n33972, A2 => n15033, ZN => n39153);
   U3403 : NAND2_X1 port map( A1 => n30056, A2 => n3818, ZN => n35095);
   U3405 : AND2_X1 port map( A1 => n29220, A2 => n18240, Z => n14421);
   U3408 : AOI21_X1 port map( A1 => n29870, A2 => n28, B => n29692, ZN => 
                           n29693);
   U3409 : INV_X2 port map( I => n29870, ZN => n33094);
   U3410 : NOR2_X1 port map( A1 => n10096, A2 => n29870, ZN => n32359);
   U3416 : OR2_X1 port map( A1 => n9214, A2 => n9235, Z => n26652);
   U3417 : AOI22_X1 port map( A1 => n38829, A2 => n33437, B1 => n30216, B2 => 
                           n38227, ZN => n38267);
   U3418 : OR2_X1 port map( A1 => n37013, A2 => n29005, Z => n5736);
   U3422 : INV_X1 port map( I => n25252, ZN => n38958);
   U3426 : CLKBUF_X4 port map( I => n30242, Z => n32415);
   U3427 : NAND2_X1 port map( A1 => n1068, A2 => n28676, ZN => n28576);
   U3428 : AOI21_X1 port map( A1 => n35199, A2 => n28591, B => n28676, ZN => 
                           n14701);
   U3429 : NOR2_X1 port map( A1 => n39126, A2 => n28141, ZN => n10756);
   U3432 : NOR2_X1 port map( A1 => n33405, A2 => n28141, ZN => n9655);
   U3440 : CLKBUF_X2 port map( I => n28141, Z => n39298);
   U3441 : NAND3_X1 port map( A1 => n30506, A2 => n35377, A3 => n36191, ZN => 
                           n23290);
   U3442 : BUF_X2 port map( I => n6640, Z => n200);
   U3444 : CLKBUF_X2 port map( I => n21792, Z => n16945);
   U3454 : NOR2_X1 port map( A1 => n2802, A2 => n2801, ZN => n8990);
   U3458 : NAND2_X1 port map( A1 => n29209, A2 => n11567, ZN => n9806);
   U3459 : NAND2_X1 port map( A1 => n37544, A2 => n14940, ZN => n14892);
   U3460 : NAND2_X1 port map( A1 => n1595, A2 => n19915, ZN => n15143);
   U3462 : OAI22_X1 port map( A1 => n26865, A2 => n39737, B1 => n39598, B2 => 
                           n36549, ZN => n16124);
   U3463 : NOR2_X1 port map( A1 => n39449, A2 => n36549, ZN => n10974);
   U3464 : NAND2_X1 port map( A1 => n17831, A2 => n18785, ZN => n3966);
   U3468 : CLKBUF_X4 port map( I => n28692, Z => n8349);
   U3469 : AOI21_X1 port map( A1 => n29185, A2 => n482, B => n1181, ZN => 
                           n11803);
   U3470 : INV_X2 port map( I => n7907, ZN => n30128);
   U3471 : CLKBUF_X2 port map( I => n7907, Z => n32508);
   U3476 : AND2_X1 port map( A1 => n39583, A2 => n27252, Z => n10581);
   U3482 : OR2_X1 port map( A1 => n27252, A2 => n39583, Z => n4105);
   U3483 : AND2_X1 port map( A1 => n5410, A2 => n8116, Z => n3133);
   U3484 : CLKBUF_X4 port map( I => n29568, Z => n29571);
   U3485 : NAND2_X1 port map( A1 => n9200, A2 => n33521, ZN => n30201);
   U3487 : NAND2_X1 port map( A1 => n28722, A2 => n28680, ZN => n2790);
   U3488 : NOR2_X1 port map( A1 => n13594, A2 => n28680, ZN => n28360);
   U3489 : CLKBUF_X4 port map( I => n15113, Z => n5093);
   U3494 : AOI21_X1 port map( A1 => n26847, A2 => n26614, B => n26849, ZN => 
                           n16941);
   U3495 : OAI21_X1 port map( A1 => n26847, A2 => n167, B => n26945, ZN => 
                           n34396);
   U3499 : INV_X2 port map( I => n14453, ZN => n26847);
   U3500 : INV_X2 port map( I => n15473, ZN => n28724);
   U3502 : NAND2_X1 port map( A1 => n37311, A2 => n15473, ZN => n28501);
   U3506 : NAND2_X1 port map( A1 => n4369, A2 => n28463, ZN => n28095);
   U3507 : NAND2_X1 port map( A1 => n19113, A2 => n28463, ZN => n19115);
   U3508 : AOI21_X1 port map( A1 => n30077, A2 => n3818, B => n31120, ZN => 
                           n6488);
   U3511 : NAND2_X1 port map( A1 => n31120, A2 => n30077, ZN => n39022);
   U3512 : INV_X2 port map( I => n28313, ZN => n1193);
   U3513 : NOR2_X1 port map( A1 => n28313, A2 => n19844, ZN => n28510);
   U3519 : NAND2_X1 port map( A1 => n22795, A2 => n35213, ZN => n16967);
   U3523 : CLKBUF_X2 port map( I => n22795, Z => n34457);
   U3525 : NAND2_X1 port map( A1 => n34014, A2 => n22795, ZN => n13688);
   U3526 : INV_X1 port map( I => n19384, ZN => n37882);
   U3527 : NOR2_X1 port map( A1 => n457, A2 => n39406, ZN => n34277);
   U3530 : NAND2_X1 port map( A1 => n39406, A2 => n9197, ZN => n33541);
   U3537 : AOI21_X1 port map( A1 => n9197, A2 => n39406, B => n39405, ZN => 
                           n37515);
   U3538 : NAND2_X1 port map( A1 => n31095, A2 => n14400, ZN => n29375);
   U3541 : NAND2_X1 port map( A1 => n14400, A2 => n9333, ZN => n38461);
   U3547 : INV_X2 port map( I => n4947, ZN => n6065);
   U3549 : NOR2_X1 port map( A1 => n4947, A2 => n1530, ZN => n7467);
   U3550 : NAND2_X1 port map( A1 => n2148, A2 => n4947, ZN => n4755);
   U3553 : NAND2_X1 port map( A1 => n3053, A2 => n3052, ZN => n34291);
   U3554 : OAI21_X1 port map( A1 => n4284, A2 => n1419, B => n34695, ZN => 
                           n3053);
   U3558 : CLKBUF_X2 port map( I => n5638, Z => n5471);
   U3559 : INV_X1 port map( I => n28465, ZN => n39365);
   U3560 : OAI21_X1 port map( A1 => n28639, A2 => n33046, B => n28465, ZN => 
                           n31030);
   U3562 : NAND2_X1 port map( A1 => n11389, A2 => n9955, ZN => n5645);
   U3563 : INV_X1 port map( I => n18004, ZN => n15591);
   U3564 : OR2_X1 port map( A1 => n14000, A2 => n18903, Z => n18904);
   U3566 : NAND2_X1 port map( A1 => n20429, A2 => n13261, ZN => n32987);
   U3567 : INV_X1 port map( I => n28638, ZN => n19113);
   U3578 : NAND2_X1 port map( A1 => n28638, A2 => n28464, ZN => n28465);
   U3579 : NAND2_X1 port map( A1 => n15573, A2 => n28638, ZN => n5009);
   U3580 : NAND2_X1 port map( A1 => n20453, A2 => n30186, ZN => n34344);
   U3583 : OAI21_X1 port map( A1 => n23469, A2 => n32930, B => n36448, ZN => 
                           n39670);
   U3584 : AOI22_X1 port map( A1 => n30417, A2 => n36448, B1 => n8680, B2 => 
                           n37839, ZN => n39333);
   U3586 : NOR2_X1 port map( A1 => n23645, A2 => n36448, ZN => n4634);
   U3587 : CLKBUF_X2 port map( I => n8026, Z => n35590);
   U3589 : OAI21_X1 port map( A1 => n29309, A2 => n31279, B => n6262, ZN => 
                           n39134);
   U3592 : AOI21_X1 port map( A1 => n18031, A2 => n25614, B => n2721, ZN => 
                           n36434);
   U3595 : CLKBUF_X4 port map( I => n26249, Z => n26970);
   U3596 : NAND2_X1 port map( A1 => n26876, A2 => n26249, ZN => n15124);
   U3598 : CLKBUF_X1 port map( I => n18186, Z => n5062);
   U3600 : NAND2_X1 port map( A1 => n23181, A2 => n22903, ZN => n20957);
   U3601 : AOI22_X1 port map( A1 => n15040, A2 => n15039, B1 => n18851, B2 => 
                           n23181, ZN => n31319);
   U3604 : NAND2_X1 port map( A1 => n28659, A2 => n31663, ZN => n28437);
   U3605 : INV_X1 port map( I => n28437, ZN => n28438);
   U3607 : NOR2_X1 port map( A1 => n28437, A2 => n28554, ZN => n35000);
   U3608 : AOI21_X1 port map( A1 => n17031, A2 => n3538, B => n28742, ZN => 
                           n11474);
   U3609 : NAND2_X1 port map( A1 => n11506, A2 => n29437, ZN => n12321);
   U3612 : NOR2_X1 port map( A1 => n1392, A2 => n29437, ZN => n14414);
   U3616 : OR2_X1 port map( A1 => n1812, A2 => n34475, Z => n15229);
   U3618 : INV_X1 port map( I => n7506, ZN => n1268);
   U3622 : NOR2_X1 port map( A1 => n7506, A2 => n24903, ZN => n24904);
   U3628 : NAND2_X1 port map( A1 => n19050, A2 => n33963, ZN => n4805);
   U3629 : NOR2_X1 port map( A1 => n33288, A2 => n20889, ZN => n20355);
   U3631 : NAND2_X1 port map( A1 => n16398, A2 => n209, ZN => n31643);
   U3632 : OAI21_X1 port map( A1 => n36465, A2 => n13404, B => n37898, ZN => 
                           n32524);
   U3633 : NAND2_X1 port map( A1 => n37898, A2 => n974, ZN => n28340);
   U3634 : AOI21_X1 port map( A1 => n19005, A2 => n33864, B => n23380, ZN => 
                           n6518);
   U3636 : INV_X1 port map( I => n11125, ZN => n33278);
   U3640 : NOR2_X1 port map( A1 => n34652, A2 => n7141, ZN => n37274);
   U3641 : AOI21_X1 port map( A1 => n28050, A2 => n28124, B => n14404, ZN => 
                           n27152);
   U3649 : INV_X2 port map( I => n14404, ZN => n983);
   U3651 : AOI22_X1 port map( A1 => n9660, A2 => n33697, B1 => n22902, B2 => 
                           n36369, ZN => n12130);
   U3654 : AOI22_X1 port map( A1 => n5982, A2 => n30883, B1 => n5981, B2 => 
                           n3345, ZN => n31630);
   U3655 : NAND2_X1 port map( A1 => n3345, A2 => n37997, ZN => n26237);
   U3656 : NAND2_X1 port map( A1 => n9694, A2 => n3345, ZN => n35947);
   U3657 : NAND2_X1 port map( A1 => n37997, A2 => n3345, ZN => n37996);
   U3658 : INV_X2 port map( I => n34265, ZN => n3345);
   U3659 : AOI21_X1 port map( A1 => n17857, A2 => n2906, B => n7044, ZN => 
                           n2905);
   U3662 : NAND2_X1 port map( A1 => n7044, A2 => n34011, ZN => n2904);
   U3668 : NOR2_X1 port map( A1 => n34011, A2 => n7044, ZN => n24601);
   U3669 : NAND2_X1 port map( A1 => n7044, A2 => n32882, ZN => n3044);
   U3670 : OAI21_X1 port map( A1 => n27377, A2 => n8137, B => n6445, ZN => 
                           n27381);
   U3671 : NAND2_X1 port map( A1 => n39153, A2 => n34131, ZN => n15452);
   U3678 : OAI21_X1 port map( A1 => n27998, A2 => n18061, B => n11461, ZN => 
                           n8524);
   U3681 : NAND2_X1 port map( A1 => n28200, A2 => n18061, ZN => n37322);
   U3682 : NOR2_X1 port map( A1 => n1022, A2 => n25695, ZN => n31131);
   U3684 : NAND2_X1 port map( A1 => n34424, A2 => n33579, ZN => n34422);
   U3685 : NOR3_X1 port map( A1 => n33579, A2 => n2192, A3 => n37107, ZN => 
                           n37439);
   U3686 : CLKBUF_X2 port map( I => n11753, Z => n37951);
   U3687 : OAI21_X1 port map( A1 => n6902, A2 => n6901, B => n4573, ZN => n6900
                           );
   U3688 : AOI21_X1 port map( A1 => n4573, A2 => n640, B => n33554, ZN => 
                           n37750);
   U3691 : OAI21_X1 port map( A1 => n4573, A2 => n640, B => n1318, ZN => n39297
                           );
   U3694 : NAND2_X1 port map( A1 => n25829, A2 => n2830, ZN => n6097);
   U3696 : INV_X2 port map( I => n18017, ZN => n25692);
   U3697 : NOR2_X1 port map( A1 => n19914, A2 => n1006, ZN => n11305);
   U3698 : OAI21_X1 port map( A1 => n1493, A2 => n14458, B => n19914, ZN => 
                           n5746);
   U3699 : NAND2_X1 port map( A1 => n13491, A2 => n281, ZN => n27935);
   U3702 : NOR2_X1 port map( A1 => n281, A2 => n12663, ZN => n13059);
   U3704 : NAND3_X1 port map( A1 => n32354, A2 => n8380, A3 => n8381, ZN => 
                           n5622);
   U3706 : INV_X1 port map( I => n32354, ZN => n37270);
   U3707 : NOR2_X1 port map( A1 => n19782, A2 => n24465, ZN => n24251);
   U3708 : OAI21_X1 port map( A1 => n24465, A2 => n24467, B => n18347, ZN => 
                           n24158);
   U3717 : NOR2_X1 port map( A1 => n18348, A2 => n24465, ZN => n7361);
   U3718 : NAND2_X1 port map( A1 => n35903, A2 => n4553, ZN => n26034);
   U3720 : NOR2_X1 port map( A1 => n26838, A2 => n1092, ZN => n3093);
   U3723 : OAI22_X1 port map( A1 => n24351, A2 => n9921, B1 => n3487, B2 => 
                           n18653, ZN => n12643);
   U3724 : AOI21_X1 port map( A1 => n5957, A2 => n18653, B => n24770, ZN => 
                           n13428);
   U3726 : NAND2_X1 port map( A1 => n18653, A2 => n3487, ZN => n39182);
   U3727 : NAND2_X1 port map( A1 => n26219, A2 => n1494, ZN => n20547);
   U3728 : NAND2_X1 port map( A1 => n9268, A2 => n11162, ZN => n8601);
   U3729 : AOI21_X1 port map( A1 => n26953, A2 => n11162, B => n30768, ZN => 
                           n11463);
   U3737 : NAND2_X1 port map( A1 => n27508, A2 => n998, ZN => n11162);
   U3741 : AOI21_X1 port map( A1 => n33935, A2 => n22129, B => n8245, ZN => 
                           n17778);
   U3743 : OAI21_X1 port map( A1 => n12630, A2 => n33935, B => n7496, ZN => 
                           n7495);
   U3745 : AOI21_X1 port map( A1 => n6366, A2 => n33935, B => n1831, ZN => 
                           n7496);
   U3746 : NAND2_X1 port map( A1 => n1831, A2 => n33935, ZN => n22909);
   U3748 : NOR2_X1 port map( A1 => n16463, A2 => n33935, ZN => n37517);
   U3751 : NOR3_X1 port map( A1 => n28023, A2 => n6643, A3 => n16065, ZN => 
                           n32150);
   U3752 : INV_X2 port map( I => n16065, ZN => n989);
   U3753 : AOI22_X1 port map( A1 => n15669, A2 => n26852, B1 => n15668, B2 => 
                           n167, ZN => n15667);
   U3754 : NOR2_X1 port map( A1 => n26852, A2 => n38797, ZN => n39257);
   U3755 : BUF_X2 port map( I => n26852, Z => n15670);
   U3756 : OAI21_X1 port map( A1 => n11432, A2 => n27337, B => n11431, ZN => 
                           n26890);
   U3757 : NAND2_X1 port map( A1 => n39417, A2 => n4886, ZN => n27218);
   U3759 : INV_X1 port map( I => n39417, ZN => n35745);
   U3761 : NAND2_X1 port map( A1 => n27069, A2 => n39417, ZN => n6013);
   U3764 : NAND2_X1 port map( A1 => n38097, A2 => n2741, ZN => n14203);
   U3765 : CLKBUF_X4 port map( I => n4378, Z => n3818);
   U3766 : INV_X1 port map( I => n17184, ZN => n17395);
   U3767 : CLKBUF_X2 port map( I => n17184, Z => n38714);
   U3769 : NAND2_X1 port map( A1 => n35523, A2 => n38327, ZN => n38056);
   U3770 : AND2_X1 port map( A1 => n5530, A2 => n29284, Z => n6843);
   U3774 : NAND3_X1 port map( A1 => n30258, A2 => n11700, A3 => n19663, ZN => 
                           n31652);
   U3775 : INV_X1 port map( I => n26660, ZN => n26697);
   U3777 : CLKBUF_X4 port map( I => n15423, Z => n8757);
   U3779 : NAND2_X1 port map( A1 => n6357, A2 => n30464, ZN => n18653);
   U3780 : OAI21_X1 port map( A1 => n13170, A2 => n35357, B => n5465, ZN => 
                           n8635);
   U3782 : NAND2_X1 port map( A1 => n35357, A2 => n19759, ZN => n31347);
   U3783 : AOI22_X1 port map( A1 => n33577, A2 => n28812, B1 => n28764, B2 => 
                           n35357, ZN => n32376);
   U3786 : OAI21_X1 port map( A1 => n28808, A2 => n35357, B => n31542, ZN => 
                           n35083);
   U3787 : NAND3_X1 port map( A1 => n30292, A2 => n35357, A3 => n28764, ZN => 
                           n33675);
   U3790 : OAI21_X1 port map( A1 => n30161, A2 => n30162, B => n1400, ZN => 
                           n11429);
   U3793 : NAND2_X1 port map( A1 => n11125, A2 => n30161, ZN => n39686);
   U3796 : OAI21_X1 port map( A1 => n2522, A2 => n35919, B => n38414, ZN => 
                           n3996);
   U3799 : CLKBUF_X2 port map( I => n4771, Z => n39448);
   U3800 : AND2_X1 port map( A1 => n8412, A2 => n4771, Z => n16144);
   U3801 : AND3_X1 port map( A1 => n27440, A2 => n27438, A3 => n4771, Z => n161
                           );
   U3804 : INV_X1 port map( I => n4771, ZN => n13992);
   U3811 : OR2_X1 port map( A1 => n4771, A2 => n27438, Z => n11638);
   U3815 : INV_X2 port map( I => n13650, ZN => n34184);
   U3817 : AOI21_X1 port map( A1 => n603, A2 => n32691, B => n25912, ZN => 
                           n32056);
   U3819 : AOI21_X1 port map( A1 => n32691, A2 => n25912, B => n32690, ZN => 
                           n32689);
   U3820 : CLKBUF_X2 port map( I => n12572, Z => n7892);
   U3821 : NOR2_X1 port map( A1 => n9444, A2 => n28533, ZN => n9443);
   U3824 : NOR2_X1 port map( A1 => n8727, A2 => n29851, ZN => n37390);
   U3828 : OAI21_X1 port map( A1 => n2969, A2 => n32168, B => n32559, ZN => 
                           n2968);
   U3830 : NAND2_X1 port map( A1 => n31716, A2 => n27049, ZN => n12745);
   U3837 : INV_X1 port map( I => n27049, ZN => n54);
   U3841 : OAI22_X1 port map( A1 => n38611, A2 => n14739, B1 => n20788, B2 => 
                           n23610, ZN => n4528);
   U3842 : INV_X1 port map( I => n856, ZN => n17158);
   U3843 : BUF_X2 port map( I => n856, Z => n11138);
   U3845 : NOR2_X1 port map( A1 => n27405, A2 => n27155, ZN => n32853);
   U3846 : OAI21_X1 port map( A1 => n29310, A2 => n12880, B => n10422, ZN => 
                           n12879);
   U3847 : AND2_X1 port map( A1 => n29384, A2 => n10422, Z => n35966);
   U3849 : OR3_X1 port map( A1 => n11084, A2 => n36426, A3 => n10422, Z => 
                           n1822);
   U3850 : INV_X1 port map( I => n11383, ZN => n37721);
   U3852 : NOR3_X1 port map( A1 => n24473, A2 => n15461, A3 => n39309, ZN => 
                           n33085);
   U3862 : CLKBUF_X1 port map( I => n24473, Z => n37916);
   U3866 : BUF_X2 port map( I => n36894, Z => n34829);
   U3869 : BUF_X2 port map( I => n9918, Z => n39576);
   U3873 : NOR2_X1 port map( A1 => n29940, A2 => n9918, ZN => n29939);
   U3874 : NAND2_X1 port map( A1 => n29940, A2 => n9918, ZN => n9143);
   U3877 : NOR2_X1 port map( A1 => n32854, A2 => n13305, ZN => n16367);
   U3878 : NAND2_X1 port map( A1 => n4805, A2 => n6938, ZN => n31025);
   U3885 : INV_X1 port map( I => n10739, ZN => n13691);
   U3887 : NAND2_X1 port map( A1 => n10739, A2 => n19389, ZN => n7820);
   U3888 : NAND2_X1 port map( A1 => n23506, A2 => n23580, ZN => n13833);
   U3890 : NAND2_X1 port map( A1 => n18453, A2 => n7023, ZN => n34819);
   U3898 : CLKBUF_X2 port map( I => n7023, Z => n1432);
   U3908 : NAND2_X1 port map( A1 => n13424, A2 => n209, ZN => n7849);
   U3913 : NAND2_X1 port map( A1 => n14752, A2 => n38491, ZN => n27013);
   U3914 : CLKBUF_X2 port map( I => n14752, Z => n7619);
   U3915 : BUF_X2 port map( I => Key(47), Z => n30169);
   U3917 : INV_X1 port map( I => n16989, ZN => n3733);
   U3918 : INV_X2 port map( I => n3840, ZN => n14027);
   U3922 : NAND2_X1 port map( A1 => n3840, A2 => n18303, ZN => n16989);
   U3929 : AND2_X1 port map( A1 => n3840, A2 => n1338, Z => n1778);
   U3930 : OR2_X1 port map( A1 => n5028, A2 => n28729, Z => n14497);
   U3934 : INV_X1 port map( I => n28729, ZN => n15649);
   U3935 : INV_X1 port map( I => n28729, ZN => n38998);
   U3940 : NAND2_X1 port map( A1 => n21770, A2 => n21768, ZN => n21605);
   U3946 : CLKBUF_X4 port map( I => n21768, Z => n19546);
   U3947 : NOR2_X1 port map( A1 => n21768, A2 => n21770, ZN => n16052);
   U3953 : INV_X2 port map( I => n21768, ZN => n19084);
   U3954 : CLKBUF_X2 port map( I => n9501, Z => n31721);
   U3955 : INV_X1 port map( I => n9501, ZN => n10563);
   U3956 : NAND2_X1 port map( A1 => n425, A2 => n25894, ZN => n5276);
   U3957 : BUF_X2 port map( I => n25894, Z => n30900);
   U3962 : INV_X2 port map( I => n25894, ZN => n1103);
   U3964 : NOR2_X1 port map( A1 => n15677, A2 => n25894, ZN => n25738);
   U3971 : NAND3_X1 port map( A1 => n28383, A2 => n20494, A3 => n31855, ZN => 
                           n28384);
   U3972 : NAND2_X1 port map( A1 => n31854, A2 => n31855, ZN => n30636);
   U3977 : NAND2_X1 port map( A1 => n29675, A2 => n29683, ZN => n29682);
   U3980 : INV_X1 port map( I => n29683, ZN => n29677);
   U3983 : OR2_X1 port map( A1 => n21885, A2 => n15839, Z => n13858);
   U3986 : NOR2_X1 port map( A1 => n18246, A2 => n11729, ZN => n37703);
   U3987 : NAND3_X1 port map( A1 => n9699, A2 => n8569, A3 => n20309, ZN => 
                           n22830);
   U3989 : NAND2_X1 port map( A1 => n20309, A2 => n19000, ZN => n22934);
   U3990 : INV_X2 port map( I => n20313, ZN => n24172);
   U3993 : NAND2_X1 port map( A1 => n20312, A2 => n20313, ZN => n263);
   U3995 : INV_X2 port map( I => n36840, ZN => n7588);
   U4005 : AOI22_X1 port map( A1 => n27255, A2 => n36840, B1 => n18716, B2 => 
                           n18195, ZN => n27256);
   U4014 : NAND2_X1 port map( A1 => n36840, A2 => n39583, ZN => n27049);
   U4017 : NAND2_X1 port map( A1 => n15911, A2 => n962, ZN => n38001);
   U4024 : OAI21_X1 port map( A1 => n8942, A2 => n962, B => n5581, ZN => n5582)
                           ;
   U4026 : INV_X2 port map( I => n14415, ZN => n1094);
   U4027 : NOR2_X1 port map( A1 => n14415, A2 => n14380, ZN => n34249);
   U4034 : AOI21_X1 port map( A1 => n11636, A2 => n14415, B => n8413, ZN => 
                           n8917);
   U4036 : OAI21_X1 port map( A1 => n39415, A2 => n21043, B => n7658, ZN => 
                           n4128);
   U4037 : OAI22_X1 port map( A1 => n1034, A2 => n24425, B1 => n17456, B2 => 
                           n21043, ZN => n298);
   U4053 : OAI21_X1 port map( A1 => n21043, A2 => n38561, B => n17456, ZN => 
                           n31252);
   U4057 : NAND2_X1 port map( A1 => n21043, A2 => n37580, ZN => n17062);
   U4061 : NAND2_X1 port map( A1 => n20643, A2 => n19518, ZN => n33015);
   U4063 : INV_X1 port map( I => n35376, ZN => n23730);
   U4065 : AOI21_X1 port map( A1 => n24738, A2 => n31722, B => n24737, ZN => 
                           n35128);
   U4069 : NAND2_X1 port map( A1 => n31722, A2 => n31679, ZN => n16671);
   U4071 : NAND2_X1 port map( A1 => n23535, A2 => n14759, ZN => n23227);
   U4072 : NOR2_X1 port map( A1 => n14759, A2 => n23535, ZN => n20100);
   U4074 : INV_X1 port map( I => n14759, ZN => n23538);
   U4075 : NAND2_X1 port map( A1 => n3907, A2 => n22113, ZN => n10154);
   U4077 : NAND3_X1 port map( A1 => n1049, A2 => n3907, A3 => n38448, ZN => 
                           n11456);
   U4078 : NAND3_X1 port map( A1 => n10930, A2 => n13191, A3 => n3907, ZN => 
                           n38484);
   U4080 : CLKBUF_X2 port map( I => n6285, Z => n33656);
   U4081 : INV_X1 port map( I => n18160, ZN => n5564);
   U4083 : AND2_X2 port map( A1 => n37922, A2 => n38229, Z => n37062);
   U4088 : INV_X1 port map( I => n10482, ZN => n14089);
   U4091 : INV_X2 port map( I => n4574, ZN => n39527);
   U4096 : AND3_X1 port map( A1 => n15455, A2 => n1046, A3 => n20267, Z => 
                           n37063);
   U4097 : CLKBUF_X4 port map( I => n4524, Z => n38408);
   U4099 : INV_X2 port map( I => n4524, ZN => n38611);
   U4104 : INV_X2 port map( I => n15299, ZN => n32424);
   U4105 : OR2_X2 port map( A1 => n7577, A2 => n15299, Z => n37064);
   U4114 : INV_X2 port map( I => n15933, ZN => n24394);
   U4115 : AND2_X1 port map( A1 => n24090, A2 => n24442, Z => n37066);
   U4116 : AND2_X2 port map( A1 => n33616, A2 => n39191, Z => n37067);
   U4119 : NAND2_X2 port map( A1 => n31143, A2 => n39731, ZN => n25085);
   U4120 : OR2_X1 port map( A1 => n25513, A2 => n25540, Z => n37069);
   U4122 : INV_X2 port map( I => n17624, ZN => n32193);
   U4124 : AND3_X1 port map( A1 => n178, A2 => n25359, A3 => n33130, Z => 
                           n37070);
   U4125 : AND2_X1 port map( A1 => n25367, A2 => n25540, Z => n37071);
   U4126 : INV_X2 port map( I => n25288, ZN => n25989);
   U4130 : CLKBUF_X4 port map( I => n25288, Z => n38548);
   U4131 : INV_X1 port map( I => n17803, ZN => n17951);
   U4133 : BUF_X4 port map( I => n17803, Z => n38168);
   U4136 : AND2_X1 port map( A1 => n9859, A2 => n25887, Z => n37073);
   U4137 : OR2_X2 port map( A1 => n38939, A2 => n38755, Z => n37075);
   U4140 : INV_X4 port map( I => n13973, ZN => n1891);
   U4141 : INV_X2 port map( I => n36050, ZN => n38690);
   U4142 : OR2_X1 port map( A1 => n27292, A2 => n6191, Z => n37077);
   U4143 : INV_X2 port map( I => n19995, ZN => n37754);
   U4144 : BUF_X2 port map( I => n27910, Z => n580);
   U4146 : OR2_X1 port map( A1 => n19541, A2 => n5525, Z => n37078);
   U4151 : XOR2_X1 port map( A1 => n3206, A2 => n35438, Z => n37079);
   U4160 : INV_X4 port map( I => n7063, ZN => n39724);
   U4161 : INV_X2 port map( I => n5028, ZN => n30805);
   U4168 : INV_X1 port map( I => n14448, ZN => n154);
   U4170 : OR2_X2 port map( A1 => n28748, A2 => n28622, Z => n37080);
   U4173 : AND2_X2 port map( A1 => n32077, A2 => n6264, Z => n37081);
   U4177 : NAND2_X2 port map( A1 => n2868, A2 => n39112, ZN => n35657);
   U4178 : INV_X2 port map( I => n20673, ZN => n19992);
   U4181 : CLKBUF_X4 port map( I => n20673, Z => n481);
   U4188 : NAND2_X2 port map( A1 => n2784, A2 => n2789, ZN => n38147);
   U4189 : OR2_X2 port map( A1 => n35551, A2 => n18288, Z => n37083);
   U4190 : NAND2_X1 port map( A1 => n17861, A2 => n20255, ZN => n21972);
   U4195 : INV_X2 port map( I => n20255, ZN => n20996);
   U4199 : BUF_X2 port map( I => n20255, Z => n7613);
   U4201 : AND2_X2 port map( A1 => n11573, A2 => n30221, Z => n9708);
   U4204 : OR2_X2 port map( A1 => n20541, A2 => n30221, Z => n30225);
   U4206 : OR2_X2 port map( A1 => n14833, A2 => n5796, Z => n5795);
   U4211 : CLKBUF_X4 port map( I => n9387, Z => n32039);
   U4212 : AOI21_X1 port map( A1 => n21726, A2 => n21727, B => n18293, ZN => 
                           n18979);
   U4218 : INV_X2 port map( I => n15868, ZN => n18408);
   U4223 : NOR2_X1 port map( A1 => n22274, A2 => n15868, ZN => n15280);
   U4224 : NAND2_X1 port map( A1 => n39059, A2 => n36908, ZN => n24687);
   U4227 : OAI22_X1 port map( A1 => n33151, A2 => n14265, B1 => n39059, B2 => 
                           n36908, ZN => n8296);
   U4233 : OR2_X2 port map( A1 => n33230, A2 => n36908, Z => n37999);
   U4237 : OR2_X2 port map( A1 => n7067, A2 => n7066, Z => n31290);
   U4240 : NOR2_X2 port map( A1 => n22146, A2 => n22240, ZN => n22145);
   U4241 : CLKBUF_X12 port map( I => n734, Z => n35216);
   U4247 : CLKBUF_X12 port map( I => n734, Z => n7583);
   U4251 : INV_X2 port map( I => n29497, ZN => n2954);
   U4252 : NAND2_X1 port map( A1 => n29389, A2 => n29497, ZN => n39274);
   U4256 : OAI21_X1 port map( A1 => n29389, A2 => n19151, B => n29497, ZN => 
                           n15876);
   U4257 : NAND2_X1 port map( A1 => n29459, A2 => n29497, ZN => n29501);
   U4258 : NOR2_X1 port map( A1 => n5127, A2 => n18929, ZN => n10092);
   U4264 : INV_X2 port map( I => n18929, ZN => n6128);
   U4275 : INV_X2 port map( I => n10047, ZN => n15455);
   U4276 : INV_X1 port map( I => n35431, ZN => n22299);
   U4279 : OAI21_X1 port map( A1 => n2341, A2 => n19422, B => n1029, ZN => 
                           n20929);
   U4282 : INV_X1 port map( I => n19422, ZN => n1576);
   U4283 : INV_X1 port map( I => n31367, ZN => n950);
   U4286 : NAND3_X1 port map( A1 => n24416, A2 => n37355, A3 => n31213, ZN => 
                           n17979);
   U4287 : INV_X2 port map( I => n24416, ZN => n19679);
   U4296 : CLKBUF_X4 port map( I => n24366, Z => n32683);
   U4297 : INV_X2 port map( I => n24366, ZN => n9135);
   U4299 : NAND2_X1 port map( A1 => n24366, A2 => n37107, ZN => n34424);
   U4303 : NOR2_X1 port map( A1 => n2084, A2 => n2085, ZN => n33775);
   U4305 : BUF_X2 port map( I => n37047, Z => n36556);
   U4310 : INV_X1 port map( I => n37047, ZN => n24426);
   U4315 : AND2_X2 port map( A1 => n29377, A2 => n20726, Z => n34973);
   U4316 : OR2_X2 port map( A1 => n36357, A2 => n39456, Z => n39535);
   U4317 : AND2_X2 port map( A1 => n33510, A2 => n36357, Z => n10288);
   U4318 : AND2_X2 port map( A1 => n20669, A2 => n12012, Z => n33633);
   U4321 : INV_X1 port map( I => n21848, ZN => n6198);
   U4322 : OAI22_X1 port map( A1 => n2643, A2 => n19133, B1 => n21944, B2 => 
                           n21605, ZN => n38836);
   U4323 : OR2_X2 port map( A1 => n5656, A2 => n10455, Z => n12245);
   U4325 : NAND2_X1 port map( A1 => n18850, A2 => n38704, ZN => n32013);
   U4326 : NAND2_X1 port map( A1 => n18850, A2 => n23310, ZN => n23606);
   U4327 : INV_X1 port map( I => n18850, ZN => n1636);
   U4329 : NAND2_X1 port map( A1 => n33168, A2 => n18998, ZN => n15852);
   U4330 : INV_X1 port map( I => n33168, ZN => n32457);
   U4331 : AOI21_X1 port map( A1 => n20376, A2 => n33168, B => n7131, ZN => 
                           n21977);
   U4332 : NOR2_X1 port map( A1 => n9422, A2 => n33168, ZN => n7216);
   U4336 : INV_X1 port map( I => n20662, ZN => n28532);
   U4339 : NAND2_X1 port map( A1 => n24565, A2 => n32637, ZN => n24566);
   U4341 : AND3_X2 port map( A1 => n24557, A2 => n24812, A3 => n32637, Z => 
                           n39713);
   U4344 : NAND2_X1 port map( A1 => n32637, A2 => n24565, ZN => n36618);
   U4345 : OAI22_X1 port map( A1 => n7878, A2 => n10158, B1 => n19637, B2 => 
                           n19636, ZN => n7877);
   U4346 : OAI21_X1 port map( A1 => n19637, A2 => n4048, B => n25387, ZN => 
                           n17231);
   U4347 : INV_X1 port map( I => n19637, ZN => n1255);
   U4352 : CLKBUF_X12 port map( I => n9824, Z => n36683);
   U4354 : AND2_X2 port map( A1 => n20194, A2 => n25694, Z => n25195);
   U4356 : CLKBUF_X4 port map( I => n6355, Z => n4743);
   U4357 : OAI21_X1 port map( A1 => n21923, A2 => n9316, B => n21924, ZN => 
                           n38898);
   U4358 : CLKBUF_X12 port map( I => n13039, Z => n37084);
   U4359 : INV_X1 port map( I => n32230, ZN => n4956);
   U4367 : BUF_X2 port map( I => n32230, Z => n32122);
   U4368 : OAI22_X1 port map( A1 => n19382, A2 => n1595, B1 => n545, B2 => 
                           n1276, ZN => n37967);
   U4369 : NAND2_X1 port map( A1 => n1276, A2 => n5985, ZN => n24102);
   U4370 : INV_X1 port map( I => n19112, ZN => n21257);
   U4373 : CLKBUF_X12 port map( I => n2145, Z => n38468);
   U4375 : INV_X1 port map( I => n3213, ZN => n6543);
   U4378 : INV_X2 port map( I => n22484, ZN => n33415);
   U4379 : CLKBUF_X4 port map( I => n21214, Z => n7916);
   U4380 : OR2_X1 port map( A1 => n24600, A2 => n18788, Z => n9073);
   U4381 : BUF_X2 port map( I => n16489, Z => n11696);
   U4383 : INV_X1 port map( I => n26435, ZN => n10878);
   U4386 : INV_X1 port map( I => n20423, ZN => n32427);
   U4387 : AND2_X1 port map( A1 => n20423, A2 => n19867, Z => n18587);
   U4392 : NOR2_X1 port map( A1 => n26972, A2 => n20423, ZN => n26815);
   U4393 : NAND2_X1 port map( A1 => n20423, A2 => n858, ZN => n15980);
   U4399 : INV_X1 port map( I => n18549, ZN => n37487);
   U4400 : NAND2_X1 port map( A1 => n19203, A2 => n18549, ZN => n19352);
   U4401 : NAND2_X1 port map( A1 => n27383, A2 => n18549, ZN => n36797);
   U4403 : NOR2_X1 port map( A1 => n1221, A2 => n18549, ZN => n27026);
   U4405 : CLKBUF_X12 port map( I => n18507, Z => n37085);
   U4407 : CLKBUF_X12 port map( I => n6347, Z => n39010);
   U4411 : INV_X1 port map( I => n6347, ZN => n2818);
   U4414 : NAND2_X1 port map( A1 => n7644, A2 => n4576, ZN => n19389);
   U4416 : NAND2_X1 port map( A1 => n7379, A2 => n7644, ZN => n31662);
   U4420 : NAND2_X1 port map( A1 => n33287, A2 => n7644, ZN => n16126);
   U4422 : NAND2_X2 port map( A1 => n21479, A2 => n2157, ZN => n2156);
   U4432 : CLKBUF_X12 port map( I => n38839, Z => n37803);
   U4435 : INV_X2 port map( I => n38839, ZN => n38302);
   U4437 : BUF_X2 port map( I => n15299, Z => n6638);
   U4438 : INV_X1 port map( I => n3003, ZN => n20799);
   U4446 : BUF_X2 port map( I => n3003, Z => n31407);
   U4453 : NAND2_X1 port map( A1 => n36058, A2 => n13300, ZN => n24605);
   U4454 : INV_X2 port map( I => n26229, ZN => n34495);
   U4455 : NAND2_X1 port map( A1 => n4149, A2 => n17887, ZN => n5371);
   U4460 : OR2_X2 port map( A1 => n19594, A2 => n35246, Z => n4340);
   U4461 : NOR2_X1 port map( A1 => n19966, A2 => n19594, ZN => n22793);
   U4463 : INV_X1 port map( I => n26048, ZN => n1242);
   U4468 : NOR2_X1 port map( A1 => n26048, A2 => n1524, ZN => n5475);
   U4469 : BUF_X2 port map( I => n37232, Z => n37086);
   U4471 : OAI21_X1 port map( A1 => n4147, A2 => n12790, B => n36263, ZN => 
                           n31951);
   U4476 : NAND2_X1 port map( A1 => n27133, A2 => n1225, ZN => n31734);
   U4478 : NAND2_X1 port map( A1 => n5027, A2 => n27133, ZN => n10066);
   U4480 : INV_X1 port map( I => n36750, ZN => n15909);
   U4485 : CLKBUF_X12 port map( I => n36750, Z => n39116);
   U4488 : AOI22_X1 port map( A1 => n37985, A2 => n30764, B1 => n9656, B2 => 
                           n24591, ZN => n819);
   U4490 : INV_X2 port map( I => n30764, ZN => n958);
   U4493 : NAND2_X1 port map( A1 => n878, A2 => n33956, ZN => n27900);
   U4499 : CLKBUF_X12 port map( I => n33956, Z => n310);
   U4500 : INV_X1 port map( I => n5274, ZN => n16663);
   U4502 : INV_X2 port map( I => n9802, ZN => n1015);
   U4504 : NAND2_X1 port map( A1 => n9802, A2 => n33997, ZN => n32035);
   U4508 : AOI22_X1 port map( A1 => n1015, A2 => n25860, B1 => n362, B2 => 
                           n9802, ZN => n12712);
   U4509 : NOR2_X1 port map( A1 => n1520, A2 => n9802, ZN => n37309);
   U4510 : OAI21_X1 port map( A1 => n14881, A2 => n31006, B => n35895, ZN => 
                           n14795);
   U4512 : OR2_X2 port map( A1 => n37662, A2 => n25636, Z => n25717);
   U4516 : CLKBUF_X2 port map( I => n25636, Z => n9132);
   U4517 : CLKBUF_X12 port map( I => n33847, Z => n37087);
   U4518 : BUF_X4 port map( I => n33847, Z => n37088);
   U4523 : INV_X1 port map( I => n10782, ZN => n20820);
   U4532 : OAI22_X1 port map( A1 => n38211, A2 => n8251, B1 => n8253, B2 => 
                           n1082, ZN => n2380);
   U4534 : AND2_X2 port map( A1 => n25481, A2 => n19928, Z => n20565);
   U4536 : INV_X1 port map( I => n7497, ZN => n6451);
   U4541 : NOR2_X1 port map( A1 => n1151, A2 => n7497, ZN => n5876);
   U4542 : INV_X1 port map( I => n8972, ZN => n37995);
   U4543 : AOI22_X1 port map( A1 => n2837, A2 => n26030, B1 => n25923, B2 => 
                           n25962, ZN => n38102);
   U4545 : OR2_X2 port map( A1 => n19478, A2 => n25553, Z => n25477);
   U4548 : OR2_X1 port map( A1 => n19992, A2 => n29781, Z => n19993);
   U4552 : INV_X1 port map( I => n25163, ZN => n10273);
   U4554 : NOR2_X1 port map( A1 => n1097, A2 => n4604, ZN => n3359);
   U4556 : NAND2_X1 port map( A1 => n4604, A2 => n38416, ZN => n25768);
   U4557 : BUF_X2 port map( I => n4604, Z => n34402);
   U4559 : CLKBUF_X12 port map( I => n24403, Z => n37904);
   U4560 : OAI22_X1 port map( A1 => n1032, A2 => n39055, B1 => n13555, B2 => 
                           n24403, ZN => n33727);
   U4563 : NAND2_X1 port map( A1 => n24403, A2 => n13443, ZN => n12366);
   U4564 : AND3_X2 port map( A1 => n20517, A2 => n24403, A3 => n13555, Z => 
                           n33500);
   U4566 : NAND2_X1 port map( A1 => n22240, A2 => n21214, ZN => n22147);
   U4567 : INV_X1 port map( I => n22240, ZN => n21821);
   U4571 : NAND2_X1 port map( A1 => n9387, A2 => n10820, ZN => n20034);
   U4576 : INV_X2 port map( I => n30210, ZN => n30214);
   U4577 : NAND2_X1 port map( A1 => n21802, A2 => n8899, ZN => n22075);
   U4588 : OR2_X2 port map( A1 => n20397, A2 => n8899, Z => n3269);
   U4589 : INV_X2 port map( I => n15515, ZN => n25527);
   U4593 : NOR2_X1 port map( A1 => n39415, A2 => n9193, ZN => n38349);
   U4594 : NAND3_X2 port map( A1 => n7472, A2 => n7471, A3 => n27149, ZN => 
                           n38277);
   U4598 : AOI22_X1 port map( A1 => n50, A2 => n14448, B1 => n28732, B2 => 
                           n36623, ZN => n15321);
   U4599 : NOR2_X1 port map( A1 => n7712, A2 => n31612, ZN => n23425);
   U4605 : INV_X1 port map( I => n31612, ZN => n7008);
   U4608 : BUF_X2 port map( I => n31612, Z => n4600);
   U4610 : NOR2_X1 port map( A1 => n12331, A2 => n14817, ZN => n22992);
   U4611 : INV_X2 port map( I => n12331, ZN => n6674);
   U4613 : NAND2_X1 port map( A1 => n22865, A2 => n12331, ZN => n16638);
   U4626 : NAND2_X1 port map( A1 => n31744, A2 => n21248, ZN => n32546);
   U4629 : INV_X2 port map( I => n13029, ZN => n23350);
   U4634 : NAND2_X1 port map( A1 => n6590, A2 => n26109, ZN => n14229);
   U4635 : INV_X2 port map( I => n6590, ZN => n951);
   U4636 : NOR2_X1 port map( A1 => n6590, A2 => n26109, ZN => n37462);
   U4642 : NOR2_X1 port map( A1 => n23303, A2 => n11970, ZN => n23420);
   U4646 : OR2_X1 port map( A1 => n29939, A2 => n1057, Z => n34086);
   U4648 : CLKBUF_X12 port map( I => n28179, Z => n18832);
   U4661 : INV_X1 port map( I => n28873, ZN => n33715);
   U4663 : INV_X1 port map( I => n8003, ZN => n39725);
   U4664 : OAI22_X1 port map( A1 => n29571, A2 => n31899, B1 => n1393, B2 => 
                           n17262, ZN => n29577);
   U4666 : OAI21_X1 port map( A1 => n30629, A2 => n17400, B => n25975, ZN => 
                           n17002);
   U4667 : AOI22_X1 port map( A1 => n5311, A2 => n27407, B1 => n27153, B2 => 
                           n27406, ZN => n5085);
   U4669 : AOI22_X1 port map( A1 => n27153, A2 => n27407, B1 => n2947, B2 => 
                           n1487, ZN => n27405);
   U4674 : NAND2_X1 port map( A1 => n17714, A2 => n28729, ZN => n38123);
   U4683 : NAND2_X1 port map( A1 => n36623, A2 => n28729, ZN => n36633);
   U4689 : OAI21_X1 port map( A1 => n28178, A2 => n28031, B => n16559, ZN => 
                           n20084);
   U4696 : OR2_X2 port map( A1 => n27964, A2 => n33960, Z => n21322);
   U4698 : AND2_X2 port map( A1 => n33960, A2 => n27964, Z => n4640);
   U4701 : NAND2_X1 port map( A1 => n13995, A2 => n2047, ZN => n23146);
   U4703 : NOR2_X1 port map( A1 => n13995, A2 => n2047, ZN => n23044);
   U4705 : INV_X2 port map( I => n13995, ZN => n37791);
   U4708 : NOR2_X1 port map( A1 => n23145, A2 => n13995, ZN => n23148);
   U4710 : NOR2_X1 port map( A1 => n27325, A2 => n35500, ZN => n17985);
   U4712 : NAND2_X1 port map( A1 => n17142, A2 => n27325, ZN => n37512);
   U4718 : NAND3_X1 port map( A1 => n11910, A2 => n17142, A3 => n27325, ZN => 
                           n38734);
   U4719 : AOI21_X1 port map( A1 => n12326, A2 => n27325, B => n11910, ZN => 
                           n27329);
   U4720 : NOR2_X1 port map( A1 => n12326, A2 => n27325, ZN => n4253);
   U4721 : INV_X1 port map( I => n29041, ZN => n5992);
   U4722 : INV_X1 port map( I => n26125, ZN => n39661);
   U4723 : NOR2_X1 port map( A1 => n14126, A2 => n30097, ZN => n2489);
   U4724 : OAI21_X1 port map( A1 => n32682, A2 => n38172, B => n9686, ZN => 
                           n4871);
   U4726 : INV_X2 port map( I => n9686, ZN => n28736);
   U4730 : NAND2_X1 port map( A1 => n9686, A2 => n17234, ZN => n28547);
   U4731 : INV_X1 port map( I => n21754, ZN => n21699);
   U4732 : NAND2_X1 port map( A1 => n14493, A2 => n21754, ZN => n21542);
   U4733 : BUF_X2 port map( I => n21754, Z => n1372);
   U4734 : NAND2_X1 port map( A1 => n26063, A2 => n25943, ZN => n35679);
   U4735 : INV_X2 port map( I => n3874, ZN => n4699);
   U4738 : NAND2_X1 port map( A1 => n31367, A2 => n3874, ZN => n25870);
   U4739 : NAND2_X1 port map( A1 => n3669, A2 => n3874, ZN => n17700);
   U4745 : NAND3_X1 port map( A1 => n15577, A2 => n27305, A3 => n27304, ZN => 
                           n10735);
   U4747 : OAI21_X1 port map( A1 => n27305, A2 => n17166, B => n35906, ZN => 
                           n12072);
   U4748 : INV_X1 port map( I => n22669, ZN => n35810);
   U4749 : OR2_X2 port map( A1 => n20896, A2 => n34120, Z => n12323);
   U4750 : INV_X2 port map( I => n27438, ZN => n19719);
   U4754 : INV_X1 port map( I => n38981, ZN => n23321);
   U4757 : CLKBUF_X4 port map( I => n38981, Z => n16047);
   U4758 : AOI21_X1 port map( A1 => n7424, A2 => n17072, B => n14881, ZN => 
                           n14796);
   U4760 : AOI21_X1 port map( A1 => n7426, A2 => n34959, B => n3708, ZN => 
                           n7425);
   U4761 : NOR2_X2 port map( A1 => n37070, A2 => n9482, ZN => n9479);
   U4762 : INV_X1 port map( I => n26364, ZN => n26366);
   U4764 : BUF_X2 port map( I => n26765, Z => n26922);
   U4765 : OAI22_X1 port map( A1 => n26765, A2 => n13543, B1 => n19371, B2 => 
                           n3606, ZN => n39758);
   U4766 : INV_X2 port map( I => n180, ZN => n1420);
   U4767 : NAND2_X1 port map( A1 => n28616, A2 => n180, ZN => n28615);
   U4769 : NOR2_X1 port map( A1 => n6147, A2 => n14126, ZN => n20099);
   U4771 : NOR2_X1 port map( A1 => n30092, A2 => n6147, ZN => n37356);
   U4772 : NAND2_X1 port map( A1 => n6147, A2 => n31601, ZN => n7600);
   U4776 : INV_X1 port map( I => n28972, ZN => n4314);
   U4777 : NOR2_X1 port map( A1 => n3434, A2 => n25800, ZN => n32233);
   U4779 : NOR2_X1 port map( A1 => n20031, A2 => n9862, ZN => n2453);
   U4787 : NAND2_X1 port map( A1 => n12952, A2 => n1145, ZN => n38513);
   U4791 : NAND3_X1 port map( A1 => n8260, A2 => n8261, A3 => n7542, ZN => 
                           n37696);
   U4798 : NAND2_X1 port map( A1 => n15135, A2 => n10171, ZN => n27305);
   U4799 : INV_X2 port map( I => n10171, ZN => n35332);
   U4802 : INV_X1 port map( I => n10611, ZN => n25037);
   U4804 : AND3_X1 port map( A1 => n1021, A2 => n17624, A3 => n11148, Z => 
                           n25781);
   U4807 : OR2_X1 port map( A1 => n11148, A2 => n15575, Z => n37213);
   U4813 : OAI22_X1 port map( A1 => n29723, A2 => n29717, B1 => n29710, B2 => 
                           n29709, ZN => n32519);
   U4814 : NOR2_X1 port map( A1 => n29723, A2 => n5951, ZN => n39101);
   U4816 : AND2_X2 port map( A1 => n22879, A2 => n5891, Z => n6009);
   U4820 : OR2_X2 port map( A1 => n22879, A2 => n5891, Z => n12032);
   U4821 : CLKBUF_X12 port map( I => n3116, Z => n37092);
   U4822 : BUF_X2 port map( I => n3116, Z => n37093);
   U4827 : AOI21_X1 port map( A1 => n38068, A2 => n4192, B => n27446, ZN => 
                           n32940);
   U4833 : NAND2_X1 port map( A1 => n27446, A2 => n38187, ZN => n5630);
   U4836 : INV_X1 port map( I => n17351, ZN => n17350);
   U4839 : CLKBUF_X12 port map( I => n11627, Z => n531);
   U4843 : NAND2_X1 port map( A1 => n23566, A2 => n3713, ZN => n5792);
   U4849 : CLKBUF_X4 port map( I => n33734, Z => n2192);
   U4857 : INV_X1 port map( I => n33734, ZN => n4243);
   U4858 : INV_X1 port map( I => n21488, ZN => n19699);
   U4860 : NAND2_X1 port map( A1 => n2765, A2 => n8679, ZN => n22144);
   U4866 : INV_X4 port map( I => n1812, ZN => n18253);
   U4872 : OAI21_X1 port map( A1 => n38973, A2 => n39059, B => n33230, ZN => 
                           n8355);
   U4875 : NAND2_X1 port map( A1 => n36908, A2 => n33230, ZN => n13554);
   U4876 : NAND2_X1 port map( A1 => n33230, A2 => n24761, ZN => n14338);
   U4881 : INV_X2 port map( I => n23482, ZN => n6303);
   U4891 : CLKBUF_X4 port map( I => n23482, Z => n9078);
   U4893 : OAI21_X1 port map( A1 => n1630, A2 => n38244, B => n23586, ZN => 
                           n34585);
   U4897 : INV_X2 port map( I => n12617, ZN => n38244);
   U4900 : AND3_X2 port map( A1 => n38976, A2 => n22196, A3 => n30800, Z => 
                           n14269);
   U4901 : OAI22_X1 port map( A1 => n38976, A2 => n1327, B1 => n8520, B2 => 
                           n22287, ZN => n5557);
   U4902 : INV_X2 port map( I => n38976, ZN => n1328);
   U4904 : OAI21_X1 port map( A1 => n5396, A2 => n39227, B => n13598, ZN => 
                           n5397);
   U4906 : INV_X1 port map( I => n19370, ZN => n21517);
   U4920 : CLKBUF_X12 port map( I => n19370, Z => n17534);
   U4923 : OR3_X2 port map( A1 => n20207, A2 => n9945, A3 => n24116, Z => n4687
                           );
   U4924 : AND2_X2 port map( A1 => n24287, A2 => n20207, Z => n11132);
   U4926 : AOI21_X1 port map( A1 => n14423, A2 => n4239, B => n34813, ZN => 
                           n2907);
   U4936 : OR2_X2 port map( A1 => n20449, A2 => n12100, Z => n22990);
   U4940 : AND2_X2 port map( A1 => n3861, A2 => n2858, Z => n29852);
   U4944 : INV_X1 port map( I => n17758, ZN => n26319);
   U4946 : NOR2_X1 port map( A1 => n18502, A2 => n29438, ZN => n17293);
   U4948 : NOR2_X1 port map( A1 => n29439, A2 => n29438, ZN => n29433);
   U4952 : INV_X1 port map( I => n31944, ZN => n23450);
   U4954 : NAND2_X1 port map( A1 => n31944, A2 => n11678, ZN => n23394);
   U4956 : AND2_X2 port map( A1 => n11585, A2 => n11586, Z => n18193);
   U4958 : NAND3_X1 port map( A1 => n21847, A2 => n19392, A3 => n21668, ZN => 
                           n16653);
   U4959 : AOI21_X1 port map( A1 => n19517, A2 => n18219, B => n21847, ZN => 
                           n6101);
   U4966 : NOR2_X1 port map( A1 => n20538, A2 => n20342, ZN => n2466);
   U4970 : NAND2_X1 port map( A1 => n5450, A2 => n4424, ZN => n3681);
   U4972 : AOI21_X1 port map( A1 => n2480, A2 => n5450, B => n18567, ZN => 
                           n4045);
   U4975 : NAND2_X1 port map( A1 => n5450, A2 => n14833, ZN => n22256);
   U4976 : INV_X1 port map( I => n5450, ZN => n22063);
   U4981 : NOR3_X1 port map( A1 => n16094, A2 => n23477, A3 => n23473, ZN => 
                           n17388);
   U4986 : NAND2_X1 port map( A1 => n16094, A2 => n1139, ZN => n12870);
   U4990 : NAND2_X1 port map( A1 => n34558, A2 => n16094, ZN => n23475);
   U4991 : OR2_X2 port map( A1 => n36442, A2 => n16094, Z => n8432);
   U5004 : NAND2_X1 port map( A1 => n25583, A2 => n24896, ZN => n20295);
   U5007 : INV_X1 port map( I => n25191, ZN => n34788);
   U5023 : NAND3_X1 port map( A1 => n28812, A2 => n33577, A3 => n19759, ZN => 
                           n8913);
   U5025 : OR2_X2 port map( A1 => n9845, A2 => n28231, Z => n27970);
   U5029 : OR2_X2 port map( A1 => n10216, A2 => n33786, Z => n8027);
   U5031 : INV_X2 port map( I => n37016, ZN => n32045);
   U5032 : INV_X1 port map( I => n9916, ZN => n14132);
   U5036 : CLKBUF_X12 port map( I => n22223, Z => n39284);
   U5040 : BUF_X4 port map( I => n21814, Z => n19768);
   U5047 : CLKBUF_X12 port map( I => n29005, Z => n621);
   U5052 : INV_X1 port map( I => n18399, ZN => n33243);
   U5053 : CLKBUF_X12 port map( I => n13794, Z => n36426);
   U5059 : OAI21_X1 port map( A1 => n31845, A2 => n39268, B => n24618, ZN => 
                           n39562);
   U5060 : NAND2_X1 port map( A1 => n37624, A2 => n39268, ZN => n24534);
   U5063 : AOI21_X1 port map( A1 => n31845, A2 => n39268, B => n1026, ZN => 
                           n6187);
   U5076 : NAND2_X1 port map( A1 => n25813, A2 => n33909, ZN => n35671);
   U5080 : INV_X1 port map( I => n25813, ZN => n32510);
   U5083 : BUF_X4 port map( I => n22623, Z => n37094);
   U5084 : CLKBUF_X4 port map( I => n24053, Z => n38813);
   U5087 : NAND2_X1 port map( A1 => n28463, A2 => n28464, ZN => n1815);
   U5093 : INV_X2 port map( I => n28464, ZN => n28637);
   U5099 : NAND3_X1 port map( A1 => n38600, A2 => n34558, A3 => n36442, ZN => 
                           n22681);
   U5101 : INV_X1 port map( I => n36442, ZN => n20343);
   U5102 : NAND2_X1 port map( A1 => n36442, A2 => n23473, ZN => n11186);
   U5103 : CLKBUF_X4 port map( I => n26272, Z => n26979);
   U5106 : NAND2_X1 port map( A1 => n37341, A2 => n12633, ZN => n39343);
   U5107 : OAI22_X1 port map( A1 => n33151, A2 => n12633, B1 => n14857, B2 => 
                           n36908, ZN => n13002);
   U5117 : INV_X1 port map( I => n17583, ZN => n14968);
   U5127 : NAND2_X1 port map( A1 => n17583, A2 => n28330, ZN => n17031);
   U5128 : OR2_X2 port map( A1 => n5732, A2 => n962, Z => n8769);
   U5133 : AND2_X2 port map( A1 => n8628, A2 => n5732, Z => n8508);
   U5136 : BUF_X1 port map( I => n21885, Z => n36754);
   U5146 : NOR3_X1 port map( A1 => n34977, A2 => n27211, A3 => n8412, ZN => 
                           n36407);
   U5149 : NAND2_X1 port map( A1 => n19719, A2 => n8412, ZN => n27097);
   U5150 : CLKBUF_X4 port map( I => n8412, Z => n7494);
   U5168 : NAND2_X1 port map( A1 => n7852, A2 => n36082, ZN => n24768);
   U5175 : AND2_X1 port map( A1 => n7852, A2 => n24764, Z => n39099);
   U5183 : OAI22_X1 port map( A1 => n21591, A2 => n21592, B1 => n38480, B2 => 
                           n21576, ZN => n20585);
   U5184 : NOR3_X1 port map( A1 => n8735, A2 => n37934, A3 => n24406, ZN => 
                           n37551);
   U5186 : INV_X1 port map( I => n6756, ZN => n30534);
   U5191 : AOI21_X1 port map( A1 => n24126, A2 => n19484, B => n6756, ZN => 
                           n24127);
   U5192 : NOR2_X1 port map( A1 => n23516, A2 => n23517, ZN => n2175);
   U5198 : OAI22_X1 port map( A1 => n7049, A2 => n18475, B1 => n23516, B2 => 
                           n39001, ZN => n38024);
   U5202 : OR2_X2 port map( A1 => n12950, A2 => n35954, Z => n24206);
   U5209 : CLKBUF_X12 port map( I => n17397, Z => n33646);
   U5210 : NAND2_X1 port map( A1 => n17397, A2 => n28207, ZN => n28361);
   U5224 : INV_X2 port map( I => n17397, ZN => n28723);
   U5225 : BUF_X4 port map( I => n35465, Z => n37096);
   U5228 : INV_X1 port map( I => n34685, ZN => n25857);
   U5232 : NOR2_X1 port map( A1 => n34685, A2 => n10404, ZN => n34206);
   U5234 : AND3_X2 port map( A1 => n15796, A2 => n25849, A3 => n34685, Z => 
                           n12063);
   U5240 : CLKBUF_X12 port map( I => n18211, Z => n5021);
   U5241 : NAND2_X1 port map( A1 => n24765, A2 => n24764, ZN => n24766);
   U5242 : AND2_X2 port map( A1 => n26195, A2 => n35750, Z => n14667);
   U5244 : NAND2_X1 port map( A1 => n35750, A2 => n5089, ZN => n34842);
   U5248 : OR2_X2 port map( A1 => n26643, A2 => n26932, Z => n26547);
   U5251 : NAND3_X1 port map( A1 => n33352, A2 => n26933, A3 => n26932, ZN => 
                           n33383);
   U5254 : INV_X1 port map( I => n26932, ZN => n35912);
   U5258 : AND2_X2 port map( A1 => n26932, A2 => n37235, Z => n14485);
   U5260 : BUF_X1 port map( I => n26818, Z => n19353);
   U5266 : NAND2_X1 port map( A1 => n10404, A2 => n25887, ZN => n26072);
   U5273 : NOR2_X1 port map( A1 => n9859, A2 => n25887, ZN => n26071);
   U5274 : OAI22_X1 port map( A1 => n23342, A2 => n23430, B1 => n15787, B2 => 
                           n23343, ZN => n1829);
   U5281 : NAND2_X1 port map( A1 => n1628, A2 => n23430, ZN => n3506);
   U5288 : NOR2_X1 port map( A1 => n9685, A2 => n22092, ZN => n22094);
   U5289 : NAND2_X1 port map( A1 => n1152, A2 => n22092, ZN => n22205);
   U5292 : NOR2_X1 port map( A1 => n4190, A2 => n6904, ZN => n17645);
   U5293 : OAI21_X1 port map( A1 => n6904, A2 => n26125, B => n5098, ZN => 
                           n38783);
   U5294 : NAND3_X1 port map( A1 => n39454, A2 => n6904, A3 => n4516, ZN => 
                           n26010);
   U5296 : NAND2_X1 port map( A1 => n39826, A2 => n27389, ZN => n27167);
   U5309 : CLKBUF_X12 port map( I => n19478, Z => n31580);
   U5311 : BUF_X2 port map( I => n25418, Z => n19495);
   U5314 : NOR2_X1 port map( A1 => n35260, A2 => n25418, ZN => n25597);
   U5317 : AOI21_X1 port map( A1 => n10623, A2 => n3840, B => n3086, ZN => 
                           n3085);
   U5318 : INV_X2 port map( I => n23076, ZN => n23181);
   U5322 : CLKBUF_X12 port map( I => n26668, Z => n19331);
   U5323 : INV_X1 port map( I => n26668, ZN => n26973);
   U5324 : AND2_X2 port map( A1 => n38901, A2 => n26668, Z => n33006);
   U5327 : NAND2_X1 port map( A1 => n26178, A2 => n26701, ZN => n4641);
   U5329 : NOR2_X1 port map( A1 => n23076, A2 => n23077, ZN => n787);
   U5331 : NOR2_X1 port map( A1 => n33933, A2 => n23076, ZN => n9841);
   U5336 : NOR2_X1 port map( A1 => n15641, A2 => n39424, ZN => n21109);
   U5339 : NOR2_X1 port map( A1 => n27221, A2 => n39424, ZN => n4627);
   U5341 : INV_X1 port map( I => n39424, ZN => n39531);
   U5346 : AOI21_X1 port map( A1 => n27292, A2 => n39424, B => n5588, ZN => 
                           n4700);
   U5347 : NAND2_X1 port map( A1 => n28748, A2 => n28622, ZN => n28747);
   U5348 : INV_X2 port map( I => n28622, ZN => n34244);
   U5349 : NAND2_X1 port map( A1 => n24829, A2 => n24802, ZN => n10161);
   U5350 : NOR2_X1 port map( A1 => n24829, A2 => n38194, ZN => n24572);
   U5358 : NAND2_X1 port map( A1 => n2018, A2 => n24829, ZN => n10160);
   U5360 : INV_X1 port map( I => n17405, ZN => n5266);
   U5369 : INV_X4 port map( I => n29617, ZN => n35405);
   U5370 : NAND2_X1 port map( A1 => n28681, A2 => n28720, ZN => n2788);
   U5378 : NOR2_X1 port map( A1 => n28720, A2 => n28722, ZN => n37560);
   U5382 : INV_X1 port map( I => n28720, ZN => n28721);
   U5383 : AND2_X2 port map( A1 => n862, A2 => n867, Z => n13489);
   U5387 : CLKBUF_X4 port map( I => n867, Z => n2451);
   U5388 : NAND2_X1 port map( A1 => n32046, A2 => n32566, ZN => n38068);
   U5391 : INV_X1 port map( I => n32566, ZN => n16782);
   U5398 : INV_X1 port map( I => n15135, ZN => n27586);
   U5400 : BUF_X2 port map( I => n15135, Z => n4781);
   U5405 : NAND3_X1 port map( A1 => n16181, A2 => n16071, A3 => n17624, ZN => 
                           n16070);
   U5407 : INV_X1 port map( I => n15754, ZN => n15751);
   U5412 : OAI21_X1 port map( A1 => n30024, A2 => n30022, B => n8039, ZN => 
                           n30011);
   U5414 : NAND2_X1 port map( A1 => n31371, A2 => n13151, ZN => n15602);
   U5416 : NAND2_X1 port map( A1 => n2534, A2 => n11034, ZN => n35099);
   U5418 : INV_X2 port map( I => n11034, ZN => n36099);
   U5426 : OR3_X2 port map( A1 => n24883, A2 => n19499, A3 => n18788, Z => 
                           n24681);
   U5428 : NOR2_X1 port map( A1 => n24753, A2 => n18788, ZN => n32099);
   U5429 : INV_X1 port map( I => n18788, ZN => n24680);
   U5432 : NAND2_X1 port map( A1 => n18788, A2 => n6756, ZN => n5137);
   U5435 : OAI22_X1 port map( A1 => n9066, A2 => n15903, B1 => n20839, B2 => 
                           n24296, ZN => n37634);
   U5436 : INV_X1 port map( I => n16864, ZN => n39468);
   U5438 : INV_X1 port map( I => n25303, ZN => n12441);
   U5439 : INV_X1 port map( I => n24741, ZN => n25386);
   U5440 : OR2_X2 port map( A1 => n18722, A2 => n32820, Z => n3215);
   U5441 : INV_X2 port map( I => n29284, ZN => n19090);
   U5447 : OR2_X2 port map( A1 => n11699, A2 => n10534, Z => n15968);
   U5451 : NAND2_X1 port map( A1 => n21882, A2 => n21883, ZN => n21576);
   U5455 : NAND3_X1 port map( A1 => n896, A2 => n2465, A3 => n11968, ZN => 
                           n37644);
   U5457 : AOI21_X1 port map( A1 => n30177, A2 => n20342, B => n30183, ZN => 
                           n7318);
   U5459 : CLKBUF_X2 port map( I => n16309, Z => n39025);
   U5465 : INV_X1 port map( I => n28365, ZN => n5738);
   U5466 : CLKBUF_X1 port map( I => n20597, Z => n39363);
   U5468 : INV_X1 port map( I => n28615, ZN => n32703);
   U5473 : CLKBUF_X1 port map( I => n5383, Z => n32178);
   U5478 : NAND2_X1 port map( A1 => n310, A2 => n16461, ZN => n4503);
   U5479 : CLKBUF_X8 port map( I => n39126, Z => n37671);
   U5481 : CLKBUF_X1 port map( I => n36463, Z => n39786);
   U5486 : CLKBUF_X2 port map( I => n8078, Z => n38762);
   U5488 : CLKBUF_X2 port map( I => n18860, Z => n38419);
   U5492 : INV_X2 port map( I => n31683, ZN => n38877);
   U5494 : NAND2_X1 port map( A1 => n37654, A2 => n37653, ZN => n37652);
   U5497 : NOR2_X1 port map( A1 => n2923, A2 => n11765, ZN => n37801);
   U5498 : INV_X2 port map( I => n18195, ZN => n9633);
   U5499 : NOR2_X1 port map( A1 => n27071, A2 => n36989, ZN => n37384);
   U5502 : INV_X2 port map( I => n27292, ZN => n38488);
   U5503 : NAND2_X1 port map( A1 => n26762, A2 => n26761, ZN => n37826);
   U5510 : CLKBUF_X1 port map( I => n5218, Z => n39262);
   U5512 : NAND2_X1 port map( A1 => n15196, A2 => n2081, ZN => n32799);
   U5513 : OR3_X1 port map( A1 => n38002, A2 => n1092, A3 => n37103, Z => 
                           n36112);
   U5514 : BUF_X2 port map( I => n26724, Z => n38928);
   U5521 : NOR2_X1 port map( A1 => n7725, A2 => n7516, ZN => n26798);
   U5526 : INV_X4 port map( I => n13770, ZN => n37098);
   U5529 : CLKBUF_X2 port map( I => n26185, Z => n39507);
   U5533 : AND2_X1 port map( A1 => n1518, A2 => n1017, Z => n37172);
   U5534 : AOI21_X1 port map( A1 => n11552, A2 => n18406, B => n9413, ZN => 
                           n11551);
   U5538 : BUF_X2 port map( I => n25860, Z => n36819);
   U5541 : BUF_X2 port map( I => n25971, Z => n39248);
   U5546 : CLKBUF_X1 port map( I => n9833, Z => n39165);
   U5547 : INV_X1 port map( I => n38004, ZN => n20628);
   U5550 : NAND2_X1 port map( A1 => n12748, A2 => n25517, ZN => n37339);
   U5551 : NOR2_X1 port map( A1 => n18294, A2 => n16264, ZN => n39251);
   U5552 : INV_X2 port map( I => n5042, ZN => n38728);
   U5553 : CLKBUF_X2 port map( I => n13811, Z => n38300);
   U5554 : NAND2_X1 port map( A1 => n32775, A2 => n10938, ZN => n25486);
   U5556 : CLKBUF_X2 port map( I => n25140, Z => n39295);
   U5560 : INV_X2 port map( I => n20128, ZN => n24832);
   U5568 : OAI21_X1 port map( A1 => n32785, A2 => n24478, B => n32784, ZN => 
                           n37504);
   U5576 : NOR2_X1 port map( A1 => n38349, A2 => n38561, ZN => n38652);
   U5580 : INV_X1 port map( I => n20119, ZN => n9723);
   U5590 : NAND2_X1 port map( A1 => n24397, A2 => n24396, ZN => n37710);
   U5592 : NOR2_X1 port map( A1 => n38812, A2 => n24123, ZN => n37891);
   U5594 : NAND2_X1 port map( A1 => n39415, A2 => n38251, ZN => n38250);
   U5602 : CLKBUF_X2 port map( I => n16366, Z => n39504);
   U5603 : NAND2_X1 port map( A1 => n39067, A2 => n17076, ZN => n24081);
   U5604 : INV_X2 port map( I => n30311, ZN => n39706);
   U5606 : BUF_X4 port map( I => n4880, Z => n39415);
   U5607 : CLKBUF_X2 port map( I => n20384, Z => n37896);
   U5608 : CLKBUF_X2 port map( I => n13395, Z => n39636);
   U5610 : CLKBUF_X2 port map( I => n18301, Z => n37842);
   U5616 : NAND2_X1 port map( A1 => n38894, A2 => n38893, ZN => n35753);
   U5617 : NAND2_X1 port map( A1 => n38792, A2 => n38299, ZN => n6520);
   U5620 : CLKBUF_X2 port map( I => n16013, Z => n37923);
   U5624 : OAI21_X1 port map( A1 => n10867, A2 => n2116, B => n19319, ZN => 
                           n13641);
   U5626 : CLKBUF_X2 port map( I => n17511, Z => n34823);
   U5628 : NAND2_X1 port map( A1 => n39601, A2 => n17009, ZN => n7491);
   U5630 : CLKBUF_X2 port map( I => n23162, Z => n19870);
   U5634 : NAND2_X1 port map( A1 => n23082, A2 => n14442, ZN => n38903);
   U5642 : INV_X1 port map( I => n14494, ZN => n23173);
   U5649 : OR2_X1 port map( A1 => n23189, A2 => n34200, Z => n23192);
   U5651 : AND2_X1 port map( A1 => n39075, A2 => n1149, Z => n37189);
   U5652 : AOI21_X1 port map( A1 => n20756, A2 => n33549, B => n37911, ZN => 
                           n38522);
   U5658 : BUF_X2 port map( I => n31202, Z => n37938);
   U5661 : CLKBUF_X2 port map( I => n36281, Z => n37775);
   U5667 : INV_X2 port map( I => n10463, ZN => n22143);
   U5668 : CLKBUF_X2 port map( I => n33993, Z => n38375);
   U5671 : OAI21_X1 port map( A1 => n21942, A2 => n16128, B => n19133, ZN => 
                           n37399);
   U5677 : INV_X1 port map( I => n21422, ZN => n20827);
   U5678 : INV_X1 port map( I => n19831, ZN => n37112);
   U5681 : BUF_X2 port map( I => n14245, Z => n39716);
   U5686 : INV_X1 port map( I => n19629, ZN => n37109);
   U5688 : INV_X1 port map( I => n29879, ZN => n37110);
   U5696 : NOR3_X1 port map( A1 => n30147, A2 => n30146, A3 => n3896, ZN => 
                           n39510);
   U5701 : NAND2_X1 port map( A1 => n29547, A2 => n6252, ZN => n9837);
   U5703 : NAND3_X1 port map( A1 => n29505, A2 => n29504, A3 => n16083, ZN => 
                           n38802);
   U5705 : NAND3_X1 port map( A1 => n10409, A2 => n10410, A3 => n10513, ZN => 
                           n37825);
   U5708 : OAI22_X1 port map( A1 => n29608, A2 => n29607, B1 => n37258, B2 => 
                           n37430, ZN => n29610);
   U5710 : NOR3_X1 port map( A1 => n2205, A2 => n2507, A3 => n1054, ZN => 
                           n39079);
   U5714 : INV_X1 port map( I => n30026, ZN => n30025);
   U5716 : CLKBUF_X2 port map( I => n85, Z => n34534);
   U5722 : INV_X2 port map( I => n29612, ZN => n29627);
   U5726 : CLKBUF_X4 port map( I => n17996, Z => n17997);
   U5727 : NAND2_X1 port map( A1 => n37531, A2 => n30432, ZN => n31499);
   U5728 : INV_X1 port map( I => n39006, ZN => n39005);
   U5738 : NAND2_X1 port map( A1 => n36994, A2 => n31279, ZN => n37359);
   U5753 : INV_X4 port map( I => n18815, ZN => n3700);
   U5758 : CLKBUF_X4 port map( I => n35551, Z => n36207);
   U5759 : CLKBUF_X2 port map( I => n29598, Z => n38420);
   U5763 : BUF_X2 port map( I => n10006, Z => n31583);
   U5764 : INV_X1 port map( I => n29498, ZN => n37376);
   U5765 : INV_X1 port map( I => n29694, ZN => n37752);
   U5768 : CLKBUF_X2 port map( I => n11783, Z => n39187);
   U5769 : INV_X4 port map( I => n18720, ZN => n37099);
   U5771 : INV_X2 port map( I => n29863, ZN => n29957);
   U5782 : BUF_X2 port map( I => n30221, Z => n6938);
   U5783 : BUF_X4 port map( I => n6449, Z => n6019);
   U5787 : BUF_X4 port map( I => n29312, Z => n37100);
   U5790 : INV_X1 port map( I => n18623, ZN => n39634);
   U5795 : BUF_X2 port map( I => n29054, Z => n6661);
   U5799 : INV_X1 port map( I => n39391, ZN => n37059);
   U5802 : CLKBUF_X2 port map( I => n6930, Z => n38703);
   U5808 : CLKBUF_X2 port map( I => n28610, Z => n38290);
   U5811 : CLKBUF_X2 port map( I => n12244, Z => n39536);
   U5812 : NAND2_X1 port map( A1 => n35875, A2 => n37615, ZN => n32758);
   U5814 : CLKBUF_X2 port map( I => n18453, Z => n38556);
   U5815 : NAND2_X1 port map( A1 => n28561, A2 => n38858, ZN => n38857);
   U5818 : NAND2_X1 port map( A1 => n28335, A2 => n33647, ZN => n38061);
   U5819 : NOR2_X1 port map( A1 => n6017, A2 => n28473, ZN => n39332);
   U5830 : OAI21_X1 port map( A1 => n33100, A2 => n28758, B => n13508, ZN => 
                           n32273);
   U5833 : INV_X1 port map( I => n28061, ZN => n37414);
   U5837 : NAND2_X1 port map( A1 => n28430, A2 => n9586, ZN => n37413);
   U5842 : NAND2_X1 port map( A1 => n28553, A2 => n1431, ZN => n28556);
   U5844 : INV_X1 port map( I => n28440, ZN => n37579);
   U5854 : INV_X1 port map( I => n28360, ZN => n20879);
   U5861 : INV_X1 port map( I => n34176, ZN => n28395);
   U5867 : BUF_X4 port map( I => n28621, Z => n11490);
   U5868 : CLKBUF_X2 port map( I => n15540, Z => n38566);
   U5872 : CLKBUF_X4 port map( I => n20662, Z => n11614);
   U5873 : AND2_X1 port map( A1 => n11831, A2 => n7221, Z => n35172);
   U5879 : CLKBUF_X2 port map( I => n33707, Z => n39425);
   U5881 : CLKBUF_X2 port map( I => n18480, Z => n37804);
   U5883 : CLKBUF_X2 port map( I => n38854, Z => n38075);
   U5885 : CLKBUF_X2 port map( I => n28753, Z => n37460);
   U5887 : INV_X1 port map( I => n38203, ZN => n37484);
   U5889 : NAND2_X1 port map( A1 => n37895, A2 => n11754, ZN => n38391);
   U5893 : NAND2_X1 port map( A1 => n37445, A2 => n13366, ZN => n18224);
   U5894 : NAND2_X1 port map( A1 => n8525, A2 => n8524, ZN => n39180);
   U5897 : NAND2_X1 port map( A1 => n15364, A2 => n16869, ZN => n37445);
   U5907 : OR2_X1 port map( A1 => n28205, A2 => n438, Z => n27891);
   U5908 : NAND2_X1 port map( A1 => n27940, A2 => n39193, ZN => n20019);
   U5912 : NAND2_X1 port map( A1 => n4502, A2 => n4503, ZN => n4508);
   U5914 : NOR2_X1 port map( A1 => n28101, A2 => n5266, ZN => n39193);
   U5917 : NAND2_X1 port map( A1 => n28180, A2 => n14389, ZN => n4766);
   U5918 : INV_X1 port map( I => n36643, ZN => n2467);
   U5922 : BUF_X1 port map( I => n17197, Z => n34668);
   U5924 : CLKBUF_X2 port map( I => n4945, Z => n39132);
   U5925 : AND2_X1 port map( A1 => n7528, A2 => n28282, Z => n37136);
   U5930 : CLKBUF_X2 port map( I => n18628, Z => n39789);
   U5934 : CLKBUF_X4 port map( I => n27624, Z => n28419);
   U5935 : BUF_X4 port map( I => n28182, Z => n14397);
   U5936 : BUF_X1 port map( I => n3159, Z => n38010);
   U5937 : BUF_X2 port map( I => n14411, Z => n16325);
   U5945 : BUF_X4 port map( I => n27604, Z => n28272);
   U5953 : AND2_X1 port map( A1 => n2868, A2 => n28224, Z => n37186);
   U5956 : CLKBUF_X2 port map( I => n18451, Z => n39574);
   U5957 : INV_X1 port map( I => n13883, ZN => n37540);
   U5960 : INV_X1 port map( I => n27723, ZN => n37427);
   U5970 : BUF_X2 port map( I => n13703, Z => n386);
   U5971 : CLKBUF_X2 port map( I => n27647, Z => n18577);
   U5977 : BUF_X2 port map( I => n4127, Z => n35350);
   U5979 : CLKBUF_X4 port map( I => n12551, Z => n37101);
   U5982 : NAND2_X1 port map( A1 => n35681, A2 => n39572, ZN => n32245);
   U5985 : NAND2_X1 port map( A1 => n20203, A2 => n27312, ZN => n38635);
   U5986 : INV_X1 port map( I => n38152, ZN => n38515);
   U5989 : INV_X1 port map( I => n37433, ZN => n37432);
   U6002 : NAND2_X1 port map( A1 => n6508, A2 => n6507, ZN => n38587);
   U6013 : NAND2_X1 port map( A1 => n26647, A2 => n38690, ZN => n38688);
   U6015 : NAND2_X1 port map( A1 => n35978, A2 => n38637, ZN => n38636);
   U6024 : INV_X1 port map( I => n27354, ZN => n39485);
   U6029 : INV_X1 port map( I => n39573, ZN => n39572);
   U6033 : NAND2_X1 port map( A1 => n27289, A2 => n37130, ZN => n18769);
   U6041 : INV_X1 port map( I => n15641, ZN => n38489);
   U6063 : NOR2_X1 port map( A1 => n37771, A2 => n37770, ZN => n8535);
   U6064 : OR2_X1 port map( A1 => n5101, A2 => n27240, Z => n37158);
   U6067 : NOR2_X1 port map( A1 => n37385, A2 => n37384, ZN => n35294);
   U6069 : OAI21_X1 port map( A1 => n27096, A2 => n13992, B => n27441, ZN => 
                           n37903);
   U6072 : NAND2_X1 port map( A1 => n38306, A2 => n38305, ZN => n31926);
   U6074 : NOR2_X1 port map( A1 => n4627, A2 => n6191, ZN => n37655);
   U6075 : OAI21_X1 port map( A1 => n19326, A2 => n27131, B => n27338, ZN => 
                           n39336);
   U6079 : OR2_X1 port map( A1 => n18195, A2 => n38193, Z => n9632);
   U6081 : NOR2_X1 port map( A1 => n38983, A2 => n27253, ZN => n27255);
   U6089 : INV_X2 port map( I => n27435, ZN => n27149);
   U6092 : INV_X1 port map( I => n12766, ZN => n37827);
   U6096 : INV_X2 port map( I => n27379, ZN => n27298);
   U6097 : CLKBUF_X2 port map( I => n39484, Z => n38571);
   U6100 : CLKBUF_X2 port map( I => n9144, Z => n33503);
   U6104 : INV_X2 port map( I => n15284, ZN => n27278);
   U6110 : AND2_X1 port map( A1 => n6908, A2 => n21272, Z => n37192);
   U6119 : CLKBUF_X4 port map( I => n36200, Z => n34387);
   U6125 : CLKBUF_X2 port map( I => n35500, Z => n39216);
   U6132 : CLKBUF_X4 port map( I => n27438, Z => n7612);
   U6139 : INV_X1 port map( I => n16835, ZN => n38983);
   U6142 : CLKBUF_X4 port map( I => n6533, Z => n39414);
   U6144 : CLKBUF_X2 port map( I => n4886, Z => n39628);
   U6145 : CLKBUF_X2 port map( I => n16736, Z => n38578);
   U6147 : NAND2_X1 port map( A1 => n38363, A2 => n38362, ZN => n26446);
   U6159 : NOR2_X1 port map( A1 => n12795, A2 => n37161, ZN => n33098);
   U6167 : AND3_X1 port map( A1 => n33849, A2 => n19179, A3 => n37098, Z => 
                           n37161);
   U6168 : AOI21_X1 port map( A1 => n26618, A2 => n34003, B => n26621, ZN => 
                           n9658);
   U6170 : NAND2_X1 port map( A1 => n26785, A2 => n26862, ZN => n4);
   U6172 : NAND2_X1 port map( A1 => n1491, A2 => n8746, ZN => n38362);
   U6174 : AND2_X1 port map( A1 => n26847, A2 => n26945, Z => n37133);
   U6175 : NAND2_X1 port map( A1 => n26443, A2 => n33689, ZN => n38363);
   U6176 : AND2_X1 port map( A1 => n32344, A2 => n7619, Z => n37131);
   U6177 : OR2_X1 port map( A1 => n10187, A2 => n8478, Z => n37188);
   U6178 : INV_X1 port map( I => n32072, ZN => n37590);
   U6181 : INV_X4 port map( I => n10338, ZN => n37102);
   U6184 : INV_X1 port map( I => n27013, ZN => n39064);
   U6187 : NAND2_X1 port map( A1 => n26769, A2 => n19442, ZN => n16939);
   U6188 : NOR2_X1 port map( A1 => n20666, A2 => n26990, ZN => n19191);
   U6189 : OR2_X1 port map( A1 => n16160, A2 => n20858, Z => n34003);
   U6190 : CLKBUF_X2 port map( I => n26837, Z => n38407);
   U6195 : OR2_X1 port map( A1 => n26876, A2 => n21099, Z => n37140);
   U6197 : CLKBUF_X2 port map( I => n34160, Z => n38483);
   U6199 : BUF_X4 port map( I => n11617, Z => n11616);
   U6200 : OR2_X1 port map( A1 => n20171, A2 => n26770, Z => n4808);
   U6204 : CLKBUF_X2 port map( I => n11948, Z => n39564);
   U6205 : BUF_X4 port map( I => n26836, Z => n37103);
   U6208 : CLKBUF_X4 port map( I => n26808, Z => n19179);
   U6209 : INV_X1 port map( I => n31546, ZN => n39602);
   U6210 : CLKBUF_X4 port map( I => n12788, Z => n37104);
   U6212 : INV_X1 port map( I => n39611, ZN => n26475);
   U6216 : CLKBUF_X2 port map( I => n26361, Z => n38896);
   U6219 : BUF_X2 port map( I => n4875, Z => n39637);
   U6220 : CLKBUF_X2 port map( I => n30913, Z => n39093);
   U6221 : NAND2_X1 port map( A1 => n37930, A2 => n35947, ZN => n30967);
   U6222 : NOR2_X1 port map( A1 => n37372, A2 => n18801, ZN => n6478);
   U6223 : NAND2_X1 port map( A1 => n14985, A2 => n38783, ZN => n14984);
   U6225 : NAND2_X2 port map( A1 => n9868, A2 => n25920, ZN => n25596);
   U6228 : INV_X1 port map( I => n38930, ZN => n34512);
   U6229 : AND2_X1 port map( A1 => n7258, A2 => n11033, Z => n37116);
   U6230 : INV_X1 port map( I => n30957, ZN => n37310);
   U6232 : BUF_X1 port map( I => n1015, Z => n37837);
   U6233 : INV_X2 port map( I => n5753, ZN => n34577);
   U6237 : CLKBUF_X1 port map( I => n9412, Z => n37819);
   U6241 : CLKBUF_X2 port map( I => n9694, Z => n39375);
   U6242 : CLKBUF_X2 port map( I => n33879, Z => n37502);
   U6246 : INV_X1 port map( I => n31367, ZN => n37746);
   U6250 : BUF_X1 port map( I => n26108, Z => n38501);
   U6253 : CLKBUF_X2 port map( I => n17696, Z => n38507);
   U6254 : CLKBUF_X2 port map( I => n17180, Z => n38760);
   U6255 : CLKBUF_X4 port map( I => n25899, Z => n38825);
   U6256 : NAND2_X1 port map( A1 => n1932, A2 => n1933, ZN => n21204);
   U6257 : CLKBUF_X2 port map( I => n26093, Z => n39729);
   U6259 : NAND2_X1 port map( A1 => n37713, A2 => n37712, ZN => n37711);
   U6262 : OAI21_X1 port map( A1 => n19829, A2 => n10444, B => n38013, ZN => 
                           n38132);
   U6268 : NAND2_X1 port map( A1 => n25645, A2 => n4467, ZN => n37616);
   U6270 : OAI21_X1 port map( A1 => n39252, A2 => n39251, B => n5051, ZN => 
                           n25635);
   U6271 : NAND2_X1 port map( A1 => n9429, A2 => n15329, ZN => n38301);
   U6272 : OR2_X1 port map( A1 => n219, A2 => n32879, Z => n38933);
   U6273 : INV_X1 port map( I => n38050, ZN => n6173);
   U6275 : OR2_X1 port map( A1 => n39328, A2 => n17029, Z => n37182);
   U6277 : AND2_X1 port map( A1 => n14436, A2 => n12533, Z => n6472);
   U6291 : CLKBUF_X2 port map( I => n31895, Z => n37748);
   U6296 : BUF_X2 port map( I => n32775, Z => n38245);
   U6299 : NAND2_X1 port map( A1 => n38863, A2 => n38862, ZN => n38113);
   U6304 : CLKBUF_X4 port map( I => n10414, Z => n39599);
   U6311 : CLKBUF_X2 port map( I => n11622, Z => n38178);
   U6328 : CLKBUF_X2 port map( I => n19582, Z => n39389);
   U6332 : CLKBUF_X4 port map( I => n25700, Z => n12675);
   U6334 : BUF_X2 port map( I => n32165, Z => n15172);
   U6335 : CLKBUF_X2 port map( I => n13873, Z => n38661);
   U6341 : CLKBUF_X2 port map( I => n32433, Z => n38560);
   U6343 : CLKBUF_X2 port map( I => n25186, Z => n39146);
   U6344 : CLKBUF_X2 port map( I => n33132, Z => n37312);
   U6346 : CLKBUF_X4 port map( I => n25269, Z => n39765);
   U6350 : CLKBUF_X2 port map( I => n25118, Z => n38665);
   U6360 : CLKBUF_X2 port map( I => n24999, Z => n38950);
   U6362 : NAND2_X1 port map( A1 => n17106, A2 => n9612, ZN => n39496);
   U6365 : NAND2_X1 port map( A1 => n11367, A2 => n38389, ZN => n4427);
   U6366 : INV_X1 port map( I => n39256, ZN => n39255);
   U6377 : NAND2_X1 port map( A1 => n10793, A2 => n37193, ZN => n24884);
   U6385 : BUF_X2 port map( I => n8605, Z => n507);
   U6387 : NAND2_X1 port map( A1 => n30700, A2 => n30698, ZN => n37664);
   U6388 : NOR2_X1 port map( A1 => n37233, A2 => n6357, ZN => n30386);
   U6397 : OR2_X1 port map( A1 => n24898, A2 => n38317, Z => n31455);
   U6405 : INV_X1 port map( I => n24776, ZN => n39540);
   U6409 : CLKBUF_X2 port map( I => n1118, Z => n38631);
   U6420 : NOR2_X1 port map( A1 => n1263, A2 => n16671, ZN => n37688);
   U6426 : NAND2_X1 port map( A1 => n38347, A2 => n24696, ZN => n23857);
   U6467 : CLKBUF_X8 port map( I => n33996, Z => n37477);
   U6475 : BUF_X4 port map( I => n39681, Z => n31845);
   U6476 : CLKBUF_X2 port map( I => n7769, Z => n37640);
   U6477 : BUF_X1 port map( I => n7770, Z => n39513);
   U6481 : BUF_X4 port map( I => n17607, Z => n37355);
   U6482 : CLKBUF_X8 port map( I => n32825, Z => n37105);
   U6485 : BUF_X2 port map( I => n24779, Z => n38658);
   U6489 : NAND2_X1 port map( A1 => n37891, A2 => n18647, ZN => n18608);
   U6491 : CLKBUF_X1 port map( I => n24753, Z => n38884);
   U6492 : INV_X2 port map( I => n24650, ZN => n36988);
   U6493 : NAND2_X1 port map( A1 => n38652, A2 => n38250, ZN => n37472);
   U6497 : NAND2_X1 port map( A1 => n39660, A2 => n39659, ZN => n18647);
   U6500 : NAND2_X1 port map( A1 => n34938, A2 => n24069, ZN => n39092);
   U6515 : NAND2_X1 port map( A1 => n37710, A2 => n24170, ZN => n38925);
   U6516 : NAND2_X1 port map( A1 => n24305, A2 => n39796, ZN => n8319);
   U6517 : NAND2_X1 port map( A1 => n24253, A2 => n19782, ZN => n39587);
   U6518 : NAND2_X1 port map( A1 => n37959, A2 => n37958, ZN => n5716);
   U6520 : NAND2_X1 port map( A1 => n18759, A2 => n7000, ZN => n6999);
   U6524 : INV_X1 port map( I => n16377, ZN => n38473);
   U6525 : NOR2_X1 port map( A1 => n6933, A2 => n24453, ZN => n37392);
   U6546 : NAND2_X1 port map( A1 => n4359, A2 => n24336, ZN => n37635);
   U6558 : NAND2_X1 port map( A1 => n9083, A2 => n9084, ZN => n39738);
   U6561 : AND2_X1 port map( A1 => n24396, A2 => n24169, Z => n37187);
   U6567 : NAND2_X1 port map( A1 => n38948, A2 => n11477, ZN => n12176);
   U6570 : NAND2_X1 port map( A1 => n16666, A2 => n24372, ZN => n37959);
   U6571 : CLKBUF_X2 port map( I => n24381, Z => n38812);
   U6582 : CLKBUF_X4 port map( I => n1129, Z => n38431);
   U6583 : INV_X1 port map( I => n24470, ZN => n38032);
   U6585 : INV_X2 port map( I => n13099, ZN => n24169);
   U6590 : CLKBUF_X2 port map( I => n18830, Z => n38487);
   U6593 : CLKBUF_X2 port map( I => n17871, Z => n37733);
   U6594 : INV_X1 port map( I => n32899, ZN => n38251);
   U6595 : BUF_X1 port map( I => n12235, Z => n37994);
   U6596 : BUF_X4 port map( I => n37267, Z => n39067);
   U6618 : CLKBUF_X2 port map( I => n11795, Z => n37480);
   U6619 : BUF_X2 port map( I => n24106, Z => n24396);
   U6620 : INV_X1 port map( I => n23565, ZN => n37352);
   U6622 : BUF_X4 port map( I => n2297, Z => n37107);
   U6625 : INV_X1 port map( I => n20384, ZN => n35134);
   U6634 : INV_X1 port map( I => n7558, ZN => n17288);
   U6637 : INV_X1 port map( I => n16833, ZN => n5667);
   U6645 : CLKBUF_X2 port map( I => n39163, Z => n37899);
   U6646 : CLKBUF_X2 port map( I => n3601, Z => n39014);
   U6651 : NAND2_X1 port map( A1 => n2960, A2 => n7389, ZN => n39506);
   U6653 : INV_X1 port map( I => n12362, ZN => n32562);
   U6657 : CLKBUF_X2 port map( I => n39038, Z => n38370);
   U6668 : NAND2_X1 port map( A1 => n32407, A2 => n32406, ZN => n37705);
   U6678 : NAND2_X1 port map( A1 => n30788, A2 => n37924, ZN => n39218);
   U6680 : CLKBUF_X2 port map( I => n23619, Z => n37431);
   U6682 : NAND2_X1 port map( A1 => n4534, A2 => n37266, ZN => n36966);
   U6687 : INV_X2 port map( I => n36859, ZN => n38894);
   U6689 : NAND2_X1 port map( A1 => n30524, A2 => n38726, ZN => n23385);
   U6704 : BUF_X2 port map( I => n18204, Z => n7387);
   U6710 : AND3_X1 port map( A1 => n23477, A2 => n1139, A3 => n15176, Z => 
                           n37135);
   U6712 : CLKBUF_X2 port map( I => n23355, Z => n39534);
   U6714 : CLKBUF_X4 port map( I => n13217, Z => n37523);
   U6715 : INV_X2 port map( I => n18199, ZN => n23355);
   U6719 : BUF_X1 port map( I => n23310, Z => n39626);
   U6721 : BUF_X1 port map( I => n23548, Z => n38656);
   U6725 : CLKBUF_X2 port map( I => n1635, Z => n37622);
   U6729 : INV_X2 port map( I => n32471, ZN => n1304);
   U6730 : CLKBUF_X2 port map( I => n23423, Z => n37814);
   U6731 : CLKBUF_X2 port map( I => n19671, Z => n37463);
   U6735 : INV_X2 port map( I => n11342, ZN => n31234);
   U6736 : CLKBUF_X2 port map( I => n30881, Z => n38042);
   U6738 : NOR2_X1 port map( A1 => n783, A2 => n37127, ZN => n37500);
   U6741 : AOI22_X1 port map( A1 => n17498, A2 => n23165, B1 => n17497, B2 => 
                           n23169, ZN => n37901);
   U6744 : NOR2_X1 port map( A1 => n37840, A2 => n14851, ZN => n20910);
   U6752 : CLKBUF_X2 port map( I => n38653, Z => n38100);
   U6755 : OAI21_X1 port map( A1 => n23061, A2 => n23000, B => n36167, ZN => 
                           n38967);
   U6762 : NAND2_X1 port map( A1 => n39297, A2 => n15032, ZN => n35067);
   U6765 : OAI21_X1 port map( A1 => n23082, A2 => n5515, B => n38903, ZN => 
                           n22910);
   U6767 : NOR2_X1 port map( A1 => n7626, A2 => n12630, ZN => n37518);
   U6774 : CLKBUF_X2 port map( I => n23173, Z => n38752);
   U6775 : NAND3_X1 port map( A1 => n23209, A2 => n23135, A3 => n19859, ZN => 
                           n23134);
   U6783 : BUF_X2 port map( I => n19731, Z => n121);
   U6784 : CLKBUF_X2 port map( I => n780, Z => n38329);
   U6788 : BUF_X2 port map( I => n22864, Z => n19288);
   U6792 : CLKBUF_X2 port map( I => n7584, Z => n38542);
   U6795 : BUF_X2 port map( I => n34200, Z => n5515);
   U6803 : CLKBUF_X2 port map( I => n1319, Z => n39034);
   U6806 : CLKBUF_X2 port map( I => n23074, Z => n31005);
   U6807 : CLKBUF_X4 port map( I => n7518, Z => n6466);
   U6818 : BUF_X2 port map( I => n22879, Z => n4682);
   U6819 : INV_X4 port map( I => n1046, ZN => n37108);
   U6821 : BUF_X4 port map( I => n22942, Z => n19586);
   U6825 : CLKBUF_X1 port map( I => n10382, Z => n38216);
   U6828 : CLKBUF_X4 port map( I => n4624, Z => n39787);
   U6835 : CLKBUF_X2 port map( I => n16798, Z => n39548);
   U6842 : CLKBUF_X2 port map( I => n9982, Z => n38330);
   U6844 : NAND2_X1 port map( A1 => n22141, A2 => n20731, ZN => n37708);
   U6845 : INV_X1 port map( I => n38522, ZN => n10996);
   U6849 : NAND2_X1 port map( A1 => n22319, A2 => n38917, ZN => n12815);
   U6853 : OAI21_X1 port map( A1 => n21963, A2 => n9987, B => n38699, ZN => 
                           n20042);
   U6854 : INV_X1 port map( I => n21972, ZN => n17636);
   U6862 : INV_X1 port map( I => n37491, ZN => n37490);
   U6863 : INV_X1 port map( I => n22282, ZN => n38105);
   U6864 : CLKBUF_X2 port map( I => n11329, Z => n37911);
   U6866 : AND3_X1 port map( A1 => n32107, A2 => n22349, A3 => n22389, Z => 
                           n2886);
   U6870 : CLKBUF_X2 port map( I => n22254, Z => n39151);
   U6871 : NAND2_X1 port map( A1 => n22205, A2 => n21288, ZN => n38931);
   U6877 : BUF_X2 port map( I => n22362, Z => n34246);
   U6882 : BUF_X2 port map( I => n22170, Z => n554);
   U6889 : BUF_X2 port map( I => n6947, Z => n6361);
   U6891 : CLKBUF_X2 port map( I => n38395, Z => n38246);
   U6892 : NAND2_X1 port map( A1 => n13239, A2 => n13240, ZN => n39746);
   U6897 : INV_X1 port map( I => n37789, ZN => n17436);
   U6900 : NAND2_X1 port map( A1 => n13345, A2 => n17161, ZN => n34683);
   U6902 : AOI22_X1 port map( A1 => n21343, A2 => n21861, B1 => n21342, B2 => 
                           n36351, ZN => n39771);
   U6907 : NAND2_X1 port map( A1 => n21649, A2 => n1157, ZN => n38547);
   U6910 : NAND2_X1 port map( A1 => n20367, A2 => n21950, ZN => n39658);
   U6915 : INV_X1 port map( I => n37399, ZN => n37398);
   U6917 : NAND2_X1 port map( A1 => n21695, A2 => n21876, ZN => n39732);
   U6918 : BUF_X2 port map( I => n21905, Z => n19647);
   U6920 : CLKBUF_X2 port map( I => n21593, Z => n38480);
   U6926 : BUF_X2 port map( I => n12754, Z => n35839);
   U6927 : NAND2_X1 port map( A1 => n19650, A2 => n21876, ZN => n21873);
   U6929 : CLKBUF_X4 port map( I => n21883, Z => n19434);
   U6935 : INV_X1 port map( I => n30170, ZN => n38261);
   U6936 : CLKBUF_X2 port map( I => n21628, Z => n32412);
   U6942 : CLKBUF_X2 port map( I => n10656, Z => n39656);
   U6944 : CLKBUF_X2 port map( I => n21641, Z => n39650);
   U6948 : INV_X1 port map( I => n19919, ZN => n38962);
   U6949 : INV_X1 port map( I => n29805, ZN => n37261);
   U6962 : BUF_X2 port map( I => n15009, Z => n37111);
   U6965 : INV_X1 port map( I => Plaintext(151), ZN => n38991);
   U6966 : INV_X1 port map( I => n4759, ZN => n37659);
   U6971 : INV_X1 port map( I => n9759, ZN => n38273);
   U6972 : NOR2_X1 port map( A1 => n20003, A2 => n18028, ZN => n16537);
   U6974 : INV_X1 port map( I => n21929, ZN => n36721);
   U6975 : NAND2_X1 port map( A1 => n21787, A2 => n18205, ZN => n17966);
   U6979 : CLKBUF_X1 port map( I => n21669, Z => n31222);
   U6983 : INV_X1 port map( I => n21582, ZN => n19579);
   U6985 : NAND2_X1 port map( A1 => n21274, A2 => n7536, ZN => n38496);
   U6988 : CLKBUF_X1 port map( I => n32820, Z => n39594);
   U6991 : CLKBUF_X2 port map( I => n33999, Z => n39192);
   U6993 : NOR2_X1 port map( A1 => n19403, A2 => n19554, ZN => n19553);
   U7000 : NAND2_X1 port map( A1 => n19084, A2 => n12754, ZN => n2643);
   U7004 : AOI21_X1 port map( A1 => n21820, A2 => n39594, B => n1349, ZN => 
                           n14734);
   U7007 : CLKBUF_X1 port map( I => n21721, Z => n32704);
   U7009 : CLKBUF_X4 port map( I => n3839, Z => n3562);
   U7010 : CLKBUF_X1 port map( I => n21644, Z => n18112);
   U7013 : NOR2_X1 port map( A1 => n21804, A2 => n36735, ZN => n10127);
   U7019 : NAND2_X1 port map( A1 => n21555, A2 => n10211, ZN => n10144);
   U7021 : NAND2_X1 port map( A1 => n21713, A2 => n19542, ZN => n21531);
   U7030 : INV_X1 port map( I => n21854, ZN => n21852);
   U7036 : NAND3_X1 port map( A1 => n1156, A2 => n38241, A3 => n1345, ZN => 
                           n7963);
   U7040 : NAND2_X1 port map( A1 => n14928, A2 => n22315, ZN => n19136);
   U7044 : INV_X1 port map( I => n37963, ZN => n37962);
   U7047 : CLKBUF_X2 port map( I => n36728, Z => n21783);
   U7054 : NAND2_X1 port map( A1 => n30824, A2 => n3564, ZN => n39785);
   U7059 : NAND2_X1 port map( A1 => n6101, A2 => n21850, ZN => n6098);
   U7061 : NAND2_X1 port map( A1 => n5391, A2 => n5392, ZN => n13438);
   U7066 : INV_X2 port map( I => n22229, ZN => n1675);
   U7067 : INV_X1 port map( I => n22316, ZN => n915);
   U7073 : CLKBUF_X4 port map( I => n21488, Z => n21893);
   U7074 : BUF_X2 port map( I => n22292, Z => n33571);
   U7079 : OAI21_X1 port map( A1 => n22176, A2 => n4613, B => n22335, ZN => 
                           n21298);
   U7083 : OAI21_X1 port map( A1 => n11091, A2 => n39075, B => n1680, ZN => 
                           n11142);
   U7084 : NAND2_X1 port map( A1 => n22365, A2 => n7357, ZN => n22007);
   U7087 : CLKBUF_X2 port map( I => n15350, Z => n36227);
   U7093 : NOR2_X1 port map( A1 => n37358, A2 => n33886, ZN => n19777);
   U7104 : CLKBUF_X4 port map( I => n5929, Z => n5075);
   U7108 : AOI21_X1 port map( A1 => n133, A2 => n17897, B => n7613, ZN => 
                           n20254);
   U7112 : INV_X2 port map( I => n4613, ZN => n22101);
   U7117 : NOR2_X1 port map( A1 => n6347, A2 => n2257, ZN => n2816);
   U7128 : AOI21_X1 port map( A1 => n915, A2 => n22317, B => n9824, ZN => 
                           n12433);
   U7131 : NAND2_X1 port map( A1 => n11171, A2 => n36397, ZN => n19385);
   U7134 : NAND2_X1 port map( A1 => n39151, A2 => n17723, ZN => n12091);
   U7137 : OAI22_X1 port map( A1 => n18429, A2 => n20623, B1 => n22365, B2 => 
                           n22366, ZN => n11878);
   U7138 : NAND2_X1 port map( A1 => n12365, A2 => n22324, ZN => n37918);
   U7141 : NAND3_X1 port map( A1 => n22061, A2 => n22178, A3 => n19261, ZN => 
                           n16259);
   U7143 : INV_X1 port map( I => n22511, ZN => n22695);
   U7146 : CLKBUF_X1 port map( I => n22621, Z => n39654);
   U7152 : INV_X1 port map( I => n15871, ZN => n22677);
   U7153 : INV_X1 port map( I => n15439, ZN => n38920);
   U7157 : OAI21_X1 port map( A1 => n16346, A2 => n16345, B => n15439, ZN => 
                           n6048);
   U7161 : NAND2_X1 port map( A1 => n22255, A2 => n20308, ZN => n17407);
   U7162 : INV_X1 port map( I => n7510, ZN => n10384);
   U7172 : INV_X1 port map( I => n22689, ZN => n3233);
   U7180 : INV_X1 port map( I => n22435, ZN => n39047);
   U7185 : NAND2_X1 port map( A1 => n33925, A2 => n14409, ZN => n19724);
   U7186 : NAND2_X1 port map( A1 => n10383, A2 => n15794, ZN => n13719);
   U7187 : NAND3_X1 port map( A1 => n20439, A2 => n17127, A3 => n1989, ZN => 
                           n3289);
   U7188 : NAND2_X1 port map( A1 => n14524, A2 => n5907, ZN => n22799);
   U7196 : NAND2_X1 port map( A1 => n20957, A2 => n23079, ZN => n32358);
   U7199 : OAI22_X1 port map( A1 => n15678, A2 => n781, B1 => n22895, B2 => 
                           n35918, ZN => n14544);
   U7201 : NAND2_X1 port map( A1 => n33935, A2 => n8197, ZN => n7804);
   U7205 : NOR2_X1 port map( A1 => n15455, A2 => n14089, ZN => n22948);
   U7208 : INV_X2 port map( I => n19966, ZN => n1648);
   U7209 : NOR2_X1 port map( A1 => n8628, A2 => n16174, ZN => n34522);
   U7215 : CLKBUF_X2 port map( I => n23080, Z => n4846);
   U7220 : INV_X1 port map( I => n38282, ZN => n22889);
   U7226 : CLKBUF_X2 port map( I => n23132, Z => n17578);
   U7230 : INV_X1 port map( I => n33972, ZN => n22931);
   U7238 : AOI21_X1 port map( A1 => n17131, A2 => n17127, B => n39810, ZN => 
                           n18481);
   U7244 : CLKBUF_X1 port map( I => n23188, Z => n39266);
   U7245 : INV_X2 port map( I => n22802, ZN => n1645);
   U7246 : NAND2_X1 port map( A1 => n22949, A2 => n37108, ZN => n22722);
   U7248 : AOI21_X1 port map( A1 => n23166, A2 => n22975, B => n36554, ZN => 
                           n22976);
   U7250 : NOR2_X1 port map( A1 => n38019, A2 => n4773, ZN => n37913);
   U7252 : INV_X2 port map( I => n14409, ZN => n13946);
   U7253 : OAI21_X1 port map( A1 => n22802, A2 => n32228, B => n19134, ZN => 
                           n9798);
   U7254 : NAND2_X1 port map( A1 => n8676, A2 => n14804, ZN => n33585);
   U7263 : NAND2_X1 port map( A1 => n9797, A2 => n20518, ZN => n14744);
   U7271 : AOI22_X1 port map( A1 => n23044, A2 => n22368, B1 => n1989, B2 => 
                           n5806, ZN => n5805);
   U7274 : AOI21_X1 port map( A1 => n10378, A2 => n10377, B => n8730, ZN => 
                           n37840);
   U7275 : NAND2_X1 port map( A1 => n22993, A2 => n22994, ZN => n23067);
   U7283 : CLKBUF_X2 port map( I => n20077, Z => n39418);
   U7286 : INV_X1 port map( I => n14561, ZN => n23212);
   U7290 : INV_X1 port map( I => n37043, ZN => n9543);
   U7305 : INV_X1 port map( I => n18481, ZN => n37792);
   U7306 : OAI22_X1 port map( A1 => n5658, A2 => n5657, B1 => n23197, B2 => 
                           n12245, ZN => n327);
   U7323 : NAND2_X1 port map( A1 => n1304, A2 => n20418, ZN => n30789);
   U7325 : INV_X1 port map( I => n9823, ZN => n18284);
   U7327 : INV_X1 port map( I => n23456, ZN => n23293);
   U7333 : NAND3_X1 port map( A1 => n1043, A2 => n1146, A3 => n31838, ZN => 
                           n13078);
   U7336 : AOI21_X1 port map( A1 => n936, A2 => n23020, B => n1046, ZN => 
                           n35939);
   U7345 : CLKBUF_X4 port map( I => n22005, Z => n23111);
   U7346 : OAI21_X1 port map( A1 => n38248, A2 => n1136, B => n9321, ZN => 
                           n38376);
   U7350 : NAND3_X1 port map( A1 => n1632, A2 => n21247, A3 => n23602, ZN => 
                           n23604);
   U7352 : INV_X2 port map( I => n10334, ZN => n1144);
   U7353 : AOI21_X1 port map( A1 => n23401, A2 => n16047, B => n38353, ZN => 
                           n12639);
   U7355 : OAI21_X1 port map( A1 => n23358, A2 => n23250, B => n33864, ZN => 
                           n31055);
   U7358 : INV_X1 port map( I => n19005, ZN => n21051);
   U7359 : INV_X1 port map( I => n37354, ZN => n36635);
   U7362 : INV_X1 port map( I => n35001, ZN => n38299);
   U7366 : NAND2_X1 port map( A1 => n16047, A2 => n23400, ZN => n37924);
   U7372 : AOI21_X1 port map( A1 => n18939, A2 => n36564, B => n30456, ZN => 
                           n38373);
   U7374 : INV_X1 port map( I => n15353, ZN => n5759);
   U7375 : NAND3_X1 port map( A1 => n23370, A2 => n9823, A3 => n1140, ZN => 
                           n4287);
   U7380 : NAND2_X1 port map( A1 => n23493, A2 => n23315, ZN => n22966);
   U7381 : NOR2_X1 port map( A1 => n38535, A2 => n37463, ZN => n20818);
   U7382 : NOR3_X1 port map( A1 => n1290, A2 => n39194, A3 => n13414, ZN => 
                           n9772);
   U7389 : OAI21_X1 port map( A1 => n1304, A2 => n30499, B => n12638, ZN => 
                           n18917);
   U7396 : NAND2_X1 port map( A1 => n19869, A2 => n18850, ZN => n23009);
   U7401 : NAND2_X1 port map( A1 => n20418, A2 => n36810, ZN => n20776);
   U7408 : CLKBUF_X2 port map( I => n12966, Z => n38881);
   U7409 : NAND2_X1 port map( A1 => n4525, A2 => n38611, ZN => n35302);
   U7410 : INV_X2 port map( I => n23749, ZN => n10763);
   U7419 : INV_X1 port map( I => n23515, ZN => n1293);
   U7423 : CLKBUF_X4 port map( I => n18681, Z => n32858);
   U7424 : NOR2_X1 port map( A1 => n16013, A2 => n23619, ZN => n23455);
   U7431 : AOI21_X1 port map( A1 => n37523, A2 => n23350, B => n31906, ZN => 
                           n38754);
   U7432 : AOI21_X1 port map( A1 => n23321, A2 => n16299, B => n23320, ZN => 
                           n23322);
   U7435 : CLKBUF_X2 port map( I => n23967, Z => n35561);
   U7441 : INV_X1 port map( I => n6559, ZN => n36143);
   U7447 : NAND2_X1 port map( A1 => n12597, A2 => n23303, ZN => n32406);
   U7449 : INV_X1 port map( I => n4117, ZN => n7833);
   U7452 : CLKBUF_X4 port map( I => n12362, Z => n5116);
   U7453 : INV_X1 port map( I => n23943, ZN => n30688);
   U7454 : INV_X1 port map( I => n23729, ZN => n36068);
   U7459 : NOR2_X1 port map( A1 => n9193, A2 => n39648, ZN => n10589);
   U7468 : INV_X1 port map( I => n12799, ZN => n11794);
   U7469 : NOR2_X1 port map( A1 => n19656, A2 => n23976, ZN => n2223);
   U7471 : CLKBUF_X2 port map( I => n24052, Z => n39310);
   U7475 : NOR2_X1 port map( A1 => n24235, A2 => n10477, ZN => n32787);
   U7478 : NAND2_X1 port map( A1 => n23819, A2 => n34561, ZN => n36003);
   U7480 : NAND2_X1 port map( A1 => n20404, A2 => n37230, ZN => n34330);
   U7481 : NAND2_X1 port map( A1 => n19857, A2 => n24271, ZN => n38595);
   U7485 : INV_X1 port map( I => n1131, ZN => n6465);
   U7486 : NAND2_X1 port map( A1 => n4880, A2 => n21043, ZN => n4286);
   U7488 : NAND2_X1 port map( A1 => n39706, A2 => n94, ZN => n7772);
   U7493 : NOR2_X1 port map( A1 => n32899, A2 => n4880, ZN => n37580);
   U7497 : INV_X1 port map( I => n39605, ZN => n37849);
   U7499 : NAND2_X1 port map( A1 => n24271, A2 => n11795, ZN => n24272);
   U7503 : NAND2_X1 port map( A1 => n38473, A2 => n1130, ZN => n38472);
   U7507 : NAND2_X1 port map( A1 => n2348, A2 => n11585, ZN => n36561);
   U7509 : NOR2_X1 port map( A1 => n24458, A2 => n38886, ZN => n35854);
   U7510 : NOR2_X1 port map( A1 => n24390, A2 => n9963, ZN => n24187);
   U7513 : INV_X1 port map( I => n24164, ZN => n24484);
   U7514 : AOI21_X1 port map( A1 => n1128, A2 => n1130, B => n38032, ZN => 
                           n8360);
   U7515 : NOR2_X1 port map( A1 => n24329, A2 => n24328, ZN => n31443);
   U7518 : INV_X1 port map( I => n24467, ZN => n1600);
   U7527 : NOR2_X1 port map( A1 => n39067, A2 => n24461, ZN => n20395);
   U7529 : NAND2_X1 port map( A1 => n2395, A2 => n2393, ZN => n2400);
   U7530 : NOR2_X1 port map( A1 => n1275, A2 => n39699, ZN => n34133);
   U7532 : OAI22_X1 port map( A1 => n1601, A2 => n24309, B1 => n19745, B2 => 
                           n24445, ZN => n24137);
   U7535 : OAI21_X1 port map( A1 => n16590, A2 => n1594, B => n24412, ZN => 
                           n12425);
   U7542 : INV_X1 port map( I => n18830, ZN => n24382);
   U7545 : INV_X1 port map( I => n12804, ZN => n24399);
   U7550 : NAND2_X1 port map( A1 => n24650, A2 => n37477, ZN => n15850);
   U7552 : INV_X2 port map( I => n17693, ZN => n1586);
   U7554 : NOR2_X1 port map( A1 => n35952, A2 => n32093, ZN => n34372);
   U7555 : NAND2_X1 port map( A1 => n18721, A2 => n33104, ZN => n17811);
   U7557 : OAI21_X1 port map( A1 => n14617, A2 => n18551, B => n24464, ZN => 
                           n18550);
   U7558 : NAND2_X1 port map( A1 => n10815, A2 => n37994, ZN => n5138);
   U7560 : NAND2_X1 port map( A1 => n19566, A2 => n205, ZN => n24157);
   U7565 : NOR2_X1 port map( A1 => n12665, A2 => n36154, ZN => n34656);
   U7566 : NAND3_X1 port map( A1 => n24442, A2 => n24443, A3 => n250, ZN => 
                           n5066);
   U7567 : NOR2_X1 port map( A1 => n3226, A2 => n24400, ZN => n32484);
   U7573 : NAND2_X1 port map( A1 => n4050, A2 => n2989, ZN => n13228);
   U7574 : AOI22_X1 port map( A1 => n14241, A2 => n36340, B1 => n24792, B2 => 
                           n19901, ZN => n15849);
   U7575 : INV_X1 port map( I => n24674, ZN => n13128);
   U7579 : NAND3_X1 port map( A1 => n958, A2 => n24717, A3 => n24719, ZN => 
                           n30507);
   U7581 : INV_X1 port map( I => n7529, ZN => n24818);
   U7582 : NOR2_X1 port map( A1 => n30554, A2 => n1577, ZN => n30947);
   U7586 : CLKBUF_X2 port map( I => n19294, Z => n36296);
   U7587 : AOI22_X1 port map( A1 => n11053, A2 => n5431, B1 => n33012, B2 => 
                           n24826, ZN => n38044);
   U7590 : NAND2_X1 port map( A1 => n32882, A2 => n24746, ZN => n13735);
   U7591 : NAND2_X1 port map( A1 => n24789, A2 => n20039, ZN => n8428);
   U7595 : NOR2_X1 port map( A1 => n24897, A2 => n38317, ZN => n38475);
   U7598 : INV_X1 port map( I => n21310, ZN => n11169);
   U7599 : INV_X2 port map( I => n7769, ZN => n38317);
   U7603 : BUF_X2 port map( I => n30464, Z => n9921);
   U7604 : NOR3_X1 port map( A1 => n1284, A2 => n24300, A3 => n8581, ZN => 
                           n24185);
   U7607 : INV_X1 port map( I => n6066, ZN => n5261);
   U7609 : INV_X1 port map( I => n7250, ZN => n11319);
   U7612 : OAI21_X1 port map( A1 => n24770, A2 => n8173, B => n5495, ZN => 
                           n5494);
   U7613 : NAND2_X1 port map( A1 => n6491, A2 => n34526, ZN => n31361);
   U7626 : INV_X1 port map( I => n25080, ZN => n25124);
   U7627 : INV_X1 port map( I => n24545, ZN => n24783);
   U7628 : OAI22_X1 port map( A1 => n24798, A2 => n33409, B1 => n24800, B2 => 
                           n24799, ZN => n3878);
   U7630 : NOR2_X1 port map( A1 => n443, A2 => n36920, ZN => n442);
   U7635 : AOI21_X1 port map( A1 => n1122, A2 => n14857, B => n14265, ZN => 
                           n32400);
   U7639 : OAI21_X1 port map( A1 => n37983, A2 => n16196, B => n39279, ZN => 
                           n7248);
   U7640 : INV_X1 port map( I => n24719, ZN => n24721);
   U7642 : NAND2_X1 port map( A1 => n1845, A2 => n933, ZN => n1844);
   U7643 : INV_X1 port map( I => n24417, ZN => n1559);
   U7646 : INV_X1 port map( I => n12233, ZN => n32896);
   U7648 : CLKBUF_X2 port map( I => n24997, Z => n38641);
   U7650 : INV_X1 port map( I => n25284, ZN => n1556);
   U7651 : INV_X1 port map( I => n25272, ZN => n39655);
   U7652 : OAI21_X1 port map( A1 => n17100, A2 => n16540, B => n16539, ZN => 
                           n2530);
   U7662 : NAND2_X1 port map( A1 => n24651, A2 => n24868, ZN => n24652);
   U7664 : NAND2_X1 port map( A1 => n21049, A2 => n24841, ZN => n16746);
   U7666 : INV_X1 port map( I => n25210, ZN => n4796);
   U7669 : INV_X1 port map( I => n25317, ZN => n38430);
   U7671 : INV_X1 port map( I => n25196, ZN => n38712);
   U7674 : INV_X1 port map( I => n32349, ZN => n5433);
   U7675 : INV_X1 port map( I => n20304, ZN => n35472);
   U7680 : INV_X1 port map( I => n36039, ZN => n12251);
   U7684 : NAND2_X1 port map( A1 => n25616, A2 => n18031, ZN => n38625);
   U7687 : INV_X1 port map( I => n18810, ZN => n38425);
   U7692 : NAND2_X1 port map( A1 => n33268, A2 => n25361, ZN => n149);
   U7698 : INV_X2 port map( I => n10055, ZN => n38686);
   U7699 : NAND2_X1 port map( A1 => n36991, A2 => n25513, ZN => n38730);
   U7700 : NOR2_X1 port map( A1 => n31359, A2 => n31358, ZN => n831);
   U7703 : INV_X1 port map( I => n12944, ZN => n12748);
   U7706 : OAI21_X1 port map( A1 => n25527, A2 => n16933, B => n19701, ZN => 
                           n10788);
   U7707 : INV_X1 port map( I => n3451, ZN => n32495);
   U7708 : NAND2_X1 port map( A1 => n25365, A2 => n2576, ZN => n20881);
   U7716 : NOR2_X1 port map( A1 => n25328, A2 => n2803, ZN => n19927);
   U7717 : NOR2_X1 port map( A1 => n1252, A2 => n24963, ZN => n39223);
   U7732 : AOI21_X1 port map( A1 => n1531, A2 => n25692, B => n8014, ZN => 
                           n12779);
   U7733 : NAND2_X1 port map( A1 => n36792, A2 => n16677, ZN => n36475);
   U7734 : NOR2_X1 port map( A1 => n1548, A2 => n32654, ZN => n16739);
   U7737 : NOR2_X1 port map( A1 => n178, A2 => n25670, ZN => n12983);
   U7742 : CLKBUF_X4 port map( I => n15566, Z => n39061);
   U7743 : INV_X2 port map( I => n826, ZN => n21302);
   U7748 : NOR3_X1 port map( A1 => n39061, A2 => n14413, A3 => n13129, ZN => 
                           n18842);
   U7751 : AOI22_X1 port map( A1 => n38732, A2 => n5042, B1 => n13461, B2 => 
                           n36486, ZN => n15790);
   U7754 : CLKBUF_X2 port map( I => n36105, Z => n34583);
   U7756 : OAI21_X1 port map( A1 => n33130, A2 => n21042, B => n39053, ZN => 
                           n25497);
   U7758 : BUF_X2 port map( I => n25322, Z => n25484);
   U7760 : INV_X1 port map( I => n13717, ZN => n35015);
   U7767 : INV_X1 port map( I => n19644, ZN => n12896);
   U7772 : OAI22_X1 port map( A1 => n25603, A2 => n14708, B1 => n8739, B2 => 
                           n10814, ZN => n35467);
   U7773 : NAND2_X1 port map( A1 => n9336, A2 => n25644, ZN => n9335);
   U7775 : AOI21_X1 port map( A1 => n541, A2 => n16114, B => n25517, ZN => 
                           n16113);
   U7777 : NAND3_X1 port map( A1 => n541, A2 => n11874, A3 => n1249, ZN => 
                           n25621);
   U7778 : NAND2_X1 port map( A1 => n16200, A2 => n26042, ZN => n32468);
   U7780 : NOR2_X1 port map( A1 => n926, A2 => n26055, ZN => n13732);
   U7781 : AOI21_X1 port map( A1 => n6844, A2 => n6845, B => n1377, ZN => n3219
                           );
   U7783 : INV_X1 port map( I => n25915, ZN => n5982);
   U7784 : NAND2_X1 port map( A1 => n24535, A2 => n25647, ZN => n33056);
   U7786 : AOI21_X1 port map( A1 => n37336, A2 => n39160, B => n911, ZN => 
                           n38477);
   U7788 : INV_X1 port map( I => n35648, ZN => n26103);
   U7795 : CLKBUF_X2 port map( I => n9743, Z => n424);
   U7797 : INV_X2 port map( I => n12548, ZN => n32690);
   U7798 : CLKBUF_X1 port map( I => n26086, Z => n4772);
   U7799 : INV_X1 port map( I => n25870, ZN => n25871);
   U7800 : NOR3_X1 port map( A1 => n36906, A2 => n7767, A3 => n37393, ZN => 
                           n30283);
   U7802 : OAI21_X1 port map( A1 => n11624, A2 => n11552, B => n18406, ZN => 
                           n11623);
   U7803 : CLKBUF_X2 port map( I => n26092, Z => n33237);
   U7806 : NAND2_X1 port map( A1 => n4512, A2 => n4511, ZN => n37821);
   U7808 : INV_X1 port map( I => n17455, ZN => n16376);
   U7812 : INV_X1 port map( I => n11533, ZN => n13391);
   U7813 : OAI21_X1 port map( A1 => n34206, A2 => n2424, B => n11858, ZN => 
                           n17188);
   U7814 : NOR2_X1 port map( A1 => n26331, A2 => n1240, ZN => n24967);
   U7816 : NAND2_X1 port map( A1 => n9294, A2 => n34743, ZN => n34742);
   U7817 : OAI22_X1 port map( A1 => n12002, A2 => n37072, B1 => n4191, B2 => 
                           n929, ZN => n4189);
   U7820 : INV_X1 port map( I => n19648, ZN => n39183);
   U7823 : INV_X2 port map( I => n37476, ZN => n1506);
   U7825 : CLKBUF_X2 port map( I => n32106, Z => n39793);
   U7827 : INV_X1 port map( I => n16294, ZN => n37448);
   U7829 : CLKBUF_X2 port map( I => n26334, Z => n38279);
   U7841 : CLKBUF_X4 port map( I => n6571, Z => n39172);
   U7844 : CLKBUF_X2 port map( I => n26161, Z => n38753);
   U7846 : INV_X1 port map( I => n26205, ZN => n38028);
   U7850 : INV_X1 port map( I => n32386, ZN => n7726);
   U7853 : CLKBUF_X2 port map( I => n34768, Z => n39032);
   U7857 : NAND2_X1 port map( A1 => n35967, A2 => n14355, ZN => n3351);
   U7860 : NAND2_X1 port map( A1 => n13110, A2 => n39825, ZN => n3368);
   U7862 : INV_X1 port map( I => n19448, ZN => n26830);
   U7867 : INV_X1 port map( I => n26385, ZN => n34648);
   U7869 : NAND3_X1 port map( A1 => n19972, A2 => n1234, A3 => n9117, ZN => 
                           n26907);
   U7871 : INV_X1 port map( I => n26627, ZN => n18226);
   U7873 : INV_X2 port map( I => n26830, ZN => n1231);
   U7876 : INV_X1 port map( I => n26877, ZN => n30724);
   U7879 : NAND2_X1 port map( A1 => n14394, A2 => n1234, ZN => n31220);
   U7880 : CLKBUF_X2 port map( I => n7742, Z => n33279);
   U7881 : INV_X1 port map( I => n10187, ZN => n38775);
   U7882 : AND3_X1 port map( A1 => n10479, A2 => n37289, A3 => n11696, Z => 
                           n37139);
   U7886 : INV_X2 port map( I => n26852, ZN => n26614);
   U7887 : OAI21_X1 port map( A1 => n26909, A2 => n26908, B => n19972, ZN => 
                           n26911);
   U7890 : NAND2_X1 port map( A1 => n14079, A2 => n39564, ZN => n15341);
   U7894 : NAND2_X1 port map( A1 => n38776, A2 => n26709, ZN => n9619);
   U7898 : BUF_X2 port map( I => n26832, Z => n19225);
   U7899 : CLKBUF_X4 port map( I => n26839, Z => n32345);
   U7901 : NAND2_X1 port map( A1 => n30724, A2 => n30725, ZN => n38778);
   U7904 : INV_X1 port map( I => n20704, ZN => n26797);
   U7906 : CLKBUF_X4 port map( I => n18135, Z => n13757);
   U7907 : AOI21_X1 port map( A1 => n26840, A2 => n37103, B => n32345, ZN => 
                           n20754);
   U7908 : OAI21_X1 port map( A1 => n948, A2 => n26696, B => n1495, ZN => 
                           n16708);
   U7910 : NOR2_X1 port map( A1 => n37289, A2 => n11696, ZN => n6312);
   U7911 : CLKBUF_X4 port map( I => n14383, Z => n36344);
   U7917 : CLKBUF_X2 port map( I => n26935, Z => n38120);
   U7918 : OAI21_X1 port map( A1 => n26758, A2 => n12755, B => n12767, ZN => 
                           n12766);
   U7924 : NAND2_X1 port map( A1 => n15411, A2 => n17158, ZN => n11467);
   U7927 : NOR2_X1 port map( A1 => n11696, A2 => n17515, ZN => n13487);
   U7930 : INV_X1 port map( I => n35485, ZN => n37654);
   U7931 : INV_X1 port map( I => n1492, ZN => n21091);
   U7938 : INV_X1 port map( I => n4272, ZN => n37653);
   U7939 : AND3_X1 port map( A1 => n18054, A2 => n36344, A3 => n2158, Z => 
                           n36583);
   U7940 : AND2_X1 port map( A1 => n1092, A2 => n38002, Z => n3962);
   U7942 : CLKBUF_X1 port map( I => n9618, Z => n38577);
   U7943 : NAND3_X1 port map( A1 => n14825, A2 => n16834, A3 => n6615, ZN => 
                           n14824);
   U7945 : NAND2_X1 port map( A1 => n26672, A2 => n3328, ZN => n17260);
   U7946 : CLKBUF_X2 port map( I => n9188, Z => n35282);
   U7948 : INV_X1 port map( I => n27363, ZN => n1484);
   U7956 : OAI21_X1 port map( A1 => n14521, A2 => n19505, B => n26804, ZN => 
                           n19504);
   U7960 : NAND2_X1 port map( A1 => n27278, A2 => n9875, ZN => n38306);
   U7962 : INV_X1 port map( I => n27131, ZN => n19557);
   U7968 : INV_X1 port map( I => n32205, ZN => n27053);
   U7970 : CLKBUF_X1 port map( I => n27213, Z => n38926);
   U7972 : INV_X1 port map( I => n27392, ZN => n13699);
   U7973 : NOR2_X1 port map( A1 => n36989, A2 => n4034, ZN => n27170);
   U7978 : NAND2_X1 port map( A1 => n27150, A2 => n27149, ZN => n32942);
   U7979 : NOR2_X1 port map( A1 => n11162, A2 => n20057, ZN => n9926);
   U7989 : NOR2_X1 port map( A1 => n2035, A2 => n27402, ZN => n11090);
   U7992 : NOR2_X1 port map( A1 => n31875, A2 => n16170, ZN => n37771);
   U7993 : NOR2_X1 port map( A1 => n13278, A2 => n4272, ZN => n27220);
   U7997 : INV_X1 port map( I => n20190, ZN => n27015);
   U7998 : CLKBUF_X4 port map( I => n36177, Z => n35990);
   U7999 : OR3_X1 port map( A1 => n27337, A2 => n19326, A3 => n7096, Z => 
                           n31735);
   U8000 : INV_X2 port map( I => n27320, ZN => n27391);
   U8001 : NAND2_X1 port map( A1 => n5027, A2 => n7096, ZN => n35681);
   U8007 : NAND2_X1 port map( A1 => n14261, A2 => n5675, ZN => n33403);
   U8008 : OAI21_X1 port map( A1 => n39532, A2 => n39531, B => n6191, ZN => 
                           n39730);
   U8010 : NOR2_X1 port map( A1 => n2522, A2 => n1891, ZN => n2304);
   U8012 : OAI21_X1 port map( A1 => n11767, A2 => n36762, B => n27449, ZN => 
                           n8644);
   U8013 : NAND2_X1 port map( A1 => n27232, A2 => n30671, ZN => n18350);
   U8014 : OAI21_X1 port map( A1 => n37801, A2 => n27092, B => n16043, ZN => 
                           n16045);
   U8015 : NAND2_X1 port map( A1 => n32631, A2 => n7312, ZN => n35158);
   U8018 : CLKBUF_X2 port map( I => n5588, Z => n35485);
   U8019 : INV_X1 port map( I => n27304, ZN => n27585);
   U8020 : BUF_X2 port map( I => n27404, Z => n33803);
   U8022 : NAND3_X1 port map( A1 => n34387, A2 => n31875, A3 => n4743, ZN => 
                           n38637);
   U8026 : NAND2_X1 port map( A1 => n27401, A2 => n33335, ZN => n26845);
   U8027 : OAI21_X1 port map( A1 => n38630, A2 => n27314, B => n4434, ZN => 
                           n4490);
   U8028 : INV_X2 port map( I => n6533, ZN => n6534);
   U8033 : NOR2_X1 port map( A1 => n13294, A2 => n39414, ZN => n3921);
   U8038 : NOR2_X1 port map( A1 => n27172, A2 => n19062, ZN => n38144);
   U8049 : CLKBUF_X2 port map( I => n37881, Z => n37499);
   U8052 : INV_X1 port map( I => n31778, ZN => n27531);
   U8054 : CLKBUF_X4 port map( I => n11694, Z => n282);
   U8057 : CLKBUF_X1 port map( I => n27810, Z => n31320);
   U8058 : INV_X1 port map( I => n27725, ZN => n37327);
   U8061 : INV_X1 port map( I => n27712, ZN => n31137);
   U8065 : INV_X1 port map( I => n762, ZN => n6365);
   U8066 : CLKBUF_X2 port map( I => n27498, Z => n37639);
   U8067 : CLKBUF_X2 port map( I => n27566, Z => n34902);
   U8068 : INV_X1 port map( I => n27547, ZN => n11155);
   U8069 : INV_X1 port map( I => n35469, ZN => n37418);
   U8070 : INV_X2 port map( I => n14426, ZN => n1759);
   U8082 : INV_X1 port map( I => n27692, ZN => n6642);
   U8085 : NOR2_X1 port map( A1 => n20053, A2 => n15925, ZN => n5940);
   U8088 : NAND2_X1 port map( A1 => n11512, A2 => n17447, ZN => n15364);
   U8090 : OR2_X1 port map( A1 => n3771, A2 => n3770, Z => n28234);
   U8094 : BUF_X2 port map( I => n20774, Z => n39571);
   U8095 : INV_X2 port map( I => n14399, ZN => n28273);
   U8098 : INV_X1 port map( I => n8078, ZN => n28220);
   U8099 : INV_X1 port map( I => n1212, ZN => n1450);
   U8100 : CLKBUF_X2 port map( I => n8080, Z => n4649);
   U8106 : NAND2_X1 port map( A1 => n288, A2 => n31571, ZN => n37784);
   U8108 : INV_X1 port map( I => n36197, ZN => n36954);
   U8110 : CLKBUF_X1 port map( I => n2980, Z => n2262);
   U8111 : NOR2_X1 port map( A1 => n28079, A2 => n7872, ZN => n28080);
   U8114 : INV_X2 port map( I => n14480, ZN => n16869);
   U8116 : CLKBUF_X2 port map( I => n9516, Z => n156);
   U8122 : NOR2_X1 port map( A1 => n36979, A2 => n14376, ZN => n35146);
   U8123 : NAND2_X1 port map( A1 => n16065, A2 => n28221, ZN => n9702);
   U8126 : CLKBUF_X4 port map( I => n33958, Z => n12260);
   U8127 : NAND2_X1 port map( A1 => n6643, A2 => n16065, ZN => n9024);
   U8129 : NOR2_X1 port map( A1 => n28212, A2 => n12192, ZN => n37642);
   U8131 : NOR3_X1 port map( A1 => n6733, A2 => n28089, A3 => n8149, ZN => 
                           n5160);
   U8133 : NAND2_X1 port map( A1 => n2982, A2 => n2740, ZN => n2981);
   U8134 : INV_X2 port map( I => n16363, ZN => n17532);
   U8136 : NAND2_X1 port map( A1 => n20663, A2 => n28269, ZN => n20470);
   U8138 : INV_X1 port map( I => n28049, ZN => n28139);
   U8145 : CLKBUF_X2 port map( I => n3158, Z => n37451);
   U8146 : CLKBUF_X2 port map( I => n16500, Z => n16154);
   U8147 : NOR2_X1 port map( A1 => n28249, A2 => n3032, ZN => n30366);
   U8148 : NOR2_X1 port map( A1 => n35694, A2 => n16576, ZN => n18379);
   U8151 : OAI21_X1 port map( A1 => n28217, A2 => n987, B => n16971, ZN => 
                           n28083);
   U8153 : AOI21_X1 port map( A1 => n1200, A2 => n12406, B => n1074, ZN => 
                           n27743);
   U8157 : OAI21_X1 port map( A1 => n10756, A2 => n13059, B => n33405, ZN => 
                           n5864);
   U8160 : NAND2_X1 port map( A1 => n15691, A2 => n15693, ZN => n34480);
   U8165 : INV_X1 port map( I => n28753, ZN => n31924);
   U8170 : NAND2_X1 port map( A1 => n3598, A2 => n28575, ZN => n2704);
   U8171 : NAND3_X1 port map( A1 => n34516, A2 => n27983, A3 => n34515, ZN => 
                           n38155);
   U8172 : NAND2_X1 port map( A1 => n35357, A2 => n28807, ZN => n8637);
   U8174 : NAND2_X1 port map( A1 => n28546, A2 => n28729, ZN => n9056);
   U8175 : CLKBUF_X1 port map( I => n28591, Z => n35888);
   U8177 : AOI21_X1 port map( A1 => n36788, A2 => n35173, B => n28611, ZN => 
                           n12891);
   U8184 : NOR2_X1 port map( A1 => n32759, A2 => n1882, ZN => n28708);
   U8185 : OAI21_X1 port map( A1 => n19946, A2 => n34170, B => n4724, ZN => 
                           n28091);
   U8192 : INV_X2 port map( I => n28620, ZN => n28339);
   U8194 : NOR2_X1 port map( A1 => n1874, A2 => n30581, ZN => n34305);
   U8195 : INV_X2 port map( I => n33765, ZN => n19349);
   U8200 : NAND2_X1 port map( A1 => n28758, A2 => n978, ZN => n9017);
   U8204 : NOR2_X1 port map( A1 => n12237, A2 => n5383, ZN => n2333);
   U8205 : CLKBUF_X4 port map( I => n9597, Z => n2022);
   U8207 : AND2_X1 port map( A1 => n13727, A2 => n13726, Z => n38172);
   U8209 : INV_X1 port map( I => n34651, ZN => n31147);
   U8210 : NOR3_X1 port map( A1 => n30953, A2 => n977, A3 => n28746, ZN => 
                           n18626);
   U8212 : NOR2_X1 port map( A1 => n28312, A2 => n5418, ZN => n4969);
   U8213 : INV_X2 port map( I => n28496, ZN => n7454);
   U8214 : INV_X1 port map( I => n28559, ZN => n28655);
   U8216 : INV_X1 port map( I => n1184, ZN => n34739);
   U8218 : OAI21_X1 port map( A1 => n13237, A2 => n34915, B => n28758, ZN => 
                           n8449);
   U8220 : NAND2_X1 port map( A1 => n38857, A2 => n38856, ZN => n28565);
   U8225 : NAND2_X1 port map( A1 => n13891, A2 => n17800, ZN => n13893);
   U8231 : NAND2_X1 port map( A1 => n28605, A2 => n8349, ZN => n10758);
   U8232 : CLKBUF_X2 port map( I => n7429, Z => n37956);
   U8233 : CLKBUF_X2 port map( I => n29057, Z => n39631);
   U8234 : CLKBUF_X2 port map( I => n28971, Z => n19405);
   U8236 : NAND2_X1 port map( A1 => n35804, A2 => n35805, ZN => n13965);
   U8238 : NOR3_X1 port map( A1 => n39332, A2 => n13598, A3 => n31888, ZN => 
                           n38608);
   U8239 : CLKBUF_X4 port map( I => n29144, Z => n36905);
   U8240 : NAND2_X1 port map( A1 => n1184, A2 => n9106, ZN => n9109);
   U8242 : INV_X1 port map( I => n20465, ZN => n38679);
   U8243 : CLKBUF_X2 port map( I => n15157, Z => n15156);
   U8248 : INV_X1 port map( I => n29645, ZN => n37304);
   U8252 : NOR2_X1 port map( A1 => n29200, A2 => n15153, ZN => n11885);
   U8254 : OAI21_X1 port map( A1 => n30238, A2 => n9394, B => n15651, ZN => 
                           n33267);
   U8255 : NAND2_X1 port map( A1 => n14449, A2 => n32906, ZN => n29265);
   U8257 : NAND2_X1 port map( A1 => n29459, A2 => n36275, ZN => n36893);
   U8258 : INV_X1 port map( I => n19896, ZN => n20429);
   U8262 : INV_X1 port map( I => n33368, ZN => n18947);
   U8264 : CLKBUF_X2 port map( I => n14403, Z => n8677);
   U8265 : INV_X2 port map( I => n14158, ZN => n1183);
   U8266 : NAND2_X1 port map( A1 => n1183, A2 => n14600, ZN => n29861);
   U8269 : CLKBUF_X2 port map( I => n12940, Z => n39585);
   U8271 : INV_X2 port map( I => n29059, ZN => n39392);
   U8276 : NAND2_X1 port map( A1 => n29452, A2 => n9993, ZN => n28900);
   U8279 : INV_X2 port map( I => n37061, ZN => n21269);
   U8281 : NOR2_X1 port map( A1 => n19734, A2 => n29642, ZN => n36102);
   U8283 : AOI21_X1 port map( A1 => n28864, A2 => n14428, B => n18947, ZN => 
                           n9885);
   U8285 : CLKBUF_X4 port map( I => n17698, Z => n1962);
   U8288 : NOR2_X1 port map( A1 => n10610, A2 => n29815, ZN => n39017);
   U8289 : INV_X1 port map( I => n16224, ZN => n29938);
   U8292 : OAI21_X1 port map( A1 => n16060, A2 => n8529, B => n4255, ZN => 
                           n37531);
   U8295 : NAND2_X1 port map( A1 => n1181, A2 => n29185, ZN => n14184);
   U8297 : CLKBUF_X2 port map( I => n29381, Z => n12876);
   U8301 : NAND2_X1 port map( A1 => n2792, A2 => n15189, ZN => n7015);
   U8302 : INV_X2 port map( I => n4083, ZN => n19476);
   U8307 : OAI21_X1 port map( A1 => n28822, A2 => n30046, B => n28825, ZN => 
                           n11404);
   U8309 : NAND2_X1 port map( A1 => n19162, A2 => n14892, ZN => n30237);
   U8310 : NAND2_X1 port map( A1 => n38163, A2 => n30128, ZN => n11845);
   U8311 : CLKBUF_X1 port map( I => n29532, Z => n39178);
   U8312 : NAND2_X1 port map( A1 => n29437, A2 => n18502, ZN => n29434);
   U8313 : NAND2_X1 port map( A1 => n36101, A2 => n36100, ZN => n19175);
   U8321 : INV_X1 port map( I => n29971, ZN => n32129);
   U8324 : NOR2_X1 port map( A1 => n11845, A2 => n17192, ZN => n35625);
   U8325 : CLKBUF_X1 port map( I => n29535, Z => n37605);
   U8326 : NOR2_X1 port map( A1 => n19090, A2 => n16233, ZN => n29275);
   U8329 : INV_X1 port map( I => n29410, ZN => n29416);
   U8335 : OAI21_X1 port map( A1 => n18793, A2 => n18794, B => n33128, ZN => 
                           n32452);
   U8338 : BUF_X2 port map( I => n18241, Z => n3896);
   U8343 : CLKBUF_X1 port map( I => Key(140), Z => n29522);
   U8345 : INV_X1 port map( I => n29680, ZN => n34239);
   U8346 : AOI22_X1 port map( A1 => n13277, A2 => n29355, B1 => n29356, B2 => 
                           n13981, ZN => n37262);
   U8350 : OAI21_X1 port map( A1 => n32768, A2 => n32767, B => n29362, ZN => 
                           n37273);
   U8355 : INV_X1 port map( I => n29334, ZN => n39482);
   U8356 : INV_X1 port map( I => n29442, ZN => n1377);
   U8361 : AOI21_X1 port map( A1 => n29790, A2 => n29791, B => n37781, ZN => 
                           n20939);
   U8362 : INV_X1 port map( I => n19674, ZN => n1051);
   U8367 : OR2_X1 port map( A1 => n14349, A2 => n11344, Z => n37113);
   U8370 : NAND2_X1 port map( A1 => n15573, A2 => n6067, ZN => n37114);
   U8373 : AND2_X2 port map( A1 => n24698, A2 => n24903, Z => n37115);
   U8381 : OR2_X2 port map( A1 => n11404, A2 => n35183, Z => n37117);
   U8383 : AND2_X2 port map( A1 => n6876, A2 => n35228, Z => n37118);
   U8384 : AND2_X1 port map( A1 => n5314, A2 => n16246, Z => n37119);
   U8389 : AND3_X1 port map( A1 => n28149, A2 => n37754, A3 => n1076, Z => 
                           n37120);
   U8391 : XNOR2_X1 port map( A1 => n15102, A2 => n19851, ZN => n37121);
   U8393 : OR2_X1 port map( A1 => n24169, A2 => n20457, Z => n37122);
   U8396 : AND2_X1 port map( A1 => n1408, A2 => n29780, Z => n37123);
   U8397 : AND2_X2 port map( A1 => n32472, A2 => n35705, Z => n37125);
   U8399 : OR2_X1 port map( A1 => n14560, A2 => n38229, Z => n37127);
   U8400 : OR2_X2 port map( A1 => n38636, A2 => n38635, Z => n37129);
   U8409 : OR2_X1 port map( A1 => n2761, A2 => n35299, Z => n37130);
   U8411 : OR2_X1 port map( A1 => n446, A2 => n14212, Z => n37132);
   U8414 : OR2_X2 port map( A1 => n2741, A2 => n37896, Z => n37134);
   U8415 : AND2_X2 port map( A1 => n31005, A2 => n33933, Z => n37137);
   U8418 : OR2_X1 port map( A1 => n22920, A2 => n9725, Z => n37138);
   U8419 : AND2_X1 port map( A1 => n22995, A2 => n19288, Z => n37141);
   U8420 : AND2_X1 port map( A1 => n27284, A2 => n30851, Z => n37143);
   U8422 : AND2_X1 port map( A1 => n38578, A2 => n27267, Z => n37144);
   U8426 : AND3_X1 port map( A1 => n15209, A2 => n1393, A3 => n29571, Z => 
                           n37145);
   U8428 : AND2_X2 port map( A1 => n29346, A2 => n29241, Z => n37146);
   U8430 : XOR2_X1 port map( A1 => n27851, A2 => n19940, Z => n37147);
   U8432 : XNOR2_X1 port map( A1 => n23933, A2 => n29432, ZN => n37148);
   U8436 : XOR2_X1 port map( A1 => n17310, A2 => n19763, Z => n37149);
   U8437 : AND2_X1 port map( A1 => n26329, A2 => n26092, Z => n37150);
   U8438 : INV_X1 port map( I => n15466, ZN => n21930);
   U8440 : OR2_X2 port map( A1 => n38507, A2 => n32691, Z => n37151);
   U8442 : AND2_X2 port map( A1 => n19434, A2 => n19238, Z => n37152);
   U8447 : OR2_X1 port map( A1 => n26901, A2 => n34005, Z => n37153);
   U8449 : AND2_X1 port map( A1 => n21893, A2 => n21894, Z => n37155);
   U8450 : AND2_X1 port map( A1 => n8155, A2 => n18870, Z => n37156);
   U8452 : NOR2_X1 port map( A1 => n1445, A2 => n17755, ZN => n37159);
   U8457 : AND2_X2 port map( A1 => n39061, A2 => n20838, Z => n37160);
   U8458 : AND2_X2 port map( A1 => n9875, A2 => n15284, Z => n37162);
   U8459 : AND2_X2 port map( A1 => n22317, A2 => n22316, Z => n37163);
   U8461 : NOR2_X1 port map( A1 => n38202, A2 => n20056, ZN => n37164);
   U8465 : CLKBUF_X2 port map( I => n19326, Z => n5027);
   U8468 : INV_X1 port map( I => n10006, ZN => n14428);
   U8472 : AND2_X1 port map( A1 => n25566, A2 => n5166, Z => n37165);
   U8474 : AND3_X1 port map( A1 => n24310, A2 => n1289, A3 => n250, Z => n37166
                           );
   U8477 : AND2_X1 port map( A1 => n23128, A2 => n5380, Z => n37167);
   U8479 : OR3_X1 port map( A1 => n34783, A2 => n24234, A3 => n30311, Z => 
                           n37168);
   U8482 : AND2_X1 port map( A1 => n5124, A2 => n5063, Z => n37169);
   U8484 : AND2_X1 port map( A1 => n39406, A2 => n35137, Z => n37171);
   U8491 : NOR2_X1 port map( A1 => n33949, A2 => n13286, ZN => n37173);
   U8492 : AND3_X1 port map( A1 => n1016, A2 => n26032, A3 => n3345, Z => 
                           n37175);
   U8496 : OR2_X1 port map( A1 => n21618, A2 => n1049, Z => n37176);
   U8499 : AND2_X1 port map( A1 => n16860, A2 => n39676, Z => n37178);
   U8500 : AND2_X1 port map( A1 => n3631, A2 => n18815, Z => n37179);
   U8501 : OR2_X2 port map( A1 => n32134, A2 => n37025, Z => n37183);
   U8502 : OR2_X2 port map( A1 => n25587, A2 => n4603, Z => n37184);
   U8503 : AND2_X1 port map( A1 => n18667, A2 => n777, Z => n37185);
   U8506 : AND2_X1 port map( A1 => n4542, A2 => n8692, Z => n37190);
   U8508 : OR2_X1 port map( A1 => n18114, A2 => n6337, Z => n37193);
   U8509 : XNOR2_X1 port map( A1 => n22492, A2 => n30101, ZN => n37194);
   U8510 : XNOR2_X1 port map( A1 => n27499, A2 => n28910, ZN => n37195);
   U8513 : INV_X1 port map( I => n18757, ZN => n19850);
   U8514 : CLKBUF_X2 port map( I => n18757, Z => n16302);
   U8519 : INV_X1 port map( I => n19677, ZN => n37443);
   U8520 : OR2_X1 port map( A1 => n17931, A2 => n13029, Z => n37196);
   U8526 : XNOR2_X1 port map( A1 => n8312, A2 => n10558, ZN => n37197);
   U8527 : OR2_X2 port map( A1 => n27153, A2 => n27408, Z => n37198);
   U8530 : CLKBUF_X2 port map( I => n21871, Z => n19650);
   U8532 : INV_X1 port map( I => n21871, ZN => n21756);
   U8534 : XOR2_X1 port map( A1 => Plaintext(64), A2 => Key(64), Z => n37200);
   U8535 : AND2_X2 port map( A1 => n5089, A2 => n34644, Z => n37201);
   U8536 : AND2_X1 port map( A1 => n28726, A2 => n12237, Z => n37203);
   U8538 : AND3_X2 port map( A1 => n34516, A2 => n27983, A3 => n34515, Z => 
                           n37204);
   U8540 : AND2_X1 port map( A1 => n27397, A2 => n2522, Z => n37205);
   U8544 : INV_X1 port map( I => n5126, ZN => n30621);
   U8547 : INV_X2 port map( I => n12754, ZN => n21942);
   U8555 : XNOR2_X1 port map( A1 => n9151, A2 => n7018, ZN => n37206);
   U8560 : NOR2_X1 port map( A1 => n20346, A2 => n7644, ZN => n37207);
   U8561 : AND2_X2 port map( A1 => n23227, A2 => n23533, Z => n37208);
   U8562 : AND2_X2 port map( A1 => n12617, A2 => n19481, Z => n37209);
   U8566 : OR2_X2 port map( A1 => n30845, A2 => n7529, Z => n37210);
   U8567 : INV_X2 port map( I => n31307, ZN => n12943);
   U8571 : INV_X1 port map( I => n38948, ZN => n15145);
   U8575 : AND3_X1 port map( A1 => n19740, A2 => n37819, A3 => n37613, Z => 
                           n37211);
   U8579 : OR2_X2 port map( A1 => n10980, A2 => n16502, Z => n37212);
   U8586 : CLKBUF_X1 port map( I => n10980, Z => n36395);
   U8590 : INV_X1 port map( I => n27820, ZN => n37855);
   U8591 : XNOR2_X1 port map( A1 => n22584, A2 => n5235, ZN => n37214);
   U8592 : NOR2_X1 port map( A1 => n3510, A2 => n32956, ZN => n39714);
   U8593 : NAND2_X1 port map( A1 => n39714, A2 => n24912, ZN => n37215);
   U8595 : AND2_X2 port map( A1 => n17074, A2 => n10632, Z => n37216);
   U8597 : OR2_X2 port map( A1 => n21370, A2 => n21369, Z => n37217);
   U8608 : INV_X1 port map( I => n23201, ZN => n19524);
   U8609 : INV_X1 port map( I => n34200, ZN => n7266);
   U8618 : XOR2_X1 port map( A1 => n5835, A2 => n35286, Z => n37218);
   U8622 : OR2_X1 port map( A1 => n23192, A2 => n1147, Z => n37219);
   U8625 : OR2_X1 port map( A1 => n9835, A2 => n23475, Z => n37220);
   U8626 : XOR2_X1 port map( A1 => n23952, A2 => n30122, Z => n37221);
   U8630 : XNOR2_X1 port map( A1 => n32239, A2 => n16320, ZN => n37222);
   U8634 : XNOR2_X1 port map( A1 => n11372, A2 => n39183, ZN => n37223);
   U8643 : XNOR2_X1 port map( A1 => n23888, A2 => n23808, ZN => n37224);
   U8646 : AND2_X1 port map( A1 => n1290, A2 => n39194, Z => n37225);
   U8647 : AND2_X1 port map( A1 => n22295, A2 => n16880, Z => n37226);
   U8651 : XNOR2_X1 port map( A1 => n6156, A2 => n30451, ZN => n37227);
   U8652 : NAND2_X1 port map( A1 => n37016, A2 => n37411, ZN => n37228);
   U8657 : INV_X1 port map( I => n25574, ZN => n1113);
   U8660 : AND2_X2 port map( A1 => n24369, A2 => n24192, Z => n37229);
   U8665 : XNOR2_X1 port map( A1 => n7920, A2 => n31869, ZN => n37230);
   U8673 : XNOR2_X1 port map( A1 => n4302, A2 => n36171, ZN => n37231);
   U8674 : XOR2_X1 port map( A1 => n37816, A2 => n39044, Z => n37232);
   U8675 : INV_X1 port map( I => n39681, ZN => n19565);
   U8677 : INV_X2 port map( I => n31722, ZN => n16990);
   U8678 : OR2_X1 port map( A1 => n3760, A2 => n30464, Z => n37233);
   U8679 : XOR2_X1 port map( A1 => n11321, A2 => n19919, Z => n37234);
   U8680 : INV_X2 port map( I => n5634, ZN => n37983);
   U8681 : CLKBUF_X1 port map( I => n36798, Z => n39048);
   U8689 : CLKBUF_X2 port map( I => n21301, Z => n15541);
   U8694 : INV_X1 port map( I => n21301, ZN => n37553);
   U8699 : INV_X2 port map( I => n840, ZN => n19889);
   U8702 : XNOR2_X1 port map( A1 => n5118, A2 => n6877, ZN => n37235);
   U8703 : XOR2_X1 port map( A1 => n34469, A2 => n29371, Z => n37236);
   U8713 : OR2_X2 port map( A1 => n33949, A2 => n25322, Z => n37237);
   U8714 : OR2_X2 port map( A1 => n14045, A2 => n730, Z => n37238);
   U8730 : AND2_X2 port map( A1 => n11003, A2 => n840, Z => n37239);
   U8731 : INV_X1 port map( I => n17237, ZN => n36391);
   U8742 : CLKBUF_X4 port map( I => n17237, Z => n38238);
   U8747 : XNOR2_X1 port map( A1 => n21044, A2 => n27634, ZN => n37240);
   U8797 : INV_X2 port map( I => n1235, ZN => n11513);
   U8800 : AND2_X2 port map( A1 => n8988, A2 => n8798, Z => n37241);
   U8801 : XNOR2_X1 port map( A1 => n27499, A2 => n27178, ZN => n37242);
   U8805 : XNOR2_X1 port map( A1 => n27681, A2 => n27680, ZN => n37243);
   U8807 : OR2_X1 port map( A1 => n33491, A2 => n35260, Z => n37244);
   U8809 : OR2_X2 port map( A1 => n9658, A2 => n32563, Z => n37245);
   U8810 : XNOR2_X1 port map( A1 => n20713, A2 => n6133, ZN => n37247);
   U8814 : OR3_X1 port map( A1 => n28683, A2 => n1414, A3 => n1196, Z => n37248
                           );
   U8821 : AND2_X1 port map( A1 => n28698, A2 => n28695, Z => n37249);
   U8822 : CLKBUF_X4 port map( I => n26906, Z => n1234);
   U8823 : INV_X1 port map( I => n13891, ZN => n6703);
   U8825 : INV_X1 port map( I => n11375, ZN => n14152);
   U8833 : INV_X1 port map( I => n14411, ZN => n13492);
   U8837 : NOR2_X1 port map( A1 => n10461, A2 => n35427, ZN => n37250);
   U8843 : AND2_X2 port map( A1 => n20056, A2 => n15047, Z => n37251);
   U8845 : XNOR2_X1 port map( A1 => n15745, A2 => n1710, ZN => n37252);
   U8848 : INV_X1 port map( I => n29247, ZN => n4905);
   U8850 : OR2_X1 port map( A1 => n31595, A2 => n30057, Z => n37253);
   U8851 : XNOR2_X1 port map( A1 => n29095, A2 => n19683, ZN => n37254);
   U8852 : AND2_X1 port map( A1 => n36935, A2 => n31554, Z => n37255);
   U8861 : AND2_X2 port map( A1 => n11491, A2 => n11492, Z => n37256);
   U8866 : INV_X1 port map( I => n10422, ZN => n14449);
   U8869 : AND2_X1 port map( A1 => n3159, A2 => n32932, Z => n37257);
   U8870 : INV_X1 port map( I => n30221, ZN => n30158);
   U8871 : AND2_X1 port map( A1 => n29627, A2 => n29626, Z => n37258);
   U8885 : XOR2_X1 port map( A1 => n13248, A2 => n13246, Z => n37259);
   U8887 : NOR3_X2 port map( A1 => n38542, A2 => n8491, A3 => n35684, ZN => 
                           n33737);
   U8889 : XOR2_X1 port map( A1 => n31775, A2 => n29282, Z => n34586);
   U8891 : NAND2_X2 port map( A1 => n35885, A2 => n3795, ZN => n31775);
   U8894 : XOR2_X1 port map( A1 => n15532, A2 => n37260, Z => n33701);
   U8895 : XOR2_X1 port map( A1 => n23973, A2 => n37261, Z => n37260);
   U8896 : NAND2_X2 port map( A1 => n3076, A2 => n31861, ZN => n31637);
   U8901 : XOR2_X1 port map( A1 => n37262, A2 => n1717, Z => Ciphertext(30));
   U8902 : XOR2_X1 port map( A1 => n4622, A2 => n37112, Z => n34165);
   U8905 : NAND2_X2 port map( A1 => n25377, A2 => n36900, ZN => n4622);
   U8906 : XOR2_X1 port map( A1 => n23700, A2 => n13074, Z => n13871);
   U8908 : XNOR2_X1 port map( A1 => n23832, A2 => n23938, ZN => n23700);
   U8909 : NAND2_X1 port map( A1 => n10404, A2 => n34685, ZN => n25370);
   U8912 : NAND2_X2 port map( A1 => n16767, A2 => n36897, ZN => n34685);
   U8914 : INV_X2 port map( I => n11145, ZN => n25513);
   U8923 : NAND2_X2 port map( A1 => n37346, A2 => n32942, ZN => n34838);
   U8927 : OAI22_X2 port map( A1 => n32255, A2 => n8221, B1 => n8223, B2 => 
                           n20648, ZN => n37378);
   U8931 : XOR2_X1 port map( A1 => n22619, A2 => n22759, Z => n8068);
   U8932 : XOR2_X1 port map( A1 => n5171, A2 => n22371, Z => n22759);
   U8934 : CLKBUF_X4 port map( I => n15218, Z => n37589);
   U8938 : NAND2_X2 port map( A1 => n29845, A2 => n37263, ZN => n2346);
   U8939 : NAND3_X2 port map( A1 => n29908, A2 => n29954, A3 => n29863, ZN => 
                           n37263);
   U8941 : XOR2_X1 port map( A1 => n30856, A2 => n8729, Z => n28970);
   U8943 : AOI21_X2 port map( A1 => n15829, A2 => n19690, B => n24219, ZN => 
                           n24565);
   U8950 : XNOR2_X1 port map( A1 => n9930, A2 => n28982, ZN => n29066);
   U8951 : NAND2_X2 port map( A1 => n4196, A2 => n4197, ZN => n28982);
   U8958 : NAND2_X1 port map( A1 => n4745, A2 => n4746, ZN => n33036);
   U8963 : BUF_X4 port map( I => n19857, Z => n37264);
   U8966 : NAND2_X1 port map( A1 => n12065, A2 => n37604, ZN => n18469);
   U8967 : XOR2_X1 port map( A1 => n15442, A2 => n37053, Z => n11927);
   U8969 : INV_X2 port map( I => n36743, ZN => n37053);
   U8973 : XOR2_X1 port map( A1 => n18012, A2 => n13155, Z => n36743);
   U8975 : NOR2_X2 port map( A1 => n38911, A2 => n2886, ZN => n37031);
   U8980 : NAND2_X2 port map( A1 => n37265, A2 => n39179, ZN => n7542);
   U8982 : NOR2_X2 port map( A1 => n36307, A2 => n36306, ZN => n37265);
   U8983 : XOR2_X1 port map( A1 => n37381, A2 => n10592, Z => n36435);
   U8984 : NAND2_X2 port map( A1 => n27233, A2 => n12306, ZN => n27434);
   U8990 : NAND2_X2 port map( A1 => n35321, A2 => n3136, ZN => n27233);
   U8993 : NAND2_X2 port map( A1 => n1294, A2 => n2182, ZN => n37266);
   U8994 : NAND2_X2 port map( A1 => n7034, A2 => n7033, ZN => n24746);
   U8997 : INV_X2 port map( I => n14353, ZN => n14668);
   U9000 : NAND2_X2 port map( A1 => n17926, A2 => n14354, ZN => n14353);
   U9001 : INV_X2 port map( I => n31673, ZN => n37267);
   U9002 : XOR2_X1 port map( A1 => n37268, A2 => n12014, Z => n35796);
   U9007 : XOR2_X1 port map( A1 => n30653, A2 => n31073, Z => n37268);
   U9008 : XOR2_X1 port map( A1 => n10792, A2 => n25303, Z => n25102);
   U9009 : OAI22_X2 port map( A1 => n24128, A2 => n18114, B1 => n24127, B2 => 
                           n6337, ZN => n10792);
   U9014 : NAND2_X2 port map( A1 => n910, A2 => n11034, ZN => n2865);
   U9015 : OAI22_X2 port map( A1 => n7513, A2 => n11548, B1 => n25365, B2 => 
                           n36345, ZN => n11034);
   U9016 : OAI21_X1 port map( A1 => n1140, A2 => n18090, B => n23299, ZN => 
                           n31052);
   U9020 : NAND2_X2 port map( A1 => n27357, A2 => n35198, ZN => n27066);
   U9021 : NAND2_X2 port map( A1 => n6376, A2 => n5560, ZN => n27357);
   U9025 : XOR2_X1 port map( A1 => n12296, A2 => n37269, Z => n35645);
   U9026 : XOR2_X1 port map( A1 => n25083, A2 => n37498, Z => n37269);
   U9028 : XOR2_X1 port map( A1 => n22549, A2 => n22647, Z => n22736);
   U9030 : NAND2_X2 port map( A1 => n22105, A2 => n22104, ZN => n22647);
   U9032 : NAND2_X1 port map( A1 => n38079, A2 => n19061, ZN => n4463);
   U9033 : NAND2_X2 port map( A1 => n37270, A2 => n5625, ZN => n5623);
   U9034 : NAND2_X2 port map( A1 => n31702, A2 => n5361, ZN => n32354);
   U9037 : OR2_X1 port map( A1 => n7317, A2 => n35138, Z => n2940);
   U9045 : NAND3_X1 port map( A1 => n25999, A2 => n2940, A3 => n19121, ZN => 
                           n38342);
   U9060 : AOI22_X2 port map( A1 => n1604, A2 => n37271, B1 => n37480, B2 => 
                           n33289, ZN => n15829);
   U9061 : NAND2_X1 port map( A1 => n35954, A2 => n12950, ZN => n37271);
   U9064 : XOR2_X1 port map( A1 => n22475, A2 => n9873, Z => n7942);
   U9071 : AOI21_X2 port map( A1 => n5878, A2 => n5877, B => n5874, ZN => 
                           n22475);
   U9073 : INV_X2 port map( I => n28163, ZN => n2877);
   U9075 : XOR2_X1 port map( A1 => n11730, A2 => n27748, Z => n31880);
   U9084 : OAI22_X1 port map( A1 => n961, A2 => n20418, B1 => n32471, B2 => 
                           n23399, ZN => n22873);
   U9085 : OAI21_X2 port map( A1 => n18413, A2 => n37272, B => n1056, ZN => 
                           n33476);
   U9087 : NOR2_X1 port map( A1 => n29998, A2 => n30041, ZN => n37272);
   U9091 : XOR2_X1 port map( A1 => n37273, A2 => n29363, Z => Ciphertext(33));
   U9093 : AOI21_X2 port map( A1 => n4075, A2 => n34652, B => n37274, ZN => 
                           n4073);
   U9096 : AND2_X1 port map( A1 => n14089, A2 => n17210, Z => n17459);
   U9097 : NOR2_X2 port map( A1 => n37275, A2 => n3624, ZN => n24813);
   U9098 : XOR2_X1 port map( A1 => n21096, A2 => n34809, Z => n19458);
   U9100 : XOR2_X1 port map( A1 => n37280, A2 => n13568, Z => n36822);
   U9106 : XOR2_X1 port map( A1 => n8865, A2 => n557, Z => n37280);
   U9108 : OAI21_X1 port map( A1 => n27951, A2 => n20739, B => n12303, ZN => 
                           n37895);
   U9109 : XOR2_X1 port map( A1 => n36522, A2 => n19933, Z => n12935);
   U9112 : NAND2_X2 port map( A1 => n8234, A2 => n8235, ZN => n36522);
   U9115 : XOR2_X1 port map( A1 => n27668, A2 => n18548, Z => n18547);
   U9118 : XOR2_X1 port map( A1 => n4934, A2 => n27802, Z => n27668);
   U9119 : INV_X2 port map( I => n26026, ZN => n26525);
   U9120 : OR2_X1 port map( A1 => n28661, A2 => n28660, Z => n34176);
   U9123 : XOR2_X1 port map( A1 => n26514, A2 => n10965, Z => n26375);
   U9126 : NOR2_X2 port map( A1 => n14722, A2 => n21307, ZN => n26514);
   U9130 : NAND2_X2 port map( A1 => n9916, A2 => n25936, ZN => n25812);
   U9131 : NAND3_X2 port map( A1 => n10936, A2 => n10935, A3 => n10313, ZN => 
                           n9916);
   U9132 : NAND2_X2 port map( A1 => n33546, A2 => n15667, ZN => n27508);
   U9133 : NOR2_X2 port map( A1 => n37281, A2 => n36801, ZN => n37522);
   U9134 : AOI21_X2 port map( A1 => n24227, A2 => n18573, B => n4601, ZN => 
                           n10648);
   U9136 : NAND2_X2 port map( A1 => n1029, A2 => n2634, ZN => n24227);
   U9141 : NAND2_X2 port map( A1 => n19438, A2 => n25567, ZN => n5356);
   U9147 : NAND2_X1 port map( A1 => n5354, A2 => n25724, ZN => n19438);
   U9149 : XOR2_X1 port map( A1 => n37593, A2 => n11105, Z => n2068);
   U9152 : NAND2_X2 port map( A1 => n10269, A2 => n10270, ZN => n37593);
   U9155 : XOR2_X1 port map( A1 => n37282, A2 => n33758, Z => n39326);
   U9158 : XOR2_X1 port map( A1 => n37855, A2 => n3114, Z => n37282);
   U9161 : AOI22_X2 port map( A1 => n37915, A2 => n37914, B1 => n38319, B2 => 
                           n30237, ZN => n38204);
   U9164 : NAND2_X2 port map( A1 => n34853, A2 => n27306, ZN => n26790);
   U9165 : XOR2_X1 port map( A1 => n34237, A2 => n26485, Z => n38968);
   U9166 : NAND3_X2 port map( A1 => n36458, A2 => n38632, A3 => n38633, ZN => 
                           n26485);
   U9168 : XOR2_X1 port map( A1 => n27655, A2 => n27654, Z => n11358);
   U9169 : XOR2_X1 port map( A1 => n27637, A2 => n27729, Z => n27655);
   U9170 : NAND2_X2 port map( A1 => n38766, A2 => n37283, ZN => n28400);
   U9171 : AOI22_X2 port map( A1 => n10084, A2 => n38666, B1 => n1202, B2 => 
                           n12038, ZN => n37283);
   U9173 : XOR2_X1 port map( A1 => n29147, A2 => n6758, Z => n29258);
   U9179 : NAND2_X2 port map( A1 => n28304, A2 => n28305, ZN => n6758);
   U9181 : XOR2_X1 port map( A1 => n27668, A2 => n7416, Z => n7864);
   U9183 : XOR2_X1 port map( A1 => n27504, A2 => n27492, Z => n7416);
   U9194 : NOR3_X2 port map( A1 => n33395, A2 => n586, A3 => n26053, ZN => 
                           n34310);
   U9196 : XNOR2_X1 port map( A1 => n25087, A2 => n14643, ZN => n38109);
   U9201 : OAI22_X2 port map( A1 => n37284, A2 => n33963, B1 => n10568, B2 => 
                           n20251, ZN => n20274);
   U9202 : NOR2_X2 port map( A1 => n14539, A2 => n18007, ZN => n37284);
   U9205 : NOR3_X1 port map( A1 => n26018, A2 => n2349, A3 => n26054, ZN => 
                           n2621);
   U9206 : NAND2_X2 port map( A1 => n9788, A2 => n37711, ZN => n26018);
   U9207 : NAND4_X2 port map( A1 => n9806, A2 => n12452, A3 => n30401, A4 => 
                           n31495, ZN => n38067);
   U9209 : NAND2_X1 port map( A1 => n35381, A2 => n6191, ZN => n35380);
   U9210 : NOR2_X1 port map( A1 => n38051, A2 => n19151, ZN => n29499);
   U9212 : XOR2_X1 port map( A1 => n15091, A2 => n15090, Z => n17425);
   U9214 : XOR2_X1 port map( A1 => n26536, A2 => n26539, Z => n8021);
   U9215 : XOR2_X1 port map( A1 => n5241, A2 => n26163, Z => n26539);
   U9218 : OR2_X1 port map( A1 => n27218, A2 => n15616, Z => n13231);
   U9220 : NAND2_X1 port map( A1 => n28724, A2 => n28360, ZN => n37285);
   U9222 : XOR2_X1 port map( A1 => n26160, A2 => n26484, Z => n13426);
   U9223 : XOR2_X1 port map( A1 => n38514, A2 => n26448, Z => n26160);
   U9225 : NAND2_X1 port map( A1 => n32861, A2 => n37002, ZN => n38482);
   U9228 : NOR2_X2 port map( A1 => n37287, A2 => n37286, ZN => n31769);
   U9234 : INV_X2 port map( I => n26893, ZN => n37289);
   U9236 : XOR2_X1 port map( A1 => n27612, A2 => n27469, Z => n37668);
   U9242 : XOR2_X1 port map( A1 => n37833, A2 => n5900, Z => n27612);
   U9245 : OAI22_X2 port map( A1 => n26700, A2 => n19951, B1 => n36244, B2 => 
                           n10440, ZN => n26178);
   U9246 : XOR2_X1 port map( A1 => n37290, A2 => n7734, Z => n9133);
   U9248 : XOR2_X1 port map( A1 => n23716, A2 => n23725, Z => n37290);
   U9249 : AOI21_X2 port map( A1 => n5906, A2 => n1440, B => n37291, ZN => 
                           n6426);
   U9250 : OAI22_X1 port map( A1 => n5905, A2 => n8522, B1 => n18696, B2 => 
                           n5266, ZN => n37291);
   U9251 : NOR2_X1 port map( A1 => n920, A2 => n37632, ZN => n11567);
   U9257 : AOI22_X2 port map( A1 => n38237, A2 => n38236, B1 => n12657, B2 => 
                           n18043, ZN => n37632);
   U9259 : NAND3_X2 port map( A1 => n38093, A2 => n27203, A3 => n37292, ZN => 
                           n27792);
   U9264 : NAND3_X1 port map( A1 => n16946, A2 => n27201, A3 => n14881, ZN => 
                           n37292);
   U9265 : NOR2_X2 port map( A1 => n39291, A2 => n25921, ZN => n34339);
   U9268 : NAND2_X2 port map( A1 => n5908, A2 => n26215, ZN => n25921);
   U9274 : NOR2_X2 port map( A1 => n14469, A2 => n37293, ZN => n7424);
   U9276 : OAI22_X2 port map( A1 => n26858, A2 => n8103, B1 => n11651, B2 => 
                           n11652, ZN => n37293);
   U9277 : INV_X4 port map( I => n23381, ZN => n33864);
   U9280 : OAI22_X2 port map( A1 => n4099, A2 => n4100, B1 => n4102, B2 => 
                           n23057, ZN => n23381);
   U9281 : XOR2_X1 port map( A1 => n22538, A2 => n37294, Z => n37459);
   U9285 : XOR2_X1 port map( A1 => n22534, A2 => n22533, Z => n37294);
   U9291 : BUF_X2 port map( I => n28772, Z => n37295);
   U9294 : XOR2_X1 port map( A1 => n4077, A2 => n26417, Z => n3161);
   U9297 : NAND2_X2 port map( A1 => n7317, A2 => n35138, ZN => n26000);
   U9303 : OR2_X2 port map( A1 => n5929, A2 => n8882, Z => n8089);
   U9307 : NAND3_X2 port map( A1 => n38481, A2 => n38482, A3 => n26789, ZN => 
                           n27542);
   U9308 : OAI21_X2 port map( A1 => n6585, A2 => n24175, B => n24228, ZN => 
                           n37601);
   U9310 : XOR2_X1 port map( A1 => n9122, A2 => n23882, Z => n9121);
   U9311 : XOR2_X1 port map( A1 => n37932, A2 => n23890, Z => n23882);
   U9316 : INV_X2 port map( I => n2030, ZN => n38282);
   U9318 : XOR2_X1 port map( A1 => n37296, A2 => n25323, Z => n25174);
   U9320 : NOR2_X2 port map( A1 => n17474, A2 => n17473, ZN => n25323);
   U9323 : INV_X2 port map( I => n24857, ZN => n37296);
   U9325 : XOR2_X1 port map( A1 => n37297, A2 => n18359, Z => n32128);
   U9326 : XOR2_X1 port map( A1 => n22627, A2 => n22628, Z => n37297);
   U9331 : OAI22_X2 port map( A1 => n33359, A2 => n17989, B1 => n4200, B2 => 
                           n17499, ZN => n4199);
   U9333 : NAND2_X1 port map( A1 => n38063, A2 => n29626, ZN => n37298);
   U9335 : NAND3_X2 port map( A1 => n28326, A2 => n30389, A3 => n28325, ZN => 
                           n3927);
   U9339 : NAND2_X2 port map( A1 => n36860, A2 => n7872, ZN => n30389);
   U9340 : XOR2_X1 port map( A1 => n26527, A2 => n37299, Z => n2754);
   U9343 : XOR2_X1 port map( A1 => n1506, A2 => n26587, Z => n37299);
   U9344 : NOR2_X2 port map( A1 => n1244, A2 => n26055, ZN => n26053);
   U9346 : OAI21_X2 port map( A1 => n1320, A2 => n8491, B => n22935, ZN => 
                           n13542);
   U9348 : INV_X2 port map( I => n31558, ZN => n8491);
   U9349 : XOR2_X1 port map( A1 => n628, A2 => n31559, Z => n31558);
   U9359 : NAND2_X2 port map( A1 => n15763, A2 => n21091, ZN => n4579);
   U9361 : OAI22_X2 port map( A1 => n12065, A2 => n7305, B1 => n2140, B2 => 
                           n33952, ZN => n15763);
   U9362 : NAND2_X2 port map( A1 => n21067, A2 => n21066, ZN => n23885);
   U9363 : NAND2_X2 port map( A1 => n23520, A2 => n10024, ZN => n21067);
   U9364 : XOR2_X1 port map( A1 => n8021, A2 => n8020, Z => n19298);
   U9366 : XOR2_X1 port map( A1 => n9861, A2 => n19751, Z => n33924);
   U9369 : OAI22_X2 port map( A1 => n24254, A2 => n34055, B1 => n34141, B2 => 
                           n21049, ZN => n9861);
   U9370 : XOR2_X1 port map( A1 => n9548, A2 => n9549, Z => n9383);
   U9371 : NAND3_X2 port map( A1 => n35145, A2 => n2495, A3 => n2496, ZN => 
                           n692);
   U9373 : NAND2_X2 port map( A1 => n20458, A2 => n15258, ZN => n37732);
   U9380 : NAND2_X1 port map( A1 => n4001, A2 => n1545, ZN => n4468);
   U9385 : XOR2_X1 port map( A1 => n37301, A2 => n38712, Z => n38711);
   U9388 : XOR2_X1 port map( A1 => n37357, A2 => n25083, Z => n37301);
   U9390 : XOR2_X1 port map( A1 => n16743, A2 => n31767, Z => n34365);
   U9391 : NAND2_X2 port map( A1 => n36467, A2 => n8485, ZN => n16743);
   U9393 : NAND3_X2 port map( A1 => n946, A2 => n26695, A3 => n10338, ZN => 
                           n142);
   U9397 : NAND2_X2 port map( A1 => n37550, A2 => n5533, ZN => n5024);
   U9398 : NAND2_X1 port map( A1 => n22323, A2 => n22322, ZN => n37302);
   U9400 : OAI22_X2 port map( A1 => n28618, A2 => n30858, B1 => n2500, B2 => 
                           n28655, ZN => n29137);
   U9401 : NOR2_X2 port map( A1 => n2678, A2 => n11034, ZN => n25925);
   U9405 : NAND2_X2 port map( A1 => n6965, A2 => n32615, ZN => n2678);
   U9407 : NAND2_X2 port map( A1 => n37305, A2 => n3722, ZN => n34603);
   U9408 : NAND3_X2 port map( A1 => n36251, A2 => n5309, A3 => n1653, ZN => 
                           n37305);
   U9410 : BUF_X2 port map( I => n37730, Z => n37306);
   U9412 : XOR2_X1 port map( A1 => n27631, A2 => n37307, Z => n31778);
   U9413 : XOR2_X1 port map( A1 => n10582, A2 => n25201, Z => n10583);
   U9414 : INV_X2 port map( I => n30279, ZN => n19466);
   U9415 : NOR2_X2 port map( A1 => n13201, A2 => n13200, ZN => n25133);
   U9418 : OR2_X1 port map( A1 => n37308, A2 => n23461, Z => n3174);
   U9419 : OAI21_X2 port map( A1 => n37310, A2 => n37309, B => n12711, ZN => 
                           n39521);
   U9420 : INV_X2 port map( I => n28680, ZN => n37311);
   U9422 : XOR2_X1 port map( A1 => n27677, A2 => n8874, Z => n8873);
   U9424 : XOR2_X1 port map( A1 => n8875, A2 => n39442, Z => n8874);
   U9426 : XOR2_X1 port map( A1 => n37313, A2 => n17646, Z => Ciphertext(168));
   U9432 : AOI22_X1 port map( A1 => n30135, A2 => n30144, B1 => n30134, B2 => 
                           n30133, ZN => n37313);
   U9434 : NOR2_X2 port map( A1 => n19657, A2 => n37251, ZN => n27686);
   U9439 : XOR2_X1 port map( A1 => n37314, A2 => n23921, Z => n32472);
   U9440 : XOR2_X1 port map( A1 => n5441, A2 => n5442, Z => n37314);
   U9442 : OAI21_X2 port map( A1 => n2464, A2 => n21148, B => n37315, ZN => 
                           n19279);
   U9449 : OAI21_X2 port map( A1 => n5572, A2 => n33077, B => n37316, ZN => 
                           n37315);
   U9450 : NOR2_X2 port map( A1 => n32507, A2 => n37125, ZN => n37316);
   U9452 : XOR2_X1 port map( A1 => n2618, A2 => n37317, Z => n30982);
   U9453 : XOR2_X1 port map( A1 => n34149, A2 => n25314, Z => n37317);
   U9454 : NAND2_X2 port map( A1 => n26608, A2 => n21317, ZN => n27449);
   U9455 : XOR2_X1 port map( A1 => n14312, A2 => n11215, Z => n5322);
   U9457 : XOR2_X1 port map( A1 => n4956, A2 => n23832, Z => n14312);
   U9458 : NAND2_X2 port map( A1 => n27263, A2 => n36969, ZN => n27265);
   U9459 : XOR2_X1 port map( A1 => n12196, A2 => n34250, Z => n15412);
   U9460 : OAI22_X2 port map( A1 => n37732, A2 => n21124, B1 => n37229, B2 => 
                           n20083, ZN => n24650);
   U9461 : AOI22_X2 port map( A1 => n9071, A2 => n9073, B1 => n18845, B2 => 
                           n355, ZN => n37498);
   U9462 : INV_X1 port map( I => n28719, ZN => n37561);
   U9463 : NOR2_X2 port map( A1 => n29413, A2 => n29409, ZN => n20724);
   U9468 : AOI22_X2 port map( A1 => n29379, A2 => n6314, B1 => n17295, B2 => 
                           n16876, ZN => n29413);
   U9470 : INV_X2 port map( I => n4322, ZN => n31192);
   U9472 : NAND2_X2 port map( A1 => n25384, A2 => n12996, ZN => n4322);
   U9475 : NOR3_X2 port map( A1 => n31483, A2 => n37318, A3 => n32504, ZN => 
                           n37989);
   U9479 : INV_X1 port map( I => n38941, ZN => n29600);
   U9489 : OAI21_X2 port map( A1 => n5035, A2 => n35663, B => n3923, ZN => 
                           n35998);
   U9499 : AOI22_X2 port map( A1 => n39448, A2 => n37598, B1 => n19719, B2 => 
                           n36203, ZN => n35663);
   U9505 : AOI22_X2 port map( A1 => n2462, A2 => n2461, B1 => n25437, B2 => 
                           n25562, ZN => n8096);
   U9506 : OAI22_X2 port map( A1 => n6505, A2 => n28376, B1 => n32012, B2 => 
                           n28448, ZN => n32866);
   U9509 : NOR2_X2 port map( A1 => n3899, A2 => n39020, ZN => n28376);
   U9510 : NOR2_X2 port map( A1 => n36583, A2 => n36582, ZN => n998);
   U9511 : AND2_X1 port map( A1 => n6892, A2 => n12527, Z => n28336);
   U9514 : XNOR2_X1 port map( A1 => n25272, A2 => n2064, ZN => n37324);
   U9516 : BUF_X4 port map( I => n18967, Z => n34000);
   U9523 : NAND3_X2 port map( A1 => n37321, A2 => n4543, A3 => n37320, ZN => 
                           n24034);
   U9525 : NAND2_X2 port map( A1 => n13603, A2 => n33080, ZN => n37321);
   U9532 : NOR2_X2 port map( A1 => n39303, A2 => n37108, ZN => n22950);
   U9534 : XOR2_X1 port map( A1 => n2065, A2 => n37324, Z => n37662);
   U9536 : XOR2_X1 port map( A1 => n37325, A2 => n287, Z => n1961);
   U9538 : XOR2_X1 port map( A1 => n38133, A2 => n33715, Z => n37325);
   U9539 : XOR2_X1 port map( A1 => n37326, A2 => n14031, Z => n38470);
   U9540 : XOR2_X1 port map( A1 => n37427, A2 => n37327, Z => n37326);
   U9541 : OAI21_X2 port map( A1 => n13536, A2 => n13538, B => n13535, ZN => 
                           n37393);
   U9545 : XOR2_X1 port map( A1 => n15686, A2 => n37328, Z => n16186);
   U9546 : XOR2_X1 port map( A1 => n25208, A2 => n17595, Z => n37328);
   U9547 : NAND3_X2 port map( A1 => n37330, A2 => n14232, A3 => n37329, ZN => 
                           n39382);
   U9548 : INV_X2 port map( I => n28272, ZN => n37329);
   U9550 : NAND2_X2 port map( A1 => n1759, A2 => n11628, ZN => n37330);
   U9551 : NAND2_X2 port map( A1 => n11252, A2 => n11251, ZN => n6904);
   U9553 : INV_X2 port map( I => n37331, ZN => n38084);
   U9566 : NAND2_X2 port map( A1 => n13780, A2 => n11613, ZN => n37331);
   U9573 : INV_X1 port map( I => n3441, ZN => n39501);
   U9575 : NOR2_X2 port map( A1 => n11560, A2 => n37332, ZN => n6559);
   U9588 : OAI22_X2 port map( A1 => n23338, A2 => n21293, B1 => n12870, B2 => 
                           n23474, ZN => n37332);
   U9592 : OAI21_X2 port map( A1 => n13206, A2 => n5569, B => n37333, ZN => 
                           n17508);
   U9597 : NAND2_X2 port map( A1 => n15743, A2 => n32590, ZN => n37333);
   U9599 : XOR2_X1 port map( A1 => n23786, A2 => n23785, Z => n6092);
   U9601 : NAND2_X2 port map( A1 => n26003, A2 => n38507, ZN => n25854);
   U9603 : NAND2_X2 port map( A1 => n37334, A2 => n34762, ZN => n3903);
   U9605 : BUF_X2 port map( I => n22849, Z => n37335);
   U9607 : AOI21_X2 port map( A1 => n13690, A2 => n10883, B => n1429, ZN => 
                           n9692);
   U9611 : INV_X4 port map( I => n27624, ZN => n35694);
   U9612 : BUF_X2 port map( I => n39061, Z => n37336);
   U9614 : NOR2_X2 port map( A1 => n38755, A2 => n38939, ZN => n38211);
   U9615 : XOR2_X1 port map( A1 => n23965, A2 => n11383, Z => n1971);
   U9621 : NAND2_X2 port map( A1 => n2950, A2 => n23345, ZN => n23965);
   U9624 : NOR2_X1 port map( A1 => n39696, A2 => n18144, ZN => n38906);
   U9625 : XOR2_X1 port map( A1 => n37337, A2 => n7729, Z => n27903);
   U9626 : XOR2_X1 port map( A1 => n37540, A2 => n1859, Z => n37337);
   U9627 : NAND3_X2 port map( A1 => n17754, A2 => n27147, A3 => n27434, ZN => 
                           n37346);
   U9628 : OR2_X1 port map( A1 => n24699, A2 => n24698, Z => n35735);
   U9637 : NAND2_X2 port map( A1 => n24712, A2 => n24903, ZN => n24699);
   U9640 : NAND2_X2 port map( A1 => n10907, A2 => n28686, ZN => n18035);
   U9641 : NAND2_X2 port map( A1 => n35496, A2 => n12349, ZN => n10907);
   U9645 : NOR2_X2 port map( A1 => n12925, A2 => n22899, ZN => n22902);
   U9646 : INV_X4 port map( I => n39127, ZN => n13491);
   U9649 : INV_X2 port map( I => n17727, ZN => n1659);
   U9652 : NAND2_X2 port map( A1 => n9391, A2 => n9392, ZN => n17727);
   U9653 : NOR2_X2 port map( A1 => n11676, A2 => n27910, ZN => n12038);
   U9662 : NAND2_X2 port map( A1 => n37669, A2 => n25608, ZN => n19258);
   U9667 : AOI22_X2 port map( A1 => n25872, A2 => n32520, B1 => n25871, B2 => 
                           n17501, ZN => n37742);
   U9668 : XOR2_X1 port map( A1 => n26340, A2 => n26227, Z => n12014);
   U9671 : NOR2_X2 port map( A1 => n12709, A2 => n12708, ZN => n26340);
   U9672 : BUF_X2 port map( I => n39442, Z => n37338);
   U9674 : NAND3_X2 port map( A1 => n37339, A2 => n5902, A3 => n5901, ZN => 
                           n17696);
   U9676 : XOR2_X1 port map( A1 => n20044, A2 => n19343, Z => n31673);
   U9679 : XOR2_X1 port map( A1 => n12299, A2 => n33120, Z => n15988);
   U9681 : XOR2_X1 port map( A1 => n12805, A2 => n37340, Z => n33934);
   U9682 : XOR2_X1 port map( A1 => n39047, A2 => n22436, Z => n37340);
   U9686 : XOR2_X1 port map( A1 => n25204, A2 => n39582, Z => n38736);
   U9689 : BUF_X2 port map( I => n10054, Z => n37341);
   U9694 : XOR2_X1 port map( A1 => n27526, A2 => n27813, Z => n3474);
   U9695 : XOR2_X1 port map( A1 => n13802, A2 => n27617, Z => n27526);
   U9697 : NAND2_X2 port map( A1 => n38604, A2 => n4997, ZN => n14234);
   U9699 : XOR2_X1 port map( A1 => n31293, A2 => n26279, Z => n10668);
   U9702 : NAND2_X2 port map( A1 => n38122, A2 => n34499, ZN => n26279);
   U9709 : INV_X2 port map( I => n37342, ZN => n3873);
   U9711 : XNOR2_X1 port map( A1 => n3732, A2 => n38706, ZN => n37342);
   U9713 : NAND2_X2 port map( A1 => n37343, A2 => n22952, ZN => n10480);
   U9715 : OAI21_X2 port map( A1 => n22948, A2 => n17459, B => n23138, ZN => 
                           n37343);
   U9716 : XOR2_X1 port map( A1 => n38639, A2 => n37344, Z => n18732);
   U9718 : XOR2_X1 port map( A1 => n10562, A2 => n8723, Z => n37344);
   U9720 : INV_X2 port map( I => n34969, ZN => n27411);
   U9722 : NAND3_X2 port map( A1 => n7362, A2 => n25428, A3 => n20358, ZN => 
                           n11148);
   U9723 : XOR2_X1 port map( A1 => n37345, A2 => n26403, Z => n26410);
   U9724 : XOR2_X1 port map( A1 => n26405, A2 => n26402, Z => n37345);
   U9725 : NAND2_X2 port map( A1 => n10480, A2 => n8668, ZN => n23620);
   U9727 : OR2_X1 port map( A1 => n23572, A2 => n12154, Z => n32362);
   U9728 : OAI21_X2 port map( A1 => n28129, A2 => n31942, B => n10287, ZN => 
                           n28464);
   U9734 : XOR2_X1 port map( A1 => n22720, A2 => n17612, Z => n37382);
   U9735 : XOR2_X1 port map( A1 => n16226, A2 => n39528, Z => n17612);
   U9739 : XOR2_X1 port map( A1 => n37347, A2 => n11072, Z => n3827);
   U9742 : XOR2_X1 port map( A1 => n14454, A2 => n23985, Z => n35601);
   U9743 : OAI21_X2 port map( A1 => n24182, A2 => n19739, B => n1587, ZN => 
                           n12279);
   U9749 : NOR2_X1 port map( A1 => n12138, A2 => n35164, ZN => n19739);
   U9753 : INV_X2 port map( I => n29377, ZN => n31521);
   U9754 : NAND2_X2 port map( A1 => n3697, A2 => n35952, ZN => n38801);
   U9756 : NAND2_X2 port map( A1 => n33529, A2 => n4184, ZN => n3697);
   U9759 : INV_X1 port map( I => n39788, ZN => n7224);
   U9761 : AND2_X1 port map( A1 => n39788, A2 => n13414, Z => n39803);
   U9764 : NAND2_X1 port map( A1 => n29611, A2 => n32980, ZN => n20126);
   U9767 : NOR2_X1 port map( A1 => n25564, A2 => n25563, ZN => n37584);
   U9773 : NAND2_X2 port map( A1 => n12363, A2 => n12364, ZN => n33132);
   U9774 : XOR2_X1 port map( A1 => n26242, A2 => n26243, Z => n37347);
   U9775 : OAI22_X2 port map( A1 => n4433, A2 => n35887, B1 => n299, B2 => 
                           n4013, ZN => n38416);
   U9778 : AOI22_X2 port map( A1 => n19495, A2 => n1254, B1 => n9815, B2 => 
                           n33491, ZN => n4013);
   U9779 : AOI22_X2 port map( A1 => n37244, A2 => n37348, B1 => n25597, B2 => 
                           n20515, ZN => n20381);
   U9780 : NOR2_X2 port map( A1 => n37350, A2 => n5503, ZN => n37559);
   U9781 : AOI21_X2 port map( A1 => n13437, A2 => n6604, B => n5392, ZN => 
                           n37350);
   U9782 : NOR3_X2 port map( A1 => n31607, A2 => n36844, A3 => n28246, ZN => 
                           n15087);
   U9783 : OAI21_X2 port map( A1 => n4152, A2 => n4153, B => n28102, ZN => 
                           n20020);
   U9794 : OAI22_X2 port map( A1 => n36574, A2 => n36575, B1 => n15183, B2 => 
                           n3356, ZN => n32253);
   U9796 : XOR2_X1 port map( A1 => n19024, A2 => n6177, Z => n17486);
   U9798 : AOI22_X2 port map( A1 => n32109, A2 => n13731, B1 => n34524, B2 => 
                           n25424, ZN => n4660);
   U9801 : XOR2_X1 port map( A1 => n25239, A2 => n19064, Z => n20365);
   U9802 : XOR2_X1 port map( A1 => n17653, A2 => n1261, Z => n19064);
   U9805 : XOR2_X1 port map( A1 => n13199, A2 => n3475, Z => n35987);
   U9806 : OR2_X1 port map( A1 => n23202, A2 => n2430, Z => n11704);
   U9809 : BUF_X2 port map( I => n686, Z => n37351);
   U9817 : NAND2_X2 port map( A1 => n38049, A2 => n36927, ZN => n23873);
   U9828 : XOR2_X1 port map( A1 => n20698, A2 => n7728, Z => n25268);
   U9834 : OAI22_X2 port map( A1 => n20806, A2 => n20696, B1 => n19507, B2 => 
                           n20807, ZN => n20698);
   U9837 : XOR2_X1 port map( A1 => n37353, A2 => n37352, Z => n791);
   U9843 : XOR2_X1 port map( A1 => n36461, A2 => n1374, Z => n37353);
   U9844 : NAND2_X1 port map( A1 => n35809, A2 => n29898, ZN => n19540);
   U9847 : NOR2_X2 port map( A1 => n38408, A2 => n1627, ZN => n37354);
   U9848 : NOR2_X1 port map( A1 => n37356, A2 => n30087, ZN => n30084);
   U9859 : BUF_X2 port map( I => n34564, Z => n37357);
   U9860 : NAND2_X2 port map( A1 => n39499, A2 => n8196, ZN => n13400);
   U9863 : OAI21_X1 port map( A1 => n33516, A2 => n12218, B => n1198, ZN => 
                           n38804);
   U9870 : XOR2_X1 port map( A1 => n8404, A2 => n8403, Z => n17755);
   U9872 : XOR2_X1 port map( A1 => n27748, A2 => n27716, Z => n8404);
   U9875 : NAND2_X2 port map( A1 => n4388, A2 => n21980, ZN => n37358);
   U9876 : NAND2_X2 port map( A1 => n37942, A2 => n37359, ZN => n29270);
   U9877 : NAND2_X2 port map( A1 => n37360, A2 => n21021, ZN => n495);
   U9878 : AOI22_X2 port map( A1 => n37549, A2 => n11336, B1 => n11339, B2 => 
                           n1093, ZN => n37360);
   U9882 : XOR2_X1 port map( A1 => n30950, A2 => n1668, Z => n17854);
   U9883 : NAND3_X1 port map( A1 => n1170, A2 => n6623, A3 => n18897, ZN => 
                           n7270);
   U9884 : NAND2_X2 port map( A1 => n35570, A2 => n37361, ZN => n12168);
   U9886 : NOR2_X2 port map( A1 => n33912, A2 => n33913, ZN => n37361);
   U9891 : AOI22_X2 port map( A1 => n1027, A2 => n24556, B1 => n24528, B2 => 
                           n12159, ZN => n39120);
   U9892 : NOR2_X2 port map( A1 => n24811, A2 => n12159, ZN => n24556);
   U9893 : XOR2_X1 port map( A1 => n11369, A2 => n37362, Z => n14332);
   U9897 : XOR2_X1 port map( A1 => n25302, A2 => n33005, Z => n37362);
   U9902 : NAND2_X2 port map( A1 => n20966, A2 => n37363, ZN => n28396);
   U9903 : NAND3_X1 port map( A1 => n11353, A2 => n9534, A3 => n27666, ZN => 
                           n37363);
   U9905 : NAND2_X1 port map( A1 => n11820, A2 => n9369, ZN => n33203);
   U9906 : NAND2_X2 port map( A1 => n11818, A2 => n37798, ZN => n11820);
   U9907 : XOR2_X1 port map( A1 => n22686, A2 => n22688, Z => n16755);
   U9908 : XOR2_X1 port map( A1 => n22657, A2 => n22776, Z => n22688);
   U9912 : NOR2_X2 port map( A1 => n15433, A2 => n15434, ZN => n15368);
   U9913 : NOR2_X2 port map( A1 => n30485, A2 => n3718, ZN => n15433);
   U9914 : NAND2_X2 port map( A1 => n37364, A2 => n16369, ZN => n10570);
   U9917 : NAND3_X2 port map( A1 => n23116, A2 => n23117, A3 => n12289, ZN => 
                           n37364);
   U9925 : OR2_X1 port map( A1 => n39678, A2 => n5227, Z => n13016);
   U9926 : NAND2_X2 port map( A1 => n20507, A2 => n37365, ZN => n9030);
   U9927 : INV_X2 port map( I => n37366, ZN => n20541);
   U9928 : XNOR2_X1 port map( A1 => n10390, A2 => n10391, ZN => n37366);
   U9930 : XOR2_X1 port map( A1 => n37367, A2 => n23954, Z => n2229);
   U9931 : XOR2_X1 port map( A1 => n14345, A2 => n18160, Z => n37367);
   U9938 : NAND2_X1 port map( A1 => n10764, A2 => n37746, ZN => n5326);
   U9940 : AOI22_X2 port map( A1 => n37177, A2 => n37368, B1 => n6496, B2 => 
                           n37021, ZN => n17980);
   U9941 : INV_X2 port map( I => n30000, ZN => n37368);
   U9943 : XOR2_X1 port map( A1 => n37369, A2 => n21226, Z => Ciphertext(5));
   U9944 : AOI22_X1 port map( A1 => n9807, A2 => n29209, B1 => n18039, B2 => 
                           n11972, ZN => n37369);
   U9948 : NAND3_X2 port map( A1 => n39402, A2 => n32235, A3 => n37370, ZN => 
                           n14193);
   U9951 : NAND3_X1 port map( A1 => n941, A2 => n18603, A3 => n34120, ZN => 
                           n37370);
   U9955 : NAND2_X2 port map( A1 => n15586, A2 => n37371, ZN => n32765);
   U9960 : NOR2_X2 port map( A1 => n39712, A2 => n39713, ZN => n37371);
   U9974 : INV_X2 port map( I => n36058, ZN => n19593);
   U9975 : NOR2_X2 port map( A1 => n31626, A2 => n26135, ZN => n37372);
   U9976 : NOR2_X1 port map( A1 => n6246, A2 => n4211, ZN => n37373);
   U9977 : XOR2_X1 port map( A1 => n31043, A2 => n881, Z => n28025);
   U9980 : XOR2_X1 port map( A1 => n37650, A2 => n11349, Z => n11482);
   U9982 : AND2_X1 port map( A1 => n37103, A2 => n26839, Z => n21171);
   U9983 : XOR2_X1 port map( A1 => n10221, A2 => n9151, Z => n26208);
   U9984 : NAND2_X2 port map( A1 => n6219, A2 => n1851, ZN => n9151);
   U9988 : XOR2_X1 port map( A1 => n38703, A2 => n39698, Z => n31582);
   U9989 : XOR2_X1 port map( A1 => n19289, A2 => n28821, Z => n26566);
   U9992 : OAI21_X2 port map( A1 => n20612, A2 => n20611, B => n11848, ZN => 
                           n8699);
   U9993 : NAND2_X2 port map( A1 => n39227, A2 => n38203, ZN => n28430);
   U9994 : NAND2_X1 port map( A1 => n28267, A2 => n1206, ZN => n18665);
   U9995 : XOR2_X1 port map( A1 => n37379, A2 => n5801, Z => n14751);
   U9996 : XOR2_X1 port map( A1 => n25161, A2 => n5800, Z => n37379);
   U10001 : XOR2_X1 port map( A1 => n27655, A2 => n11564, Z => n11563);
   U10006 : XOR2_X1 port map( A1 => n25115, A2 => n24985, Z => n25072);
   U10007 : OAI22_X2 port map( A1 => n11199, A2 => n11198, B1 => n1842, B2 => 
                           n24528, ZN => n25115);
   U10010 : INV_X2 port map( I => n29204, ZN => n29208);
   U10012 : XOR2_X1 port map( A1 => n33921, A2 => n37380, Z => n36730);
   U10017 : INV_X1 port map( I => n19894, ZN => n37380);
   U10018 : NAND2_X2 port map( A1 => n39077, A2 => n25451, ZN => n37730);
   U10019 : NOR2_X1 port map( A1 => n18077, A2 => n10004, ZN => n25045);
   U10020 : BUF_X4 port map( I => n11676, Z => n38666);
   U10023 : INV_X2 port map( I => n7099, ZN => n19465);
   U10027 : XNOR2_X1 port map( A1 => n7102, A2 => n7100, ZN => n7099);
   U10029 : NAND2_X2 port map( A1 => n18929, A2 => n5061, ZN => n22296);
   U10030 : NAND2_X2 port map( A1 => n37559, A2 => n5504, ZN => n18929);
   U10044 : XOR2_X1 port map( A1 => n37053, A2 => n3330, Z => n37381);
   U10047 : XOR2_X1 port map( A1 => n33533, A2 => n27864, Z => n27598);
   U10048 : NAND2_X2 port map( A1 => n39565, A2 => n12017, ZN => n33533);
   U10053 : XOR2_X1 port map( A1 => n36756, A2 => n37382, Z => n14381);
   U10059 : XOR2_X1 port map( A1 => n13977, A2 => n23917, Z => n6988);
   U10063 : XOR2_X1 port map( A1 => n35181, A2 => n39209, Z => n23917);
   U10067 : INV_X2 port map( I => n37383, ZN => n25611);
   U10070 : XNOR2_X1 port map( A1 => n10615, A2 => n1896, ZN => n37383);
   U10071 : OR2_X1 port map( A1 => n32898, A2 => n35686, Z => n36280);
   U10072 : NOR2_X1 port map( A1 => n27299, A2 => n34717, ZN => n37385);
   U10074 : XOR2_X1 port map( A1 => n26460, A2 => n26498, Z => n26150);
   U10075 : NAND2_X2 port map( A1 => n9983, A2 => n34481, ZN => n26460);
   U10078 : NOR2_X2 port map( A1 => n4824, A2 => n38779, ZN => n13534);
   U10081 : OAI22_X2 port map( A1 => n14736, A2 => n14696, B1 => n7904, B2 => 
                           n27902, ZN => n38220);
   U10082 : AOI22_X2 port map( A1 => n985, A2 => n1208, B1 => n759, B2 => n1439
                           , ZN => n27902);
   U10084 : XOR2_X1 port map( A1 => n19642, A2 => n14264, Z => n27712);
   U10087 : NAND2_X2 port map( A1 => n35037, A2 => n9491, ZN => n14264);
   U10091 : XOR2_X1 port map( A1 => n11372, A2 => n39073, Z => n2106);
   U10097 : NAND2_X2 port map( A1 => n18890, A2 => n18889, ZN => n39073);
   U10099 : NAND3_X2 port map( A1 => n21979, A2 => n21978, A3 => n19654, ZN => 
                           n22586);
   U10108 : NAND2_X2 port map( A1 => n36525, A2 => n37386, ZN => n12527);
   U10113 : AOI22_X2 port map( A1 => n39399, A2 => n28115, B1 => n15993, B2 => 
                           n13457, ZN => n37386);
   U10127 : NOR2_X2 port map( A1 => n37387, A2 => n21356, ZN => n22497);
   U10128 : AOI21_X2 port map( A1 => n21354, A2 => n39368, B => n39716, ZN => 
                           n37387);
   U10132 : NOR2_X2 port map( A1 => n21666, A2 => n21436, ZN => n21359);
   U10133 : XOR2_X1 port map( A1 => n27793, A2 => n27795, Z => n15723);
   U10136 : XOR2_X1 port map( A1 => n27776, A2 => n38964, Z => n27793);
   U10146 : INV_X1 port map( I => n10992, ZN => n37453);
   U10150 : INV_X1 port map( I => n37388, ZN => n5817);
   U10157 : INV_X4 port map( I => n20597, ZN => n978);
   U10158 : NAND2_X2 port map( A1 => n10720, A2 => n2023, ZN => n20597);
   U10159 : NOR2_X2 port map( A1 => n35192, A2 => n38614, ZN => n11108);
   U10163 : NAND2_X2 port map( A1 => n37516, A2 => n6860, ZN => n38614);
   U10164 : NAND2_X2 port map( A1 => n30191, A2 => n30241, ZN => n9173);
   U10173 : INV_X2 port map( I => n35893, ZN => n37389);
   U10174 : OR2_X1 port map( A1 => n35128, A2 => n37389, Z => n38634);
   U10178 : NOR2_X2 port map( A1 => n16576, A2 => n28153, ZN => n28004);
   U10182 : XOR2_X1 port map( A1 => n16342, A2 => n24049, Z => n31636);
   U10189 : INV_X2 port map( I => n3903, ZN => n28666);
   U10190 : NOR3_X2 port map( A1 => n9676, A2 => n37390, A3 => n14160, ZN => 
                           n37952);
   U10195 : NOR2_X2 port map( A1 => n11717, A2 => n28402, ZN => n28772);
   U10196 : OAI21_X2 port map( A1 => n7984, A2 => n32186, B => n7983, ZN => 
                           n11717);
   U10199 : XOR2_X1 port map( A1 => n7848, A2 => n30090, Z => n2036);
   U10201 : NAND2_X2 port map( A1 => n37719, A2 => n38818, ZN => n7848);
   U10202 : XOR2_X1 port map( A1 => n37391, A2 => n27784, Z => n11823);
   U10204 : XOR2_X1 port map( A1 => n9162, A2 => n36861, Z => n37391);
   U10206 : INV_X4 port map( I => n15573, ZN => n37981);
   U10207 : XNOR2_X1 port map( A1 => n19187, A2 => n33439, ZN => n37394);
   U10208 : NOR2_X2 port map( A1 => n37392, A2 => n7880, ZN => n7882);
   U10209 : XOR2_X1 port map( A1 => n32994, A2 => n37394, Z => n34764);
   U10214 : NAND2_X2 port map( A1 => n37396, A2 => n37395, ZN => n34141);
   U10224 : INV_X2 port map( I => n24639, ZN => n37395);
   U10225 : INV_X2 port map( I => n34906, ZN => n37396);
   U10230 : XOR2_X1 port map( A1 => n10526, A2 => n9611, Z => n37738);
   U10231 : NAND2_X2 port map( A1 => n1919, A2 => n1917, ZN => n10526);
   U10232 : NOR2_X2 port map( A1 => n2202, A2 => n3683, ZN => n39441);
   U10233 : AOI21_X1 port map( A1 => n37423, A2 => n29679, B => n9610, ZN => 
                           n36168);
   U10234 : INV_X1 port map( I => n39268, ZN => n37539);
   U10237 : XOR2_X1 port map( A1 => n22754, A2 => n7358, Z => n9449);
   U10239 : NAND3_X2 port map( A1 => n37397, A2 => n25874, A3 => n6222, ZN => 
                           n25878);
   U10243 : NAND2_X2 port map( A1 => n32974, A2 => n36546, ZN => n37397);
   U10244 : OR3_X1 port map( A1 => n10436, A2 => n37815, A3 => n8452, Z => 
                           n4566);
   U10246 : NAND2_X2 port map( A1 => n38014, A2 => n27685, ZN => n9848);
   U10249 : OAI21_X2 port map( A1 => n19546, A2 => n35839, B => n37398, ZN => 
                           n21774);
   U10251 : XOR2_X1 port map( A1 => n37400, A2 => n1738, Z => Ciphertext(184));
   U10252 : NOR2_X1 port map( A1 => n15419, A2 => n39139, ZN => n37400);
   U10254 : OAI21_X2 port map( A1 => n37401, A2 => n15605, B => n30238, ZN => 
                           n5054);
   U10257 : INV_X2 port map( I => n29200, ZN => n37401);
   U10276 : NAND2_X2 port map( A1 => n892, A2 => n30154, ZN => n29200);
   U10284 : OAI22_X2 port map( A1 => n37178, A2 => n11945, B1 => n20884, B2 => 
                           n34117, ZN => n26157);
   U10285 : OAI21_X2 port map( A1 => n4317, A2 => n4318, B => n4316, ZN => 
                           n35727);
   U10287 : NAND2_X2 port map( A1 => n5527, A2 => n33015, ZN => n4317);
   U10288 : XOR2_X1 port map( A1 => n26466, A2 => n26465, Z => n10112);
   U10290 : XOR2_X1 port map( A1 => n26394, A2 => n37024, Z => n26465);
   U10291 : NOR2_X1 port map( A1 => n37584, A2 => n25560, ZN => n37663);
   U10294 : NAND2_X2 port map( A1 => n37402, A2 => n505, ZN => n37486);
   U10295 : NAND2_X2 port map( A1 => n12428, A2 => n29451, ZN => n37402);
   U10307 : OAI21_X2 port map( A1 => n38594, A2 => n24274, B => n7279, ZN => 
                           n37717);
   U10311 : AOI21_X2 port map( A1 => n1823, A2 => n20494, B => n38970, ZN => 
                           n35549);
   U10321 : XOR2_X1 port map( A1 => n334, A2 => n16610, Z => n26497);
   U10325 : OAI21_X2 port map( A1 => n37821, A2 => n39781, B => n13756, ZN => 
                           n16610);
   U10332 : XOR2_X1 port map( A1 => n5484, A2 => n38791, Z => n2391);
   U10335 : XOR2_X1 port map( A1 => n27864, A2 => n37403, Z => n27757);
   U10337 : INV_X2 port map( I => n27738, ZN => n37403);
   U10341 : OAI22_X2 port map( A1 => n18438, A2 => n12108, B1 => n4490, B2 => 
                           n18436, ZN => n27738);
   U10355 : AOI21_X2 port map( A1 => n37918, A2 => n37919, B => n37404, ZN => 
                           n22588);
   U10366 : OAI22_X2 port map( A1 => n37113, A2 => n18253, B1 => n17976, B2 => 
                           n1683, ZN => n37404);
   U10370 : XOR2_X1 port map( A1 => n32776, A2 => n20586, Z => n17344);
   U10371 : AOI22_X2 port map( A1 => n2156, A2 => n37200, B1 => n2154, B2 => 
                           n1349, ZN => n2153);
   U10372 : NAND2_X2 port map( A1 => n37487, A2 => n18562, ZN => n37603);
   U10374 : XOR2_X1 port map( A1 => n10525, A2 => n22452, Z => n5516);
   U10377 : NAND2_X2 port map( A1 => n4495, A2 => n4494, ZN => n10525);
   U10378 : OR2_X1 port map( A1 => n11164, A2 => n8743, Z => n37557);
   U10380 : NAND2_X2 port map( A1 => n6491, A2 => n6492, ZN => n6490);
   U10381 : OAI21_X1 port map( A1 => n29884, A2 => n17286, B => n37405, ZN => 
                           n17748);
   U10382 : NAND3_X2 port map( A1 => n29883, A2 => n15773, A3 => n6720, ZN => 
                           n37405);
   U10384 : XOR2_X1 port map( A1 => n37406, A2 => n10107, Z => n23083);
   U10385 : XOR2_X1 port map( A1 => n22446, A2 => n21206, Z => n37406);
   U10386 : XOR2_X1 port map( A1 => n23946, A2 => n23947, Z => n23948);
   U10387 : XOR2_X1 port map( A1 => n35376, A2 => n10526, Z => n23947);
   U10388 : XOR2_X1 port map( A1 => n29243, A2 => n28824, Z => n3707);
   U10389 : XOR2_X1 port map( A1 => n29042, A2 => n39739, Z => n29243);
   U10391 : OR2_X1 port map( A1 => n31272, A2 => n20070, Z => n39692);
   U10393 : XOR2_X1 port map( A1 => n22710, A2 => n1322, Z => n39215);
   U10402 : XOR2_X1 port map( A1 => n37407, A2 => n19800, Z => Ciphertext(87));
   U10414 : NAND3_X1 port map( A1 => n2111, A2 => n2110, A3 => n3118, ZN => 
                           n37407);
   U10416 : NAND2_X2 port map( A1 => n37408, A2 => n7717, ZN => n28433);
   U10417 : NAND2_X2 port map( A1 => n39419, A2 => n34863, ZN => n37408);
   U10427 : OAI21_X2 port map( A1 => n1564, A2 => n24816, B => n33012, ZN => 
                           n6408);
   U10428 : INV_X2 port map( I => n36191, ZN => n1633);
   U10431 : NAND2_X2 port map( A1 => n12698, A2 => n12697, ZN => n36191);
   U10434 : NAND2_X2 port map( A1 => n37409, A2 => n27176, ZN => n27499);
   U10494 : OAI22_X2 port map( A1 => n30732, A2 => n27174, B1 => n34562, B2 => 
                           n19132, ZN => n37409);
   U10498 : NAND2_X2 port map( A1 => n37892, A2 => n37410, ZN => n39423);
   U10503 : AOI21_X2 port map( A1 => n28015, A2 => n7326, B => n20164, ZN => 
                           n37410);
   U10506 : OAI21_X1 port map( A1 => n16590, A2 => n16366, B => n18920, ZN => 
                           n24100);
   U10508 : INV_X2 port map( I => n32898, ZN => n37411);
   U10509 : AND2_X1 port map( A1 => n37016, A2 => n37411, Z => n24644);
   U10511 : XOR2_X1 port map( A1 => n10941, A2 => n37412, Z => n10940);
   U10512 : XOR2_X1 port map( A1 => n33524, A2 => n23727, Z => n37412);
   U10517 : OAI21_X1 port map( A1 => n37414, A2 => n9586, B => n37413, ZN => 
                           n28063);
   U10520 : NAND2_X1 port map( A1 => n18722, A2 => n32820, ZN => n2155);
   U10523 : XOR2_X1 port map( A1 => Plaintext(61), A2 => Key(61), Z => n32820);
   U10524 : NOR2_X2 port map( A1 => n20267, A2 => n36620, ZN => n11476);
   U10525 : XOR2_X1 port map( A1 => n20341, A2 => n37243, Z => n38381);
   U10527 : XOR2_X1 port map( A1 => n37415, A2 => n17140, Z => n38111);
   U10528 : XOR2_X1 port map( A1 => n17850, A2 => n11525, Z => n37415);
   U10530 : NAND2_X2 port map( A1 => n11697, A2 => n18036, ZN => n3664);
   U10531 : NOR2_X2 port map( A1 => n15975, A2 => n3234, ZN => n11697);
   U10533 : XOR2_X1 port map( A1 => n33252, A2 => n26379, Z => n26521);
   U10534 : NAND2_X2 port map( A1 => n38131, A2 => n5161, ZN => n33252);
   U10535 : INV_X2 port map( I => n24469, ZN => n38303);
   U10536 : AND2_X1 port map( A1 => n24469, A2 => n38839, Z => n8916);
   U10538 : NOR2_X2 port map( A1 => n26089, A2 => n37416, ZN => n5164);
   U10539 : NOR2_X1 port map( A1 => n32424, A2 => n7577, ZN => n34996);
   U10541 : NAND2_X2 port map( A1 => n37417, A2 => n1076, ZN => n11279);
   U10545 : NAND2_X2 port map( A1 => n37419, A2 => n274, ZN => n37417);
   U10548 : NAND2_X2 port map( A1 => n36954, A2 => n28278, ZN => n37419);
   U10549 : XOR2_X1 port map( A1 => n26231, A2 => n37476, Z => n26311);
   U10551 : NAND2_X2 port map( A1 => n3332, A2 => n26188, ZN => n26231);
   U10553 : XOR2_X1 port map( A1 => n37420, A2 => n24931, Z => n32639);
   U10555 : XOR2_X1 port map( A1 => n2653, A2 => n29051, Z => n37420);
   U10556 : XOR2_X1 port map( A1 => n19156, A2 => n25292, Z => n36138);
   U10557 : INV_X1 port map( I => n38909, ZN => n34156);
   U10559 : OR2_X1 port map( A1 => n38909, A2 => n25345, Z => n18217);
   U10564 : BUF_X2 port map( I => n16048, Z => n35001);
   U10566 : BUF_X2 port map( I => n19593, Z => n37421);
   U10569 : XOR2_X1 port map( A1 => n37422, A2 => n38870, Z => n38259);
   U10576 : XOR2_X1 port map( A1 => n27725, A2 => n37242, Z => n37422);
   U10577 : XOR2_X1 port map( A1 => n26569, A2 => n39691, Z => n32844);
   U10583 : NAND2_X1 port map( A1 => n37493, A2 => n18478, ZN => n32574);
   U10585 : BUF_X4 port map( I => n20936, Z => n35537);
   U10586 : NAND2_X1 port map( A1 => n29674, A2 => n14522, ZN => n37423);
   U10588 : XOR2_X1 port map( A1 => n5789, A2 => n37424, Z => n3675);
   U10601 : XOR2_X1 port map( A1 => n8003, A2 => n11102, Z => n37424);
   U10604 : AOI21_X2 port map( A1 => n10735, A2 => n27307, B => n37425, ZN => 
                           n5750);
   U10607 : NOR2_X1 port map( A1 => n14041, A2 => n17166, ZN => n37425);
   U10610 : NAND2_X2 port map( A1 => n36222, A2 => n27306, ZN => n14041);
   U10620 : NAND2_X2 port map( A1 => n16129, A2 => n14420, ZN => n22277);
   U10623 : OR2_X1 port map( A1 => n309, A2 => n28771, Z => n35776);
   U10624 : XOR2_X1 port map( A1 => n23563, A2 => n37426, Z => n35300);
   U10627 : XOR2_X1 port map( A1 => n39239, A2 => n23562, Z => n37426);
   U10628 : XOR2_X1 port map( A1 => n35220, A2 => n10791, Z => n3589);
   U10629 : NAND2_X2 port map( A1 => n14874, A2 => n24754, ZN => n10791);
   U10634 : NOR2_X1 port map( A1 => n3169, A2 => n3170, ZN => n38757);
   U10637 : NAND2_X2 port map( A1 => n14082, A2 => n25674, ZN => n14083);
   U10638 : NOR2_X2 port map( A1 => n11596, A2 => n11594, ZN => n12141);
   U10640 : AOI21_X2 port map( A1 => n11597, A2 => n29317, B => n29263, ZN => 
                           n11596);
   U10644 : AND3_X1 port map( A1 => n12235, A2 => n18466, A3 => n19658, Z => 
                           n4785);
   U10645 : XOR2_X1 port map( A1 => n27549, A2 => n27679, Z => n27725);
   U10647 : NAND2_X2 port map( A1 => n16751, A2 => n15945, ZN => n25097);
   U10649 : NAND3_X2 port map( A1 => n16990, A2 => n38738, A3 => n38942, ZN => 
                           n16751);
   U10652 : XOR2_X1 port map( A1 => n19561, A2 => n27823, Z => n13035);
   U10653 : NAND2_X2 port map( A1 => n34989, A2 => n33016, ZN => n19561);
   U10655 : BUF_X2 port map( I => n18595, Z => n37428);
   U10656 : XOR2_X1 port map( A1 => n31240, A2 => n23937, Z => n34439);
   U10658 : XOR2_X1 port map( A1 => n39412, A2 => n23938, Z => n31240);
   U10660 : NAND2_X2 port map( A1 => n37429, A2 => n22032, ZN => n22348);
   U10661 : OAI21_X2 port map( A1 => n19012, A2 => n7916, B => n19011, ZN => 
                           n37429);
   U10662 : OAI21_X1 port map( A1 => n36548, A2 => n29627, B => n35405, ZN => 
                           n37430);
   U10665 : NAND2_X2 port map( A1 => n12543, A2 => n18960, ZN => n28652);
   U10672 : AOI21_X2 port map( A1 => n27115, A2 => n33088, B => n19334, ZN => 
                           n37433);
   U10674 : NOR2_X2 port map( A1 => n37435, A2 => n16132, ZN => n12396);
   U10675 : XOR2_X1 port map( A1 => n37874, A2 => n31515, Z => n21186);
   U10679 : AOI21_X2 port map( A1 => n13028, A2 => n28653, B => n13027, ZN => 
                           n37874);
   U10681 : NAND3_X2 port map( A1 => n38536, A2 => n38534, A3 => n38252, ZN => 
                           n21066);
   U10689 : XOR2_X1 port map( A1 => n31137, A2 => n18650, Z => n5566);
   U10691 : XOR2_X1 port map( A1 => n27687, A2 => n19606, Z => n18650);
   U10692 : XOR2_X1 port map( A1 => n22635, A2 => n37434, Z => n17430);
   U10693 : XOR2_X1 port map( A1 => n36641, A2 => n22620, Z => n37434);
   U10694 : AOI21_X2 port map( A1 => n2751, A2 => n5674, B => n34310, ZN => 
                           n37476);
   U10695 : OR2_X2 port map( A1 => n37104, A2 => n26988, Z => n26989);
   U10697 : OR2_X1 port map( A1 => n29885, A2 => n6720, Z => n29884);
   U10701 : OAI22_X2 port map( A1 => n32539, A2 => n35342, B1 => n17148, B2 => 
                           n19093, ZN => n6720);
   U10702 : NAND2_X2 port map( A1 => n30191, A2 => n30245, ZN => n35391);
   U10703 : INV_X2 port map( I => n883, ZN => n1070);
   U10704 : XNOR2_X1 port map( A1 => n4362, A2 => n4364, ZN => n883);
   U10708 : XOR2_X1 port map( A1 => n39100, A2 => n30648, Z => n33621);
   U10709 : AOI22_X2 port map( A1 => n33510, A2 => n14480, B1 => n17447, B2 => 
                           n28093, ZN => n28129);
   U10710 : OAI22_X2 port map( A1 => n18527, A2 => n14594, B1 => n20230, B2 => 
                           n33196, ZN => n37435);
   U10711 : NAND2_X2 port map( A1 => n38435, A2 => n34799, ZN => n12306);
   U10714 : XOR2_X1 port map( A1 => n37436, A2 => n37380, Z => Ciphertext(35));
   U10715 : NOR2_X1 port map( A1 => n15957, A2 => n15956, ZN => n37436);
   U10719 : XOR2_X1 port map( A1 => n17159, A2 => n12231, Z => n13724);
   U10720 : XOR2_X1 port map( A1 => n37437, A2 => n19681, Z => Ciphertext(14));
   U10721 : NAND2_X1 port map( A1 => n15027, A2 => n15026, ZN => n37437);
   U10723 : INV_X4 port map( I => n25611, ZN => n34010);
   U10724 : XOR2_X1 port map( A1 => n15078, A2 => n26260, Z => n15077);
   U10725 : INV_X2 port map( I => n26412, ZN => n15078);
   U10727 : XOR2_X1 port map( A1 => n26519, A2 => n26259, Z => n26412);
   U10729 : XOR2_X1 port map( A1 => n37438, A2 => n9315, Z => n37829);
   U10730 : XOR2_X1 port map( A1 => n27774, A2 => n13703, Z => n37438);
   U10737 : NOR2_X2 port map( A1 => n35434, A2 => n37439, ZN => n4184);
   U10738 : AOI21_X2 port map( A1 => n10013, A2 => n24847, B => n19630, ZN => 
                           n24730);
   U10740 : NAND2_X2 port map( A1 => n37168, A2 => n13625, ZN => n24847);
   U10749 : AOI21_X2 port map( A1 => n36590, A2 => n1408, B => n37440, ZN => 
                           n2013);
   U10757 : NOR3_X1 port map( A1 => n1962, A2 => n20866, A3 => n20673, ZN => 
                           n37440);
   U10758 : XOR2_X1 port map( A1 => n26379, A2 => n19902, Z => n26380);
   U10760 : NAND2_X2 port map( A1 => n21265, A2 => n34742, ZN => n26379);
   U10763 : XOR2_X1 port map( A1 => n9858, A2 => n17890, Z => n26376);
   U10764 : NAND2_X2 port map( A1 => n10016, A2 => n12941, ZN => n9858);
   U10766 : NAND2_X2 port map( A1 => n34217, A2 => n16250, ZN => n25990);
   U10771 : NAND2_X2 port map( A1 => n20337, A2 => n37441, ZN => n25951);
   U10772 : NAND2_X2 port map( A1 => n25564, A2 => n39458, ZN => n37441);
   U10773 : XOR2_X1 port map( A1 => n4624, A2 => n22488, Z => n22760);
   U10776 : NAND2_X2 port map( A1 => n3267, A2 => n3265, ZN => n4624);
   U10779 : XOR2_X1 port map( A1 => n37442, A2 => n8826, Z => n37587);
   U10783 : XOR2_X1 port map( A1 => n31773, A2 => n23801, Z => n37442);
   U10785 : NOR3_X1 port map( A1 => n27288, A2 => n34279, A3 => n39417, ZN => 
                           n36314);
   U10786 : NAND2_X2 port map( A1 => n4641, A2 => n36538, ZN => n39417);
   U10787 : NOR2_X2 port map( A1 => n35119, A2 => n35118, ZN => n15945);
   U10791 : OR2_X1 port map( A1 => n31760, A2 => n13872, Z => n39273);
   U10793 : XOR2_X1 port map( A1 => n36423, A2 => n38569, Z => n31760);
   U10795 : INV_X2 port map( I => n38880, ZN => n1612);
   U10797 : XOR2_X1 port map( A1 => n38880, A2 => n37443, Z => n23357);
   U10802 : NAND2_X2 port map( A1 => n39276, A2 => n2933, ZN => n38880);
   U10805 : NOR2_X2 port map( A1 => n12966, A2 => n7225, ZN => n39788);
   U10810 : NOR2_X2 port map( A1 => n23137, A2 => n23136, ZN => n12966);
   U10814 : OAI22_X2 port map( A1 => n7209, A2 => n17067, B1 => n20795, B2 => 
                           n7210, ZN => n35893);
   U10815 : NAND2_X1 port map( A1 => n14900, A2 => n2500, ZN => n14001);
   U10817 : AOI22_X2 port map( A1 => n31353, A2 => n15792, B1 => n28560, B2 => 
                           n28617, ZN => n2500);
   U10818 : OAI21_X2 port map( A1 => n37444, A2 => n36643, B => n31942, ZN => 
                           n18223);
   U10820 : NOR2_X2 port map( A1 => n13366, A2 => n36517, ZN => n37444);
   U10821 : NAND2_X1 port map( A1 => n8651, A2 => n19448, ZN => n16049);
   U10823 : XOR2_X1 port map( A1 => n10076, A2 => n26520, Z => n26258);
   U10824 : OAI21_X2 port map( A1 => n14579, A2 => n15177, B => n33764, ZN => 
                           n10076);
   U10830 : AND2_X1 port map( A1 => n37934, A2 => n37651, Z => n14645);
   U10831 : AOI21_X2 port map( A1 => n7239, A2 => n7237, B => n7234, ZN => 
                           n33263);
   U10832 : XOR2_X1 port map( A1 => n37446, A2 => n29282, Z => Ciphertext(21));
   U10837 : NAND3_X1 port map( A1 => n29280, A2 => n29281, A3 => n29279, ZN => 
                           n37446);
   U10839 : XOR2_X1 port map( A1 => n8402, A2 => n35986, Z => n27716);
   U10840 : XOR2_X1 port map( A1 => n37447, A2 => n1714, Z => Ciphertext(121));
   U10841 : AOI22_X1 port map( A1 => n29877, A2 => n29876, B1 => n29880, B2 => 
                           n29889, ZN => n37447);
   U10842 : INV_X4 port map( I => n1548, ZN => n33022);
   U10851 : NAND2_X1 port map( A1 => n1284, A2 => n17081, ZN => n38097);
   U10854 : XOR2_X1 port map( A1 => n35721, A2 => n37448, Z => n39611);
   U10856 : INV_X4 port map( I => n2678, ZN => n2534);
   U10859 : INV_X4 port map( I => n32802, ZN => n39258);
   U10860 : INV_X4 port map( I => n8131, ZN => n35357);
   U10862 : NAND2_X2 port map( A1 => n33059, A2 => n6588, ZN => n8131);
   U10864 : XOR2_X1 port map( A1 => n10329, A2 => n25180, Z => n10333);
   U10879 : XOR2_X1 port map( A1 => n1259, A2 => n11698, Z => n10329);
   U10880 : NAND2_X1 port map( A1 => n38906, A2 => n30799, ZN => n28184);
   U10881 : OR2_X1 port map( A1 => n10266, A2 => n19435, Z => n12349);
   U10889 : NAND2_X1 port map( A1 => n33646, A2 => n20879, ZN => n34285);
   U10890 : NOR2_X1 port map( A1 => n38568, A2 => n37903, ZN => n12776);
   U10891 : NAND2_X1 port map( A1 => n24273, A2 => n24272, ZN => n35959);
   U10895 : XOR2_X1 port map( A1 => n22748, A2 => n12901, Z => n12898);
   U10899 : XOR2_X1 port map( A1 => n22411, A2 => n22430, Z => n22748);
   U10900 : NAND2_X2 port map( A1 => n19476, A2 => n1755, ZN => n30720);
   U10901 : NAND2_X2 port map( A1 => n31312, A2 => n37449, ZN => n34533);
   U10904 : OR2_X1 port map( A1 => n26019, A2 => n26020, Z => n37449);
   U10905 : NAND3_X2 port map( A1 => n37450, A2 => n2130, A3 => n2129, ZN => 
                           n36496);
   U10906 : NAND2_X1 port map( A1 => n26624, A2 => n35764, ZN => n37450);
   U10910 : XOR2_X1 port map( A1 => n17908, A2 => n22486, Z => n19781);
   U10911 : XOR2_X1 port map( A1 => n22485, A2 => n22484, Z => n17908);
   U10912 : INV_X1 port map( I => n39769, ZN => n34070);
   U10913 : NAND2_X2 port map( A1 => n19544, A2 => n12081, ZN => n39769);
   U10914 : XOR2_X1 port map( A1 => n22392, A2 => n1660, Z => n38118);
   U10916 : NAND3_X2 port map( A1 => n37453, A2 => n38855, A3 => n37452, ZN => 
                           n37927);
   U10919 : NAND2_X1 port map( A1 => n5383, A2 => n12527, ZN => n37452);
   U10929 : NAND3_X2 port map( A1 => n32283, A2 => n34664, A3 => n2356, ZN => 
                           n16094);
   U10934 : NAND2_X2 port map( A1 => n14052, A2 => n8499, ZN => n35981);
   U10935 : AOI22_X2 port map( A1 => n38047, A2 => n20981, B1 => n27286, B2 => 
                           n10284, ZN => n27501);
   U10938 : NAND2_X2 port map( A1 => n465, A2 => n8758, ZN => n15423);
   U10939 : OAI22_X2 port map( A1 => n10487, A2 => n22344, B1 => n22170, B2 => 
                           n22342, ZN => n347);
   U10941 : NAND2_X2 port map( A1 => n37455, A2 => n26835, ZN => n8105);
   U10942 : NAND2_X2 port map( A1 => n26722, A2 => n9269, ZN => n37455);
   U10945 : INV_X1 port map( I => n2437, ZN => n38076);
   U10948 : NOR2_X1 port map( A1 => n34430, A2 => n24394, ZN => n21319);
   U10949 : XOR2_X1 port map( A1 => n19536, A2 => n23861, Z => n23688);
   U10951 : AOI21_X2 port map( A1 => n23447, A2 => n2084, B => n10078, ZN => 
                           n23861);
   U10952 : NAND3_X1 port map( A1 => n30230, A2 => n30228, A3 => n30229, ZN => 
                           n37636);
   U10953 : NAND2_X2 port map( A1 => n36243, A2 => n35535, ZN => n19203);
   U10956 : XOR2_X1 port map( A1 => n37456, A2 => n9994, Z => n4786);
   U10957 : XOR2_X1 port map( A1 => n13176, A2 => n11479, Z => n37456);
   U10959 : NAND2_X2 port map( A1 => n24138, A2 => n24139, ZN => n39279);
   U10960 : OR2_X1 port map( A1 => n24639, A2 => n24250, Z => n20800);
   U10962 : NOR2_X1 port map( A1 => n9758, A2 => n30445, ZN => n14916);
   U10965 : OAI22_X2 port map( A1 => n2769, A2 => n2768, B1 => n2767, B2 => 
                           n36225, ZN => n16180);
   U10969 : XOR2_X1 port map( A1 => n38989, A2 => n21154, Z => n233);
   U10978 : OAI22_X2 port map( A1 => n36624, A2 => n4636, B1 => n4132, B2 => 
                           n17353, ZN => n17624);
   U10981 : INV_X4 port map( I => n2747, ZN => n38794);
   U10983 : XOR2_X1 port map( A1 => n20501, A2 => n37457, Z => n14000);
   U10984 : XOR2_X1 port map( A1 => n10153, A2 => n31999, Z => n37457);
   U10986 : NOR2_X2 port map( A1 => n21627, A2 => n10085, ZN => n7357);
   U10987 : XOR2_X1 port map( A1 => n18051, A2 => n8833, Z => n4077);
   U10991 : NOR2_X2 port map( A1 => n38672, A2 => n31831, ZN => n8833);
   U10993 : AOI21_X1 port map( A1 => n5424, A2 => n3538, B => n17583, ZN => 
                           n39555);
   U10994 : NAND3_X2 port map( A1 => n32374, A2 => n3461, A3 => n28075, ZN => 
                           n17583);
   U10995 : INV_X2 port map( I => n16180, ZN => n30111);
   U10996 : XOR2_X1 port map( A1 => n23885, A2 => n24025, Z => n23743);
   U11002 : AOI21_X2 port map( A1 => n22873, A2 => n16047, B => n37458, ZN => 
                           n23623);
   U11004 : OAI22_X2 port map( A1 => n22872, A2 => n16047, B1 => n20776, B2 => 
                           n961, ZN => n37458);
   U11007 : INV_X2 port map( I => n37459, ZN => n23162);
   U11008 : XOR2_X1 port map( A1 => n37461, A2 => n10396, Z => n13862);
   U11010 : XOR2_X1 port map( A1 => n15164, A2 => n36656, Z => n37461);
   U11014 : XOR2_X1 port map( A1 => n27580, A2 => n29805, Z => n10399);
   U11016 : NAND2_X2 port map( A1 => n37978, A2 => n33160, ZN => n27580);
   U11019 : NAND2_X2 port map( A1 => n31362, A2 => n692, ZN => n25954);
   U11027 : NOR3_X1 port map( A1 => n39048, A2 => n31133, A3 => n25820, ZN => 
                           n25821);
   U11029 : NOR2_X2 port map( A1 => n37464, A2 => n36682, ZN => n7291);
   U11030 : NOR2_X1 port map( A1 => n2967, A2 => n2968, ZN => n37464);
   U11036 : XNOR2_X1 port map( A1 => n15368, A2 => n6026, ZN => n39259);
   U11037 : NAND2_X1 port map( A1 => n9415, A2 => n27428, ZN => n17718);
   U11038 : INV_X2 port map( I => n35427, ZN => n27428);
   U11042 : NAND2_X2 port map( A1 => n37766, A2 => n39508, ZN => n35427);
   U11051 : NAND2_X2 port map( A1 => n37734, A2 => n30220, ZN => n29202);
   U11053 : OAI21_X2 port map( A1 => n37250, A2 => n37465, B => n27228, ZN => 
                           n27592);
   U11054 : OR2_X1 port map( A1 => n29208, A2 => n15535, Z => n29207);
   U11055 : XNOR2_X1 port map( A1 => n38192, A2 => n7247, ZN => n9960);
   U11056 : NAND2_X2 port map( A1 => n7243, A2 => n7241, ZN => n7247);
   U11059 : INV_X2 port map( I => n38848, ZN => n34720);
   U11061 : NAND2_X2 port map( A1 => n37975, A2 => n37472, ZN => n38848);
   U11062 : XOR2_X1 port map( A1 => n25206, A2 => n25208, Z => n6658);
   U11063 : BUF_X2 port map( I => n34345, Z => n37466);
   U11068 : NAND2_X2 port map( A1 => n39533, A2 => n38373, ZN => n23982);
   U11071 : OR2_X2 port map( A1 => n39639, A2 => n20361, Z => n21854);
   U11080 : NAND2_X1 port map( A1 => n15376, A2 => n19599, ZN => n39740);
   U11083 : INV_X2 port map( I => n9387, ZN => n8792);
   U11084 : NAND2_X2 port map( A1 => n7998, A2 => n7999, ZN => n9387);
   U11086 : NAND2_X1 port map( A1 => n10019, A2 => n37999, ZN => n24689);
   U11087 : NAND2_X2 port map( A1 => n37468, A2 => n37467, ZN => n24412);
   U11090 : INV_X1 port map( I => n31403, ZN => n37467);
   U11093 : INV_X2 port map( I => n24408, ZN => n37468);
   U11097 : XOR2_X1 port map( A1 => n19600, A2 => n7032, Z => n7031);
   U11098 : NAND2_X2 port map( A1 => n37114, A2 => n37469, ZN => n6068);
   U11108 : NOR2_X2 port map( A1 => n4369, A2 => n37470, ZN => n37469);
   U11111 : NOR2_X2 port map( A1 => n28639, A2 => n39355, ZN => n37470);
   U11112 : NOR2_X2 port map( A1 => n37471, A2 => n8963, ZN => n4584);
   U11116 : NOR2_X2 port map( A1 => n1495, A2 => n8311, ZN => n37471);
   U11125 : NAND2_X2 port map( A1 => n9218, A2 => n20326, ZN => n20605);
   U11127 : XOR2_X1 port map( A1 => n25164, A2 => n8240, Z => n31151);
   U11132 : XOR2_X1 port map( A1 => n13076, A2 => n15625, Z => n25164);
   U11133 : XOR2_X1 port map( A1 => n29140, A2 => n29139, Z => n5347);
   U11138 : OAI22_X1 port map( A1 => n30080, A2 => n30070, B1 => n6453, B2 => 
                           n30066, ZN => n30730);
   U11143 : NOR2_X2 port map( A1 => n4168, A2 => n4379, ZN => n30080);
   U11145 : NAND2_X2 port map( A1 => n39194, A2 => n9862, ZN => n23441);
   U11148 : NAND2_X2 port map( A1 => n3047, A2 => n3046, ZN => n39194);
   U11152 : NAND2_X1 port map( A1 => n36669, A2 => n13610, ZN => n39735);
   U11157 : AOI21_X1 port map( A1 => n7797, A2 => n37473, B => n7792, ZN => 
                           n32903);
   U11159 : NAND2_X1 port map( A1 => n7795, A2 => n7796, ZN => n37473);
   U11160 : AND2_X1 port map( A1 => n18164, A2 => n32622, Z => n11646);
   U11161 : XOR2_X1 port map( A1 => n4341, A2 => n29289, Z => n17957);
   U11163 : NAND2_X2 port map( A1 => n6093, A2 => n12342, ZN => n4341);
   U11166 : NAND2_X1 port map( A1 => n38595, A2 => n38115, ZN => n38594);
   U11174 : NOR2_X2 port map( A1 => n39513, A2 => n37475, ZN => n37474);
   U11182 : INV_X2 port map( I => n38674, ZN => n37475);
   U11183 : BUF_X4 port map( I => n3455, Z => n38437);
   U11184 : NOR2_X2 port map( A1 => n4155, A2 => n19750, ZN => n4927);
   U11187 : NAND2_X2 port map( A1 => n11890, A2 => n10254, ZN => n4155);
   U11188 : NAND2_X2 port map( A1 => n6913, A2 => n6912, ZN => n39196);
   U11192 : INV_X4 port map( I => n19465, ZN => n37604);
   U11199 : XOR2_X1 port map( A1 => n6535, A2 => n6537, Z => n11428);
   U11201 : AOI21_X1 port map( A1 => n37819, A2 => n37613, B => n19740, ZN => 
                           n12526);
   U11202 : OAI21_X2 port map( A1 => n20628, A2 => n20626, B => n14486, ZN => 
                           n37613);
   U11209 : NOR2_X1 port map( A1 => n9547, A2 => n626, ZN => n6483);
   U11210 : INV_X2 port map( I => n32518, ZN => n626);
   U11211 : XOR2_X1 port map( A1 => n6988, A2 => n6985, Z => n32518);
   U11214 : NAND2_X1 port map( A1 => n6645, A2 => n37478, ZN => n3723);
   U11220 : NAND2_X2 port map( A1 => n6646, A2 => n38725, ZN => n37478);
   U11224 : XOR2_X1 port map( A1 => n25089, A2 => n37479, Z => n36537);
   U11226 : XOR2_X1 port map( A1 => n39320, A2 => n15912, Z => n37479);
   U11227 : XOR2_X1 port map( A1 => n1555, A2 => n25241, Z => n25089);
   U11232 : XOR2_X1 port map( A1 => n38710, A2 => n29817, Z => n29936);
   U11233 : XOR2_X1 port map( A1 => n29043, A2 => n31782, Z => n29817);
   U11234 : XOR2_X1 port map( A1 => n23776, A2 => n23829, Z => n24058);
   U11236 : NAND3_X2 port map( A1 => n23239, A2 => n23241, A3 => n23240, ZN => 
                           n23776);
   U11237 : NAND2_X2 port map( A1 => n9823, A2 => n23238, ZN => n23460);
   U11239 : NAND2_X2 port map( A1 => n35347, A2 => n14875, ZN => n9823);
   U11240 : NAND2_X2 port map( A1 => n30775, A2 => n23873, ZN => n6583);
   U11242 : NAND2_X2 port map( A1 => n35278, A2 => n35279, ZN => n30775);
   U11247 : NAND2_X2 port map( A1 => n11852, A2 => n4058, ZN => n21925);
   U11249 : XOR2_X1 port map( A1 => n11099, A2 => n32127, Z => n36253);
   U11251 : XOR2_X1 port map( A1 => n18498, A2 => n39614, Z => n11099);
   U11253 : XOR2_X1 port map( A1 => n1895, A2 => n11950, Z => n1897);
   U11254 : NAND2_X2 port map( A1 => n198, A2 => n199, ZN => n1895);
   U11255 : NOR2_X2 port map( A1 => n37482, A2 => n37481, ZN => n7144);
   U11258 : NOR2_X2 port map( A1 => n23229, A2 => n23749, ZN => n37481);
   U11261 : XOR2_X1 port map( A1 => n22601, A2 => n37466, Z => n13652);
   U11263 : AOI21_X2 port map( A1 => n5557, A2 => n8518, B => n5556, ZN => 
                           n34345);
   U11266 : NAND2_X1 port map( A1 => n39638, A2 => n14170, ZN => n26860);
   U11269 : XOR2_X1 port map( A1 => n39612, A2 => n39611, Z => n39638);
   U11270 : INV_X2 port map( I => n37483, ZN => n10642);
   U11273 : XNOR2_X1 port map( A1 => n11099, A2 => n32127, ZN => n37483);
   U11274 : NAND2_X2 port map( A1 => n37485, A2 => n37506, ZN => n9859);
   U11275 : AND2_X1 port map( A1 => n14840, A2 => n25369, Z => n37485);
   U11279 : NAND2_X2 port map( A1 => n37486, A2 => n2132, ZN => n29473);
   U11281 : INV_X2 port map( I => n36177, ZN => n27372);
   U11283 : NAND2_X2 port map( A1 => n33853, A2 => n3255, ZN => n36177);
   U11285 : NAND3_X1 port map( A1 => n24788, A2 => n8430, A3 => n18148, ZN => 
                           n18564);
   U11287 : XOR2_X1 port map( A1 => n6403, A2 => n33231, Z => n6402);
   U11288 : NOR3_X2 port map( A1 => n3644, A2 => n38448, A3 => n1049, ZN => 
                           n10743);
   U11289 : INV_X4 port map( I => n2654, ZN => n3644);
   U11290 : NOR2_X2 port map( A1 => n34059, A2 => n35860, ZN => n2654);
   U11291 : NAND2_X2 port map( A1 => n32614, A2 => n38967, ZN => n18850);
   U11292 : XOR2_X1 port map( A1 => n5116, A2 => n24076, Z => n10683);
   U11295 : NAND2_X1 port map( A1 => n11196, A2 => n24447, ZN => n38312);
   U11297 : NAND3_X2 port map( A1 => n35753, A2 => n10842, A3 => n10841, ZN => 
                           n12362);
   U11300 : XOR2_X1 port map( A1 => n37489, A2 => n15311, Z => n10860);
   U11302 : XOR2_X1 port map( A1 => n13236, A2 => n10862, Z => n37489);
   U11303 : AOI22_X2 port map( A1 => n30862, A2 => n24723, B1 => n32398, B2 => 
                           n4323, ZN => n18600);
   U11304 : OAI22_X2 port map( A1 => n24723, A2 => n24717, B1 => n5056, B2 => 
                           n24719, ZN => n4323);
   U11308 : NAND2_X2 port map( A1 => n34317, A2 => n37490, ZN => n16226);
   U11309 : OAI21_X2 port map( A1 => n22235, A2 => n19261, B => n18064, ZN => 
                           n37491);
   U11310 : XOR2_X1 port map( A1 => n37492, A2 => n29157, Z => n8443);
   U11317 : XOR2_X1 port map( A1 => n16334, A2 => n5041, Z => n37492);
   U11320 : OAI22_X2 port map( A1 => n38357, A2 => n39800, B1 => n25379, B2 => 
                           n19863, ZN => n38356);
   U11325 : XOR2_X1 port map( A1 => n23685, A2 => n19953, Z => n4327);
   U11327 : NAND3_X2 port map( A1 => n4287, A2 => n4290, A3 => n4288, ZN => 
                           n23685);
   U11336 : XOR2_X1 port map( A1 => n26324, A2 => n26247, Z => n2069);
   U11345 : XOR2_X1 port map( A1 => n26554, A2 => n7402, Z => n26247);
   U11346 : NAND2_X2 port map( A1 => n23333, A2 => n17167, ZN => n37493);
   U11347 : AND2_X1 port map( A1 => n36685, A2 => n28591, Z => n4833);
   U11352 : NAND3_X2 port map( A1 => n17, A2 => n28162, A3 => n11742, ZN => 
                           n36685);
   U11355 : XOR2_X1 port map( A1 => n17462, A2 => n23675, Z => n24019);
   U11356 : NAND2_X2 port map( A1 => n10570, A2 => n23118, ZN => n17462);
   U11358 : NAND2_X2 port map( A1 => n23094, A2 => n6466, ZN => n7026);
   U11362 : NOR2_X2 port map( A1 => n9586, A2 => n28430, ZN => n39190);
   U11364 : INV_X2 port map( I => n32472, ZN => n585);
   U11365 : XOR2_X1 port map( A1 => n38781, A2 => n37494, Z => n38597);
   U11366 : XOR2_X1 port map( A1 => n742, A2 => n37223, Z => n37494);
   U11368 : AOI21_X2 port map( A1 => n1521, A2 => n930, B => n7258, ZN => 
                           n36568);
   U11374 : XOR2_X1 port map( A1 => n10926, A2 => n10928, Z => n20838);
   U11377 : NAND2_X1 port map( A1 => n18694, A2 => n38477, ZN => n38476);
   U11380 : XOR2_X1 port map( A1 => n2896, A2 => n24552, Z => n33946);
   U11381 : NAND2_X2 port map( A1 => n4159, A2 => n31080, ZN => n16182);
   U11382 : INV_X1 port map( I => n29856, ZN => n37497);
   U11384 : NAND2_X2 port map( A1 => n23390, A2 => n16013, ZN => n23453);
   U11389 : XOR2_X1 port map( A1 => n37495, A2 => n18751, Z => n22781);
   U11393 : XOR2_X1 port map( A1 => n33862, A2 => n22776, Z => n37495);
   U11395 : XOR2_X1 port map( A1 => n10370, A2 => n10722, Z => n10371);
   U11403 : AOI21_X2 port map( A1 => n12638, A2 => n12639, B => n36241, ZN => 
                           n10370);
   U11408 : INV_X2 port map( I => n13379, ZN => n3988);
   U11410 : OAI21_X2 port map( A1 => n36914, A2 => n34470, B => n27982, ZN => 
                           n13379);
   U11415 : NOR3_X1 port map( A1 => n22925, A2 => n6327, A3 => n38229, ZN => 
                           n32753);
   U11416 : XOR2_X1 port map( A1 => n17159, A2 => n17493, Z => n9923);
   U11420 : XOR2_X1 port map( A1 => n1065, A2 => n15581, Z => n17493);
   U11423 : XOR2_X1 port map( A1 => n36916, A2 => n10132, Z => n28262);
   U11427 : OAI21_X2 port map( A1 => n33706, A2 => n23084, B => n37496, ZN => 
                           n3713);
   U11431 : AOI22_X2 port map( A1 => n23184, A2 => n14396, B1 => n14725, B2 => 
                           n35567, ZN => n37496);
   U11434 : AOI22_X1 port map( A1 => n37497, A2 => n1054, B1 => n5579, B2 => 
                           n29858, ZN => n19872);
   U11438 : NAND2_X2 port map( A1 => n2347, A2 => n3861, ZN => n29856);
   U11442 : NAND2_X2 port map( A1 => n39538, A2 => n31937, ZN => n36058);
   U11443 : NAND2_X2 port map( A1 => n6921, A2 => n6920, ZN => n30033);
   U11445 : XOR2_X1 port map( A1 => n23590, A2 => n39209, Z => n17775);
   U11446 : NAND2_X2 port map( A1 => n38025, A2 => n38024, ZN => n39209);
   U11449 : XOR2_X1 port map( A1 => n27837, A2 => n27719, Z => n18048);
   U11450 : XOR2_X1 port map( A1 => n1468, A2 => n35229, Z => n27719);
   U11452 : NAND2_X1 port map( A1 => n21039, A2 => n17400, ZN => n25958);
   U11457 : NAND3_X1 port map( A1 => n35333, A2 => n5908, A3 => n26039, ZN => 
                           n36766);
   U11460 : NAND2_X2 port map( A1 => n25464, A2 => n34877, ZN => n35333);
   U11462 : AOI22_X2 port map( A1 => n17191, A2 => n28755, B1 => n32791, B2 => 
                           n16691, ZN => n14971);
   U11467 : AOI22_X2 port map( A1 => n34465, A2 => n34464, B1 => n1546, B2 => 
                           n25501, ZN => n25288);
   U11469 : OAI22_X2 port map( A1 => n6592, A2 => n37025, B1 => n14081, B2 => 
                           n25434, ZN => n25501);
   U11474 : NAND3_X2 port map( A1 => n2682, A2 => n2683, A3 => n23386, ZN => 
                           n2685);
   U11475 : XOR2_X1 port map( A1 => n6984, A2 => n25, Z => n34397);
   U11478 : XOR2_X1 port map( A1 => n27698, A2 => n27667, Z => n27001);
   U11483 : XOR2_X1 port map( A1 => n19396, A2 => n9315, Z => n27698);
   U11484 : INV_X2 port map( I => n28089, ZN => n8207);
   U11485 : NOR3_X1 port map( A1 => n36796, A2 => n11614, A3 => n8743, ZN => 
                           n27653);
   U11486 : INV_X4 port map( I => n3669, ZN => n17501);
   U11488 : NAND2_X2 port map( A1 => n35710, A2 => n39486, ZN => n3669);
   U11490 : NAND2_X2 port map( A1 => n37643, A2 => n19615, ZN => n26824);
   U11494 : INV_X2 port map( I => n37501, ZN => n12663);
   U11495 : XNOR2_X1 port map( A1 => n11235, A2 => n11237, ZN => n37501);
   U11496 : INV_X2 port map( I => n26328, ZN => n1515);
   U11498 : NAND2_X2 port map( A1 => n11533, A2 => n33258, ZN => n26328);
   U11500 : NAND2_X1 port map( A1 => n15290, A2 => n23173, ZN => n6645);
   U11504 : NAND2_X2 port map( A1 => n36911, A2 => n5101, ZN => n8260);
   U11510 : INV_X2 port map( I => n28389, ZN => n34702);
   U11511 : NOR2_X1 port map( A1 => n28081, A2 => n28080, ZN => n28082);
   U11512 : NAND2_X2 port map( A1 => n37503, A2 => n3904, ZN => n39020);
   U11513 : NAND3_X2 port map( A1 => n37960, A2 => n15334, A3 => n39235, ZN => 
                           n37503);
   U11515 : NAND2_X2 port map( A1 => n37504, A2 => n24481, ZN => n19713);
   U11518 : XOR2_X1 port map( A1 => n4436, A2 => n37505, Z => n39427);
   U11519 : XOR2_X1 port map( A1 => n22600, A2 => n3528, Z => n37505);
   U11521 : XOR2_X1 port map( A1 => n1616, A2 => n38468, Z => n6468);
   U11522 : NOR2_X2 port map( A1 => n38794, A2 => n934, ZN => n15527);
   U11525 : NAND2_X1 port map( A1 => n25368, A2 => n17855, ZN => n37506);
   U11526 : NAND3_X2 port map( A1 => n36918, A2 => n37507, A3 => n34881, ZN => 
                           n33038);
   U11530 : NAND2_X1 port map( A1 => n18325, A2 => n18326, ZN => n37507);
   U11537 : NAND2_X1 port map( A1 => n29380, A2 => n13302, ZN => n13942);
   U11538 : BUF_X2 port map( I => n27395, Z => n37508);
   U11539 : INV_X2 port map( I => n8899, ZN => n22300);
   U11541 : NAND2_X2 port map( A1 => n21, A2 => n4391, ZN => n8899);
   U11542 : NOR2_X2 port map( A1 => n35560, A2 => n32045, ZN => n24612);
   U11547 : NAND2_X2 port map( A1 => n37509, A2 => n34811, ZN => n2305);
   U11549 : NAND2_X2 port map( A1 => n9202, A2 => n1890, ZN => n37509);
   U11552 : XOR2_X1 port map( A1 => n23714, A2 => n2145, Z => n23725);
   U11553 : NOR2_X2 port map( A1 => n33775, A2 => n2086, ZN => n2145);
   U11554 : NAND2_X2 port map( A1 => n39668, A2 => n9941, ZN => n22298);
   U11556 : AOI21_X2 port map( A1 => n28399, A2 => n28755, B => n37510, ZN => 
                           n28610);
   U11558 : AOI21_X2 port map( A1 => n12312, A2 => n12313, B => n28755, ZN => 
                           n37510);
   U11559 : NAND3_X2 port map( A1 => n35963, A2 => n23444, A3 => n4207, ZN => 
                           n2087);
   U11561 : XOR2_X1 port map( A1 => n29306, A2 => n28948, Z => n29257);
   U11562 : OAI21_X2 port map( A1 => n27958, A2 => n28490, B => n27957, ZN => 
                           n29306);
   U11567 : XOR2_X1 port map( A1 => n33645, A2 => n26487, Z => n26370);
   U11569 : NAND2_X2 port map( A1 => n39633, A2 => n39822, ZN => n26487);
   U11570 : XOR2_X1 port map( A1 => n23952, A2 => n23775, Z => n23904);
   U11572 : AOI21_X2 port map( A1 => n6052, A2 => n23394, B => n23393, ZN => 
                           n23952);
   U11573 : XOR2_X1 port map( A1 => n37511, A2 => n10478, Z => n14463);
   U11575 : XOR2_X1 port map( A1 => n10887, A2 => n10888, Z => n37511);
   U11581 : AND2_X1 port map( A1 => n15359, A2 => n7696, Z => n17948);
   U11585 : XOR2_X1 port map( A1 => n38054, A2 => n18923, Z => n34120);
   U11589 : NOR2_X2 port map( A1 => n12663, A2 => n16500, ZN => n39127);
   U11590 : INV_X2 port map( I => n16489, ZN => n26639);
   U11591 : XOR2_X1 port map( A1 => n3995, A2 => n35017, Z => n16489);
   U11592 : NAND2_X2 port map( A1 => n26109, A2 => n13712, ZN => n16860);
   U11595 : XOR2_X1 port map( A1 => n26495, A2 => n11935, Z => n4205);
   U11598 : NAND2_X2 port map( A1 => n38249, A2 => n1647, ZN => n3813);
   U11599 : XNOR2_X1 port map( A1 => n25026, A2 => n18600, ZN => n25166);
   U11600 : XOR2_X1 port map( A1 => n37513, A2 => n4238, Z => n3229);
   U11602 : INV_X1 port map( I => n17837, ZN => n37513);
   U11603 : XOR2_X1 port map( A1 => n1261, A2 => n15102, Z => n17837);
   U11605 : NAND2_X1 port map( A1 => n1094, A2 => n37054, ZN => n26858);
   U11606 : INV_X1 port map( I => n25198, ZN => n37658);
   U11609 : NOR2_X2 port map( A1 => n37135, A2 => n37514, ZN => n38397);
   U11611 : NAND2_X2 port map( A1 => n6466, A2 => n31183, ZN => n22836);
   U11613 : OAI22_X2 port map( A1 => n39317, A2 => n37515, B1 => n24547, B2 => 
                           n37067, ZN => n19691);
   U11614 : NOR2_X2 port map( A1 => n37717, A2 => n11494, ZN => n32091);
   U11615 : NAND2_X1 port map( A1 => n33289, A2 => n12950, ZN => n24205);
   U11617 : NOR2_X2 port map( A1 => n37518, A2 => n37517, ZN => n37516);
   U11619 : NAND3_X2 port map( A1 => n37519, A2 => n19111, A3 => n31583, ZN => 
                           n19109);
   U11625 : NAND2_X2 port map( A1 => n38580, A2 => n32720, ZN => n37519);
   U11626 : XOR2_X1 port map( A1 => n17566, A2 => n22449, Z => n17565);
   U11634 : XOR2_X1 port map( A1 => n33736, A2 => n22743, Z => n22449);
   U11635 : OAI21_X1 port map( A1 => n31598, A2 => n967, B => n10848, ZN => 
                           n10847);
   U11640 : XOR2_X1 port map( A1 => n15912, A2 => n25182, Z => n19072);
   U11641 : NAND2_X2 port map( A1 => n18458, A2 => n24652, ZN => n15912);
   U11642 : CLKBUF_X4 port map( I => n17114, Z => n37661);
   U11645 : OAI22_X2 port map( A1 => n25927, A2 => n2029, B1 => n25928, B2 => 
                           n2561, ZN => n26084);
   U11646 : AOI22_X2 port map( A1 => n30059, A2 => n30000, B1 => n16353, B2 => 
                           n30057, ZN => n32548);
   U11649 : XOR2_X1 port map( A1 => n37520, A2 => n710, Z => n10181);
   U11653 : XOR2_X1 port map( A1 => n23671, A2 => n37521, Z => n37520);
   U11659 : INV_X2 port map( I => n7148, ZN => n37521);
   U11660 : XOR2_X1 port map( A1 => n37874, A2 => n296, Z => n29043);
   U11666 : OAI21_X2 port map( A1 => n28177, A2 => n38311, B => n35961, ZN => 
                           n296);
   U11670 : XOR2_X1 port map( A1 => n4077, A2 => n7101, Z => n7100);
   U11671 : NOR2_X1 port map( A1 => n8599, A2 => n8600, ZN => n8598);
   U11675 : NAND2_X2 port map( A1 => n37522, A2 => n37140, ZN => n14496);
   U11677 : NAND2_X2 port map( A1 => n37604, A2 => n37524, ZN => n10901);
   U11678 : INV_X1 port map( I => n26885, ZN => n37524);
   U11679 : BUF_X2 port map( I => n20128, Z => n37525);
   U11680 : AND2_X1 port map( A1 => n23060, A2 => n37922, Z => n39004);
   U11681 : XOR2_X1 port map( A1 => n11752, A2 => n6523, Z => n8502);
   U11683 : OAI21_X2 port map( A1 => n2421, A2 => n4854, B => n8161, ZN => 
                           n6523);
   U11684 : XOR2_X1 port map( A1 => n37526, A2 => n39245, Z => n34587);
   U11685 : XOR2_X1 port map( A1 => n11502, A2 => n27790, Z => n37526);
   U11687 : XOR2_X1 port map( A1 => n37527, A2 => n29168, Z => n33716);
   U11688 : XOR2_X1 port map( A1 => n32073, A2 => n29167, Z => n37527);
   U11689 : AND2_X1 port map( A1 => n19326, A2 => n27131, Z => n8486);
   U11692 : NAND2_X2 port map( A1 => n14216, A2 => n13607, ZN => n17287);
   U11694 : XOR2_X1 port map( A1 => n37529, A2 => n29206, Z => Ciphertext(4));
   U11698 : NAND2_X1 port map( A1 => n2569, A2 => n36862, ZN => n37529);
   U11704 : INV_X4 port map( I => n28400, ZN => n12537);
   U11705 : NOR2_X1 port map( A1 => n974, A2 => n28400, ZN => n36465);
   U11708 : XOR2_X1 port map( A1 => n37530, A2 => n23943, Z => n15860);
   U11711 : XOR2_X1 port map( A1 => n39408, A2 => n36461, Z => n37530);
   U11712 : XOR2_X1 port map( A1 => n33473, A2 => n37532, Z => n9214);
   U11713 : XOR2_X1 port map( A1 => n26522, A2 => n26344, Z => n37532);
   U11714 : XOR2_X1 port map( A1 => n37533, A2 => n36040, Z => Ciphertext(51));
   U11719 : AOI22_X1 port map( A1 => n6340, A2 => n6343, B1 => n6339, B2 => 
                           n13433, ZN => n37533);
   U11721 : XOR2_X1 port map( A1 => n10214, A2 => n10939, Z => n36002);
   U11725 : NOR2_X2 port map( A1 => n37534, A2 => n12239, ZN => n39588);
   U11726 : NOR3_X2 port map( A1 => n1146, A2 => n8569, A3 => n9699, ZN => 
                           n37534);
   U11729 : OAI22_X2 port map( A1 => n1337, A2 => n2709, B1 => n22022, B2 => 
                           n32434, ZN => n39455);
   U11733 : INV_X2 port map( I => n22086, ZN => n1337);
   U11734 : OAI21_X2 port map( A1 => n21491, A2 => n3670, B => n38091, ZN => 
                           n22086);
   U11735 : XOR2_X1 port map( A1 => n31568, A2 => n37038, Z => n15978);
   U11736 : NOR2_X2 port map( A1 => n15525, A2 => n15526, ZN => n37038);
   U11737 : NAND4_X1 port map( A1 => n29472, A2 => n29473, A3 => n29469, A4 => 
                           n29470, ZN => n6342);
   U11744 : XOR2_X1 port map( A1 => n10794, A2 => n29833, Z => n32200);
   U11746 : AOI22_X2 port map( A1 => n7869, A2 => n28539, B1 => n4228, B2 => 
                           n28538, ZN => n10794);
   U11753 : NAND2_X2 port map( A1 => n5304, A2 => n5303, ZN => n38976);
   U11754 : AOI22_X2 port map( A1 => n5551, A2 => n5132, B1 => n21916, B2 => 
                           n5391, ZN => n5304);
   U11759 : XOR2_X1 port map( A1 => n26569, A2 => n26466, Z => n26313);
   U11761 : XOR2_X1 port map( A1 => n26421, A2 => n20600, Z => n26466);
   U11764 : NAND2_X2 port map( A1 => n17826, A2 => n32797, ZN => n38466);
   U11766 : NOR2_X2 port map( A1 => n37535, A2 => n9233, ZN => n36889);
   U11768 : AOI21_X2 port map( A1 => n29993, A2 => n4095, B => n3693, ZN => 
                           n37535);
   U11771 : OAI22_X2 port map( A1 => n37536, A2 => n3363, B1 => n23525, B2 => 
                           n36103, ZN => n18540);
   U11775 : NAND2_X2 port map( A1 => n3366, A2 => n30835, ZN => n37536);
   U11776 : OAI21_X2 port map( A1 => n37538, A2 => n31845, B => n37537, ZN => 
                           n23859);
   U11777 : NOR2_X2 port map( A1 => n957, A2 => n38777, ZN => n37538);
   U11779 : NAND2_X2 port map( A1 => n37541, A2 => n16121, ZN => n15841);
   U11782 : NAND2_X1 port map( A1 => n36968, A2 => n16252, ZN => n37541);
   U11783 : NAND2_X2 port map( A1 => n3862, A2 => n19288, ZN => n17928);
   U11791 : OAI22_X2 port map( A1 => n14817, A2 => n22993, B1 => n22929, B2 => 
                           n20449, ZN => n3862);
   U11793 : NAND2_X2 port map( A1 => n30107, A2 => n35187, ZN => n30112);
   U11802 : NAND2_X2 port map( A1 => n33070, A2 => n4073, ZN => n30107);
   U11804 : XOR2_X1 port map( A1 => n26155, A2 => n26503, Z => n17171);
   U11812 : OR2_X1 port map( A1 => n875, A2 => n26934, Z => n34918);
   U11813 : AOI21_X1 port map( A1 => n9512, A2 => n30986, B => n9454, ZN => 
                           n37760);
   U11815 : INV_X2 port map( I => n8050, ZN => n451);
   U11816 : NAND2_X2 port map( A1 => n14278, A2 => n11956, ZN => n8050);
   U11818 : NAND2_X2 port map( A1 => n28344, A2 => n28346, ZN => n28716);
   U11822 : NOR2_X2 port map( A1 => n24328, A2 => n1607, ZN => n6585);
   U11826 : NAND2_X2 port map( A1 => n39664, A2 => n37460, ZN => n16921);
   U11829 : NAND2_X2 port map( A1 => n27346, A2 => n27345, ZN => n9185);
   U11835 : OAI21_X2 port map( A1 => n4668, A2 => n5027, B => n4667, ZN => 
                           n27346);
   U11839 : AOI22_X2 port map( A1 => n3708, A2 => n23523, B1 => n34959, B2 => 
                           n5258, ZN => n23589);
   U11841 : NAND2_X2 port map( A1 => n35361, A2 => n30815, ZN => n3708);
   U11844 : XOR2_X1 port map( A1 => n26462, A2 => n19973, Z => n10113);
   U11847 : XOR2_X1 port map( A1 => n1505, A2 => n12649, Z => n26462);
   U11849 : XOR2_X1 port map( A1 => n3501, A2 => n27745, Z => n14977);
   U11852 : XOR2_X1 port map( A1 => n37542, A2 => n25185, Z => n10926);
   U11855 : XOR2_X1 port map( A1 => n25184, A2 => n39146, Z => n37542);
   U11858 : XOR2_X1 port map( A1 => n10100, A2 => n1614, Z => n39344);
   U11860 : NAND2_X1 port map( A1 => n15919, A2 => n32690, ZN => n38866);
   U11862 : INV_X2 port map( I => n11219, ZN => n39126);
   U11865 : NAND3_X2 port map( A1 => n38734, A2 => n34535, A3 => n27398, ZN => 
                           n35243);
   U11869 : NAND2_X2 port map( A1 => n10856, A2 => n37543, ZN => n29050);
   U11873 : AOI22_X2 port map( A1 => n38275, A2 => n18996, B1 => n36663, B2 => 
                           n36076, ZN => n37543);
   U11874 : NAND2_X2 port map( A1 => n37545, A2 => n37544, ZN => n37915);
   U11877 : INV_X2 port map( I => n777, ZN => n37544);
   U11878 : XOR2_X1 port map( A1 => n11250, A2 => n37546, Z => n32474);
   U11890 : XOR2_X1 port map( A1 => n27812, A2 => n27813, Z => n37546);
   U11893 : NAND2_X1 port map( A1 => n20923, A2 => n12754, ZN => n21606);
   U11895 : NAND2_X2 port map( A1 => n37548, A2 => n37547, ZN => n36810);
   U11897 : OAI21_X2 port map( A1 => n22869, A2 => n22870, B => n16963, ZN => 
                           n37547);
   U11901 : XOR2_X1 port map( A1 => n26205, A2 => n26462, Z => n3780);
   U11904 : AOI21_X2 port map( A1 => n14146, A2 => n10290, B => n13677, ZN => 
                           n14145);
   U11906 : NOR2_X2 port map( A1 => n1014, A2 => n31205, ZN => n10290);
   U11910 : AND2_X1 port map( A1 => n23493, A2 => n34603, Z => n37906);
   U11911 : NOR2_X1 port map( A1 => n9452, A2 => n37760, ZN => n9513);
   U11912 : NOR2_X1 port map( A1 => n12331, A2 => n22929, ZN => n22991);
   U11916 : INV_X2 port map( I => n12100, ZN => n12331);
   U11917 : XOR2_X1 port map( A1 => n12102, A2 => n9595, Z => n12100);
   U11919 : NAND2_X1 port map( A1 => n37557, A2 => n28503, ZN => n37556);
   U11920 : NOR2_X2 port map( A1 => n36912, A2 => n39426, ZN => n37550);
   U11921 : NOR2_X2 port map( A1 => n35781, A2 => n37551, ZN => n38478);
   U11926 : AND2_X1 port map( A1 => n25882, A2 => n840, Z => n31471);
   U11927 : XOR2_X1 port map( A1 => n38022, A2 => n5841, Z => n23807);
   U11928 : NAND2_X2 port map( A1 => n37625, A2 => n10853, ZN => n9875);
   U11930 : OR2_X1 port map( A1 => n39417, A2 => n39628, Z => n36984);
   U11933 : NAND3_X2 port map( A1 => n17191, A2 => n28756, A3 => n28398, ZN => 
                           n17190);
   U11934 : INV_X1 port map( I => n14369, ZN => n1552);
   U11936 : AND2_X2 port map( A1 => n14369, A2 => n37553, Z => n25603);
   U11942 : XOR2_X1 port map( A1 => n8713, A2 => n31075, Z => n14369);
   U11943 : OAI21_X1 port map( A1 => n17369, A2 => n29662, B => n29660, ZN => 
                           n32290);
   U11945 : INV_X1 port map( I => n29641, ZN => n17369);
   U11947 : AOI22_X2 port map( A1 => n29638, A2 => n29761, B1 => n29637, B2 => 
                           n1178, ZN => n29641);
   U11948 : XOR2_X1 port map( A1 => n9939, A2 => n15592, Z => n7076);
   U11949 : XOR2_X1 port map( A1 => n589, A2 => n14835, Z => n14834);
   U11954 : XOR2_X1 port map( A1 => n3342, A2 => n34375, Z => n589);
   U11955 : XOR2_X1 port map( A1 => n37554, A2 => n14147, Z => n13091);
   U11959 : XOR2_X1 port map( A1 => n27790, A2 => n39410, Z => n37554);
   U11962 : XOR2_X1 port map( A1 => n26356, A2 => n26357, Z => n20082);
   U11970 : NAND2_X2 port map( A1 => n1849, A2 => n1850, ZN => n26356);
   U11971 : AND2_X1 port map( A1 => n6056, A2 => n4382, Z => n25792);
   U11973 : OAI22_X2 port map( A1 => n37555, A2 => n6698, B1 => n6697, B2 => 
                           n28178, ZN => n28966);
   U11980 : NAND2_X2 port map( A1 => n6684, A2 => n1637, ZN => n9346);
   U11981 : XOR2_X1 port map( A1 => n25280, A2 => n6185, Z => n10582);
   U11982 : AOI21_X2 port map( A1 => n20505, A2 => n3630, B => n3629, ZN => 
                           n25280);
   U11983 : XOR2_X1 port map( A1 => n36366, A2 => n26502, Z => n26512);
   U11984 : OAI22_X2 port map( A1 => n38084, A2 => n13891, B1 => n37558, B2 => 
                           n37556, ZN => n29041);
   U11988 : NAND2_X2 port map( A1 => n36798, A2 => n598, ZN => n25822);
   U11990 : AOI22_X2 port map( A1 => n12931, A2 => n9439, B1 => n9440, B2 => 
                           n38338, ZN => n598);
   U11992 : NOR2_X2 port map( A1 => n4941, A2 => n30837, ZN => n28503);
   U11995 : NAND2_X2 port map( A1 => n18131, A2 => n31087, ZN => n4941);
   U12003 : NAND2_X1 port map( A1 => n12675, A2 => n13811, ZN => n38959);
   U12006 : AND2_X2 port map( A1 => n18342, A2 => n24271, Z => n18698);
   U12009 : NOR2_X2 port map( A1 => n2522, A2 => n1081, ZN => n2519);
   U12015 : NOR2_X2 port map( A1 => n12081, A2 => n19544, ZN => n39393);
   U12016 : NAND2_X2 port map( A1 => n37788, A2 => n37562, ZN => n27438);
   U12022 : NAND2_X2 port map( A1 => n34820, A2 => n37563, ZN => n8966);
   U12024 : OAI21_X2 port map( A1 => n30944, A2 => n31490, B => n305, ZN => 
                           n37563);
   U12026 : XOR2_X1 port map( A1 => n26246, A2 => n26245, Z => n26324);
   U12027 : NOR2_X2 port map( A1 => n4884, A2 => n25531, ZN => n26246);
   U12028 : NAND3_X2 port map( A1 => n37028, A2 => n25916, A3 => n1016, ZN => 
                           n25917);
   U12029 : BUF_X2 port map( I => n3937, Z => n4001);
   U12032 : OAI21_X1 port map( A1 => n25644, A2 => n25666, B => n4468, ZN => 
                           n4466);
   U12034 : OR2_X1 port map( A1 => n5062, A2 => n28197, Z => n33804);
   U12036 : OR2_X1 port map( A1 => n12924, A2 => n36396, Z => n18997);
   U12037 : XOR2_X1 port map( A1 => n29829, A2 => n29081, Z => n28893);
   U12038 : OAI21_X2 port map( A1 => n27033, A2 => n37205, B => n27032, ZN => 
                           n27774);
   U12042 : NAND2_X1 port map( A1 => n35380, A2 => n4700, ZN => n37657);
   U12046 : OAI21_X2 port map( A1 => n299, A2 => n17613, B => n20381, ZN => 
                           n35903);
   U12051 : XOR2_X1 port map( A1 => n37564, A2 => n19498, Z => Ciphertext(100))
                           ;
   U12053 : NAND2_X1 port map( A1 => n29749, A2 => n31477, ZN => n37564);
   U12054 : NAND2_X1 port map( A1 => n32802, A2 => n24900, ZN => n17475);
   U12059 : NAND2_X1 port map( A1 => n29632, A2 => n1398, ZN => n37565);
   U12064 : XOR2_X1 port map( A1 => n26141, A2 => n21086, Z => n34966);
   U12065 : OAI21_X2 port map( A1 => n3044, A2 => n38073, B => n37566, ZN => 
                           n35925);
   U12066 : NAND3_X2 port map( A1 => n37737, A2 => n39279, A3 => n34011, ZN => 
                           n37566);
   U12067 : NAND3_X2 port map( A1 => n19400, A2 => n39389, A3 => n37051, ZN => 
                           n13535);
   U12069 : NAND2_X1 port map( A1 => n36177, A2 => n9267, ZN => n38788);
   U12079 : XOR2_X1 port map( A1 => n37567, A2 => n31062, Z => Ciphertext(62));
   U12083 : NAND3_X2 port map( A1 => n28905, A2 => n28906, A3 => n28907, ZN => 
                           n37567);
   U12085 : XOR2_X1 port map( A1 => n35062, A2 => n23930, Z => n23787);
   U12086 : NOR2_X1 port map( A1 => n14278, A2 => n11956, ZN => n34567);
   U12089 : OAI21_X2 port map( A1 => n6160, A2 => n31275, B => n31785, ZN => 
                           n11956);
   U12093 : NAND2_X2 port map( A1 => n4579, A2 => n4580, ZN => n15135);
   U12099 : XOR2_X1 port map( A1 => n37568, A2 => n34017, Z => Ciphertext(11));
   U12100 : AOI22_X1 port map( A1 => n29226, A2 => n35264, B1 => n1378, B2 => 
                           n12691, ZN => n37568);
   U12121 : XOR2_X1 port map( A1 => n9874, A2 => n22572, Z => n22625);
   U12125 : XOR2_X1 port map( A1 => n33194, A2 => n26548, Z => n26408);
   U12129 : NAND2_X2 port map( A1 => n25984, A2 => n25983, ZN => n26548);
   U12130 : XOR2_X1 port map( A1 => n6559, A2 => n6560, Z => n23785);
   U12134 : OAI21_X2 port map( A1 => n37569, A2 => n17674, B => n10763, ZN => 
                           n17673);
   U12140 : XOR2_X1 port map( A1 => n37038, A2 => n31181, Z => n25180);
   U12141 : NAND2_X2 port map( A1 => n37570, A2 => n19702, ZN => n38713);
   U12143 : AOI21_X2 port map( A1 => n25527, A2 => n19701, B => n1539, ZN => 
                           n37570);
   U12148 : NOR2_X1 port map( A1 => n33266, A2 => n39026, ZN => n38257);
   U12150 : NOR2_X2 port map( A1 => n3190, A2 => n7950, ZN => n3441);
   U12151 : XOR2_X1 port map( A1 => n1260, A2 => n12297, Z => n12296);
   U12161 : AOI22_X2 port map( A1 => n24701, A2 => n6791, B1 => n24270, B2 => 
                           n24530, ZN => n25259);
   U12163 : XOR2_X1 port map( A1 => n29096, A2 => n37571, Z => n12157);
   U12168 : INV_X2 port map( I => n14956, ZN => n37571);
   U12169 : OAI21_X2 port map( A1 => n37572, A2 => n23372, B => n38623, ZN => 
                           n13395);
   U12173 : OAI21_X2 port map( A1 => n34386, A2 => n32061, B => n37573, ZN => 
                           n37572);
   U12174 : NAND2_X2 port map( A1 => n34386, A2 => n23370, ZN => n37573);
   U12177 : NOR2_X1 port map( A1 => n13432, A2 => n13431, ZN => n37620);
   U12179 : XOR2_X1 port map( A1 => n16805, A2 => n37574, Z => n32822);
   U12180 : XOR2_X1 port map( A1 => n37860, A2 => n767, Z => n37574);
   U12182 : NOR2_X2 port map( A1 => n11470, A2 => n11208, ZN => n18960);
   U12186 : NAND3_X2 port map( A1 => n9303, A2 => n25756, A3 => n12931, ZN => 
                           n37949);
   U12188 : XOR2_X1 port map( A1 => n25324, A2 => n24931, Z => n24946);
   U12190 : NAND2_X2 port map( A1 => n19356, A2 => n24706, ZN => n25324);
   U12193 : NAND2_X2 port map( A1 => n37575, A2 => n7488, ZN => n32691);
   U12196 : NOR2_X2 port map( A1 => n36302, A2 => n19927, ZN => n37575);
   U12209 : XOR2_X1 port map( A1 => n38455, A2 => n11402, Z => n3785);
   U12211 : XOR2_X1 port map( A1 => n27483, A2 => n27535, Z => n36628);
   U12212 : NAND2_X2 port map( A1 => n29895, A2 => n37576, ZN => n19097);
   U12213 : OAI21_X2 port map( A1 => n32498, A2 => n32499, B => n17240, ZN => 
                           n37576);
   U12217 : NOR2_X1 port map( A1 => n30747, A2 => n1178, ZN => n15376);
   U12219 : BUF_X4 port map( I => n25324, Z => n37943);
   U12221 : XOR2_X1 port map( A1 => n18498, A2 => n27865, Z => n33642);
   U12229 : XOR2_X1 port map( A1 => n27737, A2 => n27736, Z => n27865);
   U12230 : AOI21_X2 port map( A1 => n37578, A2 => n37577, B => n14652, ZN => 
                           n28896);
   U12231 : NOR2_X2 port map( A1 => n28438, A2 => n37579, ZN => n37578);
   U12232 : NAND2_X2 port map( A1 => n35123, A2 => n38078, ZN => n38816);
   U12233 : XOR2_X1 port map( A1 => n27722, A2 => n27721, Z => n36603);
   U12237 : XOR2_X1 port map( A1 => n27593, A2 => n27703, Z => n27722);
   U12238 : OAI21_X2 port map( A1 => n1011, A2 => n1243, B => n30629, ZN => 
                           n11980);
   U12247 : OAI21_X2 port map( A1 => n13534, A2 => n13533, B => n12705, ZN => 
                           n30629);
   U12249 : XOR2_X1 port map( A1 => n27777, A2 => n27511, Z => n608);
   U12254 : NAND2_X2 port map( A1 => n27052, A2 => n27051, ZN => n27777);
   U12258 : NAND2_X1 port map( A1 => n8820, A2 => n8822, ZN => n11514);
   U12262 : NAND2_X2 port map( A1 => n17231, A2 => n17232, ZN => n25801);
   U12264 : OAI21_X2 port map( A1 => n36344, A2 => n26857, B => n1491, ZN => 
                           n34985);
   U12266 : XOR2_X1 port map( A1 => n33578, A2 => n2222, Z => n6226);
   U12268 : NAND2_X2 port map( A1 => n19636, A2 => n19637, ZN => n25387);
   U12270 : NAND2_X2 port map( A1 => n11496, A2 => n24741, ZN => n19636);
   U12272 : XOR2_X1 port map( A1 => n1184, A2 => n14941, Z => n29126);
   U12273 : BUF_X4 port map( I => n15988, Z => n1006);
   U12276 : NOR2_X2 port map( A1 => n37581, A2 => n6423, ZN => n23310);
   U12278 : NOR2_X2 port map( A1 => n16416, A2 => n23013, ZN => n37581);
   U12280 : BUF_X2 port map( I => n36571, Z => n37582);
   U12281 : NAND2_X2 port map( A1 => n37583, A2 => n6509, ZN => n7565);
   U12283 : NOR2_X2 port map( A1 => n18698, A2 => n37264, ZN => n37583);
   U12284 : XOR2_X1 port map( A1 => n25016, A2 => n35900, Z => n9939);
   U12288 : NAND2_X2 port map( A1 => n8108, A2 => n11738, ZN => n25016);
   U12291 : BUF_X2 port map( I => n19728, Z => n37585);
   U12297 : NOR2_X2 port map( A1 => n29468, A2 => n9105, ZN => n12369);
   U12299 : NOR2_X2 port map( A1 => n39060, A2 => n8924, ZN => n29468);
   U12301 : OAI21_X2 port map( A1 => n12167, A2 => n29644, B => n37586, ZN => 
                           n10030);
   U12305 : NAND2_X2 port map( A1 => n37743, A2 => n29645, ZN => n37586);
   U12312 : INV_X2 port map( I => n37587, ZN => n35233);
   U12315 : XOR2_X1 port map( A1 => n9555, A2 => n6455, Z => n37588);
   U12319 : XOR2_X1 port map( A1 => n10498, A2 => n8793, Z => n9266);
   U12322 : AOI22_X2 port map( A1 => n10901, A2 => n10903, B1 => n39302, B2 => 
                           n10902, ZN => n37625);
   U12325 : XOR2_X1 port map( A1 => n17757, A2 => n26463, Z => n12145);
   U12326 : NOR3_X2 port map( A1 => n13440, A2 => n18314, A3 => n17297, ZN => 
                           n26463);
   U12327 : NOR2_X2 port map( A1 => n37591, A2 => n37590, ZN => n38965);
   U12328 : NAND3_X1 port map( A1 => n16633, A2 => n4410, A3 => n37235, ZN => 
                           n37592);
   U12330 : AND2_X1 port map( A1 => n26642, A2 => n26644, Z => n39179);
   U12334 : NAND2_X2 port map( A1 => n9694, A2 => n26031, ZN => n25915);
   U12338 : NAND2_X2 port map( A1 => n34260, A2 => n25605, ZN => n9694);
   U12339 : AOI21_X2 port map( A1 => n31516, A2 => n30747, B => n19599, ZN => 
                           n30746);
   U12341 : NOR2_X1 port map( A1 => n9893, A2 => n14369, ZN => n12616);
   U12342 : XOR2_X1 port map( A1 => n25102, A2 => n10611, Z => n37998);
   U12348 : NOR2_X2 port map( A1 => n3509, A2 => n36450, ZN => n2561);
   U12351 : NAND2_X2 port map( A1 => n7466, A2 => n39380, ZN => n3509);
   U12353 : NAND2_X2 port map( A1 => n167, A2 => n19425, ZN => n26943);
   U12354 : INV_X2 port map( I => n35176, ZN => n19272);
   U12357 : XOR2_X1 port map( A1 => n37594, A2 => n37639, Z => n39750);
   U12359 : XOR2_X1 port map( A1 => n33587, A2 => n27556, Z => n37594);
   U12361 : INV_X2 port map( I => n5745, ZN => n11083);
   U12362 : OR2_X1 port map( A1 => n17119, A2 => n39810, Z => n17128);
   U12364 : OR2_X1 port map( A1 => n18682, A2 => n16528, Z => n18478);
   U12367 : XOR2_X1 port map( A1 => n37595, A2 => n1371, Z => Ciphertext(112));
   U12369 : NOR3_X1 port map( A1 => n36410, A2 => n36365, A3 => n6650, ZN => 
                           n37595);
   U12372 : NAND2_X2 port map( A1 => n12178, A2 => n20845, ZN => n28500);
   U12375 : OR2_X1 port map( A1 => n12682, A2 => n3873, Z => n26859);
   U12381 : XOR2_X1 port map( A1 => n26486, A2 => n10668, Z => n3732);
   U12382 : XOR2_X1 port map( A1 => n26542, A2 => n35214, Z => n26486);
   U12384 : OAI21_X2 port map( A1 => n3631, A2 => n3699, B => n3698, ZN => 
                           n28924);
   U12391 : NAND2_X2 port map( A1 => n37596, A2 => n30372, ZN => n31362);
   U12392 : XOR2_X1 port map( A1 => n11116, A2 => n15202, Z => n11115);
   U12394 : XOR2_X1 port map( A1 => n25166, A2 => n25007, Z => n3495);
   U12401 : INV_X2 port map( I => n18870, ZN => n17346);
   U12403 : NOR2_X1 port map( A1 => n35881, A2 => n5392, ZN => n21916);
   U12418 : NAND2_X2 port map( A1 => n37597, A2 => n12249, ZN => n14283);
   U12419 : NAND2_X2 port map( A1 => n37967, A2 => n1127, ZN => n37597);
   U12422 : OR2_X1 port map( A1 => n38976, A2 => n30800, Z => n20756);
   U12424 : BUF_X2 port map( I => n34977, Z => n37598);
   U12429 : NAND2_X2 port map( A1 => n19340, A2 => n37599, ZN => n25924);
   U12435 : NAND2_X2 port map( A1 => n25803, A2 => n16407, ZN => n37599);
   U12437 : XOR2_X1 port map( A1 => n37600, A2 => n20819, Z => n29196);
   U12440 : XOR2_X1 port map( A1 => n28502, A2 => n29105, Z => n37600);
   U12441 : INV_X2 port map( I => n29626, ZN => n29618);
   U12442 : NAND3_X2 port map( A1 => n34097, A2 => n8996, A3 => n8999, ZN => 
                           n29626);
   U12448 : NAND2_X2 port map( A1 => n36986, A2 => n2774, ZN => n34599);
   U12450 : NAND2_X2 port map( A1 => n37601, A2 => n24167, ZN => n10980);
   U12456 : XOR2_X1 port map( A1 => n10215, A2 => n21253, Z => n8923);
   U12467 : AOI22_X2 port map( A1 => n29557, A2 => n29558, B1 => n29559, B2 => 
                           n29560, ZN => n21158);
   U12468 : XOR2_X1 port map( A1 => n28835, A2 => n29816, Z => n10899);
   U12469 : XOR2_X1 port map( A1 => n36928, A2 => n296, Z => n28835);
   U12471 : XOR2_X1 port map( A1 => n23732, A2 => n714, Z => n37834);
   U12474 : XOR2_X1 port map( A1 => n23888, A2 => n23886, Z => n23732);
   U12475 : INV_X2 port map( I => n29124, ZN => n38610);
   U12478 : NAND2_X2 port map( A1 => n37759, A2 => n36313, ZN => n29124);
   U12481 : NOR2_X2 port map( A1 => n10171, A2 => n15135, ZN => n26791);
   U12483 : XOR2_X1 port map( A1 => n26441, A2 => n4622, Z => n26254);
   U12484 : NOR2_X2 port map( A1 => n34413, A2 => n11010, ZN => n26441);
   U12485 : XOR2_X1 port map( A1 => n37602, A2 => n26374, Z => n26272);
   U12488 : XOR2_X1 port map( A1 => n32442, A2 => n13814, Z => n37602);
   U12490 : OR2_X2 port map( A1 => n2616, A2 => n17351, Z => n7267);
   U12493 : OAI21_X2 port map( A1 => n27026, A2 => n27174, B => n37603, ZN => 
                           n7808);
   U12495 : AND2_X1 port map( A1 => n5392, A2 => n21912, Z => n21913);
   U12497 : OAI22_X1 port map( A1 => n30110, A2 => n10118, B1 => n30111, B2 => 
                           n30112, ZN => n39578);
   U12498 : OAI22_X2 port map( A1 => n37604, A2 => n12066, B1 => n12065, B2 => 
                           n2140, ZN => n7861);
   U12499 : BUF_X4 port map( I => n15579, Z => n34386);
   U12503 : OR3_X1 port map( A1 => n27969, A2 => n14451, A3 => n19366, Z => 
                           n20919);
   U12512 : XOR2_X1 port map( A1 => n7061, A2 => n7059, Z => n19764);
   U12513 : XOR2_X1 port map( A1 => n27842, A2 => n27754, Z => n27524);
   U12514 : NOR2_X2 port map( A1 => n27060, A2 => n27061, ZN => n27842);
   U12515 : NAND3_X1 port map( A1 => n28498, A2 => n33591, A3 => n28497, ZN => 
                           n12178);
   U12529 : NAND2_X2 port map( A1 => n35491, A2 => n1882, ZN => n28498);
   U12530 : NOR2_X2 port map( A1 => n37607, A2 => n37606, ZN => n20454);
   U12536 : OAI22_X2 port map( A1 => n19276, A2 => n7676, B1 => n27118, B2 => 
                           n32976, ZN => n37606);
   U12538 : AOI21_X1 port map( A1 => n20455, A2 => n27006, B => n35184, ZN => 
                           n37607);
   U12543 : XOR2_X1 port map( A1 => n8474, A2 => n28988, Z => n10541);
   U12544 : XOR2_X1 port map( A1 => n31615, A2 => n28500, Z => n28988);
   U12545 : NAND2_X2 port map( A1 => n26657, A2 => n37608, ZN => n7975);
   U12553 : AOI22_X2 port map( A1 => n13645, A2 => n26701, B1 => n13644, B2 => 
                           n36244, ZN => n37608);
   U12558 : XOR2_X1 port map( A1 => n10153, A2 => n37609, Z => n7980);
   U12560 : XOR2_X1 port map( A1 => n33812, A2 => n38209, Z => n37609);
   U12562 : XOR2_X1 port map( A1 => n10792, A2 => n16900, Z => n25251);
   U12573 : AOI22_X2 port map( A1 => n35180, A2 => n29525, B1 => n29527, B2 => 
                           n29531, ZN => n29536);
   U12574 : AOI21_X2 port map( A1 => n14780, A2 => n24275, B => n364, ZN => 
                           n2616);
   U12576 : NAND2_X2 port map( A1 => n39250, A2 => n10321, ZN => n26097);
   U12578 : XOR2_X1 port map( A1 => n5609, A2 => n37610, Z => n5732);
   U12579 : XOR2_X1 port map( A1 => n17910, A2 => n3734, Z => n37610);
   U12580 : XOR2_X1 port map( A1 => n37611, A2 => n39103, Z => n13429);
   U12581 : XOR2_X1 port map( A1 => n5913, A2 => n5915, Z => n37611);
   U12582 : BUF_X2 port map( I => n7935, Z => n37612);
   U12584 : XOR2_X1 port map( A1 => n22774, A2 => n22494, Z => n387);
   U12585 : XOR2_X1 port map( A1 => n22600, A2 => n13704, Z => n22774);
   U12588 : XOR2_X1 port map( A1 => n12069, A2 => n13800, Z => n39171);
   U12595 : NAND3_X2 port map( A1 => n3221, A2 => n11465, A3 => n16791, ZN => 
                           n29289);
   U12597 : XOR2_X1 port map( A1 => n36743, A2 => n26184, Z => n32339);
   U12601 : XOR2_X1 port map( A1 => n17048, A2 => n26567, Z => n26184);
   U12606 : AND2_X1 port map( A1 => n32284, A2 => n35777, Z => n37615);
   U12607 : OAI22_X2 port map( A1 => n29541, A2 => n1394, B1 => n29546, B2 => 
                           n29558, ZN => n29560);
   U12619 : NAND2_X2 port map( A1 => n37645, A2 => n37616, ZN => n25971);
   U12621 : XOR2_X1 port map( A1 => n18975, A2 => n26386, Z => n18974);
   U12628 : XOR2_X1 port map( A1 => n26511, A2 => n26224, Z => n26386);
   U12631 : INV_X2 port map( I => n20877, ZN => n24017);
   U12635 : XOR2_X1 port map( A1 => n23778, A2 => n37617, Z => n20877);
   U12636 : INV_X2 port map( I => n23899, ZN => n37617);
   U12640 : XOR2_X1 port map( A1 => n8303, A2 => n28886, Z => n29151);
   U12641 : OAI21_X2 port map( A1 => n21026, A2 => n28298, B => n21024, ZN => 
                           n8303);
   U12646 : XOR2_X1 port map( A1 => n31524, A2 => n31127, Z => n38772);
   U12647 : NAND2_X2 port map( A1 => n32758, A2 => n11719, ZN => n31524);
   U12654 : OR2_X2 port map( A1 => n10111, A2 => n20891, Z => n26926);
   U12655 : XOR2_X1 port map( A1 => n16647, A2 => n9590, Z => n39443);
   U12657 : NAND3_X2 port map( A1 => n18352, A2 => n37618, A3 => n18353, ZN => 
                           n33645);
   U12658 : NAND2_X2 port map( A1 => n37619, A2 => n12537, ZN => n34171);
   U12659 : INV_X2 port map( I => n32146, ZN => n37619);
   U12663 : XOR2_X1 port map( A1 => n37620, A2 => n33184, Z => Ciphertext(48));
   U12667 : OAI22_X2 port map( A1 => n17066, A2 => n24383, B1 => n18907, B2 => 
                           n18402, ZN => n20795);
   U12669 : OAI21_X2 port map( A1 => n30357, A2 => n15389, B => n37621, ZN => 
                           n28245);
   U12671 : NAND2_X2 port map( A1 => n15389, A2 => n28240, ZN => n37621);
   U12673 : NOR2_X1 port map( A1 => n39554, A2 => n18668, ZN => n19034);
   U12675 : BUF_X2 port map( I => n28159, Z => n37623);
   U12680 : XOR2_X1 port map( A1 => n4999, A2 => n5646, Z => n11543);
   U12685 : XOR2_X1 port map( A1 => n17563, A2 => n8113, Z => n6403);
   U12688 : OAI22_X2 port map( A1 => n27057, A2 => n27368, B1 => n27056, B2 => 
                           n33050, ZN => n27511);
   U12689 : NOR2_X1 port map( A1 => n31788, A2 => n30154, ZN => n34065);
   U12690 : AOI21_X2 port map( A1 => n28149, A2 => n27622, B => n17753, ZN => 
                           n37626);
   U12698 : NAND2_X2 port map( A1 => n21144, A2 => n27276, ZN => n27059);
   U12703 : XOR2_X1 port map( A1 => n27645, A2 => n27494, Z => n10498);
   U12704 : XOR2_X1 port map( A1 => n14808, A2 => n10997, Z => n27645);
   U12713 : INV_X2 port map( I => n11126, ZN => n37624);
   U12717 : NAND2_X2 port map( A1 => n13179, A2 => n37626, ZN => n8743);
   U12718 : XOR2_X1 port map( A1 => n12865, A2 => n37627, Z => n5291);
   U12719 : XOR2_X1 port map( A1 => n16857, A2 => n33587, Z => n37627);
   U12720 : NOR3_X1 port map( A1 => n15004, A2 => n8493, A3 => n19604, ZN => 
                           n31369);
   U12721 : NOR2_X2 port map( A1 => n19454, A2 => n37628, ZN => n34378);
   U12724 : OAI22_X1 port map( A1 => n6692, A2 => n8529, B1 => n29937, B2 => 
                           n29935, ZN => n37628);
   U12725 : OR2_X1 port map( A1 => n3873, A2 => n14415, Z => n5263);
   U12727 : XOR2_X1 port map( A1 => n34812, A2 => n27554, Z => n11236);
   U12729 : NAND2_X2 port map( A1 => n2303, A2 => n2305, ZN => n27554);
   U12732 : NAND2_X1 port map( A1 => n34008, A2 => n27932, ZN => n8056);
   U12737 : NAND3_X2 port map( A1 => n37630, A2 => n11455, A3 => n11456, ZN => 
                           n22740);
   U12739 : NAND2_X1 port map( A1 => n3137, A2 => n11234, ZN => n37630);
   U12743 : XOR2_X1 port map( A1 => n37631, A2 => n39071, Z => n13540);
   U12745 : XOR2_X1 port map( A1 => n3932, A2 => n8884, Z => n37631);
   U12748 : INV_X2 port map( I => n3937, ZN => n20441);
   U12750 : NAND2_X2 port map( A1 => n37633, A2 => n8289, ZN => n31663);
   U12753 : OAI21_X2 port map( A1 => n33020, A2 => n33981, B => n28265, ZN => 
                           n37633);
   U12755 : AOI22_X2 port map( A1 => n9068, A2 => n24297, B1 => n12248, B2 => 
                           n37634, ZN => n19499);
   U12759 : NAND3_X2 port map( A1 => n37635, A2 => n4360, A3 => n4361, ZN => 
                           n15266);
   U12762 : INV_X4 port map( I => n19771, ZN => n28742);
   U12764 : NAND2_X2 port map( A1 => n34965, A2 => n406, ZN => n19771);
   U12765 : NAND3_X2 port map( A1 => n20994, A2 => n30231, A3 => n37636, ZN => 
                           n30249);
   U12766 : XOR2_X1 port map( A1 => n37899, A2 => n17850, Z => n17518);
   U12767 : OAI21_X1 port map( A1 => n36649, A2 => n38830, B => n37805, ZN => 
                           n38832);
   U12768 : NAND2_X1 port map( A1 => n38832, A2 => n38746, ZN => n9734);
   U12770 : XNOR2_X1 port map( A1 => n27703, A2 => n27595, ZN => n27831);
   U12773 : NAND2_X2 port map( A1 => n8601, A2 => n13792, ZN => n27595);
   U12774 : OAI22_X2 port map( A1 => n2338, A2 => n37671, B1 => n3235, B2 => 
                           n39298, ZN => n6160);
   U12777 : NAND3_X1 port map( A1 => n2803, A2 => n25484, A3 => n3985, ZN => 
                           n36459);
   U12778 : XOR2_X1 port map( A1 => n28967, A2 => n9035, Z => n37973);
   U12782 : NOR2_X2 port map( A1 => n37638, A2 => n37637, ZN => n28967);
   U12785 : INV_X2 port map( I => n17132, ZN => n38060);
   U12787 : NAND2_X2 port map( A1 => n7914, A2 => n28547, ZN => n35326);
   U12788 : NAND2_X2 port map( A1 => n7251, A2 => n11956, ZN => n7914);
   U12790 : BUF_X2 port map( I => n14415, Z => n278);
   U12791 : INV_X2 port map( I => n35657, ZN => n2870);
   U12792 : NAND2_X1 port map( A1 => n12869, A2 => n12552, ZN => n34826);
   U12794 : AOI21_X2 port map( A1 => n5365, A2 => n7612, B => n36407, ZN => 
                           n31702);
   U12798 : INV_X1 port map( I => n27390, ZN => n37641);
   U12800 : NOR2_X1 port map( A1 => n30358, A2 => n37641, ZN => n38146);
   U12802 : BUF_X2 port map( I => n38742, Z => n37643);
   U12803 : OAI22_X2 port map( A1 => n6691, A2 => n23060, B1 => n37629, B2 => 
                           n22925, ZN => n14743);
   U12805 : XOR2_X1 port map( A1 => n37644, A2 => n30170, Z => Ciphertext(175))
                           ;
   U12806 : NOR2_X2 port map( A1 => n38029, A2 => n7339, ZN => n37645);
   U12810 : XOR2_X1 port map( A1 => n8505, A2 => n37646, Z => n9945);
   U12811 : XOR2_X1 port map( A1 => n33248, A2 => n24055, Z => n37646);
   U12812 : NAND2_X2 port map( A1 => n25667, A2 => n37647, ZN => n25936);
   U12814 : INV_X2 port map( I => n5768, ZN => n5124);
   U12815 : NAND2_X2 port map( A1 => n24584, A2 => n24583, ZN => n5768);
   U12816 : NAND3_X1 port map( A1 => n37648, A2 => n10642, A3 => n28074, ZN => 
                           n3461);
   U12817 : NAND2_X2 port map( A1 => n28273, A2 => n988, ZN => n37648);
   U12834 : NOR2_X1 port map( A1 => n19615, A2 => n38742, ZN => n26769);
   U12836 : XOR2_X1 port map( A1 => n35222, A2 => n29088, Z => n29001);
   U12837 : NAND2_X2 port map( A1 => n6370, A2 => n6371, ZN => n29088);
   U12838 : NAND2_X2 port map( A1 => n13213, A2 => n19918, ZN => n27118);
   U12840 : NAND2_X2 port map( A1 => n38871, A2 => n13890, ZN => n29820);
   U12841 : NOR2_X2 port map( A1 => n38924, A2 => n36834, ZN => n38871);
   U12842 : XOR2_X1 port map( A1 => n3560, A2 => n1938, Z => n3559);
   U12844 : XOR2_X1 port map( A1 => n28987, A2 => n39233, Z => n37650);
   U12845 : XOR2_X1 port map( A1 => n7374, A2 => n36510, Z => n36931);
   U12847 : NAND2_X2 port map( A1 => n13860, A2 => n37030, ZN => n1746);
   U12853 : INV_X2 port map( I => n5227, ZN => n12394);
   U12857 : XNOR2_X1 port map( A1 => n5228, A2 => n5229, ZN => n5227);
   U12859 : NAND2_X2 port map( A1 => n23225, A2 => n14365, ZN => n37851);
   U12860 : XOR2_X1 port map( A1 => n19071, A2 => n37221, Z => n16942);
   U12863 : XOR2_X1 port map( A1 => n35936, A2 => n15202, Z => n19071);
   U12865 : BUF_X2 port map( I => n24408, Z => n37651);
   U12870 : INV_X2 port map( I => n37656, ZN => n38130);
   U12871 : NAND3_X2 port map( A1 => n23169, A2 => n36554, A3 => n23167, ZN => 
                           n37656);
   U12876 : NAND2_X2 port map( A1 => n37657, A2 => n17500, ZN => n21110);
   U12878 : XOR2_X1 port map( A1 => n8302, A2 => n35241, Z => n9947);
   U12879 : NAND2_X2 port map( A1 => n23081, A2 => n3145, ZN => n23566);
   U12883 : XOR2_X1 port map( A1 => n37658, A2 => n37037, Z => n32118);
   U12884 : XOR2_X1 port map( A1 => n3110, A2 => n25151, Z => n25198);
   U12888 : NOR3_X2 port map( A1 => n21887, A2 => n21889, A3 => n16302, ZN => 
                           n15812);
   U12889 : XOR2_X1 port map( A1 => n25063, A2 => n18543, Z => n3292);
   U12891 : XOR2_X1 port map( A1 => n25133, A2 => n24857, Z => n18543);
   U12893 : AOI22_X2 port map( A1 => n5791, A2 => n31829, B1 => n5790, B2 => 
                           n17556, ZN => n2932);
   U12901 : NAND2_X2 port map( A1 => n20153, A2 => n13545, ZN => n25483);
   U12906 : AOI22_X1 port map( A1 => n23256, A2 => n23515, B1 => n4638, B2 => 
                           n4637, ZN => n36279);
   U12908 : XNOR2_X1 port map( A1 => n15368, A2 => n37833, ZN => n39186);
   U12920 : XOR2_X1 port map( A1 => n13852, A2 => n8475, Z => n8474);
   U12923 : AOI21_X2 port map( A1 => n35621, A2 => n10758, B => n10757, ZN => 
                           n13852);
   U12926 : BUF_X2 port map( I => n35920, Z => n37660);
   U12928 : NOR2_X2 port map( A1 => n35449, A2 => n18909, ZN => n4636);
   U12933 : XOR2_X1 port map( A1 => n38581, A2 => n24924, Z => n25191);
   U12936 : NAND2_X2 port map( A1 => n39496, A2 => n17267, ZN => n38581);
   U12937 : AOI21_X1 port map( A1 => n29593, A2 => n38420, B => n31374, ZN => 
                           n38941);
   U12940 : NOR2_X1 port map( A1 => n63, A2 => n29946, ZN => n14592);
   U12945 : INV_X2 port map( I => n2792, ZN => n6652);
   U12948 : INV_X2 port map( I => n37662, ZN => n25718);
   U12956 : NAND2_X2 port map( A1 => n37663, A2 => n1855, ZN => n26125);
   U12957 : NAND2_X2 port map( A1 => n1425, A2 => n5418, ZN => n28365);
   U12960 : AOI21_X2 port map( A1 => n37664, A2 => n38073, B => n35925, ZN => 
                           n10012);
   U12962 : NAND3_X2 port map( A1 => n28146, A2 => n28145, A3 => n28144, ZN => 
                           n28686);
   U12970 : XOR2_X1 port map( A1 => n22391, A2 => n22542, Z => n20294);
   U12974 : NAND2_X2 port map( A1 => n10744, A2 => n10742, ZN => n22391);
   U12981 : INV_X2 port map( I => n16237, ZN => n1477);
   U12982 : NAND2_X2 port map( A1 => n30617, A2 => n39542, ZN => n16237);
   U12983 : XOR2_X1 port map( A1 => n6318, A2 => n37666, Z => n20726);
   U12987 : XOR2_X1 port map( A1 => n37665, A2 => n19786, Z => Ciphertext(148))
                           ;
   U12990 : NAND4_X2 port map( A1 => n30075, A2 => n30072, A3 => n30074, A4 => 
                           n30073, ZN => n37665);
   U12992 : OAI21_X2 port map( A1 => n30043, A2 => n29998, B => n29997, ZN => 
                           n35649);
   U12993 : OAI21_X2 port map( A1 => n35653, A2 => n20125, B => n35649, ZN => 
                           n6919);
   U12994 : INV_X2 port map( I => n3815, ZN => n30077);
   U12995 : NAND2_X2 port map( A1 => n34378, A2 => n31499, ZN => n3815);
   U13000 : XOR2_X1 port map( A1 => n6316, A2 => n20727, Z => n37666);
   U13006 : OR2_X1 port map( A1 => n25309, A2 => n825, Z => n18233);
   U13014 : XOR2_X1 port map( A1 => n37667, A2 => n27706, Z => n20511);
   U13016 : XOR2_X1 port map( A1 => n20513, A2 => n35177, Z => n37667);
   U13018 : XOR2_X1 port map( A1 => n37668, A2 => n6991, Z => n5899);
   U13019 : XOR2_X1 port map( A1 => n6522, A2 => n26500, Z => n3995);
   U13021 : NAND2_X1 port map( A1 => n18234, A2 => n18233, ZN => n37669);
   U13031 : XOR2_X1 port map( A1 => n9030, A2 => n30913, Z => n6522);
   U13032 : XOR2_X1 port map( A1 => n22789, A2 => n20335, Z => n22522);
   U13035 : NOR2_X2 port map( A1 => n11440, A2 => n11439, ZN => n22789);
   U13038 : NOR2_X2 port map( A1 => n31769, A2 => n18776, ZN => n39424);
   U13053 : NAND3_X2 port map( A1 => n39083, A2 => n30213, A3 => n14387, ZN => 
                           n39142);
   U13060 : NAND2_X2 port map( A1 => n13488, A2 => n36769, ZN => n6533);
   U13063 : OAI21_X2 port map( A1 => n18743, A2 => n32131, B => n19061, ZN => 
                           n39249);
   U13067 : NAND2_X2 port map( A1 => n39249, A2 => n4570, ZN => n30908);
   U13070 : XOR2_X1 port map( A1 => n5395, A2 => n37786, Z => n8148);
   U13071 : NAND2_X2 port map( A1 => n39222, A2 => n37670, ZN => n27211);
   U13073 : NAND2_X1 port map( A1 => n35612, A2 => n35613, ZN => n37670);
   U13074 : NOR2_X2 port map( A1 => n33407, A2 => n3057, ZN => n38398);
   U13076 : INV_X4 port map( I => n3697, ZN => n4225);
   U13078 : NAND3_X1 port map( A1 => n6839, A2 => n12975, A3 => n19942, ZN => 
                           n24088);
   U13087 : XOR2_X1 port map( A1 => n22763, A2 => n9982, Z => n22713);
   U13091 : AOI22_X2 port map( A1 => n22186, A2 => n35652, B1 => n22188, B2 => 
                           n22187, ZN => n22763);
   U13092 : NOR2_X2 port map( A1 => n23162, A2 => n23163, ZN => n22869);
   U13096 : XOR2_X1 port map( A1 => n2370, A2 => n2372, Z => n11573);
   U13099 : NOR2_X2 port map( A1 => n39264, A2 => n13197, ZN => n13196);
   U13102 : NOR2_X2 port map( A1 => n5140, A2 => n37672, ZN => n6756);
   U13103 : OAI21_X2 port map( A1 => n1054, A2 => n29859, B => n11898, ZN => 
                           n11897);
   U13104 : XOR2_X1 port map( A1 => n37673, A2 => n22457, Z => n19002);
   U13107 : XOR2_X1 port map( A1 => n36641, A2 => n1656, Z => n37673);
   U13111 : BUF_X2 port map( I => n23149, Z => n37674);
   U13112 : XOR2_X1 port map( A1 => n37675, A2 => n9994, Z => n10959);
   U13113 : XOR2_X1 port map( A1 => n39520, A2 => n29098, Z => n37675);
   U13117 : XOR2_X1 port map( A1 => n437, A2 => n32959, Z => n35260);
   U13122 : XOR2_X1 port map( A1 => n19074, A2 => n19073, Z => n32959);
   U13126 : XOR2_X1 port map( A1 => n37676, A2 => n35969, Z => n30736);
   U13127 : XOR2_X1 port map( A1 => n16523, A2 => n23961, Z => n37676);
   U13128 : NAND2_X1 port map( A1 => n28626, A2 => n7914, ZN => n18125);
   U13135 : NAND2_X2 port map( A1 => n38065, A2 => n32681, ZN => n28626);
   U13137 : INV_X4 port map( I => n3642, ZN => n7258);
   U13143 : NAND2_X2 port map( A1 => n14300, A2 => n34297, ZN => n3642);
   U13144 : NAND2_X2 port map( A1 => n15896, A2 => n37677, ZN => n18743);
   U13150 : AOI22_X2 port map( A1 => n9423, A2 => n18870, B1 => n17346, B2 => 
                           n8155, ZN => n37677);
   U13153 : NOR2_X2 port map( A1 => n37589, A2 => n4473, ZN => n22683);
   U13154 : XOR2_X1 port map( A1 => n28990, A2 => n9787, Z => n9786);
   U13159 : XOR2_X1 port map( A1 => n10080, A2 => n10079, Z => n28990);
   U13160 : INV_X2 port map( I => n7703, ZN => n37678);
   U13161 : OR2_X1 port map( A1 => n13359, A2 => n37678, Z => n9466);
   U13162 : NAND2_X2 port map( A1 => n37679, A2 => n38010, ZN => n13458);
   U13164 : OAI21_X2 port map( A1 => n21223, A2 => n28249, B => n28115, ZN => 
                           n37679);
   U13165 : OAI21_X1 port map( A1 => n12189, A2 => n10677, B => n6648, ZN => 
                           n10177);
   U13167 : XOR2_X1 port map( A1 => n12441, A2 => n19096, Z => n24560);
   U13168 : XOR2_X1 port map( A1 => n37680, A2 => n19342, Z => n11627);
   U13170 : XOR2_X1 port map( A1 => n7118, A2 => n7119, Z => n37680);
   U13171 : XOR2_X1 port map( A1 => n8670, A2 => n33851, Z => n13099);
   U13174 : XOR2_X1 port map( A1 => n37681, A2 => n15046, Z => Ciphertext(69));
   U13176 : NOR3_X1 port map( A1 => n39340, A2 => n29569, A3 => n37145, ZN => 
                           n37681);
   U13180 : XOR2_X1 port map( A1 => n6435, A2 => n34492, Z => n28040);
   U13182 : NAND2_X2 port map( A1 => n14788, A2 => n31717, ZN => n5457);
   U13186 : OAI22_X2 port map( A1 => n18616, A2 => n15062, B1 => n38320, B2 => 
                           n38319, ZN => n14788);
   U13187 : NAND2_X2 port map( A1 => n18166, A2 => n22408, ZN => n7644);
   U13195 : XOR2_X1 port map( A1 => n37682, A2 => n29169, Z => n16371);
   U13199 : XOR2_X1 port map( A1 => n38058, A2 => n29038, Z => n37682);
   U13202 : XOR2_X1 port map( A1 => n26302, A2 => n26303, Z => n38188);
   U13203 : XOR2_X1 port map( A1 => n26449, A2 => n26301, Z => n26302);
   U13204 : BUF_X2 port map( I => n7660, Z => n37683);
   U13211 : NAND3_X2 port map( A1 => n5775, A2 => n5774, A3 => n5771, ZN => 
                           n27537);
   U13212 : OAI22_X2 port map( A1 => n13275, A2 => n2254, B1 => n38492, B2 => 
                           n2253, ZN => n16048);
   U13216 : INV_X2 port map( I => n7500, ZN => n14473);
   U13222 : NAND2_X2 port map( A1 => n12290, A2 => n26688, ZN => n26982);
   U13226 : OAI21_X2 port map( A1 => n37684, A2 => n24862, B => n524, ZN => 
                           n15001);
   U13229 : NAND2_X2 port map( A1 => n37685, A2 => n8217, ZN => n8475);
   U13233 : NAND2_X1 port map( A1 => n31077, A2 => n8216, ZN => n37685);
   U13235 : XOR2_X1 port map( A1 => n37686, A2 => n19808, Z => Ciphertext(109))
                           ;
   U13237 : OAI22_X1 port map( A1 => n39062, A2 => n3612, B1 => n3611, B2 => 
                           n29813, ZN => n37686);
   U13239 : BUF_X2 port map( I => n24589, Z => n37687);
   U13249 : XOR2_X1 port map( A1 => n39163, A2 => n38175, Z => n13074);
   U13256 : INV_X4 port map( I => n24590, ZN => n24717);
   U13258 : NAND2_X2 port map( A1 => n16882, A2 => n16881, ZN => n24590);
   U13260 : NOR2_X2 port map( A1 => n37688, A2 => n19278, ZN => n20657);
   U13261 : NAND2_X2 port map( A1 => n19942, A2 => n24221, ZN => n20119);
   U13264 : NOR2_X2 port map( A1 => n4686, A2 => n6891, ZN => n34658);
   U13271 : NOR2_X2 port map( A1 => n14377, A2 => n19179, ZN => n4686);
   U13272 : NAND2_X2 port map( A1 => n38141, A2 => n2792, ZN => n29800);
   U13277 : AOI22_X2 port map( A1 => n6649, A2 => n19393, B1 => n28960, B2 => 
                           n972, ZN => n15189);
   U13278 : XOR2_X1 port map( A1 => n30776, A2 => n37689, Z => n26665);
   U13280 : XOR2_X1 port map( A1 => n26375, A2 => n26166, Z => n37689);
   U13282 : XNOR2_X1 port map( A1 => n25310, A2 => n6996, ZN => n37968);
   U13284 : NOR2_X1 port map( A1 => n32111, A2 => n8784, ZN => n31079);
   U13285 : AOI21_X2 port map( A1 => n15767, A2 => n31133, B => n37690, ZN => 
                           n16525);
   U13286 : OAI21_X2 port map( A1 => n31626, A2 => n31133, B => n25822, ZN => 
                           n37690);
   U13300 : NAND2_X2 port map( A1 => n17616, A2 => n7585, ZN => n27395);
   U13304 : NAND3_X1 port map( A1 => n19362, A2 => n29517, A3 => n18384, ZN => 
                           n29521);
   U13307 : XOR2_X1 port map( A1 => n10611, A2 => n18428, Z => n32126);
   U13310 : OR2_X1 port map( A1 => n27624, A2 => n31121, Z => n18131);
   U13311 : NAND2_X2 port map( A1 => n17538, A2 => n5405, ZN => n32851);
   U13316 : OAI22_X2 port map( A1 => n6606, A2 => n26932, B1 => n4411, B2 => 
                           n5274, ZN => n17538);
   U13317 : XOR2_X1 port map( A1 => n23737, A2 => n37691, Z => n34933);
   U13318 : INV_X2 port map( I => n23709, ZN => n37691);
   U13323 : XOR2_X1 port map( A1 => n13617, A2 => n14289, Z => n23709);
   U13329 : OR2_X1 port map( A1 => n18790, A2 => n10810, Z => n24371);
   U13331 : NAND2_X2 port map( A1 => n37692, A2 => n23539, ZN => n5181);
   U13334 : OAI22_X2 port map( A1 => n23537, A2 => n31332, B1 => n23538, B2 => 
                           n12289, ZN => n37692);
   U13338 : NAND2_X2 port map( A1 => n37693, A2 => n35005, ZN => n28621);
   U13342 : OR2_X1 port map( A1 => n28232, A2 => n876, Z => n37693);
   U13345 : BUF_X4 port map( I => n5554, Z => n36911);
   U13346 : CLKBUF_X4 port map( I => n11569, Z => n6747);
   U13349 : XOR2_X1 port map( A1 => n7125, A2 => n7128, Z => n32010);
   U13352 : NAND2_X2 port map( A1 => n37694, A2 => n39128, ZN => n6355);
   U13353 : NOR2_X1 port map( A1 => n34028, A2 => n36052, ZN => n36004);
   U13354 : NOR2_X2 port map( A1 => n23476, A2 => n21293, ZN => n35917);
   U13359 : NAND2_X2 port map( A1 => n15176, A2 => n38600, ZN => n23476);
   U13361 : NAND3_X2 port map( A1 => n4857, A2 => n37897, A3 => n37695, ZN => 
                           n9108);
   U13362 : NAND2_X1 port map( A1 => n11490, A2 => n12537, ZN => n37695);
   U13364 : NAND2_X2 port map( A1 => n446, A2 => n38953, ZN => n25988);
   U13369 : NOR2_X2 port map( A1 => n36720, A2 => n23505, ZN => n7885);
   U13372 : NAND2_X2 port map( A1 => n37696, A2 => n8263, ZN => n35795);
   U13373 : INV_X2 port map( I => n37697, ZN => n19990);
   U13374 : XNOR2_X1 port map( A1 => n8937, A2 => n38000, ZN => n37697);
   U13376 : NAND2_X2 port map( A1 => n19175, A2 => n38101, ZN => n31899);
   U13377 : BUF_X2 port map( I => n18209, Z => n6691);
   U13379 : AOI22_X2 port map( A1 => n35048, A2 => n35049, B1 => n24743, B2 => 
                           n24744, ZN => n3111);
   U13380 : NOR2_X2 port map( A1 => n16999, A2 => n39317, ZN => n24744);
   U13385 : NOR2_X2 port map( A1 => n14993, A2 => n23597, ZN => n23680);
   U13386 : NAND2_X2 port map( A1 => n12373, A2 => n26639, ZN => n3992);
   U13391 : NAND2_X2 port map( A1 => n36726, A2 => n37698, ZN => n20418);
   U13394 : NAND3_X2 port map( A1 => n23061, A2 => n18637, A3 => n20518, ZN => 
                           n37698);
   U13395 : BUF_X4 port map( I => n23142, Z => n37984);
   U13396 : NAND2_X2 port map( A1 => n3077, A2 => n3561, ZN => n33609);
   U13401 : NAND2_X2 port map( A1 => n8766, A2 => n37948, ZN => n3077);
   U13404 : NOR2_X2 port map( A1 => n10474, A2 => n35956, ZN => n10473);
   U13412 : BUF_X2 port map( I => n19152, Z => n37699);
   U13417 : OAI21_X2 port map( A1 => n34000, A2 => n1962, B => n37700, ZN => 
                           n39736);
   U13421 : AOI21_X2 port map( A1 => n1962, A2 => n20673, B => n29781, ZN => 
                           n37700);
   U13423 : XOR2_X1 port map( A1 => n39760, A2 => n33672, Z => n23781);
   U13424 : INV_X4 port map( I => n8287, ZN => n1385);
   U13425 : OR2_X1 port map( A1 => n19713, A2 => n37016, Z => n7830);
   U13427 : BUF_X2 port map( I => n23714, Z => n37701);
   U13442 : XOR2_X1 port map( A1 => n33041, A2 => n1184, Z => n2032);
   U13443 : XOR2_X1 port map( A1 => n12534, A2 => n19862, Z => n25046);
   U13446 : NAND3_X2 port map( A1 => n38331, A2 => n24534, A3 => n37931, ZN => 
                           n19862);
   U13450 : NOR2_X1 port map( A1 => n37724, A2 => n10813, ZN => n37988);
   U13455 : INV_X1 port map( I => n14742, ZN => n38335);
   U13457 : INV_X1 port map( I => n29009, ZN => n37729);
   U13460 : XOR2_X1 port map( A1 => n22752, A2 => n22581, Z => n5233);
   U13462 : XNOR2_X1 port map( A1 => n5849, A2 => n5851, ZN => n38445);
   U13464 : XOR2_X1 port map( A1 => n14285, A2 => n14533, Z => n5851);
   U13466 : NOR2_X2 port map( A1 => n38695, A2 => n37702, ZN => n32136);
   U13468 : OAI22_X2 port map( A1 => n4702, A2 => n9101, B1 => n16902, B2 => 
                           n1035, ZN => n37702);
   U13470 : XOR2_X1 port map( A1 => n11695, A2 => n28997, Z => n29294);
   U13471 : NAND2_X2 port map( A1 => n39104, A2 => n13784, ZN => n28997);
   U13476 : OAI21_X1 port map( A1 => n26819, A2 => n7195, B => n30859, ZN => 
                           n26283);
   U13478 : NAND2_X2 port map( A1 => n37705, A2 => n23305, ZN => n18849);
   U13479 : XOR2_X1 port map( A1 => n11161, A2 => n39719, Z => n36064);
   U13481 : NAND2_X2 port map( A1 => n37706, A2 => n19460, ZN => n32646);
   U13484 : NAND2_X1 port map( A1 => n30615, A2 => n30613, ZN => n37706);
   U13486 : XOR2_X1 port map( A1 => n27679, A2 => n27633, Z => n27765);
   U13489 : NAND2_X2 port map( A1 => n27038, A2 => n18861, ZN => n27679);
   U13490 : XOR2_X1 port map( A1 => n16085, A2 => n27726, Z => n8563);
   U13492 : XOR2_X1 port map( A1 => n12556, A2 => n4885, Z => n27726);
   U13494 : BUF_X4 port map( I => n2046, Z => n1989);
   U13499 : XOR2_X1 port map( A1 => n7942, A2 => n37707, Z => n3476);
   U13501 : XOR2_X1 port map( A1 => n3478, A2 => n359, Z => n37707);
   U13502 : NAND2_X2 port map( A1 => n15946, A2 => n39521, ZN => n30913);
   U13508 : NOR2_X1 port map( A1 => n29810, A2 => n29803, ZN => n3614);
   U13509 : NAND2_X2 port map( A1 => n28923, A2 => n28924, ZN => n29810);
   U13511 : NAND2_X2 port map( A1 => n37708, A2 => n38640, ZN => n17756);
   U13515 : OAI21_X2 port map( A1 => n37803, A2 => n31270, B => n6849, ZN => 
                           n30684);
   U13519 : NAND2_X2 port map( A1 => n37709, A2 => n38484, ZN => n22376);
   U13526 : NAND2_X1 port map( A1 => n36090, A2 => n7852, ZN => n8580);
   U13536 : NAND2_X1 port map( A1 => n10004, A2 => n1257, ZN => n37712);
   U13549 : INV_X1 port map( I => n18249, ZN => n37713);
   U13551 : XOR2_X1 port map( A1 => n14264, A2 => n13245, Z => n10129);
   U13552 : INV_X1 port map( I => n38785, ZN => n38784);
   U13553 : XOR2_X1 port map( A1 => n28842, A2 => n8371, Z => n1914);
   U13558 : XOR2_X1 port map( A1 => n29147, A2 => n1915, Z => n8371);
   U13559 : NAND2_X2 port map( A1 => n37714, A2 => n2342, ZN => n2634);
   U13561 : NOR2_X2 port map( A1 => n15898, A2 => n33500, ZN => n37714);
   U13565 : NAND2_X2 port map( A1 => n9508, A2 => n19508, ZN => n33855);
   U13571 : XOR2_X1 port map( A1 => n37715, A2 => n23921, Z => n11699);
   U13572 : XOR2_X1 port map( A1 => n8904, A2 => n39177, Z => n37715);
   U13574 : XOR2_X1 port map( A1 => n4123, A2 => n4210, Z => n4209);
   U13576 : NAND2_X2 port map( A1 => n30877, A2 => n30354, ZN => n4210);
   U13577 : NAND2_X2 port map( A1 => n33461, A2 => n5619, ZN => n31612);
   U13579 : AND2_X2 port map( A1 => n25639, A2 => n25669, Z => n3101);
   U13580 : XOR2_X1 port map( A1 => n39219, A2 => n29294, Z => n15091);
   U13591 : XOR2_X1 port map( A1 => n2126, A2 => n5246, Z => n7582);
   U13595 : NAND2_X2 port map( A1 => n36795, A2 => n3909, ZN => n2126);
   U13600 : AOI21_X1 port map( A1 => n14337, A2 => n29722, B => n29719, ZN => 
                           n29705);
   U13604 : AOI22_X2 port map( A1 => n32192, A2 => n4448, B1 => n29703, B2 => 
                           n4447, ZN => n29722);
   U13607 : INV_X1 port map( I => n32228, ZN => n1655);
   U13608 : AND2_X1 port map( A1 => n32228, A2 => n19840, Z => n32202);
   U13609 : OAI22_X2 port map( A1 => n2772, A2 => n8942, B1 => n5628, B2 => 
                           n8707, ZN => n31325);
   U13613 : AOI22_X2 port map( A1 => n29430, A2 => n37716, B1 => n35517, B2 => 
                           n34194, ZN => n18502);
   U13617 : NAND2_X1 port map( A1 => n15089, A2 => n29497, ZN => n37716);
   U13623 : XOR2_X1 port map( A1 => n37718, A2 => n38875, Z => n9791);
   U13625 : XOR2_X1 port map( A1 => n11730, A2 => n39515, Z => n37718);
   U13632 : INV_X2 port map( I => n10216, ZN => n2182);
   U13633 : NAND3_X2 port map( A1 => n39588, A2 => n13077, A3 => n13078, ZN => 
                           n10216);
   U13634 : INV_X2 port map( I => n33949, ZN => n36162);
   U13637 : OAI21_X2 port map( A1 => n35788, A2 => n35789, B => n19827, ZN => 
                           n37719);
   U13641 : XOR2_X1 port map( A1 => n4077, A2 => n37720, Z => n4081);
   U13643 : XOR2_X1 port map( A1 => n30913, A2 => n1238, Z => n37720);
   U13651 : XOR2_X1 port map( A1 => n37721, A2 => n12972, Z => n10872);
   U13655 : NAND2_X2 port map( A1 => n36966, A2 => n31446, ZN => n12972);
   U13659 : NAND2_X2 port map( A1 => n29781, A2 => n29777, ZN => n39154);
   U13660 : NAND2_X2 port map( A1 => n39154, A2 => n29779, ZN => n38574);
   U13662 : XOR2_X1 port map( A1 => n37723, A2 => n37722, Z => n12334);
   U13663 : XOR2_X1 port map( A1 => n4815, A2 => n27641, Z => n37722);
   U13666 : XOR2_X1 port map( A1 => n27642, A2 => n20641, Z => n37723);
   U13667 : OAI22_X2 port map( A1 => n17502, A2 => n7915, B1 => n32747, B2 => 
                           n32520, ZN => n10458);
   U13672 : XOR2_X1 port map( A1 => n29037, A2 => n37725, Z => n38136);
   U13674 : XOR2_X1 port map( A1 => n37726, A2 => n14956, Z => n37725);
   U13679 : AOI21_X2 port map( A1 => n36701, A2 => n36011, B => n1695, ZN => 
                           n37763);
   U13682 : XNOR2_X1 port map( A1 => n33756, A2 => n32646, ZN => n514);
   U13683 : NAND2_X2 port map( A1 => n29010, A2 => n37728, ZN => n37727);
   U13684 : INV_X2 port map( I => n20525, ZN => n37728);
   U13687 : BUF_X4 port map( I => n25319, Z => n39491);
   U13688 : INV_X2 port map( I => n37731, ZN => n21768);
   U13691 : XNOR2_X1 port map( A1 => Key(161), A2 => Plaintext(161), ZN => 
                           n37731);
   U13694 : OAI21_X2 port map( A1 => n23302, A2 => n32017, B => n23489, ZN => 
                           n529);
   U13699 : BUF_X2 port map( I => n30186, Z => n37734);
   U13702 : NAND2_X2 port map( A1 => n34205, A2 => n37735, ZN => n30358);
   U13706 : OAI21_X2 port map( A1 => n37173, A2 => n37736, B => n36133, ZN => 
                           n36460);
   U13708 : NOR2_X2 port map( A1 => n36162, A2 => n3985, ZN => n37736);
   U13709 : INV_X4 port map( I => n36385, ZN => n1271);
   U13712 : NAND2_X2 port map( A1 => n13706, A2 => n13709, ZN => n36385);
   U13713 : XOR2_X1 port map( A1 => n27723, A2 => n27635, Z => n7022);
   U13715 : XOR2_X1 port map( A1 => n27829, A2 => n27595, Z => n27723);
   U13717 : NAND3_X2 port map( A1 => n38960, A2 => n19584, A3 => n24443, ZN => 
                           n24313);
   U13731 : XOR2_X1 port map( A1 => n37738, A2 => n23789, Z => n23926);
   U13737 : NAND2_X2 port map( A1 => n32025, A2 => n23093, ZN => n23568);
   U13739 : NOR2_X2 port map( A1 => n12050, A2 => n37739, ZN => n24668);
   U13756 : AND2_X1 port map( A1 => n13040, A2 => n5954, Z => n37739);
   U13760 : NOR2_X2 port map( A1 => n31144, A2 => n37740, ZN => n31143);
   U13761 : NOR3_X2 port map( A1 => n1570, A2 => n24750, A3 => n38182, ZN => 
                           n37740);
   U13763 : XOR2_X1 port map( A1 => n24039, A2 => n24028, Z => n36760);
   U13765 : XOR2_X1 port map( A1 => n17925, A2 => n35235, Z => n24028);
   U13775 : AOI22_X2 port map( A1 => n39260, A2 => n37102, B1 => n38138, B2 => 
                           n10340, ZN => n35750);
   U13777 : AOI21_X2 port map( A1 => n23360, A2 => n23359, B => n31594, ZN => 
                           n38650);
   U13778 : INV_X2 port map( I => n281, ZN => n28143);
   U13779 : XOR2_X1 port map( A1 => n11856, A2 => n37741, Z => n16699);
   U13780 : XOR2_X1 port map( A1 => n25251, A2 => n10215, Z => n37741);
   U13782 : NAND2_X2 port map( A1 => n9499, A2 => n37742, ZN => n10225);
   U13783 : XOR2_X1 port map( A1 => n29824, A2 => n28852, Z => n13381);
   U13786 : NAND2_X2 port map( A1 => n35574, A2 => n12607, ZN => n29824);
   U13789 : NAND3_X1 port map( A1 => n28671, A2 => n28674, A3 => n18883, ZN => 
                           n15959);
   U13791 : XOR2_X1 port map( A1 => n20095, A2 => n15545, Z => n38081);
   U13793 : NOR2_X1 port map( A1 => n35368, A2 => n13620, ZN => n13618);
   U13798 : XOR2_X1 port map( A1 => n27759, A2 => n27760, Z => n36863);
   U13801 : XOR2_X1 port map( A1 => n38937, A2 => n17349, Z => n27759);
   U13804 : OR2_X1 port map( A1 => n26724, A2 => n26832, Z => n26679);
   U13805 : OAI21_X2 port map( A1 => n21587, A2 => n14499, B => n8597, ZN => 
                           n21413);
   U13808 : NOR2_X2 port map( A1 => n20979, A2 => n29642, ZN => n37743);
   U13809 : XOR2_X1 port map( A1 => n37744, A2 => n8502, Z => n39027);
   U13812 : XOR2_X1 port map( A1 => n33812, A2 => n38495, Z => n37744);
   U13814 : INV_X2 port map( I => n32134, ZN => n6592);
   U13821 : XOR2_X1 port map( A1 => n13920, A2 => n6595, Z => n32134);
   U13822 : OAI22_X2 port map( A1 => n19590, A2 => n16200, B1 => n1518, B2 => 
                           n32469, ZN => n37745);
   U13827 : XOR2_X1 port map( A1 => n29098, A2 => n28916, Z => n28878);
   U13829 : XOR2_X1 port map( A1 => n18305, A2 => n15745, Z => n29098);
   U13832 : XOR2_X1 port map( A1 => n27459, A2 => n27715, Z => n14359);
   U13837 : XOR2_X1 port map( A1 => n31551, A2 => n34963, Z => n27459);
   U13838 : XOR2_X1 port map( A1 => n23878, A2 => n20877, Z => n2596);
   U13840 : XOR2_X1 port map( A1 => n1617, A2 => n24079, Z => n23878);
   U13844 : NAND2_X2 port map( A1 => n31640, A2 => n5787, ZN => n10764);
   U13847 : XOR2_X1 port map( A1 => n26558, A2 => n3152, Z => n3151);
   U13848 : NAND2_X2 port map( A1 => n37747, A2 => n35670, ZN => n31937);
   U13850 : NAND2_X2 port map( A1 => n34504, A2 => n1602, ZN => n37747);
   U13855 : XOR2_X1 port map( A1 => n23975, A2 => n23742, Z => n11119);
   U13859 : OAI21_X2 port map( A1 => n19246, A2 => n39045, B => n37749, ZN => 
                           n17931);
   U13860 : NOR2_X2 port map( A1 => n37750, A2 => n15452, ZN => n1627);
   U13861 : XOR2_X1 port map( A1 => n25144, A2 => n25318, Z => n32532);
   U13864 : NAND3_X1 port map( A1 => n38012, A2 => n5038, A3 => n39350, ZN => 
                           n20191);
   U13865 : XNOR2_X1 port map( A1 => n22470, A2 => n22567, ZN => n37869);
   U13878 : AOI22_X2 port map( A1 => n20013, A2 => n24664, B1 => n37751, B2 => 
                           n2340, ZN => n16051);
   U13879 : NOR2_X2 port map( A1 => n35578, A2 => n38523, ZN => n37751);
   U13883 : XOR2_X1 port map( A1 => n16900, A2 => n33271, Z => n10611);
   U13884 : NAND2_X2 port map( A1 => n7396, A2 => n4729, ZN => n16900);
   U13885 : INV_X1 port map( I => n20010, ZN => n37753);
   U13886 : NOR3_X2 port map( A1 => n36662, A2 => n3411, A3 => n3410, ZN => 
                           n3409);
   U13891 : XOR2_X1 port map( A1 => n7553, A2 => n26570, Z => n18738);
   U13894 : XOR2_X1 port map( A1 => n26571, A2 => n6177, Z => n7553);
   U13895 : AOI22_X2 port map( A1 => n7479, A2 => n10702, B1 => n19544, B2 => 
                           n11677, ZN => n3463);
   U13905 : NOR2_X2 port map( A1 => n34264, A2 => n4215, ZN => n26029);
   U13906 : XOR2_X1 port map( A1 => n11050, A2 => n37755, Z => n38026);
   U13910 : XOR2_X1 port map( A1 => n37889, A2 => n35257, Z => n37755);
   U13919 : XOR2_X1 port map( A1 => n7981, A2 => n37756, Z => n23682);
   U13920 : XOR2_X1 port map( A1 => n24058, A2 => n17398, Z => n37756);
   U13928 : INV_X2 port map( I => n4599, ZN => n33561);
   U13930 : OR2_X1 port map( A1 => n1265, A2 => n24737, Z => n38738);
   U13937 : OAI21_X2 port map( A1 => n2581, A2 => n25466, B => n35271, ZN => 
                           n36499);
   U13948 : NOR2_X2 port map( A1 => n220, A2 => n591, ZN => n2581);
   U13949 : BUF_X2 port map( I => n35534, Z => n37757);
   U13953 : OAI22_X2 port map( A1 => n33325, A2 => n28457, B1 => n1823, B2 => 
                           n28458, ZN => n37759);
   U13954 : NAND3_X1 port map( A1 => n25999, A2 => n31362, A3 => n35138, ZN => 
                           n2493);
   U13958 : OAI21_X2 port map( A1 => n8698, A2 => n35749, B => n14041, ZN => 
                           n8697);
   U13959 : NAND2_X1 port map( A1 => n34069, A2 => n28276, ZN => n35844);
   U13964 : OR2_X1 port map( A1 => n2654, A2 => n36371, Z => n30893);
   U13965 : OAI21_X2 port map( A1 => n8154, A2 => n17194, B => n19222, ZN => 
                           n9367);
   U13967 : BUF_X4 port map( I => n39477, Z => n38519);
   U13969 : XOR2_X1 port map( A1 => n37761, A2 => n39559, Z => Ciphertext(46));
   U13971 : AOI22_X1 port map( A1 => n15132, A2 => n15131, B1 => n15128, B2 => 
                           n15127, ZN => n37761);
   U13975 : XOR2_X1 port map( A1 => n23891, A2 => n23892, Z => n23897);
   U13977 : XOR2_X1 port map( A1 => n24061, A2 => n23808, Z => n23891);
   U13978 : NOR2_X2 port map( A1 => n11247, A2 => n25759, ZN => n38584);
   U13989 : NAND2_X2 port map( A1 => n37762, A2 => n25443, ZN => n11734);
   U13996 : NAND3_X2 port map( A1 => n37949, A2 => n30399, A3 => n9305, ZN => 
                           n37762);
   U13997 : INV_X1 port map( I => n37763, ZN => n11987);
   U13999 : XOR2_X1 port map( A1 => n37765, A2 => n37764, Z => n18220);
   U14000 : XOR2_X1 port map( A1 => n487, A2 => n7337, Z => n37765);
   U14008 : XOR2_X1 port map( A1 => n22527, A2 => n1368, Z => n39693);
   U14012 : OAI22_X2 port map( A1 => n7105, A2 => n20376, B1 => n31953, B2 => 
                           n7104, ZN => n22527);
   U14018 : XOR2_X1 port map( A1 => n17606, A2 => n13935, Z => n24955);
   U14022 : INV_X2 port map( I => n38385, ZN => n38905);
   U14032 : XOR2_X1 port map( A1 => n3917, A2 => n38385, Z => n3773);
   U14062 : NOR2_X2 port map( A1 => n35018, A2 => n31816, ZN => n38385);
   U14072 : XOR2_X1 port map( A1 => n26254, A2 => n15010, Z => n21085);
   U14074 : XOR2_X1 port map( A1 => n8634, A2 => n23807, Z => n30891);
   U14075 : XOR2_X1 port map( A1 => n24030, A2 => n238, Z => n8634);
   U14078 : AOI22_X2 port map( A1 => n9672, A2 => n23522, B1 => n36878, B2 => 
                           n9190, ZN => n35885);
   U14079 : XOR2_X1 port map( A1 => n37767, A2 => n4270, Z => n3585);
   U14083 : XOR2_X1 port map( A1 => n3475, A2 => n22711, Z => n37767);
   U14085 : INV_X4 port map( I => n2616, ZN => n16841);
   U14097 : AOI21_X2 port map( A1 => n37142, A2 => n21472, B => n37768, ZN => 
                           n22250);
   U14101 : AOI22_X1 port map( A1 => n21617, A2 => n18293, B1 => n19372, B2 => 
                           n917, ZN => n37768);
   U14106 : XOR2_X1 port map( A1 => n26518, A2 => n31293, Z => n26221);
   U14108 : NAND2_X2 port map( A1 => n16952, A2 => n25914, ZN => n26518);
   U14111 : XOR2_X1 port map( A1 => n11602, A2 => n34911, Z => n15566);
   U14116 : INV_X2 port map( I => n37769, ZN => n38166);
   U14117 : NAND3_X2 port map( A1 => n29597, A2 => n29596, A3 => n29595, ZN => 
                           n37769);
   U14126 : INV_X1 port map( I => n19997, ZN => n37770);
   U14127 : NOR2_X2 port map( A1 => n38368, A2 => n5385, ZN => n34632);
   U14129 : INV_X4 port map( I => n29452, ZN => n14151);
   U14131 : XOR2_X1 port map( A1 => n29041, A2 => n28966, Z => n29090);
   U14132 : XOR2_X1 port map( A1 => n31599, A2 => n23965, Z => n8400);
   U14133 : AOI21_X2 port map( A1 => n23356, A2 => n39534, B => n33696, ZN => 
                           n31599);
   U14134 : XOR2_X1 port map( A1 => n17703, A2 => n14603, Z => n8888);
   U14135 : XOR2_X1 port map( A1 => n6435, A2 => n37951, Z => n17703);
   U14140 : NAND2_X2 port map( A1 => n5209, A2 => n10373, ZN => n7328);
   U14147 : NAND2_X2 port map( A1 => n35248, A2 => n36105, ZN => n12944);
   U14148 : NOR2_X2 port map( A1 => n12406, A2 => n14397, ZN => n27870);
   U14153 : NAND2_X2 port map( A1 => n7751, A2 => n19168, ZN => n33747);
   U14161 : XOR2_X1 port map( A1 => n35222, A2 => n18362, Z => n3140);
   U14166 : BUF_X2 port map( I => n14260, Z => n37833);
   U14167 : XOR2_X1 port map( A1 => n18808, A2 => n37772, Z => n36962);
   U14169 : XOR2_X1 port map( A1 => n31293, A2 => n39662, Z => n37772);
   U14171 : BUF_X2 port map( I => n10764, Z => n32520);
   U14172 : XOR2_X1 port map( A1 => n16566, A2 => n26508, Z => n4572);
   U14176 : NAND2_X2 port map( A1 => n37773, A2 => n29771, ZN => n15867);
   U14181 : NAND2_X1 port map( A1 => n20895, A2 => n20894, ZN => n37773);
   U14190 : AND2_X1 port map( A1 => n11970, A2 => n37774, Z => n11969);
   U14193 : XOR2_X1 port map( A1 => n37995, A2 => n26510, Z => n33750);
   U14194 : NAND2_X2 port map( A1 => n25918, A2 => n25917, ZN => n26510);
   U14197 : XOR2_X1 port map( A1 => n24023, A2 => n24065, Z => n17563);
   U14201 : NOR2_X2 port map( A1 => n37777, A2 => n37776, ZN => n34639);
   U14202 : INV_X2 port map( I => n39423, ZN => n37776);
   U14204 : NOR2_X2 port map( A1 => n37976, A2 => n11797, ZN => n16057);
   U14205 : XOR2_X1 port map( A1 => n25315, A2 => n17606, Z => n2618);
   U14208 : XOR2_X1 port map( A1 => n25296, A2 => n25196, Z => n25315);
   U14210 : NOR2_X2 port map( A1 => n6747, A2 => n1545, ZN => n25666);
   U14212 : NAND2_X1 port map( A1 => n37539, A2 => n39196, ZN => n6186);
   U14213 : XOR2_X1 port map( A1 => n37778, A2 => n4564, Z => n16445);
   U14214 : XOR2_X1 port map( A1 => n21257, A2 => n4563, Z => n37778);
   U14215 : XOR2_X1 port map( A1 => n14297, A2 => n12101, Z => n30842);
   U14218 : XOR2_X1 port map( A1 => n22439, A2 => n1668, Z => n14297);
   U14219 : AOI21_X2 port map( A1 => n6184, A2 => n6183, B => n6189, ZN => 
                           n6185);
   U14221 : NAND2_X2 port map( A1 => n31200, A2 => n37779, ZN => n23976);
   U14222 : AND2_X1 port map( A1 => n9694, A2 => n4553, Z => n19898);
   U14226 : XOR2_X1 port map( A1 => n9274, A2 => n2815, Z => n18383);
   U14230 : OAI21_X2 port map( A1 => n29775, A2 => n18222, B => n37780, ZN => 
                           n29797);
   U14232 : NOR2_X2 port map( A1 => n18221, A2 => n17912, ZN => n37780);
   U14235 : NAND2_X1 port map( A1 => n28017, A2 => n31494, ZN => n37785);
   U14236 : XOR2_X1 port map( A1 => n27718, A2 => n5394, Z => n37786);
   U14242 : XOR2_X1 port map( A1 => n404, A2 => n37787, Z => n20945);
   U14243 : XOR2_X1 port map( A1 => n29000, A2 => n37256, Z => n37787);
   U14249 : OAI21_X2 port map( A1 => n3742, A2 => n34249, B => n32256, ZN => 
                           n37788);
   U14250 : NAND2_X1 port map( A1 => n30465, A2 => n6747, ZN => n20440);
   U14252 : AOI21_X2 port map( A1 => n8752, A2 => n22401, B => n8750, ZN => 
                           n35824);
   U14253 : OAI21_X2 port map( A1 => n21497, A2 => n38878, B => n21309, ZN => 
                           n37789);
   U14254 : XOR2_X1 port map( A1 => n9576, A2 => n2055, Z => n19973);
   U14255 : NAND2_X2 port map( A1 => n5679, A2 => n5683, ZN => n2055);
   U14257 : XOR2_X1 port map( A1 => n37790, A2 => n33429, Z => n19170);
   U14262 : XOR2_X1 port map( A1 => n3787, A2 => n38440, Z => n37790);
   U14266 : NAND3_X2 port map( A1 => n7014, A2 => n7012, A3 => n7013, ZN => 
                           n35232);
   U14267 : NAND2_X2 port map( A1 => n38574, A2 => n481, ZN => n2560);
   U14274 : AOI22_X2 port map( A1 => n37792, A2 => n37791, B1 => n22368, B2 => 
                           n17319, ZN => n16528);
   U14279 : XOR2_X1 port map( A1 => n28888, A2 => n17325, Z => n39247);
   U14281 : INV_X2 port map( I => n8787, ZN => n28494);
   U14282 : NAND3_X2 port map( A1 => n28352, A2 => n12885, A3 => n28349, ZN => 
                           n8787);
   U14283 : NAND2_X1 port map( A1 => n35551, A2 => n19693, ZN => n35695);
   U14284 : NOR2_X1 port map( A1 => n20943, A2 => n20351, ZN => n37793);
   U14287 : XOR2_X1 port map( A1 => n26255, A2 => n5848, Z => n26417);
   U14291 : NAND2_X2 port map( A1 => n30967, A2 => n31630, ZN => n5241);
   U14293 : BUF_X2 port map( I => n2803, Z => n37795);
   U14294 : XOR2_X1 port map( A1 => n24061, A2 => n23762, Z => n23944);
   U14295 : OAI22_X2 port map( A1 => n17787, A2 => n14649, B1 => n17788, B2 => 
                           n38252, ZN => n24061);
   U14297 : XOR2_X1 port map( A1 => n27542, A2 => n13374, Z => n27654);
   U14298 : AOI22_X2 port map( A1 => n10356, A2 => n10357, B1 => n10358, B2 => 
                           n1474, ZN => n13374);
   U14299 : XOR2_X1 port map( A1 => n28878, A2 => n34773, Z => n18967);
   U14302 : AOI22_X2 port map( A1 => n15918, A2 => n4434, B1 => n27410, B2 => 
                           n15917, ZN => n4462);
   U14306 : NAND2_X1 port map( A1 => n1414, A2 => n38629, ZN => n28480);
   U14312 : NAND2_X2 port map( A1 => n20020, A2 => n28104, ZN => n38629);
   U14316 : AOI22_X2 port map( A1 => n24165, A2 => n39156, B1 => n1282, B2 => 
                           n23704, ZN => n24584);
   U14321 : NOR2_X1 port map( A1 => n6331, A2 => n20601, ZN => n23704);
   U14325 : XOR2_X1 port map( A1 => n2445, A2 => n39550, Z => n7500);
   U14326 : XOR2_X1 port map( A1 => n6987, A2 => n37796, Z => n15935);
   U14329 : XOR2_X1 port map( A1 => n1614, A2 => n13978, Z => n37796);
   U14331 : XOR2_X1 port map( A1 => n25173, A2 => n25172, Z => n36959);
   U14332 : XOR2_X1 port map( A1 => n25214, A2 => n8183, Z => n25173);
   U14335 : XOR2_X1 port map( A1 => n26399, A2 => n15595, Z => n13658);
   U14336 : XOR2_X1 port map( A1 => n26117, A2 => n31965, Z => n15595);
   U14341 : AND2_X1 port map( A1 => n15284, A2 => n39484, Z => n26694);
   U14355 : NAND2_X2 port map( A1 => n38232, A2 => n31406, ZN => n15284);
   U14356 : NAND2_X2 port map( A1 => n38805, A2 => n37797, ZN => n29439);
   U14358 : OAI21_X2 port map( A1 => n25347, A2 => n4013, B => n25346, ZN => 
                           n31115);
   U14359 : NAND2_X2 port map( A1 => n3337, A2 => n13861, ZN => n13860);
   U14365 : NOR2_X2 port map( A1 => n3784, A2 => n13855, ZN => n3337);
   U14373 : NAND2_X2 port map( A1 => n26928, A2 => n26927, ZN => n37798);
   U14374 : AOI21_X2 port map( A1 => n19993, A2 => n16790, B => n34000, ZN => 
                           n16845);
   U14378 : NAND3_X2 port map( A1 => n4931, A2 => n5702, A3 => n33972, ZN => 
                           n37982);
   U14379 : XOR2_X1 port map( A1 => n37799, A2 => n19890, Z => Ciphertext(43));
   U14387 : NAND3_X1 port map( A1 => n12340, A2 => n12339, A3 => n12321, ZN => 
                           n37799);
   U14390 : XOR2_X1 port map( A1 => n37800, A2 => n14715, Z => n25598);
   U14392 : XOR2_X1 port map( A1 => n720, A2 => n25002, Z => n37800);
   U14394 : OAI21_X1 port map( A1 => n4576, A2 => n23426, B => n32024, ZN => 
                           n37802);
   U14397 : XOR2_X1 port map( A1 => n27501, A2 => n12341, Z => n27760);
   U14400 : AOI22_X2 port map( A1 => n8268, A2 => n1625, B1 => n23531, B2 => 
                           n8269, ZN => n33462);
   U14403 : AND2_X1 port map( A1 => n25597, A2 => n1254, Z => n33407);
   U14408 : NAND2_X1 port map( A1 => n4613, A2 => n4342, ZN => n37805);
   U14410 : INV_X2 port map( I => n6691, ZN => n36724);
   U14413 : XOR2_X1 port map( A1 => n37806, A2 => n29974, Z => Ciphertext(135))
                           ;
   U14415 : NAND3_X2 port map( A1 => n32570, A2 => n7270, A3 => n7271, ZN => 
                           n37806);
   U14423 : XOR2_X1 port map( A1 => n29094, A2 => n29255, Z => n14981);
   U14424 : NAND3_X2 port map( A1 => n7752, A2 => n9269, A3 => n16970, ZN => 
                           n20094);
   U14426 : AND2_X1 port map( A1 => n4613, A2 => n22337, Z => n22102);
   U14428 : OAI21_X1 port map( A1 => n19442, A2 => n14000, B => n35197, ZN => 
                           n11421);
   U14430 : XOR2_X1 port map( A1 => n37807, A2 => n27844, Z => n38054);
   U14437 : XOR2_X1 port map( A1 => n15421, A2 => n27554, Z => n37807);
   U14441 : OR2_X1 port map( A1 => n23517, A2 => n39001, Z => n38536);
   U14445 : XOR2_X1 port map( A1 => n37808, A2 => n26201, Z => n26770);
   U14446 : XOR2_X1 port map( A1 => n32934, A2 => n26200, Z => n37808);
   U14450 : OR2_X1 port map( A1 => n24747, A2 => n24601, Z => n19999);
   U14453 : NAND2_X2 port map( A1 => n16196, A2 => n37983, ZN => n24747);
   U14454 : NOR2_X2 port map( A1 => n23201, A2 => n35576, ZN => n15200);
   U14455 : NAND2_X2 port map( A1 => n37810, A2 => n3437, ZN => n22196);
   U14458 : NAND2_X1 port map( A1 => n20844, A2 => n9316, ZN => n37810);
   U14459 : XOR2_X1 port map( A1 => n31445, A2 => n37811, Z => n10665);
   U14462 : XOR2_X1 port map( A1 => n25171, A2 => n16555, Z => n37811);
   U14463 : AOI21_X2 port map( A1 => n29202, A2 => n33488, B => n37813, ZN => 
                           n39829);
   U14464 : NOR2_X1 port map( A1 => n10779, A2 => n1436, ZN => n38764);
   U14465 : BUF_X2 port map( I => n36150, Z => n37815);
   U14466 : XOR2_X1 port map( A1 => n4305, A2 => n39725, Z => n37816);
   U14467 : OR2_X1 port map( A1 => n5886, A2 => n26048, Z => n8898);
   U14474 : INV_X2 port map( I => n29220, ZN => n13107);
   U14475 : NAND2_X2 port map( A1 => n32189, A2 => n38071, ZN => n29220);
   U14476 : NAND2_X2 port map( A1 => n16348, A2 => n16347, ZN => n19094);
   U14478 : NAND2_X2 port map( A1 => n17557, A2 => n2458, ZN => n16348);
   U14480 : AOI22_X2 port map( A1 => n9508, A2 => n5471, B1 => n18816, B2 => 
                           n5570, ZN => n3247);
   U14481 : XOR2_X1 port map( A1 => n3015, A2 => n25292, Z => n8003);
   U14483 : NOR2_X2 port map( A1 => n2905, A2 => n2903, ZN => n25292);
   U14487 : AND2_X1 port map( A1 => n11145, A2 => n14332, Z => n32536);
   U14488 : NAND3_X1 port map( A1 => n32783, A2 => n13714, A3 => n15597, ZN => 
                           n32235);
   U14491 : AND2_X1 port map( A1 => n2117, A2 => n32310, Z => n24314);
   U14494 : NOR2_X1 port map( A1 => n13005, A2 => n19249, ZN => n38995);
   U14500 : INV_X2 port map( I => n25860, ZN => n1520);
   U14501 : XOR2_X1 port map( A1 => n17399, A2 => n3126, Z => n3117);
   U14505 : XOR2_X1 port map( A1 => n29045, A2 => n30964, Z => n17399);
   U14508 : XOR2_X1 port map( A1 => n37817, A2 => n23913, Z => n31505);
   U14509 : XOR2_X1 port map( A1 => n10312, A2 => n1619, Z => n37817);
   U14512 : AOI21_X2 port map( A1 => n34608, A2 => n37818, B => n36314, ZN => 
                           n38318);
   U14515 : NAND2_X2 port map( A1 => n35745, A2 => n31433, ZN => n37818);
   U14516 : XOR2_X1 port map( A1 => n16296, A2 => n23939, Z => n8904);
   U14519 : NAND2_X2 port map( A1 => n39218, A2 => n23322, ZN => n16296);
   U14521 : OR2_X1 port map( A1 => n8395, A2 => n8604, Z => n8291);
   U14522 : OAI21_X1 port map( A1 => n38830, A2 => n20391, B => n22058, ZN => 
                           n16403);
   U14525 : XOR2_X1 port map( A1 => n34544, A2 => n27646, Z => n18474);
   U14526 : XOR2_X1 port map( A1 => n6960, A2 => n37820, Z => n36847);
   U14527 : XOR2_X1 port map( A1 => n26234, A2 => n17396, Z => n37820);
   U14529 : NAND3_X2 port map( A1 => n8491, A2 => n1042, A3 => n35684, ZN => 
                           n10437);
   U14536 : NAND2_X2 port map( A1 => n23255, A2 => n33702, ZN => n19536);
   U14537 : NAND2_X1 port map( A1 => n24371, A2 => n24370, ZN => n13070);
   U14538 : XOR2_X1 port map( A1 => n39804, A2 => n16898, Z => n14106);
   U14539 : NOR2_X2 port map( A1 => n21338, A2 => n19216, ZN => n39804);
   U14542 : XOR2_X1 port map( A1 => n8852, A2 => n31127, Z => n29153);
   U14544 : OAI21_X2 port map( A1 => n38127, A2 => n28759, B => n8449, ZN => 
                           n8852);
   U14545 : XOR2_X1 port map( A1 => n34998, A2 => n5703, Z => n35724);
   U14546 : XOR2_X1 port map( A1 => n37998, A2 => n39744, Z => n32556);
   U14547 : XOR2_X1 port map( A1 => n38585, A2 => n2712, Z => n30503);
   U14548 : XOR2_X1 port map( A1 => n6719, A2 => n14307, Z => n29038);
   U14549 : NAND2_X2 port map( A1 => n38077, A2 => n4005, ZN => n14307);
   U14550 : XNOR2_X1 port map( A1 => n1010, A2 => n5084, ZN => n26420);
   U14554 : NAND2_X2 port map( A1 => n8380, A2 => n8381, ZN => n5625);
   U14556 : NAND2_X2 port map( A1 => n8383, A2 => n8385, ZN => n8380);
   U14562 : NOR2_X2 port map( A1 => n37823, A2 => n37822, ZN => n17249);
   U14564 : INV_X1 port map( I => n5131, ZN => n37822);
   U14566 : INV_X2 port map( I => n21912, ZN => n37823);
   U14571 : NAND2_X2 port map( A1 => n37824, A2 => n15201, ZN => n8693);
   U14575 : OAI21_X2 port map( A1 => n15200, A2 => n15199, B => n22849, ZN => 
                           n37824);
   U14577 : XOR2_X1 port map( A1 => n37825, A2 => n19676, Z => Ciphertext(177))
                           ;
   U14579 : XOR2_X1 port map( A1 => n13917, A2 => n25267, Z => n14955);
   U14589 : OAI21_X2 port map( A1 => n36485, A2 => n24113, B => n24101, ZN => 
                           n13316);
   U14593 : OAI21_X2 port map( A1 => n16890, A2 => n2498, B => n692, ZN => 
                           n39164);
   U14594 : XOR2_X1 port map( A1 => n4929, A2 => n14953, Z => n11092);
   U14595 : INV_X2 port map( I => n38630, ZN => n35287);
   U14596 : NAND2_X2 port map( A1 => n37827, A2 => n37826, ZN => n38630);
   U14598 : OAI21_X2 port map( A1 => n30699, A2 => n37737, B => n2549, ZN => 
                           n10894);
   U14599 : BUF_X2 port map( I => n28219, Z => n37828);
   U14600 : NAND2_X2 port map( A1 => n8817, A2 => n8814, ZN => n13056);
   U14605 : INV_X2 port map( I => n32622, ZN => n841);
   U14608 : NAND2_X2 port map( A1 => n38397, A2 => n37220, ZN => n11383);
   U14609 : AOI21_X1 port map( A1 => n24467, A2 => n18345, B => n37259, ZN => 
                           n35774);
   U14610 : XOR2_X1 port map( A1 => n37829, A2 => n16806, Z => n16804);
   U14611 : XOR2_X1 port map( A1 => n25113, A2 => n25189, Z => n25208);
   U14612 : OAI22_X2 port map( A1 => n14797, A2 => n14796, B1 => n37246, B2 => 
                           n14795, ZN => n37881);
   U14614 : XOR2_X1 port map( A1 => n11887, A2 => n11615, Z => n9023);
   U14615 : XOR2_X1 port map( A1 => n13617, A2 => n23903, Z => n11887);
   U14618 : OAI22_X2 port map( A1 => n36021, A2 => n33449, B1 => n37831, B2 => 
                           n37830, ZN => n3649);
   U14624 : NOR2_X2 port map( A1 => n24609, A2 => n39704, ZN => n37831);
   U14626 : XOR2_X1 port map( A1 => n25257, A2 => n37832, Z => n25122);
   U14635 : XOR2_X1 port map( A1 => n25224, A2 => n25116, Z => n37832);
   U14646 : NOR2_X2 port map( A1 => n24327, A2 => n2396, ZN => n24175);
   U14648 : XOR2_X1 port map( A1 => n37834, A2 => n2402, Z => n39362);
   U14649 : NAND2_X2 port map( A1 => n36945, A2 => n39670, ZN => n37957);
   U14650 : NAND2_X2 port map( A1 => n37835, A2 => n32999, ZN => n26498);
   U14651 : NOR2_X1 port map( A1 => n37893, A2 => n17954, ZN => n37835);
   U14655 : NOR2_X2 port map( A1 => n37836, A2 => n31074, ZN => n16524);
   U14656 : NOR2_X2 port map( A1 => n31951, A2 => n36888, ZN => n37836);
   U14657 : NOR2_X2 port map( A1 => n18540, A2 => n19227, ZN => n10722);
   U14660 : INV_X2 port map( I => n39401, ZN => n37839);
   U14665 : XOR2_X1 port map( A1 => n16054, A2 => n38147, Z => n34649);
   U14666 : AOI22_X2 port map( A1 => n37733, A2 => n37841, B1 => n24314, B2 => 
                           n7883, ZN => n8961);
   U14667 : NAND2_X2 port map( A1 => n38366, A2 => n33077, ZN => n37841);
   U14668 : INV_X4 port map( I => n12931, ZN => n38338);
   U14669 : XOR2_X1 port map( A1 => n35707, A2 => n33038, Z => n828);
   U14678 : AOI21_X2 port map( A1 => n11942, A2 => n3879, B => n3878, ZN => 
                           n35707);
   U14679 : OAI22_X2 port map( A1 => n24755, A2 => n37852, B1 => n19420, B2 => 
                           n1577, ZN => n17963);
   U14684 : NOR2_X2 port map( A1 => n933, A2 => n36385, ZN => n37852);
   U14685 : XOR2_X1 port map( A1 => n23697, A2 => n31775, Z => n23913);
   U14686 : NAND2_X2 port map( A1 => n22825, A2 => n22824, ZN => n23697);
   U14687 : XOR2_X1 port map( A1 => n34440, A2 => n32646, Z => n17651);
   U14690 : INV_X2 port map( I => n37843, ZN => n35954);
   U14697 : XNOR2_X1 port map( A1 => n12921, A2 => n12920, ZN => n37843);
   U14699 : NAND2_X1 port map( A1 => n22823, A2 => n1630, ZN => n38266);
   U14700 : INV_X4 port map( I => n6945, ZN => n13150);
   U14704 : XOR2_X1 port map( A1 => n22669, A2 => n30406, Z => n30898);
   U14705 : XOR2_X1 port map( A1 => n18595, A2 => n22728, Z => n22669);
   U14710 : NAND2_X2 port map( A1 => n5330, A2 => n37846, ZN => n7445);
   U14711 : NAND2_X2 port map( A1 => n32322, A2 => n37847, ZN => n37846);
   U14712 : NAND2_X2 port map( A1 => n37849, A2 => n37848, ZN => n37847);
   U14713 : INV_X2 port map( I => n1125, ZN => n37848);
   U14716 : INV_X4 port map( I => n30059, ZN => n1403);
   U14717 : XOR2_X1 port map( A1 => n37850, A2 => n11976, Z => n12187);
   U14719 : XOR2_X1 port map( A1 => n27790, A2 => n27789, Z => n37850);
   U14720 : XOR2_X1 port map( A1 => n29039, A2 => n29108, Z => n28895);
   U14721 : XOR2_X1 port map( A1 => n973, A2 => n17039, Z => n29108);
   U14723 : OAI21_X2 port map( A1 => n37851, A2 => n23335, B => n20421, ZN => 
                           n19846);
   U14733 : XOR2_X1 port map( A1 => n26376, A2 => n20425, Z => n20424);
   U14734 : XOR2_X1 port map( A1 => n33178, A2 => n2281, Z => n19652);
   U14735 : NAND2_X2 port map( A1 => n13196, A2 => n13194, ZN => n11533);
   U14737 : NAND3_X2 port map( A1 => n21501, A2 => n39705, A3 => n37853, ZN => 
                           n22332);
   U14738 : NAND2_X1 port map( A1 => n39627, A2 => n21499, ZN => n37853);
   U14740 : NOR2_X2 port map( A1 => n33561, A2 => n26818, ZN => n39054);
   U14741 : XOR2_X1 port map( A1 => n39058, A2 => n33486, Z => n4599);
   U14744 : INV_X1 port map( I => n10213, ZN => n34553);
   U14746 : XNOR2_X1 port map( A1 => n19152, A2 => n10213, ZN => n10939);
   U14749 : NOR2_X2 port map( A1 => n39801, A2 => n4479, ZN => n10213);
   U14750 : NAND2_X2 port map( A1 => n1944, A2 => n28612, ZN => n5928);
   U14753 : XOR2_X1 port map( A1 => n32106, A2 => n26278, Z => n7661);
   U14761 : NAND2_X2 port map( A1 => n5101, A2 => n37854, ZN => n38689);
   U14763 : INV_X4 port map( I => n34217, ZN => n38953);
   U14764 : NOR2_X2 port map( A1 => n28093, A2 => n9266, ZN => n36643);
   U14765 : NAND2_X2 port map( A1 => n26759, A2 => n12755, ZN => n12767);
   U14768 : NOR2_X2 port map( A1 => n37098, A2 => n37856, ZN => n26759);
   U14771 : NOR2_X2 port map( A1 => n19232, A2 => n34603, ZN => n4149);
   U14778 : NAND2_X2 port map( A1 => n21195, A2 => n37857, ZN => n29336);
   U14781 : OR2_X2 port map( A1 => n11657, A2 => n7923, Z => n25625);
   U14783 : XOR2_X1 port map( A1 => n27477, A2 => n35190, Z => n37860);
   U14785 : XOR2_X1 port map( A1 => n22710, A2 => n10558, Z => n35835);
   U14787 : OR2_X1 port map( A1 => n19142, A2 => n6402, Z => n16902);
   U14788 : OAI21_X2 port map( A1 => n31921, A2 => n5953, B => n39413, ZN => 
                           n24583);
   U14790 : XOR2_X1 port map( A1 => n6559, A2 => n37861, Z => n18080);
   U14795 : NOR2_X2 port map( A1 => n31404, A2 => n37862, ZN => n10343);
   U14801 : XOR2_X1 port map( A1 => n11721, A2 => n3488, Z => n39552);
   U14802 : INV_X4 port map( I => n21401, ZN => n20037);
   U14805 : NAND2_X2 port map( A1 => n36275, A2 => n37614, ZN => n18216);
   U14808 : AOI21_X2 port map( A1 => n5124, A2 => n37640, B => n37475, ZN => 
                           n6619);
   U14809 : BUF_X2 port map( I => n31664, Z => n37863);
   U14814 : XOR2_X1 port map( A1 => n3824, A2 => n37864, Z => n38770);
   U14816 : XOR2_X1 port map( A1 => n10083, A2 => n16368, Z => n37864);
   U14817 : NOR2_X2 port map( A1 => n34892, A2 => n3449, ZN => n26952);
   U14824 : XOR2_X1 port map( A1 => n37865, A2 => n26338, Z => n38009);
   U14827 : XOR2_X1 port map( A1 => n10965, A2 => n19681, Z => n37865);
   U14828 : NAND3_X2 port map( A1 => n34116, A2 => n1777, A3 => n1781, ZN => 
                           n31565);
   U14837 : XOR2_X1 port map( A1 => n18490, A2 => n29509, Z => n20956);
   U14838 : NAND3_X2 port map( A1 => n18745, A2 => n25896, A3 => n34565, ZN => 
                           n18490);
   U14840 : NAND3_X2 port map( A1 => n35398, A2 => n35397, A3 => n5839, ZN => 
                           n23714);
   U14843 : INV_X1 port map( I => n8080, ZN => n16115);
   U14847 : NOR2_X1 port map( A1 => n37867, A2 => n37866, ZN => n11650);
   U14848 : INV_X1 port map( I => n20632, ZN => n37866);
   U14849 : NAND2_X1 port map( A1 => n20774, A2 => n8080, ZN => n37867);
   U14851 : XOR2_X1 port map( A1 => n7864, A2 => n7865, Z => n8080);
   U14852 : NAND2_X2 port map( A1 => n5231, A2 => n37868, ZN => n12324);
   U14853 : NAND2_X1 port map( A1 => n39075, A2 => n37226, ZN => n37868);
   U14854 : NAND3_X2 port map( A1 => n27381, A2 => n27382, A3 => n32913, ZN => 
                           n4934);
   U14857 : NOR2_X2 port map( A1 => n1962, A2 => n33964, ZN => n2456);
   U14860 : XOR2_X1 port map( A1 => n37870, A2 => n37869, Z => n37929);
   U14863 : XOR2_X1 port map( A1 => n32972, A2 => n11437, Z => n37870);
   U14866 : INV_X4 port map( I => n35932, ZN => n23505);
   U14868 : XOR2_X1 port map( A1 => n26432, A2 => n32095, Z => n26454);
   U14869 : NAND2_X2 port map( A1 => n11270, A2 => n11269, ZN => n26432);
   U14871 : NAND2_X2 port map( A1 => n18729, A2 => n37871, ZN => n11974);
   U14875 : AOI22_X2 port map( A1 => n18728, A2 => n36237, B1 => n22229, B2 => 
                           n22230, ZN => n37871);
   U14877 : NOR2_X1 port map( A1 => n30629, A2 => n36404, ZN => n8377);
   U14882 : OAI21_X2 port map( A1 => n28594, A2 => n31088, B => n37872, ZN => 
                           n6810);
   U14883 : NAND2_X2 port map( A1 => n28700, A2 => n38669, ZN => n37872);
   U14887 : XOR2_X1 port map( A1 => n22500, A2 => n22509, Z => n22635);
   U14890 : NAND2_X2 port map( A1 => n39275, A2 => n19284, ZN => n22500);
   U14891 : XOR2_X1 port map( A1 => n10658, A2 => n35027, Z => n7666);
   U14895 : XOR2_X1 port map( A1 => n15157, A2 => n28943, Z => n3126);
   U14899 : NAND3_X2 port map( A1 => n16183, A2 => n3128, A3 => n28709, ZN => 
                           n15157);
   U14901 : AND2_X1 port map( A1 => n3850, A2 => n1890, Z => n38910);
   U14902 : NAND2_X1 port map( A1 => n38345, A2 => n8085, ZN => n34891);
   U14905 : NAND2_X2 port map( A1 => n31364, A2 => n11588, ZN => n7225);
   U14907 : XOR2_X1 port map( A1 => n4366, A2 => n38816, Z => n16085);
   U14909 : NOR2_X1 port map( A1 => n2500, A2 => n28442, ZN => n14002);
   U14913 : NAND2_X2 port map( A1 => n14660, A2 => n37873, ZN => n26223);
   U14923 : AOI22_X2 port map( A1 => n11633, A2 => n31133, B1 => n7732, B2 => 
                           n1018, ZN => n37873);
   U14926 : OAI21_X2 port map( A1 => n34601, A2 => n37875, B => n5263, ZN => 
                           n1788);
   U14934 : NOR2_X2 port map( A1 => n32256, A2 => n2735, ZN => n37875);
   U14936 : OAI21_X2 port map( A1 => n12926, A2 => n15755, B => n33944, ZN => 
                           n36016);
   U14939 : NAND2_X2 port map( A1 => n20572, A2 => n38365, ZN => n28285);
   U14941 : INV_X1 port map( I => n9956, ZN => n38414);
   U14943 : NAND2_X2 port map( A1 => n11736, A2 => n33417, ZN => n19061);
   U14944 : NOR2_X2 port map( A1 => n14201, A2 => n32917, ZN => n33417);
   U14945 : XOR2_X1 port map( A1 => n37876, A2 => n37240, Z => n34610);
   U14946 : XOR2_X1 port map( A1 => n27635, A2 => n379, Z => n37876);
   U14949 : XOR2_X1 port map( A1 => n22600, A2 => n22561, Z => n22609);
   U14950 : AOI22_X2 port map( A1 => n9523, A2 => n22239, B1 => n16888, B2 => 
                           n9521, ZN => n22600);
   U14951 : NOR2_X1 port map( A1 => n32594, A2 => n38611, ZN => n38892);
   U14962 : XOR2_X1 port map( A1 => n37877, A2 => n4064, Z => n8057);
   U14963 : XOR2_X1 port map( A1 => n27459, A2 => n38121, Z => n37877);
   U14964 : NAND2_X2 port map( A1 => n7, A2 => n39036, ZN => n31767);
   U14967 : NAND2_X2 port map( A1 => n29644, A2 => n37878, ZN => n33643);
   U14969 : NAND2_X2 port map( A1 => n29643, A2 => n37879, ZN => n37878);
   U14971 : NAND2_X2 port map( A1 => n33630, A2 => n25907, ZN => n26402);
   U14974 : NAND2_X2 port map( A1 => n32574, A2 => n32573, ZN => n15202);
   U14978 : NOR2_X1 port map( A1 => n15174, A2 => n29551, ZN => n21177);
   U14981 : BUF_X2 port map( I => n33047, Z => n37880);
   U14984 : OR2_X2 port map( A1 => n14383, A2 => n860, Z => n26946);
   U14987 : INV_X4 port map( I => n17887, ZN => n6514);
   U14989 : NAND2_X2 port map( A1 => n3545, A2 => n3544, ZN => n17887);
   U14990 : NAND2_X1 port map( A1 => n11521, A2 => n8194, ZN => n36584);
   U14994 : XOR2_X1 port map( A1 => n38180, A2 => n37882, Z => n751);
   U14998 : NOR2_X2 port map( A1 => n12456, A2 => n12458, ZN => n38180);
   U15000 : XOR2_X1 port map( A1 => n24926, A2 => n25181, Z => n6352);
   U15007 : NOR2_X2 port map( A1 => n7350, A2 => n12643, ZN => n24926);
   U15010 : XOR2_X1 port map( A1 => n5473, A2 => n5472, Z => n5518);
   U15011 : AOI22_X2 port map( A1 => n31030, A2 => n28463, B1 => n34312, B2 => 
                           n30757, ZN => n28791);
   U15012 : NAND2_X2 port map( A1 => n33022, A2 => n19452, ZN => n25697);
   U15013 : XOR2_X1 port map( A1 => n11189, A2 => n37094, Z => n11192);
   U15015 : XOR2_X1 port map( A1 => n37884, A2 => n20536, Z => n11188);
   U15018 : XOR2_X1 port map( A1 => n5553, A2 => n39512, Z => n37884);
   U15019 : NAND2_X2 port map( A1 => n11669, A2 => n7577, ZN => n32832);
   U15022 : OAI22_X2 port map( A1 => n30145, A2 => n35234, B1 => n18241, B2 => 
                           n30132, ZN => n29015);
   U15024 : NAND2_X2 port map( A1 => n7366, A2 => n22896, ZN => n23456);
   U15033 : NOR2_X1 port map( A1 => n3356, A2 => n1106, ZN => n3360);
   U15035 : NOR2_X2 port map( A1 => n37120, A2 => n37885, ZN => n36705);
   U15036 : NOR2_X1 port map( A1 => n274, A2 => n28150, ZN => n37885);
   U15037 : NOR2_X1 port map( A1 => n28616, A2 => n180, ZN => n28454);
   U15040 : NAND2_X2 port map( A1 => n34871, A2 => n14330, ZN => n180);
   U15041 : NAND2_X2 port map( A1 => n38957, A2 => n28170, ZN => n28676);
   U15044 : XOR2_X1 port map( A1 => n28891, A2 => n6433, Z => n29159);
   U15047 : NAND3_X2 port map( A1 => n15630, A2 => n28678, A3 => n15629, ZN => 
                           n6433);
   U15053 : NAND2_X2 port map( A1 => n1445, A2 => n34166, ZN => n38743);
   U15057 : AOI21_X2 port map( A1 => n16353, A2 => n30057, B => n30059, ZN => 
                           n3045);
   U15060 : XOR2_X1 port map( A1 => n4413, A2 => n22741, Z => n7358);
   U15064 : NAND2_X2 port map( A1 => n35727, A2 => n20123, ZN => n4413);
   U15068 : INV_X2 port map( I => n26255, ZN => n1505);
   U15071 : NAND3_X2 port map( A1 => n38866, A2 => n30468, A3 => n16612, ZN => 
                           n26255);
   U15073 : AOI21_X2 port map( A1 => n15790, A2 => n15791, B => n15789, ZN => 
                           n12548);
   U15078 : OAI21_X2 port map( A1 => n38387, A2 => n9888, B => n37886, ZN => 
                           n7852);
   U15080 : NAND2_X1 port map( A1 => n37887, A2 => n2597, ZN => n37886);
   U15082 : NOR2_X1 port map( A1 => n15049, A2 => n38702, ZN => n37887);
   U15083 : XOR2_X1 port map( A1 => n14136, A2 => n37888, Z => n16907);
   U15085 : XOR2_X1 port map( A1 => n29055, A2 => n29056, Z => n37888);
   U15086 : NAND2_X1 port map( A1 => n29265, A2 => n1406, ZN => n37942);
   U15091 : XOR2_X1 port map( A1 => n16610, A2 => n29432, Z => n37889);
   U15094 : XOR2_X1 port map( A1 => n15916, A2 => n16324, Z => n23954);
   U15097 : AOI21_X2 port map( A1 => n15799, A2 => n18762, B => n15949, ZN => 
                           n15916);
   U15098 : NOR2_X1 port map( A1 => n17692, A2 => n17691, ZN => n39645);
   U15107 : NAND3_X1 port map( A1 => n6487, A2 => n3947, A3 => n6486, ZN => 
                           n32460);
   U15114 : AOI22_X2 port map( A1 => n31498, A2 => n9295, B1 => n27374, B2 => 
                           n27266, ZN => n27749);
   U15120 : XOR2_X1 port map( A1 => n3889, A2 => n27677, Z => n3886);
   U15121 : NAND3_X1 port map( A1 => n13191, A2 => n36371, A3 => n2654, ZN => 
                           n11455);
   U15122 : BUF_X4 port map( I => n1033, Z => n39156);
   U15124 : NAND2_X2 port map( A1 => n17227, A2 => n27046, ZN => n18195);
   U15125 : AOI22_X2 port map( A1 => n34170, A2 => n19946, B1 => n37186, B2 => 
                           n28131, ZN => n37892);
   U15129 : OAI21_X2 port map( A1 => n37167, A2 => n23127, B => n34124, ZN => 
                           n9862);
   U15133 : NAND2_X2 port map( A1 => n1302, A2 => n5487, ZN => n18312);
   U15134 : NAND2_X1 port map( A1 => n26902, A2 => n19673, ZN => n37900);
   U15135 : NAND2_X1 port map( A1 => n37077, A2 => n27018, ZN => n39503);
   U15137 : OAI21_X2 port map( A1 => n13261, A2 => n29377, B => n29453, ZN => 
                           n29379);
   U15139 : XOR2_X1 port map( A1 => n13703, A2 => n27631, Z => n31731);
   U15142 : AOI21_X2 port map( A1 => n30678, A2 => n4231, B => n30416, ZN => 
                           n27631);
   U15144 : XOR2_X1 port map( A1 => n26571, A2 => n12838, Z => n26197);
   U15147 : NOR2_X2 port map( A1 => n18631, A2 => n18630, ZN => n12838);
   U15148 : AND2_X1 port map( A1 => n32377, A2 => n6945, Z => n13830);
   U15149 : XOR2_X1 port map( A1 => n32660, A2 => n30976, Z => n37934);
   U15153 : BUF_X4 port map( I => n26556, Z => n11667);
   U15155 : NOR2_X1 port map( A1 => n36352, A2 => n3013, ZN => n37893);
   U15156 : NAND2_X2 port map( A1 => n37894, A2 => n39566, ZN => n27858);
   U15158 : NAND2_X1 port map( A1 => n17718, A2 => n17719, ZN => n37894);
   U15162 : XOR2_X1 port map( A1 => n25318, A2 => n25320, Z => n12330);
   U15166 : NAND2_X2 port map( A1 => n33043, A2 => n2530, ZN => n25318);
   U15174 : NAND2_X2 port map( A1 => n13782, A2 => n30766, ZN => n30845);
   U15175 : XOR2_X1 port map( A1 => n24036, A2 => n18849, Z => n23756);
   U15176 : OAI22_X2 port map( A1 => n21040, A2 => n17458, B1 => n15524, B2 => 
                           n4382, ZN => n11668);
   U15177 : OR2_X1 port map( A1 => n23198, A2 => n32856, Z => n8462);
   U15179 : NAND3_X1 port map( A1 => n9107, A2 => n9878, A3 => n37619, ZN => 
                           n37897);
   U15183 : OAI22_X2 port map( A1 => n22275, A2 => n35771, B1 => n16772, B2 => 
                           n14196, ZN => n13785);
   U15194 : BUF_X2 port map( I => n32535, Z => n37898);
   U15195 : AOI21_X1 port map( A1 => n34299, A2 => n8988, B => n35767, ZN => 
                           n6383);
   U15197 : INV_X2 port map( I => n19477, ZN => n35767);
   U15202 : NAND2_X2 port map( A1 => n11514, A2 => n11516, ZN => n19477);
   U15204 : OAI21_X2 port map( A1 => n10753, A2 => n31780, B => n1548, ZN => 
                           n32481);
   U15207 : INV_X2 port map( I => n26808, ZN => n26810);
   U15208 : XOR2_X1 port map( A1 => n6033, A2 => n29666, Z => n13229);
   U15213 : NAND2_X2 port map( A1 => n38318, A2 => n13231, ZN => n6033);
   U15214 : NOR2_X1 port map( A1 => n35264, A2 => n36910, ZN => n36976);
   U15215 : INV_X4 port map( I => n16559, ZN => n19893);
   U15216 : AOI22_X2 port map( A1 => n7945, A2 => n1072, B1 => n6788, B2 => 
                           n7946, ZN => n7324);
   U15217 : XOR2_X1 port map( A1 => n8897, A2 => n33133, Z => n10009);
   U15221 : AND2_X1 port map( A1 => n32566, A2 => n33593, Z => n3690);
   U15227 : NAND2_X2 port map( A1 => n3102, A2 => n8685, ZN => n32566);
   U15228 : NAND2_X2 port map( A1 => n16182, A2 => n23482, ZN => n38691);
   U15229 : NAND2_X2 port map( A1 => n19414, A2 => n14632, ZN => n9686);
   U15231 : XOR2_X1 port map( A1 => n38815, A2 => n38814, Z => n13872);
   U15234 : NAND2_X2 port map( A1 => n31079, A2 => n15534, ZN => n39163);
   U15235 : NOR2_X2 port map( A1 => n37900, A2 => n35311, ZN => n9956);
   U15236 : NAND2_X1 port map( A1 => n39569, A2 => n929, ZN => n4512);
   U15241 : NAND2_X2 port map( A1 => n8843, A2 => n15365, ZN => n31679);
   U15243 : OAI21_X2 port map( A1 => n38527, A2 => n38528, B => n35761, ZN => 
                           n8843);
   U15246 : INV_X2 port map( I => n28758, ZN => n1426);
   U15247 : OR2_X1 port map( A1 => n28758, A2 => n20597, Z => n8850);
   U15249 : INV_X4 port map( I => n9855, ZN => n11807);
   U15250 : NAND2_X2 port map( A1 => n32826, A2 => n32827, ZN => n9855);
   U15251 : NAND2_X2 port map( A1 => n36374, A2 => n37901, ZN => n32854);
   U15255 : NAND3_X2 port map( A1 => n13585, A2 => n25762, A3 => n25761, ZN => 
                           n19450);
   U15256 : OAI22_X2 port map( A1 => n548, A2 => n33401, B1 => n1119, B2 => 
                           n18858, ZN => n13637);
   U15259 : AOI22_X2 port map( A1 => n17754, A2 => n27235, B1 => n36234, B2 => 
                           n27233, ZN => n35902);
   U15260 : XOR2_X1 port map( A1 => n26411, A2 => n16216, Z => n14770);
   U15261 : XOR2_X1 port map( A1 => n26532, A2 => n26591, Z => n26411);
   U15265 : XOR2_X1 port map( A1 => n34800, A2 => n33364, Z => n3771);
   U15266 : XOR2_X1 port map( A1 => n828, A2 => n25191, Z => n15686);
   U15267 : XOR2_X1 port map( A1 => n140, A2 => n36363, Z => n34213);
   U15271 : XOR2_X1 port map( A1 => n29126, A2 => n2142, Z => n2005);
   U15272 : AND2_X1 port map( A1 => n23613, A2 => n1627, Z => n32294);
   U15276 : NAND2_X1 port map( A1 => n30453, A2 => n33356, ZN => n35018);
   U15278 : OAI21_X1 port map( A1 => n39806, A2 => n2830, B => n32193, ZN => 
                           n1743);
   U15280 : NAND2_X2 port map( A1 => n15579, A2 => n23237, ZN => n23459);
   U15284 : NOR2_X2 port map( A1 => n327, A2 => n32850, ZN => n15579);
   U15285 : XOR2_X1 port map( A1 => n23794, A2 => n23671, Z => n17398);
   U15287 : NAND2_X2 port map( A1 => n6141, A2 => n6139, ZN => n23671);
   U15291 : NOR2_X1 port map( A1 => n39510, A2 => n37902, ZN => n38462);
   U15292 : OAI22_X1 port map( A1 => n18424, A2 => n30144, B1 => n30143, B2 => 
                           n18588, ZN => n37902);
   U15293 : OAI21_X2 port map( A1 => n37981, A2 => n37880, B => n4369, ZN => 
                           n38504);
   U15295 : XOR2_X1 port map( A1 => n32239, A2 => n17463, Z => n8299);
   U15297 : NAND2_X2 port map( A1 => n36429, A2 => n3031, ZN => n32239);
   U15298 : NAND2_X1 port map( A1 => n15575, A2 => n18827, ZN => n25866);
   U15301 : NAND2_X2 port map( A1 => n32658, A2 => n17740, ZN => n15575);
   U15304 : XOR2_X1 port map( A1 => n15676, A2 => n35240, Z => n36383);
   U15306 : INV_X2 port map( I => n17989, ZN => n14024);
   U15313 : NAND2_X1 port map( A1 => n20555, A2 => n35687, ZN => n22809);
   U15315 : INV_X4 port map( I => n23198, ZN => n38283);
   U15321 : BUF_X2 port map( I => n2576, Z => n37905);
   U15327 : NOR2_X2 port map( A1 => n39584, A2 => n34399, ZN => n38956);
   U15328 : XOR2_X1 port map( A1 => n31633, A2 => n17581, Z => n12138);
   U15330 : NAND2_X2 port map( A1 => n1177, A2 => n1399, ZN => n12955);
   U15334 : OAI22_X2 port map( A1 => n37906, A2 => n23416, B1 => n23418, B2 => 
                           n36130, ZN => n3521);
   U15339 : XOR2_X1 port map( A1 => n23677, A2 => n23947, Z => n1791);
   U15341 : NAND2_X1 port map( A1 => n15223, A2 => n16430, ZN => n38182);
   U15343 : NAND2_X2 port map( A1 => n5146, A2 => n39174, ZN => n5171);
   U15346 : NOR2_X2 port map( A1 => n7170, A2 => n37907, ZN => n7168);
   U15347 : NOR2_X2 port map( A1 => n8120, A2 => n11807, ZN => n37907);
   U15348 : XOR2_X1 port map( A1 => n13531, A2 => n25316, Z => n39315);
   U15356 : XOR2_X1 port map( A1 => n4592, A2 => n32190, Z => n18655);
   U15357 : INV_X2 port map( I => n29803, ZN => n966);
   U15363 : INV_X2 port map( I => n5869, ZN => n4411);
   U15370 : XOR2_X1 port map( A1 => n5312, A2 => n32915, Z => n5869);
   U15372 : NAND3_X2 port map( A1 => n8041, A2 => n18721, A3 => n8042, ZN => 
                           n33102);
   U15376 : XOR2_X1 port map( A1 => n27642, A2 => n27861, Z => n17276);
   U15378 : XOR2_X1 port map( A1 => n27828, A2 => n27766, Z => n27861);
   U15380 : XOR2_X1 port map( A1 => n37908, A2 => n13172, Z => n23132);
   U15382 : XOR2_X1 port map( A1 => n13174, A2 => n22658, Z => n37908);
   U15385 : XOR2_X1 port map( A1 => n17612, A2 => n37909, Z => n32662);
   U15386 : XOR2_X1 port map( A1 => n2585, A2 => n963, Z => n37909);
   U15387 : XOR2_X1 port map( A1 => n29297, A2 => n28967, Z => n29033);
   U15392 : XOR2_X1 port map( A1 => n7848, A2 => n29166, Z => n29297);
   U15396 : XOR2_X1 port map( A1 => n16709, A2 => n37910, Z => n6848);
   U15397 : XOR2_X1 port map( A1 => n282, A2 => n27825, Z => n37910);
   U15398 : NAND2_X2 port map( A1 => n15701, A2 => n15775, ZN => n13386);
   U15402 : XOR2_X1 port map( A1 => n22703, A2 => n17756, Z => n18001);
   U15403 : NAND2_X2 port map( A1 => n21452, A2 => n21453, ZN => n22703);
   U15404 : XOR2_X1 port map( A1 => n12570, A2 => n37912, Z => n12200);
   U15407 : XOR2_X1 port map( A1 => n20509, A2 => n23894, Z => n12570);
   U15408 : INV_X1 port map( I => n24039, ZN => n37912);
   U15415 : OR2_X1 port map( A1 => n24271, A2 => n18342, Z => n38115);
   U15416 : NAND2_X2 port map( A1 => n37970, A2 => n37913, ZN => n23251);
   U15420 : AND2_X1 port map( A1 => n2840, A2 => n22042, Z => n10623);
   U15429 : NOR2_X2 port map( A1 => n7636, A2 => n37920, ZN => n37919);
   U15437 : INV_X2 port map( I => n18253, ZN => n37920);
   U15441 : NOR2_X2 port map( A1 => n18637, A2 => n23060, ZN => n18636);
   U15446 : NAND2_X2 port map( A1 => n37922, A2 => n37921, ZN => n18637);
   U15448 : INV_X1 port map( I => n18209, ZN => n37921);
   U15454 : XOR2_X1 port map( A1 => n15532, A2 => n23971, Z => n20615);
   U15460 : AOI21_X2 port map( A1 => n28216, A2 => n28219, B => n28217, ZN => 
                           n16467);
   U15461 : NAND2_X2 port map( A1 => n987, A2 => n16631, ZN => n28219);
   U15462 : NOR2_X2 port map( A1 => n23522, A2 => n3708, ZN => n23318);
   U15464 : AOI21_X1 port map( A1 => n16869, A2 => n33510, B => n28214, ZN => 
                           n16868);
   U15467 : XOR2_X1 port map( A1 => n4136, A2 => n13939, Z => n4135);
   U15471 : NAND2_X2 port map( A1 => n11491, A2 => n11492, ZN => n31515);
   U15478 : XOR2_X1 port map( A1 => n28500, A2 => n28886, Z => n29105);
   U15480 : OAI21_X2 port map( A1 => n3877, A2 => n8878, B => n37925, ZN => 
                           n3874);
   U15481 : OAI21_X2 port map( A1 => n15620, A2 => n34060, B => n10882, ZN => 
                           n37925);
   U15483 : BUF_X2 port map( I => n31305, Z => n37926);
   U15484 : XOR2_X1 port map( A1 => n37247, A2 => n6134, Z => n38467);
   U15486 : XOR2_X1 port map( A1 => n11319, A2 => n15930, Z => n6458);
   U15488 : AND2_X2 port map( A1 => n8479, A2 => n35476, Z => n26805);
   U15492 : XOR2_X1 port map( A1 => n3320, A2 => n27475, Z => n18846);
   U15493 : XOR2_X1 port map( A1 => n7910, A2 => n16162, Z => n27475);
   U15495 : NOR3_X1 port map( A1 => n26220, A2 => n2000, A3 => n26839, ZN => 
                           n16298);
   U15496 : OAI22_X1 port map( A1 => n29276, A2 => n17773, B1 => n13886, B2 => 
                           n29275, ZN => n5088);
   U15500 : NAND2_X2 port map( A1 => n7088, A2 => n29125, ZN => n33833);
   U15501 : NAND2_X2 port map( A1 => n37248, A2 => n13823, ZN => n29125);
   U15502 : NAND3_X2 port map( A1 => n37927, A2 => n38062, A3 => n38061, ZN => 
                           n29057);
   U15505 : XOR2_X1 port map( A1 => n8003, A2 => n37928, Z => n135);
   U15508 : XOR2_X1 port map( A1 => n16673, A2 => n25225, Z => n37928);
   U15509 : AOI21_X2 port map( A1 => n37890, A2 => n27372, B => n16042, ZN => 
                           n13526);
   U15511 : INV_X2 port map( I => n16040, ZN => n16042);
   U15513 : NOR2_X2 port map( A1 => n17795, A2 => n27123, ZN => n16040);
   U15515 : NOR2_X2 port map( A1 => n20035, A2 => n31798, ZN => n23590);
   U15519 : NAND2_X1 port map( A1 => n4190, A2 => n10834, ZN => n26012);
   U15521 : NAND2_X2 port map( A1 => n4018, A2 => n9335, ZN => n4190);
   U15523 : INV_X2 port map( I => n37929, ZN => n33972);
   U15524 : XOR2_X1 port map( A1 => n5289, A2 => n15960, Z => n5320);
   U15528 : NAND2_X2 port map( A1 => n5287, A2 => n33190, ZN => n5289);
   U15529 : NAND2_X2 port map( A1 => n7892, A2 => n14869, ZN => n16548);
   U15530 : NAND3_X1 port map( A1 => n24806, A2 => n1026, A3 => n19565, ZN => 
                           n37931);
   U15531 : INV_X2 port map( I => n18035, ZN => n28425);
   U15534 : BUF_X4 port map( I => n21660, Z => n39627);
   U15535 : NOR2_X2 port map( A1 => n209, A2 => n1424, ZN => n12398);
   U15536 : NAND2_X2 port map( A1 => n14107, A2 => n23252, ZN => n23890);
   U15540 : INV_X2 port map( I => n32239, ZN => n37932);
   U15545 : XOR2_X1 port map( A1 => n25204, A2 => n25114, Z => n15758);
   U15550 : NOR2_X2 port map( A1 => n13637, A2 => n13638, ZN => n25204);
   U15552 : XOR2_X1 port map( A1 => n5761, A2 => n5760, Z => n12758);
   U15556 : NAND2_X2 port map( A1 => n31862, A2 => n32607, ZN => n27383);
   U15558 : NAND2_X2 port map( A1 => n37933, A2 => n39734, ZN => n10118);
   U15559 : NAND3_X2 port map( A1 => n39416, A2 => n3958, A3 => n38883, ZN => 
                           n37933);
   U15561 : NAND2_X2 port map( A1 => n39216, A2 => n20671, ZN => n27205);
   U15568 : NOR2_X2 port map( A1 => n27139, A2 => n27140, ZN => n27197);
   U15570 : OAI22_X2 port map( A1 => n19433, A2 => n26692, B1 => n26691, B2 => 
                           n39825, ZN => n27139);
   U15571 : XOR2_X1 port map( A1 => n37935, A2 => n19815, Z => Ciphertext(151))
                           ;
   U15574 : OAI22_X1 port map( A1 => n28658, A2 => n28657, B1 => n17977, B2 => 
                           n1197, ZN => n31705);
   U15579 : NAND3_X2 port map( A1 => n2338, A2 => n20184, A3 => n16154, ZN => 
                           n2023);
   U15580 : XOR2_X1 port map( A1 => n4282, A2 => n38659, Z => n16931);
   U15582 : NAND2_X1 port map( A1 => n36060, A2 => n36059, ZN => n39388);
   U15583 : OAI21_X2 port map( A1 => n29867, A2 => n29843, B => n29869, ZN => 
                           n20894);
   U15589 : XOR2_X1 port map( A1 => n1503, A2 => n26584, Z => n26482);
   U15591 : NAND3_X2 port map( A1 => n13103, A2 => n25827, A3 => n25828, ZN => 
                           n26584);
   U15593 : INV_X2 port map( I => n37937, ZN => n26249);
   U15597 : XNOR2_X1 port map( A1 => n2069, A2 => n2066, ZN => n37937);
   U15601 : OAI22_X2 port map( A1 => n20370, A2 => n29629, B1 => n20371, B2 => 
                           n13441, ZN => n20369);
   U15607 : CLKBUF_X4 port map( I => n33424, Z => n38275);
   U15608 : INV_X1 port map( I => n21790, ZN => n37939);
   U15616 : XNOR2_X1 port map( A1 => n17804, A2 => n8796, ZN => n38558);
   U15617 : NAND2_X2 port map( A1 => n38737, A2 => n29103, ZN => n29236);
   U15619 : NAND2_X2 port map( A1 => n38034, A2 => n33102, ZN => n38918);
   U15622 : INV_X1 port map( I => n9935, ZN => n37940);
   U15623 : NAND2_X1 port map( A1 => n37940, A2 => n36076, ZN => n5642);
   U15624 : XOR2_X1 port map( A1 => n17957, A2 => n37941, Z => n10812);
   U15628 : XOR2_X1 port map( A1 => n3223, A2 => n29050, Z => n37941);
   U15632 : OR2_X1 port map( A1 => n26029, A2 => n18320, Z => n25804);
   U15634 : NAND2_X2 port map( A1 => n8407, A2 => n26041, ZN => n25825);
   U15635 : NAND2_X2 port map( A1 => n25814, A2 => n25813, ZN => n26023);
   U15636 : NAND3_X1 port map( A1 => n29278, A2 => n29284, A3 => n1379, ZN => 
                           n29279);
   U15648 : INV_X2 port map( I => n19518, ZN => n35618);
   U15652 : NAND3_X2 port map( A1 => n5024, A2 => n5023, A3 => n13438, ZN => 
                           n19518);
   U15655 : NAND2_X1 port map( A1 => n7305, A2 => n19465, ZN => n14427);
   U15656 : XOR2_X1 port map( A1 => n3703, A2 => n3668, Z => n31725);
   U15658 : XOR2_X1 port map( A1 => n15013, A2 => n22664, Z => n15012);
   U15659 : XOR2_X1 port map( A1 => n37944, A2 => n3404, Z => n18860);
   U15672 : XOR2_X1 port map( A1 => n27765, A2 => n37991, Z => n37944);
   U15673 : XOR2_X1 port map( A1 => n20303, A2 => n24949, Z => n25158);
   U15674 : XOR2_X1 port map( A1 => n20304, A2 => n24946, Z => n20303);
   U15679 : XOR2_X1 port map( A1 => n35243, A2 => n20483, Z => n38069);
   U15684 : NAND2_X2 port map( A1 => n24875, A2 => n1580, ZN => n9213);
   U15686 : XOR2_X1 port map( A1 => n37945, A2 => n29411, Z => Ciphertext(40));
   U15691 : NAND3_X2 port map( A1 => n7733, A2 => n15042, A3 => n14517, ZN => 
                           n37945);
   U15693 : INV_X2 port map( I => n25177, ZN => n1557);
   U15695 : NAND2_X2 port map( A1 => n32268, A2 => n24871, ZN => n25177);
   U15698 : AOI21_X2 port map( A1 => n11094, A2 => n28772, B => n37946, ZN => 
                           n11389);
   U15703 : NOR3_X2 port map( A1 => n5662, A2 => n31418, A3 => n10618, ZN => 
                           n37946);
   U15704 : XOR2_X1 port map( A1 => n17250, A2 => n37947, Z => n5317);
   U15705 : XOR2_X1 port map( A1 => n31550, A2 => n29070, Z => n37947);
   U15711 : NAND3_X2 port map( A1 => n8769, A2 => n38001, A3 => n2771, ZN => 
                           n37948);
   U15712 : AND2_X1 port map( A1 => n12682, A2 => n3873, Z => n2735);
   U15713 : NAND2_X2 port map( A1 => n37950, A2 => n14192, ZN => n35151);
   U15714 : AND2_X1 port map( A1 => n14262, A2 => n25643, Z => n37950);
   U15719 : NOR2_X2 port map( A1 => n6127, A2 => n15268, ZN => n12628);
   U15721 : NAND2_X1 port map( A1 => n32418, A2 => n18529, ZN => n27873);
   U15722 : AOI21_X2 port map( A1 => n36269, A2 => n37368, B => n3045, ZN => 
                           n3600);
   U15728 : XNOR2_X1 port map( A1 => n27516, A2 => n27566, ZN => n13883);
   U15732 : XOR2_X1 port map( A1 => n37952, A2 => n20420, Z => Ciphertext(117))
                           ;
   U15733 : BUF_X4 port map( I => n16040, Z => n1475);
   U15734 : XOR2_X1 port map( A1 => n11739, A2 => n19851, Z => n6746);
   U15736 : NAND2_X2 port map( A1 => n3348, A2 => n430, ZN => n11739);
   U15737 : NOR2_X2 port map( A1 => n39235, A2 => n17770, ZN => n34446);
   U15748 : NAND2_X2 port map( A1 => n9514, A2 => n7904, ZN => n17770);
   U15749 : INV_X2 port map( I => n26015, ZN => n26120);
   U15750 : OAI22_X2 port map( A1 => n15254, A2 => n25501, B1 => n15647, B2 => 
                           n37183, ZN => n26015);
   U15759 : XOR2_X1 port map( A1 => n37953, A2 => n28793, Z => n28796);
   U15760 : XOR2_X1 port map( A1 => n29260, A2 => n36990, Z => n37953);
   U15766 : OR2_X1 port map( A1 => n686, A2 => n21912, Z => n3692);
   U15767 : OR2_X1 port map( A1 => n39444, A2 => n19223, Z => n25502);
   U15771 : XOR2_X1 port map( A1 => n27749, A2 => n27537, Z => n27665);
   U15773 : NOR2_X2 port map( A1 => n38860, A2 => n36791, ZN => n31371);
   U15782 : XOR2_X1 port map( A1 => n28873, A2 => n10430, Z => n13315);
   U15785 : XNOR2_X1 port map( A1 => n25170, A2 => n25285, ZN => n31445);
   U15791 : XOR2_X1 port map( A1 => n25284, A2 => n9701, Z => n25170);
   U15792 : NAND2_X2 port map( A1 => n12733, A2 => n37954, ZN => n30379);
   U15793 : INV_X2 port map( I => n2394, ZN => n37954);
   U15799 : XOR2_X1 port map( A1 => n35177, A2 => n38964, Z => n10866);
   U15803 : NAND2_X2 port map( A1 => n36639, A2 => n35603, ZN => n35177);
   U15805 : INV_X2 port map( I => n26946, ZN => n14135);
   U15806 : XOR2_X1 port map( A1 => n6774, A2 => n15782, Z => n29943);
   U15807 : XOR2_X1 port map( A1 => n15930, A2 => n17078, Z => n13763);
   U15809 : AOI22_X2 port map( A1 => n38424, A2 => n33705, B1 => n21028, B2 => 
                           n24750, ZN => n15930);
   U15811 : AND2_X1 port map( A1 => n15049, A2 => n2597, Z => n36621);
   U15812 : NOR2_X2 port map( A1 => n10883, A2 => n28685, ZN => n9935);
   U15813 : INV_X4 port map( I => n7291, ZN => n38305);
   U15814 : NAND2_X2 port map( A1 => n32206, A2 => n5665, ZN => n10883);
   U15815 : NAND2_X2 port map( A1 => n1441, A2 => n1438, ZN => n37960);
   U15817 : NAND2_X2 port map( A1 => n33713, A2 => n31202, ZN => n22293);
   U15818 : NAND2_X2 port map( A1 => n3323, A2 => n3327, ZN => n20397);
   U15819 : XOR2_X1 port map( A1 => n26313, A2 => n26312, Z => n26809);
   U15821 : XOR2_X1 port map( A1 => n34686, A2 => n13608, Z => n13787);
   U15826 : AND2_X2 port map( A1 => n37961, A2 => n7245, Z => n7250);
   U15827 : OAI21_X1 port map( A1 => n3374, A2 => n16745, B => n7044, ZN => 
                           n37961);
   U15835 : NAND3_X2 port map( A1 => n19575, A2 => n26946, A3 => n26857, ZN => 
                           n36942);
   U15836 : NAND2_X2 port map( A1 => n23767, A2 => n23796, ZN => n33987);
   U15839 : AOI21_X2 port map( A1 => n37962, A2 => n4298, B => n9040, ZN => 
                           n4297);
   U15840 : OAI21_X2 port map( A1 => n19545, A2 => n21804, B => n36735, ZN => 
                           n37963);
   U15845 : NAND2_X2 port map( A1 => n12620, A2 => n12618, ZN => n12617);
   U15850 : NAND2_X2 port map( A1 => n7008, A2 => n35232, ZN => n21213);
   U15851 : NOR2_X1 port map( A1 => n24829, A2 => n20128, ZN => n15688);
   U15852 : NAND2_X2 port map( A1 => n24625, A2 => n10421, ZN => n20128);
   U15854 : XOR2_X1 port map( A1 => n37964, A2 => n13313, Z => n13312);
   U15856 : XOR2_X1 port map( A1 => n38290, A2 => n37965, Z => n37964);
   U15857 : INV_X2 port map( I => n19035, ZN => n37965);
   U15858 : INV_X4 port map( I => n15049, ZN => n38404);
   U15859 : XOR2_X1 port map( A1 => n28830, A2 => n7744, Z => n29029);
   U15860 : NAND2_X2 port map( A1 => n34753, A2 => n31887, ZN => n28830);
   U15864 : OR2_X1 port map( A1 => n21497, A2 => n14418, Z => n15707);
   U15865 : BUF_X2 port map( I => n33514, Z => n37966);
   U15866 : NAND3_X2 port map( A1 => n25435, A2 => n39269, A3 => n4467, ZN => 
                           n12893);
   U15867 : OR2_X2 port map( A1 => n13561, A2 => n14381, Z => n22816);
   U15868 : NAND2_X2 port map( A1 => n34883, A2 => n38102, ZN => n26532);
   U15869 : XOR2_X1 port map( A1 => n24935, A2 => n24999, Z => n20618);
   U15870 : NAND3_X2 port map( A1 => n14782, A2 => n9912, A3 => n15689, ZN => 
                           n24999);
   U15872 : XOR2_X1 port map( A1 => n821, A2 => n37968, Z => n35077);
   U15876 : XOR2_X1 port map( A1 => n37969, A2 => n32309, Z => n39710);
   U15882 : XOR2_X1 port map( A1 => n5848, A2 => n29602, Z => n37969);
   U15887 : OR2_X1 port map( A1 => n19590, A2 => n26042, Z => n25828);
   U15889 : NAND3_X2 port map( A1 => n22962, A2 => n23020, A3 => n10507, ZN => 
                           n37970);
   U15890 : INV_X1 port map( I => n28647, ZN => n30951);
   U15891 : OAI21_X2 port map( A1 => n9099, A2 => n37971, B => n9098, ZN => 
                           n7974);
   U15895 : AOI22_X2 port map( A1 => n14807, A2 => n26661, B1 => n39342, B2 => 
                           n14458, ZN => n37971);
   U15900 : NAND2_X1 port map( A1 => n6876, A2 => n21101, ZN => n5773);
   U15903 : NAND2_X2 port map( A1 => n34001, A2 => n27363, ZN => n6876);
   U15904 : NAND2_X2 port map( A1 => n37972, A2 => n19812, ZN => n22573);
   U15909 : NAND2_X2 port map( A1 => n17896, A2 => n17898, ZN => n37972);
   U15913 : XOR2_X1 port map( A1 => n37973, A2 => n29001, Z => n32718);
   U15914 : NAND2_X1 port map( A1 => n18199, A2 => n13029, ZN => n23351);
   U15915 : NAND2_X2 port map( A1 => n35067, A2 => n22846, ZN => n18199);
   U15918 : XOR2_X1 port map( A1 => n12393, A2 => n37974, Z => n22639);
   U15931 : INV_X2 port map( I => n8312, ZN => n37974);
   U15932 : OAI22_X2 port map( A1 => n7816, A2 => n916, B1 => n7815, B2 => 
                           n7814, ZN => n8312);
   U15939 : XOR2_X1 port map( A1 => n25189, A2 => n20707, Z => n25317);
   U15944 : NAND2_X2 port map( A1 => n38083, A2 => n471, ZN => n25189);
   U15946 : AOI21_X2 port map( A1 => n5254, A2 => n1034, B => n7657, ZN => 
                           n37975);
   U15947 : NAND2_X2 port map( A1 => n37977, A2 => n20583, ZN => n36908);
   U15950 : XOR2_X1 port map( A1 => n36515, A2 => n24054, Z => n798);
   U15955 : NAND3_X1 port map( A1 => n7251, A2 => n32682, A3 => n36935, ZN => 
                           n8048);
   U15956 : XOR2_X1 port map( A1 => n26597, A2 => n13232, Z => n11600);
   U15957 : XOR2_X1 port map( A1 => n38137, A2 => n10776, Z => n26597);
   U15960 : NAND2_X2 port map( A1 => n35709, A2 => n31060, ZN => n29803);
   U15962 : NAND3_X1 port map( A1 => n23013, A2 => n4573, A3 => n39527, ZN => 
                           n16400);
   U15963 : XOR2_X1 port map( A1 => n26574, A2 => n26575, Z => n36864);
   U15966 : AND2_X1 port map( A1 => n21232, A2 => n27028, Z => n37978);
   U15967 : NAND3_X1 port map( A1 => n18408, A2 => n22274, A3 => n22151, ZN => 
                           n22152);
   U15968 : XOR2_X1 port map( A1 => n37979, A2 => n12322, Z => n36868);
   U15971 : XOR2_X1 port map( A1 => n39118, A2 => n35639, Z => n37979);
   U15974 : NOR2_X2 port map( A1 => n19228, A2 => n37980, ZN => n2273);
   U15976 : NAND2_X2 port map( A1 => n5249, A2 => n5248, ZN => n26031);
   U15977 : XOR2_X1 port map( A1 => n5241, A2 => n37261, Z => n484);
   U15978 : NOR2_X2 port map( A1 => n37981, A2 => n28639, ZN => n35788);
   U15983 : XOR2_X1 port map( A1 => n9185, A2 => n3963, Z => n3501);
   U15987 : XOR2_X1 port map( A1 => n12310, A2 => n12311, Z => n25421);
   U15989 : NAND3_X2 port map( A1 => n6900, A2 => n6903, A3 => n37982, ZN => 
                           n38981);
   U15990 : XOR2_X1 port map( A1 => n27688, A2 => n27502, Z => n10540);
   U15991 : XOR2_X1 port map( A1 => n20706, A2 => n13245, Z => n27688);
   U15993 : NOR2_X2 port map( A1 => n30778, A2 => n13034, ZN => n39486);
   U16002 : OR2_X1 port map( A1 => n31014, A2 => n17095, Z => n27334);
   U16007 : NAND2_X2 port map( A1 => n34309, A2 => n12391, ZN => n26329);
   U16008 : NAND2_X2 port map( A1 => n15867, A2 => n29792, ZN => n29795);
   U16010 : OAI22_X2 port map( A1 => n3693, A2 => n3986, B1 => n20616, B2 => 
                           n775, ZN => n31326);
   U16019 : NOR3_X1 port map( A1 => n1531, A2 => n33446, A3 => n39678, ZN => 
                           n9944);
   U16022 : XOR2_X1 port map( A1 => n18399, A2 => n1051, Z => n295);
   U16030 : NAND2_X2 port map( A1 => n6785, A2 => n6784, ZN => n18399);
   U16032 : OAI21_X2 port map( A1 => n9656, A2 => n24717, B => n24719, ZN => 
                           n37985);
   U16034 : NAND2_X2 port map( A1 => n37986, A2 => n19951, ZN => n36538);
   U16038 : NAND2_X2 port map( A1 => n30539, A2 => n26702, ZN => n37986);
   U16039 : NOR2_X1 port map( A1 => n26872, A2 => n5935, ZN => n35345);
   U16046 : NAND2_X1 port map( A1 => n37988, A2 => n37987, ZN => n372);
   U16047 : NAND2_X1 port map( A1 => n1385, A2 => n30128, ZN => n37987);
   U16048 : NOR3_X2 port map( A1 => n707, A2 => n7315, A3 => n684, ZN => n10650
                           );
   U16050 : AOI21_X1 port map( A1 => n12617, A2 => n35534, B => n19481, ZN => 
                           n34373);
   U16051 : NAND2_X2 port map( A1 => n39492, A2 => n11156, ZN => n19481);
   U16053 : NAND2_X2 port map( A1 => n31253, A2 => n7397, ZN => n6191);
   U16054 : NAND2_X2 port map( A1 => n37989, A2 => n6934, ZN => n25086);
   U16055 : OAI21_X2 port map( A1 => n34047, A2 => n31743, B => n37990, ZN => 
                           n3082);
   U16056 : XOR2_X1 port map( A1 => n31807, A2 => n38069, Z => n37991);
   U16057 : OR2_X2 port map( A1 => n11481, A2 => n12770, Z => n9080);
   U16060 : OR2_X1 port map( A1 => n20596, A2 => n293, Z => n19756);
   U16063 : NAND2_X1 port map( A1 => n23131, A2 => n22674, ZN => n22800);
   U16068 : NAND2_X2 port map( A1 => n23226, A2 => n23337, ZN => n23534);
   U16071 : NAND3_X2 port map( A1 => n20191, A2 => n22708, A3 => n16400, ZN => 
                           n23226);
   U16075 : INV_X2 port map( I => n19094, ZN => n38921);
   U16079 : NAND2_X2 port map( A1 => n5716, A2 => n37992, ZN => n31722);
   U16081 : NOR2_X2 port map( A1 => n4784, A2 => n4785, ZN => n37992);
   U16091 : BUF_X2 port map( I => n37051, Z => n37993);
   U16092 : INV_X2 port map( I => n33750, ZN => n16566);
   U16099 : OAI22_X2 port map( A1 => n33001, A2 => n32948, B1 => n36711, B2 => 
                           n38092, ZN => n38187);
   U16101 : INV_X2 port map( I => n25978, ZN => n37997);
   U16105 : CLKBUF_X4 port map( I => n36509, Z => n39632);
   U16113 : NAND3_X1 port map( A1 => n37153, A2 => n38643, A3 => n26645, ZN => 
                           n38831);
   U16121 : XOR2_X1 port map( A1 => n38736, A2 => n25207, Z => n31724);
   U16123 : XOR2_X1 port map( A1 => n25241, A2 => n25181, Z => n25183);
   U16127 : AOI21_X2 port map( A1 => n24657, A2 => n24656, B => n14781, ZN => 
                           n25241);
   U16129 : NAND2_X1 port map( A1 => n10940, A2 => n15873, ZN => n31184);
   U16131 : XOR2_X1 port map( A1 => n24055, A2 => n14312, Z => n38000);
   U16133 : BUF_X2 port map( I => n26625, Z => n38002);
   U16137 : XOR2_X1 port map( A1 => n7416, A2 => n869, Z => n34358);
   U16138 : NAND2_X1 port map( A1 => n4772, A2 => n36546, ZN => n6831);
   U16148 : NAND2_X2 port map( A1 => n7540, A2 => n12995, ZN => n36546);
   U16149 : XOR2_X1 port map( A1 => n38003, A2 => n1050, Z => Ciphertext(180));
   U16153 : AOI22_X1 port map( A1 => n30201, A2 => n14387, B1 => n32263, B2 => 
                           n36738, ZN => n38003);
   U16157 : AND2_X1 port map( A1 => n26933, A2 => n4411, Z => n5720);
   U16161 : XOR2_X1 port map( A1 => n38005, A2 => n29239, Z => Ciphertext(17));
   U16163 : AOI22_X1 port map( A1 => n35185, A2 => n15482, B1 => n15483, B2 => 
                           n29237, ZN => n38005);
   U16164 : OR2_X1 port map( A1 => n29241, A2 => n13815, Z => n9716);
   U16169 : OAI22_X2 port map( A1 => n6619, A2 => n5030, B1 => n37640, B2 => 
                           n37212, ZN => n8605);
   U16170 : INV_X2 port map( I => n27774, ZN => n4366);
   U16171 : NAND2_X2 port map( A1 => n4120, A2 => n4119, ZN => n13807);
   U16177 : XOR2_X1 port map( A1 => n4560, A2 => n38006, Z => n19167);
   U16190 : XOR2_X1 port map( A1 => n4558, A2 => n4559, Z => n38006);
   U16191 : INV_X2 port map( I => n17876, ZN => n20498);
   U16205 : OAI22_X2 port map( A1 => n29693, A2 => n29843, B1 => n17877, B2 => 
                           n29867, ZN => n17876);
   U16209 : OAI21_X2 port map( A1 => n38008, A2 => n38007, B => n8623, ZN => 
                           n57);
   U16210 : NOR2_X2 port map( A1 => n8621, A2 => n8622, ZN => n38008);
   U16212 : INV_X2 port map( I => n30217, ZN => n14869);
   U16214 : OAI22_X2 port map( A1 => n31025, A2 => n4807, B1 => n2322, B2 => 
                           n2321, ZN => n30217);
   U16215 : XOR2_X1 port map( A1 => n20715, A2 => n24060, Z => n20516);
   U16216 : NOR2_X1 port map( A1 => n27199, A2 => n4353, ZN => n27030);
   U16217 : INV_X2 port map( I => n27395, ZN => n27199);
   U16218 : NOR2_X1 port map( A1 => n24279, A2 => n17911, ZN => n34046);
   U16219 : XOR2_X1 port map( A1 => n38009, A2 => n26419, Z => n34580);
   U16221 : NAND2_X1 port map( A1 => n35098, A2 => n33514, ZN => n36007);
   U16223 : OAI21_X2 port map( A1 => n7890, A2 => n25366, B => n38662, ZN => 
                           n33514);
   U16230 : NAND3_X2 port map( A1 => n34654, A2 => n17813, A3 => n22029, ZN => 
                           n9127);
   U16231 : NOR2_X2 port map( A1 => n1535, A2 => n32775, ZN => n25466);
   U16239 : BUF_X2 port map( I => n19587, Z => n38011);
   U16243 : NAND2_X1 port map( A1 => n22931, A2 => n7160, ZN => n38012);
   U16245 : BUF_X2 port map( I => n25487, Z => n38013);
   U16246 : XOR2_X1 port map( A1 => n23685, A2 => n14289, Z => n16833);
   U16251 : NAND2_X2 port map( A1 => n5181, A2 => n5183, ZN => n14289);
   U16252 : XOR2_X1 port map( A1 => n12690, A2 => n15844, Z => n9400);
   U16255 : XOR2_X1 port map( A1 => n9757, A2 => n27746, Z => n12690);
   U16257 : NOR2_X2 port map( A1 => n21521, A2 => n21587, ZN => n8600);
   U16258 : NAND2_X2 port map( A1 => n1081, A2 => n37508, ZN => n9082);
   U16262 : AOI21_X2 port map( A1 => n27686, A2 => n28193, B => n37164, ZN => 
                           n38014);
   U16264 : INV_X2 port map( I => n38015, ZN => n34987);
   U16265 : XOR2_X1 port map( A1 => n31485, A2 => n12084, Z => n38015);
   U16278 : NAND2_X1 port map( A1 => n11067, A2 => n37095, ZN => n29372);
   U16282 : OAI22_X2 port map( A1 => n29345, A2 => n39647, B1 => n12479, B2 => 
                           n19896, ZN => n35465);
   U16283 : INV_X2 port map( I => n19846, ZN => n35936);
   U16284 : NAND2_X2 port map( A1 => n5768, A2 => n7770, ZN => n24898);
   U16287 : NOR3_X2 port map( A1 => n34071, A2 => n35297, A3 => n32797, ZN => 
                           n27140);
   U16290 : XOR2_X1 port map( A1 => n25, A2 => n25148, Z => n33527);
   U16291 : XOR2_X1 port map( A1 => n18366, A2 => n38016, Z => n26995);
   U16300 : XOR2_X1 port map( A1 => n26434, A2 => n31414, Z => n38016);
   U16308 : OR2_X1 port map( A1 => n35300, A2 => n32010, Z => n24370);
   U16309 : OAI21_X2 port map( A1 => n11133, A2 => n24119, B => n11131, ZN => 
                           n7529);
   U16310 : NOR2_X2 port map( A1 => n35360, A2 => n38017, ZN => n32608);
   U16314 : XOR2_X1 port map( A1 => n20424, A2 => n38018, Z => n33895);
   U16317 : XOR2_X1 port map( A1 => n20730, A2 => n26222, Z => n38018);
   U16322 : NAND2_X2 port map( A1 => n18788, A2 => n19499, ZN => n39232);
   U16324 : XNOR2_X1 port map( A1 => n38208, A2 => n16618, ZN => n39239);
   U16329 : XOR2_X1 port map( A1 => n20586, A2 => n24052, Z => n19188);
   U16336 : NAND2_X2 port map( A1 => n39581, A2 => n39333, ZN => n24052);
   U16338 : OAI21_X2 port map( A1 => n13445, A2 => n37904, B => n12307, ZN => 
                           n9847);
   U16339 : XOR2_X1 port map( A1 => n32895, A2 => n4900, Z => n7140);
   U16340 : NOR2_X1 port map( A1 => n21047, A2 => n23020, ZN => n38019);
   U16341 : XOR2_X1 port map( A1 => n33322, A2 => n29463, Z => n5094);
   U16348 : OAI22_X2 port map( A1 => n23593, A2 => n4148, B1 => n4149, B2 => 
                           n23594, ZN => n33322);
   U16350 : OAI21_X2 port map( A1 => n17863, A2 => n17862, B => n10894, ZN => 
                           n25113);
   U16355 : INV_X2 port map( I => n5063, ZN => n38668);
   U16356 : NAND2_X1 port map( A1 => n26918, A2 => n13392, ZN => n33062);
   U16357 : NAND2_X2 port map( A1 => n10461, A2 => n35427, ZN => n27009);
   U16358 : XOR2_X1 port map( A1 => n13439, A2 => n9246, Z => n23802);
   U16360 : NAND2_X2 port map( A1 => n33698, A2 => n23584, ZN => n13439);
   U16365 : OAI21_X2 port map( A1 => n23578, A2 => n6945, B => n1138, ZN => 
                           n21296);
   U16366 : NAND2_X2 port map( A1 => n38576, A2 => n38020, ZN => n36634);
   U16369 : OAI21_X2 port map( A1 => n33101, A2 => n36556, B => n34044, ZN => 
                           n38020);
   U16370 : NAND2_X2 port map( A1 => n1759, A2 => n33516, ZN => n28066);
   U16376 : NOR2_X2 port map( A1 => n37105, A2 => n36634, ZN => n38916);
   U16382 : NAND2_X2 port map( A1 => n16579, A2 => n12160, ZN => n13516);
   U16392 : OAI21_X2 port map( A1 => n28623, A2 => n33283, B => n19161, ZN => 
                           n33519);
   U16393 : NAND2_X2 port map( A1 => n33283, A2 => n2147, ZN => n19161);
   U16394 : AND2_X1 port map( A1 => n35427, A2 => n9369, Z => n27430);
   U16395 : BUF_X2 port map( I => n15037, Z => n36549);
   U16398 : NOR3_X2 port map( A1 => n33513, A2 => n39605, A3 => n24282, ZN => 
                           n32542);
   U16399 : NAND2_X2 port map( A1 => n29862, A2 => n9649, ZN => n29908);
   U16400 : XOR2_X1 port map( A1 => n24938, A2 => n25030, Z => n38992);
   U16401 : NOR2_X2 port map( A1 => n24607, A2 => n12846, ZN => n25030);
   U16403 : NAND3_X2 port map( A1 => n23511, A2 => n23510, A3 => n11245, ZN => 
                           n15299);
   U16405 : NAND2_X2 port map( A1 => n12156, A2 => n35427, ZN => n11256);
   U16407 : OR2_X1 port map( A1 => n30156, A2 => n14254, Z => n31357);
   U16408 : XOR2_X1 port map( A1 => n29100, A2 => n38384, Z => n30156);
   U16412 : OR2_X1 port map( A1 => n5282, A2 => n24515, Z => n34143);
   U16415 : NAND2_X1 port map( A1 => n38023, A2 => n1536, ZN => n5292);
   U16417 : OAI22_X1 port map( A1 => n1531, A2 => n25692, B1 => n8014, B2 => 
                           n12500, ZN => n38023);
   U16421 : AOI22_X2 port map( A1 => n8946, A2 => n33867, B1 => n27652, B2 => 
                           n13955, ZN => n8944);
   U16423 : AOI21_X1 port map( A1 => n28235, A2 => n28234, B => n11283, ZN => 
                           n38512);
   U16424 : XOR2_X1 port map( A1 => n19862, A2 => n19902, Z => n6923);
   U16425 : XOR2_X1 port map( A1 => n27594, A2 => n27796, Z => n27753);
   U16427 : NAND3_X2 port map( A1 => n17151, A2 => n15275, A3 => n15277, ZN => 
                           n27796);
   U16435 : XOR2_X1 port map( A1 => n38026, A2 => n2176, Z => n8526);
   U16436 : NAND2_X2 port map( A1 => n36849, A2 => n32081, ZN => n22488);
   U16438 : XOR2_X1 port map( A1 => n9036, A2 => n29282, Z => n13700);
   U16439 : NAND2_X2 port map( A1 => n137, A2 => n6039, ZN => n9036);
   U16440 : NOR2_X1 port map( A1 => n36854, A2 => n28234, ZN => n4415);
   U16442 : NOR2_X1 port map( A1 => n2573, A2 => n4531, ZN => n12379);
   U16444 : NAND2_X2 port map( A1 => n4244, A2 => n38027, ZN => n15716);
   U16445 : NAND2_X1 port map( A1 => n33061, A2 => n18116, ZN => n38027);
   U16448 : NAND2_X1 port map( A1 => n39017, A2 => n15358, ZN => n35709);
   U16452 : NAND2_X2 port map( A1 => n14216, A2 => n7643, ZN => n31486);
   U16453 : XOR2_X1 port map( A1 => n31541, A2 => n4301, Z => n22233);
   U16456 : XOR2_X1 port map( A1 => n38028, A2 => n26204, Z => n33067);
   U16463 : XNOR2_X1 port map( A1 => n16610, A2 => n9576, ZN => n26204);
   U16465 : NOR2_X2 port map( A1 => n149, A2 => n4467, ZN => n38029);
   U16475 : OAI21_X2 port map( A1 => n31177, A2 => n31175, B => n38030, ZN => 
                           n39268);
   U16482 : AOI22_X2 port map( A1 => n14645, A2 => n8735, B1 => n16590, B2 => 
                           n15872, ZN => n38030);
   U16483 : XOR2_X1 port map( A1 => n13569, A2 => n27470, Z => n13568);
   U16484 : OR2_X1 port map( A1 => n10375, A2 => n33431, Z => n22834);
   U16486 : XOR2_X1 port map( A1 => n22651, A2 => n12267, Z => n22463);
   U16488 : OAI21_X2 port map( A1 => n16624, A2 => n16623, B => n22081, ZN => 
                           n22651);
   U16497 : OAI22_X2 port map( A1 => n1234, A2 => n14394, B1 => n26719, B2 => 
                           n735, ZN => n11248);
   U16499 : XOR2_X1 port map( A1 => n38427, A2 => n33576, Z => n10686);
   U16504 : NAND2_X2 port map( A1 => n16325, A2 => n14461, ZN => n5509);
   U16510 : XOR2_X1 port map( A1 => n28827, A2 => n29052, Z => n8909);
   U16512 : NAND2_X2 port map( A1 => n8910, A2 => n8911, ZN => n28827);
   U16513 : XOR2_X1 port map( A1 => n38031, A2 => n1700, Z => Ciphertext(6));
   U16515 : NOR2_X1 port map( A1 => n9606, A2 => n9607, ZN => n38031);
   U16516 : XOR2_X1 port map( A1 => n10406, A2 => n10407, Z => n11657);
   U16517 : OAI21_X2 port map( A1 => n24355, A2 => n8359, B => n19818, ZN => 
                           n35666);
   U16519 : NOR2_X2 port map( A1 => n39074, A2 => n32069, ZN => n24355);
   U16521 : INV_X2 port map( I => n13761, ZN => n29219);
   U16522 : NAND3_X2 port map( A1 => n35502, A2 => n30655, A3 => n32267, ZN => 
                           n13761);
   U16524 : NAND3_X2 port map( A1 => n25360, A2 => n19971, A3 => n19311, ZN => 
                           n39108);
   U16525 : NAND2_X1 port map( A1 => n13663, A2 => n17248, ZN => n39402);
   U16526 : INV_X4 port map( I => n24709, ZN => n6491);
   U16527 : NAND2_X2 port map( A1 => n12422, A2 => n12424, ZN => n24709);
   U16537 : XOR2_X1 port map( A1 => n21079, A2 => n38033, Z => n19948);
   U16541 : XOR2_X1 port map( A1 => n31692, A2 => n28853, Z => n38033);
   U16546 : NOR2_X2 port map( A1 => n27341, A2 => n32205, ZN => n27133);
   U16561 : INV_X2 port map( I => n26888, ZN => n27341);
   U16564 : NAND3_X2 port map( A1 => n26698, A2 => n142, A3 => n26699, ZN => 
                           n26888);
   U16565 : NAND3_X2 port map( A1 => n36556, A2 => n19070, A3 => n17810, ZN => 
                           n38034);
   U16566 : XOR2_X1 port map( A1 => n38035, A2 => n19128, Z => Ciphertext(20));
   U16567 : NAND3_X1 port map( A1 => n17955, A2 => n6841, A3 => n6842, ZN => 
                           n38035);
   U16568 : XOR2_X1 port map( A1 => n11794, A2 => n23869, Z => n15114);
   U16571 : NOR2_X2 port map( A1 => n38036, A2 => n24154, ZN => n24698);
   U16572 : XOR2_X1 port map( A1 => n13703, A2 => n13877, Z => n39613);
   U16574 : OAI22_X2 port map( A1 => n4089, A2 => n4253, B1 => n38572, B2 => 
                           n4254, ZN => n13877);
   U16576 : XOR2_X1 port map( A1 => n20294, A2 => n18153, Z => n31752);
   U16577 : NOR2_X2 port map( A1 => n23616, A2 => n38037, ZN => n24038);
   U16581 : AOI21_X2 port map( A1 => n36635, A2 => n39434, B => n23614, ZN => 
                           n38037);
   U16587 : XOR2_X1 port map( A1 => n38038, A2 => n18993, Z => Ciphertext(15));
   U16590 : NOR2_X1 port map( A1 => n14200, A2 => n14197, ZN => n38038);
   U16593 : NAND2_X1 port map( A1 => n26761, A2 => n26810, ZN => n11515);
   U16595 : INV_X1 port map( I => n24974, ZN => n35339);
   U16596 : XOR2_X1 port map( A1 => n36748, A2 => n23609, Z => n23677);
   U16599 : XOR2_X1 port map( A1 => n30610, A2 => n30609, Z => n5274);
   U16602 : XOR2_X1 port map( A1 => n26321, A2 => n39667, Z => n26630);
   U16604 : NAND2_X2 port map( A1 => n38040, A2 => n38039, ZN => n18303);
   U16607 : OAI21_X2 port map( A1 => n13421, A2 => n21892, B => n21893, ZN => 
                           n38039);
   U16613 : OAI21_X2 port map( A1 => n21896, A2 => n15528, B => n21895, ZN => 
                           n38040);
   U16614 : XOR2_X1 port map( A1 => n10562, A2 => n27859, Z => n10483);
   U16615 : XOR2_X1 port map( A1 => n27779, A2 => n27778, Z => n27859);
   U16618 : BUF_X2 port map( I => n38619, Z => n38041);
   U16620 : INV_X4 port map( I => n26935, ZN => n1093);
   U16625 : INV_X2 port map( I => n29070, ZN => n7489);
   U16643 : XOR2_X1 port map( A1 => n8634, A2 => n23950, Z => n636);
   U16645 : XOR2_X1 port map( A1 => n33322, A2 => n23680, Z => n23950);
   U16646 : XOR2_X1 port map( A1 => n25179, A2 => n25096, Z => n31563);
   U16647 : NAND2_X2 port map( A1 => n12832, A2 => n24085, ZN => n25096);
   U16648 : NAND2_X2 port map( A1 => n7892, A2 => n33437, ZN => n9200);
   U16649 : NAND2_X2 port map( A1 => n2684, A2 => n2685, ZN => n23889);
   U16651 : NOR2_X2 port map( A1 => n24802, A2 => n35901, ZN => n15414);
   U16656 : XOR2_X1 port map( A1 => n6130, A2 => n26026, Z => n26399);
   U16664 : NOR2_X2 port map( A1 => n33950, A2 => n25692, ZN => n8222);
   U16667 : XOR2_X1 port map( A1 => n32349, A2 => n38043, Z => n9986);
   U16668 : INV_X2 port map( I => n25200, ZN => n38043);
   U16669 : XOR2_X1 port map( A1 => n25296, A2 => n24991, Z => n25200);
   U16676 : NAND2_X2 port map( A1 => n11614, A2 => n1433, ZN => n13780);
   U16681 : XOR2_X1 port map( A1 => n39378, A2 => n30849, Z => n38048);
   U16682 : NAND2_X2 port map( A1 => n17335, A2 => n2458, ZN => n17333);
   U16687 : OR3_X2 port map( A1 => n15515, A2 => n25480, A3 => n16933, Z => 
                           n25529);
   U16690 : OAI22_X2 port map( A1 => n17225, A2 => n1061, B1 => n1062, B2 => 
                           n20566, ZN => n39240);
   U16691 : NAND3_X2 port map( A1 => n29370, A2 => n39677, A3 => n4669, ZN => 
                           n39208);
   U16692 : OAI21_X2 port map( A1 => n11054, A2 => n37106, B => n38044, ZN => 
                           n8542);
   U16694 : XOR2_X1 port map( A1 => n38045, A2 => n38711, Z => n25544);
   U16697 : XOR2_X1 port map( A1 => n5433, A2 => n38458, Z => n38045);
   U16699 : XOR2_X1 port map( A1 => n5803, A2 => n5804, Z => n39353);
   U16702 : XOR2_X1 port map( A1 => n38046, A2 => n19738, Z => Ciphertext(92));
   U16703 : NAND4_X2 port map( A1 => n29714, A2 => n29716, A3 => n29713, A4 => 
                           n29715, ZN => n38046);
   U16706 : NAND2_X2 port map( A1 => n31960, A2 => n19911, ZN => n15868);
   U16710 : XOR2_X1 port map( A1 => n38048, A2 => n23410, Z => n34473);
   U16713 : XOR2_X1 port map( A1 => n8852, A2 => n18430, Z => n29024);
   U16716 : NAND2_X2 port map( A1 => n8854, A2 => n8853, ZN => n18430);
   U16718 : XOR2_X1 port map( A1 => n12840, A2 => n798, Z => n19295);
   U16719 : NAND3_X2 port map( A1 => n20177, A2 => n22819, A3 => n20176, ZN => 
                           n38724);
   U16725 : AOI22_X2 port map( A1 => n3309, A2 => n5591, B1 => n23412, B2 => 
                           n1636, ZN => n38049);
   U16726 : OAI21_X2 port map( A1 => n38782, A2 => n19941, B => n16677, ZN => 
                           n38050);
   U16732 : XOR2_X1 port map( A1 => n26590, A2 => n19450, Z => n13496);
   U16735 : INV_X2 port map( I => n26272, ZN => n26687);
   U16737 : XOR2_X1 port map( A1 => n29057, A2 => n18133, Z => n19428);
   U16738 : NAND2_X2 port map( A1 => n28338, A2 => n9442, ZN => n18133);
   U16739 : XOR2_X1 port map( A1 => n35065, A2 => n23982, Z => n14386);
   U16743 : OAI22_X2 port map( A1 => n10495, A2 => n10494, B1 => n5049, B2 => 
                           n1134, ZN => n35065);
   U16747 : XOR2_X1 port map( A1 => n26389, A2 => n26436, Z => n26508);
   U16749 : NAND2_X2 port map( A1 => n25926, A2 => n9226, ZN => n26389);
   U16750 : XOR2_X1 port map( A1 => n1661, A2 => n3953, Z => n13842);
   U16751 : XOR2_X1 port map( A1 => n22534, A2 => n22520, Z => n22524);
   U16753 : XOR2_X1 port map( A1 => n22628, A2 => n1662, Z => n22534);
   U16755 : INV_X2 port map( I => n38052, ZN => n15466);
   U16760 : XOR2_X1 port map( A1 => Plaintext(168), A2 => Key(168), Z => n38052
                           );
   U16762 : NAND2_X2 port map( A1 => n11337, A2 => n26935, ZN => n11336);
   U16764 : NAND3_X2 port map( A1 => n28491, A2 => n28490, A3 => n28489, ZN => 
                           n28492);
   U16766 : BUF_X2 port map( I => n29344, Z => n29458);
   U16767 : INV_X2 port map( I => n38053, ZN => n17307);
   U16770 : NOR2_X2 port map( A1 => n21460, A2 => n21459, ZN => n38053);
   U16776 : OAI21_X2 port map( A1 => n21539, A2 => n21542, B => n9424, ZN => 
                           n21459);
   U16782 : NOR2_X2 port map( A1 => n12191, A2 => n5487, ZN => n5490);
   U16783 : INV_X2 port map( I => n18681, ZN => n12191);
   U16784 : NAND2_X2 port map( A1 => n35006, A2 => n17201, ZN => n18681);
   U16787 : XOR2_X1 port map( A1 => n2627, A2 => n269, Z => n3207);
   U16790 : NAND2_X2 port map( A1 => n1834, A2 => n32184, ZN => n2627);
   U16791 : NAND2_X2 port map( A1 => n11225, A2 => n36483, ZN => n27435);
   U16794 : INV_X1 port map( I => n19279, ZN => n38626);
   U16795 : XOR2_X1 port map( A1 => n12145, A2 => n39579, Z => n36239);
   U16796 : NAND2_X2 port map( A1 => n11279, A2 => n11280, ZN => n35203);
   U16801 : AOI22_X2 port map( A1 => n37225, A2 => n38055, B1 => n2012, B2 => 
                           n17960, ZN => n2009);
   U16804 : INV_X2 port map( I => n1036, ZN => n38055);
   U16805 : NAND2_X2 port map( A1 => n38949, A2 => n39748, ZN => n34350);
   U16808 : NOR2_X1 port map( A1 => n15048, A2 => n11737, ZN => n38765);
   U16818 : NAND2_X2 port map( A1 => n38056, A2 => n27543, ZN => n16853);
   U16828 : NAND2_X2 port map( A1 => n38057, A2 => n13093, ZN => n13414);
   U16832 : OAI21_X2 port map( A1 => n32873, A2 => n32872, B => n37883, ZN => 
                           n38057);
   U16833 : NAND2_X2 port map( A1 => n14833, A2 => n4424, ZN => n2480);
   U16838 : XOR2_X1 port map( A1 => n38352, A2 => n39698, Z => n38058);
   U16846 : INV_X2 port map( I => n5282, ZN => n24603);
   U16849 : XOR2_X1 port map( A1 => n5625, A2 => n17884, Z => n27496);
   U16854 : NOR2_X1 port map( A1 => n22265, A2 => n22267, ZN => n11684);
   U16856 : OAI21_X1 port map( A1 => n36910, A2 => n9914, B => n29224, ZN => 
                           n13771);
   U16857 : INV_X1 port map( I => n29220, ZN => n36910);
   U16863 : AND2_X1 port map( A1 => n31357, A2 => n35870, Z => n38236);
   U16865 : OAI21_X2 port map( A1 => n38059, A2 => n34817, B => n28212, ZN => 
                           n39087);
   U16869 : NOR2_X2 port map( A1 => n28213, A2 => n16950, ZN => n38059);
   U16880 : INV_X2 port map( I => n8475, ZN => n38799);
   U16881 : XOR2_X1 port map( A1 => n27516, A2 => n19800, Z => n31070);
   U16883 : NAND2_X2 port map( A1 => n14058, A2 => n14057, ZN => n27516);
   U16884 : OAI21_X2 port map( A1 => n32343, A2 => n32344, B => n11679, ZN => 
                           n20190);
   U16886 : NOR2_X2 port map( A1 => n6615, A2 => n38284, ZN => n32343);
   U16888 : NAND3_X2 port map( A1 => n6195, A2 => n32545, A3 => n6192, ZN => 
                           n36386);
   U16890 : AOI21_X2 port map( A1 => n29873, A2 => n29869, B => n33297, ZN => 
                           n38217);
   U16893 : NAND3_X2 port map( A1 => n38757, A2 => n31170, A3 => n35547, ZN => 
                           n30095);
   U16896 : INV_X2 port map( I => n13333, ZN => n32555);
   U16897 : NOR3_X2 port map( A1 => n30694, A2 => n25622, A3 => n33785, ZN => 
                           n3010);
   U16903 : OR2_X1 port map( A1 => n6932, A2 => n16619, Z => n4949);
   U16904 : XOR2_X1 port map( A1 => n6727, A2 => n25263, Z => n25153);
   U16909 : NOR2_X1 port map( A1 => n29627, A2 => n29617, ZN => n38063);
   U16911 : XOR2_X1 port map( A1 => n26437, A2 => n26009, Z => n26528);
   U16914 : OR2_X2 port map( A1 => n27875, A2 => n17378, Z => n28199);
   U16915 : XOR2_X1 port map( A1 => n16054, A2 => n6758, Z => n29060);
   U16919 : AOI21_X2 port map( A1 => n6789, A2 => n6788, B => n38064, ZN => 
                           n6786);
   U16920 : NOR3_X1 port map( A1 => n5239, A2 => n5352, A3 => n34008, ZN => 
                           n38064);
   U16922 : INV_X2 port map( I => n27588, ZN => n27587);
   U16923 : NAND2_X2 port map( A1 => n35332, A2 => n2722, ZN => n27588);
   U16930 : NAND2_X2 port map( A1 => n10231, A2 => n11616, ZN => n26899);
   U16938 : INV_X2 port map( I => n38066, ZN => n16174);
   U16941 : XNOR2_X1 port map( A1 => n32431, A2 => n32432, ZN => n38066);
   U16947 : NAND3_X1 port map( A1 => n14375, A2 => n38168, A3 => n35855, ZN => 
                           n18352);
   U16950 : XOR2_X1 port map( A1 => n10233, A2 => n5584, Z => n20960);
   U16951 : NAND3_X2 port map( A1 => n9142, A2 => n29180, A3 => n7933, ZN => 
                           n30117);
   U16952 : OR2_X1 port map( A1 => n23468, A2 => n23467, Z => n7534);
   U16954 : AND2_X1 port map( A1 => n19782, A2 => n24465, Z => n35873);
   U16956 : NAND2_X2 port map( A1 => n38437, A2 => n26042, ZN => n17178);
   U16957 : AND2_X1 port map( A1 => n36810, A2 => n32471, Z => n16299);
   U16965 : INV_X2 port map( I => n24827, ZN => n11271);
   U16968 : NAND3_X2 port map( A1 => n1877, A2 => n1875, A3 => n5432, ZN => 
                           n24827);
   U16979 : XOR2_X1 port map( A1 => n27480, A2 => n20167, Z => n20166);
   U16982 : XOR2_X1 port map( A1 => n27851, A2 => n5750, Z => n27480);
   U16985 : XOR2_X1 port map( A1 => n38067, A2 => n29295, Z => Ciphertext(3));
   U16987 : XOR2_X1 port map( A1 => n28783, A2 => n12989, Z => n29128);
   U16990 : NAND2_X2 port map( A1 => n5397, A2 => n5398, ZN => n28783);
   U17001 : NAND2_X2 port map( A1 => n910, A2 => n2678, ZN => n25977);
   U17004 : NOR2_X2 port map( A1 => n19544, A2 => n7790, ZN => n9025);
   U17007 : XOR2_X1 port map( A1 => n14353, A2 => n17925, Z => n14454);
   U17012 : INV_X1 port map( I => n38070, ZN => n35360);
   U17013 : OAI21_X1 port map( A1 => n34567, A2 => n34568, B => n28735, ZN => 
                           n38070);
   U17015 : INV_X2 port map( I => n12572, ZN => n30211);
   U17016 : NAND3_X2 port map( A1 => n39432, A2 => n7893, A3 => n39431, ZN => 
                           n12572);
   U17017 : INV_X4 port map( I => n17685, ZN => n937);
   U17022 : AOI22_X2 port map( A1 => n17794, A2 => n29263, B1 => n37185, B2 => 
                           n16123, ZN => n38071);
   U17024 : NAND2_X1 port map( A1 => n38072, A2 => n10703, ZN => n39551);
   U17025 : NOR2_X1 port map( A1 => n39393, A2 => n39392, ZN => n38072);
   U17026 : XOR2_X1 port map( A1 => n23874, A2 => n19608, Z => n23876);
   U17029 : INV_X2 port map( I => n24887, ZN => n38073);
   U17033 : AND2_X1 port map( A1 => n7044, A2 => n38073, Z => n17863);
   U17044 : XOR2_X1 port map( A1 => n22789, A2 => n22728, Z => n22581);
   U17048 : NOR2_X2 port map( A1 => n39190, A2 => n34433, ZN => n34753);
   U17049 : AND2_X1 port map( A1 => n19560, A2 => n24872, Z => n30422);
   U17050 : NAND2_X2 port map( A1 => n31161, A2 => n18148, ZN => n19560);
   U17053 : NAND2_X2 port map( A1 => n4246, A2 => n4247, ZN => n38619);
   U17058 : XOR2_X1 port map( A1 => n36617, A2 => n38076, Z => n35544);
   U17070 : XNOR2_X1 port map( A1 => n27845, A2 => n8875, ZN => n2437);
   U17074 : NOR2_X2 port map( A1 => n38247, A2 => n25820, ZN => n31473);
   U17075 : NAND2_X2 port map( A1 => n18686, A2 => n18685, ZN => n5819);
   U17078 : AOI22_X2 port map( A1 => n21943, A2 => n20923, B1 => n16128, B2 => 
                           n16052, ZN => n18685);
   U17081 : INV_X4 port map( I => n3293, ZN => n21583);
   U17085 : NAND2_X1 port map( A1 => n31461, A2 => n8349, ZN => n38077);
   U17086 : XOR2_X1 port map( A1 => n8654, A2 => n37252, Z => n9590);
   U17087 : XNOR2_X1 port map( A1 => n39391, A2 => n8532, ZN => n8654);
   U17088 : NOR2_X2 port map( A1 => n35377, A2 => n34962, ZN => n31945);
   U17089 : BUF_X2 port map( I => n27314, Z => n38079);
   U17090 : XOR2_X1 port map( A1 => n10636, A2 => n38080, Z => n10733);
   U17098 : XOR2_X1 port map( A1 => n12026, A2 => n12480, Z => n38080);
   U17104 : INV_X2 port map( I => n38081, ZN => n6640);
   U17115 : OAI21_X1 port map( A1 => n12675, A2 => n10563, B => n38959, ZN => 
                           n9439);
   U17117 : NAND3_X2 port map( A1 => n3583, A2 => n20472, A3 => n32927, ZN => 
                           n39161);
   U17122 : OAI21_X2 port map( A1 => n33437, A2 => n39083, B => n30204, ZN => 
                           n30206);
   U17132 : XOR2_X1 port map( A1 => n15904, A2 => n38082, Z => n32821);
   U17135 : XOR2_X1 port map( A1 => n23809, A2 => n37224, Z => n38082);
   U17138 : XOR2_X1 port map( A1 => n11870, A2 => n11871, Z => n13499);
   U17146 : BUF_X4 port map( I => n17095, Z => n33335);
   U17148 : OAI21_X2 port map( A1 => n10902, A2 => n31157, B => n37524, ZN => 
                           n26151);
   U17152 : XOR2_X1 port map( A1 => n27787, A2 => n27632, Z => n27527);
   U17156 : NAND2_X2 port map( A1 => n27023, A2 => n27024, ZN => n27787);
   U17167 : AOI21_X1 port map( A1 => n39584, A2 => n9743, B => n949, ZN => 
                           n5162);
   U17172 : XOR2_X1 port map( A1 => n24001, A2 => n33232, Z => n33231);
   U17175 : OAI21_X2 port map( A1 => n5591, A2 => n38085, B => n23606, ZN => 
                           n9331);
   U17180 : OR2_X1 port map( A1 => n23308, A2 => n18850, Z => n38085);
   U17182 : XOR2_X1 port map( A1 => n10767, A2 => n12003, Z => n3392);
   U17186 : XOR2_X1 port map( A1 => n16096, A2 => n7464, Z => n10767);
   U17187 : XOR2_X1 port map( A1 => n29068, A2 => n38086, Z => n21323);
   U17191 : XOR2_X1 port map( A1 => n34178, A2 => n38087, Z => n38086);
   U17195 : AND2_X1 port map( A1 => n11150, A2 => n36708, Z => n832);
   U17196 : NAND2_X2 port map( A1 => n39290, A2 => n38088, ZN => n3510);
   U17198 : NAND3_X1 port map( A1 => n224, A2 => n34374, A3 => n9193, ZN => 
                           n38088);
   U17213 : AND2_X1 port map( A1 => n2597, A2 => n39699, Z => n2595);
   U17214 : XOR2_X1 port map( A1 => n10488, A2 => n22643, Z => n10705);
   U17215 : AOI21_X2 port map( A1 => n16027, A2 => n7771, B => n347, ZN => 
                           n22643);
   U17219 : AND2_X1 port map( A1 => n28676, A2 => n28578, Z => n9951);
   U17220 : OR2_X1 port map( A1 => n9801, A2 => n11784, Z => n13004);
   U17222 : XOR2_X1 port map( A1 => n35105, A2 => n2196, Z => n9801);
   U17223 : INV_X2 port map( I => n38089, ZN => n18920);
   U17227 : XOR2_X1 port map( A1 => n18922, A2 => n18921, Z => n38089);
   U17229 : NAND2_X1 port map( A1 => n38090, A2 => n19521, ZN => n13913);
   U17231 : OAI21_X1 port map( A1 => n34401, A2 => n14483, B => n22901, ZN => 
                           n38090);
   U17234 : INV_X2 port map( I => n14502, ZN => n23201);
   U17235 : XOR2_X1 port map( A1 => n10502, A2 => n10501, Z => n14502);
   U17240 : XOR2_X1 port map( A1 => n24033, A2 => n2220, Z => n33578);
   U17241 : AOI22_X2 port map( A1 => n3821, A2 => n33885, B1 => n21892, B2 => 
                           n21489, ZN => n38091);
   U17249 : NOR2_X2 port map( A1 => n32683, A2 => n11796, ZN => n35434);
   U17251 : BUF_X4 port map( I => n5745, Z => n5675);
   U17253 : NAND2_X2 port map( A1 => n34632, A2 => n14506, ZN => n15581);
   U17255 : NOR2_X2 port map( A1 => n27484, A2 => n39296, ZN => n11041);
   U17256 : NAND2_X2 port map( A1 => n35576, A2 => n14502, ZN => n3683);
   U17257 : INV_X2 port map( I => n14833, ZN => n22128);
   U17258 : NAND2_X1 port map( A1 => n30060, A2 => n30793, ZN => n30062);
   U17259 : XOR2_X1 port map( A1 => n4828, A2 => n31965, Z => n26503);
   U17264 : OAI21_X2 port map( A1 => n3519, A2 => n3518, B => n3516, ZN => 
                           n31965);
   U17266 : BUF_X2 port map( I => n3449, Z => n38092);
   U17267 : NAND3_X2 port map( A1 => n27200, A2 => n17298, A3 => n32961, ZN => 
                           n38093);
   U17270 : NOR2_X2 port map( A1 => n22927, A2 => n8141, ZN => n20788);
   U17272 : AND2_X2 port map( A1 => n8142, A2 => n22917, Z => n8141);
   U17273 : NAND2_X2 port map( A1 => n36527, A2 => n8507, ZN => n38704);
   U17274 : INV_X2 port map( I => n21167, ZN => n8445);
   U17275 : XOR2_X1 port map( A1 => n38094, A2 => n22590, Z => n22678);
   U17276 : XOR2_X1 port map( A1 => n22529, A2 => n22528, Z => n38094);
   U17286 : XOR2_X1 port map( A1 => n7936, A2 => n38095, Z => n3705);
   U17290 : XOR2_X1 port map( A1 => n3703, A2 => n31547, Z => n38095);
   U17296 : XOR2_X1 port map( A1 => n21036, A2 => n38096, Z => n11250);
   U17297 : XOR2_X1 port map( A1 => n34531, A2 => n31320, Z => n38096);
   U17299 : XOR2_X1 port map( A1 => n3610, A2 => n15346, Z => n9205);
   U17305 : NAND3_X2 port map( A1 => n2588, A2 => n2589, A3 => n2590, ZN => 
                           n3610);
   U17306 : NAND2_X1 port map( A1 => n2765, A2 => n10463, ZN => n4865);
   U17308 : NAND2_X2 port map( A1 => n6099, A2 => n6098, ZN => n2765);
   U17310 : XOR2_X1 port map( A1 => n12741, A2 => n8940, Z => n19374);
   U17312 : NAND2_X2 port map( A1 => n11536, A2 => n11534, ZN => n8940);
   U17313 : NAND2_X2 port map( A1 => n17792, A2 => n21587, ZN => n21520);
   U17315 : NAND2_X2 port map( A1 => n38098, A2 => n6734, ZN => n29555);
   U17317 : NAND2_X1 port map( A1 => n20426, A2 => n32987, ZN => n38098);
   U17318 : NAND2_X2 port map( A1 => n3050, A2 => n27972, ZN => n28948);
   U17326 : AND2_X1 port map( A1 => n7901, A2 => n33644, Z => n18354);
   U17328 : XOR2_X1 port map( A1 => n22563, A2 => n16667, Z => n7038);
   U17331 : NOR2_X2 port map( A1 => n8947, A2 => n9485, ZN => n8744);
   U17332 : INV_X2 port map( I => n38099, ZN => n8947);
   U17333 : NAND2_X2 port map( A1 => n8948, A2 => n22222, ZN => n38099);
   U17335 : NAND3_X1 port map( A1 => n7373, A2 => n18120, A3 => n30680, ZN => 
                           n38101);
   U17342 : INV_X4 port map( I => n27064, ZN => n1221);
   U17345 : NAND3_X1 port map( A1 => n17365, A2 => n15308, A3 => n15209, ZN => 
                           n15307);
   U17349 : NAND2_X2 port map( A1 => n10883, A2 => n28685, ZN => n11030);
   U17352 : NOR3_X2 port map( A1 => n20578, A2 => n26841, A3 => n36392, ZN => 
                           n36647);
   U17357 : AND2_X1 port map( A1 => n39054, A2 => n17022, Z => n38234);
   U17360 : XOR2_X1 port map( A1 => n38103, A2 => n4397, Z => n18853);
   U17361 : XOR2_X1 port map( A1 => n5655, A2 => n6795, Z => n38103);
   U17365 : XOR2_X1 port map( A1 => n34513, A2 => n26262, Z => n13171);
   U17368 : XOR2_X1 port map( A1 => n13802, A2 => n8059, Z => n27832);
   U17369 : NAND3_X2 port map( A1 => n27040, A2 => n27039, A3 => n27041, ZN => 
                           n13802);
   U17372 : AOI21_X2 port map( A1 => n18901, A2 => n26825, B => n38104, ZN => 
                           n35036);
   U17373 : NOR2_X2 port map( A1 => n26823, A2 => n26824, ZN => n38104);
   U17387 : INV_X2 port map( I => n38106, ZN => n10261);
   U17388 : NOR2_X1 port map( A1 => n38106, A2 => n38105, ZN => n6724);
   U17389 : NAND2_X2 port map( A1 => n18686, A2 => n18685, ZN => n38106);
   U17396 : XOR2_X1 port map( A1 => n38107, A2 => n39259, Z => n38554);
   U17398 : XOR2_X1 port map( A1 => n27643, A2 => n37147, Z => n38107);
   U17399 : NAND2_X1 port map( A1 => n10210, A2 => n35869, ZN => n3430);
   U17406 : INV_X2 port map( I => n38108, ZN => n8604);
   U17408 : XNOR2_X1 port map( A1 => n18663, A2 => n33831, ZN => n38108);
   U17409 : OAI21_X2 port map( A1 => n38338, A2 => n1110, B => n25754, ZN => 
                           n9305);
   U17410 : XOR2_X1 port map( A1 => n25146, A2 => n25026, Z => n25239);
   U17412 : NAND2_X2 port map( A1 => n10876, A2 => n7495, ZN => n23303);
   U17414 : XOR2_X1 port map( A1 => n38344, A2 => n3151, Z => n5558);
   U17416 : NAND3_X2 port map( A1 => n13665, A2 => n18196, A3 => n37525, ZN => 
                           n9912);
   U17419 : NOR2_X2 port map( A1 => n22935, A2 => n8491, ZN => n8386);
   U17420 : NAND2_X1 port map( A1 => n6226, A2 => n36992, ZN => n224);
   U17425 : NAND2_X1 port map( A1 => n34068, A2 => n38114, ZN => n31200);
   U17429 : XOR2_X1 port map( A1 => n16765, A2 => n16766, Z => n24164);
   U17430 : NOR2_X2 port map( A1 => n28728, A2 => n28473, ZN => n8092);
   U17434 : NAND2_X2 port map( A1 => n27878, A2 => n4788, ZN => n28728);
   U17435 : NAND2_X2 port map( A1 => n37028, A2 => n37300, ZN => n26236);
   U17436 : XOR2_X1 port map( A1 => n22439, A2 => n22531, Z => n22640);
   U17439 : NAND2_X2 port map( A1 => n13614, A2 => n31476, ZN => n22531);
   U17445 : INV_X2 port map( I => n8430, ZN => n24789);
   U17447 : NAND2_X2 port map( A1 => n39354, A2 => n32057, ZN => n8430);
   U17451 : INV_X4 port map( I => n1755, ZN => n34389);
   U17453 : XOR2_X1 port map( A1 => n38110, A2 => n38109, Z => n2778);
   U17457 : XOR2_X1 port map( A1 => n2184, A2 => n2185, Z => n38110);
   U17460 : BUF_X4 port map( I => n8205, Z => n38609);
   U17463 : INV_X2 port map( I => n19930, ZN => n1439);
   U17471 : XOR2_X1 port map( A1 => n6848, A2 => n6796, Z => n19930);
   U17472 : NAND2_X2 port map( A1 => n30132, A2 => n18241, ZN => n19098);
   U17474 : NAND3_X2 port map( A1 => n26422, A2 => n3449, A3 => n37055, ZN => 
                           n38394);
   U17477 : XOR2_X1 port map( A1 => n36645, A2 => n6475, Z => n32537);
   U17478 : XOR2_X1 port map( A1 => n38111, A2 => n24015, Z => n24317);
   U17485 : BUF_X4 port map( I => n12237, Z => n38855);
   U17490 : NAND2_X2 port map( A1 => n17989, A2 => n17499, ZN => n34283);
   U17491 : NAND2_X2 port map( A1 => n33359, A2 => n34283, ZN => n38339);
   U17492 : INV_X2 port map( I => n27244, ZN => n34606);
   U17495 : NAND3_X2 port map( A1 => n15495, A2 => n20954, A3 => n23232, ZN => 
                           n24079);
   U17497 : AOI21_X2 port map( A1 => n20399, A2 => n1089, B => n36549, ZN => 
                           n36711);
   U17501 : NOR2_X1 port map( A1 => n33289, A2 => n19857, ZN => n8987);
   U17502 : NAND3_X2 port map( A1 => n38112, A2 => n11501, A3 => n39786, ZN => 
                           n17);
   U17508 : NAND2_X2 port map( A1 => n33603, A2 => n11375, ZN => n38112);
   U17509 : XOR2_X1 port map( A1 => n16336, A2 => n16334, Z => n33777);
   U17510 : NAND2_X2 port map( A1 => n15733, A2 => n36473, ZN => n16334);
   U17516 : AND2_X1 port map( A1 => n23102, A2 => n9677, Z => n3411);
   U17519 : OAI21_X2 port map( A1 => n15459, A2 => n5051, B => n38113, ZN => 
                           n11241);
   U17521 : NOR2_X1 port map( A1 => n38119, A2 => n23358, ZN => n38114);
   U17522 : AOI21_X2 port map( A1 => n28415, A2 => n34667, B => n35199, ZN => 
                           n38311);
   U17523 : NAND4_X2 port map( A1 => n34192, A2 => n9364, A3 => n9357, A4 => 
                           n7595, ZN => n18211);
   U17526 : NAND2_X2 port map( A1 => n26125, A2 => n4190, ZN => n39569);
   U17527 : NAND2_X1 port map( A1 => n38116, A2 => n23487, ZN => n23305);
   U17533 : OAI22_X1 port map( A1 => n23488, A2 => n1632, B1 => n32017, B2 => 
                           n37774, ZN => n38116);
   U17534 : XOR2_X1 port map( A1 => n10616, A2 => n38117, Z => n4059);
   U17535 : XOR2_X1 port map( A1 => n18600, A2 => n25214, Z => n38117);
   U17536 : XOR2_X1 port map( A1 => n8546, A2 => n38118, Z => n8544);
   U17541 : NOR2_X1 port map( A1 => n33263, A2 => n37393, ZN => n38432);
   U17544 : BUF_X4 port map( I => n29936, Z => n16224);
   U17547 : INV_X4 port map( I => n4190, ZN => n39454);
   U17548 : XOR2_X1 port map( A1 => n27749, A2 => n37812, Z => n38121);
   U17550 : XOR2_X1 port map( A1 => n19642, A2 => n27738, Z => n27502);
   U17552 : AOI22_X2 port map( A1 => n7079, A2 => n2888, B1 => n25743, B2 => 
                           n33795, ZN => n7080);
   U17553 : NAND2_X2 port map( A1 => n18213, A2 => n18215, ZN => n38122);
   U17555 : NAND3_X2 port map( A1 => n38123, A2 => n17715, A3 => n30805, ZN => 
                           n39104);
   U17556 : INV_X4 port map( I => n12306, ZN => n36234);
   U17557 : OAI21_X2 port map( A1 => n22969, A2 => n45, B => n38124, ZN => 
                           n23592);
   U17559 : OAI21_X1 port map( A1 => n35994, A2 => n6009, B => n13572, ZN => 
                           n38124);
   U17560 : NAND2_X1 port map( A1 => n34685, A2 => n25888, ZN => n25850);
   U17570 : NAND2_X2 port map( A1 => n7583, A2 => n33346, ZN => n25489);
   U17571 : NAND2_X2 port map( A1 => n38125, A2 => n34395, ZN => n14956);
   U17572 : AOI21_X2 port map( A1 => n37128, A2 => n7486, B => n38126, ZN => 
                           n38125);
   U17575 : NOR2_X2 port map( A1 => n7486, A2 => n28073, ZN => n38126);
   U17581 : NAND2_X2 port map( A1 => n4584, A2 => n4581, ZN => n10171);
   U17585 : NOR2_X1 port map( A1 => n21840, A2 => n21903, ZN => n21624);
   U17587 : OR2_X1 port map( A1 => n17217, A2 => n856, Z => n9061);
   U17592 : AND2_X1 port map( A1 => n8849, A2 => n8850, Z => n38127);
   U17593 : AOI21_X2 port map( A1 => n24832, A2 => n24573, B => n38128, ZN => 
                           n16864);
   U17594 : OAI21_X2 port map( A1 => n16208, A2 => n24832, B => n24574, ZN => 
                           n38128);
   U17595 : XNOR2_X1 port map( A1 => n17310, A2 => n22552, ZN => n6630);
   U17596 : OAI21_X2 port map( A1 => n6582, A2 => n36946, B => n22159, ZN => 
                           n22552);
   U17599 : AOI21_X2 port map( A1 => n38129, A2 => n19734, B => n19962, ZN => 
                           n2243);
   U17600 : NAND2_X1 port map( A1 => n8229, A2 => n38429, ZN => n39522);
   U17601 : NOR2_X2 port map( A1 => n16733, A2 => n38130, ZN => n16732);
   U17602 : NAND2_X2 port map( A1 => n26870, A2 => n7975, ZN => n27006);
   U17605 : XOR2_X1 port map( A1 => n36778, A2 => n22580, Z => n2471);
   U17607 : XOR2_X1 port map( A1 => n20454, A2 => n27687, Z => n27490);
   U17608 : XOR2_X1 port map( A1 => n11399, A2 => n32505, Z => n16425);
   U17610 : NAND2_X2 port map( A1 => n19435, A2 => n20157, ZN => n11526);
   U17614 : XOR2_X1 port map( A1 => n27758, A2 => n27534, Z => n3557);
   U17620 : NAND2_X2 port map( A1 => n13400, A2 => n35790, ZN => n27758);
   U17622 : XOR2_X1 port map( A1 => n27667, A2 => n31061, Z => n12304);
   U17623 : NAND2_X2 port map( A1 => n15768, A2 => n37096, ZN => n29361);
   U17640 : XOR2_X1 port map( A1 => n22748, A2 => n22747, Z => n5338);
   U17642 : XOR2_X1 port map( A1 => n16804, A2 => n16805, Z => n18186);
   U17643 : XOR2_X1 port map( A1 => n27541, A2 => n34986, Z => n16805);
   U17645 : OR2_X1 port map( A1 => n25836, A2 => n19580, Z => n18214);
   U17647 : AOI22_X2 port map( A1 => n5164, A2 => n927, B1 => n26090, B2 => 
                           n37239, ZN => n38131);
   U17650 : XOR2_X1 port map( A1 => n1886, A2 => n1883, Z => n10938);
   U17652 : NAND2_X2 port map( A1 => n25975, A2 => n6056, ZN => n15524);
   U17654 : NOR3_X2 port map( A1 => n10882, A2 => n1548, A3 => n31780, ZN => 
                           n32011);
   U17656 : NAND2_X2 port map( A1 => n38132, A2 => n39622, ZN => n25836);
   U17657 : XOR2_X1 port map( A1 => n2782, A2 => n38181, Z => n38133);
   U17661 : NAND2_X2 port map( A1 => n24740, A2 => n24821, ZN => n35785);
   U17662 : OAI21_X2 port map( A1 => n14167, A2 => n24820, B => n14166, ZN => 
                           n24740);
   U17663 : BUF_X4 port map( I => n9920, Z => n9321);
   U17666 : NAND2_X2 port map( A1 => n28748, A2 => n9917, ZN => n28623);
   U17670 : NAND2_X2 port map( A1 => n8535, A2 => n8534, ZN => n27633);
   U17671 : NAND2_X2 port map( A1 => n23505, A2 => n20276, ZN => n23596);
   U17672 : NOR2_X2 port map( A1 => n23051, A2 => n4565, ZN => n35932);
   U17675 : OR2_X1 port map( A1 => n13717, A2 => n26001, Z => n2657);
   U17683 : XOR2_X1 port map( A1 => n38134, A2 => n30126, Z => Ciphertext(166))
                           ;
   U17685 : NAND3_X2 port map( A1 => n36005, A2 => n36420, A3 => n9261, ZN => 
                           n38134);
   U17687 : BUF_X4 port map( I => n26459, Z => n26909);
   U17688 : INV_X2 port map( I => n38135, ZN => n39815);
   U17689 : XOR2_X1 port map( A1 => n8567, A2 => n8565, Z => n38135);
   U17694 : XOR2_X1 port map( A1 => n38136, A2 => n1769, Z => n32985);
   U17700 : BUF_X2 port map( I => n17890, Z => n38137);
   U17701 : NOR2_X2 port map( A1 => n31264, A2 => n37102, ZN => n38138);
   U17705 : INV_X2 port map( I => n22510, ZN => n22778);
   U17713 : NAND2_X2 port map( A1 => n20256, A2 => n33655, ZN => n22510);
   U17718 : AOI22_X1 port map( A1 => n30098, A2 => n2489, B1 => n2484, B2 => 
                           n35175, ZN => n36182);
   U17719 : NAND2_X2 port map( A1 => n36736, A2 => n8730, ZN => n38653);
   U17722 : XOR2_X1 port map( A1 => n15305, A2 => n38139, Z => n20883);
   U17725 : XOR2_X1 port map( A1 => n15303, A2 => n15304, Z => n38139);
   U17726 : XOR2_X1 port map( A1 => n23973, A2 => n18175, Z => n23937);
   U17727 : NAND2_X2 port map( A1 => n39506, A2 => n32487, ZN => n23973);
   U17729 : XOR2_X1 port map( A1 => n35878, A2 => n22727, Z => n13561);
   U17734 : INV_X1 port map( I => n38512, ZN => n35374);
   U17738 : OAI21_X1 port map( A1 => n33104, A2 => n12146, B => n2091, ZN => 
                           n36444);
   U17739 : INV_X2 port map( I => n17653, ZN => n2848);
   U17740 : NAND2_X2 port map( A1 => n32391, A2 => n5282, ZN => n17891);
   U17741 : NOR3_X2 port map( A1 => n35313, A2 => n31661, A3 => n36885, ZN => 
                           n32054);
   U17753 : NAND3_X2 port map( A1 => n20498, A2 => n29722, A3 => n17708, ZN => 
                           n29714);
   U17754 : AND2_X1 port map( A1 => n30184, A2 => n17996, Z => n12301);
   U17762 : NAND2_X2 port map( A1 => n23255, A2 => n33702, ZN => n38175);
   U17763 : INV_X2 port map( I => n25813, ZN => n1014);
   U17765 : OAI21_X2 port map( A1 => n38775, A2 => n35580, B => n38774, ZN => 
                           n26650);
   U17773 : NOR2_X2 port map( A1 => n15623, A2 => n3983, ZN => n36224);
   U17774 : AOI22_X2 port map( A1 => n26132, A2 => n1014, B1 => n6749, B2 => 
                           n25936, ZN => n39625);
   U17775 : INV_X2 port map( I => n26459, ZN => n26719);
   U17782 : NAND2_X2 port map( A1 => n988, A2 => n27894, ZN => n13955);
   U17793 : INV_X2 port map( I => n8412, ZN => n27440);
   U17796 : AOI21_X2 port map( A1 => n2868, A2 => n28224, B => n28229, ZN => 
                           n15571);
   U17797 : OAI22_X2 port map( A1 => n33001, A2 => n32948, B1 => n36711, B2 => 
                           n38092, ZN => n38402);
   U17801 : BUF_X4 port map( I => n38402, Z => n32926);
   U17804 : NAND2_X2 port map( A1 => n2740, A2 => n12443, ZN => n12488);
   U17805 : NAND2_X2 port map( A1 => n691, A2 => n29555, ZN => n29547);
   U17806 : OR2_X1 port map( A1 => n29437, A2 => n29438, Z => n18495);
   U17814 : INV_X4 port map( I => n13366, ZN => n28213);
   U17815 : OAI21_X1 port map( A1 => n8307, A2 => n1198, B => n38804, ZN => 
                           n33161);
   U17818 : AOI22_X2 port map( A1 => n12478, A2 => n7866, B1 => n1531, B2 => 
                           n25692, ZN => n8223);
   U17819 : AOI22_X2 port map( A1 => n8965, A2 => n38119, B1 => n8757, B2 => 
                           n23358, ZN => n6517);
   U17820 : NAND2_X2 port map( A1 => n8407, A2 => n25782, ZN => n35786);
   U17822 : INV_X2 port map( I => n30257, ZN => n30258);
   U17828 : INV_X2 port map( I => n23540, ZN => n10495);
   U17829 : NAND2_X1 port map( A1 => n38266, A2 => n36654, ZN => n22825);
   U17832 : NAND2_X2 port map( A1 => n945, A2 => n27233, ZN => n7471);
   U17833 : AOI21_X2 port map( A1 => n986, A2 => n20977, B => n38443, ZN => 
                           n8993);
   U17835 : NAND2_X2 port map( A1 => n34740, A2 => n34739, ZN => n34738);
   U17836 : NOR2_X2 port map( A1 => n20010, A2 => n28279, ZN => n30773);
   U17837 : AOI21_X2 port map( A1 => n38404, A2 => n38702, B => n2597, ZN => 
                           n30550);
   U17838 : NOR3_X2 port map( A1 => n310, A2 => n16461, A3 => n28200, ZN => 
                           n35309);
   U17840 : NAND2_X2 port map( A1 => n25692, A2 => n12478, ZN => n12382);
   U17847 : NAND2_X2 port map( A1 => n31486, A2 => n39768, ZN => n38143);
   U17848 : OAI21_X1 port map( A1 => n6204, A2 => n1407, B => n31444, ZN => 
                           n29194);
   U17857 : BUF_X4 port map( I => n28231, Z => n19366);
   U17858 : INV_X2 port map( I => n29998, ZN => n29949);
   U17859 : OAI22_X2 port map( A1 => n30365, A2 => n1093, B1 => n38824, B2 => 
                           n38120, ZN => n18023);
   U17861 : INV_X2 port map( I => n29781, ZN => n1408);
   U17863 : NAND2_X1 port map( A1 => n6831, A2 => n36375, ZN => n38632);
   U17866 : NAND2_X2 port map( A1 => n13151, A2 => n36791, ZN => n13372);
   U17868 : OR2_X1 port map( A1 => n5881, A2 => n5884, Z => n38140);
   U17870 : INV_X1 port map( I => n25246, ZN => n38895);
   U17872 : INV_X1 port map( I => n39793, ZN => n25848);
   U17876 : NOR2_X1 port map( A1 => n20157, A2 => n32977, ZN => n30370);
   U17882 : NOR3_X1 port map( A1 => n32977, A2 => n28049, A3 => n20157, ZN => 
                           n10166);
   U17884 : NAND2_X1 port map( A1 => n36391, A2 => n14601, ZN => n12986);
   U17893 : INV_X1 port map( I => n29559, ZN => n39003);
   U17895 : AOI21_X1 port map( A1 => n27416, A2 => n19564, B => n27110, ZN => 
                           n27111);
   U17896 : NOR2_X1 port map( A1 => n28131, A2 => n2868, ZN => n15568);
   U17900 : CLKBUF_X4 port map( I => n20522, Z => n33784);
   U17902 : NAND2_X1 port map( A1 => n30241, A2 => n20525, ZN => n31237);
   U17903 : NAND2_X1 port map( A1 => n859, A2 => n26935, ZN => n13777);
   U17910 : NAND2_X1 port map( A1 => n29354, A2 => n29422, ZN => n6865);
   U17914 : CLKBUF_X4 port map( I => n33961, Z => n2782);
   U17915 : INV_X1 port map( I => n27802, ZN => n1457);
   U17917 : NOR2_X1 port map( A1 => n19475, A2 => n20160, ZN => n38142);
   U17918 : INV_X1 port map( I => n29204, ZN => n15601);
   U17920 : NAND2_X1 port map( A1 => n25962, A2 => n16407, ZN => n26027);
   U17922 : NAND3_X1 port map( A1 => n27866, A2 => n19657, A3 => n9553, ZN => 
                           n27685);
   U17932 : OR2_X1 port map( A1 => n29869, A2 => n773, Z => n5973);
   U17933 : NAND2_X1 port map( A1 => n38506, A2 => n14030, ZN => n38145);
   U17934 : NOR2_X1 port map( A1 => n28142, A2 => n20184, ZN => n20500);
   U17935 : CLKBUF_X4 port map( I => n28473, Z => n5396);
   U17936 : CLKBUF_X4 port map( I => n17777, Z => n11676);
   U17945 : NAND2_X1 port map( A1 => n9802, A2 => n19580, ZN => n30957);
   U17948 : NAND2_X1 port map( A1 => n29701, A2 => n29700, ZN => n16385);
   U17951 : OAI21_X1 port map( A1 => n29699, A2 => n29700, B => n29698, ZN => 
                           n28513);
   U17953 : NAND2_X1 port map( A1 => n30034, A2 => n30024, ZN => n10942);
   U17954 : INV_X2 port map( I => n4879, ZN => n29843);
   U17955 : NOR2_X1 port map( A1 => n4879, A2 => n20793, ZN => n3379);
   U17958 : OR2_X1 port map( A1 => n39126, A2 => n32822, Z => n5863);
   U17961 : NOR2_X1 port map( A1 => n16154, A2 => n28143, ZN => n7255);
   U17962 : AOI22_X1 port map( A1 => n25420, A2 => n18031, B1 => n12381, B2 => 
                           n13166, ZN => n38628);
   U17967 : INV_X1 port map( I => n21546, ZN => n1692);
   U17972 : INV_X2 port map( I => n19696, ZN => n19452);
   U17975 : BUF_X2 port map( I => n4382, Z => n32385);
   U17976 : NOR2_X1 port map( A1 => n39334, A2 => n28738, ZN => n28743);
   U17988 : INV_X1 port map( I => n28286, ZN => n28161);
   U17992 : NAND2_X1 port map( A1 => n31143, A2 => n39731, ZN => n38148);
   U17993 : NAND3_X1 port map( A1 => n29712, A2 => n29719, A3 => n14337, ZN => 
                           n29716);
   U17994 : OR2_X2 port map( A1 => n9118, A2 => n26459, Z => n26927);
   U17995 : AND2_X1 port map( A1 => n33960, A2 => n15774, Z => n33185);
   U17997 : CLKBUF_X1 port map( I => n7464, Z => n34492);
   U18000 : NOR2_X1 port map( A1 => n24169, A2 => n24396, ZN => n23844);
   U18001 : NAND3_X1 port map( A1 => n1142, A2 => n11307, A3 => n20782, ZN => 
                           n23086);
   U18002 : NOR2_X1 port map( A1 => n25942, A2 => n6579, ZN => n9714);
   U18004 : OAI21_X1 port map( A1 => n10800, A2 => n35690, B => n10046, ZN => 
                           n10799);
   U18006 : INV_X1 port map( I => n36571, ZN => n34482);
   U18007 : INV_X2 port map( I => n26780, ZN => n26948);
   U18010 : NOR2_X1 port map( A1 => n28478, A2 => n1196, ZN => n28479);
   U18011 : NAND2_X1 port map( A1 => n1414, A2 => n1196, ZN => n33229);
   U18014 : OAI21_X2 port map( A1 => n20050, A2 => n20051, B => n20049, ZN => 
                           n38149);
   U18026 : OAI21_X1 port map( A1 => n20050, A2 => n20051, B => n20049, ZN => 
                           n20210);
   U18044 : OR2_X1 port map( A1 => n24536, A2 => n7705, Z => n19532);
   U18053 : AND3_X1 port map( A1 => n19398, A2 => n7705, A3 => n25683, Z => 
                           n34025);
   U18054 : NAND2_X1 port map( A1 => n29375, A2 => n37100, ZN => n19244);
   U18055 : NAND2_X1 port map( A1 => n29310, A2 => n29384, ZN => n36994);
   U18056 : NAND2_X1 port map( A1 => n35508, A2 => n36133, ZN => n25534);
   U18057 : NOR2_X1 port map( A1 => n32366, A2 => n1294, ZN => n8214);
   U18058 : NAND2_X1 port map( A1 => n11491, A2 => n11492, ZN => n38150);
   U18059 : INV_X1 port map( I => n36523, ZN => n36050);
   U18063 : INV_X1 port map( I => n7106, ZN => n31425);
   U18064 : NAND3_X1 port map( A1 => n7106, A2 => n12415, A3 => n26967, ZN => 
                           n6797);
   U18066 : OR2_X1 port map( A1 => n14387, A2 => n30217, Z => n36739);
   U18076 : INV_X2 port map( I => n33963, ZN => n10569);
   U18079 : NAND2_X1 port map( A1 => n13370, A2 => n14856, ZN => n13834);
   U18080 : OAI21_X1 port map( A1 => n27927, A2 => n27926, B => n36414, ZN => 
                           n8910);
   U18081 : OR2_X1 port map( A1 => n12371, A2 => n12372, Z => n38151);
   U18083 : NAND2_X1 port map( A1 => n11787, A2 => n11785, ZN => n35029);
   U18084 : OAI21_X2 port map( A1 => n27258, A2 => n27257, B => n27256, ZN => 
                           n38152);
   U18085 : OAI21_X1 port map( A1 => n27258, A2 => n27257, B => n27256, ZN => 
                           n38153);
   U18087 : OAI21_X1 port map( A1 => n27258, A2 => n27257, B => n27256, ZN => 
                           n27717);
   U18089 : NOR2_X2 port map( A1 => n32697, A2 => n7588, ZN => n27257);
   U18093 : CLKBUF_X4 port map( I => n26888, Z => n27337);
   U18108 : AND2_X1 port map( A1 => n2792, A2 => n29810, Z => n14009);
   U18111 : NAND2_X2 port map( A1 => n33563, A2 => n21164, ZN => n38154);
   U18114 : INV_X1 port map( I => n18908, ZN => n2113);
   U18117 : INV_X2 port map( I => n378, ZN => n14793);
   U18120 : NAND2_X1 port map( A1 => n378, A2 => n36922, ZN => n36815);
   U18121 : NOR2_X1 port map( A1 => n36922, A2 => n378, ZN => n30644);
   U18122 : NAND2_X1 port map( A1 => n378, A2 => n33293, ZN => n7404);
   U18124 : OAI21_X1 port map( A1 => n10338, A2 => n10524, B => n8311, ZN => 
                           n26270);
   U18135 : NOR2_X1 port map( A1 => n27141, A2 => n10338, ZN => n38494);
   U18136 : INV_X2 port map( I => n8000, ZN => n10338);
   U18137 : OR3_X1 port map( A1 => n8960, A2 => n27624, A3 => n16576, Z => 
                           n7983);
   U18138 : NOR2_X1 port map( A1 => n32186, A2 => n16576, ZN => n28422);
   U18139 : OAI21_X1 port map( A1 => n28328, A2 => n28327, B => n39423, ZN => 
                           n38970);
   U18144 : NOR2_X1 port map( A1 => n39423, A2 => n39422, ZN => n35548);
   U18145 : INV_X1 port map( I => n38461, ZN => n5334);
   U18148 : NAND2_X1 port map( A1 => n34386, A2 => n9823, ZN => n38623);
   U18162 : INV_X1 port map( I => n15625, ZN => n25277);
   U18165 : OR2_X2 port map( A1 => n37079, A2 => n8395, Z => n28043);
   U18168 : NOR2_X1 port map( A1 => n27250, A2 => n33503, ZN => n11854);
   U18169 : AOI21_X1 port map( A1 => n13907, A2 => n310, B => n13906, ZN => 
                           n13905);
   U18175 : INV_X1 port map( I => n35705, ZN => n1605);
   U18182 : NAND2_X1 port map( A1 => n609, A2 => n35705, ZN => n24451);
   U18185 : OR2_X1 port map( A1 => n16459, A2 => n35705, Z => n6933);
   U18187 : INV_X1 port map( I => n29336, ZN => n38156);
   U18191 : AND2_X1 port map( A1 => n32790, A2 => n14858, Z => n29328);
   U18197 : CLKBUF_X12 port map( I => n29336, Z => n32790);
   U18198 : OAI21_X1 port map( A1 => n19669, A2 => n20691, B => n27498, ZN => 
                           n16856);
   U18200 : OAI21_X1 port map( A1 => n6975, A2 => n27027, B => n27251, ZN => 
                           n33160);
   U18202 : NAND2_X1 port map( A1 => n13088, A2 => n26988, ZN => n6261);
   U18207 : NAND2_X1 port map( A1 => n29800, A2 => n29799, ZN => n5145);
   U18208 : NOR2_X1 port map( A1 => n29800, A2 => n3614, ZN => n39062);
   U18214 : NAND2_X1 port map( A1 => n35273, A2 => n29616, ZN => n29624);
   U18216 : NAND3_X2 port map( A1 => n8031, A2 => n37728, A3 => n8030, ZN => 
                           n10978);
   U18219 : CLKBUF_X4 port map( I => n833, Z => n7284);
   U18220 : XNOR2_X1 port map( A1 => n23832, A2 => n24050, ZN => n17140);
   U18231 : XOR2_X1 port map( A1 => n2805, A2 => n38157, Z => n36380);
   U18246 : XOR2_X1 port map( A1 => n23887, A2 => n678, Z => n38157);
   U18248 : NOR2_X1 port map( A1 => n28163, A2 => n5988, ZN => n885);
   U18249 : BUF_X2 port map( I => n28163, Z => n32705);
   U18251 : AOI21_X1 port map( A1 => n28163, A2 => n16363, B => n27979, ZN => 
                           n35931);
   U18252 : CLKBUF_X1 port map( I => n30184, Z => n31846);
   U18256 : AOI21_X1 port map( A1 => n38683, A2 => n15317, B => n26901, ZN => 
                           n5589);
   U18258 : NAND3_X1 port map( A1 => n26903, A2 => n26901, A3 => n11616, ZN => 
                           n34843);
   U18259 : NAND2_X1 port map( A1 => n34000, A2 => n1402, ZN => n39312);
   U18260 : NOR2_X1 port map( A1 => n39313, A2 => n34000, ZN => n32335);
   U18261 : NAND2_X1 port map( A1 => n8519, A2 => n22196, ZN => n3435);
   U18266 : OAI21_X1 port map( A1 => n5509, A2 => n13851, B => n13322, ZN => 
                           n13321);
   U18270 : NAND2_X1 port map( A1 => n15963, A2 => n3988, ZN => n35030);
   U18273 : AOI22_X1 port map( A1 => n33139, A2 => n9627, B1 => n29333, B2 => 
                           n29340, ZN => n31801);
   U18279 : INV_X2 port map( I => n12543, ZN => n4950);
   U18282 : NOR2_X1 port map( A1 => n26841, A2 => n36392, ZN => n38798);
   U18284 : CLKBUF_X4 port map( I => n20595, Z => n1548);
   U18287 : OAI22_X1 port map( A1 => n19452, A2 => n1548, B1 => n16836, B2 => 
                           n16246, ZN => n25402);
   U18304 : OAI21_X1 port map( A1 => n1548, A2 => n953, B => n16246, ZN => 
                           n3877);
   U18305 : NAND2_X2 port map( A1 => n32755, A2 => n38333, ZN => n38158);
   U18309 : NOR2_X2 port map( A1 => n4941, A2 => n30837, ZN => n38159);
   U18311 : NAND2_X1 port map( A1 => n32755, A2 => n38333, ZN => n38964);
   U18312 : NAND2_X2 port map( A1 => n32756, A2 => n32757, ZN => n32755);
   U18315 : CLKBUF_X12 port map( I => n20883, Z => n10346);
   U18318 : NOR2_X1 port map( A1 => n13442, A2 => n35179, ZN => n29566);
   U18324 : INV_X1 port map( I => n5031, ZN => n26117);
   U18329 : NAND2_X1 port map( A1 => n29889, A2 => n29888, ZN => n11787);
   U18330 : NAND2_X1 port map( A1 => n26905, A2 => n26564, ZN => n15880);
   U18335 : NAND3_X1 port map( A1 => n30858, A2 => n28444, A3 => n30857, ZN => 
                           n27972);
   U18339 : NOR2_X1 port map( A1 => n10746, A2 => n2456, ZN => n9064);
   U18340 : NAND2_X1 port map( A1 => n38871, A2 => n13890, ZN => n38160);
   U18345 : AND2_X1 port map( A1 => n26048, A2 => n26019, Z => n26050);
   U18357 : NOR2_X1 port map( A1 => n18281, A2 => n7905, ZN => n28705);
   U18360 : NOR2_X1 port map( A1 => n39019, A2 => n17286, ZN => n29877);
   U18362 : NAND4_X1 port map( A1 => n1560, A2 => n11601, A3 => n14874, A4 => 
                           n24754, ZN => n11605);
   U18363 : OAI21_X1 port map( A1 => n3631, A2 => n2121, B => n38784, ZN => 
                           n28923);
   U18364 : NAND2_X1 port map( A1 => n9328, A2 => n9327, ZN => n38162);
   U18370 : NAND2_X2 port map( A1 => n27906, A2 => n9897, ZN => n9327);
   U18372 : OR2_X2 port map( A1 => n139, A2 => n32925, Z => n38163);
   U18376 : OR2_X2 port map( A1 => n139, A2 => n32925, Z => n38164);
   U18377 : INV_X1 port map( I => n26591, ZN => n15676);
   U18378 : NAND2_X1 port map( A1 => n33200, A2 => n33199, ZN => n27890);
   U18380 : NOR2_X1 port map( A1 => n6892, A2 => n28609, ZN => n28335);
   U18381 : OAI21_X1 port map( A1 => n12238, A2 => n12611, B => n28609, ZN => 
                           n35574);
   U18382 : NAND3_X1 port map( A1 => n178, A2 => n25670, A3 => n18164, ZN => 
                           n10936);
   U18383 : NOR2_X1 port map( A1 => n1066, A2 => n16559, ZN => n35997);
   U18385 : INV_X1 port map( I => n9246, ZN => n8045);
   U18389 : NAND2_X1 port map( A1 => n12943, A2 => n9839, ZN => n29365);
   U18393 : INV_X2 port map( I => n9839, ZN => n13981);
   U18399 : AOI21_X2 port map( A1 => n28623, A2 => n19161, B => n977, ZN => 
                           n13656);
   U18400 : INV_X2 port map( I => n28745, ZN => n977);
   U18404 : INV_X1 port map( I => n36275, ZN => n18190);
   U18407 : INV_X1 port map( I => n11939, ZN => n31912);
   U18408 : OR3_X1 port map( A1 => n968, A2 => n939, A3 => n3462, Z => n30401);
   U18413 : CLKBUF_X4 port map( I => n28130, Z => n2868);
   U18418 : INV_X1 port map( I => n39456, ZN => n34479);
   U18421 : OAI21_X1 port map( A1 => n21724, A2 => n4925, B => n4924, ZN => 
                           n21725);
   U18425 : INV_X1 port map( I => n12537, ZN => n10058);
   U18426 : NOR2_X1 port map( A1 => n11443, A2 => n27010, ZN => n32490);
   U18427 : INV_X2 port map( I => n14557, ZN => n30047);
   U18428 : CLKBUF_X4 port map( I => n14557, Z => n36850);
   U18437 : AOI21_X2 port map( A1 => n3798, A2 => n3799, B => n33519, ZN => 
                           n38165);
   U18443 : NAND2_X2 port map( A1 => n977, A2 => n28746, ZN => n3798);
   U18454 : INV_X2 port map( I => n29777, ZN => n39313);
   U18457 : INV_X2 port map( I => n28398, ZN => n16691);
   U18460 : NAND2_X1 port map( A1 => n28398, A2 => n16303, ZN => n16304);
   U18463 : NAND2_X1 port map( A1 => n28398, A2 => n28755, ZN => n27909);
   U18465 : OR2_X1 port map( A1 => n16039, A2 => n15466, Z => n21617);
   U18466 : NAND2_X1 port map( A1 => n28422, A2 => n27624, ZN => n31087);
   U18469 : INV_X1 port map( I => n16324, ZN => n5290);
   U18470 : XNOR2_X1 port map( A1 => n36254, A2 => n36255, ZN => n38167);
   U18474 : NAND2_X1 port map( A1 => n3944, A2 => n14448, ZN => n38727);
   U18475 : NAND2_X1 port map( A1 => n12488, A2 => n982, ZN => n3981);
   U18477 : NAND2_X1 port map( A1 => n12488, A2 => n2262, ZN => n12487);
   U18494 : OAI21_X1 port map( A1 => n33107, A2 => n33106, B => n30953, ZN => 
                           n18624);
   U18496 : CLKBUF_X12 port map( I => n2147, Z => n30953);
   U18498 : NAND2_X1 port map( A1 => n8314, A2 => n36385, ZN => n1845);
   U18500 : OR2_X2 port map( A1 => n26779, A2 => n20063, Z => n26848);
   U18501 : NAND2_X1 port map( A1 => n34857, A2 => n39140, ZN => n39822);
   U18502 : NOR2_X1 port map( A1 => n27963, A2 => n28050, ZN => n10515);
   U18503 : NAND2_X1 port map( A1 => n37754, A2 => n28279, ZN => n27621);
   U18504 : INV_X1 port map( I => n12081, ZN => n1397);
   U18508 : XOR2_X1 port map( A1 => n38169, A2 => n38170, Z => n34251);
   U18509 : XNOR2_X1 port map( A1 => n27773, A2 => n19561, ZN => n38169);
   U18511 : XOR2_X1 port map( A1 => n9315, A2 => n15273, Z => n38170);
   U18512 : NOR2_X1 port map( A1 => n773, A2 => n1063, ZN => n34858);
   U18520 : OR2_X1 port map( A1 => n13758, A2 => n26219, Z => n14862);
   U18522 : NAND2_X1 port map( A1 => n27412, A2 => n36200, ZN => n6353);
   U18524 : NOR2_X1 port map( A1 => n21401, A2 => n21644, ZN => n21720);
   U18530 : AOI21_X1 port map( A1 => n21401, A2 => n32704, B => n21909, ZN => 
                           n13239);
   U18534 : NAND2_X1 port map( A1 => n20120, A2 => n2752, ZN => n38774);
   U18535 : BUF_X2 port map( I => n20120, Z => n35580);
   U18539 : NAND2_X1 port map( A1 => n15594, A2 => n20120, ZN => n26748);
   U18542 : INV_X1 port map( I => n20120, ZN => n8478);
   U18545 : AOI22_X1 port map( A1 => n29796, A2 => n36096, B1 => n29798, B2 => 
                           n29797, ZN => n36808);
   U18548 : AOI22_X1 port map( A1 => n29784, A2 => n29783, B1 => n29798, B2 => 
                           n29789, ZN => n39278);
   U18552 : OR3_X2 port map( A1 => n30195, A2 => n35551, A3 => n4083, Z => 
                           n35329);
   U18555 : NAND2_X1 port map( A1 => n21759, A2 => n21545, ZN => n21549);
   U18556 : OAI21_X1 port map( A1 => n17997, A2 => n31846, B => n2466, ZN => 
                           n2465);
   U18560 : OR2_X2 port map( A1 => n37896, A2 => n12519, Z => n24401);
   U18563 : CLKBUF_X4 port map( I => n29452, Z => n505);
   U18565 : INV_X2 port map( I => n29869, ZN => n972);
   U18576 : AOI21_X1 port map( A1 => n36225, A2 => n19476, B => n11826, ZN => 
                           n2769);
   U18587 : AOI21_X1 port map( A1 => n1802, A2 => n21017, B => n33945, ZN => 
                           n38171);
   U18589 : AOI21_X1 port map( A1 => n1802, A2 => n21017, B => n33945, ZN => 
                           n35317);
   U18593 : NOR2_X1 port map( A1 => n37619, A2 => n12537, ZN => n13403);
   U18594 : NAND2_X1 port map( A1 => n35745, A2 => n15616, ZN => n31146);
   U18603 : NAND3_X1 port map( A1 => n17661, A2 => n27218, A3 => n15616, ZN => 
                           n4948);
   U18606 : NOR2_X1 port map( A1 => n4649, A2 => n1209, ZN => n10084);
   U18612 : NOR2_X1 port map( A1 => n22295, A2 => n5061, ZN => n5127);
   U18613 : INV_X1 port map( I => n8988, ZN => n38853);
   U18617 : INV_X1 port map( I => n12707, ZN => n14128);
   U18619 : CLKBUF_X12 port map( I => n39528, Z => n38951);
   U18634 : AOI21_X1 port map( A1 => n37075, A2 => n8253, B => n33662, ZN => 
                           n2381);
   U18635 : AOI21_X1 port map( A1 => n33082, A2 => n22907, B => n22906, ZN => 
                           n23391);
   U18641 : NAND2_X1 port map( A1 => n6691, A2 => n14560, ZN => n32042);
   U18646 : INV_X1 port map( I => n28484, ZN => n28391);
   U18652 : NAND2_X1 port map( A1 => n11089, A2 => n11087, ZN => n38174);
   U18654 : INV_X1 port map( I => n11330, ZN => n28609);
   U18659 : INV_X1 port map( I => n32623, ZN => n3328);
   U18661 : NAND2_X1 port map( A1 => n30244, A2 => n30245, ZN => n30246);
   U18668 : NOR2_X1 port map( A1 => n30245, A2 => n39187, ZN => n10977);
   U18669 : NAND2_X1 port map( A1 => n29815, A2 => n8677, ZN => n29774);
   U18670 : NAND2_X1 port map( A1 => n4520, A2 => n18601, ZN => n4519);
   U18671 : INV_X2 port map( I => n5457, ZN => n18601);
   U18677 : INV_X1 port map( I => n25700, ZN => n31895);
   U18681 : NAND2_X1 port map( A1 => n1944, A2 => n7454, ZN => n28359);
   U18684 : NAND2_X1 port map( A1 => n20830, A2 => n29458, ZN => n20427);
   U18685 : OAI21_X1 port map( A1 => n10648, A2 => n10988, B => n17653, ZN => 
                           n10645);
   U18687 : OR2_X2 port map( A1 => n19543, A2 => n20778, Z => n6349);
   U18688 : CLKBUF_X4 port map( I => n33086, Z => n38337);
   U18689 : NAND2_X1 port map( A1 => n28563, A2 => n1197, ZN => n38856);
   U18690 : INV_X1 port map( I => n1197, ZN => n38858);
   U18696 : AND2_X2 port map( A1 => n2153, A2 => n33748, Z => n14250);
   U18698 : NAND2_X2 port map( A1 => n8145, A2 => n38651, ZN => n23255);
   U18702 : INV_X2 port map( I => n17598, ZN => n9553);
   U18703 : NOR2_X2 port map( A1 => n33752, A2 => n6589, ZN => n38176);
   U18706 : XOR2_X1 port map( A1 => n9989, A2 => n26481, Z => n38177);
   U18715 : XOR2_X1 port map( A1 => n6630, A2 => n17513, Z => n38179);
   U18718 : OR3_X2 port map( A1 => n13300, A2 => n38749, A3 => n24515, Z => 
                           n24777);
   U18720 : OR2_X2 port map( A1 => n37245, A2 => n34977, Z => n30412);
   U18722 : NAND2_X1 port map( A1 => n8262, A2 => n7542, ZN => n26647);
   U18723 : NAND2_X1 port map( A1 => n1107, A2 => n25860, ZN => n25708);
   U18727 : OAI21_X2 port map( A1 => n4429, A2 => n4428, B => n4076, ZN => 
                           n38181);
   U18728 : NAND2_X1 port map( A1 => n7497, A2 => n20351, ZN => n22235);
   U18730 : OR2_X2 port map( A1 => n4291, A2 => n8544, Z => n23106);
   U18734 : NAND2_X1 port map( A1 => n31234, A2 => n23349, ZN => n2692);
   U18738 : NAND2_X1 port map( A1 => n19332, A2 => n20995, ZN => n26709);
   U18742 : INV_X1 port map( I => n2273, ZN => n23317);
   U18743 : BUF_X2 port map( I => n29137, Z => n30856);
   U18751 : NAND3_X1 port map( A1 => n15327, A2 => n15328, A3 => n30057, ZN => 
                           n32668);
   U18753 : INV_X1 port map( I => n29236, ZN => n38945);
   U18757 : NAND2_X1 port map( A1 => n39300, A2 => n20276, ZN => n39299);
   U18758 : INV_X2 port map( I => n20276, ZN => n23504);
   U18777 : NOR2_X1 port map( A1 => n8190, A2 => n20276, ZN => n8212);
   U18794 : NAND2_X1 port map( A1 => n33455, A2 => n39477, ZN => n26634);
   U18796 : INV_X1 port map( I => n16080, ZN => n8305);
   U18797 : NAND2_X1 port map( A1 => n3513, A2 => n34717, ZN => n4033);
   U18798 : NOR2_X1 port map( A1 => n1224, A2 => n34717, ZN => n3514);
   U18804 : INV_X1 port map( I => n25558, ZN => n38183);
   U18813 : NAND3_X1 port map( A1 => n24763, A2 => n1269, A3 => n39098, ZN => 
                           n24767);
   U18816 : AND2_X2 port map( A1 => n199, A2 => n198, Z => n38184);
   U18822 : OR2_X2 port map( A1 => n15135, A2 => n2722, Z => n27584);
   U18825 : NAND2_X1 port map( A1 => n15135, A2 => n11020, ZN => n36222);
   U18829 : NOR2_X1 port map( A1 => n6218, A2 => n36539, ZN => n8268);
   U18837 : NOR3_X1 port map( A1 => n18907, A2 => n18402, A3 => n24203, ZN => 
                           n34673);
   U18841 : NAND2_X1 port map( A1 => n18907, A2 => n18402, ZN => n39659);
   U18855 : NAND2_X1 port map( A1 => n35985, A2 => n18907, ZN => n16982);
   U18858 : CLKBUF_X12 port map( I => n13365, Z => n7789);
   U18859 : INV_X2 port map( I => n21666, ZN => n21834);
   U18861 : AOI21_X2 port map( A1 => n2542, A2 => n25858, B => n2541, ZN => 
                           n12221);
   U18863 : INV_X2 port map( I => n13213, ZN => n27251);
   U18864 : OAI21_X1 port map( A1 => n24608, A2 => n19255, B => n31161, ZN => 
                           n36021);
   U18872 : OAI21_X1 port map( A1 => n19255, A2 => n31161, B => n9257, ZN => 
                           n9256);
   U18875 : INV_X2 port map( I => n24232, ZN => n24176);
   U18878 : OR2_X1 port map( A1 => n37632, A2 => n12726, Z => n11981);
   U18880 : OR2_X1 port map( A1 => n15535, A2 => n12726, Z => n280);
   U18882 : OAI22_X1 port map( A1 => n34004, A2 => n39823, B1 => n31526, B2 => 
                           n17237, ZN => n26843);
   U18883 : OAI21_X1 port map( A1 => n29219, A2 => n31772, B => n29222, ZN => 
                           n12979);
   U18891 : XOR2_X1 port map( A1 => n266, A2 => n17737, Z => n38186);
   U18893 : OR2_X1 port map( A1 => n38186, A2 => n29495, Z => n20113);
   U18900 : OAI21_X1 port map( A1 => n31179, A2 => n23237, B => n23238, ZN => 
                           n4288);
   U18901 : INV_X2 port map( I => n5554, ZN => n8262);
   U18902 : NOR2_X1 port map( A1 => n15579, A2 => n23461, ZN => n31179);
   U18903 : INV_X2 port map( I => n15579, ZN => n23462);
   U18906 : INV_X2 port map( I => n3649, ZN => n25224);
   U18907 : NAND2_X1 port map( A1 => n21476, A2 => n21587, ZN => n21477);
   U18912 : NAND3_X1 port map( A1 => n29677, A2 => n29667, A3 => n31538, ZN => 
                           n29669);
   U18913 : NAND2_X1 port map( A1 => n13804, A2 => n15768, ZN => n13803);
   U18915 : INV_X1 port map( I => n11102, ZN => n34894);
   U18918 : NAND2_X1 port map( A1 => n34154, A2 => n7317, ZN => n25807);
   U18920 : NOR2_X1 port map( A1 => n22170, A2 => n21966, ZN => n39173);
   U18931 : INV_X2 port map( I => n22170, ZN => n20238);
   U18939 : INV_X2 port map( I => n38188, ZN => n26918);
   U18942 : AOI21_X1 port map( A1 => n5758, A2 => n5890, B => n5757, ZN => 
                           n38189);
   U18943 : AOI21_X1 port map( A1 => n5758, A2 => n5890, B => n5757, ZN => 
                           n38190);
   U18944 : AOI21_X1 port map( A1 => n5758, A2 => n5890, B => n5757, ZN => 
                           n5755);
   U18945 : NAND2_X1 port map( A1 => n28725, A2 => n17801, ZN => n5758);
   U18947 : XOR2_X1 port map( A1 => n38813, A2 => n30612, Z => n38191);
   U18955 : NAND2_X2 port map( A1 => n38847, A2 => n8406, ZN => n38192);
   U18956 : OAI21_X1 port map( A1 => n28179, A2 => n14389, B => n28181, ZN => 
                           n32418);
   U18961 : NAND2_X2 port map( A1 => n18605, A2 => n30585, ZN => n38193);
   U18963 : BUF_X2 port map( I => n36150, Z => n35684);
   U18969 : OR2_X2 port map( A1 => n8889, A2 => n37815, Z => n5111);
   U18975 : NOR2_X1 port map( A1 => n4434, A2 => n27314, ZN => n15917);
   U18980 : NOR2_X1 port map( A1 => n18711, A2 => n31202, ZN => n22138);
   U18989 : INV_X1 port map( I => n36509, ZN => n27455);
   U18991 : OAI21_X2 port map( A1 => n13445, A2 => n37904, B => n12307, ZN => 
                           n38194);
   U18994 : INV_X1 port map( I => n24106, ZN => n24168);
   U18995 : NAND2_X2 port map( A1 => n28305, A2 => n28304, ZN => n38195);
   U18997 : NOR2_X1 port map( A1 => n27097, A2 => n4771, ZN => n38568);
   U19000 : NAND2_X1 port map( A1 => n33950, A2 => n12478, ZN => n12368);
   U19005 : OAI21_X1 port map( A1 => n8608, A2 => n8607, B => n25114, ZN => 
                           n8606);
   U19008 : NAND3_X1 port map( A1 => n30805, A2 => n14448, A3 => n28546, ZN => 
                           n28470);
   U19009 : XOR2_X1 port map( A1 => n3187, A2 => n3188, Z => n38197);
   U19010 : NAND2_X2 port map( A1 => n36535, A2 => n38841, ZN => n38198);
   U19011 : NOR2_X2 port map( A1 => n16911, A2 => n34581, ZN => n38841);
   U19012 : NAND3_X1 port map( A1 => n32960, A2 => n32962, A3 => n7424, ZN => 
                           n30939);
   U19014 : OAI21_X1 port map( A1 => n35508, A2 => n25484, B => n611, ZN => 
                           n25537);
   U19015 : OR2_X2 port map( A1 => n3873, A2 => n30503, Z => n11726);
   U19018 : INV_X2 port map( I => n24805, ZN => n1026);
   U19019 : INV_X1 port map( I => n24805, ZN => n38347);
   U19020 : INV_X1 port map( I => n11105, ZN => n3100);
   U19021 : XOR2_X1 port map( A1 => n5177, A2 => n5176, Z => n38199);
   U19022 : NAND2_X2 port map( A1 => n29472, A2 => n29469, ZN => n38200);
   U19026 : OR2_X1 port map( A1 => n38199, A2 => n20960, Z => n15317);
   U19039 : INV_X1 port map( I => n31627, ZN => n7714);
   U19040 : NAND2_X1 port map( A1 => n11150, A2 => n138, ZN => n39328);
   U19041 : NAND2_X1 port map( A1 => n1108, A2 => n11150, ZN => n15173);
   U19043 : NAND3_X2 port map( A1 => n3399, A2 => n24907, A3 => n812, ZN => 
                           n38201);
   U19045 : NAND3_X1 port map( A1 => n3399, A2 => n24907, A3 => n812, ZN => 
                           n25151);
   U19046 : XOR2_X1 port map( A1 => n33722, A2 => n39115, Z => n38202);
   U19049 : NAND2_X2 port map( A1 => n31098, A2 => n3846, ZN => n38203);
   U19053 : OAI21_X1 port map( A1 => n35663, A2 => n5035, B => n3923, ZN => 
                           n38205);
   U19054 : NAND2_X1 port map( A1 => n9250, A2 => n9248, ZN => n38206);
   U19055 : INV_X2 port map( I => n17447, ZN => n28212);
   U19057 : INV_X2 port map( I => n34479, ZN => n33510);
   U19059 : INV_X1 port map( I => n2947, ZN => n39203);
   U19061 : NOR2_X1 port map( A1 => n495, A2 => n2947, ZN => n459);
   U19069 : CLKBUF_X4 port map( I => n17833, Z => n17792);
   U19071 : AOI21_X1 port map( A1 => n32974, A2 => n25874, B => n3575, ZN => 
                           n36375);
   U19072 : NAND2_X1 port map( A1 => n18866, A2 => n5258, ZN => n7427);
   U19073 : INV_X2 port map( I => n5258, ZN => n7426);
   U19077 : NAND2_X1 port map( A1 => n30299, A2 => n15423, ZN => n16213);
   U19080 : INV_X1 port map( I => n30299, ZN => n23379);
   U19086 : NAND3_X2 port map( A1 => n6195, A2 => n32545, A3 => n6192, ZN => 
                           n38207);
   U19098 : INV_X2 port map( I => n16048, ZN => n1039);
   U19101 : NAND2_X1 port map( A1 => n30574, A2 => n16048, ZN => n22987);
   U19102 : INV_X2 port map( I => n5211, ZN => n9193);
   U19104 : AOI21_X2 port map( A1 => n8238, A2 => n16575, B => n34472, ZN => 
                           n38208);
   U19107 : AOI21_X2 port map( A1 => n2542, A2 => n25858, B => n2541, ZN => 
                           n38209);
   U19108 : AOI21_X1 port map( A1 => n8238, A2 => n16575, B => n34472, ZN => 
                           n36842);
   U19111 : AOI21_X1 port map( A1 => n38141, A2 => n29802, B => n2792, ZN => 
                           n5880);
   U19113 : INV_X1 port map( I => n4353, ZN => n27318);
   U19114 : NAND2_X1 port map( A1 => n4353, A2 => n13973, ZN => n4345);
   U19117 : NAND3_X1 port map( A1 => n35963, A2 => n31931, A3 => n39316, ZN => 
                           n10841);
   U19120 : OAI22_X1 port map( A1 => n12212, A2 => n35545, B1 => n10122, B2 => 
                           n31931, ZN => n10078);
   U19121 : NAND2_X1 port map( A1 => n35545, A2 => n31931, ZN => n9350);
   U19126 : XNOR2_X1 port map( A1 => n3292, A2 => n25065, ZN => n38210);
   U19133 : INV_X2 port map( I => n8728, ZN => n1388);
   U19134 : NAND2_X1 port map( A1 => n8728, A2 => n29231, ZN => n38944);
   U19139 : AOI21_X1 port map( A1 => n35184, A2 => n7975, B => n1480, ZN => 
                           n2563);
   U19140 : CLKBUF_X12 port map( I => n20778, Z => n9809);
   U19141 : INV_X2 port map( I => n10764, ZN => n33815);
   U19146 : CLKBUF_X12 port map( I => n19930, Z => n438);
   U19149 : NOR2_X1 port map( A1 => n28546, A2 => n3944, ZN => n17073);
   U19150 : INV_X2 port map( I => n3944, ZN => n28643);
   U19153 : NAND2_X1 port map( A1 => n28546, A2 => n3944, ZN => n28647);
   U19154 : NOR2_X1 port map( A1 => n9530, A2 => n25943, ZN => n9529);
   U19157 : OAI21_X1 port map( A1 => n22173, A2 => n5450, B => n14833, ZN => 
                           n14903);
   U19161 : NAND3_X1 port map( A1 => n35901, A2 => n14064, A3 => n20128, ZN => 
                           n17765);
   U19165 : NOR2_X1 port map( A1 => n31433, A2 => n34279, ZN => n35608);
   U19168 : NAND2_X1 port map( A1 => n34279, A2 => n31433, ZN => n39159);
   U19175 : OAI21_X2 port map( A1 => n11735, A2 => n4463, B => n4462, ZN => 
                           n38212);
   U19177 : OAI21_X1 port map( A1 => n7922, A2 => n5941, B => n39417, ZN => 
                           n36805);
   U19178 : NAND2_X2 port map( A1 => n26648, A2 => n36953, ZN => n38213);
   U19182 : NAND2_X2 port map( A1 => n26641, A2 => n36911, ZN => n36953);
   U19183 : INV_X2 port map( I => n939, ZN => n920);
   U19186 : NAND2_X1 port map( A1 => n9682, A2 => n4516, ZN => n14985);
   U19187 : NAND2_X1 port map( A1 => n39454, A2 => n4516, ZN => n4511);
   U19192 : XOR2_X1 port map( A1 => n36468, A2 => n14302, Z => n38214);
   U19194 : INV_X1 port map( I => n25669, ZN => n38963);
   U19196 : CLKBUF_X12 port map( I => n25669, Z => n178);
   U19197 : XOR2_X1 port map( A1 => n2215, A2 => n2214, Z => n38215);
   U19198 : NAND3_X1 port map( A1 => n999, A2 => n495, A3 => n27153, ZN => 
                           n39707);
   U19200 : CLKBUF_X4 port map( I => n7654, Z => n21804);
   U19203 : INV_X1 port map( I => n7654, ZN => n21806);
   U19204 : INV_X1 port map( I => n28182, ZN => n4457);
   U19206 : AND2_X1 port map( A1 => n38199, A2 => n20960, Z => n26752);
   U19209 : NOR2_X1 port map( A1 => n27221, A2 => n5588, ZN => n27224);
   U19210 : INV_X1 port map( I => n11569, ZN => n25665);
   U19224 : OR3_X1 port map( A1 => n17180, A2 => n25782, A3 => n8407, Z => 
                           n25826);
   U19225 : NAND2_X1 port map( A1 => n7096, A2 => n19326, ZN => n27054);
   U19233 : INV_X1 port map( I => n19326, ZN => n27343);
   U19234 : OAI21_X1 port map( A1 => n27341, A2 => n27131, B => n19326, ZN => 
                           n4667);
   U19237 : INV_X1 port map( I => n6282, ZN => n1104);
   U19243 : NAND2_X1 port map( A1 => n32682, A2 => n36935, ZN => n32681);
   U19247 : NOR2_X1 port map( A1 => n11770, A2 => n2546, ZN => n38218);
   U19249 : NOR2_X1 port map( A1 => n11770, A2 => n2546, ZN => n38219);
   U19251 : NOR2_X1 port map( A1 => n11770, A2 => n2546, ZN => n2443);
   U19253 : INV_X2 port map( I => n23472, ZN => n23749);
   U19254 : AND2_X2 port map( A1 => n39820, A2 => n14332, Z => n25542);
   U19255 : CLKBUF_X12 port map( I => n5514, Z => n31283);
   U19261 : INV_X1 port map( I => n5514, ZN => n18816);
   U19262 : CLKBUF_X2 port map( I => n29678, Z => n33128);
   U19264 : NOR2_X1 port map( A1 => n36969, A2 => n33893, ZN => n2922);
   U19265 : XOR2_X1 port map( A1 => n1775, A2 => n16357, Z => n38221);
   U19268 : NOR2_X1 port map( A1 => n34008, A2 => n27985, ZN => n28105);
   U19269 : NOR2_X1 port map( A1 => n27484, A2 => n30758, ZN => n31000);
   U19277 : NAND3_X1 port map( A1 => n35115, A2 => n13753, A3 => n27484, ZN => 
                           n4741);
   U19278 : INV_X1 port map( I => n25289, ZN => n38511);
   U19279 : INV_X1 port map( I => n1234, ZN => n26908);
   U19280 : NAND3_X2 port map( A1 => n5344, A2 => n5342, A3 => n8048, ZN => 
                           n38222);
   U19281 : XOR2_X1 port map( A1 => n5731, A2 => n36339, Z => n38223);
   U19284 : INV_X1 port map( I => n7990, ZN => n7992);
   U19293 : XOR2_X1 port map( A1 => n16696, A2 => n16698, Z => n38224);
   U19299 : AOI21_X1 port map( A1 => n27287, A2 => n1080, B => n6010, ZN => 
                           n38225);
   U19300 : AOI21_X1 port map( A1 => n27287, A2 => n1080, B => n6010, ZN => 
                           n38226);
   U19305 : INV_X1 port map( I => n14869, ZN => n38227);
   U19306 : NAND3_X2 port map( A1 => n38516, A2 => n38525, A3 => n27242, ZN => 
                           n38228);
   U19307 : NAND3_X2 port map( A1 => n27238, A2 => n27237, A3 => n38690, ZN => 
                           n38516);
   U19309 : NAND2_X1 port map( A1 => n17685, A2 => n32675, ZN => n21503);
   U19311 : NOR3_X1 port map( A1 => n10242, A2 => n17685, A3 => n12077, ZN => 
                           n12040);
   U19312 : CLKBUF_X12 port map( I => n29199, Z => n30193);
   U19319 : INV_X1 port map( I => n29199, ZN => n30229);
   U19320 : INV_X1 port map( I => n32043, ZN => n12303);
   U19322 : AOI21_X1 port map( A1 => n4008, A2 => n39098, B => n5896, ZN => 
                           n18326);
   U19323 : NOR2_X1 port map( A1 => n35138, A2 => n692, ZN => n2311);
   U19327 : AND2_X2 port map( A1 => n22925, A2 => n18209, Z => n22999);
   U19336 : INV_X1 port map( I => n35242, ZN => n20041);
   U19339 : NOR2_X1 port map( A1 => n1420, A2 => n38155, ZN => n15963);
   U19340 : XOR2_X1 port map( A1 => n38564, A2 => n3232, Z => n38229);
   U19341 : INV_X1 port map( I => n8093, ZN => n38230);
   U19342 : NOR2_X1 port map( A1 => n28704, A2 => n38220, ZN => n27897);
   U19344 : INV_X1 port map( I => n26558, ZN => n35746);
   U19350 : NOR2_X1 port map( A1 => n35254, A2 => n12198, ZN => n30176);
   U19351 : INV_X1 port map( I => n28686, ZN => n31045);
   U19366 : OAI21_X1 port map( A1 => n1527, A2 => n38168, B => n14375, ZN => 
                           n3433);
   U19368 : INV_X2 port map( I => n5383, ZN => n28608);
   U19372 : NAND2_X1 port map( A1 => n5383, A2 => n36588, ZN => n3637);
   U19374 : NAND2_X1 port map( A1 => n7769, A2 => n10980, ZN => n39076);
   U19375 : NOR2_X1 port map( A1 => n16213, A2 => n23358, ZN => n462);
   U19378 : NAND2_X1 port map( A1 => n23379, A2 => n23358, ZN => n23359);
   U19379 : NAND2_X1 port map( A1 => n23358, A2 => n23250, ZN => n31199);
   U19381 : NAND2_X2 port map( A1 => n12660, A2 => n12661, ZN => n10558);
   U19384 : NAND3_X2 port map( A1 => n22048, A2 => n37199, A3 => n19089, ZN => 
                           n12660);
   U19386 : INV_X2 port map( I => n38235, ZN => n11363);
   U19387 : NOR2_X2 port map( A1 => n25539, A2 => n39820, ZN => n38235);
   U19388 : INV_X1 port map( I => n14282, ZN => n38237);
   U19389 : INV_X2 port map( I => n38239, ZN => n39810);
   U19390 : XOR2_X1 port map( A1 => n7199, A2 => n7201, Z => n38239);
   U19391 : XOR2_X1 port map( A1 => n25172, A2 => n18428, Z => n11369);
   U19393 : XOR2_X1 port map( A1 => n26261, A2 => n31537, Z => n9762);
   U19398 : XOR2_X1 port map( A1 => n14353, A2 => n23710, Z => n23887);
   U19403 : XOR2_X1 port map( A1 => n35070, A2 => n38179, Z => n17119);
   U19405 : NOR2_X1 port map( A1 => n16948, A2 => n16949, ZN => n17936);
   U19406 : XOR2_X1 port map( A1 => n23666, A2 => n38240, Z => n36272);
   U19413 : XOR2_X1 port map( A1 => n23729, A2 => n12799, Z => n38240);
   U19414 : AOI21_X1 port map( A1 => n6581, A2 => n37589, B => n14561, ZN => 
                           n13206);
   U19415 : OAI21_X2 port map( A1 => n11598, A2 => n21439, B => n6690, ZN => 
                           n33738);
   U19416 : AOI22_X2 port map( A1 => n693, A2 => n21692, B1 => n21339, B2 => 
                           n21687, ZN => n21439);
   U19419 : NAND2_X2 port map( A1 => n21993, A2 => n21992, ZN => n17310);
   U19422 : BUF_X2 port map( I => n39639, Z => n38241);
   U19425 : OR2_X2 port map( A1 => n18998, A2 => n8071, Z => n22272);
   U19427 : AOI22_X1 port map( A1 => n29599, A2 => n31667, B1 => n4786, B2 => 
                           n38420, ZN => n33746);
   U19430 : XOR2_X1 port map( A1 => n1618, A2 => n23686, Z => n24033);
   U19432 : NAND2_X2 port map( A1 => n34662, A2 => n37395, ZN => n38242);
   U19434 : NOR2_X2 port map( A1 => n38390, A2 => n7491, ZN => n16013);
   U19440 : XOR2_X1 port map( A1 => n36057, A2 => n38243, Z => n14110);
   U19442 : XOR2_X1 port map( A1 => n22454, A2 => n22766, Z => n38243);
   U19448 : NAND2_X2 port map( A1 => n38508, A2 => n35697, ZN => n3015);
   U19451 : AND2_X1 port map( A1 => n8604, A2 => n8395, Z => n18628);
   U19454 : XOR2_X1 port map( A1 => n5322, A2 => n6516, Z => n24195);
   U19455 : BUF_X2 port map( I => n18425, Z => n38248);
   U19459 : NAND2_X2 port map( A1 => n22843, A2 => n2163, ZN => n38249);
   U19469 : OAI21_X2 port map( A1 => n13121, A2 => n19218, B => n18162, ZN => 
                           n32897);
   U19473 : XOR2_X1 port map( A1 => n792, A2 => n3824, Z => n3823);
   U19476 : XNOR2_X1 port map( A1 => n3503, A2 => n18175, ZN => n3824);
   U19477 : XOR2_X1 port map( A1 => n14113, A2 => n38253, Z => n7674);
   U19478 : XOR2_X1 port map( A1 => n22603, A2 => n14112, Z => n38253);
   U19482 : XOR2_X1 port map( A1 => n27530, A2 => n38254, Z => n27875);
   U19483 : XOR2_X1 port map( A1 => n27527, A2 => n39465, Z => n38254);
   U19484 : XOR2_X1 port map( A1 => n18175, A2 => n32122, Z => n23863);
   U19487 : AND2_X1 port map( A1 => n740, A2 => n8556, Z => n8652);
   U19494 : NAND2_X2 port map( A1 => n36623, A2 => n5028, ZN => n28730);
   U19499 : NAND2_X2 port map( A1 => n31042, A2 => n38923, ZN => n36623);
   U19508 : XOR2_X1 port map( A1 => n4440, A2 => n16199, Z => n4438);
   U19511 : XOR2_X1 port map( A1 => n15346, A2 => n16226, Z => n16199);
   U19514 : NAND2_X2 port map( A1 => n39262, A2 => n27064, ZN => n8372);
   U19517 : AND2_X1 port map( A1 => n9118, A2 => n735, Z => n6501);
   U19519 : XOR2_X1 port map( A1 => n13369, A2 => n13367, Z => n18156);
   U19522 : XOR2_X1 port map( A1 => n8408, A2 => n8410, Z => n32806);
   U19524 : OR2_X1 port map( A1 => n38255, A2 => n30198, Z => n2767);
   U19525 : NOR2_X2 port map( A1 => n33861, A2 => n1755, ZN => n30198);
   U19528 : INV_X1 port map( I => n29222, ZN => n29224);
   U19530 : NAND2_X1 port map( A1 => n29222, A2 => n6002, ZN => n3415);
   U19532 : NOR2_X2 port map( A1 => n38257, A2 => n38256, ZN => n29222);
   U19534 : INV_X1 port map( I => n36694, ZN => n38256);
   U19541 : OAI21_X1 port map( A1 => n18278, A2 => n18039, B => n38258, ZN => 
                           n36862);
   U19543 : NAND2_X1 port map( A1 => n29205, A2 => n18039, ZN => n38258);
   U19544 : NAND2_X2 port map( A1 => n10595, A2 => n34897, ZN => n19326);
   U19548 : XOR2_X1 port map( A1 => n26429, A2 => n12300, Z => n12299);
   U19549 : XOR2_X1 port map( A1 => n33027, A2 => n38619, Z => n26429);
   U19550 : OAI21_X2 port map( A1 => n11886, A2 => n29201, B => n34983, ZN => 
                           n29204);
   U19551 : NAND2_X2 port map( A1 => n7745, A2 => n3945, ZN => n3944);
   U19553 : XOR2_X1 port map( A1 => n34491, A2 => n11814, Z => n16500);
   U19557 : NOR2_X2 port map( A1 => n7872, A2 => n28215, ZN => n38443);
   U19567 : INV_X2 port map( I => n38259, ZN => n20860);
   U19569 : OAI21_X1 port map( A1 => n16577, A2 => n17708, B => n38260, ZN => 
                           n5778);
   U19575 : AOI22_X1 port map( A1 => n5779, A2 => n20498, B1 => n29717, B2 => 
                           n29722, ZN => n38260);
   U19576 : XOR2_X1 port map( A1 => n22668, A2 => n38261, Z => n649);
   U19586 : NAND2_X2 port map( A1 => n17901, A2 => n17902, ZN => n35241);
   U19594 : NOR2_X2 port map( A1 => n14626, A2 => n16953, ZN => n17901);
   U19596 : OAI21_X2 port map( A1 => n8105, A2 => n26726, B => n26725, ZN => 
                           n27269);
   U19599 : XOR2_X1 port map( A1 => n2005, A2 => n2002, Z => n9649);
   U19601 : BUF_X2 port map( I => n20018, Z => n38262);
   U19603 : XOR2_X1 port map( A1 => n24017, A2 => n24016, Z => n14719);
   U19605 : XOR2_X1 port map( A1 => n24026, A2 => n38263, Z => n39591);
   U19607 : XOR2_X1 port map( A1 => n10722, A2 => n11180, Z => n38263);
   U19608 : AOI21_X2 port map( A1 => n36287, A2 => n34570, B => n27103, ZN => 
                           n27802);
   U19610 : NOR2_X1 port map( A1 => n9489, A2 => n9487, ZN => n5458);
   U19612 : XOR2_X1 port map( A1 => n38264, A2 => n18316, Z => n18315);
   U19616 : XOR2_X1 port map( A1 => n18319, A2 => n30925, Z => n38264);
   U19617 : XOR2_X1 port map( A1 => n1262, A2 => n25086, Z => n8240);
   U19629 : OAI22_X2 port map( A1 => n14538, A2 => n15826, B1 => n20119, B2 => 
                           n1608, ZN => n32637);
   U19634 : XOR2_X1 port map( A1 => n27640, A2 => n38265, Z => n39742);
   U19638 : INV_X1 port map( I => n29920, ZN => n38265);
   U19639 : NAND2_X2 port map( A1 => n14586, A2 => n38873, ZN => n27640);
   U19647 : NAND2_X1 port map( A1 => n19420, A2 => n8966, ZN => n24500);
   U19652 : NOR2_X2 port map( A1 => n38835, A2 => n32690, ZN => n30696);
   U19653 : NAND2_X2 port map( A1 => n9173, A2 => n35673, ZN => n35187);
   U19654 : XOR2_X1 port map( A1 => n23736, A2 => n23913, Z => n12921);
   U19659 : XOR2_X1 port map( A1 => n38267, A2 => n27465, Z => Ciphertext(185))
                           ;
   U19665 : NAND2_X1 port map( A1 => n27456, A2 => n37158, ZN => n26641);
   U19668 : XOR2_X1 port map( A1 => n26257, A2 => n13131, Z => n17063);
   U19676 : XOR2_X1 port map( A1 => n26381, A2 => n9870, Z => n13131);
   U19678 : NAND2_X2 port map( A1 => n2316, A2 => n25755, ZN => n35138);
   U19679 : BUF_X2 port map( I => n32095, Z => n38269);
   U19681 : NAND2_X2 port map( A1 => n28256, A2 => n3989, ZN => n28047);
   U19683 : XNOR2_X1 port map( A1 => n10520, A2 => n6185, ZN => n25222);
   U19684 : NAND2_X2 port map( A1 => n38296, A2 => n38270, ZN => n25813);
   U19687 : AOI22_X2 port map( A1 => n12404, A2 => n1117, B1 => n19863, B2 => 
                           n25660, ZN => n38270);
   U19688 : OAI21_X2 port map( A1 => n37123, A2 => n9064, B => n9063, ZN => 
                           n29794);
   U19689 : XOR2_X1 port map( A1 => n38271, A2 => n38969, Z => n27919);
   U19692 : XOR2_X1 port map( A1 => n33883, A2 => n27788, Z => n38271);
   U19698 : NAND2_X2 port map( A1 => n959, A2 => n626, ZN => n33586);
   U19699 : NAND2_X2 port map( A1 => n6054, A2 => n6053, ZN => n23775);
   U19700 : AOI22_X2 port map( A1 => n38274, A2 => n38272, B1 => n21527, B2 => 
                           n39627, ZN => n39616);
   U19701 : NOR2_X2 port map( A1 => n39627, A2 => n38273, ZN => n38272);
   U19704 : INV_X2 port map( I => n35071, ZN => n38274);
   U19706 : XOR2_X1 port map( A1 => n29071, A2 => n28886, Z => n28914);
   U19710 : NAND3_X2 port map( A1 => n35415, A2 => n35414, A3 => n16632, ZN => 
                           n11831);
   U19712 : XOR2_X1 port map( A1 => n8183, A2 => n25252, Z => n21253);
   U19715 : NAND2_X2 port map( A1 => n12676, A2 => n35688, ZN => n8183);
   U19717 : NAND2_X2 port map( A1 => n4990, A2 => n30595, ZN => n32748);
   U19718 : XOR2_X1 port map( A1 => n35218, A2 => n8302, Z => n36637);
   U19719 : NOR2_X2 port map( A1 => n1333, A2 => n3003, ZN => n22230);
   U19722 : INV_X2 port map( I => n31271, ZN => n38839);
   U19724 : XOR2_X1 port map( A1 => n5179, A2 => n36540, Z => n31271);
   U19725 : NAND2_X2 port map( A1 => n10128, A2 => n10126, ZN => n38395);
   U19728 : XOR2_X1 port map( A1 => n28971, A2 => n13639, Z => n29123);
   U19729 : NAND2_X2 port map( A1 => n28648, A2 => n18891, ZN => n13639);
   U19730 : NAND2_X2 port map( A1 => n34579, A2 => n38276, ZN => n27023);
   U19742 : XOR2_X1 port map( A1 => n6317, A2 => n6196, Z => n20727);
   U19743 : NAND2_X2 port map( A1 => n28416, A2 => n28417, ZN => n6196);
   U19744 : NOR2_X2 port map( A1 => n34685, A2 => n34350, ZN => n25737);
   U19745 : XOR2_X1 port map( A1 => n27807, A2 => n20846, Z => n32647);
   U19746 : XOR2_X1 port map( A1 => n33197, A2 => n25252, Z => n25302);
   U19753 : NAND2_X1 port map( A1 => n4516, A2 => n6904, ZN => n12569);
   U19757 : NAND2_X2 port map( A1 => n9540, A2 => n25559, ZN => n4516);
   U19759 : NAND2_X2 port map( A1 => n5675, A2 => n27274, ZN => n27085);
   U19760 : NAND3_X2 port map( A1 => n38277, A2 => n27151, A3 => n27148, ZN => 
                           n27778);
   U19761 : AOI22_X2 port map( A1 => n33910, A2 => n38278, B1 => n28401, B2 => 
                           n11490, ZN => n11492);
   U19765 : NAND2_X2 port map( A1 => n2937, A2 => n12537, ZN => n38278);
   U19767 : AOI21_X2 port map( A1 => n11591, A2 => n943, B => n11590, ZN => 
                           n13245);
   U19768 : INV_X2 port map( I => n38280, ZN => n37054);
   U19779 : XOR2_X1 port map( A1 => n3459, A2 => n3456, Z => n38280);
   U19782 : NOR3_X1 port map( A1 => n1429, A2 => n10907, A3 => n18871, ZN => 
                           n32075);
   U19783 : XOR2_X1 port map( A1 => n29050, A2 => n29125, Z => n29158);
   U19786 : XOR2_X1 port map( A1 => n38605, A2 => n21271, Z => n36396);
   U19791 : XOR2_X1 port map( A1 => n30502, A2 => n38890, Z => n38781);
   U19795 : OAI22_X2 port map( A1 => n924, A2 => n3388, B1 => n38214, B2 => 
                           n14458, ZN => n8686);
   U19806 : OAI21_X2 port map( A1 => n35295, A2 => n35296, B => n32714, ZN => 
                           n29438);
   U19808 : XOR2_X1 port map( A1 => n22657, A2 => n22761, Z => n22608);
   U19816 : NAND2_X2 port map( A1 => n16548, A2 => n30212, ZN => n38829);
   U19819 : NAND3_X2 port map( A1 => n17648, A2 => n32598, A3 => n2632, ZN => 
                           n39481);
   U19823 : NAND2_X2 port map( A1 => n2633, A2 => n1633, ZN => n17648);
   U19825 : NAND2_X2 port map( A1 => n39503, A2 => n38281, ZN => n27683);
   U19826 : AOI22_X1 port map( A1 => n27017, A2 => n39424, B1 => n27224, B2 => 
                           n13278, ZN => n38281);
   U19827 : NOR2_X2 port map( A1 => n38283, A2 => n38282, ZN => n22803);
   U19828 : INV_X1 port map( I => n14752, ZN => n38284);
   U19829 : BUF_X2 port map( I => n24712, Z => n38285);
   U19830 : AND2_X1 port map( A1 => n20541, A2 => n33963, Z => n38919);
   U19831 : NAND2_X2 port map( A1 => n38286, A2 => n38354, ZN => n16526);
   U19835 : XOR2_X1 port map( A1 => n16552, A2 => n16554, Z => n32750);
   U19841 : AOI21_X2 port map( A1 => n37141, A2 => n32084, B => n34643, ZN => 
                           n16636);
   U19848 : NAND2_X2 port map( A1 => n30311, A2 => n94, ZN => n33944);
   U19857 : XOR2_X1 port map( A1 => n6571, A2 => n11105, Z => n26490);
   U19858 : NAND2_X2 port map( A1 => n32380, A2 => n39777, ZN => n11105);
   U19861 : XOR2_X1 port map( A1 => n26567, A2 => n26334, Z => n35721);
   U19868 : NAND2_X2 port map( A1 => n9377, A2 => n31883, ZN => n26567);
   U19871 : NOR2_X2 port map( A1 => n33289, A2 => n35954, ZN => n24219);
   U19872 : NOR2_X2 port map( A1 => n22019, A2 => n2818, ZN => n38287);
   U19877 : NAND2_X2 port map( A1 => n38391, A2 => n38288, ZN => n11120);
   U19880 : XOR2_X1 port map( A1 => n38289, A2 => n1160, Z => Ciphertext(22));
   U19887 : NOR2_X1 port map( A1 => n38348, A2 => n30577, ZN => n38289);
   U19889 : NAND2_X2 port map( A1 => n35158, A2 => n17420, ZN => n27779);
   U19891 : OAI21_X2 port map( A1 => n25838, A2 => n38982, B => n25837, ZN => 
                           n9989);
   U19900 : XOR2_X1 port map( A1 => n33010, A2 => n38291, Z => n23921);
   U19904 : INV_X2 port map( I => n24049, ZN => n38291);
   U19906 : BUF_X2 port map( I => n388, Z => n38292);
   U19907 : XOR2_X1 port map( A1 => n38294, A2 => n20400, Z => n18188);
   U19909 : XOR2_X1 port map( A1 => n36628, A2 => n27648, Z => n38294);
   U19910 : NAND2_X2 port map( A1 => n35750, A2 => n34644, ZN => n10032);
   U19911 : AOI22_X2 port map( A1 => n18484, A2 => n2396, B1 => n24331, B2 => 
                           n24330, ZN => n34263);
   U19915 : NOR2_X2 port map( A1 => n12733, A2 => n24328, ZN => n18484);
   U19916 : XOR2_X1 port map( A1 => n38958, A2 => n38192, Z => n38809);
   U19917 : NAND2_X2 port map( A1 => n38847, A2 => n8406, ZN => n7990);
   U19918 : XOR2_X1 port map( A1 => n38295, A2 => n2351, Z => n23202);
   U19921 : XOR2_X1 port map( A1 => n14297, A2 => n2354, Z => n38295);
   U19924 : OAI21_X2 port map( A1 => n34099, A2 => n229, B => n25662, ZN => 
                           n38296);
   U19925 : XOR2_X1 port map( A1 => n29039, A2 => n28920, Z => n8678);
   U19926 : XOR2_X1 port map( A1 => n9106, A2 => n12989, Z => n28920);
   U19927 : XOR2_X1 port map( A1 => n24019, A2 => n23676, Z => n5255);
   U19930 : NAND2_X2 port map( A1 => n38298, A2 => n38297, ZN => n20255);
   U19931 : AOI22_X1 port map( A1 => n32372, A2 => n12144, B1 => n17233, B2 => 
                           n14418, ZN => n38297);
   U19933 : OAI21_X2 port map( A1 => n21535, A2 => n21536, B => n14501, ZN => 
                           n38298);
   U19941 : XNOR2_X1 port map( A1 => n26391, A2 => n19450, ZN => n26449);
   U19943 : NAND3_X2 port map( A1 => n38301, A2 => n37182, A3 => n9427, ZN => 
                           n18994);
   U19944 : NAND2_X2 port map( A1 => n28429, A2 => n12797, ZN => n8729);
   U19946 : OAI21_X1 port map( A1 => n37126, A2 => n4347, B => n38308, ZN => 
                           n8328);
   U19948 : XOR2_X1 port map( A1 => n16109, A2 => n16110, Z => n15865);
   U19949 : NAND2_X1 port map( A1 => n22206, A2 => n19837, ZN => n38932);
   U19953 : NAND2_X1 port map( A1 => n38932, A2 => n38931, ZN => n22211);
   U19959 : NOR2_X2 port map( A1 => n12063, A2 => n6150, ZN => n26334);
   U19964 : XOR2_X1 port map( A1 => n23868, A2 => n675, Z => n20485);
   U19968 : XOR2_X1 port map( A1 => n36842, A2 => n19656, Z => n23868);
   U19972 : NAND2_X2 port map( A1 => n18170, A2 => n18171, ZN => n20589);
   U19973 : XOR2_X1 port map( A1 => n12215, A2 => n38309, Z => n21116);
   U19977 : XOR2_X1 port map( A1 => n31582, A2 => n28986, Z => n38309);
   U19978 : OAI22_X2 port map( A1 => n13427, A2 => n33849, B1 => n26811, B2 => 
                           n26810, ZN => n12756);
   U19985 : INV_X2 port map( I => n38310, ZN => n13427);
   U19996 : NOR2_X2 port map( A1 => n12755, A2 => n13770, ZN => n38310);
   U19997 : NAND2_X2 port map( A1 => n17583, A2 => n5424, ZN => n8423);
   U20002 : AND2_X1 port map( A1 => n10940, A2 => n24408, Z => n39271);
   U20003 : INV_X2 port map( I => n10520, ZN => n25256);
   U20004 : NAND2_X2 port map( A1 => n35664, A2 => n19559, ZN => n23302);
   U20009 : INV_X1 port map( I => n2283, ZN => n27520);
   U20023 : OR2_X1 port map( A1 => n36371, A2 => n3644, Z => n17998);
   U20028 : XOR2_X1 port map( A1 => n18423, A2 => n18421, Z => n34956);
   U20029 : NAND3_X2 port map( A1 => n38312, A2 => n39324, A3 => n39325, ZN => 
                           n35813);
   U20031 : XOR2_X1 port map( A1 => n12520, A2 => n36389, Z => n38486);
   U20033 : XNOR2_X1 port map( A1 => n10683, A2 => n10684, ZN => n38465);
   U20034 : NOR3_X2 port map( A1 => n37108, A2 => n39303, A3 => n39752, ZN => 
                           n35950);
   U20035 : XOR2_X1 port map( A1 => n39804, A2 => n17310, Z => n18239);
   U20040 : XOR2_X1 port map( A1 => n26229, A2 => n38313, Z => n38842);
   U20041 : XOR2_X1 port map( A1 => n11298, A2 => n26525, Z => n38313);
   U20042 : XOR2_X1 port map( A1 => n38314, A2 => n20748, Z => Ciphertext(165))
                           ;
   U20046 : NOR4_X2 port map( A1 => n34706, A2 => n34707, A3 => n35625, A4 => 
                           n35624, ZN => n38314);
   U20049 : NAND2_X2 port map( A1 => n36099, A2 => n26113, ZN => n39066);
   U20050 : NAND3_X2 port map( A1 => n36678, A2 => n31004, A3 => n371, ZN => 
                           n35665);
   U20054 : NAND2_X1 port map( A1 => n1948, A2 => n15427, ZN => n16146);
   U20055 : XOR2_X1 port map( A1 => n38316, A2 => n38315, Z => n31485);
   U20057 : XOR2_X1 port map( A1 => n17189, A2 => n31576, Z => n38315);
   U20061 : XOR2_X1 port map( A1 => n1323, A2 => n31504, Z => n38316);
   U20062 : AND2_X1 port map( A1 => n5768, A2 => n38317, Z => n12680);
   U20063 : XOR2_X1 port map( A1 => n3976, A2 => n3975, Z => n38742);
   U20064 : INV_X1 port map( I => n19783, ZN => n38319);
   U20066 : INV_X1 port map( I => n14789, ZN => n38320);
   U20068 : NAND3_X1 port map( A1 => n11453, A2 => n38656, A3 => n19068, ZN => 
                           n12746);
   U20069 : XOR2_X1 port map( A1 => n38321, A2 => n23985, Z => n23991);
   U20070 : XOR2_X1 port map( A1 => n23984, A2 => n35235, Z => n38321);
   U20073 : NAND2_X1 port map( A1 => n3593, A2 => n38960, ZN => n39016);
   U20075 : XOR2_X1 port map( A1 => n38322, A2 => n11570, Z => n32994);
   U20077 : XOR2_X1 port map( A1 => n33924, A2 => n25197, Z => n38322);
   U20078 : OAI22_X1 port map( A1 => n21983, A2 => n3907, B1 => n3644, B2 => 
                           n38323, ZN => n11440);
   U20080 : OR2_X1 port map( A1 => n3907, A2 => n21982, Z => n38323);
   U20081 : XOR2_X1 port map( A1 => n38324, A2 => n19648, Z => Ciphertext(99));
   U20085 : NAND2_X1 port map( A1 => n29736, A2 => n19369, ZN => n38324);
   U20086 : XOR2_X1 port map( A1 => n24074, A2 => n20973, Z => n20550);
   U20089 : XOR2_X1 port map( A1 => n23898, A2 => n23955, Z => n24074);
   U20092 : NAND2_X2 port map( A1 => n33161, A2 => n13755, ZN => n38669);
   U20093 : XOR2_X1 port map( A1 => n25234, A2 => n14214, Z => n12997);
   U20096 : XOR2_X1 port map( A1 => n38325, A2 => n19534, Z => Ciphertext(113))
                           ;
   U20098 : NAND2_X1 port map( A1 => n6441, A2 => n6438, ZN => n38325);
   U20099 : XOR2_X1 port map( A1 => n18335, A2 => n38326, Z => n850);
   U20105 : XOR2_X1 port map( A1 => n35202, A2 => n33735, Z => n38326);
   U20107 : XOR2_X1 port map( A1 => n29041, A2 => n31547, Z => n28873);
   U20116 : OAI21_X2 port map( A1 => n2335, A2 => n2334, B => n33649, ZN => 
                           n31547);
   U20117 : NAND2_X2 port map( A1 => n31027, A2 => n30668, ZN => n5424);
   U20120 : XOR2_X1 port map( A1 => n18813, A2 => n7070, Z => n39516);
   U20126 : BUF_X2 port map( I => n16123, Z => n38328);
   U20132 : AND2_X1 port map( A1 => n5514, A2 => n39011, Z => n39110);
   U20134 : NAND3_X1 port map( A1 => n24532, A2 => n6169, A3 => n957, ZN => 
                           n38331);
   U20135 : NAND2_X2 port map( A1 => n7487, A2 => n38332, ZN => n24002);
   U20136 : AOI22_X2 port map( A1 => n30460, A2 => n1644, B1 => n33080, B2 => 
                           n605, ZN => n38332);
   U20140 : NAND2_X2 port map( A1 => n27116, A2 => n7588, ZN => n38333);
   U20150 : OR2_X1 port map( A1 => n18619, A2 => n19949, Z => n17586);
   U20151 : XOR2_X1 port map( A1 => n26539, A2 => n26513, Z => n5225);
   U20155 : XOR2_X1 port map( A1 => n38619, A2 => n26161, Z => n26513);
   U20159 : XNOR2_X1 port map( A1 => n22551, A2 => n5463, ZN => n39040);
   U20164 : XOR2_X1 port map( A1 => n22586, A2 => n20392, Z => n5463);
   U20166 : NOR2_X2 port map( A1 => n14746, A2 => n20788, ZN => n38334);
   U20167 : XOR2_X1 port map( A1 => n25079, A2 => n38336, Z => n39563);
   U20168 : NAND2_X2 port map( A1 => n6574, A2 => n6837, ZN => n25079);
   U20169 : NOR2_X1 port map( A1 => n20739, A2 => n32043, ZN => n28324);
   U20179 : INV_X1 port map( I => n39140, ZN => n34524);
   U20188 : OAI21_X2 port map( A1 => n36433, A2 => n36434, B => n38642, ZN => 
                           n39140);
   U20198 : AND3_X1 port map( A1 => n3988, A2 => n28616, A3 => n6287, Z => 
                           n5385);
   U20201 : AOI22_X2 port map( A1 => n37181, A2 => n38338, B1 => n25627, B2 => 
                           n37748, ZN => n31082);
   U20204 : NOR2_X2 port map( A1 => n11476, A2 => n2272, ZN => n38400);
   U20207 : AOI22_X2 port map( A1 => n16206, A2 => n35326, B1 => n4871, B2 => 
                           n28548, ZN => n35262);
   U20212 : NAND2_X2 port map( A1 => n32651, A2 => n32637, ZN => n16579);
   U20215 : NOR2_X1 port map( A1 => n10913, A2 => n26978, ZN => n34868);
   U20223 : NOR2_X2 port map( A1 => n852, A2 => n17097, ZN => n10913);
   U20228 : XOR2_X1 port map( A1 => n39215, A2 => n10525, Z => n34616);
   U20230 : NAND2_X2 port map( A1 => n21245, A2 => n10472, ZN => n19559);
   U20240 : INV_X2 port map( I => n19671, ZN => n1299);
   U20243 : NAND2_X2 port map( A1 => n13087, A2 => n39819, ZN => n19671);
   U20244 : NAND2_X2 port map( A1 => n4010, A2 => n10729, ZN => n4301);
   U20245 : OAI22_X2 port map( A1 => n7107, A2 => n33359, B1 => n7108, B2 => 
                           n38339, ZN => n22659);
   U20247 : NAND2_X2 port map( A1 => n38663, A2 => n39782, ZN => n7512);
   U20248 : XOR2_X1 port map( A1 => n10647, A2 => n4734, Z => n11062);
   U20249 : NAND2_X2 port map( A1 => n10646, A2 => n10645, ZN => n10647);
   U20253 : NOR2_X2 port map( A1 => n23072, A2 => n22919, ZN => n36230);
   U20255 : NAND2_X2 port map( A1 => n38634, A2 => n2850, ZN => n17653);
   U20262 : NAND2_X2 port map( A1 => n38340, A2 => n16763, ZN => n21543);
   U20264 : XOR2_X1 port map( A1 => n16627, A2 => n1558, Z => n11570);
   U20265 : INV_X2 port map( I => n38341, ZN => n21117);
   U20267 : NOR2_X2 port map( A1 => n2654, A2 => n21982, ZN => n38341);
   U20268 : NAND2_X2 port map( A1 => n38342, A2 => n2941, ZN => n18012);
   U20278 : XOR2_X1 port map( A1 => n29029, A2 => n29030, Z => n9768);
   U20279 : XOR2_X1 port map( A1 => n15780, A2 => n29818, Z => n29030);
   U20296 : XOR2_X1 port map( A1 => n38343, A2 => n23876, Z => n1923);
   U20298 : XOR2_X1 port map( A1 => n13224, A2 => n36143, Z => n38343);
   U20300 : XOR2_X1 port map( A1 => n12014, A2 => n3150, Z => n38344);
   U20303 : AND2_X2 port map( A1 => n34134, A2 => n11657, Z => n25364);
   U20304 : XOR2_X1 port map( A1 => n17567, A2 => n35320, Z => n21108);
   U20305 : NAND2_X2 port map( A1 => n38469, A2 => n8320, ZN => n17567);
   U20306 : XOR2_X1 port map( A1 => n15517, A2 => n15516, Z => n19928);
   U20308 : NAND2_X2 port map( A1 => n8314, A2 => n1579, ZN => n8317);
   U20311 : OAI21_X2 port map( A1 => n28727, A2 => n8094, B => n34525, ZN => 
                           n8090);
   U20316 : INV_X2 port map( I => n39227, ZN => n28727);
   U20318 : NAND3_X2 port map( A1 => n27868, A2 => n27867, A3 => n18149, ZN => 
                           n39227);
   U20319 : OAI21_X2 port map( A1 => n1074, A2 => n12406, B => n1200, ZN => 
                           n38345);
   U20320 : NAND3_X2 port map( A1 => n31695, A2 => n24957, A3 => n38346, ZN => 
                           n26092);
   U20321 : NAND3_X1 port map( A1 => n38338, A2 => n25756, A3 => n12675, ZN => 
                           n38346);
   U20324 : INV_X2 port map( I => n26432, ZN => n12934);
   U20325 : NOR2_X1 port map( A1 => n20889, A2 => n35399, ZN => n14777);
   U20326 : NAND2_X2 port map( A1 => n21774, A2 => n21773, ZN => n20889);
   U20328 : NAND2_X1 port map( A1 => n25261, A2 => n11727, ZN => n34411);
   U20331 : NAND2_X1 port map( A1 => n11394, A2 => n11395, ZN => n38348);
   U20335 : NAND2_X1 port map( A1 => n38686, A2 => n33495, ZN => n12704);
   U20339 : XOR2_X1 port map( A1 => n23970, A2 => n23967, Z => n23869);
   U20340 : NAND2_X2 port map( A1 => n23301, A2 => n31052, ZN => n23967);
   U20349 : OR2_X1 port map( A1 => n33980, A2 => n28250, Z => n28247);
   U20351 : XOR2_X1 port map( A1 => n15995, A2 => n15994, Z => n33980);
   U20353 : XOR2_X1 port map( A1 => n23764, A2 => n38350, Z => n37044);
   U20359 : INV_X2 port map( I => n23654, ZN => n38350);
   U20360 : XOR2_X1 port map( A1 => n38351, A2 => n6531, Z => n6528);
   U20361 : XOR2_X1 port map( A1 => n1620, A2 => n5699, Z => n38351);
   U20362 : XOR2_X1 port map( A1 => n29819, A2 => n29506, Z => n38352);
   U20364 : OAI21_X2 port map( A1 => n39034, A2 => n22863, B => n9472, ZN => 
                           n6213);
   U20366 : AND2_X2 port map( A1 => n3839, A2 => n7696, Z => n21461);
   U20368 : NAND2_X2 port map( A1 => n16123, A2 => n14940, ZN => n7207);
   U20369 : NOR2_X2 port map( A1 => n961, A2 => n23401, ZN => n38353);
   U20371 : OAI21_X2 port map( A1 => n6744, A2 => n2898, B => n37212, ZN => 
                           n38354);
   U20372 : OAI21_X2 port map( A1 => n3981, A2 => n9688, B => n37006, ZN => 
                           n2147);
   U20374 : XOR2_X1 port map( A1 => n3652, A2 => n3650, Z => n33446);
   U20381 : XOR2_X1 port map( A1 => n9469, A2 => n9468, Z => n39155);
   U20382 : OAI21_X2 port map( A1 => n32937, A2 => n12146, B => n38355, ZN => 
                           n17806);
   U20384 : AOI21_X2 port map( A1 => n36556, A2 => n19070, B => n17810, ZN => 
                           n38355);
   U20386 : NAND2_X1 port map( A1 => n1211, A2 => n5402, ZN => n6119);
   U20388 : NOR2_X2 port map( A1 => n32325, A2 => n38356, ZN => n18320);
   U20394 : NOR2_X2 port map( A1 => n38359, A2 => n38358, ZN => n38357);
   U20395 : INV_X2 port map( I => n25379, ZN => n38358);
   U20397 : INV_X2 port map( I => n10674, ZN => n38359);
   U20400 : XOR2_X1 port map( A1 => n38361, A2 => n38360, Z => n13759);
   U20404 : XOR2_X1 port map( A1 => n26539, A2 => n15508, Z => n38360);
   U20406 : XOR2_X1 port map( A1 => n39743, A2 => n26419, Z => n38361);
   U20409 : NAND2_X2 port map( A1 => n14618, A2 => n19852, ZN => n12227);
   U20419 : OR2_X2 port map( A1 => n25355, A2 => n24896, Z => n25389);
   U20420 : OAI22_X2 port map( A1 => n3962, A2 => n37103, B1 => n3135, B2 => 
                           n1090, ZN => n38435);
   U20421 : XOR2_X1 port map( A1 => n6658, A2 => n31724, Z => n32622);
   U20424 : INV_X2 port map( I => n5637, ZN => n12231);
   U20425 : XOR2_X1 port map( A1 => n28791, A2 => n6317, Z => n5637);
   U20428 : XOR2_X1 port map( A1 => n10401, A2 => n23945, Z => n10400);
   U20430 : NAND3_X1 port map( A1 => n33795, A2 => n2888, A3 => n3575, ZN => 
                           n38633);
   U20435 : XOR2_X1 port map( A1 => n33961, A2 => n20465, Z => n7936);
   U20437 : NAND3_X2 port map( A1 => n28521, A2 => n12947, A3 => n28520, ZN => 
                           n20465);
   U20439 : NAND2_X1 port map( A1 => n5671, A2 => n28285, ZN => n34516);
   U20440 : XOR2_X1 port map( A1 => n29049, A2 => n16355, Z => n4393);
   U20442 : XOR2_X1 port map( A1 => n1775, A2 => n16357, Z => n16355);
   U20445 : XOR2_X1 port map( A1 => n19608, A2 => n35196, Z => n3929);
   U20446 : XOR2_X1 port map( A1 => n19513, A2 => n29034, Z => n15216);
   U20447 : AOI22_X2 port map( A1 => n16474, A2 => n37311, B1 => n18836, B2 => 
                           n16475, ZN => n19513);
   U20448 : XOR2_X1 port map( A1 => n25046, A2 => n14563, Z => n5033);
   U20449 : AOI21_X2 port map( A1 => n6696, A2 => n1873, B => n38364, ZN => 
                           n39622);
   U20455 : XNOR2_X1 port map( A1 => n5208, A2 => n29538, ZN => n39720);
   U20456 : INV_X2 port map( I => n15922, ZN => n38365);
   U20462 : NAND2_X1 port map( A1 => n38367, A2 => n32472, ZN => n38366);
   U20463 : NOR2_X1 port map( A1 => n10272, A2 => n30716, ZN => n38368);
   U20464 : BUF_X2 port map( I => n933, Z => n38369);
   U20465 : XOR2_X1 port map( A1 => n38371, A2 => n1370, Z => Ciphertext(176));
   U20470 : OAI21_X2 port map( A1 => n13113, A2 => n13112, B => n1771, ZN => 
                           n23767);
   U20472 : NAND2_X2 port map( A1 => n35690, A2 => n14206, ZN => n1771);
   U20476 : XOR2_X1 port map( A1 => n8324, A2 => n38430, Z => n4894);
   U20478 : OAI21_X2 port map( A1 => n19707, A2 => n1372, B => n38372, ZN => 
                           n22234);
   U20483 : NAND2_X2 port map( A1 => n1372, A2 => n21755, ZN => n38372);
   U20485 : OAI21_X2 port map( A1 => n37143, A2 => n27163, B => n27164, ZN => 
                           n16997);
   U20486 : NOR2_X2 port map( A1 => n15391, A2 => n38374, ZN => n39200);
   U20492 : INV_X2 port map( I => n32107, ZN => n7955);
   U20495 : OAI22_X2 port map( A1 => n21553, A2 => n9886, B1 => n7954, B2 => 
                           n21719, ZN => n32107);
   U20499 : XNOR2_X1 port map( A1 => n21217, A2 => n20048, ZN => n38763);
   U20500 : NAND2_X1 port map( A1 => n22804, A2 => n14409, ZN => n32676);
   U20504 : OAI21_X2 port map( A1 => n8239, A2 => n13752, B => n38376, ZN => 
                           n10208);
   U20508 : BUF_X2 port map( I => n32623, Z => n38377);
   U20514 : XOR2_X1 port map( A1 => n32190, A2 => n18807, Z => n2526);
   U20515 : NAND2_X2 port map( A1 => n26113, A2 => n3642, ZN => n17269);
   U20522 : NAND2_X2 port map( A1 => n38476, A2 => n18349, ZN => n26113);
   U20528 : OAI22_X2 port map( A1 => n35902, A2 => n30671, B1 => n26966, B2 => 
                           n36234, ZN => n27825);
   U20531 : NAND3_X2 port map( A1 => n16621, A2 => n16634, A3 => n38378, ZN => 
                           n22744);
   U20532 : NAND2_X2 port map( A1 => n22136, A2 => n14196, ZN => n38378);
   U20533 : NOR2_X2 port map( A1 => n13601, A2 => n30304, ZN => n13598);
   U20534 : NAND3_X2 port map( A1 => n13600, A2 => n13599, A3 => n27874, ZN => 
                           n30304);
   U20535 : NOR2_X2 port map( A1 => n17869, A2 => n15868, ZN => n22275);
   U20536 : OAI22_X1 port map( A1 => n7515, A2 => n1121, B1 => n16210, B2 => 
                           n14283, ZN => n24780);
   U20537 : NAND3_X2 port map( A1 => n34167, A2 => n36159, A3 => n12326, ZN => 
                           n34535);
   U20542 : NAND2_X2 port map( A1 => n445, A2 => n5253, ZN => n39038);
   U20544 : XOR2_X1 port map( A1 => n7276, A2 => n38379, Z => n22879);
   U20548 : XOR2_X1 port map( A1 => n22745, A2 => n7275, Z => n38379);
   U20550 : XOR2_X1 port map( A1 => n6768, A2 => n39408, Z => n39008);
   U20553 : OR2_X1 port map( A1 => n36191, A2 => n34962, Z => n38380);
   U20556 : XOR2_X1 port map( A1 => n7288, A2 => n20460, Z => n9787);
   U20558 : NAND2_X1 port map( A1 => n5149, A2 => n20986, ZN => n39174);
   U20560 : INV_X2 port map( I => n38381, ZN => n36838);
   U20566 : NAND2_X2 port map( A1 => n38450, A2 => n34930, ZN => n38837);
   U20570 : AOI21_X2 port map( A1 => n37255, A2 => n32682, B => n38382, ZN => 
                           n38717);
   U20571 : NOR3_X2 port map( A1 => n7251, A2 => n36935, A3 => n9686, ZN => 
                           n38382);
   U20572 : NOR2_X2 port map( A1 => n38877, A2 => n27403, ZN => n34036);
   U20575 : AND2_X1 port map( A1 => n7485, A2 => n23577, Z => n38726);
   U20582 : XOR2_X1 port map( A1 => n38383, A2 => n13514, Z => n14758);
   U20583 : XOR2_X1 port map( A1 => n22518, A2 => n22519, Z => n38383);
   U20584 : XOR2_X1 port map( A1 => n29099, A2 => n12796, Z => n38384);
   U20585 : NAND2_X1 port map( A1 => n38751, A2 => n33384, ZN => n2062);
   U20588 : BUF_X4 port map( I => n33993, Z => n38448);
   U20589 : NAND2_X2 port map( A1 => n13494, A2 => n14768, ZN => n25179);
   U20594 : OAI21_X1 port map( A1 => n33128, A2 => n29676, B => n18042, ZN => 
                           n29679);
   U20595 : XOR2_X1 port map( A1 => n24014, A2 => n38385, Z => n13654);
   U20596 : NAND2_X2 port map( A1 => n38386, A2 => n16813, ZN => n26571);
   U20602 : NOR3_X2 port map( A1 => n38405, A2 => n38404, A3 => n34133, ZN => 
                           n38387);
   U20603 : NOR2_X1 port map( A1 => n5570, A2 => n921, ZN => n9249);
   U20607 : INV_X2 port map( I => n5638, ZN => n5570);
   U20611 : XOR2_X1 port map( A1 => n1914, A2 => n1911, Z => n5638);
   U20612 : NAND2_X2 port map( A1 => n38388, A2 => n23041, ZN => n23764);
   U20613 : NOR2_X2 port map( A1 => n32060, A2 => n4707, ZN => n38388);
   U20617 : OAI21_X2 port map( A1 => n38493, A2 => n38494, B => n21191, ZN => 
                           n13213);
   U20619 : NOR2_X2 port map( A1 => n23595, A2 => n23504, ZN => n38929);
   U20620 : NOR2_X2 port map( A1 => n24589, A2 => n31679, ZN => n24538);
   U20628 : NAND2_X2 port map( A1 => n5712, A2 => n5713, ZN => n24589);
   U20633 : XOR2_X1 port map( A1 => n9036, A2 => n33509, Z => n29087);
   U20634 : MUX2_X1 port map( I0 => n27897, I1 => n32002, S => n31664, Z => 
                           n27898);
   U20636 : NAND2_X2 port map( A1 => n16706, A2 => n7190, ZN => n31664);
   U20638 : XOR2_X1 port map( A1 => n10939, A2 => n10239, Z => n36406);
   U20640 : NAND2_X2 port map( A1 => n9166, A2 => n11248, ZN => n11818);
   U20641 : XOR2_X1 port map( A1 => n26302, A2 => n26303, Z => n26765);
   U20642 : XOR2_X1 port map( A1 => n7475, A2 => n30094, Z => n10100);
   U20645 : OAI22_X2 port map( A1 => n35477, A2 => n36103, B1 => n23589, B2 => 
                           n2273, ZN => n7475);
   U20649 : XOR2_X1 port map( A1 => n26391, A2 => n38140, Z => n7854);
   U20650 : NAND2_X2 port map( A1 => n32897, A2 => n13118, ZN => n26391);
   U20653 : NOR3_X1 port map( A1 => n22940, A2 => n33969, A3 => n6646, ZN => 
                           n38390);
   U20654 : XOR2_X1 port map( A1 => n33863, A2 => n22508, Z => n22765);
   U20657 : NOR2_X2 port map( A1 => n14957, A2 => n667, ZN => n22508);
   U20663 : XOR2_X1 port map( A1 => n38392, A2 => n39049, Z => n5211);
   U20671 : XOR2_X1 port map( A1 => n39344, A2 => n5667, Z => n38392);
   U20674 : NOR2_X2 port map( A1 => n26092, A2 => n26093, ZN => n25852);
   U20675 : NAND2_X2 port map( A1 => n4595, A2 => n31165, ZN => n26093);
   U20676 : NAND2_X2 port map( A1 => n10216, A2 => n32366, ZN => n23595);
   U20681 : NAND2_X2 port map( A1 => n400, A2 => n15492, ZN => n29231);
   U20682 : NAND2_X2 port map( A1 => n25047, A2 => n36690, ZN => n13843);
   U20684 : NAND2_X2 port map( A1 => n25048, A2 => n3510, ZN => n25047);
   U20685 : NAND2_X2 port map( A1 => n23502, A2 => n32366, ZN => n23374);
   U20687 : NAND2_X2 port map( A1 => n12254, A2 => n12253, ZN => n23502);
   U20692 : NAND2_X2 port map( A1 => n38394, A2 => n39051, ZN => n39050);
   U20698 : NAND2_X1 port map( A1 => n36623, A2 => n3944, ZN => n17715);
   U20701 : OAI21_X2 port map( A1 => n10587, A2 => n9648, B => n38396, ZN => 
                           n28521);
   U20702 : AOI21_X2 port map( A1 => n38529, A2 => n16295, B => n37081, ZN => 
                           n38396);
   U20707 : XOR2_X1 port map( A1 => n18991, A2 => n32765, Z => n14023);
   U20708 : NOR2_X2 port map( A1 => n12504, A2 => n12503, ZN => n18991);
   U20714 : NAND2_X2 port map( A1 => n38398, A2 => n36277, ZN => n26054);
   U20716 : XNOR2_X1 port map( A1 => n1790, A2 => n24062, ZN => n38975);
   U20717 : XOR2_X1 port map( A1 => n23898, A2 => n23968, Z => n23812);
   U20721 : NAND2_X2 port map( A1 => n23224, A2 => n23223, ZN => n23898);
   U20724 : INV_X2 port map( I => n17844, ZN => n20839);
   U20727 : XOR2_X1 port map( A1 => n32096, A2 => n18935, Z => n17844);
   U20733 : OAI21_X2 port map( A1 => n38400, A2 => n35880, B => n23141, ZN => 
                           n31908);
   U20734 : NAND3_X2 port map( A1 => n36911, A2 => n39414, A3 => n27240, ZN => 
                           n38525);
   U20736 : NAND2_X2 port map( A1 => n38401, A2 => n16305, ZN => n4391);
   U20740 : OAI21_X2 port map( A1 => n21570, A2 => n21599, B => n21870, ZN => 
                           n38401);
   U20757 : XOR2_X1 port map( A1 => n26595, A2 => n7018, Z => n26491);
   U20767 : XOR2_X1 port map( A1 => n4330, A2 => n32954, Z => n867);
   U20769 : XOR2_X1 port map( A1 => n29246, A2 => n38403, Z => n12069);
   U20773 : XOR2_X1 port map( A1 => n29832, A2 => n4905, Z => n38403);
   U20776 : XOR2_X1 port map( A1 => n29021, A2 => n29142, Z => n10430);
   U20779 : NAND3_X2 port map( A1 => n7849, A2 => n15602, A3 => n13422, ZN => 
                           n29021);
   U20780 : NOR2_X2 port map( A1 => n39366, A2 => n39365, ZN => n39364);
   U20781 : INV_X2 port map( I => n38406, ZN => n14179);
   U20784 : XNOR2_X1 port map( A1 => n9435, A2 => n38567, ZN => n38406);
   U20785 : NAND3_X2 port map( A1 => n32833, A2 => n19391, A3 => n1417, ZN => 
                           n1741);
   U20788 : NAND3_X2 port map( A1 => n39736, A2 => n5924, A3 => n5923, ZN => 
                           n17730);
   U20792 : AOI22_X2 port map( A1 => n31603, A2 => n12081, B1 => n39280, B2 => 
                           n19544, ZN => n3464);
   U20793 : AOI22_X2 port map( A1 => n31764, A2 => n12156, B1 => n27226, B2 => 
                           n10461, ZN => n5983);
   U20796 : NOR2_X2 port map( A1 => n10051, A2 => n27184, ZN => n27226);
   U20797 : OR2_X1 port map( A1 => n25782, A2 => n26106, Z => n11581);
   U20800 : OAI21_X2 port map( A1 => n11442, A2 => n11589, B => n11441, ZN => 
                           n25782);
   U20807 : AOI22_X2 port map( A1 => n3899, A2 => n28570, B1 => n3903, B2 => 
                           n33995, ZN => n4002);
   U20808 : XOR2_X1 port map( A1 => n24053, A2 => n23963, Z => n23928);
   U20814 : NAND2_X2 port map( A1 => n34421, A2 => n38859, ZN => n24053);
   U20816 : NAND2_X2 port map( A1 => n31719, A2 => n26122, ZN => n38409);
   U20820 : XOR2_X1 port map( A1 => n38410, A2 => n16268, Z => n36463);
   U20825 : XOR2_X1 port map( A1 => n36687, A2 => n6795, Z => n38410);
   U20827 : XOR2_X1 port map( A1 => n10226, A2 => n38411, Z => n39511);
   U20830 : XOR2_X1 port map( A1 => n27531, A2 => n27505, Z => n38411);
   U20832 : XOR2_X1 port map( A1 => n24064, A2 => n24002, Z => n11267);
   U20837 : NAND2_X2 port map( A1 => n23019, A2 => n23018, ZN => n24064);
   U20838 : NOR2_X2 port map( A1 => n196, A2 => n1688, ZN => n13009);
   U20841 : OR2_X2 port map( A1 => n38412, A2 => n10821, Z => n10820);
   U20843 : AOI21_X1 port map( A1 => n9466, A2 => n10875, B => n20810, ZN => 
                           n38412);
   U20844 : AOI21_X2 port map( A1 => n2339, A2 => n8154, B => n38413, ZN => 
                           n38908);
   U20847 : NOR2_X1 port map( A1 => n13371, A2 => n4748, ZN => n38413);
   U20862 : NAND4_X2 port map( A1 => n26913, A2 => n26914, A3 => n26915, A4 => 
                           n18749, ZN => n27700);
   U20868 : NAND2_X2 port map( A1 => n1891, A2 => n38414, ZN => n18749);
   U20870 : INV_X2 port map( I => n38415, ZN => n21644);
   U20872 : XNOR2_X1 port map( A1 => n21399, A2 => Key(183), ZN => n38415);
   U20877 : INV_X2 port map( I => n9303, ZN => n25753);
   U20879 : NAND2_X2 port map( A1 => n25754, A2 => n25699, ZN => n9303);
   U20881 : XOR2_X1 port map( A1 => n14218, A2 => n13883, Z => n12884);
   U20885 : XOR2_X1 port map( A1 => n36566, A2 => n27767, Z => n14218);
   U20886 : XOR2_X1 port map( A1 => n9001, A2 => n17263, Z => n26570);
   U20891 : NOR2_X2 port map( A1 => n13387, A2 => n13388, ZN => n9001);
   U20897 : XOR2_X1 port map( A1 => n35257, A2 => n30063, Z => n18736);
   U20898 : OAI21_X1 port map( A1 => n3361, A2 => n3360, B => n35646, ZN => 
                           n35257);
   U20899 : INV_X2 port map( I => n29160, ZN => n973);
   U20900 : NAND2_X2 port map( A1 => n39364, A2 => n35351, ZN => n29160);
   U20902 : AOI21_X2 port map( A1 => n24175, A2 => n24328, B => n6585, ZN => 
                           n11373);
   U20904 : NAND2_X2 port map( A1 => n38417, A2 => n14006, ZN => n15373);
   U20905 : NAND3_X2 port map( A1 => n1653, A2 => n6646, A3 => n38725, ZN => 
                           n38417);
   U20911 : INV_X2 port map( I => n9108, ZN => n1184);
   U20912 : XNOR2_X1 port map( A1 => n25298, A2 => n25113, ZN => n25144);
   U20916 : NOR2_X1 port map( A1 => n38418, A2 => n2785, ZN => n2784);
   U20917 : NOR2_X1 port map( A1 => n2788, A2 => n33646, ZN => n38418);
   U20919 : NAND2_X1 port map( A1 => n3443, A2 => n7935, ZN => n4058);
   U20920 : XOR2_X1 port map( A1 => Plaintext(186), A2 => Key(186), Z => n7935)
                           ;
   U20921 : NAND2_X2 port map( A1 => n33224, A2 => n38421, ZN => n32831);
   U20926 : NOR2_X2 port map( A1 => n38423, A2 => n38422, ZN => n38421);
   U20927 : NOR2_X2 port map( A1 => n24155, A2 => n9101, ZN => n38423);
   U20932 : OAI21_X1 port map( A1 => n21464, A2 => n21463, B => n21645, ZN => 
                           n9495);
   U20933 : OAI21_X2 port map( A1 => n8264, A2 => n1570, B => n30843, ZN => 
                           n38424);
   U20934 : NAND2_X2 port map( A1 => n20122, A2 => n39690, ZN => n3575);
   U20936 : XOR2_X1 port map( A1 => n19071, A2 => n23696, Z => n6943);
   U20940 : BUF_X4 port map( I => n39648, Z => n38561);
   U20943 : NAND3_X2 port map( A1 => n38426, A2 => n25416, A3 => n38425, ZN => 
                           n25509);
   U20945 : NAND2_X2 port map( A1 => n9740, A2 => n38178, ZN => n38426);
   U20947 : INV_X4 port map( I => n26029, ZN => n16867);
   U20948 : NOR2_X2 port map( A1 => n23120, A2 => n15947, ZN => n31364);
   U20949 : NOR3_X2 port map( A1 => n37074, A2 => n26799, A3 => n35282, ZN => 
                           n38755);
   U20956 : NOR2_X2 port map( A1 => n849, A2 => n4138, ZN => n26799);
   U20960 : NAND3_X2 port map( A1 => n36393, A2 => n23627, A3 => n36394, ZN => 
                           n33672);
   U20961 : NAND2_X2 port map( A1 => n2560, A2 => n2557, ZN => n29617);
   U20966 : NAND2_X2 port map( A1 => n23303, A2 => n11970, ZN => n23489);
   U20971 : XOR2_X1 port map( A1 => n34788, A2 => n24970, Z => n38427);
   U20972 : INV_X2 port map( I => n38428, ZN => n25307);
   U20976 : XNOR2_X1 port map( A1 => n12592, A2 => n12594, ZN => n38428);
   U20977 : NAND3_X1 port map( A1 => n36737, A2 => n36739, A3 => n30211, ZN => 
                           n38429);
   U20979 : OAI21_X2 port map( A1 => n11714, A2 => n10013, B => n24638, ZN => 
                           n11713);
   U20980 : NAND2_X2 port map( A1 => n35960, A2 => n3120, ZN => n24638);
   U20981 : XOR2_X1 port map( A1 => n1561, A2 => n25301, Z => n8324);
   U20986 : XOR2_X1 port map( A1 => n36138, A2 => n20333, Z => n33505);
   U20991 : NAND2_X1 port map( A1 => n3568, A2 => n25728, ZN => n25729);
   U20993 : NOR2_X1 port map( A1 => n14337, A2 => n29722, ZN => n29709);
   U20996 : NAND2_X2 port map( A1 => n1082, A2 => n38211, ZN => n26807);
   U21000 : XOR2_X1 port map( A1 => n10012, A2 => n25136, Z => n25272);
   U21003 : XOR2_X1 port map( A1 => n29045, A2 => n29040, Z => n18813);
   U21005 : NOR2_X2 port map( A1 => n21145, A2 => n20735, ZN => n29040);
   U21010 : AOI21_X1 port map( A1 => n28079, A2 => n987, B => n883, ZN => n7220
                           );
   U21011 : NAND2_X2 port map( A1 => n1252, A2 => n7986, ZN => n39294);
   U21029 : XOR2_X1 port map( A1 => n16833, A2 => n15974, Z => n15973);
   U21030 : XOR2_X1 port map( A1 => n38433, A2 => n34223, Z => n8184);
   U21035 : XOR2_X1 port map( A1 => n16019, A2 => n35728, Z => n38433);
   U21039 : OR2_X1 port map( A1 => n19135, A2 => n39050, Z => n35617);
   U21041 : XOR2_X1 port map( A1 => n20706, A2 => n38620, Z => n2283);
   U21047 : XOR2_X1 port map( A1 => n3035, A2 => n38434, Z => n3974);
   U21049 : XOR2_X1 port map( A1 => n14784, A2 => n26483, Z => n38434);
   U21052 : INV_X2 port map( I => n4008, ZN => n1120);
   U21083 : NAND2_X2 port map( A1 => n32018, A2 => n36542, ZN => n4008);
   U21084 : NOR2_X1 port map( A1 => n17934, A2 => n10523, ZN => n10524);
   U21085 : XOR2_X1 port map( A1 => n17920, A2 => n17922, Z => n17934);
   U21089 : XOR2_X1 port map( A1 => n26391, A2 => n10225, Z => n15288);
   U21099 : AOI22_X2 port map( A1 => n21421, A2 => n10924, B1 => n21983, B2 => 
                           n37176, ZN => n33736);
   U21102 : XOR2_X1 port map( A1 => n13978, A2 => n16324, Z => n13977);
   U21112 : NAND2_X2 port map( A1 => n11529, A2 => n11530, ZN => n16324);
   U21113 : NAND2_X2 port map( A1 => n30795, A2 => n7978, ZN => n30539);
   U21114 : NOR2_X2 port map( A1 => n36626, A2 => n38436, ZN => n39098);
   U21115 : AOI22_X2 port map( A1 => n626, A2 => n10342, B1 => n11673, B2 => 
                           n3398, ZN => n38436);
   U21116 : XOR2_X1 port map( A1 => n27809, A2 => n27615, Z => n8336);
   U21117 : XOR2_X1 port map( A1 => n27542, A2 => n6033, Z => n27809);
   U21118 : NAND2_X2 port map( A1 => n39357, A2 => n4339, ZN => n34195);
   U21129 : NAND2_X2 port map( A1 => n38439, A2 => n38438, ZN => n9539);
   U21130 : INV_X1 port map( I => n7982, ZN => n38438);
   U21131 : XOR2_X1 port map( A1 => n37338, A2 => n16162, Z => n38440);
   U21133 : OR2_X2 port map( A1 => n36868, A2 => n36355, Z => n3574);
   U21135 : XOR2_X1 port map( A1 => n19830, A2 => n20779, Z => n9780);
   U21137 : INV_X1 port map( I => n23349, ZN => n38441);
   U21140 : NOR2_X2 port map( A1 => n10724, A2 => n38953, ZN => n4248);
   U21141 : INV_X2 port map( I => n20691, ZN => n39023);
   U21143 : NAND2_X2 port map( A1 => n38618, A2 => n4014, ZN => n20691);
   U21145 : OAI21_X2 port map( A1 => n37203, A2 => n38463, B => n38442, ZN => 
                           n12741);
   U21151 : AOI22_X2 port map( A1 => n10910, A2 => n34737, B1 => n10908, B2 => 
                           n28608, ZN => n38442);
   U21156 : NAND3_X1 port map( A1 => n11039, A2 => n13753, A3 => n35114, ZN => 
                           n26844);
   U21157 : XOR2_X1 port map( A1 => n13193, A2 => n6561, Z => n31581);
   U21158 : NAND2_X2 port map( A1 => n12822, A2 => n9968, ZN => n13193);
   U21159 : OAI22_X2 port map( A1 => n10458, A2 => n10457, B1 => n17502, B2 => 
                           n12522, ZN => n31293);
   U21170 : AOI21_X2 port map( A1 => n33264, A2 => n34598, B => n38444, ZN => 
                           n24661);
   U21171 : OAI22_X2 port map( A1 => n7086, A2 => n15968, B1 => n14004, B2 => 
                           n24403, ZN => n38444);
   U21176 : NAND2_X2 port map( A1 => n35258, A2 => n36865, ZN => n38638);
   U21177 : AOI22_X2 port map( A1 => n25445, A2 => n32520, B1 => n33011, B2 => 
                           n33815, ZN => n38672);
   U21179 : XOR2_X1 port map( A1 => n3609, A2 => n5323, Z => n23959);
   U21182 : NAND2_X2 port map( A1 => n35864, A2 => n4251, ZN => n3609);
   U21184 : INV_X2 port map( I => n38445, ZN => n1230);
   U21185 : AND2_X1 port map( A1 => n32043, A2 => n9958, Z => n36995);
   U21188 : XOR2_X1 port map( A1 => n18547, A2 => n12304, Z => n32043);
   U21189 : XNOR2_X1 port map( A1 => n12969, A2 => n15500, ZN => n39245);
   U21190 : NAND2_X2 port map( A1 => n33187, A2 => n38446, ZN => n32898);
   U21194 : NAND2_X1 port map( A1 => n367, A2 => n39176, ZN => n4495);
   U21196 : AOI21_X2 port map( A1 => n22262, A2 => n33738, B => n33086, ZN => 
                           n4339);
   U21199 : INV_X4 port map( I => n33748, ZN => n33086);
   U21200 : AOI22_X2 port map( A1 => n36578, A2 => n15099, B1 => n34048, B2 => 
                           n15096, ZN => n33748);
   U21202 : OAI22_X2 port map( A1 => n31147, A2 => n32012, B1 => n28614, B2 => 
                           n4002, ZN => n5115);
   U21203 : XOR2_X1 port map( A1 => n39282, A2 => n5114, Z => n31329);
   U21204 : OR2_X1 port map( A1 => n5112, A2 => n3675, Z => n32449);
   U21207 : OR2_X2 port map( A1 => n21722, A2 => n3507, Z => n11852);
   U21209 : OAI22_X2 port map( A1 => n28652, A2 => n35830, B1 => n28650, B2 => 
                           n30931, ZN => n13027);
   U21210 : NAND3_X2 port map( A1 => n14750, A2 => n14749, A3 => n22995, ZN => 
                           n14748);
   U21212 : NAND2_X2 port map( A1 => n6674, A2 => n20449, ZN => n14750);
   U21218 : AOI22_X2 port map( A1 => n11331, A2 => n4642, B1 => n11333, B2 => 
                           n13015, ZN => n31367);
   U21220 : AOI22_X2 port map( A1 => n39226, A2 => n579, B1 => n32684, B2 => 
                           n31721, ZN => n5787);
   U21222 : NOR2_X2 port map( A1 => n12675, A2 => n12931, ZN => n579);
   U21223 : NAND3_X2 port map( A1 => n26979, A2 => n17252, A3 => n17097, ZN => 
                           n38450);
   U21228 : XOR2_X1 port map( A1 => n28933, A2 => n28869, Z => n36706);
   U21231 : XOR2_X1 port map( A1 => n18785, A2 => n29070, Z => n28933);
   U21235 : OAI21_X2 port map( A1 => n23182, A2 => n32270, B => n37137, ZN => 
                           n23183);
   U21239 : NAND2_X2 port map( A1 => n38451, A2 => n15583, ZN => n31751);
   U21243 : NAND3_X2 port map( A1 => n39585, A2 => n38834, A3 => n38328, ZN => 
                           n38451);
   U21246 : OR2_X1 port map( A1 => n24473, A2 => n7240, Z => n38474);
   U21252 : NAND2_X2 port map( A1 => n28066, A2 => n14500, ZN => n5430);
   U21254 : AND2_X1 port map( A1 => n20077, A2 => n32537, Z => n22940);
   U21255 : CLKBUF_X4 port map( I => n26833, Z => n38852);
   U21263 : INV_X4 port map( I => n38452, ZN => n15573);
   U21265 : AND3_X2 port map( A1 => n11648, A2 => n11649, A3 => n15446, Z => 
                           n38452);
   U21266 : XOR2_X1 port map( A1 => n34876, A2 => n36114, Z => n38453);
   U21269 : XOR2_X1 port map( A1 => n28949, A2 => n28950, Z => n33434);
   U21271 : XOR2_X1 port map( A1 => n38454, A2 => n19810, Z => n26803);
   U21273 : XOR2_X1 port map( A1 => n25986, A2 => n25985, Z => n38454);
   U21274 : XOR2_X1 port map( A1 => n32613, A2 => n11401, Z => n38455);
   U21279 : AOI21_X2 port map( A1 => n7978, A2 => n30795, B => n26700, ZN => 
                           n32262);
   U21280 : NAND2_X2 port map( A1 => n39144, A2 => n38456, ZN => n33258);
   U21282 : OAI21_X2 port map( A1 => n39223, A2 => n39224, B => n7986, ZN => 
                           n38456);
   U21287 : NOR2_X2 port map( A1 => n4427, A2 => n4062, ZN => n25146);
   U21290 : XOR2_X1 port map( A1 => n31227, A2 => n476, Z => n4612);
   U21292 : XOR2_X1 port map( A1 => n13649, A2 => n38457, Z => n19658);
   U21293 : XOR2_X1 port map( A1 => n23723, A2 => n23741, Z => n38457);
   U21294 : XOR2_X1 port map( A1 => n24992, A2 => n15186, Z => n38458);
   U21295 : XOR2_X1 port map( A1 => n39163, A2 => n23675, Z => n34269);
   U21299 : NAND2_X2 port map( A1 => n34884, A2 => n20984, ZN => n23675);
   U21303 : NAND2_X1 port map( A1 => n20619, A2 => n24470, ZN => n36790);
   U21304 : NAND2_X2 port map( A1 => n39643, A2 => n28392, ZN => n6093);
   U21305 : NOR2_X2 port map( A1 => n38460, A2 => n38459, ZN => n19260);
   U21307 : AOI21_X2 port map( A1 => n18997, A2 => n31583, B => n29587, ZN => 
                           n38459);
   U21308 : AOI21_X2 port map( A1 => n20371, A2 => n29630, B => n21264, ZN => 
                           n38460);
   U21309 : XOR2_X1 port map( A1 => n37874, A2 => n15682, Z => n28845);
   U21310 : XNOR2_X1 port map( A1 => n29048, A2 => n19843, ZN => n38606);
   U21311 : NAND2_X2 port map( A1 => n1904, A2 => n21287, ZN => n6601);
   U21312 : OAI22_X2 port map( A1 => n11861, A2 => n29946, B1 => n16510, B2 => 
                           n17240, ZN => n1904);
   U21315 : XOR2_X1 port map( A1 => n18001, A2 => n14173, Z => n9943);
   U21321 : XOR2_X1 port map( A1 => n27777, A2 => n38158, Z => n5524);
   U21342 : XOR2_X1 port map( A1 => n18160, A2 => n23707, Z => n23997);
   U21343 : AOI21_X2 port map( A1 => n9971, A2 => n1307, B => n23442, ZN => 
                           n18160);
   U21347 : AOI22_X2 port map( A1 => n22977, A2 => n10828, B1 => n10470, B2 => 
                           n7266, ZN => n10469);
   U21350 : NAND3_X2 port map( A1 => n33669, A2 => n17532, A3 => n28163, ZN => 
                           n31882);
   U21355 : NOR2_X1 port map( A1 => n4713, A2 => n38513, ZN => n15947);
   U21356 : AOI21_X1 port map( A1 => n7789, A2 => n10702, B => n29059, ZN => 
                           n11777);
   U21358 : NAND2_X2 port map( A1 => n2182, A2 => n36720, ZN => n23373);
   U21361 : XOR2_X1 port map( A1 => n38462, A2 => n1161, Z => Ciphertext(171));
   U21366 : OAI21_X1 port map( A1 => n39079, A2 => n2506, B => n2945, ZN => 
                           n2203);
   U21370 : INV_X2 port map( I => n35813, ZN => n24788);
   U21371 : OR2_X1 port map( A1 => n12246, A2 => n31682, Z => n12192);
   U21372 : XOR2_X1 port map( A1 => n38464, A2 => n25090, Z => n25159);
   U21374 : INV_X2 port map( I => n25133, ZN => n38464);
   U21379 : NAND2_X2 port map( A1 => n7064, A2 => n31290, ZN => n25090);
   U21380 : XOR2_X1 port map( A1 => n14719, A2 => n38465, Z => n39277);
   U21386 : NAND2_X2 port map( A1 => n38466, A2 => n13870, ZN => n34644);
   U21387 : NOR2_X2 port map( A1 => n31705, A2 => n11800, ZN => n11695);
   U21388 : AOI22_X2 port map( A1 => n1077, A2 => n9315, B1 => n20976, B2 => 
                           n10573, ZN => n10579);
   U21389 : NAND2_X2 port map( A1 => n1570, A2 => n257, ZN => n12124);
   U21392 : XOR2_X1 port map( A1 => n24711, A2 => n25192, Z => n20554);
   U21395 : INV_X2 port map( I => n38467, ZN => n8479);
   U21396 : NAND2_X2 port map( A1 => n39131, A2 => n12133, ZN => n11698);
   U21405 : NOR2_X2 port map( A1 => n36964, A2 => n10708, ZN => n35181);
   U21408 : XOR2_X1 port map( A1 => n22635, A2 => n22633, Z => n32847);
   U21410 : XOR2_X1 port map( A1 => n22776, A2 => n22731, Z => n22633);
   U21411 : NOR2_X1 port map( A1 => n36786, A2 => n36787, ZN => n39731);
   U21419 : AOI21_X2 port map( A1 => n11424, A2 => n20336, B => n11423, ZN => 
                           n26278);
   U21426 : NAND3_X2 port map( A1 => n20470, A2 => n39382, A3 => n27620, ZN => 
                           n20662);
   U21428 : INV_X2 port map( I => n38470, ZN => n28188);
   U21429 : NAND2_X1 port map( A1 => n5101, A2 => n7542, ZN => n36981);
   U21437 : AOI21_X2 port map( A1 => n10521, A2 => n20064, B => n10159, ZN => 
                           n10520);
   U21439 : XOR2_X1 port map( A1 => n18133, A2 => n38471, Z => n38927);
   U21440 : XOR2_X1 port map( A1 => n29113, A2 => n29983, Z => n38471);
   U21442 : XOR2_X1 port map( A1 => n29105, A2 => n16529, Z => n12402);
   U21443 : NAND2_X1 port map( A1 => n32649, A2 => n32648, ZN => n39722);
   U21444 : NAND2_X2 port map( A1 => n38474, A2 => n38472, ZN => n10626);
   U21447 : NAND2_X2 port map( A1 => n1081, A2 => n3851, ZN => n3850);
   U21452 : OR2_X2 port map( A1 => n28204, A2 => n21159, Z => n9089);
   U21457 : XOR2_X1 port map( A1 => n38205, A2 => n15219, Z => n10412);
   U21460 : NOR2_X2 port map( A1 => n38910, A2 => n3849, ZN => n15219);
   U21461 : XOR2_X1 port map( A1 => n5412, A2 => n33701, Z => n5410);
   U21463 : NOR2_X2 port map( A1 => n12447, A2 => n24174, ZN => n39480);
   U21465 : NAND2_X2 port map( A1 => n1607, A2 => n37954, ZN => n12447);
   U21467 : NOR2_X2 port map( A1 => n38475, A2 => n34042, ZN => n12676);
   U21471 : XOR2_X1 port map( A1 => n12973, A2 => n24058, Z => n9548);
   U21473 : XOR2_X1 port map( A1 => n2443, A2 => n1502, Z => n2545);
   U21479 : OAI21_X2 port map( A1 => n32712, A2 => n15284, B => n12031, ZN => 
                           n21140);
   U21494 : AOI21_X2 port map( A1 => n8393, A2 => n2629, B => n1742, ZN => 
                           n35209);
   U21498 : AOI21_X2 port map( A1 => n2865, A2 => n17269, B => n930, ZN => 
                           n1742);
   U21500 : NAND2_X2 port map( A1 => n38478, A2 => n30850, ZN => n24799);
   U21504 : XOR2_X1 port map( A1 => n27760, A2 => n27413, Z => n38624);
   U21505 : XOR2_X1 port map( A1 => n27731, A2 => n7755, Z => n27413);
   U21507 : NAND2_X2 port map( A1 => n38479, A2 => n39592, ZN => n2668);
   U21509 : XOR2_X1 port map( A1 => n27778, A2 => n21093, Z => n27515);
   U21516 : NAND2_X2 port map( A1 => n10953, A2 => n36492, ZN => n21093);
   U21520 : XOR2_X1 port map( A1 => n29257, A2 => n29085, Z => n17659);
   U21522 : XOR2_X1 port map( A1 => n24030, A2 => n23883, Z => n24001);
   U21525 : NOR2_X2 port map( A1 => n1302, A2 => n1297, ZN => n8390);
   U21526 : NAND2_X2 port map( A1 => n23467, A2 => n16528, ZN => n18989);
   U21528 : NOR2_X2 port map( A1 => n38559, A2 => n6970, ZN => n23467);
   U21529 : NAND2_X2 port map( A1 => n14496, A2 => n20576, ZN => n36969);
   U21530 : XOR2_X1 port map( A1 => n20695, A2 => n24056, Z => n39201);
   U21531 : XOR2_X1 port map( A1 => n1613, A2 => n16138, Z => n20695);
   U21533 : XOR2_X1 port map( A1 => n39078, A2 => n17650, Z => n19443);
   U21541 : OAI21_X2 port map( A1 => n31470, A2 => n31471, B => n10511, ZN => 
                           n17650);
   U21542 : XOR2_X1 port map( A1 => n38485, A2 => n22506, Z => n2046);
   U21557 : XOR2_X1 port map( A1 => n16912, A2 => n22701, Z => n38485);
   U21561 : XOR2_X1 port map( A1 => n20205, A2 => n24011, Z => n23729);
   U21564 : NAND2_X2 port map( A1 => n7482, A2 => n23422, ZN => n20205);
   U21566 : XOR2_X1 port map( A1 => n38510, A2 => n15857, Z => n39285);
   U21568 : XOR2_X1 port map( A1 => n38486, A2 => n7558, Z => n12519);
   U21569 : XOR2_X1 port map( A1 => n25031, A2 => n32433, Z => n25167);
   U21572 : NAND2_X2 port map( A1 => n17916, A2 => n4937, ZN => n38493);
   U21573 : BUF_X2 port map( I => n17263, Z => n38495);
   U21578 : NAND2_X1 port map( A1 => n9836, A2 => n11777, ZN => n39586);
   U21581 : OAI21_X2 port map( A1 => n123, A2 => n683, B => n38496, ZN => 
                           n32763);
   U21585 : XOR2_X1 port map( A1 => n3495, A2 => n38497, Z => n8128);
   U21592 : XOR2_X1 port map( A1 => n32346, A2 => n3493, Z => n38497);
   U21595 : NAND2_X2 port map( A1 => n9242, A2 => n36197, ZN => n3983);
   U21596 : BUF_X1 port map( I => n6002, Z => n35264);
   U21598 : INV_X2 port map( I => n38854, ZN => n3899);
   U21602 : AOI22_X2 port map( A1 => n2614, A2 => n17532, B1 => n33669, B2 => 
                           n2613, ZN => n38596);
   U21604 : INV_X2 port map( I => n23550, ZN => n38499);
   U21616 : AOI21_X2 port map( A1 => n35191, A2 => n38499, B => n37814, ZN => 
                           n38615);
   U21620 : INV_X2 port map( I => n30981, ZN => n27366);
   U21621 : NAND2_X2 port map( A1 => n21101, A2 => n27363, ZN => n30981);
   U21622 : XOR2_X1 port map( A1 => n8059, A2 => n27862, Z => n27642);
   U21625 : BUF_X2 port map( I => n26551, Z => n38502);
   U21626 : OAI21_X2 port map( A1 => n37249, A2 => n38503, B => n9598, ZN => 
                           n34463);
   U21627 : AND2_X1 port map( A1 => n32080, A2 => n36463, Z => n28288);
   U21628 : NOR2_X2 port map( A1 => n33752, A2 => n6589, ZN => n26481);
   U21629 : OAI21_X2 port map( A1 => n4371, A2 => n4369, B => n38504, ZN => 
                           n28305);
   U21634 : XOR2_X1 port map( A1 => n38624, A2 => n38505, Z => n17777);
   U21639 : XOR2_X1 port map( A1 => n12165, A2 => n27495, Z => n38505);
   U21650 : INV_X2 port map( I => n24812, ZN => n32651);
   U21651 : XOR2_X1 port map( A1 => n10767, A2 => n13483, Z => n13090);
   U21654 : XOR2_X1 port map( A1 => n6384, A2 => n11753, Z => n13483);
   U21660 : AOI22_X2 port map( A1 => n28282, A2 => n28283, B1 => n36877, B2 => 
                           n16544, ZN => n12787);
   U21664 : NAND2_X2 port map( A1 => n33314, A2 => n38487, ZN => n24121);
   U21666 : XOR2_X1 port map( A1 => n27749, A2 => n38225, Z => n3889);
   U21674 : XOR2_X1 port map( A1 => n33645, A2 => n30170, Z => n10492);
   U21676 : INV_X4 port map( I => n19255, ZN => n31698);
   U21677 : NAND2_X2 port map( A1 => n24455, A2 => n24456, ZN => n19255);
   U21678 : NAND2_X2 port map( A1 => n5264, A2 => n16859, ZN => n27379);
   U21684 : AND2_X1 port map( A1 => n585, A2 => n17871, Z => n35075);
   U21693 : OAI22_X2 port map( A1 => n15445, A2 => n25362, B1 => n15444, B2 => 
                           n19095, ZN => n35003);
   U21694 : OAI21_X2 port map( A1 => n28187, A2 => n14642, B => n33002, ZN => 
                           n38506);
   U21696 : NOR2_X2 port map( A1 => n9969, A2 => n28191, ZN => n28187);
   U21697 : NAND2_X2 port map( A1 => n38506, A2 => n14030, ZN => n13594);
   U21698 : NAND2_X2 port map( A1 => n13492, A2 => n38947, ZN => n38946);
   U21700 : XOR2_X1 port map( A1 => n24961, A2 => n13634, Z => n25262);
   U21701 : NAND2_X2 port map( A1 => n62, A2 => n35022, ZN => n13634);
   U21702 : XOR2_X1 port map( A1 => n12749, A2 => n15265, Z => n15261);
   U21707 : NAND2_X1 port map( A1 => n3016, A2 => n24178, ZN => n38508);
   U21708 : NAND3_X2 port map( A1 => n18202, A2 => n28746, A3 => n18201, ZN => 
                           n19408);
   U21710 : XOR2_X1 port map( A1 => n19561, A2 => n35229, Z => n4266);
   U21711 : XOR2_X1 port map( A1 => n23688, A2 => n34435, Z => n2695);
   U21712 : NOR2_X2 port map( A1 => n38509, A2 => n35944, ZN => n12910);
   U21718 : XOR2_X1 port map( A1 => n25154, A2 => n38511, Z => n38510);
   U21720 : XOR2_X1 port map( A1 => n11756, A2 => n12233, Z => n24610);
   U21723 : NAND3_X1 port map( A1 => n15541, A2 => n37050, A3 => n826, ZN => 
                           n12578);
   U21725 : CLKBUF_X2 port map( I => n22929, Z => n39518);
   U21729 : NAND2_X2 port map( A1 => n38549, A2 => n13454, ZN => n8412);
   U21731 : NAND2_X2 port map( A1 => n30302, A2 => n2029, ZN => n26114);
   U21740 : NAND2_X2 port map( A1 => n31964, A2 => n31963, ZN => n2029);
   U21747 : BUF_X2 port map( I => n26530, Z => n38514);
   U21751 : XOR2_X1 port map( A1 => n15401, A2 => n38515, Z => n27474);
   U21755 : NAND2_X2 port map( A1 => n11855, A2 => n13211, ZN => n15401);
   U21757 : XOR2_X1 port map( A1 => n27542, A2 => n37101, Z => n39515);
   U21760 : NAND2_X1 port map( A1 => n16444, A2 => n25767, ZN => n34595);
   U21765 : NAND2_X1 port map( A1 => n28322, A2 => n14448, ZN => n30380);
   U21766 : OAI21_X1 port map( A1 => n25488, A2 => n32775, B => n25487, ZN => 
                           n32879);
   U21767 : XOR2_X1 port map( A1 => n16696, A2 => n16698, Z => n34561);
   U21768 : NAND3_X2 port map( A1 => n38516, A2 => n38525, A3 => n27242, ZN => 
                           n27528);
   U21769 : XOR2_X1 port map( A1 => n38517, A2 => n38518, Z => n28182);
   U21770 : XOR2_X1 port map( A1 => n15844, A2 => n15785, Z => n38517);
   U21772 : XOR2_X1 port map( A1 => n27515, A2 => n763, Z => n38518);
   U21773 : NAND2_X2 port map( A1 => n12287, A2 => n24159, ZN => n24903);
   U21777 : OAI21_X2 port map( A1 => n30388, A2 => n25566, B => n38520, ZN => 
                           n14212);
   U21779 : OAI21_X2 port map( A1 => n33897, A2 => n15459, B => n10723, ZN => 
                           n38520);
   U21780 : INV_X1 port map( I => n25170, ZN => n1930);
   U21784 : BUF_X2 port map( I => n17101, Z => n38523);
   U21786 : BUF_X2 port map( I => n23190, Z => n38524);
   U21787 : NAND2_X2 port map( A1 => n18632, A2 => n38526, ZN => n17607);
   U21792 : NOR2_X2 port map( A1 => n35314, A2 => n9135, ZN => n38528);
   U21798 : NAND2_X2 port map( A1 => n12074, A2 => n8696, ZN => n32588);
   U21801 : INV_X2 port map( I => n14349, ZN => n22323);
   U21802 : NAND2_X2 port map( A1 => n21516, A2 => n16961, ZN => n14349);
   U21804 : XOR2_X1 port map( A1 => n11881, A2 => n38530, Z => n11880);
   U21807 : BUF_X2 port map( I => n5859, Z => n38531);
   U21808 : OAI22_X2 port map( A1 => n14535, A2 => n17537, B1 => n17536, B2 => 
                           n37920, ZN => n22411);
   U21813 : XOR2_X1 port map( A1 => n29092, A2 => n29096, Z => n29027);
   U21814 : NAND2_X2 port map( A1 => n35583, A2 => n14929, ZN => n29092);
   U21816 : XOR2_X1 port map( A1 => n32608, A2 => n28851, Z => n29073);
   U21817 : OAI21_X2 port map( A1 => n12608, A2 => n12609, B => n28524, ZN => 
                           n28851);
   U21818 : XOR2_X1 port map( A1 => n557, A2 => n34963, Z => n11828);
   U21819 : INV_X2 port map( I => n39810, ZN => n19082);
   U21827 : XOR2_X1 port map( A1 => n4658, A2 => n35129, Z => n33808);
   U21828 : AOI21_X2 port map( A1 => n1966, A2 => n22148, B => n1965, ZN => 
                           n359);
   U21833 : XOR2_X1 port map( A1 => n38532, A2 => n11922, Z => n11350);
   U21834 : XOR2_X1 port map( A1 => n9777, A2 => n5542, Z => n38532);
   U21835 : XOR2_X1 port map( A1 => n23835, A2 => n20486, Z => n17492);
   U21840 : NOR2_X1 port map( A1 => n32043, A2 => n36136, ZN => n28028);
   U21841 : XOR2_X1 port map( A1 => n23743, A2 => n18980, Z => n1969);
   U21842 : NOR3_X2 port map( A1 => n33793, A2 => n30334, A3 => n38533, ZN => 
                           n33116);
   U21847 : NOR3_X2 port map( A1 => n33629, A2 => n18281, A3 => n17735, ZN => 
                           n38533);
   U21856 : XOR2_X1 port map( A1 => n29294, A2 => n28957, Z => n5782);
   U21859 : XOR2_X1 port map( A1 => n16771, A2 => n29242, Z => n28957);
   U21864 : NAND2_X1 port map( A1 => n38535, A2 => n39001, ZN => n38534);
   U21866 : INV_X2 port map( I => n12396, ZN => n38535);
   U21874 : OAI21_X2 port map( A1 => n38537, A2 => n3899, B => n39020, ZN => 
                           n3390);
   U21876 : INV_X2 port map( I => n33995, ZN => n38537);
   U21883 : NAND2_X2 port map( A1 => n38713, A2 => n36472, ZN => n9802);
   U21884 : NAND2_X1 port map( A1 => n214, A2 => n38538, ZN => n2630);
   U21886 : NAND2_X1 port map( A1 => n20418, A2 => n38981, ZN => n38538);
   U21888 : OAI21_X1 port map( A1 => n27403, A2 => n36865, B => n994, ZN => 
                           n33887);
   U21890 : INV_X4 port map( I => n13730, ZN => n27403);
   U21892 : NAND3_X2 port map( A1 => n33567, A2 => n26816, A3 => n16573, ZN => 
                           n13730);
   U21893 : XOR2_X1 port map( A1 => n18600, A2 => n38192, Z => n16133);
   U21898 : XOR2_X1 port map( A1 => n33582, A2 => n38539, Z => n33601);
   U21902 : INV_X1 port map( I => n29043, ZN => n38539);
   U21906 : NAND2_X2 port map( A1 => n14286, A2 => n9714, ZN => n5848);
   U21911 : NAND2_X2 port map( A1 => n10323, A2 => n38540, ZN => n22353);
   U21918 : OAI22_X1 port map( A1 => n21867, A2 => n17948, B1 => n19549, B2 => 
                           n21868, ZN => n38540);
   U21920 : OAI22_X2 port map( A1 => n16887, A2 => n38541, B1 => n39526, B2 => 
                           n23056, ZN => n35915);
   U21922 : OAI22_X2 port map( A1 => n12710, A2 => n25862, B1 => n12712, B2 => 
                           n12711, ZN => n26227);
   U21926 : NOR2_X2 port map( A1 => n21181, A2 => n36846, ZN => n27484);
   U21927 : OAI22_X1 port map( A1 => n27332, A2 => n27333, B1 => n35115, B2 => 
                           n27331, ZN => n27336);
   U21928 : XOR2_X1 port map( A1 => n6427, A2 => n6430, Z => n20080);
   U21929 : AOI22_X2 port map( A1 => n7255, A2 => n39298, B1 => n37661, B2 => 
                           n9655, ZN => n31785);
   U21930 : OAI21_X2 port map( A1 => n5642, A2 => n14398, B => n34774, ZN => 
                           n33509);
   U21933 : NAND2_X2 port map( A1 => n15713, A2 => n15716, ZN => n39406);
   U21948 : NAND2_X2 port map( A1 => n35301, A2 => n2953, ZN => n23419);
   U21949 : XOR2_X1 port map( A1 => n751, A2 => n38543, Z => n851);
   U21950 : XOR2_X1 port map( A1 => n26441, A2 => n29718, Z => n38543);
   U21953 : NOR2_X2 port map( A1 => n39618, A2 => n38544, ZN => n18656);
   U21961 : NAND2_X2 port map( A1 => n38547, A2 => n38545, ZN => n38544);
   U21963 : XOR2_X1 port map( A1 => n20392, A2 => n11974, Z => n22452);
   U21965 : XOR2_X1 port map( A1 => n35209, A2 => n14346, Z => n5688);
   U21966 : NOR2_X2 port map( A1 => n14226, A2 => n14224, ZN => n14346);
   U21968 : NOR2_X2 port map( A1 => n20566, A2 => n29346, ZN => n39033);
   U21971 : INV_X2 port map( I => n13815, ZN => n20566);
   U21982 : XOR2_X1 port map( A1 => n9972, A2 => n11946, Z => n13815);
   U21985 : NOR2_X2 port map( A1 => n38551, A2 => n38550, ZN => n14088);
   U21986 : INV_X2 port map( I => n12199, ZN => n38551);
   U21987 : NAND2_X2 port map( A1 => n38552, A2 => n26090, ZN => n39158);
   U21991 : NAND2_X2 port map( A1 => n4852, A2 => n25882, ZN => n38552);
   U21993 : NOR2_X1 port map( A1 => n32682, A2 => n9686, ZN => n28625);
   U21997 : XOR2_X1 port map( A1 => n38553, A2 => n30781, Z => n31426);
   U21998 : XOR2_X1 port map( A1 => n27709, A2 => n27718, Z => n38553);
   U22000 : INV_X2 port map( I => n38554, ZN => n27894);
   U22002 : NAND2_X1 port map( A1 => n38611, A2 => n1627, ZN => n14746);
   U22007 : NOR2_X2 port map( A1 => n436, A2 => n39318, ZN => n6405);
   U22009 : XOR2_X1 port map( A1 => n38796, A2 => n12322, Z => n10029);
   U22010 : XOR2_X1 port map( A1 => n26288, A2 => n38753, Z => n12322);
   U22017 : NAND2_X2 port map( A1 => n25836, A2 => n19580, ZN => n25808);
   U22019 : XOR2_X1 port map( A1 => n24947, A2 => n24948, Z => n24949);
   U22021 : XOR2_X1 port map( A1 => n23902, A2 => n18160, Z => n6987);
   U22022 : AOI21_X2 port map( A1 => n4528, A2 => n1132, B => n4526, ZN => 
                           n23902);
   U22023 : XOR2_X1 port map( A1 => n8324, A2 => n15011, Z => n4869);
   U22035 : XNOR2_X1 port map( A1 => n25221, A2 => n31579, ZN => n38563);
   U22036 : BUF_X2 port map( I => n4108, Z => n38555);
   U22038 : NAND2_X2 port map( A1 => n38557, A2 => n22834, ZN => n33257);
   U22040 : INV_X2 port map( I => n22829, ZN => n38557);
   U22047 : NOR2_X2 port map( A1 => n39096, A2 => n33431, ZN => n22829);
   U22051 : INV_X4 port map( I => n38907, ZN => n13973);
   U22052 : XOR2_X1 port map( A1 => n28845, A2 => n38885, Z => n34477);
   U22053 : XNOR2_X1 port map( A1 => n38212, A2 => n1375, ZN => n39335);
   U22056 : INV_X1 port map( I => n6591, ZN => n37025);
   U22062 : XOR2_X1 port map( A1 => n6593, A2 => n38558, Z => n6591);
   U22063 : XOR2_X1 port map( A1 => n9979, A2 => n24070, Z => n208);
   U22064 : NAND2_X2 port map( A1 => n18485, A2 => n39056, ZN => n9979);
   U22073 : NOR2_X1 port map( A1 => n29752, A2 => n29751, ZN => n29758);
   U22075 : XOR2_X1 port map( A1 => n7710, A2 => n29833, Z => n7004);
   U22078 : AOI22_X2 port map( A1 => n2125, A2 => n2124, B1 => n32385, B2 => 
                           n36722, ZN => n19384);
   U22079 : NAND3_X1 port map( A1 => n24098, A2 => n20517, A3 => n20041, ZN => 
                           n6912);
   U22082 : XOR2_X1 port map( A1 => n35842, A2 => n38562, Z => n38966);
   U22083 : XOR2_X1 port map( A1 => n25222, A2 => n38563, Z => n38562);
   U22084 : XOR2_X1 port map( A1 => n3232, A2 => n38564, Z => n32599);
   U22085 : XOR2_X1 port map( A1 => n22690, A2 => n32331, Z => n38564);
   U22086 : NAND2_X2 port map( A1 => n38565, A2 => n27102, ZN => n36287);
   U22087 : XOR2_X1 port map( A1 => n28951, A2 => n5862, Z => n38567);
   U22090 : NOR2_X1 port map( A1 => n36633, A2 => n30805, ZN => n38924);
   U22091 : XOR2_X1 port map( A1 => n25249, A2 => n17623, Z => n38569);
   U22094 : NOR2_X2 port map( A1 => n36850, A2 => n2160, ZN => n12272);
   U22097 : INV_X1 port map( I => n29968, ZN => n5678);
   U22101 : NAND2_X2 port map( A1 => n34460, A2 => n39525, ZN => n29968);
   U22104 : NAND2_X2 port map( A1 => n38570, A2 => n31606, ZN => n9917);
   U22105 : NOR2_X2 port map( A1 => n32657, A2 => n33292, ZN => n38570);
   U22106 : NOR2_X1 port map( A1 => n25665, A2 => n20441, ZN => n19336);
   U22107 : XOR2_X1 port map( A1 => n11425, A2 => n3413, Z => n20540);
   U22111 : NOR2_X2 port map( A1 => n12456, A2 => n12458, ZN => n11425);
   U22112 : OAI21_X2 port map( A1 => n31530, A2 => n3112, B => n3111, ZN => 
                           n3110);
   U22114 : OAI21_X2 port map( A1 => n38060, A2 => n18228, B => n20671, ZN => 
                           n38572);
   U22117 : XOR2_X1 port map( A1 => n762, A2 => n2437, Z => n2436);
   U22119 : XOR2_X1 port map( A1 => n27546, A2 => n35998, Z => n762);
   U22120 : NOR2_X2 port map( A1 => n38573, A2 => n5738, ZN => n31656);
   U22134 : NOR2_X2 port map( A1 => n28712, A2 => n36414, ZN => n38573);
   U22142 : NAND2_X1 port map( A1 => n34254, A2 => n32468, ZN => n39777);
   U22144 : NOR2_X2 port map( A1 => n16682, A2 => n15867, ZN => n3377);
   U22148 : XOR2_X1 port map( A1 => n23997, A2 => n36233, Z => n39665);
   U22150 : INV_X2 port map( I => n38575, ZN => n34178);
   U22152 : XOR2_X1 port map( A1 => n38575, A2 => n29054, Z => n34091);
   U22157 : NAND2_X2 port map( A1 => n36585, A2 => n15312, ZN => n38575);
   U22162 : OAI21_X2 port map( A1 => n36342, A2 => n33101, B => n36341, ZN => 
                           n38576);
   U22163 : NAND2_X1 port map( A1 => n20793, A2 => n29769, ZN => n29770);
   U22164 : NAND2_X2 port map( A1 => n17373, A2 => n13389, ZN => n17263);
   U22165 : NOR2_X2 port map( A1 => n31393, A2 => n39453, ZN => n33961);
   U22169 : AND2_X1 port map( A1 => n7993, A2 => n14463, Z => n14655);
   U22173 : OR2_X2 port map( A1 => n38214, A2 => n14061, Z => n16773);
   U22177 : NAND2_X2 port map( A1 => n39464, A2 => n9608, ZN => n23535);
   U22178 : OAI21_X1 port map( A1 => n24764, A2 => n39098, B => n7852, ZN => 
                           n32221);
   U22179 : NAND2_X2 port map( A1 => n32035, A2 => n25808, ZN => n15298);
   U22182 : NAND2_X1 port map( A1 => n10141, A2 => n24793, ZN => n17106);
   U22184 : AOI22_X2 port map( A1 => n38582, A2 => n36920, B1 => n7261, B2 => 
                           n5888, ZN => n14874);
   U22185 : INV_X2 port map( I => n24579, ZN => n38582);
   U22190 : NAND2_X2 port map( A1 => n5137, A2 => n32091, ZN => n24579);
   U22191 : NAND2_X2 port map( A1 => n30173, A2 => n30172, ZN => n4368);
   U22192 : NAND2_X2 port map( A1 => n5139, A2 => n5138, ZN => n18788);
   U22195 : NAND2_X2 port map( A1 => n38583, A2 => n18915, ZN => n23884);
   U22206 : OAI21_X2 port map( A1 => n38499, A2 => n17521, B => n36212, ZN => 
                           n38583);
   U22211 : NOR2_X1 port map( A1 => n21269, A2 => n33368, ZN => n38864);
   U22213 : INV_X2 port map( I => n12924, ZN => n33368);
   U22215 : XOR2_X1 port map( A1 => n8888, A2 => n35142, Z => n12924);
   U22218 : XOR2_X1 port map( A1 => n26483, A2 => n12683, Z => n38585);
   U22222 : INV_X2 port map( I => n38586, ZN => n12049);
   U22228 : XNOR2_X1 port map( A1 => n9768, A2 => n12039, ZN => n38586);
   U22229 : XOR2_X1 port map( A1 => n1065, A2 => n15617, Z => n29056);
   U22236 : NAND2_X2 port map( A1 => n13962, A2 => n13965, ZN => n15617);
   U22237 : XOR2_X1 port map( A1 => n22424, A2 => n22425, Z => n22943);
   U22238 : XOR2_X1 port map( A1 => n17838, A2 => n17839, Z => n11622);
   U22240 : OAI21_X2 port map( A1 => n31926, A2 => n31925, B => n38587, ZN => 
                           n7106);
   U22243 : XOR2_X1 port map( A1 => n38588, A2 => n19825, Z => Ciphertext(32));
   U22247 : AOI22_X1 port map( A1 => n13274, A2 => n15958, B1 => n13273, B2 => 
                           n13803, ZN => n38588);
   U22249 : NOR2_X2 port map( A1 => n38589, A2 => n29350, ZN => n9839);
   U22251 : OAI22_X2 port map( A1 => n4790, A2 => n5334, B1 => n5336, B2 => 
                           n1401, ZN => n38589);
   U22254 : XOR2_X1 port map( A1 => n28837, A2 => n11922, Z => n3081);
   U22256 : XOR2_X1 port map( A1 => n28925, A2 => n3082, Z => n28837);
   U22258 : XOR2_X1 port map( A1 => n29243, A2 => n38590, Z => n37034);
   U22260 : XOR2_X1 port map( A1 => n17243, A2 => n3665, Z => n38590);
   U22266 : NAND3_X1 port map( A1 => n1193, A2 => n5418, A3 => n31015, ZN => 
                           n10361);
   U22268 : INV_X2 port map( I => n10980, ZN => n38674);
   U22279 : XOR2_X1 port map( A1 => n25324, A2 => n37110, Z => n813);
   U22281 : NOR2_X1 port map( A1 => n36422, A2 => n14439, ZN => n22792);
   U22284 : NAND2_X1 port map( A1 => n38592, A2 => n38591, ZN => n18054);
   U22286 : NAND2_X2 port map( A1 => n39361, A2 => n34220, ZN => n10463);
   U22293 : NAND2_X2 port map( A1 => n38593, A2 => n19109, ZN => n29559);
   U22296 : NAND2_X1 port map( A1 => n34804, A2 => n34806, ZN => n38593);
   U22297 : OR2_X1 port map( A1 => n38358, A2 => n25660, Z => n25576);
   U22301 : NOR2_X1 port map( A1 => n24608, A2 => n39704, ZN => n7067);
   U22309 : NAND2_X2 port map( A1 => n3794, A2 => n38596, ZN => n11330);
   U22315 : INV_X1 port map( I => n34134, ZN => n39021);
   U22318 : XNOR2_X1 port map( A1 => n7076, A2 => n31289, ZN => n34134);
   U22319 : INV_X2 port map( I => n38597, ZN => n24404);
   U22321 : XOR2_X1 port map( A1 => n13568, A2 => n3447, Z => n3446);
   U22322 : XOR2_X1 port map( A1 => n26197, A2 => n26225, Z => n32839);
   U22323 : XOR2_X1 port map( A1 => n15034, A2 => n38598, Z => n15036);
   U22324 : XOR2_X1 port map( A1 => n24641, A2 => n37231, Z => n38598);
   U22325 : OAI21_X2 port map( A1 => n38599, A2 => n1940, B => n1939, ZN => 
                           n1938);
   U22347 : NOR2_X1 port map( A1 => n3690, A2 => n2502, ZN => n38599);
   U22348 : AND2_X1 port map( A1 => n22347, A2 => n22346, Z => n10037);
   U22351 : NAND2_X2 port map( A1 => n36753, A2 => n10630, ZN => n22347);
   U22353 : INV_X2 port map( I => n32601, ZN => n38600);
   U22354 : INV_X4 port map( I => n39663, ZN => n2416);
   U22366 : XOR2_X1 port map( A1 => n38602, A2 => n20257, Z => n26921);
   U22368 : XOR2_X1 port map( A1 => n20260, A2 => n32175, Z => n38602);
   U22371 : XOR2_X1 port map( A1 => n24039, A2 => n38603, Z => n2168);
   U22372 : XOR2_X1 port map( A1 => n36748, A2 => n36895, Z => n38603);
   U22373 : XOR2_X1 port map( A1 => n38988, A2 => n18491, Z => n18525);
   U22374 : OR2_X1 port map( A1 => n33483, A2 => n24192, Z => n15258);
   U22376 : XOR2_X1 port map( A1 => n15250, A2 => n7359, Z => n33483);
   U22381 : AOI22_X2 port map( A1 => n2520, A2 => n1890, B1 => n9201, B2 => 
                           n2519, ZN => n2518);
   U22383 : XOR2_X1 port map( A1 => n29158, A2 => n38606, Z => n38605);
   U22384 : NAND2_X2 port map( A1 => n28258, A2 => n27884, ZN => n28171);
   U22386 : XOR2_X1 port map( A1 => n27537, A2 => n34963, Z => n27805);
   U22391 : NOR2_X2 port map( A1 => n5769, A2 => n5770, ZN => n34963);
   U22393 : XOR2_X1 port map( A1 => n18785, A2 => n29104, Z => n28603);
   U22396 : NAND3_X2 port map( A1 => n28601, A2 => n34463, A3 => n34462, ZN => 
                           n29104);
   U22406 : NAND2_X2 port map( A1 => n27870, A2 => n19743, ZN => n27871);
   U22409 : NAND2_X2 port map( A1 => n14829, A2 => n14828, ZN => n33307);
   U22410 : AOI21_X2 port map( A1 => n21025, A2 => n16691, B => n38607, ZN => 
                           n21024);
   U22413 : NOR3_X2 port map( A1 => n36814, A2 => n31924, A3 => n28299, ZN => 
                           n38607);
   U22414 : NOR2_X2 port map( A1 => n8090, A2 => n38608, ZN => n11753);
   U22416 : INV_X2 port map( I => n26157, ZN => n26394);
   U22426 : XOR2_X1 port map( A1 => n38610, A2 => n39025, Z => n33387);
   U22428 : NAND2_X1 port map( A1 => n38408, A2 => n37088, ZN => n31739);
   U22431 : AOI22_X2 port map( A1 => n28513, A2 => n29702, B1 => n34793, B2 => 
                           n35858, ZN => n29568);
   U22435 : XOR2_X1 port map( A1 => n12865, A2 => n27480, Z => n11237);
   U22437 : NAND2_X2 port map( A1 => n5695, A2 => n16856, ZN => n12865);
   U22440 : NOR2_X2 port map( A1 => n38612, A2 => n556, ZN => n27498);
   U22442 : AOI21_X2 port map( A1 => n27205, A2 => n27206, B => n27400, ZN => 
                           n38612);
   U22443 : NAND2_X2 port map( A1 => n38615, A2 => n38613, ZN => n17745);
   U22447 : NAND2_X1 port map( A1 => n38614, A2 => n23550, ZN => n38613);
   U22448 : XOR2_X1 port map( A1 => n24013, A2 => n38616, Z => n39590);
   U22455 : XOR2_X1 port map( A1 => n24012, A2 => n35640, Z => n38616);
   U22457 : XOR2_X1 port map( A1 => n31565, A2 => n31863, Z => n11233);
   U22461 : NAND2_X2 port map( A1 => n8213, A2 => n8211, ZN => n24076);
   U22464 : AOI22_X2 port map( A1 => n33667, A2 => n23505, B1 => n8214, B2 => 
                           n8190, ZN => n8213);
   U22468 : INV_X2 port map( I => n21461, ZN => n38617);
   U22473 : NOR2_X2 port map( A1 => n38617, A2 => n21869, ZN => n32114);
   U22474 : NAND2_X2 port map( A1 => n56, A2 => n38621, ZN => n34609);
   U22476 : NAND3_X2 port map( A1 => n12704, A2 => n12705, A3 => n1115, ZN => 
                           n38621);
   U22478 : XOR2_X1 port map( A1 => n19632, A2 => n38622, Z => n26931);
   U22479 : XOR2_X1 port map( A1 => n26558, A2 => n26557, Z => n38622);
   U22481 : NOR2_X2 port map( A1 => n5311, A2 => n27407, ZN => n5059);
   U22486 : XOR2_X1 port map( A1 => n6066, A2 => n24959, Z => n25257);
   U22488 : NOR2_X2 port map( A1 => n38867, A2 => n30413, ZN => n24959);
   U22490 : XOR2_X1 port map( A1 => n23396, A2 => n37148, Z => n7734);
   U22492 : XOR2_X1 port map( A1 => n24023, A2 => n23764, Z => n23396);
   U22493 : NAND2_X2 port map( A1 => n34895, A2 => n11170, ZN => n24712);
   U22496 : AOI21_X2 port map( A1 => n1453, A2 => n2262, B => n12443, ZN => 
                           n4151);
   U22497 : XOR2_X1 port map( A1 => n29167, A2 => n6719, Z => n28909);
   U22501 : NOR2_X2 port map( A1 => n35823, A2 => n16036, ZN => n6719);
   U22502 : INV_X2 port map( I => n38627, ZN => n35792);
   U22503 : NAND3_X2 port map( A1 => n23160, A2 => n35684, A3 => n10436, ZN => 
                           n38627);
   U22505 : NAND2_X2 port map( A1 => n14794, A2 => n38628, ZN => n378);
   U22509 : XOR2_X1 port map( A1 => n27464, A2 => n27492, Z => n27847);
   U22511 : NOR2_X2 port map( A1 => n19803, A2 => n19802, ZN => n27464);
   U22513 : NAND2_X2 port map( A1 => n16535, A2 => n10209, ZN => n17996);
   U22516 : NAND2_X2 port map( A1 => n31425, A2 => n12556, ZN => n4529);
   U22523 : OR2_X1 port map( A1 => n6533, A2 => n36509, Z => n27237);
   U22524 : NAND2_X2 port map( A1 => n7800, A2 => n24240, ZN => n24243);
   U22527 : XOR2_X1 port map( A1 => n4086, A2 => n4085, Z => n8452);
   U22528 : AND2_X1 port map( A1 => n24898, A2 => n39505, Z => n5030);
   U22535 : AOI22_X2 port map( A1 => n10069, A2 => n20058, B1 => n14156, B2 => 
                           n6215, ZN => n6214);
   U22542 : OAI21_X2 port map( A1 => n33995, A2 => n38075, B => n3903, ZN => 
                           n6505);
   U22546 : NAND2_X1 port map( A1 => n3373, A2 => n19098, ZN => n3372);
   U22548 : OAI22_X2 port map( A1 => n1079, A2 => n38638, B1 => n8453, B2 => 
                           n10946, ZN => n15465);
   U22550 : XOR2_X1 port map( A1 => n12971, A2 => n33334, Z => n38639);
   U22563 : AOI22_X2 port map( A1 => n22138, A2 => n22246, B1 => n22139, B2 => 
                           n35290, ZN => n38640);
   U22565 : NAND2_X1 port map( A1 => n19514, A2 => n25420, ZN => n38642);
   U22567 : NAND2_X1 port map( A1 => n38644, A2 => n34005, ZN => n38643);
   U22569 : INV_X2 port map( I => n19821, ZN => n38644);
   U22570 : NAND2_X2 port map( A1 => n34683, A2 => n38645, ZN => n22228);
   U22573 : AOI21_X2 port map( A1 => n38647, A2 => n1351, B => n38646, ZN => 
                           n38645);
   U22574 : NOR2_X1 port map( A1 => n17160, A2 => n1351, ZN => n38646);
   U22575 : INV_X1 port map( I => n13348, ZN => n38647);
   U22579 : XOR2_X1 port map( A1 => n31352, A2 => n22605, Z => n2030);
   U22587 : XOR2_X1 port map( A1 => n38648, A2 => n11755, Z => n36880);
   U22588 : NAND2_X2 port map( A1 => n38780, A2 => n10949, ZN => n11755);
   U22602 : XOR2_X1 port map( A1 => n38649, A2 => n20674, Z => n20677);
   U22603 : XOR2_X1 port map( A1 => n21157, A2 => n10258, Z => n38649);
   U22604 : NOR2_X2 port map( A1 => n38650, A2 => n15969, ZN => n23929);
   U22612 : INV_X2 port map( I => n33786, ZN => n39300);
   U22613 : NAND2_X2 port map( A1 => n13406, A2 => n13407, ZN => n33786);
   U22615 : XOR2_X1 port map( A1 => n1557, A2 => n25079, Z => n25148);
   U22617 : NAND2_X1 port map( A1 => n23342, A2 => n23343, ZN => n23344);
   U22620 : NAND2_X2 port map( A1 => n33894, A2 => n23624, ZN => n23342);
   U22621 : XOR2_X1 port map( A1 => n23982, A2 => n5290, Z => n36079);
   U22622 : OR2_X1 port map( A1 => n39265, A2 => n24868, Z => n32268);
   U22623 : NAND2_X2 port map( A1 => n4452, A2 => n4453, ZN => n26098);
   U22624 : NAND2_X2 port map( A1 => n20642, A2 => n28297, ZN => n16096);
   U22630 : NAND3_X2 port map( A1 => n20111, A2 => n27317, A3 => n27316, ZN => 
                           n7549);
   U22634 : OAI21_X2 port map( A1 => n8993, A2 => n38868, B => n37828, ZN => 
                           n32146);
   U22635 : XOR2_X1 port map( A1 => n38654, A2 => n11210, Z => n34218);
   U22642 : XOR2_X1 port map( A1 => n27841, A2 => n27740, Z => n38654);
   U22644 : AOI22_X2 port map( A1 => n6314, A2 => n29453, B1 => n39647, B2 => 
                           n29378, ZN => n39060);
   U22648 : XOR2_X1 port map( A1 => n18930, A2 => n18705, Z => n19478);
   U22661 : INV_X1 port map( I => n38843, ZN => n17894);
   U22665 : OR2_X1 port map( A1 => n38843, A2 => n34010, Z => n17038);
   U22666 : XOR2_X1 port map( A1 => n3320, A2 => n38655, Z => n3885);
   U22671 : XOR2_X1 port map( A1 => n33310, A2 => n38261, Z => n38655);
   U22672 : NAND2_X2 port map( A1 => n3964, A2 => n3966, ZN => n29085);
   U22676 : NAND2_X2 port map( A1 => n988, A2 => n10642, ZN => n28276);
   U22677 : AOI21_X2 port map( A1 => n14543, A2 => n28808, B => n38657, ZN => 
                           n16658);
   U22680 : XOR2_X1 port map( A1 => n12401, A2 => n12400, Z => n12399);
   U22683 : NOR2_X2 port map( A1 => n27371, A2 => n31672, ZN => n12374);
   U22685 : NAND2_X2 port map( A1 => n27372, A2 => n27267, ZN => n27371);
   U22690 : XOR2_X1 port map( A1 => n24938, A2 => n25176, Z => n25246);
   U22694 : NOR2_X2 port map( A1 => n24815, A2 => n7321, ZN => n25176);
   U22695 : XOR2_X1 port map( A1 => n5731, A2 => n36339, Z => n30465);
   U22698 : NAND2_X1 port map( A1 => n39013, A2 => n36560, ZN => n39131);
   U22700 : XOR2_X1 port map( A1 => n10782, A2 => n27793, Z => n8958);
   U22702 : XOR2_X1 port map( A1 => n3163, A2 => n4734, Z => n38659);
   U22704 : XOR2_X1 port map( A1 => n28855, A2 => n28545, Z => n12455);
   U22707 : XOR2_X1 port map( A1 => n29067, A2 => n29819, Z => n28855);
   U22709 : NAND2_X2 port map( A1 => n10807, A2 => n37172, ZN => n25827);
   U22710 : INV_X2 port map( I => n3496, ZN => n33894);
   U22715 : NAND3_X2 port map( A1 => n32909, A2 => n10437, A3 => n10438, ZN => 
                           n3496);
   U22719 : XOR2_X1 port map( A1 => n38660, A2 => n2159, Z => n31107);
   U22720 : XOR2_X1 port map( A1 => n3559, A2 => n27791, Z => n38660);
   U22721 : XOR2_X1 port map( A1 => n4412, A2 => n33039, Z => n4409);
   U22722 : NAND2_X1 port map( A1 => n23272, A2 => n18199, ZN => n18198);
   U22726 : OR2_X1 port map( A1 => n29199, A2 => n11348, Z => n35869);
   U22727 : AOI22_X2 port map( A1 => n25538, A2 => n13461, B1 => n39327, B2 => 
                           n12908, ZN => n38663);
   U22731 : XOR2_X1 port map( A1 => n38664, A2 => n18270, Z => Ciphertext(16));
   U22733 : NAND4_X2 port map( A1 => n29233, A2 => n36232, A3 => n39306, A4 => 
                           n29234, ZN => n38664);
   U22738 : XOR2_X1 port map( A1 => n37129, A2 => n7549, Z => n27817);
   U22742 : NOR2_X2 port map( A1 => n14614, A2 => n6648, ZN => n20112);
   U22748 : NOR2_X2 port map( A1 => n32131, A2 => n7706, ZN => n14614);
   U22749 : NAND3_X1 port map( A1 => n5282, A2 => n24683, A3 => n13300, ZN => 
                           n17893);
   U22755 : NAND2_X2 port map( A1 => n8925, A2 => n33493, ZN => n5282);
   U22756 : NAND3_X1 port map( A1 => n20174, A2 => n20590, A3 => n19966, ZN => 
                           n2356);
   U22757 : OR2_X1 port map( A1 => n6515, A2 => n33599, Z => n35150);
   U22758 : OAI21_X2 port map( A1 => n38667, A2 => n34524, B => n1020, ZN => 
                           n3380);
   U22759 : NOR2_X2 port map( A1 => n1104, A2 => n26055, ZN => n38667);
   U22762 : XOR2_X1 port map( A1 => n22509, A2 => n22510, Z => n22661);
   U22766 : NAND3_X2 port map( A1 => n24121, A2 => n17066, A3 => n35253, ZN => 
                           n34693);
   U22770 : XOR2_X1 port map( A1 => n6277, A2 => n38670, Z => n24196);
   U22772 : XOR2_X1 port map( A1 => n23711, A2 => n23865, Z => n38670);
   U22774 : XOR2_X1 port map( A1 => n9577, A2 => n7371, Z => n26808);
   U22778 : XOR2_X1 port map( A1 => n27613, A2 => n27614, Z => n28157);
   U22780 : NAND2_X2 port map( A1 => n24345, A2 => n5953, ZN => n39413);
   U22786 : XOR2_X1 port map( A1 => n26435, A2 => n26387, Z => n26527);
   U22788 : NOR2_X2 port map( A1 => n16525, A2 => n25821, ZN => n26435);
   U22790 : AOI22_X2 port map( A1 => n23297, A2 => n23462, B1 => n23298, B2 => 
                           n23460, ZN => n23301);
   U22801 : NAND2_X1 port map( A1 => n38727, A2 => n28546, ZN => n19043);
   U22802 : AOI21_X2 port map( A1 => n9375, A2 => n9380, B => n38671, ZN => 
                           n31883);
   U22805 : INV_X2 port map( I => n25532, ZN => n38671);
   U22809 : NAND2_X2 port map( A1 => n15085, A2 => n33440, ZN => n25532);
   U22812 : XOR2_X1 port map( A1 => n4081, A2 => n39119, Z => n26651);
   U22815 : OAI22_X2 port map( A1 => n4455, A2 => n4454, B1 => n32722, B2 => 
                           n25514, ZN => n4453);
   U22816 : AOI22_X2 port map( A1 => n30397, A2 => n21900, B1 => n21901, B2 => 
                           n275, ZN => n15468);
   U22817 : NOR2_X2 port map( A1 => n21840, A2 => n1348, ZN => n21901);
   U22818 : BUF_X2 port map( I => n36371, Z => n38673);
   U22820 : NAND2_X1 port map( A1 => n29208, A2 => n15535, ZN => n29205);
   U22828 : AOI21_X2 port map( A1 => n38676, A2 => n23100, B => n11659, ZN => 
                           n13087);
   U22830 : NOR2_X2 port map( A1 => n15330, A2 => n33082, ZN => n38676);
   U22835 : NAND2_X2 port map( A1 => n38677, A2 => n11260, ZN => n24817);
   U22844 : NAND2_X1 port map( A1 => n10219, A2 => n36872, ZN => n38677);
   U22848 : XOR2_X1 port map( A1 => n29088, A2 => n2392, Z => n10185);
   U22849 : AND2_X1 port map( A1 => n18827, A2 => n35648, Z => n39806);
   U22853 : NAND3_X2 port map( A1 => n5864, A2 => n5863, A3 => n38678, ZN => 
                           n7023);
   U22857 : XOR2_X1 port map( A1 => n14039, A2 => n38679, Z => n30925);
   U22868 : NAND2_X2 port map( A1 => n12046, A2 => n12045, ZN => n14039);
   U22869 : AOI22_X2 port map( A1 => n27344, A2 => n1225, B1 => n27342, B2 => 
                           n27343, ZN => n27345);
   U22878 : OAI21_X2 port map( A1 => n1029, A2 => n9825, B => n17101, ZN => 
                           n10654);
   U22880 : NAND2_X2 port map( A1 => n24108, A2 => n24109, ZN => n9825);
   U22884 : CLKBUF_X4 port map( I => n966, Z => n39018);
   U22890 : OR2_X2 port map( A1 => n2416, A2 => n39021, Z => n36345);
   U22896 : NAND2_X2 port map( A1 => n9835, A2 => n23475, ZN => n19633);
   U22900 : NAND2_X1 port map( A1 => n38223, A2 => n3937, ZN => n9337);
   U22908 : XOR2_X1 port map( A1 => n28967, A2 => n10328, Z => n36746);
   U22911 : XOR2_X1 port map( A1 => n26531, A2 => n32253, Z => n12411);
   U22919 : OAI21_X2 port map( A1 => n3244, A2 => n7699, B => n39625, ZN => 
                           n26531);
   U22920 : XOR2_X1 port map( A1 => n36804, A2 => n38680, Z => n12298);
   U22930 : XOR2_X1 port map( A1 => n9184, A2 => n6688, Z => n38680);
   U22934 : XOR2_X1 port map( A1 => n18327, A2 => n38682, Z => n39263);
   U22945 : XOR2_X1 port map( A1 => n24702, A2 => n37121, Z => n38682);
   U22954 : NAND2_X1 port map( A1 => n38644, A2 => n11616, ZN => n38683);
   U22956 : NAND2_X1 port map( A1 => n1235, A2 => n38684, ZN => n32725);
   U22957 : NAND2_X2 port map( A1 => n12392, A2 => n23111, ZN => n3119);
   U22959 : AOI21_X2 port map( A1 => n38686, A2 => n38685, B => n1115, ZN => 
                           n34272);
   U22963 : INV_X2 port map( I => n34010, ZN => n38685);
   U22971 : BUF_X2 port map( I => n35431, Z => n38687);
   U22972 : NAND2_X2 port map( A1 => n38689, A2 => n38688, ZN => n26648);
   U22973 : XOR2_X1 port map( A1 => n26262, A2 => n35212, Z => n844);
   U22976 : OAI21_X2 port map( A1 => n16239, A2 => n7888, B => n25807, ZN => 
                           n26262);
   U22977 : OAI21_X2 port map( A1 => n16182, A2 => n6176, B => n38691, ZN => 
                           n15353);
   U22983 : NAND2_X2 port map( A1 => n4160, A2 => n4161, ZN => n6176);
   U22984 : NAND2_X2 port map( A1 => n13233, A2 => n10346, ZN => n29630);
   U22985 : XOR2_X1 port map( A1 => n9894, A2 => n38692, Z => n2052);
   U22986 : XOR2_X1 port map( A1 => n11938, A2 => n36067, Z => n38692);
   U22992 : AND2_X1 port map( A1 => n36509, A2 => n36523, Z => n32950);
   U22994 : INV_X2 port map( I => n18175, ZN => n23757);
   U23000 : NAND2_X2 port map( A1 => n38693, A2 => n36091, ZN => n18175);
   U23009 : OR2_X1 port map( A1 => n20818, A2 => n18389, Z => n38693);
   U23014 : XOR2_X1 port map( A1 => n17360, A2 => n17361, Z => n36970);
   U23015 : NOR2_X2 port map( A1 => n8641, A2 => n8640, ZN => n39442);
   U23022 : NOR2_X2 port map( A1 => n13308, A2 => n24301, ZN => n38749);
   U23028 : AOI21_X2 port map( A1 => n29781, A2 => n1402, B => n481, ZN => 
                           n2017);
   U23029 : NAND3_X1 port map( A1 => n23518, A2 => n39001, A3 => n6373, ZN => 
                           n38806);
   U23031 : AOI22_X2 port map( A1 => n38800, A2 => n35288, B1 => n17778, B2 => 
                           n7902, ZN => n39001);
   U23035 : OR2_X1 port map( A1 => n20566, A2 => n29241, Z => n38823);
   U23037 : AOI22_X2 port map( A1 => n35369, A2 => n1186, B1 => n20621, B2 => 
                           n7486, ZN => n20314);
   U23038 : BUF_X2 port map( I => n6056, Z => n38694);
   U23039 : AND2_X1 port map( A1 => n37188, A2 => n6136, Z => n39530);
   U23044 : NAND2_X2 port map( A1 => n6390, A2 => n6180, ZN => n7961);
   U23045 : INV_X2 port map( I => n27314, ZN => n27409);
   U23046 : OAI22_X2 port map( A1 => n12714, A2 => n12713, B1 => n26766, B2 => 
                           n12078, ZN => n27314);
   U23048 : NAND2_X2 port map( A1 => n8253, A2 => n32191, ZN => n27084);
   U23050 : NAND2_X2 port map( A1 => n33098, A2 => n33097, ZN => n8253);
   U23059 : AOI21_X2 port map( A1 => n24155, A2 => n10220, B => n2595, ZN => 
                           n38695);
   U23060 : NAND2_X1 port map( A1 => n25486, A2 => n18207, ZN => n25305);
   U23062 : AOI22_X2 port map( A1 => n38696, A2 => n24655, B1 => n24507, B2 => 
                           n33409, ZN => n4729);
   U23065 : NOR2_X2 port map( A1 => n19679, A2 => n37355, ZN => n38696);
   U23066 : AND2_X1 port map( A1 => n5383, A2 => n39435, Z => n39473);
   U23081 : XOR2_X1 port map( A1 => n38697, A2 => n19805, Z => Ciphertext(76));
   U23085 : NAND2_X2 port map( A1 => n38698, A2 => n35762, ZN => n29616);
   U23089 : XOR2_X1 port map( A1 => n22659, A2 => n19128, Z => n19127);
   U23094 : XNOR2_X1 port map( A1 => n22702, A2 => n644, ZN => n39039);
   U23109 : NAND3_X1 port map( A1 => n9987, A2 => n5819, A3 => n21961, ZN => 
                           n38699);
   U23111 : XOR2_X1 port map( A1 => n31492, A2 => n39654, Z => n11810);
   U23113 : NOR2_X1 port map( A1 => n38701, A2 => n38700, ZN => n39007);
   U23116 : INV_X1 port map( I => n5819, ZN => n38701);
   U23122 : INV_X2 port map( I => n19142, ZN => n38702);
   U23130 : NAND2_X2 port map( A1 => n15811, A2 => n15814, ZN => n17499);
   U23132 : INV_X1 port map( I => n5340, ZN => n8703);
   U23134 : NOR2_X2 port map( A1 => n12784, A2 => n28282, ZN => n28167);
   U23138 : OR2_X1 port map( A1 => n14212, A2 => n10986, Z => n12552);
   U23141 : XOR2_X1 port map( A1 => n27785, A2 => n20721, Z => n32807);
   U23144 : OAI21_X1 port map( A1 => n27282, A2 => n1227, B => n38705, ZN => 
                           n3718);
   U23145 : NAND2_X1 port map( A1 => n27282, A2 => n3313, ZN => n38705);
   U23148 : XOR2_X1 port map( A1 => n3731, A2 => n18887, Z => n38706);
   U23153 : XOR2_X1 port map( A1 => n311, A2 => n10014, Z => n11586);
   U23155 : NAND2_X2 port map( A1 => n32883, A2 => n2182, ZN => n9968);
   U23158 : NAND2_X2 port map( A1 => n38708, A2 => n38707, ZN => n29189);
   U23165 : NAND2_X2 port map( A1 => n29187, A2 => n3631, ZN => n38707);
   U23181 : NAND2_X2 port map( A1 => n29188, A2 => n38709, ZN => n38708);
   U23182 : NOR2_X1 port map( A1 => n24091, A2 => n37066, ZN => n39191);
   U23184 : XOR2_X1 port map( A1 => n38820, A2 => n29816, Z => n38710);
   U23187 : INV_X4 port map( I => n7445, ZN => n24646);
   U23189 : NAND2_X2 port map( A1 => n28087, A2 => n28086, ZN => n33047);
   U23193 : XOR2_X1 port map( A1 => n24997, A2 => n2653, Z => n25210);
   U23201 : NAND2_X2 port map( A1 => n16668, A2 => n14681, ZN => n24997);
   U23204 : NAND2_X2 port map( A1 => n15670, A2 => n26944, ZN => n38715);
   U23205 : NAND2_X1 port map( A1 => n19367, A2 => n12162, ZN => n38716);
   U23209 : OAI21_X2 port map( A1 => n36295, A2 => n13516, B => n24616, ZN => 
                           n34564);
   U23210 : OAI21_X2 port map( A1 => n2331, A2 => n14278, B => n38717, ZN => 
                           n16017);
   U23212 : OAI22_X2 port map( A1 => n22246, A2 => n38718, B1 => n35290, B2 => 
                           n9265, ZN => n22036);
   U23213 : INV_X2 port map( I => n33713, ZN => n38719);
   U23215 : NAND2_X2 port map( A1 => n38721, A2 => n38720, ZN => n23778);
   U23226 : NAND2_X1 port map( A1 => n19633, A2 => n12011, ZN => n38720);
   U23227 : OAI21_X2 port map( A1 => n12008, A2 => n12009, B => n34823, ZN => 
                           n38721);
   U23231 : XOR2_X1 port map( A1 => n29093, A2 => n1411, Z => n28984);
   U23234 : INV_X2 port map( I => n31396, ZN => n1411);
   U23237 : NOR2_X2 port map( A1 => n34266, A2 => n18103, ZN => n31396);
   U23239 : OAI21_X2 port map( A1 => n2062, A2 => n17075, B => n38722, ZN => 
                           n39030);
   U23240 : AOI22_X2 port map( A1 => n33113, A2 => n33115, B1 => n1984, B2 => 
                           n33114, ZN => n38722);
   U23249 : XOR2_X1 port map( A1 => n38723, A2 => n16975, Z => n29768);
   U23253 : XOR2_X1 port map( A1 => n20006, A2 => n489, Z => n38723);
   U23256 : BUF_X2 port map( I => n34757, Z => n38725);
   U23259 : INV_X4 port map( I => n24896, ZN => n38782);
   U23269 : OR2_X1 port map( A1 => n23489, A2 => n23602, Z => n30631);
   U23270 : NOR2_X1 port map( A1 => n5598, A2 => n21914, ZN => n20832);
   U23272 : AND2_X1 port map( A1 => n33316, A2 => n23444, Z => n38893);
   U23276 : NAND2_X2 port map( A1 => n38729, A2 => n38728, ZN => n30372);
   U23277 : NAND2_X2 port map( A1 => n38731, A2 => n38730, ZN => n38729);
   U23285 : INV_X2 port map( I => n25542, ZN => n38731);
   U23286 : BUF_X2 port map( I => n39820, Z => n38732);
   U23289 : NAND3_X2 port map( A1 => n38733, A2 => n36098, A3 => n36097, ZN => 
                           n9310);
   U23301 : OAI21_X2 port map( A1 => n37156, A2 => n7511, B => n26564, ZN => 
                           n38733);
   U23303 : XOR2_X1 port map( A1 => n12534, A2 => n19359, Z => n25152);
   U23309 : NAND3_X2 port map( A1 => n5123, A2 => n5122, A3 => n31455, ZN => 
                           n12534);
   U23311 : XOR2_X1 port map( A1 => n38735, A2 => n26584, Z => n11374);
   U23312 : XOR2_X1 port map( A1 => n26365, A2 => n12667, Z => n38735);
   U23314 : OAI21_X2 port map( A1 => n20584, A2 => n31966, B => n11518, ZN => 
                           n14448);
   U23315 : NAND2_X2 port map( A1 => n10469, A2 => n10471, ZN => n11970);
   U23316 : OAI21_X2 port map( A1 => n34618, A2 => n34619, B => n9872, ZN => 
                           n38737);
   U23319 : XOR2_X1 port map( A1 => n35089, A2 => n36211, Z => n34876);
   U23320 : INV_X1 port map( I => n38739, ZN => n8210);
   U23322 : OAI21_X2 port map( A1 => n31234, A2 => n31235, B => n30274, ZN => 
                           n13306);
   U23323 : NAND2_X2 port map( A1 => n18330, A2 => n18331, ZN => n11342);
   U23326 : OAI21_X2 port map( A1 => n26220, A2 => n1494, B => n38740, ZN => 
                           n6376);
   U23327 : NOR2_X2 port map( A1 => n34224, A2 => n37103, ZN => n38740);
   U23328 : XOR2_X1 port map( A1 => n27475, A2 => n38741, Z => n34491);
   U23335 : INV_X2 port map( I => n8874, ZN => n38741);
   U23340 : XOR2_X1 port map( A1 => n26278, A2 => n35214, Z => n11399);
   U23341 : NAND3_X2 port map( A1 => n13184, A2 => n13182, A3 => n36801, ZN => 
                           n20576);
   U23343 : INV_X2 port map( I => n38743, ZN => n17390);
   U23347 : NOR2_X2 port map( A1 => n38745, A2 => n38744, ZN => n36408);
   U23357 : NOR2_X2 port map( A1 => n10654, A2 => n2341, ZN => n38745);
   U23366 : BUF_X2 port map( I => n20391, Z => n38746);
   U23368 : NOR2_X2 port map( A1 => n33036, A2 => n38747, ZN => n12393);
   U23376 : NAND2_X2 port map( A1 => n20405, A2 => n34389, ZN => n6045);
   U23377 : BUF_X2 port map( I => n23550, Z => n38748);
   U23378 : NOR2_X2 port map( A1 => n31601, A2 => n30097, ZN => n30087);
   U23381 : AOI21_X2 port map( A1 => n3527, A2 => n19476, B => n6044, ZN => 
                           n31601);
   U23383 : XOR2_X1 port map( A1 => n38750, A2 => n15331, Z => n4016);
   U23386 : XOR2_X1 port map( A1 => n3386, A2 => n20719, Z => n38750);
   U23387 : XOR2_X1 port map( A1 => n5603, A2 => n39028, Z => n34757);
   U23395 : INV_X2 port map( I => n38751, ZN => n1984);
   U23397 : NAND2_X2 port map( A1 => n2416, A2 => n37086, ZN => n38751);
   U23398 : NAND2_X2 port map( A1 => n34326, A2 => n20084, ZN => n29071);
   U23399 : OR2_X1 port map( A1 => n1448, A2 => n28079, Z => n7219);
   U23408 : OAI21_X2 port map( A1 => n19006, A2 => n38754, B => n23259, ZN => 
                           n23910);
   U23411 : XOR2_X1 port map( A1 => n25186, A2 => n25118, Z => n11102);
   U23414 : NAND2_X2 port map( A1 => n819, A2 => n24210, ZN => n25118);
   U23419 : NAND2_X2 port map( A1 => n21662, A2 => n21951, ZN => n20367);
   U23421 : NAND2_X2 port map( A1 => n32113, A2 => n17991, ZN => n17989);
   U23423 : AOI21_X2 port map( A1 => n23201, A2 => n38756, B => n22850, ZN => 
                           n2413);
   U23425 : NOR2_X1 port map( A1 => n2350, A2 => n36369, ZN => n38756);
   U23426 : XOR2_X1 port map( A1 => n4354, A2 => n4355, Z => n4356);
   U23427 : INV_X1 port map( I => n33883, ZN => n27727);
   U23437 : XNOR2_X1 port map( A1 => n27683, A2 => n27858, ZN => n33883);
   U23439 : XOR2_X1 port map( A1 => n38758, A2 => n34933, Z => n18790);
   U23443 : XOR2_X1 port map( A1 => n23549, A2 => n21045, Z => n38758);
   U23445 : XOR2_X1 port map( A1 => n23979, A2 => n23715, Z => n23563);
   U23446 : XOR2_X1 port map( A1 => n7498, A2 => n9911, Z => n12631);
   U23447 : XOR2_X1 port map( A1 => n11600, A2 => n20268, Z => n20704);
   U23448 : XOR2_X1 port map( A1 => n38759, A2 => n28787, Z => n20453);
   U23449 : XOR2_X1 port map( A1 => n2431, A2 => n29128, Z => n38759);
   U23450 : XOR2_X1 port map( A1 => n22561, A2 => n3528, Z => n22758);
   U23451 : NOR2_X2 port map( A1 => n637, A2 => n12155, ZN => n22561);
   U23461 : OR2_X1 port map( A1 => n29737, A2 => n19348, Z => n19369);
   U23463 : NAND2_X2 port map( A1 => n16057, A2 => n16056, ZN => n24023);
   U23467 : XOR2_X1 port map( A1 => n23786, A2 => n15777, Z => n20602);
   U23469 : XOR2_X1 port map( A1 => n11098, A2 => n23880, Z => n15777);
   U23471 : OAI21_X2 port map( A1 => n20863, A2 => n38302, B => n14699, ZN => 
                           n13351);
   U23473 : NAND3_X2 port map( A1 => n31331, A2 => n31332, A3 => n15953, ZN => 
                           n14365);
   U23474 : NAND2_X2 port map( A1 => n39255, A2 => n38761, ZN => n8163);
   U23477 : AOI22_X2 port map( A1 => n24771, A2 => n24770, B1 => n24769, B2 => 
                           n11846, ZN => n38761);
   U23478 : XOR2_X1 port map( A1 => n38763, A2 => n6324, Z => n39043);
   U23481 : OAI21_X2 port map( A1 => n38765, A2 => n38764, B => n27911, ZN => 
                           n18480);
   U23486 : NAND2_X1 port map( A1 => n22316, A2 => n3863, ZN => n22270);
   U23487 : NAND2_X2 port map( A1 => n2403, A2 => n5417, ZN => n22316);
   U23488 : NAND2_X2 port map( A1 => n32727, A2 => n32728, ZN => n38766);
   U23494 : NAND2_X2 port map( A1 => n37014, A2 => n23456, ZN => n17995);
   U23497 : NAND2_X2 port map( A1 => n18819, A2 => n32397, ZN => n37014);
   U23499 : NOR2_X2 port map( A1 => n24336, A2 => n24232, ZN => n12250);
   U23501 : INV_X4 port map( I => n38768, ZN => n22222);
   U23505 : OR2_X2 port map( A1 => n33051, A2 => n21679, Z => n38768);
   U23508 : NAND2_X2 port map( A1 => n38769, A2 => n8058, ZN => n23337);
   U23512 : NAND2_X2 port map( A1 => n22705, A2 => n22926, ZN => n38769);
   U23513 : NOR2_X2 port map( A1 => n37106, A2 => n6822, ZN => n34303);
   U23514 : XOR2_X1 port map( A1 => n38770, A2 => n3571, Z => n23827);
   U23517 : AOI22_X2 port map( A1 => n23496, A2 => n5357, B1 => n23592, B2 => 
                           n34603, ZN => n23594);
   U23522 : NAND2_X2 port map( A1 => n29426, A2 => n29424, ZN => n6314);
   U23523 : NAND2_X1 port map( A1 => n5500, A2 => n38771, ZN => n39775);
   U23524 : NAND2_X1 port map( A1 => n7992, A2 => n4736, ZN => n38771);
   U23529 : AND2_X1 port map( A1 => n11831, A2 => n28484, Z => n3019);
   U23535 : AOI22_X2 port map( A1 => n34112, A2 => n14081, B1 => n18058, B2 => 
                           n25502, ZN => n35453);
   U23538 : INV_X2 port map( I => n38772, ZN => n3488);
   U23539 : OR2_X2 port map( A1 => n1454, A2 => n18689, Z => n28175);
   U23548 : XOR2_X1 port map( A1 => n3320, A2 => n6365, Z => n32293);
   U23550 : NAND2_X2 port map( A1 => n27392, A2 => n35895, ZN => n27393);
   U23555 : AOI21_X2 port map( A1 => n38773, A2 => n14435, B => n12954, ZN => 
                           n15535);
   U23559 : NAND2_X2 port map( A1 => n27661, A2 => n27557, ZN => n10801);
   U23561 : NAND3_X2 port map( A1 => n36250, A2 => n27431, A3 => n10755, ZN => 
                           n27661);
   U23562 : NAND2_X2 port map( A1 => n7619, A2 => n6615, ZN => n38776);
   U23575 : INV_X2 port map( I => n39268, ZN => n38777);
   U23576 : NAND2_X2 port map( A1 => n36521, A2 => n36520, ZN => n7096);
   U23590 : NAND3_X2 port map( A1 => n20217, A2 => n26817, A3 => n26626, ZN => 
                           n27095);
   U23592 : OAI21_X2 port map( A1 => n38811, A2 => n36821, B => n38848, ZN => 
                           n31797);
   U23595 : XOR2_X1 port map( A1 => n6825, A2 => n18428, Z => n32734);
   U23599 : XOR2_X1 port map( A1 => n25104, A2 => n17184, Z => n18428);
   U23602 : NAND2_X2 port map( A1 => n38778, A2 => n30726, ZN => n12485);
   U23603 : OR2_X1 port map( A1 => n25412, A2 => n25307, Z => n38779);
   U23620 : NOR2_X2 port map( A1 => n28643, A2 => n14448, ZN => n28732);
   U23621 : NAND2_X1 port map( A1 => n34111, A2 => n31185, ZN => n38780);
   U23628 : NOR2_X2 port map( A1 => n23119, A2 => n1145, ZN => n23120);
   U23632 : NAND2_X1 port map( A1 => n5570, A2 => n921, ZN => n38785);
   U23641 : XOR2_X1 port map( A1 => n18180, A2 => n26438, Z => n26155);
   U23647 : NAND2_X2 port map( A1 => n38786, A2 => n6105, ZN => n36579);
   U23648 : OAI21_X2 port map( A1 => n7293, A2 => n2625, B => n7292, ZN => 
                           n38786);
   U23653 : INV_X2 port map( I => n27102, ZN => n38787);
   U23654 : NAND2_X2 port map( A1 => n19030, A2 => n38787, ZN => n27038);
   U23655 : AOI21_X1 port map( A1 => n5471, A2 => n18816, B => n39110, ZN => 
                           n4449);
   U23656 : XOR2_X1 port map( A1 => n2527, A2 => n2524, Z => n5717);
   U23658 : INV_X2 port map( I => n9020, ZN => n24136);
   U23662 : INV_X2 port map( I => n19233, ZN => n38886);
   U23665 : XOR2_X1 port map( A1 => n36760, A2 => n36759, Z => n19233);
   U23666 : OAI21_X2 port map( A1 => n944, A2 => n27269, B => n38788, ZN => 
                           n27374);
   U23667 : OAI21_X2 port map( A1 => n36224, A2 => n28281, B => n15622, ZN => 
                           n38854);
   U23669 : XOR2_X1 port map( A1 => n26413, A2 => n26412, Z => n7374);
   U23670 : XOR2_X1 port map( A1 => n26290, A2 => n39662, Z => n26413);
   U23671 : NAND2_X2 port map( A1 => n20988, A2 => n34693, ZN => n24812);
   U23675 : XOR2_X1 port map( A1 => n10706, A2 => n5486, Z => n38791);
   U23681 : AOI22_X2 port map( A1 => n34822, A2 => n22288, B1 => n22286, B2 => 
                           n22287, ZN => n9486);
   U23685 : XOR2_X1 port map( A1 => n21108, A2 => n28775, Z => n19047);
   U23686 : NOR2_X2 port map( A1 => n17849, A2 => n35272, ZN => n19157);
   U23690 : NAND2_X2 port map( A1 => n29401, A2 => n29402, ZN => n35272);
   U23692 : NAND2_X2 port map( A1 => n27298, A2 => n7757, ZN => n27070);
   U23696 : XOR2_X1 port map( A1 => n7737, A2 => n17579, Z => n31633);
   U23703 : XOR2_X1 port map( A1 => n27841, A2 => n38793, Z => n9039);
   U23704 : XOR2_X1 port map( A1 => n33398, A2 => n31620, Z => n38793);
   U23708 : OAI22_X2 port map( A1 => n38795, A2 => n38794, B1 => n18115, B2 => 
                           n1118, ZN => n15525);
   U23709 : OAI21_X1 port map( A1 => n9016, A2 => n10712, B => n36595, ZN => 
                           n3083);
   U23710 : XOR2_X1 port map( A1 => n26450, A2 => n31154, Z => n38796);
   U23714 : INV_X2 port map( I => n19425, ZN => n38797);
   U23715 : XOR2_X1 port map( A1 => n35241, A2 => n11755, Z => n27636);
   U23723 : OR2_X1 port map( A1 => n12334, A2 => n13082, Z => n28074);
   U23726 : INV_X1 port map( I => n15019, ZN => n21949);
   U23727 : NAND2_X2 port map( A1 => n2555, A2 => n2554, ZN => n29612);
   U23735 : NOR3_X2 port map( A1 => n38238, A2 => n38798, A3 => n34061, ZN => 
                           n32444);
   U23743 : XOR2_X1 port map( A1 => n16096, A2 => n38799, Z => n7766);
   U23744 : NOR2_X1 port map( A1 => n14408, A2 => n30942, ZN => n15142);
   U23747 : NAND2_X2 port map( A1 => n14408, A2 => n1006, ZN => n26661);
   U23749 : XOR2_X1 port map( A1 => n3474, A2 => n3471, Z => n17378);
   U23753 : INV_X2 port map( I => n38801, ZN => n34123);
   U23757 : OAI22_X2 port map( A1 => n9331, A2 => n23608, B1 => n32246, B2 => 
                           n98, ZN => n24030);
   U23758 : XOR2_X1 port map( A1 => n38802, A2 => n29506, Z => Ciphertext(54));
   U23771 : INV_X4 port map( I => n9333, ZN => n9733);
   U23772 : NAND2_X2 port map( A1 => n38803, A2 => n16231, ZN => n9970);
   U23773 : OAI21_X2 port map( A1 => n16016, A2 => n5980, B => n5979, ZN => 
                           n38803);
   U23775 : NOR2_X2 port map( A1 => n38807, A2 => n46, ZN => n10015);
   U23779 : AOI21_X2 port map( A1 => n11363, A2 => n16825, B => n38728, ZN => 
                           n38807);
   U23780 : XOR2_X1 port map( A1 => n28763, A2 => n36545, Z => n21162);
   U23785 : NAND3_X1 port map( A1 => n39206, A2 => n5311, A3 => n7606, ZN => 
                           n16517);
   U23788 : XOR2_X1 port map( A1 => n38808, A2 => n36284, Z => n39608);
   U23789 : XOR2_X1 port map( A1 => n39685, A2 => n37236, Z => n38808);
   U23791 : XOR2_X1 port map( A1 => n5323, A2 => n9518, Z => n11215);
   U23792 : OR2_X1 port map( A1 => n2416, A2 => n10665, Z => n31619);
   U23795 : INV_X2 port map( I => n29439, ZN => n1392);
   U23796 : AOI22_X1 port map( A1 => n7154, A2 => n38848, B1 => n31986, B2 => 
                           n24792, ZN => n9008);
   U23799 : XOR2_X1 port map( A1 => n25253, A2 => n38809, Z => n38815);
   U23800 : XOR2_X1 port map( A1 => n7250, A2 => n25104, Z => n25253);
   U23801 : INV_X2 port map( I => n38810, ZN => n15549);
   U23804 : AOI21_X2 port map( A1 => n26950, A2 => n13056, B => n1236, ZN => 
                           n38810);
   U23809 : OAI21_X2 port map( A1 => n32640, A2 => n17897, B => n20996, ZN => 
                           n17896);
   U23810 : NOR2_X2 port map( A1 => n19901, A2 => n37477, ZN => n38811);
   U23819 : XOR2_X1 port map( A1 => n35590, A2 => n39136, Z => n11311);
   U23823 : NAND2_X2 port map( A1 => n32282, A2 => n21959, ZN => n39136);
   U23825 : XOR2_X1 port map( A1 => n25251, A2 => n13763, Z => n38814);
   U23832 : NOR2_X2 port map( A1 => n26788, A2 => n1234, ZN => n2362);
   U23838 : OAI21_X2 port map( A1 => n19972, A2 => n1234, B => n26909, ZN => 
                           n26788);
   U23844 : OAI21_X2 port map( A1 => n24429, A2 => n10815, B => n38817, ZN => 
                           n39253);
   U23847 : OAI21_X2 port map( A1 => n18466, A2 => n14478, B => n24373, ZN => 
                           n38817);
   U23849 : NAND2_X2 port map( A1 => n16224, A2 => n30047, ZN => n11111);
   U23850 : NOR2_X2 port map( A1 => n26682, A2 => n30500, ZN => n32984);
   U23851 : OAI22_X2 port map( A1 => n38819, A2 => n30550, B1 => n6715, B2 => 
                           n38404, ZN => n35250);
   U23856 : AOI21_X2 port map( A1 => n16141, A2 => n6715, B => n10220, ZN => 
                           n38819);
   U23860 : XOR2_X1 port map( A1 => n2036, A2 => n38181, Z => n38820);
   U23863 : NAND2_X2 port map( A1 => n36016, A2 => n38821, ZN => n7769);
   U23865 : AOI21_X2 port map( A1 => n38823, A2 => n38822, B => n1061, ZN => 
                           n9869);
   U23867 : AOI21_X2 port map( A1 => n3988, A2 => n28568, B => n38826, ZN => 
                           n19571);
   U23868 : NAND2_X2 port map( A1 => n36124, A2 => n13378, ZN => n38826);
   U23876 : XOR2_X1 port map( A1 => n17342, A2 => n19825, Z => n5610);
   U23880 : AOI22_X2 port map( A1 => n17309, A2 => n32385, B1 => n11980, B2 => 
                           n38694, ZN => n17342);
   U23885 : NAND3_X2 port map( A1 => n27978, A2 => n27976, A3 => n37035, ZN => 
                           n28616);
   U23889 : XOR2_X1 port map( A1 => n12976, A2 => n38827, Z => n24431);
   U23891 : XOR2_X1 port map( A1 => n12798, A2 => n31466, Z => n38827);
   U23893 : NAND2_X2 port map( A1 => n38828, A2 => n17665, ZN => n3840);
   U23894 : NAND3_X1 port map( A1 => n12333, A2 => n9592, A3 => n35999, ZN => 
                           n38828);
   U23899 : NOR2_X2 port map( A1 => n20802, A2 => n25746, ZN => n26026);
   U23900 : XOR2_X1 port map( A1 => n542, A2 => n34391, Z => n5993);
   U23901 : OAI21_X2 port map( A1 => n35549, A2 => n35548, B => n32983, ZN => 
                           n542);
   U23902 : NAND3_X2 port map( A1 => n11286, A2 => n34416, A3 => n11776, ZN => 
                           n23903);
   U23905 : NAND3_X2 port map( A1 => n38831, A2 => n36957, A3 => n5172, ZN => 
                           n36509);
   U23911 : NAND3_X2 port map( A1 => n18945, A2 => n34847, A3 => n18944, ZN => 
                           n39772);
   U23912 : XOR2_X1 port map( A1 => n1660, A2 => n22656, Z => n13174);
   U23914 : NAND2_X2 port map( A1 => n18124, A2 => n10366, ZN => n31620);
   U23916 : AOI22_X2 port map( A1 => n38833, A2 => n22326, B1 => n22249, B2 => 
                           n31383, ZN => n13161);
   U23919 : INV_X2 port map( I => n13163, ZN => n38833);
   U23920 : NOR2_X2 port map( A1 => n30722, A2 => n37131, ZN => n26744);
   U23926 : XOR2_X1 port map( A1 => n28896, A2 => n28972, Z => n16336);
   U23929 : BUF_X2 port map( I => n30232, Z => n38834);
   U23947 : NAND2_X2 port map( A1 => n33703, A2 => n36810, ZN => n23400);
   U23949 : OAI21_X2 port map( A1 => n7629, A2 => n7630, B => n16058, ZN => 
                           n24065);
   U23951 : BUF_X2 port map( I => n39030, Z => n38835);
   U23952 : XOR2_X1 port map( A1 => n12145, A2 => n26150, Z => n7102);
   U23956 : INV_X2 port map( I => n22659, ZN => n1669);
   U23967 : XNOR2_X1 port map( A1 => Plaintext(93), A2 => Key(93), ZN => n33147
                           );
   U23973 : AOI21_X2 port map( A1 => n2644, A2 => n21944, B => n38836, ZN => 
                           n4342);
   U23982 : NOR2_X2 port map( A1 => n38837, A2 => n4982, ZN => n5439);
   U23990 : INV_X2 port map( I => n22729, ZN => n22628);
   U23992 : XOR2_X1 port map( A1 => n22729, A2 => n38838, Z => n509);
   U23993 : NOR2_X2 port map( A1 => n32551, A2 => n20239, ZN => n22729);
   U23994 : INV_X2 port map( I => n20352, ZN => n38838);
   U23995 : NAND2_X1 port map( A1 => n38840, A2 => n29210, ZN => n29102);
   U23998 : NAND2_X1 port map( A1 => n19765, A2 => n35870, ZN => n38840);
   U24002 : XOR2_X1 port map( A1 => n19571, A2 => n29254, Z => n29094);
   U24004 : NOR2_X2 port map( A1 => n19191, A2 => n34669, ZN => n34371);
   U24007 : XOR2_X1 port map( A1 => n8313, A2 => n17852, Z => n18229);
   U24010 : NAND2_X2 port map( A1 => n36535, A2 => n38841, ZN => n6282);
   U24011 : NAND2_X2 port map( A1 => n5928, A2 => n31424, ZN => n29142);
   U24012 : XOR2_X1 port map( A1 => n31599, A2 => n38021, Z => n2476);
   U24016 : XOR2_X1 port map( A1 => n38842, A2 => n1978, Z => n11297);
   U24017 : XOR2_X1 port map( A1 => n3157, A2 => n36529, Z => n28117);
   U24019 : XOR2_X1 port map( A1 => n33690, A2 => n3258, Z => n36529);
   U24021 : NOR2_X2 port map( A1 => n15159, A2 => n830, ZN => n38843);
   U24027 : XOR2_X1 port map( A1 => n38845, A2 => n37261, Z => Ciphertext(110))
                           ;
   U24030 : OAI22_X1 port map( A1 => n32466, A2 => n32467, B1 => n13606, B2 => 
                           n29812, ZN => n38845);
   U24038 : OR2_X1 port map( A1 => n37061, A2 => n33368, Z => n20370);
   U24045 : XOR2_X1 port map( A1 => n23952, A2 => n24002, Z => n14220);
   U24046 : XOR2_X1 port map( A1 => n38846, A2 => n22638, Z => n12760);
   U24047 : XNOR2_X1 port map( A1 => n22562, A2 => n22775, ZN => n22638);
   U24049 : XOR2_X1 port map( A1 => n34188, A2 => n37660, Z => n38846);
   U24054 : NAND2_X2 port map( A1 => n39182, A2 => n5494, ZN => n38847);
   U24056 : NOR2_X2 port map( A1 => n32745, A2 => n875, ZN => n30365);
   U24064 : INV_X1 port map( I => n16053, ZN => n22893);
   U24066 : NAND2_X1 port map( A1 => n35246, A2 => n19594, ZN => n16053);
   U24068 : XOR2_X1 port map( A1 => n16526, A2 => n19527, Z => n12297);
   U24070 : OAI21_X1 port map( A1 => n37734, A2 => n30220, B => n30158, ZN => 
                           n2322);
   U24072 : XOR2_X1 port map( A1 => n29057, A2 => n38962, Z => n9131);
   U24083 : XOR2_X1 port map( A1 => n12839, A2 => n30006, Z => n10598);
   U24084 : NAND2_X2 port map( A1 => n36949, A2 => n36951, ZN => n12839);
   U24086 : NAND2_X2 port map( A1 => n34010, A2 => n9526, ZN => n19785);
   U24088 : XNOR2_X1 port map( A1 => n13138, A2 => n18544, ZN => n38849);
   U24091 : NOR2_X2 port map( A1 => n6347, A2 => n22019, ZN => n7355);
   U24092 : INV_X2 port map( I => n22574, ZN => n35446);
   U24094 : BUF_X2 port map( I => n15439, Z => n38850);
   U24099 : BUF_X2 port map( I => n15794, Z => n38851);
   U24107 : XOR2_X1 port map( A1 => n27830, A2 => n15776, Z => n27635);
   U24108 : NAND2_X2 port map( A1 => n26890, A2 => n34113, ZN => n15776);
   U24109 : INV_X4 port map( I => n19998, ZN => n997);
   U24110 : NAND2_X2 port map( A1 => n3349, A2 => n19172, ZN => n19998);
   U24113 : NOR2_X1 port map( A1 => n13298, A2 => n34033, ZN => n39436);
   U24117 : AND2_X1 port map( A1 => n27137, A2 => n38853, Z => n34660);
   U24122 : NAND2_X2 port map( A1 => n34738, A2 => n9109, ZN => n2431);
   U24123 : NAND2_X2 port map( A1 => n31679, A2 => n35893, ZN => n7846);
   U24125 : NAND2_X2 port map( A1 => n3664, A2 => n28560, ZN => n28563);
   U24127 : XOR2_X1 port map( A1 => n2943, A2 => n16017, Z => n16019);
   U24138 : NAND2_X2 port map( A1 => n18625, A2 => n18624, ZN => n2943);
   U24142 : NAND2_X1 port map( A1 => n30548, A2 => n14845, ZN => n38859);
   U24143 : NAND2_X1 port map( A1 => n38614, A2 => n23423, ZN => n14163);
   U24144 : NAND2_X2 port map( A1 => n25635, A2 => n25634, ZN => n13712);
   U24146 : XOR2_X1 port map( A1 => n17727, A2 => n31214, Z => n22438);
   U24147 : NAND2_X2 port map( A1 => n3967, A2 => n3969, ZN => n31214);
   U24152 : XOR2_X1 port map( A1 => n12104, A2 => n12103, Z => n31784);
   U24161 : INV_X2 port map( I => n10940, ZN => n16590);
   U24163 : BUF_X2 port map( I => n14193, Z => n38860);
   U24168 : NOR2_X2 port map( A1 => n5156, A2 => n38861, ZN => n5154);
   U24171 : INV_X2 port map( I => n25261, ZN => n38862);
   U24183 : NOR2_X1 port map( A1 => n37052, A2 => n11727, ZN => n38863);
   U24190 : NOR2_X1 port map( A1 => n12370, A2 => n5456, ZN => n18670);
   U24191 : XOR2_X1 port map( A1 => n27541, A2 => n27581, Z => n32015);
   U24193 : NAND2_X2 port map( A1 => n16997, A2 => n17829, ZN => n27541);
   U24195 : OAI21_X2 port map( A1 => n38865, A2 => n38864, B => n21264, ZN => 
                           n11001);
   U24196 : NOR2_X2 port map( A1 => n32720, A2 => n29587, ZN => n38865);
   U24198 : XOR2_X1 port map( A1 => n11746, A2 => n11747, Z => n19783);
   U24204 : AOI22_X2 port map( A1 => n20791, A2 => n18920, B1 => n37468, B2 => 
                           n8735, ZN => n24113);
   U24207 : XOR2_X1 port map( A1 => n26489, A2 => n26553, Z => n12300);
   U24226 : NAND2_X2 port map( A1 => n7168, A2 => n7171, ZN => n26489);
   U24227 : AOI21_X2 port map( A1 => n32367, A2 => n32368, B => n1567, ZN => 
                           n38867);
   U24236 : OR2_X2 port map( A1 => n32854, A2 => n11342, Z => n30274);
   U24243 : NAND2_X2 port map( A1 => n10996, A2 => n38869, ZN => n22599);
   U24246 : XOR2_X1 port map( A1 => n39742, A2 => n27169, Z => n38870);
   U24249 : XOR2_X1 port map( A1 => n38872, A2 => n34152, Z => n34957);
   U24254 : XOR2_X1 port map( A1 => n15529, A2 => n26601, Z => n38872);
   U24257 : XNOR2_X1 port map( A1 => n36386, A2 => n27534, ZN => n479);
   U24261 : NAND2_X2 port map( A1 => n31302, A2 => n36805, ZN => n27534);
   U24265 : XOR2_X1 port map( A1 => n5516, A2 => n709, Z => n34200);
   U24266 : INV_X2 port map( I => n13311, ZN => n36251);
   U24267 : NOR2_X2 port map( A1 => n15289, A2 => n15290, ZN => n13311);
   U24283 : NOR2_X1 port map( A1 => n38874, A2 => n20053, ZN => n1997);
   U24289 : INV_X2 port map( I => n15925, ZN => n38874);
   U24290 : NAND2_X2 port map( A1 => n24795, A2 => n35981, ZN => n24597);
   U24293 : NAND2_X2 port map( A1 => n14051, A2 => n14050, ZN => n24795);
   U24294 : XOR2_X1 port map( A1 => n6717, A2 => n15162, Z => n38875);
   U24295 : XOR2_X1 port map( A1 => n820, A2 => n38876, Z => n13873);
   U24308 : XOR2_X1 port map( A1 => n14350, A2 => n25260, Z => n38876);
   U24314 : XOR2_X1 port map( A1 => n26590, A2 => n26357, Z => n26558);
   U24315 : OAI21_X2 port map( A1 => n12895, A2 => n4801, B => n25766, ZN => 
                           n26590);
   U24318 : BUF_X2 port map( I => n19202, Z => n38878);
   U24319 : AOI21_X2 port map( A1 => n15943, A2 => n1119, B => n38879, ZN => 
                           n16581);
   U24320 : NOR3_X2 port map( A1 => n38182, A2 => n3076, A3 => n30843, ZN => 
                           n38879);
   U24322 : XOR2_X1 port map( A1 => n23830, A2 => n38882, Z => n5086);
   U24323 : XOR2_X1 port map( A1 => n5959, A2 => n1612, Z => n38882);
   U24324 : XOR2_X1 port map( A1 => n23973, A2 => n9043, Z => n23850);
   U24334 : MUX2_X1 port map( I0 => n25931, I1 => n11888, S => n38247, Z => 
                           n15834);
   U24340 : XOR2_X1 port map( A1 => n33511, A2 => n7288, Z => n15810);
   U24341 : OR2_X1 port map( A1 => n19424, A2 => n29900, Z => n15358);
   U24342 : AND2_X1 port map( A1 => n28079, A2 => n20860, Z => n5022);
   U24344 : AOI21_X1 port map( A1 => n8520, A2 => n38976, B => n1687, ZN => 
                           n7897);
   U24345 : XOR2_X1 port map( A1 => n11308, A2 => n19221, Z => n22650);
   U24346 : NAND2_X2 port map( A1 => n7895, A2 => n11047, ZN => n11308);
   U24347 : XOR2_X1 port map( A1 => n28844, A2 => n2392, Z => n38885);
   U24348 : NOR2_X2 port map( A1 => n39687, A2 => n25450, ZN => n26048);
   U24349 : OAI22_X2 port map( A1 => n33459, A2 => n4957, B1 => n24172, B2 => 
                           n2268, ZN => n24625);
   U24352 : NAND2_X2 port map( A1 => n15559, A2 => n15558, ZN => n20346);
   U24353 : XOR2_X1 port map( A1 => n21036, A2 => n21149, Z => n21035);
   U24355 : INV_X2 port map( I => n38887, ZN => n39816);
   U24359 : XOR2_X1 port map( A1 => n11119, A2 => n11118, Z => n38887);
   U24362 : NOR2_X2 port map( A1 => n1635, A2 => n30881, ZN => n23256);
   U24363 : OAI22_X2 port map( A1 => n3803, A2 => n20840, B1 => n34013, B2 => 
                           n13635, ZN => n4143);
   U24372 : INV_X2 port map( I => n16265, ZN => n30315);
   U24376 : OAI22_X2 port map( A1 => n32663, A2 => n15926, B1 => n15929, B2 => 
                           n21694, ZN => n16265);
   U24377 : INV_X2 port map( I => n33258, ZN => n8006);
   U24380 : NAND3_X1 port map( A1 => n3906, A2 => n962, A3 => n15911, ZN => 
                           n12696);
   U24382 : OAI21_X2 port map( A1 => n19564, A2 => n27180, B => n33773, ZN => 
                           n27110);
   U24387 : OR2_X1 port map( A1 => n7843, A2 => n30800, Z => n22199);
   U24391 : NAND3_X2 port map( A1 => n20975, A2 => n4188, A3 => n17765, ZN => 
                           n24924);
   U24396 : XOR2_X1 port map( A1 => n38888, A2 => n3427, Z => n3424);
   U24404 : XOR2_X1 port map( A1 => n8183, A2 => n3426, Z => n38888);
   U24407 : XOR2_X1 port map( A1 => n38889, A2 => n25202, Z => n320);
   U24409 : XOR2_X1 port map( A1 => n38992, A2 => n25256, Z => n38889);
   U24410 : NAND2_X1 port map( A1 => n33879, A2 => n7901, ZN => n31432);
   U24421 : NAND2_X2 port map( A1 => n18599, A2 => n12416, ZN => n33879);
   U24422 : XOR2_X1 port map( A1 => n16556, A2 => n16558, Z => n38901);
   U24426 : XOR2_X1 port map( A1 => n5116, A2 => n23659, Z => n38890);
   U24427 : NAND2_X2 port map( A1 => n38891, A2 => n32789, ZN => n34692);
   U24428 : NAND3_X2 port map( A1 => n34940, A2 => n260, A3 => n34087, ZN => 
                           n38891);
   U24431 : AOI22_X2 port map( A1 => n38892, A2 => n23234, B1 => n20450, B2 => 
                           n23292, ZN => n35301);
   U24439 : XOR2_X1 port map( A1 => n25185, A2 => n38895, Z => n1817);
   U24442 : OAI21_X2 port map( A1 => n9367, A2 => n26929, B => n38912, ZN => 
                           n9369);
   U24446 : NAND2_X2 port map( A1 => n27562, A2 => n27078, ZN => n27731);
   U24452 : NAND2_X2 port map( A1 => n33908, A2 => n14086, ZN => n27562);
   U24458 : NAND2_X2 port map( A1 => n34913, A2 => n27085, ZN => n14058);
   U24472 : XOR2_X1 port map( A1 => n18807, A2 => n23814, Z => n19991);
   U24473 : NAND3_X2 port map( A1 => n15604, A2 => n15603, A3 => n14576, ZN => 
                           n18807);
   U24475 : NAND2_X2 port map( A1 => n38897, A2 => n2404, ZN => n22317);
   U24485 : OAI21_X2 port map( A1 => n2628, A2 => n21924, B => n38898, ZN => 
                           n38897);
   U24487 : OAI22_X2 port map( A1 => n35160, A2 => n16072, B1 => n16073, B2 => 
                           n34436, ZN => n35648);
   U24488 : BUF_X2 port map( I => n6390, Z => n38899);
   U24497 : XOR2_X1 port map( A1 => n33083, A2 => n29887, Z => n39141);
   U24503 : BUF_X2 port map( I => n14153, Z => n38900);
   U24505 : XOR2_X1 port map( A1 => n38902, A2 => n3701, Z => n15794);
   U24514 : XOR2_X1 port map( A1 => n39145, A2 => n10384, Z => n38902);
   U24528 : NAND2_X2 port map( A1 => n38904, A2 => n6048, ZN => n22574);
   U24536 : NAND2_X2 port map( A1 => n38921, A2 => n38920, ZN => n38904);
   U24542 : XOR2_X1 port map( A1 => n20152, A2 => n20151, Z => n20153);
   U24543 : NAND2_X1 port map( A1 => n39527, A2 => n32981, ZN => n34131);
   U24546 : XOR2_X1 port map( A1 => n6165, A2 => n30661, Z => n32981);
   U24547 : XOR2_X1 port map( A1 => n23936, A2 => n38905, Z => n7558);
   U24548 : XOR2_X1 port map( A1 => n25146, A2 => n38192, Z => n32346);
   U24551 : AOI21_X1 port map( A1 => n425, A2 => n15677, B => n11734, ZN => 
                           n25739);
   U24556 : INV_X2 port map( I => n34692, ZN => n425);
   U24560 : NOR2_X2 port map( A1 => n13607, A2 => n14600, ZN => n10606);
   U24562 : INV_X2 port map( I => n7643, ZN => n14600);
   U24567 : XOR2_X1 port map( A1 => n17906, A2 => n17905, Z => n7643);
   U24569 : NAND2_X2 port map( A1 => n7625, A2 => n38908, ZN => n38907);
   U24570 : NAND2_X2 port map( A1 => n26063, A2 => n25941, ZN => n38909);
   U24571 : AOI21_X2 port map( A1 => n7454, A2 => n28494, B => n35173, ZN => 
                           n1944);
   U24581 : NOR2_X2 port map( A1 => n9366, A2 => n7523, ZN => n38912);
   U24588 : XOR2_X1 port map( A1 => n28909, A2 => n38913, Z => n31089);
   U24590 : XOR2_X1 port map( A1 => n248, A2 => n17784, Z => n38913);
   U24594 : XOR2_X1 port map( A1 => n34752, A2 => n8844, Z => n19226);
   U24595 : NAND2_X2 port map( A1 => n3429, A2 => n12358, ZN => n34813);
   U24597 : OAI21_X2 port map( A1 => n23154, A2 => n22919, B => n14738, ZN => 
                           n33847);
   U24598 : NOR2_X2 port map( A1 => n8173, A2 => n5957, ZN => n24769);
   U24600 : OAI21_X2 port map( A1 => n33598, A2 => n30339, B => n28193, ZN => 
                           n31098);
   U24602 : OAI22_X2 port map( A1 => n36175, A2 => n3091, B1 => n26835, B2 => 
                           n16970, ZN => n31014);
   U24605 : NAND3_X2 port map( A1 => n23266, A2 => n23265, A3 => n23267, ZN => 
                           n23905);
   U24607 : AOI21_X2 port map( A1 => n17397, A2 => n7541, B => n28681, ZN => 
                           n28362);
   U24617 : INV_X2 port map( I => n13594, ZN => n28681);
   U24622 : NOR2_X2 port map( A1 => n2416, A2 => n37086, ZN => n25366);
   U24623 : NAND2_X1 port map( A1 => n28034, A2 => n36979, ZN => n27956);
   U24628 : BUF_X2 port map( I => n34350, Z => n38914);
   U24632 : NAND2_X2 port map( A1 => n38915, A2 => n36767, ZN => n34541);
   U24633 : NAND2_X2 port map( A1 => n19785, A2 => n17894, ZN => n38915);
   U24644 : NAND2_X2 port map( A1 => n928, A2 => n38914, ZN => n33109);
   U24650 : INV_X2 port map( I => n38916, ZN => n24910);
   U24651 : NAND2_X1 port map( A1 => n825, A2 => n25309, ZN => n19968);
   U24652 : XOR2_X1 port map( A1 => n25062, A2 => n25061, Z => n25309);
   U24653 : INV_X1 port map( I => n39460, ZN => n24073);
   U24660 : XOR2_X1 port map( A1 => n26381, A2 => n26516, Z => n21142);
   U24662 : NAND2_X2 port map( A1 => n25655, A2 => n34486, ZN => n26381);
   U24665 : XOR2_X1 port map( A1 => n23623, A2 => n24012, Z => n20777);
   U24667 : NAND2_X2 port map( A1 => n18123, A2 => n18370, ZN => n24012);
   U24668 : NOR2_X2 port map( A1 => n32483, A2 => n38918, ZN => n30504);
   U24670 : INV_X2 port map( I => n38922, ZN => n34040);
   U24672 : NAND2_X2 port map( A1 => n35443, A2 => n31986, ZN => n38922);
   U24676 : NAND2_X2 port map( A1 => n12279, A2 => n38925, ZN => n24545);
   U24681 : NAND2_X1 port map( A1 => n25943, A2 => n25345, ZN => n3926);
   U24685 : OAI22_X2 port map( A1 => n34083, A2 => n12599, B1 => n34487, B2 => 
                           n12601, ZN => n25943);
   U24690 : NAND2_X2 port map( A1 => n16250, A2 => n25989, ZN => n26081);
   U24692 : NAND2_X2 port map( A1 => n9479, A2 => n17173, ZN => n16250);
   U24694 : AND2_X2 port map( A1 => n14601, A2 => n35269, Z => n30348);
   U24697 : AOI22_X2 port map( A1 => n35137, A2 => n39317, B1 => n39406, B2 => 
                           n24879, ZN => n24547);
   U24705 : XOR2_X1 port map( A1 => n38927, A2 => n9436, Z => n9435);
   U24709 : NAND3_X1 port map( A1 => n36775, A2 => n19349, A3 => n38220, ZN => 
                           n7480);
   U24713 : NOR2_X2 port map( A1 => n35594, A2 => n38929, ZN => n13075);
   U24715 : NOR2_X1 port map( A1 => n25544, A2 => n15515, ZN => n9816);
   U24719 : OAI21_X1 port map( A1 => n25966, A2 => n18320, B => n25962, ZN => 
                           n38930);
   U24724 : NAND2_X2 port map( A1 => n38933, A2 => n35448, ZN => n5753);
   U24728 : NOR2_X2 port map( A1 => n26, A2 => n22317, ZN => n2028);
   U24742 : XOR2_X1 port map( A1 => n26475, A2 => n34630, Z => n14752);
   U24745 : XNOR2_X1 port map( A1 => n29242, A2 => n9035, ZN => n18526);
   U24746 : OAI22_X2 port map( A1 => n4878, A2 => n28664, B1 => n15580, B2 => 
                           n12990, ZN => n29242);
   U24747 : XOR2_X1 port map( A1 => n11867, A2 => n20692, Z => n35324);
   U24759 : XOR2_X1 port map( A1 => n3161, A2 => n38934, Z => n13039);
   U24783 : XOR2_X1 port map( A1 => n3778, A2 => n3777, Z => n38934);
   U24788 : NAND2_X2 port map( A1 => n37080, A2 => n18990, ZN => n19409);
   U24790 : NAND2_X2 port map( A1 => n1444, A2 => n33955, ZN => n28240);
   U24791 : INV_X4 port map( I => n38965, ZN => n34001);
   U24792 : XOR2_X1 port map( A1 => n29108, A2 => n38167, Z => n9972);
   U24795 : XOR2_X1 port map( A1 => n36255, A2 => n36254, Z => n2142);
   U24797 : AOI22_X2 port map( A1 => n12745, A2 => n9756, B1 => n12744, B2 => 
                           n7588, ZN => n17349);
   U24799 : XOR2_X1 port map( A1 => n5843, A2 => n38935, Z => n39570);
   U24800 : XOR2_X1 port map( A1 => n13935, A2 => n39609, Z => n38935);
   U24809 : XOR2_X1 port map( A1 => n20589, A2 => n4127, Z => n27692);
   U24813 : NAND2_X2 port map( A1 => n11089, A2 => n11087, ZN => n4127);
   U24826 : XOR2_X1 port map( A1 => n2170, A2 => n2168, Z => n10559);
   U24828 : NAND2_X2 port map( A1 => n39502, A2 => n38936, ZN => n15792);
   U24836 : OAI21_X2 port map( A1 => n10518, A2 => n10519, B => n11891, ZN => 
                           n38936);
   U24837 : INV_X2 port map( I => n20589, ZN => n38937);
   U24839 : XOR2_X1 port map( A1 => n8741, A2 => n33373, Z => n17064);
   U24841 : XOR2_X1 port map( A1 => n21077, A2 => n4856, Z => n21074);
   U24842 : NAND2_X1 port map( A1 => n3944, A2 => n5028, ZN => n28644);
   U24846 : XOR2_X1 port map( A1 => n523, A2 => n4393, Z => n3526);
   U24851 : OAI21_X2 port map( A1 => n38938, A2 => n14846, B => n21406, ZN => 
                           n22155);
   U24852 : NAND2_X2 port map( A1 => n19210, A2 => n16177, ZN => n38939);
   U24853 : XOR2_X1 port map( A1 => n25154, A2 => n38940, Z => n33058);
   U24861 : XOR2_X1 port map( A1 => n36980, A2 => n33208, Z => n38940);
   U24865 : XOR2_X1 port map( A1 => Plaintext(155), A2 => Key(155), Z => n39519
                           );
   U24869 : NAND2_X1 port map( A1 => n1265, A2 => n35893, ZN => n38942);
   U24870 : XOR2_X1 port map( A1 => n2436, A2 => n35425, Z => n16631);
   U24876 : XOR2_X1 port map( A1 => n4592, A2 => n9043, Z => n23961);
   U24880 : NAND2_X2 port map( A1 => n35285, A2 => n23648, ZN => n4592);
   U24883 : INV_X4 port map( I => n25956, ZN => n19740);
   U24885 : NAND2_X2 port map( A1 => n34541, A2 => n11954, ZN => n25956);
   U24889 : NAND2_X2 port map( A1 => n14896, A2 => n14897, ZN => n33996);
   U24893 : XOR2_X1 port map( A1 => n38943, A2 => n19677, Z => Ciphertext(163))
                           ;
   U24894 : OAI21_X1 port map( A1 => n21006, A2 => n21005, B => n30127, ZN => 
                           n38943);
   U24895 : OAI21_X1 port map( A1 => n8728, A2 => n38945, B => n38944, ZN => 
                           n29230);
   U24897 : AOI21_X2 port map( A1 => n36979, A2 => n14376, B => n38946, ZN => 
                           n13323);
   U24898 : NAND2_X2 port map( A1 => n28189, A2 => n16327, ZN => n38947);
   U24901 : XOR2_X1 port map( A1 => n10129, A2 => n27520, Z => n13751);
   U24904 : NAND2_X2 port map( A1 => n20245, A2 => n26806, ZN => n32191);
   U24905 : OAI22_X1 port map( A1 => n28736, A2 => n36935, B1 => n34861, B2 => 
                           n9686, ZN => n28059);
   U24907 : NAND2_X2 port map( A1 => n36209, A2 => n36640, ZN => n35901);
   U24910 : NAND2_X2 port map( A1 => n6800, A2 => n6799, ZN => n39489);
   U24911 : NAND3_X2 port map( A1 => n2417, A2 => n20881, A3 => n30694, ZN => 
                           n38949);
   U24918 : XOR2_X1 port map( A1 => n38209, A2 => n7481, Z => n13324);
   U24923 : NAND2_X1 port map( A1 => n29596, A2 => n29592, ZN => n9865);
   U24925 : XOR2_X1 port map( A1 => n25139, A2 => n25138, Z => n25619);
   U24931 : NAND2_X2 port map( A1 => n38952, A2 => n34967, ZN => n4246);
   U24935 : NAND2_X2 port map( A1 => n26081, A2 => n38953, ZN => n38952);
   U24936 : NOR2_X1 port map( A1 => n9135, A2 => n35314, ZN => n15715);
   U24943 : XOR2_X1 port map( A1 => n19374, A2 => n29151, Z => n16193);
   U24949 : XOR2_X1 port map( A1 => n38954, A2 => n14866, Z => n30946);
   U24950 : XOR2_X1 port map( A1 => n26508, A2 => n39596, Z => n38954);
   U24958 : NOR2_X1 port map( A1 => n19700, A2 => n19364, ZN => n35297);
   U24963 : NAND2_X2 port map( A1 => n5983, A2 => n31110, ZN => n31535);
   U24967 : XOR2_X1 port map( A1 => n22749, A2 => n22580, Z => n22752);
   U24976 : NOR2_X2 port map( A1 => n17637, A2 => n17634, ZN => n22749);
   U24977 : AOI21_X2 port map( A1 => n37104, A2 => n30859, B => n26990, ZN => 
                           n38955);
   U24982 : XOR2_X1 port map( A1 => n5233, A2 => n37214, Z => n39347);
   U24986 : NAND2_X2 port map( A1 => n8977, A2 => n11924, ZN => n19580);
   U24988 : INV_X2 port map( I => n20297, ZN => n29346);
   U24989 : XOR2_X1 port map( A1 => n13358, A2 => n13052, Z => n20297);
   U24990 : OAI21_X2 port map( A1 => n38956, A2 => n37239, B => n424, ZN => 
                           n6845);
   U24992 : INV_X2 port map( I => n27137, ZN => n27350);
   U24993 : NAND2_X2 port map( A1 => n39041, A2 => n34974, ZN => n27137);
   U24996 : NAND2_X2 port map( A1 => n3263, A2 => n14933, ZN => n18070);
   U24998 : OR2_X1 port map( A1 => n17197, A2 => n20056, Z => n27929);
   U25007 : AOI21_X2 port map( A1 => n1108, A2 => n952, B => n17029, ZN => 
                           n10530);
   U25010 : NAND3_X2 port map( A1 => n3806, A2 => n3807, A3 => n32035, ZN => 
                           n8972);
   U25022 : AOI22_X2 port map( A1 => n5020, A2 => n28168, B1 => n28167, B2 => 
                           n7528, ZN => n38957);
   U25023 : AOI22_X2 port map( A1 => n8355, A2 => n14857, B1 => n12633, B2 => 
                           n12632, ZN => n25252);
   U25032 : NAND2_X1 port map( A1 => n9633, A2 => n38193, ZN => n27114);
   U25033 : INV_X1 port map( I => n18526, ZN => n31822);
   U25036 : AOI21_X2 port map( A1 => n9599, A2 => n35888, B => n4992, ZN => 
                           n4991);
   U25037 : XOR2_X1 port map( A1 => n7328, A2 => n25319, Z => n36039);
   U25042 : BUF_X2 port map( I => n30494, Z => n38960);
   U25047 : INV_X2 port map( I => n8423, ZN => n35369);
   U25050 : NAND3_X2 port map( A1 => n14116, A2 => n14115, A3 => n10032, ZN => 
                           n27810);
   U25055 : AOI22_X2 port map( A1 => n6097, A2 => n2835, B1 => n5327, B2 => 
                           n1519, ZN => n26365);
   U25065 : XOR2_X1 port map( A1 => n31617, A2 => n22203, Z => n780);
   U25069 : NAND2_X2 port map( A1 => n30603, A2 => n34252, ZN => n30764);
   U25072 : NAND2_X2 port map( A1 => n36187, A2 => n38961, ZN => n11003);
   U25091 : NAND3_X1 port map( A1 => n34103, A2 => n34411, A3 => n13943, ZN => 
                           n38961);
   U25092 : XOR2_X1 port map( A1 => n36497, A2 => n4540, Z => n33848);
   U25093 : XOR2_X1 port map( A1 => n34718, A2 => n38962, Z => n660);
   U25096 : XOR2_X1 port map( A1 => n1238, A2 => n26476, Z => n26522);
   U25097 : NAND2_X2 port map( A1 => n35992, A2 => n8133, ZN => n26476);
   U25109 : NAND2_X2 port map( A1 => n39002, A2 => n35839, ZN => n18686);
   U25113 : OR2_X1 port map( A1 => n25639, A2 => n38963, Z => n39053);
   U25114 : NAND2_X2 port map( A1 => n2798, A2 => n39401, ZN => n10739);
   U25122 : OR2_X2 port map( A1 => n20945, A2 => n10816, Z => n13607);
   U25125 : XOR2_X1 port map( A1 => n20618, A2 => n34856, Z => n2209);
   U25126 : XOR2_X1 port map( A1 => n36668, A2 => n29820, Z => n17159);
   U25131 : INV_X2 port map( I => n38966, ZN => n14081);
   U25133 : XOR2_X1 port map( A1 => n8887, A2 => n29258, Z => n35142);
   U25136 : XOR2_X1 port map( A1 => n38968, A2 => n19217, Z => n26545);
   U25139 : XOR2_X1 port map( A1 => n27193, A2 => n27194, Z => n38969);
   U25142 : OAI21_X2 port map( A1 => n19379, A2 => n16774, B => n38971, ZN => 
                           n1919);
   U25145 : OAI21_X2 port map( A1 => n19070, A2 => n8041, B => n24257, ZN => 
                           n23652);
   U25146 : NAND2_X2 port map( A1 => n33104, A2 => n38972, ZN => n24257);
   U25158 : INV_X2 port map( I => n18269, ZN => n38972);
   U25164 : XOR2_X1 port map( A1 => n38974, A2 => n13967, Z => n33576);
   U25173 : XOR2_X1 port map( A1 => n39582, A2 => n25238, Z => n38974);
   U25175 : XOR2_X1 port map( A1 => n26529, A2 => n26527, Z => n5312);
   U25177 : XOR2_X1 port map( A1 => n1986, A2 => n39529, Z => n15853);
   U25180 : XOR2_X1 port map( A1 => n1791, A2 => n38975, Z => n39433);
   U25182 : NAND2_X2 port map( A1 => n32524, A2 => n34301, ZN => n7744);
   U25196 : AOI22_X2 port map( A1 => n39283, A2 => n4781, B1 => n27306, B2 => 
                           n26791, ZN => n32248);
   U25198 : XOR2_X1 port map( A1 => n38977, A2 => n18700, Z => Ciphertext(45));
   U25203 : NOR2_X1 port map( A1 => n19689, A2 => n29436, ZN => n38977);
   U25205 : XOR2_X1 port map( A1 => n27717, A2 => n37881, Z => n10562);
   U25208 : NAND2_X2 port map( A1 => n36343, A2 => n30373, ZN => n24802);
   U25209 : NAND2_X2 port map( A1 => n25954, A2 => n365, ZN => n36008);
   U25213 : NAND2_X1 port map( A1 => n22473, A2 => n34131, ZN => n39199);
   U25217 : BUF_X2 port map( I => n26421, Z => n38979);
   U25219 : AOI21_X2 port map( A1 => n38980, A2 => n18877, B => n12142, ZN => 
                           n22292);
   U25227 : NAND2_X2 port map( A1 => n36358, A2 => n15626, ZN => n38980);
   U25237 : OR2_X1 port map( A1 => n25861, A2 => n1107, Z => n12710);
   U25239 : INV_X1 port map( I => n33997, ZN => n38982);
   U25240 : NAND2_X2 port map( A1 => n4150, A2 => n4151, ZN => n28104);
   U25242 : NAND2_X2 port map( A1 => n3914, A2 => n34939, ZN => n7018);
   U25247 : NAND2_X2 port map( A1 => n12171, A2 => n12170, ZN => n14153);
   U25249 : NOR2_X2 port map( A1 => n31876, A2 => n32869, ZN => n1882);
   U25251 : NOR2_X2 port map( A1 => n15890, A2 => n33792, ZN => n39528);
   U25254 : NOR3_X2 port map( A1 => n38600, A2 => n15176, A3 => n17511, ZN => 
                           n35322);
   U25256 : XOR2_X1 port map( A1 => n38985, A2 => n701, Z => n12471);
   U25258 : XOR2_X1 port map( A1 => n13652, A2 => n22520, Z => n38985);
   U25262 : INV_X2 port map( I => n20570, ZN => n38986);
   U25264 : AOI21_X2 port map( A1 => n18484, A2 => n24228, B => n38987, ZN => 
                           n20229);
   U25268 : OAI21_X2 port map( A1 => n30379, A2 => n2396, B => n2400, ZN => 
                           n38987);
   U25269 : XOR2_X1 port map( A1 => n18493, A2 => n29119, Z => n38988);
   U25271 : XOR2_X1 port map( A1 => n6989, A2 => n26599, Z => n26288);
   U25280 : XOR2_X1 port map( A1 => n34653, A2 => n14374, Z => n38989);
   U25281 : AOI22_X2 port map( A1 => n24113, A2 => n18615, B1 => n24112, B2 => 
                           n24111, ZN => n15281);
   U25282 : XOR2_X1 port map( A1 => n38990, A2 => n1356, Z => Ciphertext(95));
   U25287 : NOR2_X2 port map( A1 => n39101, A2 => n5949, ZN => n38990);
   U25289 : XOR2_X1 port map( A1 => n9930, A2 => n29092, Z => n12562);
   U25290 : NAND2_X1 port map( A1 => n33964, A2 => n17698, ZN => n29694);
   U25292 : NAND2_X2 port map( A1 => n33843, A2 => n15022, ZN => n13879);
   U25293 : NAND2_X2 port map( A1 => n5994, A2 => n34836, ZN => n3963);
   U25294 : XOR2_X1 port map( A1 => n38991, A2 => Key(151), Z => n39031);
   U25300 : XOR2_X1 port map( A1 => n39024, A2 => n18452, Z => n6449);
   U25313 : OAI21_X2 port map( A1 => n18501, A2 => n23193, B => n23192, ZN => 
                           n39070);
   U25320 : OAI21_X2 port map( A1 => n26619, A2 => n1236, B => n14271, ZN => 
                           n26618);
   U25326 : BUF_X2 port map( I => n25006, Z => n38993);
   U25329 : XOR2_X1 port map( A1 => n34902, A2 => n38994, Z => n3404);
   U25336 : XOR2_X1 port map( A1 => n990, A2 => n31602, Z => n38994);
   U25338 : XOR2_X1 port map( A1 => n7689, A2 => n39766, Z => n13062);
   U25344 : NOR2_X2 port map( A1 => n38995, A2 => n18538, ZN => n23912);
   U25347 : NOR3_X1 port map( A1 => n29813, A2 => n38141, A3 => n2792, ZN => 
                           n6650);
   U25358 : XOR2_X1 port map( A1 => n16019, A2 => n28947, Z => n31031);
   U25365 : NAND2_X2 port map( A1 => n38999, A2 => n38998, ZN => n38997);
   U25367 : NAND2_X1 port map( A1 => n28644, A2 => n28729, ZN => n39000);
   U25372 : OAI21_X1 port map( A1 => n20368, A2 => n21950, B => n39658, ZN => 
                           n21786);
   U25375 : NAND2_X1 port map( A1 => n6405, A2 => n39423, ZN => n28382);
   U25376 : NAND2_X2 port map( A1 => n12751, A2 => n12752, ZN => n39002);
   U25382 : OR2_X1 port map( A1 => n29543, A2 => n39003, Z => n7437);
   U25385 : OAI22_X2 port map( A1 => n14744, A2 => n39004, B1 => n14743, B2 => 
                           n9797, ZN => n23613);
   U25388 : NAND2_X2 port map( A1 => n6254, A2 => n39005, ZN => n6253);
   U25391 : OAI21_X2 port map( A1 => n21001, A2 => n19486, B => n39007, ZN => 
                           n22284);
   U25392 : AOI22_X2 port map( A1 => n24290, A2 => n7949, B1 => n1274, B2 => 
                           n8690, ZN => n39538);
   U25395 : NOR2_X2 port map( A1 => n13970, A2 => n232, ZN => n24290);
   U25398 : INV_X4 port map( I => n39108, ZN => n840);
   U25403 : XOR2_X1 port map( A1 => n39008, A2 => n24057, Z => n36066);
   U25406 : XOR2_X1 port map( A1 => n14023, A2 => n8920, Z => n24930);
   U25409 : AOI22_X2 port map( A1 => n5921, A2 => n14337, B1 => n29719, B2 => 
                           n29720, ZN => n29723);
   U25411 : NAND2_X2 port map( A1 => n27343, A2 => n39009, ZN => n34113);
   U25420 : NOR2_X2 port map( A1 => n27344, A2 => n7620, ZN => n39009);
   U25432 : NAND2_X2 port map( A1 => n13875, A2 => n14277, ZN => n36827);
   U25439 : INV_X2 port map( I => n39011, ZN => n921);
   U25441 : XOR2_X1 port map( A1 => n2547, A2 => n30578, Z => n39011);
   U25447 : BUF_X2 port map( I => n36539, Z => n39012);
   U25453 : XOR2_X1 port map( A1 => n39665, A2 => n9243, Z => n24318);
   U25455 : XOR2_X1 port map( A1 => n32298, A2 => n27796, Z => n32149);
   U25456 : AOI21_X2 port map( A1 => n2377, A2 => n26871, B => n36806, ZN => 
                           n32298);
   U25466 : OAI21_X2 port map( A1 => n30421, A2 => n24658, B => n1121, ZN => 
                           n39013);
   U25468 : NAND2_X2 port map( A1 => n2796, A2 => n31657, ZN => n36539);
   U25471 : NOR2_X2 port map( A1 => n10030, A2 => n30675, ZN => n197);
   U25472 : OR2_X1 port map( A1 => n1109, A2 => n19153, Z => n39800);
   U25480 : XOR2_X1 port map( A1 => n20794, A2 => n32083, Z => n20591);
   U25483 : OAI22_X2 port map( A1 => n22127, A2 => n22255, B1 => n31481, B2 => 
                           n937, ZN => n22731);
   U25485 : NAND2_X2 port map( A1 => n24440, A2 => n19584, ZN => n33457);
   U25486 : BUF_X2 port map( I => n18661, Z => n39015);
   U25489 : NAND2_X2 port map( A1 => n1949, A2 => n39016, ZN => n15426);
   U25493 : AOI21_X2 port map( A1 => n31913, A2 => n20157, B => n39069, ZN => 
                           n13727);
   U25495 : XOR2_X1 port map( A1 => n13736, A2 => n16175, Z => n10769);
   U25497 : OAI22_X2 port map( A1 => n39248, A2 => n26111, B1 => n16860, B2 => 
                           n26112, ZN => n14226);
   U25515 : BUF_X2 port map( I => n16803, Z => n39019);
   U25519 : NOR2_X1 port map( A1 => n16931, A2 => n32486, ZN => n25641);
   U25529 : NAND2_X2 port map( A1 => n39749, A2 => n32871, ZN => n6590);
   U25530 : NAND2_X2 port map( A1 => n14759, A2 => n15953, ZN => n23117);
   U25534 : NAND2_X2 port map( A1 => n32133, A2 => n18034, ZN => n14759);
   U25535 : XOR2_X1 port map( A1 => n33470, A2 => n38144, Z => n16218);
   U25539 : NAND2_X2 port map( A1 => n5377, A2 => n31273, ZN => n33470);
   U25544 : NAND4_X2 port map( A1 => n34292, A2 => n30062, A3 => n35095, A4 => 
                           n39022, ZN => n39695);
   U25545 : NAND2_X2 port map( A1 => n39023, A2 => n16848, ZN => n27854);
   U25546 : NOR2_X2 port map( A1 => n16211, A2 => n24545, ZN => n24658);
   U25557 : XOR2_X1 port map( A1 => n29001, A2 => n29000, Z => n39024);
   U25562 : XOR2_X1 port map( A1 => n27626, A2 => n11236, Z => n18094);
   U25567 : XOR2_X1 port map( A1 => n35270, A2 => n13289, Z => n27626);
   U25573 : AOI21_X1 port map( A1 => n34534, A2 => n29477, B => n1396, ZN => 
                           n12150);
   U25574 : INV_X2 port map( I => n29468, ZN => n1396);
   U25576 : NOR2_X2 port map( A1 => n23250, A2 => n30299, ZN => n7631);
   U25579 : NAND2_X2 port map( A1 => n33526, A2 => n32943, ZN => n30299);
   U25580 : XOR2_X1 port map( A1 => n12798, A2 => n24045, Z => n16765);
   U25584 : XOR2_X1 port map( A1 => n23697, A2 => n476, Z => n24045);
   U25590 : AND2_X1 port map( A1 => n36995, A2 => n28024, Z => n20968);
   U25593 : NAND3_X1 port map( A1 => n34482, A2 => n1101, A3 => n7110, ZN => 
                           n17312);
   U25598 : NOR3_X2 port map( A1 => n33081, A2 => n15651, A3 => n4893, ZN => 
                           n39026);
   U25601 : XOR2_X1 port map( A1 => n39027, A2 => n8119, Z => n35143);
   U25603 : NAND2_X2 port map( A1 => n12176, A2 => n11373, ZN => n18110);
   U25608 : NAND2_X2 port map( A1 => n30853, A2 => n35967, ZN => n26627);
   U25610 : XOR2_X1 port map( A1 => n22771, A2 => n13961, Z => n39028);
   U25611 : XOR2_X1 port map( A1 => n27804, A2 => n39029, Z => n4362);
   U25613 : XOR2_X1 port map( A1 => n1464, A2 => n35190, Z => n39029);
   U25616 : INV_X2 port map( I => n7846, ZN => n14523);
   U25621 : INV_X2 port map( I => n39031, ZN => n35116);
   U25626 : OAI21_X2 port map( A1 => n13351, A2 => n13350, B => n5613, ZN => 
                           n37016);
   U25627 : NAND2_X2 port map( A1 => n34715, A2 => n32032, ZN => n15558);
   U25631 : XOR2_X1 port map( A1 => n16898, A2 => n22563, Z => n22712);
   U25633 : NOR2_X2 port map( A1 => n35668, A2 => n6557, ZN => n16898);
   U25634 : NAND2_X1 port map( A1 => n6949, A2 => n39152, ZN => n22330);
   U25637 : INV_X2 port map( I => n39033, ZN => n34064);
   U25641 : OAI21_X2 port map( A1 => n34387, A2 => n4743, B => n16263, ZN => 
                           n10356);
   U25642 : AOI21_X2 port map( A1 => n10352, A2 => n10351, B => n39035, ZN => 
                           n10349);
   U25653 : NOR2_X2 port map( A1 => n30338, A2 => n28024, ZN => n39035);
   U25657 : OAI21_X2 port map( A1 => n35075, A2 => n34690, B => n33077, ZN => 
                           n24455);
   U25659 : NAND2_X2 port map( A1 => n23766, A2 => n23765, ZN => n13045);
   U25663 : NOR2_X1 port map( A1 => n38728, A2 => n38732, ZN => n34076);
   U25665 : NAND3_X2 port map( A1 => n4038, A2 => n1217, A3 => n37076, ZN => 
                           n39036);
   U25667 : XOR2_X1 port map( A1 => n13914, A2 => n5003, Z => n26625);
   U25668 : XOR2_X1 port map( A1 => n15093, A2 => n2782, Z => n39219);
   U25671 : BUF_X2 port map( I => n15737, Z => n39037);
   U25673 : XOR2_X1 port map( A1 => n39040, A2 => n39039, Z => n39472);
   U25675 : NOR2_X2 port map( A1 => n32016, A2 => n31018, ZN => n39041);
   U25684 : INV_X4 port map( I => n27338, ZN => n1225);
   U25693 : NAND2_X2 port map( A1 => n81, A2 => n35772, ZN => n27338);
   U25695 : OAI22_X2 port map( A1 => n25491, A2 => n9594, B1 => n16113, B2 => 
                           n20924, ZN => n33997);
   U25697 : XOR2_X1 port map( A1 => n39447, A2 => n39042, Z => n4291);
   U25698 : XOR2_X1 port map( A1 => n22394, A2 => n22557, Z => n39042);
   U25702 : INV_X2 port map( I => n39043, ZN => n22925);
   U25705 : XOR2_X1 port map( A1 => n25167, A2 => n30330, Z => n39044);
   U25706 : NAND2_X2 port map( A1 => n39046, A2 => n22926, ZN => n39045);
   U25708 : NAND2_X2 port map( A1 => n1235, A2 => n9618, ZN => n14825);
   U25715 : NOR2_X2 port map( A1 => n18055, A2 => n18056, ZN => n20806);
   U25716 : INV_X4 port map( I => n8942, ZN => n8707);
   U25718 : AND2_X1 port map( A1 => n13492, A2 => n12909, Z => n28035);
   U25724 : NAND2_X2 port map( A1 => n6556, A2 => n14233, ZN => n22563);
   U25729 : XOR2_X1 port map( A1 => n24037, A2 => n18849, Z => n39049);
   U25734 : OAI22_X2 port map( A1 => n2491, A2 => n13588, B1 => n34892, B2 => 
                           n26727, ZN => n39051);
   U25735 : INV_X2 port map( I => n39052, ZN => n19410);
   U25736 : XNOR2_X1 port map( A1 => n27646, A2 => n8424, ZN => n39052);
   U25741 : AOI21_X2 port map( A1 => n22999, A2 => n9797, B => n37062, ZN => 
                           n32614);
   U25743 : XOR2_X1 port map( A1 => n37498, A2 => n25123, Z => n13935);
   U25746 : OAI22_X2 port map( A1 => n24744, A2 => n24547, B1 => n11751, B2 => 
                           n11642, ZN => n25123);
   U25747 : AOI22_X2 port map( A1 => n10698, A2 => n37674, B1 => n23052, B2 => 
                           n14556, ZN => n33087);
   U25761 : XOR2_X1 port map( A1 => n23781, A2 => n24073, Z => n2107);
   U25763 : INV_X2 port map( I => n39054, ZN => n30285);
   U25764 : NOR2_X2 port map( A1 => n12360, A2 => n39055, ZN => n32152);
   U25769 : NAND2_X1 port map( A1 => n4525, A2 => n37088, ZN => n39434);
   U25772 : XOR2_X1 port map( A1 => n27707, A2 => n29394, Z => n7651);
   U25777 : NAND2_X2 port map( A1 => n20914, A2 => n32245, ZN => n27707);
   U25779 : NAND2_X1 port map( A1 => n2630, A2 => n32471, ZN => n39056);
   U25780 : AND2_X1 port map( A1 => n23682, A2 => n2394, Z => n39057);
   U25785 : XOR2_X1 port map( A1 => n12300, A2 => n33233, Z => n39058);
   U25787 : NAND2_X1 port map( A1 => n39059, A2 => n37341, ZN => n13901);
   U25789 : AOI21_X2 port map( A1 => n12802, A2 => n12804, B => n12800, ZN => 
                           n10054);
   U25792 : INV_X2 port map( I => n24761, ZN => n39059);
   U25793 : XOR2_X1 port map( A1 => n22629, A2 => n22652, Z => n22787);
   U25796 : OAI22_X2 port map( A1 => n22077, A2 => n20354, B1 => n20355, B2 => 
                           n22078, ZN => n22629);
   U25803 : NAND2_X2 port map( A1 => n13727, A2 => n13726, ZN => n36935);
   U25809 : BUF_X2 port map( I => n26180, Z => n39063);
   U25813 : NAND2_X2 port map( A1 => n39730, A2 => n8208, ZN => n27581);
   U25822 : INV_X1 port map( I => n3499, ZN => n39115);
   U25827 : NOR3_X1 port map( A1 => n39271, A2 => n24410, A3 => n37467, ZN => 
                           n32818);
   U25828 : INV_X2 port map( I => n10559, ZN => n39648);
   U25839 : NOR2_X2 port map( A1 => n39480, A2 => n31443, ZN => n39138);
   U25843 : AOI21_X2 port map( A1 => n11513, A2 => n17047, B => n39064, ZN => 
                           n26353);
   U25846 : INV_X2 port map( I => n34279, ZN => n39065);
   U25849 : INV_X2 port map( I => n27546, ZN => n20829);
   U25854 : OAI22_X2 port map( A1 => n3920, A2 => n27240, B1 => n3921, B2 => 
                           n35466, ZN => n27546);
   U25857 : AOI22_X1 port map( A1 => n24302, A2 => n24461, B1 => n14509, B2 => 
                           n19990, ZN => n39796);
   U25861 : AOI21_X2 port map( A1 => n39066, A2 => n17269, B => n25925, ZN => 
                           n18630);
   U25866 : AOI21_X2 port map( A1 => n39068, A2 => n31603, B => n9025, ZN => 
                           n7893);
   U25868 : NOR2_X2 port map( A1 => n10702, A2 => n30240, ZN => n39068);
   U25871 : INV_X4 port map( I => n30211, ZN => n39083);
   U25874 : NOR2_X1 port map( A1 => n28119, A2 => n28049, ZN => n39069);
   U25876 : OAI22_X1 port map( A1 => n1126, A2 => n37267, B1 => n19864, B2 => 
                           n30279, ZN => n31916);
   U25877 : XOR2_X1 port map( A1 => n27710, A2 => n27781, Z => n11730);
   U25879 : XOR2_X1 port map( A1 => n23684, A2 => n23683, Z => n39071);
   U25882 : NAND2_X2 port map( A1 => n2628, A2 => n9316, ZN => n3429);
   U25890 : NOR2_X2 port map( A1 => n18657, A2 => n33899, ZN => n2628);
   U25895 : NAND2_X2 port map( A1 => n39072, A2 => n35729, ZN => n27755);
   U25907 : MUX2_X1 port map( I0 => n27119, I1 => n27118, S => n32976, Z => 
                           n39072);
   U25913 : NAND2_X2 port map( A1 => n39501, A2 => n24673, ZN => n18115);
   U25915 : OAI21_X2 port map( A1 => n39165, A2 => n692, B => n13971, ZN => 
                           n17374);
   U25917 : NOR2_X2 port map( A1 => n2798, A2 => n10143, ZN => n8680);
   U25926 : BUF_X2 port map( I => n24470, Z => n39074);
   U25933 : OAI22_X2 port map( A1 => n18862, A2 => n26038, B1 => n18863, B2 => 
                           n25921, ZN => n26511);
   U25935 : XOR2_X1 port map( A1 => n36851, A2 => n8177, Z => n8176);
   U25938 : XOR2_X1 port map( A1 => n6746, A2 => n24075, Z => n31655);
   U25942 : AND2_X1 port map( A1 => n25490, A2 => n34427, Z => n4715);
   U25947 : AOI22_X1 port map( A1 => n5723, A2 => n36965, B1 => n35963, B2 => 
                           n31931, ZN => n8052);
   U25954 : NAND2_X2 port map( A1 => n33087, A2 => n8101, ZN => n31931);
   U25955 : BUF_X4 port map( I => n36281, Z => n39075);
   U25958 : INV_X1 port map( I => n39076, ZN => n2898);
   U25960 : INV_X2 port map( I => n23918, ZN => n36497);
   U25968 : XOR2_X1 port map( A1 => n24034, A2 => n6560, Z => n23918);
   U25970 : OAI21_X1 port map( A1 => n20242, A2 => n21782, B => n32123, ZN => 
                           n21663);
   U25981 : OAI22_X2 port map( A1 => n32202, A2 => n9798, B1 => n13451, B2 => 
                           n13450, ZN => n23580);
   U25985 : OAI21_X2 port map( A1 => n34081, A2 => n13320, B => n35419, ZN => 
                           n39077);
   U25987 : INV_X2 port map( I => n26361, ZN => n39078);
   U25988 : NAND2_X2 port map( A1 => n10510, A2 => n10509, ZN => n26361);
   U25992 : NOR2_X1 port map( A1 => n20242, A2 => n32123, ZN => n20241);
   U25993 : OAI21_X1 port map( A1 => n14438, A2 => n3700, B => n3631, ZN => 
                           n2859);
   U25999 : XOR2_X1 port map( A1 => n39080, A2 => n29036, Z => n2122);
   U26000 : XOR2_X1 port map( A1 => n29095, A2 => n19309, Z => n39080);
   U26003 : XOR2_X1 port map( A1 => n22482, A2 => n39081, Z => n130);
   U26007 : XOR2_X1 port map( A1 => n22768, A2 => n33990, Z => n39081);
   U26008 : XOR2_X1 port map( A1 => n3649, A2 => n39082, Z => n30330);
   U26019 : INV_X1 port map( I => n19953, ZN => n39082);
   U26039 : AOI21_X2 port map( A1 => n21505, A2 => n10345, B => n32319, ZN => 
                           n22254);
   U26045 : OAI21_X2 port map( A1 => n31696, A2 => n30155, B => n32777, ZN => 
                           n18589);
   U26049 : OAI21_X2 port map( A1 => n39107, A2 => n787, B => n39084, ZN => 
                           n11678);
   U26050 : OAI21_X2 port map( A1 => n10018, A2 => n9841, B => n20873, ZN => 
                           n39084);
   U26051 : NOR2_X2 port map( A1 => n35116, A2 => n37111, ZN => n15019);
   U26052 : XOR2_X1 port map( A1 => n27664, A2 => n27574, Z => n27495);
   U26055 : NOR2_X2 port map( A1 => n13721, A2 => n20149, ZN => n27664);
   U26057 : AND2_X1 port map( A1 => n22294, A2 => n22292, Z => n22139);
   U26058 : XOR2_X1 port map( A1 => n39086, A2 => n34152, Z => n19459);
   U26060 : XOR2_X1 port map( A1 => n36508, A2 => n21142, Z => n39086);
   U26067 : NAND2_X2 port map( A1 => n8350, A2 => n39087, ZN => n28692);
   U26069 : NAND2_X2 port map( A1 => n36404, A2 => n2625, ZN => n31665);
   U26071 : XOR2_X1 port map( A1 => n13115, A2 => n29038, Z => n39088);
   U26072 : XOR2_X1 port map( A1 => n1258, A2 => n14385, Z => n25063);
   U26073 : XOR2_X1 port map( A1 => n29096, A2 => n29063, Z => n19600);
   U26074 : NAND3_X2 port map( A1 => n14049, A2 => n6068, A3 => n6071, ZN => 
                           n29096);
   U26076 : NAND2_X1 port map( A1 => n13384, A2 => n38163, ZN => n9263);
   U26080 : XOR2_X1 port map( A1 => n2637, A2 => n39088, Z => n29184);
   U26081 : XOR2_X1 port map( A1 => n18620, A2 => n39089, Z => n35164);
   U26082 : XOR2_X1 port map( A1 => n23833, A2 => n18622, Z => n39089);
   U26084 : NAND2_X2 port map( A1 => n39498, A2 => n6541, ZN => n25319);
   U26087 : XOR2_X1 port map( A1 => n39090, A2 => n39310, Z => n3804);
   U26089 : XOR2_X1 port map( A1 => n23885, A2 => n1622, Z => n39090);
   U26095 : NAND2_X1 port map( A1 => n39091, A2 => n1451, ZN => n19413);
   U26096 : OAI22_X1 port map( A1 => n983, A2 => n28050, B1 => n14404, B2 => 
                           n28124, ZN => n39091);
   U26100 : XOR2_X1 port map( A1 => n18239, A2 => n22427, Z => n34468);
   U26104 : NAND2_X2 port map( A1 => n24624, A2 => n24734, ZN => n25196);
   U26107 : NAND2_X2 port map( A1 => n31712, A2 => n24769, ZN => n8406);
   U26113 : AOI21_X2 port map( A1 => n39092, A2 => n24083, B => n24082, ZN => 
                           n24735);
   U26119 : INV_X2 port map( I => n39094, ZN => n19153);
   U26121 : XOR2_X1 port map( A1 => n19154, A2 => n24633, Z => n39094);
   U26126 : NAND2_X2 port map( A1 => n39095, A2 => n2152, ZN => n26263);
   U26133 : NAND2_X2 port map( A1 => n39386, A2 => n26325, ZN => n39095);
   U26134 : BUF_X2 port map( I => n10379, Z => n39096);
   U26136 : INV_X2 port map( I => n39097, ZN => n14638);
   U26137 : XOR2_X1 port map( A1 => n10343, A2 => n28940, Z => n39097);
   U26139 : XOR2_X1 port map( A1 => n28978, A2 => n29081, Z => n2004);
   U26142 : XOR2_X1 port map( A1 => n29303, A2 => n14956, Z => n29836);
   U26144 : OAI21_X2 port map( A1 => n16920, A2 => n17007, B => n28757, ZN => 
                           n29303);
   U26146 : NAND2_X2 port map( A1 => n959, A2 => n33712, ZN => n18328);
   U26147 : NAND2_X2 port map( A1 => n19965, A2 => n19964, ZN => n25433);
   U26148 : AOI22_X2 port map( A1 => n24363, A2 => n38984, B1 => n36082, B2 => 
                           n39099, ZN => n24364);
   U26150 : XOR2_X1 port map( A1 => n8277, A2 => n8276, Z => n39100);
   U26154 : INV_X2 port map( I => n39073, ZN => n23914);
   U26158 : NOR2_X2 port map( A1 => n1270, A2 => n5282, ZN => n24775);
   U26164 : XOR2_X1 port map( A1 => n3885, A2 => n3886, Z => n28204);
   U26167 : XOR2_X1 port map( A1 => n13797, A2 => n39102, Z => n29312);
   U26168 : XOR2_X1 port map( A1 => n11346, A2 => n11922, Z => n39102);
   U26169 : XOR2_X1 port map( A1 => n23737, A2 => n14140, Z => n39103);
   U26174 : XOR2_X1 port map( A1 => n29058, A2 => n12244, Z => n29304);
   U26178 : NAND2_X2 port map( A1 => n28761, A2 => n19794, ZN => n29058);
   U26191 : XOR2_X1 port map( A1 => n10647, A2 => n10644, Z => n11402);
   U26195 : OAI21_X2 port map( A1 => n6293, A2 => n14915, B => n14914, ZN => 
                           n26055);
   U26197 : NAND2_X2 port map( A1 => n34613, A2 => n5672, ZN => n6293);
   U26202 : XOR2_X1 port map( A1 => n39105, A2 => n1322, Z => n34202);
   U26203 : XOR2_X1 port map( A1 => n22588, A2 => n22531, Z => n39105);
   U26205 : INV_X2 port map( I => n39106, ZN => n26988);
   U26209 : XNOR2_X1 port map( A1 => n13244, A2 => n7720, ZN => n39106);
   U26213 : NOR2_X1 port map( A1 => n23181, A2 => n22903, ZN => n39107);
   U26216 : XOR2_X1 port map( A1 => n26550, A2 => n26551, Z => n26601);
   U26218 : OAI21_X2 port map( A1 => n15552, A2 => n15551, B => n25784, ZN => 
                           n26551);
   U26221 : OAI22_X2 port map( A1 => n4991, A2 => n3598, B1 => n39761, B2 => 
                           n34667, ZN => n39189);
   U26224 : NAND2_X2 port map( A1 => n4492, A2 => n39109, ZN => n27690);
   U26226 : NAND3_X1 port map( A1 => n27070, A2 => n36989, A3 => n27071, ZN => 
                           n39109);
   U26227 : NAND2_X2 port map( A1 => n6844, A2 => n6845, ZN => n35654);
   U26234 : INV_X2 port map( I => n7023, ZN => n10544);
   U26235 : OAI21_X2 port map( A1 => n39150, A2 => n15986, B => n27235, ZN => 
                           n5994);
   U26239 : XOR2_X1 port map( A1 => n27778, A2 => n27746, Z => n27788);
   U26245 : OAI21_X2 port map( A1 => n5461, A2 => n5462, B => n39111, ZN => 
                           n20392);
   U26251 : XOR2_X1 port map( A1 => n27466, A2 => n32354, Z => n20846);
   U26254 : NAND2_X2 port map( A1 => n37163, A2 => n12814, ZN => n5408);
   U26260 : INV_X2 port map( I => n39113, ZN => n36361);
   U26267 : XOR2_X1 port map( A1 => Plaintext(139), A2 => Key(139), Z => n39113
                           );
   U26279 : XOR2_X1 port map( A1 => n15723, A2 => n39114, Z => n32932);
   U26282 : XOR2_X1 port map( A1 => n15721, A2 => n15722, Z => n39114);
   U26284 : XOR2_X1 port map( A1 => n33722, A2 => n39115, Z => n15692);
   U26285 : XOR2_X1 port map( A1 => n32135, A2 => n30169, Z => n22627);
   U26290 : AOI22_X2 port map( A1 => n4199, A2 => n35755, B1 => n4198, B2 => 
                           n31651, ZN => n32135);
   U26300 : BUF_X4 port map( I => n13686, Z => n39117);
   U26307 : NAND2_X2 port map( A1 => n28245, A2 => n28244, ZN => n28748);
   U26314 : XOR2_X1 port map( A1 => n484, A2 => n343, Z => n39118);
   U26332 : XOR2_X1 port map( A1 => n4079, A2 => n4080, Z => n39119);
   U26333 : OAI21_X2 port map( A1 => n2017, A2 => n2016, B => n2013, ZN => 
                           n31538);
   U26335 : NAND3_X2 port map( A1 => n10048, A2 => n14901, A3 => n11436, ZN => 
                           n34421);
   U26338 : NAND2_X2 port map( A1 => n8645, A2 => n8644, ZN => n8875);
   U26342 : NAND2_X2 port map( A1 => n12161, A2 => n39120, ZN => n25263);
   U26364 : XOR2_X1 port map( A1 => n39121, A2 => n18014, Z => n18017);
   U26371 : XOR2_X1 port map( A1 => n8240, A2 => n39544, Z => n39121);
   U26372 : BUF_X2 port map( I => n30183, Z => n39122);
   U26374 : INV_X2 port map( I => n39123, ZN => n8205);
   U26384 : XNOR2_X1 port map( A1 => n7115, A2 => n7112, ZN => n39123);
   U26385 : NAND2_X1 port map( A1 => n23247, A2 => n35232, ZN => n13578);
   U26388 : OAI22_X2 port map( A1 => n39124, A2 => n39714, B1 => n15633, B2 => 
                           n24910, ZN => n24994);
   U26402 : INV_X2 port map( I => n13843, ZN => n39124);
   U26413 : INV_X2 port map( I => n39125, ZN => n22962);
   U26419 : NOR2_X2 port map( A1 => n10047, A2 => n1046, ZN => n39125);
   U26425 : NAND2_X1 port map( A1 => n13105, A2 => n13104, ZN => n39170);
   U26427 : NAND2_X1 port map( A1 => n12694, A2 => n12505, ZN => n39128);
   U26434 : XOR2_X1 port map( A1 => n34414, A2 => n39130, Z => n35395);
   U26435 : XOR2_X1 port map( A1 => n2317, A2 => n25304, Z => n39130);
   U26440 : XOR2_X1 port map( A1 => n12999, A2 => n27773, Z => n27751);
   U26441 : BUF_X2 port map( I => n30574, Z => n39133);
   U26449 : NAND2_X2 port map( A1 => n24779, A2 => n24545, ZN => n24659);
   U26455 : OAI21_X2 port map( A1 => n16069, A2 => n18479, B => n16068, ZN => 
                           n24779);
   U26460 : XOR2_X1 port map( A1 => n39468, A2 => n25226, Z => n15316);
   U26462 : NOR2_X2 port map( A1 => n39134, A2 => n21196, ZN => n29341);
   U26463 : AOI22_X2 port map( A1 => n28510, A2 => n28509, B1 => n36414, B2 => 
                           n8218, ZN => n8217);
   U26476 : XOR2_X1 port map( A1 => n39135, A2 => n26262, Z => n13853);
   U26480 : AND2_X1 port map( A1 => n13278, A2 => n4272, Z => n39532);
   U26484 : NOR2_X2 port map( A1 => n8319, A2 => n24304, ZN => n12686);
   U26492 : XOR2_X1 port map( A1 => n39137, A2 => n6544, Z => n4997);
   U26499 : XOR2_X1 port map( A1 => n37149, A2 => n6546, Z => n39137);
   U26502 : NAND2_X2 port map( A1 => n39138, A2 => n34263, ZN => n3760);
   U26504 : NAND2_X1 port map( A1 => n39142, A2 => n31987, ZN => n39139);
   U26508 : NAND2_X2 port map( A1 => n21300, A2 => n33651, ZN => n14387);
   U26517 : XOR2_X1 port map( A1 => n11059, A2 => n39141, Z => n31125);
   U26519 : XOR2_X1 port map( A1 => n1506, A2 => n26511, Z => n11059);
   U26521 : AND2_X1 port map( A1 => n2001, A2 => n29956, Z => n32539);
   U26525 : OR2_X1 port map( A1 => n39140, A2 => n26055, Z => n13168);
   U26535 : NOR2_X2 port map( A1 => n20061, A2 => n39143, ZN => n20059);
   U26543 : XOR2_X1 port map( A1 => n3663, A2 => n35247, Z => n35246);
   U26546 : XOR2_X1 port map( A1 => n9719, A2 => n39136, Z => n39145);
   U26548 : NOR2_X2 port map( A1 => n10515, A2 => n10516, ZN => n39502);
   U26554 : INV_X4 port map( I => n4576, ZN => n7379);
   U26555 : OAI21_X2 port map( A1 => n7934, A2 => n8498, B => n35827, ZN => 
                           n7253);
   U26556 : INV_X2 port map( I => n39148, ZN => n7934);
   U26560 : NAND2_X2 port map( A1 => n2717, A2 => n2716, ZN => n39148);
   U26561 : XOR2_X1 port map( A1 => n39149, A2 => n33954, Z => n12673);
   U26563 : XOR2_X1 port map( A1 => n20820, A2 => n16549, Z => n39149);
   U26566 : XOR2_X1 port map( A1 => n22599, A2 => n22656, Z => n33177);
   U26567 : OAI21_X2 port map( A1 => n8028, A2 => n1047, B => n6032, ZN => 
                           n22656);
   U26570 : XOR2_X1 port map( A1 => n25247, A2 => n25175, Z => n25185);
   U26579 : NOR3_X1 port map( A1 => n12309, A2 => n18121, A3 => n13166, ZN => 
                           n31745);
   U26583 : NAND2_X2 port map( A1 => n29627, A2 => n29617, ZN => n29611);
   U26602 : AOI22_X1 port map( A1 => n6948, A2 => n9165, B1 => n10681, B2 => 
                           n4108, ZN => n39152);
   U26604 : NAND2_X2 port map( A1 => n1147, A2 => n5515, ZN => n30594);
   U26608 : NAND2_X2 port map( A1 => n23518, A2 => n19671, ZN => n20817);
   U26609 : NAND2_X2 port map( A1 => n6919, A2 => n37082, ZN => n8039);
   U26615 : NAND2_X2 port map( A1 => n39158, A2 => n19368, ZN => n26599);
   U26618 : OR2_X1 port map( A1 => n13686, A2 => n17034, Z => n32527);
   U26621 : XOR2_X1 port map( A1 => n39162, A2 => n17872, Z => n7319);
   U26623 : XOR2_X1 port map( A1 => n8884, A2 => n17874, Z => n39162);
   U26626 : XOR2_X1 port map( A1 => n26503, A2 => n26348, Z => n11620);
   U26627 : INV_X4 port map( I => n7542, ZN => n13294);
   U26631 : NAND2_X2 port map( A1 => n2493, A2 => n39164, ZN => n11247);
   U26638 : INV_X2 port map( I => n39166, ZN => n253);
   U26639 : XOR2_X1 port map( A1 => n10769, A2 => n10770, Z => n39166);
   U26643 : XOR2_X1 port map( A1 => n32685, A2 => n39167, Z => n34427);
   U26646 : XOR2_X1 port map( A1 => n25129, A2 => n25128, Z => n39167);
   U26651 : XOR2_X1 port map( A1 => n39168, A2 => n34955, Z => n20958);
   U26653 : XOR2_X1 port map( A1 => n22759, A2 => n20865, Z => n39168);
   U26654 : XOR2_X1 port map( A1 => n33870, A2 => n39169, Z => n19266);
   U26656 : XOR2_X1 port map( A1 => n14218, A2 => n1456, Z => n39169);
   U26657 : XOR2_X1 port map( A1 => n39170, A2 => n29221, Z => Ciphertext(9));
   U26658 : OAI21_X2 port map( A1 => n1034, A2 => n305, B => n38561, ZN => 
                           n34711);
   U26661 : INV_X2 port map( I => n39171, ZN => n9333);
   U26663 : NAND2_X2 port map( A1 => n37219, A2 => n39204, ZN => n4576);
   U26667 : AOI21_X2 port map( A1 => n19270, A2 => n554, B => n39173, ZN => 
                           n19268);
   U26673 : XOR2_X1 port map( A1 => n25010, A2 => n35339, Z => n31281);
   U26675 : INV_X2 port map( I => n39175, ZN => n7982);
   U26680 : XOR2_X1 port map( A1 => Plaintext(41), A2 => Key(41), Z => n39175);
   U26693 : AOI21_X2 port map( A1 => n34195, A2 => n4337, B => n4336, ZN => 
                           n4493);
   U26700 : XOR2_X1 port map( A1 => n15648, A2 => n9154, Z => n39177);
   U26708 : XOR2_X1 port map( A1 => n5381, A2 => n34722, Z => n5382);
   U26712 : BUF_X2 port map( I => n10429, Z => n9914);
   U26713 : NAND2_X2 port map( A1 => n4888, A2 => n25473, ZN => n35059);
   U26717 : XOR2_X1 port map( A1 => n13483, A2 => n8602, Z => n2161);
   U26718 : XOR2_X1 port map( A1 => n16054, A2 => n28850, Z => n8602);
   U26723 : NAND2_X2 port map( A1 => n35420, A2 => n32411, ZN => n28660);
   U26730 : OAI21_X2 port map( A1 => n24346, A2 => n7834, B => n1033, ZN => 
                           n7800);
   U26732 : NAND2_X1 port map( A1 => n3863, A2 => n22317, ZN => n22319);
   U26735 : XOR2_X1 port map( A1 => n36386, A2 => n27690, Z => n3258);
   U26742 : OAI21_X2 port map( A1 => n36099, A2 => n2534, B => n910, ZN => 
                           n2629);
   U26747 : NAND2_X2 port map( A1 => n39180, A2 => n28403, ZN => n31378);
   U26748 : NOR2_X1 port map( A1 => n902, A2 => n35777, ZN => n11094);
   U26750 : OAI21_X2 port map( A1 => n39181, A2 => n21564, B => n21562, ZN => 
                           n35431);
   U26754 : INV_X1 port map( I => n21560, ZN => n39181);
   U26763 : NAND2_X2 port map( A1 => n17792, A2 => n19543, ZN => n21560);
   U26768 : XOR2_X1 port map( A1 => n29121, A2 => n3280, Z => n11479);
   U26771 : AOI21_X2 port map( A1 => n13807, A2 => n28614, B => n13806, ZN => 
                           n3280);
   U26780 : XOR2_X1 port map( A1 => n36329, A2 => n15757, Z => n878);
   U26783 : AOI22_X2 port map( A1 => n6501, A2 => n26909, B1 => n1234, B2 => 
                           n26718, ZN => n35794);
   U26788 : NOR2_X1 port map( A1 => n26459, A2 => n20891, ZN => n26718);
   U26790 : NAND2_X2 port map( A1 => n2009, A2 => n12982, ZN => n11372);
   U26798 : NAND2_X2 port map( A1 => n39184, A2 => n31634, ZN => n17791);
   U26799 : NOR2_X2 port map( A1 => n18842, A2 => n37160, ZN => n39184);
   U26804 : XOR2_X1 port map( A1 => n39185, A2 => n3726, Z => n36338);
   U26807 : XOR2_X1 port map( A1 => n27673, A2 => n39186, Z => n39185);
   U26808 : NOR2_X1 port map( A1 => n13414, A2 => n12966, ZN => n2012);
   U26822 : NAND2_X2 port map( A1 => n18883, A2 => n36685, ZN => n28590);
   U26832 : XOR2_X1 port map( A1 => n6729, A2 => n6728, Z => n11145);
   U26840 : OR2_X1 port map( A1 => n28047, A2 => n39188, Z => n34340);
   U26849 : NAND2_X2 port map( A1 => n39189, A2 => n28592, ZN => n28865);
   U26852 : AND2_X1 port map( A1 => n4515, A2 => n32979, Z => n39781);
   U26854 : XOR2_X1 port map( A1 => n16755, A2 => n33182, Z => n35080);
   U26856 : OR2_X1 port map( A1 => n6945, A2 => n13370, Z => n10432);
   U26862 : NOR2_X2 port map( A1 => n18505, A2 => n22801, ZN => n6945);
   U26875 : NAND3_X2 port map( A1 => n24772, A2 => n24343, A3 => n3487, ZN => 
                           n11601);
   U26878 : NAND2_X2 port map( A1 => n25433, A2 => n7391, ZN => n15991);
   U26884 : AOI21_X1 port map( A1 => n14228, A2 => n951, B => n39015, ZN => 
                           n18464);
   U26886 : NAND2_X2 port map( A1 => n10836, A2 => n11048, ZN => n28051);
   U26887 : OAI21_X2 port map( A1 => n6807, A2 => n19211, B => n22262, ZN => 
                           n32081);
   U26891 : XOR2_X1 port map( A1 => n36305, A2 => n1969, Z => n24276);
   U26893 : XOR2_X1 port map( A1 => n39195, A2 => n24679, Z => n10309);
   U26894 : XOR2_X1 port map( A1 => n24676, A2 => n10199, Z => n39195);
   U26895 : BUF_X4 port map( I => n985, Z => n39235);
   U26902 : OAI21_X2 port map( A1 => n32260, A2 => n23569, B => n5792, ZN => 
                           n5791);
   U26910 : OR3_X1 port map( A1 => n21687, A2 => n7982, A3 => n21688, Z => 
                           n7965);
   U26913 : XOR2_X1 port map( A1 => n19112, A2 => n5802, Z => n3141);
   U26924 : XOR2_X1 port map( A1 => n20347, A2 => n25255, Z => n33759);
   U26925 : NAND2_X2 port map( A1 => n39197, A2 => n17062, ZN => n15069);
   U26927 : NAND2_X2 port map( A1 => n34268, A2 => n39415, ZN => n39197);
   U26929 : NOR2_X2 port map( A1 => n35917, A2 => n17388, ZN => n39770);
   U26930 : XOR2_X1 port map( A1 => n31348, A2 => n6456, Z => n32534);
   U26931 : INV_X1 port map( I => n2947, ZN => n999);
   U26939 : AOI21_X1 port map( A1 => n39405, A2 => n39406, B => n39317, ZN => 
                           n15553);
   U26946 : NAND2_X2 port map( A1 => n17806, A2 => n31650, ZN => n39317);
   U26954 : OAI21_X1 port map( A1 => n39261, A2 => n7387, B => n34373, ZN => 
                           n321);
   U26955 : AOI22_X2 port map( A1 => n39199, A2 => n23013, B1 => n39198, B2 => 
                           n1318, ZN => n23482);
   U26956 : OAI21_X2 port map( A1 => n16678, A2 => n5702, B => n33972, ZN => 
                           n39198);
   U26957 : NOR2_X2 port map( A1 => n32654, A2 => n31780, ZN => n20683);
   U26960 : XOR2_X1 port map( A1 => n26261, A2 => n26145, Z => n26146);
   U26961 : NAND2_X2 port map( A1 => n39200, A2 => n18309, ZN => n1414);
   U26970 : AND3_X1 port map( A1 => n28637, A2 => n39355, A3 => n33047, Z => 
                           n39366);
   U26972 : XOR2_X1 port map( A1 => n39201, A2 => n6780, Z => n24280);
   U26975 : NAND2_X1 port map( A1 => n29380, A2 => n14151, ZN => n28901);
   U26979 : NAND2_X2 port map( A1 => n1301, A2 => n35963, ZN => n20998);
   U26987 : OAI21_X2 port map( A1 => n39206, A2 => n39203, B => n27154, ZN => 
                           n3672);
   U26989 : NOR2_X2 port map( A1 => n22456, A2 => n39205, ZN => n39204);
   U26993 : XOR2_X1 port map( A1 => n27496, A2 => n27654, Z => n2042);
   U27000 : BUF_X2 port map( I => n27408, Z => n39206);
   U27005 : XOR2_X1 port map( A1 => n11740, A2 => n17657, Z => n39207);
   U27012 : INV_X2 port map( I => n18998, ZN => n9422);
   U27014 : NAND3_X2 port map( A1 => n7964, A2 => n7963, A3 => n7965, ZN => 
                           n18998);
   U27018 : XOR2_X1 port map( A1 => n39208, A2 => n29371, Z => Ciphertext(34));
   U27021 : OR2_X1 port map( A1 => n9604, A2 => n36361, Z => n15626);
   U27023 : XOR2_X1 port map( A1 => n1656, A2 => n22762, Z => n6224);
   U27026 : INV_X2 port map( I => n22228, ZN => n1331);
   U27034 : NOR2_X2 port map( A1 => n20423, A2 => n5935, ZN => n14921);
   U27037 : XOR2_X1 port map( A1 => n22750, A2 => n3172, Z => n2473);
   U27041 : XOR2_X1 port map( A1 => n22492, A2 => n22491, Z => n22750);
   U27042 : NAND2_X2 port map( A1 => n13066, A2 => n13068, ZN => n26357);
   U27043 : XOR2_X1 port map( A1 => n33807, A2 => n39210, Z => n34802);
   U27044 : XOR2_X1 port map( A1 => n61, A2 => n39211, Z => n39210);
   U27050 : INV_X2 port map( I => n31579, ZN => n39211);
   U27054 : XOR2_X1 port map( A1 => n39212, A2 => n15227, Z => n17604);
   U27055 : XOR2_X1 port map( A1 => n25200, A2 => n15226, Z => n39212);
   U27064 : INV_X2 port map( I => n39213, ZN => n34167);
   U27077 : NOR2_X2 port map( A1 => n27399, A2 => n12327, ZN => n39213);
   U27078 : OAI21_X2 port map( A1 => n15249, A2 => n28111, B => n15389, ZN => 
                           n20200);
   U27084 : NOR2_X2 port map( A1 => n8368, A2 => n4306, ZN => n15249);
   U27087 : NAND2_X2 port map( A1 => n12604, A2 => n19892, ZN => n11868);
   U27094 : NAND2_X2 port map( A1 => n2022, A2 => n3014, ZN => n19892);
   U27101 : XOR2_X1 port map( A1 => n17957, A2 => n29076, Z => n5129);
   U27102 : XOR2_X1 port map( A1 => n5130, A2 => n29082, Z => n29076);
   U27106 : AOI22_X2 port map( A1 => n11293, A2 => n37582, B1 => n11292, B2 => 
                           n7110, ZN => n17890);
   U27109 : NAND2_X1 port map( A1 => n17978, A2 => n28559, ZN => n17977);
   U27111 : XOR2_X1 port map( A1 => n38979, A2 => n26568, Z => n39685);
   U27118 : XOR2_X1 port map( A1 => n39217, A2 => n15421, Z => n14608);
   U27119 : XOR2_X1 port map( A1 => n36317, A2 => n27754, Z => n39217);
   U27120 : XOR2_X1 port map( A1 => n25243, A2 => n8163, Z => n25032);
   U27121 : INV_X2 port map( I => n30619, ZN => n29074);
   U27122 : XOR2_X1 port map( A1 => n28874, A2 => n39220, Z => n30619);
   U27123 : INV_X2 port map( I => n16309, ZN => n39220);
   U27124 : XOR2_X1 port map( A1 => n25217, A2 => n39221, Z => n25062);
   U27129 : XOR2_X1 port map( A1 => n25316, A2 => n19670, Z => n39221);
   U27130 : XOR2_X1 port map( A1 => n22443, A2 => n22527, Z => n7510);
   U27131 : INV_X4 port map( I => n31955, ZN => n27306);
   U27137 : NAND2_X1 port map( A1 => n1086, A2 => n35332, ZN => n15577);
   U27138 : NOR2_X2 port map( A1 => n35038, A2 => n34057, ZN => n31955);
   U27142 : AOI21_X2 port map( A1 => n15941, A2 => n37014, B => n1039, ZN => 
                           n15949);
   U27144 : INV_X2 port map( I => n5363, ZN => n39305);
   U27149 : NAND2_X2 port map( A1 => n39646, A2 => n15999, ZN => n5363);
   U27155 : NOR2_X2 port map( A1 => n5798, A2 => n14472, ZN => n39224);
   U27160 : NAND3_X2 port map( A1 => n12893, A2 => n9146, A3 => n9145, ZN => 
                           n10986);
   U27168 : XOR2_X1 port map( A1 => n8300, A2 => n8298, Z => n15873);
   U27169 : XOR2_X1 port map( A1 => n23781, A2 => n23878, Z => n6379);
   U27175 : NAND2_X2 port map( A1 => n39225, A2 => n37217, ZN => n39697);
   U27177 : NAND2_X2 port map( A1 => n11511, A2 => n29, ZN => n39225);
   U27178 : BUF_X2 port map( I => n25754, Z => n39226);
   U27180 : OR2_X1 port map( A1 => n9333, A2 => n37100, Z => n5335);
   U27195 : XOR2_X1 port map( A1 => n4612, A2 => n39228, Z => n7115);
   U27197 : XOR2_X1 port map( A1 => n39229, A2 => n38385, Z => n39228);
   U27204 : INV_X2 port map( I => n17937, ZN => n39229);
   U27210 : NOR2_X2 port map( A1 => n39230, A2 => n8763, ZN => n33563);
   U27215 : OR2_X1 port map( A1 => n9839, A2 => n31307, Z => n13839);
   U27221 : BUF_X2 port map( I => n36595, Z => n39231);
   U27223 : INV_X2 port map( I => n39232, ZN => n39817);
   U27229 : XOR2_X1 port map( A1 => n7929, A2 => n28925, Z => n39233);
   U27232 : XOR2_X1 port map( A1 => n8301, A2 => n8396, Z => n8395);
   U27237 : NAND2_X1 port map( A1 => n26098, A2 => n10764, ZN => n4990);
   U27246 : NOR2_X2 port map( A1 => n39236, A2 => n33376, ZN => n3071);
   U27251 : NAND2_X2 port map( A1 => n14737, A2 => n14735, ZN => n28594);
   U27252 : NAND2_X2 port map( A1 => n38220, A2 => n31664, ZN => n14735);
   U27254 : NAND2_X1 port map( A1 => n36530, A2 => n12289, ZN => n20421);
   U27255 : OAI21_X2 port map( A1 => n39237, A2 => n35290, B => n9265, ZN => 
                           n18872);
   U27266 : OAI21_X2 port map( A1 => n25845, A2 => n25844, B => n39238, ZN => 
                           n32106);
   U27283 : NAND3_X2 port map( A1 => n25842, A2 => n25954, A3 => n37966, ZN => 
                           n39238);
   U27284 : NAND2_X2 port map( A1 => n30833, A2 => n253, ZN => n24444);
   U27289 : XOR2_X1 port map( A1 => n12586, A2 => n36803, Z => n26919);
   U27292 : NOR2_X1 port map( A1 => n36361, A2 => n35455, ZN => n21780);
   U27293 : NAND2_X2 port map( A1 => n35362, A2 => n6424, ZN => n36226);
   U27297 : AOI22_X2 port map( A1 => n29349, A2 => n1062, B1 => n29348, B2 => 
                           n39240, ZN => n31307);
   U27298 : OR2_X1 port map( A1 => n807, A2 => n24266, Z => n11196);
   U27307 : NOR2_X1 port map( A1 => n29421, A2 => n32946, ZN => n12054);
   U27311 : INV_X2 port map( I => n39241, ZN => n5836);
   U27312 : XOR2_X1 port map( A1 => n8083, A2 => n35920, Z => n39241);
   U27314 : BUF_X2 port map( I => n33738, Z => n39242);
   U27317 : AOI21_X2 port map( A1 => n7986, A2 => n6064, B => n35962, ZN => 
                           n36450);
   U27321 : NOR2_X1 port map( A1 => n18601, A2 => n29338, ZN => n18671);
   U27327 : NAND2_X2 port map( A1 => n12060, A2 => n31810, ZN => n14858);
   U27329 : OAI21_X2 port map( A1 => n28287, A2 => n28288, B => n28161, ZN => 
                           n32077);
   U27335 : XOR2_X1 port map( A1 => n31240, A2 => n37222, Z => n16318);
   U27351 : XOR2_X1 port map( A1 => n24056, A2 => n24057, Z => n14821);
   U27352 : XOR2_X1 port map( A1 => n10722, A2 => n23794, Z => n24057);
   U27353 : OAI21_X2 port map( A1 => n39244, A2 => n39243, B => n3619, ZN => 
                           n19294);
   U27354 : OAI21_X1 port map( A1 => n9385, A2 => n24732, B => n35250, ZN => 
                           n3792);
   U27355 : OR2_X1 port map( A1 => n26688, A2 => n26665, Z => n18357);
   U27368 : NAND2_X2 port map( A1 => n34311, A2 => n113, ZN => n39484);
   U27375 : XOR2_X1 port map( A1 => n5225, A2 => n5226, Z => n20613);
   U27379 : NAND2_X2 port map( A1 => n23389, A2 => n4525, ZN => n23234);
   U27383 : XOR2_X1 port map( A1 => n30838, A2 => n39246, Z => n820);
   U27396 : XOR2_X1 port map( A1 => n25216, A2 => n25258, Z => n39246);
   U27407 : XOR2_X1 port map( A1 => n6681, A2 => n34351, Z => n31840);
   U27408 : XOR2_X1 port map( A1 => n11201, A2 => n22645, Z => n37023);
   U27411 : NAND2_X2 port map( A1 => n12567, A2 => n22162, ZN => n11201);
   U27418 : NOR2_X2 port map( A1 => n3685, A2 => n2336, ZN => n10065);
   U27419 : XOR2_X1 port map( A1 => n17326, A2 => n39247, Z => n29424);
   U27422 : OAI21_X2 port map( A1 => n25727, A2 => n16264, B => n39273, ZN => 
                           n10723);
   U27435 : OAI21_X1 port map( A1 => n31555, A2 => n26609, B => n39825, ZN => 
                           n34642);
   U27439 : XOR2_X1 port map( A1 => n25243, A2 => n29838, Z => n9325);
   U27444 : NAND3_X2 port map( A1 => n24766, A2 => n24767, A3 => n24768, ZN => 
                           n25243);
   U27445 : NOR2_X1 port map( A1 => n13524, A2 => n30283, ZN => n13523);
   U27448 : XOR2_X1 port map( A1 => n27665, A2 => n27835, Z => n18512);
   U27451 : INV_X1 port map( I => n35256, ZN => n39449);
   U27458 : XOR2_X1 port map( A1 => n10002, A2 => n27462, Z => n27985);
   U27463 : INV_X2 port map( I => n18257, ZN => n19716);
   U27466 : NAND2_X2 port map( A1 => n9569, A2 => n9570, ZN => n18257);
   U27480 : NAND2_X2 port map( A1 => n17917, A2 => n22891, ZN => n33163);
   U27481 : OAI22_X2 port map( A1 => n7537, A2 => n22920, B1 => n19945, B2 => 
                           n22682, ZN => n22891);
   U27484 : INV_X1 port map( I => n15459, ZN => n39252);
   U27489 : NAND2_X2 port map( A1 => n39253, A2 => n14895, ZN => n31986);
   U27492 : XOR2_X1 port map( A1 => n6571, A2 => n19816, Z => n6572);
   U27494 : NOR2_X2 port map( A1 => n4400, A2 => n4401, ZN => n6571);
   U27501 : NAND2_X2 port map( A1 => n17096, A2 => n19976, ZN => n4139);
   U27511 : OAI21_X2 port map( A1 => n19975, A2 => n17001, B => n39242, ZN => 
                           n17096);
   U27512 : XOR2_X1 port map( A1 => n39254, A2 => n34145, Z => n34351);
   U27523 : XOR2_X1 port map( A1 => n37593, A2 => n33308, Z => n39254);
   U27525 : NOR2_X2 port map( A1 => n6282, A2 => n2349, ZN => n25424);
   U27526 : NAND2_X2 port map( A1 => n24536, A2 => n19418, ZN => n25682);
   U27527 : OAI21_X2 port map( A1 => n24772, A2 => n24686, B => n5401, ZN => 
                           n39256);
   U27528 : AOI21_X2 port map( A1 => n20316, A2 => n38797, B => n39257, ZN => 
                           n16859);
   U27536 : XOR2_X1 port map( A1 => n7018, A2 => n26596, Z => n26261);
   U27546 : NAND2_X2 port map( A1 => n33517, A2 => n35568, ZN => n33030);
   U27550 : AOI22_X2 port map( A1 => n3949, A2 => n24467, B1 => n24466, B2 => 
                           n1280, ZN => n39354);
   U27554 : NOR2_X2 port map( A1 => n19566, A2 => n37259, ZN => n24466);
   U27558 : NOR2_X1 port map( A1 => n15299, A2 => n388, ZN => n4638);
   U27564 : OAI22_X2 port map( A1 => n22851, A2 => n22859, B1 => n5436, B2 => 
                           n383, ZN => n388);
   U27567 : INV_X4 port map( I => n33277, ZN => n39416);
   U27571 : XOR2_X1 port map( A1 => n17563, A2 => n638, Z => n2398);
   U27575 : XOR2_X1 port map( A1 => n35654, A2 => n26595, Z => n26358);
   U27578 : NOR2_X2 port map( A1 => n4460, A2 => n6178, ZN => n26595);
   U27580 : NOR2_X2 port map( A1 => n25661, A2 => n19153, ZN => n25383);
   U27583 : NAND2_X2 port map( A1 => n32929, A2 => n32928, ZN => n39260);
   U27585 : XOR2_X1 port map( A1 => n23712, A2 => n23893, Z => n23734);
   U27588 : NAND3_X2 port map( A1 => n23408, A2 => n23407, A3 => n23406, ZN => 
                           n23893);
   U27591 : BUF_X2 port map( I => n12617, Z => n39261);
   U27594 : INV_X2 port map( I => n33786, ZN => n1133);
   U27595 : NOR2_X2 port map( A1 => n36686, A2 => n31156, ZN => n36187);
   U27596 : XOR2_X1 port map( A1 => n12854, A2 => n12855, Z => n7865);
   U27599 : AND2_X1 port map( A1 => n24586, A2 => n10980, Z => n39505);
   U27608 : NOR2_X2 port map( A1 => n28626, A2 => n28625, ZN => n14712);
   U27624 : INV_X2 port map( I => n39263, ZN => n25498);
   U27626 : XOR2_X1 port map( A1 => n10153, A2 => n39694, Z => n12835);
   U27629 : XOR2_X1 port map( A1 => n6177, A2 => n7481, Z => n10153);
   U27632 : NAND2_X2 port map( A1 => n4823, A2 => n14848, ZN => n8493);
   U27634 : NAND2_X2 port map( A1 => n8160, A2 => n24233, ZN => n39370);
   U27640 : NAND2_X2 port map( A1 => n3869, A2 => n1609, ZN => n24233);
   U27651 : NOR2_X2 port map( A1 => n13988, A2 => n7236, ZN => n39264);
   U27653 : NOR2_X2 port map( A1 => n2832, A2 => n30656, ZN => n26591);
   U27654 : XOR2_X1 port map( A1 => n3893, A2 => n39267, Z => n3937);
   U27659 : XOR2_X1 port map( A1 => n11570, A2 => n1556, Z => n39267);
   U27667 : NAND2_X1 port map( A1 => n14587, A2 => n21391, ZN => n16289);
   U27672 : NAND2_X2 port map( A1 => n4001, A2 => n25361, ZN => n39269);
   U27686 : NOR2_X2 port map( A1 => n1676, A2 => n17207, ZN => n22136);
   U27691 : NAND3_X1 port map( A1 => n33747, A2 => n6235, A3 => n23574, ZN => 
                           n32927);
   U27692 : NAND3_X2 port map( A1 => n7825, A2 => n30631, A3 => n30276, ZN => 
                           n23970);
   U27693 : INV_X2 port map( I => n39270, ZN => n34073);
   U27694 : XOR2_X1 port map( A1 => n19015, A2 => n31849, Z => n39270);
   U27700 : XOR2_X1 port map( A1 => n208, A2 => n32441, Z => n17776);
   U27707 : XOR2_X1 port map( A1 => n25153, A2 => n21259, Z => n5629);
   U27713 : AOI22_X2 port map( A1 => n11159, A2 => n3803, B1 => n11160, B2 => 
                           n121, ZN => n39492);
   U27714 : XOR2_X1 port map( A1 => n34409, A2 => n27806, Z => n34408);
   U27725 : XOR2_X1 port map( A1 => n12411, A2 => n7726, Z => n32375);
   U27730 : XOR2_X1 port map( A1 => n39272, A2 => n27791, Z => n3157);
   U27734 : XOR2_X1 port map( A1 => n13448, A2 => n20659, Z => n39272);
   U27738 : XOR2_X1 port map( A1 => n13700, A2 => n2392, Z => n33582);
   U27741 : INV_X2 port map( I => n11601, ZN => n7350);
   U27750 : INV_X2 port map( I => n14193, ZN => n15737);
   U27752 : NAND2_X2 port map( A1 => n8845, A2 => n21211, ZN => n24683);
   U27759 : NAND2_X2 port map( A1 => n34577, A2 => n13717, ZN => n8858);
   U27761 : NAND2_X2 port map( A1 => n36693, A2 => n8863, ZN => n13717);
   U27763 : OR2_X1 port map( A1 => n33939, A2 => n13453, Z => n8847);
   U27768 : NOR2_X1 port map( A1 => n33516, A2 => n28272, ZN => n8308);
   U27771 : NAND3_X2 port map( A1 => n31358, A2 => n25467, A3 => n25469, ZN => 
                           n17329);
   U27773 : INV_X1 port map( I => n13554, ZN => n12387);
   U27775 : XOR2_X1 port map( A1 => n15348, A2 => n30626, Z => n15410);
   U27782 : XOR2_X1 port map( A1 => n24417, A2 => n9113, Z => n34347);
   U27783 : NAND3_X2 port map( A1 => n9416, A2 => n24493, A3 => n9418, ZN => 
                           n9113);
   U27788 : XOR2_X1 port map( A1 => n27817, A2 => n14325, Z => n27818);
   U27806 : OAI21_X2 port map( A1 => n18272, A2 => n18271, B => n6127, ZN => 
                           n39275);
   U27815 : XOR2_X1 port map( A1 => n28970, A2 => n34787, Z => n2218);
   U27818 : INV_X2 port map( I => n39277, ZN => n807);
   U27825 : XOR2_X1 port map( A1 => n39278, A2 => n1711, Z => Ciphertext(103));
   U27826 : BUF_X2 port map( I => n17412, Z => n39280);
   U27829 : NOR3_X2 port map( A1 => n39281, A2 => n32054, A3 => n34942, ZN => 
                           n16929);
   U27832 : XOR2_X1 port map( A1 => n25262, A2 => n39600, Z => n39282);
   U27833 : XOR2_X1 port map( A1 => n19374, A2 => n35468, Z => n3393);
   U27837 : INV_X2 port map( I => n39285, ZN => n5042);
   U27838 : NAND2_X1 port map( A1 => n39287, A2 => n39286, ZN => n5070);
   U27839 : NOR2_X1 port map( A1 => n9235, A2 => n20960, ZN => n39286);
   U27842 : XOR2_X1 port map( A1 => n35163, A2 => n39288, Z => n16110);
   U27849 : XOR2_X1 port map( A1 => n38385, A2 => n23957, Z => n39288);
   U27850 : BUF_X2 port map( I => n6145, Z => n39289);
   U27853 : AOI21_X2 port map( A1 => n12227, A2 => n28023, B => n27711, ZN => 
                           n27908);
   U27866 : XOR2_X1 port map( A1 => n35076, A2 => n5867, Z => n10251);
   U27874 : XOR2_X1 port map( A1 => n24047, A2 => n23969, Z => n23936);
   U27877 : NAND3_X2 port map( A1 => n31786, A2 => n1034, A3 => n24425, ZN => 
                           n39290);
   U27878 : OAI22_X2 port map( A1 => n39292, A2 => n39291, B1 => n2326, B2 => 
                           n1529, ZN => n33027);
   U27879 : INV_X2 port map( I => n35333, ZN => n39291);
   U27882 : INV_X2 port map( I => n26038, ZN => n39292);
   U27885 : NAND2_X2 port map( A1 => n39293, A2 => n30817, ZN => n15439);
   U27886 : NOR2_X2 port map( A1 => n14508, A2 => n15134, ZN => n39293);
   U27889 : NAND2_X1 port map( A1 => n39294, A2 => n24963, ZN => n4756);
   U27891 : XOR2_X1 port map( A1 => n19035, A2 => n16771, Z => n29119);
   U27893 : NAND3_X2 port map( A1 => n20878, A2 => n28410, A3 => n104, ZN => 
                           n19035);
   U27896 : NAND3_X2 port map( A1 => n23248, A2 => n12094, A3 => n23270, ZN => 
                           n39533);
   U27908 : BUF_X2 port map( I => n3977, Z => n39296);
   U27914 : XOR2_X1 port map( A1 => n23961, A2 => n8904, Z => n5179);
   U27915 : XOR2_X1 port map( A1 => n14393, A2 => n19835, Z => n19472);
   U27917 : NAND2_X2 port map( A1 => n7080, A2 => n14253, ZN => n14393);
   U27920 : OAI21_X2 port map( A1 => n36703, A2 => n20500, B => n2338, ZN => 
                           n28344);
   U27922 : INV_X2 port map( I => n253, ZN => n24440);
   U27923 : OAI21_X2 port map( A1 => n39301, A2 => n1133, B => n39299, ZN => 
                           n23377);
   U27924 : NOR2_X2 port map( A1 => n31157, A2 => n33952, ZN => n39302);
   U27925 : INV_X2 port map( I => n21144, ZN => n32712);
   U27928 : OAI22_X2 port map( A1 => n1076, A2 => n20010, B1 => n36197, B2 => 
                           n35469, ZN => n28281);
   U27930 : NAND2_X2 port map( A1 => n39414, A2 => n8262, ZN => n8261);
   U27941 : XOR2_X1 port map( A1 => n18049, A2 => n18048, Z => n20070);
   U27942 : INV_X2 port map( I => n3977, ZN => n35115);
   U27946 : NAND2_X2 port map( A1 => n35036, A2 => n4098, ZN => n3977);
   U27948 : XOR2_X1 port map( A1 => n28976, A2 => n28975, Z => n29907);
   U27960 : BUF_X2 port map( I => n10482, Z => n39303);
   U27968 : OAI21_X1 port map( A1 => n33369, A2 => n27385, B => n1471, ZN => 
                           n27384);
   U27971 : NAND2_X2 port map( A1 => n10693, A2 => n10689, ZN => n24529);
   U27972 : NAND2_X2 port map( A1 => n6027, A2 => n39304, ZN => n27672);
   U27975 : AOI22_X2 port map( A1 => n4610, A2 => n33336, B1 => n33369, B2 => 
                           n13222, ZN => n39304);
   U27981 : XOR2_X1 port map( A1 => n6905, A2 => n6906, Z => n19982);
   U27982 : NAND3_X1 port map( A1 => n31534, A2 => n29237, A3 => n14933, ZN => 
                           n39306);
   U28007 : NAND2_X2 port map( A1 => n39307, A2 => n13419, ZN => n32282);
   U28011 : OAI21_X2 port map( A1 => n3733, A2 => n7434, B => n2840, ZN => 
                           n39307);
   U28019 : NAND3_X1 port map( A1 => n781, A2 => n20173, A3 => n19594, ZN => 
                           n32283);
   U28020 : INV_X2 port map( I => n35246, ZN => n781);
   U28021 : INV_X2 port map( I => n39308, ZN => n29430);
   U28023 : OAI21_X2 port map( A1 => n15089, A2 => n14873, B => n36275, ZN => 
                           n39308);
   U28025 : INV_X2 port map( I => n20619, ZN => n24473);
   U28029 : NAND2_X1 port map( A1 => n39309, A2 => n20619, ZN => n4666);
   U28031 : XOR2_X1 port map( A1 => n20615, A2 => n23864, Z => n20619);
   U28033 : INV_X2 port map( I => n16816, ZN => n39309);
   U28040 : XOR2_X1 port map( A1 => n29111, A2 => n20727, Z => n16584);
   U28041 : XOR2_X1 port map( A1 => n8729, A2 => n29167, Z => n29111);
   U28051 : OAI21_X2 port map( A1 => n2731, A2 => n934, B => n24674, ZN => 
                           n31124);
   U28057 : OAI22_X2 port map( A1 => n36665, A2 => n31827, B1 => n1103, B2 => 
                           n26129, ZN => n5684);
   U28058 : NAND2_X2 port map( A1 => n5277, A2 => n12778, ZN => n25894);
   U28066 : XOR2_X1 port map( A1 => n36206, A2 => n17288, Z => n18830);
   U28072 : XOR2_X1 port map( A1 => n39311, A2 => n3304, Z => n13745);
   U28073 : XOR2_X1 port map( A1 => n3301, A2 => n3303, Z => n39311);
   U28083 : NAND2_X1 port map( A1 => n7300, A2 => n39485, ZN => n36526);
   U28092 : NOR2_X1 port map( A1 => n19992, A2 => n39312, ZN => n14432);
   U28100 : XOR2_X1 port map( A1 => n23780, A2 => n39314, Z => n39460);
   U28101 : AOI21_X2 port map( A1 => n13627, A2 => n34920, B => n13626, ZN => 
                           n5498);
   U28104 : XOR2_X1 port map( A1 => n25217, A2 => n39315, Z => n25220);
   U28106 : XOR2_X1 port map( A1 => n11267, A2 => n6051, Z => n6389);
   U28107 : AOI21_X2 port map( A1 => n4825, A2 => n9024, B => n7635, ZN => 
                           n39318);
   U28108 : BUF_X4 port map( I => n542, Z => n39739);
   U28110 : AND2_X1 port map( A1 => n892, A2 => n14405, Z => n31696);
   U28111 : XOR2_X1 port map( A1 => n16066, A2 => n27709, Z => n6395);
   U28112 : XOR2_X1 port map( A1 => n6033, A2 => n27787, Z => n27709);
   U28122 : XOR2_X1 port map( A1 => n22429, A2 => n18153, Z => n6369);
   U28123 : XOR2_X1 port map( A1 => n39319, A2 => n12853, Z => n33326);
   U28124 : XOR2_X1 port map( A1 => n21007, A2 => n33650, Z => n39319);
   U28125 : OR3_X1 port map( A1 => n39061, A2 => n25696, A3 => n20838, Z => 
                           n2495);
   U28126 : INV_X2 port map( I => n23571, ZN => n30524);
   U28127 : NOR2_X2 port map( A1 => n28771, A2 => n9290, ZN => n888);
   U28134 : OAI21_X2 port map( A1 => n5910, A2 => n37164, B => n34668, ZN => 
                           n9328);
   U28135 : INV_X2 port map( I => n39323, ZN => n18467);
   U28136 : XOR2_X1 port map( A1 => Plaintext(6), A2 => Key(6), Z => n39323);
   U28149 : NOR2_X2 port map( A1 => n11595, A2 => n11635, ZN => n11594);
   U28156 : NAND2_X1 port map( A1 => n24266, A2 => n24309, ZN => n39324);
   U28171 : NAND2_X1 port map( A1 => n11194, A2 => n24448, ZN => n39325);
   U28181 : XOR2_X1 port map( A1 => n18180, A2 => n34148, Z => n4918);
   U28182 : NAND2_X2 port map( A1 => n9140, A2 => n12152, ZN => n18180);
   U28219 : XOR2_X1 port map( A1 => n12014, A2 => n34214, Z => n26303);
   U28223 : XOR2_X1 port map( A1 => n12455, A2 => n12453, Z => n28550);
   U28224 : NAND2_X2 port map( A1 => n3844, A2 => n3843, ZN => n28473);
   U28234 : NAND2_X2 port map( A1 => n8157, A2 => n9585, ZN => n9035);
   U28244 : AOI22_X2 port map( A1 => n34585, A2 => n38724, B1 => n8046, B2 => 
                           n1630, ZN => n9246);
   U28256 : AND2_X2 port map( A1 => n16080, A2 => n7500, Z => n25427);
   U28266 : INV_X2 port map( I => n39326, ZN => n28093);
   U28281 : INV_X2 port map( I => n36634, ZN => n25053);
   U28284 : XOR2_X1 port map( A1 => n27758, A2 => n27647, Z => n27713);
   U28296 : OAI21_X2 port map( A1 => n39329, A2 => n10974, B => n26773, ZN => 
                           n39542);
   U28298 : NOR2_X2 port map( A1 => n26866, A2 => n1089, ZN => n39329);
   U28307 : OAI21_X2 port map( A1 => n39330, A2 => n21494, B => n21493, ZN => 
                           n22019);
   U28308 : OAI21_X2 port map( A1 => n35043, A2 => n21804, B => n35042, ZN => 
                           n39330);
   U28309 : XOR2_X1 port map( A1 => n27433, A2 => n34050, Z => n34650);
   U28314 : XOR2_X1 port map( A1 => n2515, A2 => n39331, Z => n30597);
   U28316 : XOR2_X1 port map( A1 => n26411, A2 => n37206, Z => n39331);
   U28317 : XOR2_X1 port map( A1 => n3665, A2 => n21056, Z => n21055);
   U28333 : XOR2_X1 port map( A1 => n16524, A2 => n23861, Z => n24055);
   U28334 : NAND3_X2 port map( A1 => n10123, A2 => n36903, A3 => n18499, ZN => 
                           n35331);
   U28337 : NOR2_X1 port map( A1 => n1186, A2 => n5424, ZN => n39334);
   U28351 : XOR2_X1 port map( A1 => n2041, A2 => n39335, Z => n35957);
   U28352 : INV_X1 port map( I => n39535, ZN => n28128);
   U28353 : AND2_X1 port map( A1 => n39535, A2 => n28093, Z => n8788);
   U28358 : INV_X1 port map( I => n39336, ZN => n36152);
   U28359 : NOR2_X2 port map( A1 => n34656, A2 => n3336, ZN => n34995);
   U28386 : OAI21_X1 port map( A1 => n39337, A2 => n29210, B => n30193, ZN => 
                           n16535);
   U28388 : NOR2_X1 port map( A1 => n17238, A2 => n35210, ZN => n39337);
   U28400 : AOI21_X2 port map( A1 => n12199, A2 => n38548, B => n37132, ZN => 
                           n3659);
   U28407 : BUF_X2 port map( I => n4034, Z => n39338);
   U28408 : INV_X2 port map( I => n39339, ZN => n640);
   U28409 : XOR2_X1 port map( A1 => n9687, A2 => n699, Z => n39339);
   U28410 : XNOR2_X1 port map( A1 => n23930, A2 => n24005, ZN => n39378);
   U28421 : XOR2_X1 port map( A1 => n18807, A2 => n19761, Z => n10083);
   U28445 : NOR2_X1 port map( A1 => n13926, A2 => n29566, ZN => n39340);
   U28463 : XOR2_X1 port map( A1 => n15973, A2 => n39341, Z => n23934);
   U28471 : XOR2_X1 port map( A1 => n15971, A2 => n15972, Z => n39341);
   U28474 : BUF_X2 port map( I => n14408, Z => n39342);
   U28476 : NOR2_X2 port map( A1 => n39343, A2 => n10019, ZN => n10193);
   U28488 : NOR2_X2 port map( A1 => n38166, A2 => n39345, ZN => n39379);
   U28489 : NOR2_X2 port map( A1 => n29444, A2 => n29595, ZN => n39345);
   U28493 : NAND2_X2 port map( A1 => n39616, A2 => n21529, ZN => n17861);
   U28522 : XOR2_X1 port map( A1 => n39346, A2 => n13288, Z => n13799);
   U28523 : XOR2_X1 port map( A1 => n29257, A2 => n13287, Z => n39346);
   U28526 : INV_X2 port map( I => n39347, ZN => n5976);
   U28531 : BUF_X2 port map( I => n32608, Z => n39348);
   U28536 : OAI22_X2 port map( A1 => n17716, A2 => n8711, B1 => n10062, B2 => 
                           n26030, ZN => n8708);
   U28538 : NAND2_X2 port map( A1 => n16407, A2 => n16867, ZN => n17716);
   U28539 : NAND2_X2 port map( A1 => n39349, A2 => n34257, ZN => n11729);
   U28556 : NOR2_X2 port map( A1 => n4656, A2 => n20549, ZN => n39349);
   U28561 : XOR2_X1 port map( A1 => n26384, A2 => n34648, Z => n19448);
   U28572 : OR2_X1 port map( A1 => n33455, A2 => n18741, Z => n13371);
   U28575 : XOR2_X1 port map( A1 => n26577, A2 => n36864, Z => n33455);
   U28576 : BUF_X2 port map( I => n4574, Z => n39350);
   U28577 : NOR2_X2 port map( A1 => n11364, A2 => n31383, ZN => n39808);
   U28582 : BUF_X2 port map( I => n950, Z => n39351);
   U28583 : NAND2_X2 port map( A1 => n34846, A2 => n39352, ZN => n10223);
   U28584 : NOR2_X1 port map( A1 => n15509, A2 => n939, ZN => n18278);
   U28592 : NOR2_X2 port map( A1 => n31751, A2 => n19706, ZN => n15509);
   U28600 : AND3_X1 port map( A1 => n28109, A2 => n8368, A3 => n33955, Z => 
                           n15391);
   U28601 : NAND2_X2 port map( A1 => n32469, A2 => n26108, ZN => n26107);
   U28602 : XOR2_X1 port map( A1 => n25010, A2 => n25011, Z => n18705);
   U28606 : XOR2_X1 port map( A1 => n25080, A2 => n35722, Z => n25010);
   U28612 : BUF_X2 port map( I => n6067, Z => n39355);
   U28616 : BUF_X2 port map( I => n22129, Z => n39356);
   U28630 : XOR2_X1 port map( A1 => n18498, A2 => n39358, Z => n8897);
   U28631 : XOR2_X1 port map( A1 => n35318, A2 => n39359, Z => n39358);
   U28632 : INV_X1 port map( I => n30120, ZN => n39359);
   U28634 : NAND2_X2 port map( A1 => n33438, A2 => n12080, ZN => n22401);
   U28638 : NAND2_X2 port map( A1 => n12776, A2 => n27099, ZN => n13703);
   U28640 : XOR2_X1 port map( A1 => n35445, A2 => n39360, Z => n31207);
   U28641 : XOR2_X1 port map( A1 => n660, A2 => n17988, Z => n39360);
   U28642 : XOR2_X1 port map( A1 => n27842, A2 => n1467, Z => n27469);
   U28645 : NAND2_X1 port map( A1 => n39126, A2 => n17114, ZN => n10721);
   U28648 : NAND2_X1 port map( A1 => n32294, A2 => n23610, ZN => n33356);
   U28652 : XOR2_X1 port map( A1 => n32765, A2 => n7990, Z => n24561);
   U28654 : AOI22_X2 port map( A1 => n10464, A2 => n919, B1 => n21836, B2 => 
                           n19620, ZN => n39361);
   U28655 : INV_X2 port map( I => n39362, ZN => n2393);
   U28679 : XOR2_X1 port map( A1 => n26363, A2 => n26184, Z => n17935);
   U28684 : XOR2_X1 port map( A1 => n39621, A2 => n20892, Z => n21301);
   U28688 : NOR2_X2 port map( A1 => n39367, A2 => n10354, ZN => n7243);
   U28693 : NOR2_X2 port map( A1 => n30282, A2 => n24691, ZN => n39367);
   U28697 : XOR2_X1 port map( A1 => n22712, A2 => n22564, Z => n5609);
   U28699 : NAND2_X2 port map( A1 => n6293, A2 => n32580, ZN => n7323);
   U28704 : OR2_X1 port map( A1 => n33249, A2 => n20694, Z => n21482);
   U28711 : XOR2_X1 port map( A1 => n9007, A2 => n39369, Z => n9338);
   U28726 : XOR2_X1 port map( A1 => n34901, A2 => n9005, Z => n39369);
   U28727 : OR2_X1 port map( A1 => n12447, A2 => n24328, Z => n20227);
   U28741 : NOR2_X2 port map( A1 => n21666, A2 => n21435, ZN => n21836);
   U28747 : NAND2_X2 port map( A1 => n34406, A2 => n34407, ZN => n34405);
   U28763 : NAND2_X2 port map( A1 => n32763, A2 => n10914, ZN => n33993);
   U28772 : NAND2_X2 port map( A1 => n39370, A2 => n23694, ZN => n423);
   U28784 : OAI21_X2 port map( A1 => n5621, A2 => n34030, B => n5380, ZN => 
                           n33461);
   U28786 : NAND2_X2 port map( A1 => n21478, A2 => n19388, ZN => n3618);
   U28788 : AOI21_X2 port map( A1 => n3620, A2 => n33240, B => n39372, ZN => 
                           n3619);
   U28793 : NOR2_X2 port map( A1 => n39373, A2 => n39381, ZN => n39372);
   U28799 : NAND2_X2 port map( A1 => n33579, A2 => n37107, ZN => n39381);
   U28800 : AND2_X1 port map( A1 => n894, A2 => n39374, Z => n36469);
   U28801 : NAND3_X1 port map( A1 => n1404, A2 => n29596, A3 => n14417, ZN => 
                           n39374);
   U28811 : NAND2_X2 port map( A1 => n1006, A2 => n924, ZN => n7596);
   U28814 : AOI21_X2 port map( A1 => n39377, A2 => n39376, B => n20357, ZN => 
                           n13922);
   U28815 : NAND2_X2 port map( A1 => n4388, A2 => n19778, ZN => n39376);
   U28819 : OAI21_X2 port map( A1 => n2410, A2 => n14417, B => n39379, ZN => 
                           n29475);
   U28820 : NAND2_X1 port map( A1 => n24963, A2 => n1530, ZN => n39380);
   U28821 : NAND2_X2 port map( A1 => n28478, A2 => n1196, ZN => n28370);
   U28826 : NAND2_X2 port map( A1 => n3533, A2 => n3534, ZN => n28478);
   U28829 : NAND2_X2 port map( A1 => n24261, A2 => n39381, ZN => n24263);
   U28833 : XOR2_X1 port map( A1 => n39383, A2 => n15700, Z => Ciphertext(169))
                           ;
   U28842 : AOI22_X1 port map( A1 => n29015, A2 => n18424, B1 => n30139, B2 => 
                           n30146, ZN => n39383);
   U28852 : AOI22_X2 port map( A1 => n27348, A2 => n33146, B1 => n27351, B2 => 
                           n27350, ZN => n10366);
   U28853 : NOR2_X1 port map( A1 => n8798, A2 => n8988, ZN => n27348);
   U28857 : XOR2_X1 port map( A1 => n39384, A2 => n28782, Z => n36514);
   U28859 : XOR2_X1 port map( A1 => n28780, A2 => n32465, Z => n39384);
   U28860 : NOR2_X2 port map( A1 => n26737, A2 => n17024, ZN => n17023);
   U28863 : XOR2_X1 port map( A1 => n25237, A2 => n25179, Z => n25188);
   U28870 : XOR2_X1 port map( A1 => n39385, A2 => n36456, Z => n34828);
   U28885 : XOR2_X1 port map( A1 => n39651, A2 => n19025, Z => n39385);
   U28887 : NAND2_X2 port map( A1 => n31048, A2 => n12936, ZN => n39583);
   U28893 : NOR3_X2 port map( A1 => n8803, A2 => n8804, A3 => n24794, ZN => 
                           n32019);
   U28894 : NAND2_X2 port map( A1 => n11614, A2 => n8944, ZN => n28505);
   U28895 : INV_X1 port map( I => n26325, ZN => n1237);
   U28896 : NOR2_X2 port map( A1 => n20851, A2 => n20852, ZN => n26325);
   U28897 : NAND2_X2 port map( A1 => n39387, A2 => n31180, ZN => n16260);
   U28907 : OAI21_X2 port map( A1 => n29383, A2 => n17444, B => n29382, ZN => 
                           n39387);
   U28908 : XOR2_X1 port map( A1 => n13852, A2 => n8939, Z => n17250);
   U28913 : NAND2_X2 port map( A1 => n34781, A2 => n8934, ZN => n8939);
   U28914 : NAND2_X2 port map( A1 => n39388, A2 => n4028, ZN => n28622);
   U28928 : OAI21_X2 port map( A1 => n14378, A2 => n17711, B => n24180, ZN => 
                           n364);
   U28937 : NAND2_X2 port map( A1 => n14378, A2 => n24142, ZN => n24180);
   U28945 : XOR2_X1 port map( A1 => n29296, A2 => n28610, Z => n29140);
   U28946 : NAND2_X2 port map( A1 => n20314, A2 => n28331, ZN => n29296);
   U28947 : OAI21_X2 port map( A1 => n1095, A2 => n1094, B => n1787, ZN => 
                           n26728);
   U28948 : XOR2_X1 port map( A1 => n17569, A2 => n30409, Z => n15118);
   U28958 : XOR2_X1 port map( A1 => n22453, A2 => n9116, Z => n17569);
   U28974 : NAND2_X2 port map( A1 => n31795, A2 => n26887, ZN => n27703);
   U28989 : XOR2_X1 port map( A1 => n21268, A2 => n182, Z => n24224);
   U28990 : NAND2_X2 port map( A1 => n33209, A2 => n33328, ZN => n1010);
   U28997 : NAND2_X2 port map( A1 => n8659, A2 => n14237, ZN => n39391);
   U29001 : AOI21_X2 port map( A1 => n36777, A2 => n7905, B => n39394, ZN => 
                           n34751);
   U29034 : INV_X2 port map( I => n14735, ZN => n39394);
   U29035 : OR2_X1 port map( A1 => n24432, A2 => n19576, Z => n20458);
   U29044 : XOR2_X1 port map( A1 => n359, A2 => n22476, Z => n22754);
   U29055 : XOR2_X1 port map( A1 => n39395, A2 => n33320, Z => Ciphertext(66));
   U29064 : AOI22_X1 port map( A1 => n31284, A2 => n29570, B1 => n13442, B2 => 
                           n20701, ZN => n39395);
   U29065 : NAND2_X2 port map( A1 => n39396, A2 => n16737, ZN => n7317);
   U29079 : OAI21_X2 port map( A1 => n14625, A2 => n16739, B => n31780, ZN => 
                           n39396);
   U29085 : BUF_X2 port map( I => n28114, Z => n39399);
   U29089 : OR2_X2 port map( A1 => n19821, A2 => n19423, Z => n39824);
   U29090 : INV_X2 port map( I => n39400, ZN => n14103);
   U29093 : NOR2_X2 port map( A1 => n5427, A2 => n1198, ZN => n39400);
   U29094 : XOR2_X1 port map( A1 => n11479, A2 => n29002, Z => n16601);
   U29096 : XOR2_X1 port map( A1 => n28971, A2 => n28896, Z => n29002);
   U29097 : XOR2_X1 port map( A1 => n31215, A2 => n14802, Z => n20171);
   U29103 : XOR2_X1 port map( A1 => n26572, A2 => n39032, Z => n14802);
   U29108 : AOI21_X2 port map( A1 => n34484, A2 => n11421, B => n35988, ZN => 
                           n614);
   U29116 : OAI22_X2 port map( A1 => n4808, A2 => n16686, B1 => n26824, B2 => 
                           n14488, ZN => n35988);
   U29117 : INV_X2 port map( I => n39403, ZN => n39811);
   U29118 : XOR2_X1 port map( A1 => n11498, A2 => n7341, Z => n39403);
   U29120 : NAND2_X2 port map( A1 => n19914, A2 => n1006, ZN => n14807);
   U29121 : INV_X2 port map( I => n39404, ZN => n24140);
   U29124 : XNOR2_X1 port map( A1 => n35481, A2 => n35480, ZN => n39404);
   U29125 : INV_X2 port map( I => n24879, ZN => n39405);
   U29126 : BUF_X2 port map( I => n9231, Z => n39407);
   U29133 : AND2_X1 port map( A1 => n15566, A2 => n34764, Z => n9293);
   U29136 : XOR2_X1 port map( A1 => n25232, A2 => n21154, Z => n2662);
   U29140 : XOR2_X1 port map( A1 => n28955, A2 => n39409, Z => n33890);
   U29142 : XOR2_X1 port map( A1 => n28951, A2 => n37254, Z => n39409);
   U29145 : XOR2_X1 port map( A1 => n32647, A2 => n39780, Z => n28130);
   U29147 : INV_X1 port map( I => n27728, ZN => n39410);
   U29153 : XOR2_X1 port map( A1 => n17417, A2 => n27779, Z => n27728);
   U29167 : OAI21_X2 port map( A1 => n26053, A2 => n34153, B => n33395, ZN => 
                           n1760);
   U29173 : INV_X2 port map( I => n39411, ZN => n21767);
   U29174 : XNOR2_X1 port map( A1 => Plaintext(132), A2 => Key(132), ZN => 
                           n39411);
   U29175 : NAND2_X2 port map( A1 => n3744, A2 => n3745, ZN => n23938);
   U29183 : XOR2_X1 port map( A1 => n8894, A2 => n27758, Z => n10539);
   U29198 : XOR2_X1 port map( A1 => n36706, A2 => n15393, Z => n17726);
   U29199 : XOR2_X1 port map( A1 => n31535, A2 => n27470, Z => n27715);
   U29202 : AOI22_X2 port map( A1 => n33278, A2 => n33277, B1 => n33276, B2 => 
                           n1400, ZN => n39734);
   U29207 : NOR2_X1 port map( A1 => n22068, A2 => n32318, ZN => n39801);
   U29227 : NAND3_X2 port map( A1 => n17236, A2 => n28052, A3 => n10443, ZN => 
                           n17234);
   U29237 : XOR2_X1 port map( A1 => n7069, A2 => n27662, Z => n7068);
   U29239 : NAND2_X2 port map( A1 => n33563, A2 => n21164, ZN => n27662);
   U29241 : NAND2_X2 port map( A1 => n34866, A2 => n1436, ZN => n39419);
   U29251 : NOR2_X2 port map( A1 => n21114, A2 => n8840, ZN => n24737);
   U29255 : AOI21_X2 port map( A1 => n24217, A2 => n24218, B => n20839, ZN => 
                           n21114);
   U29263 : NAND2_X2 port map( A1 => n28435, A2 => n8321, ZN => n35320);
   U29264 : NOR2_X2 port map( A1 => n3634, A2 => n31036, ZN => n36595);
   U29265 : XOR2_X1 port map( A1 => n28940, A2 => n29818, Z => n29168);
   U29266 : NOR2_X2 port map( A1 => n31608, A2 => n16503, ZN => n28940);
   U29269 : NAND2_X1 port map( A1 => n34476, A2 => n39421, ZN => n30512);
   U29271 : AOI22_X1 port map( A1 => n30070, A2 => n30076, B1 => n3815, B2 => 
                           n6687, ZN => n39421);
   U29272 : NOR2_X1 port map( A1 => n3927, A2 => n6405, ZN => n39422);
   U29273 : OR2_X1 port map( A1 => n39769, A2 => n29059, Z => n39432);
   U29277 : OR2_X1 port map( A1 => n2798, A2 => n39401, Z => n16842);
   U29279 : XOR2_X1 port map( A1 => n4438, A2 => n39427, Z => n5975);
   U29281 : XOR2_X1 port map( A1 => n28839, A2 => n28838, Z => n2547);
   U29282 : XOR2_X1 port map( A1 => n16357, A2 => n29828, Z => n28839);
   U29283 : OAI21_X2 port map( A1 => n2453, A2 => n2454, B => n39428, ZN => 
                           n14272);
   U29284 : AOI22_X2 port map( A1 => n34073, A2 => n14390, B1 => n19823, B2 => 
                           n17464, ZN => n23154);
   U29285 : XOR2_X1 port map( A1 => n26555, A2 => n39429, Z => n157);
   U29290 : XOR2_X1 port map( A1 => n26194, A2 => n8002, Z => n39429);
   U29292 : NAND3_X1 port map( A1 => n13876, A2 => n876, A3 => n27970, ZN => 
                           n13875);
   U29293 : OAI21_X2 port map( A1 => n26353, A2 => n17786, B => n20190, ZN => 
                           n4272);
   U29303 : OAI21_X2 port map( A1 => n27587, A2 => n27306, B => n4781, ZN => 
                           n27040);
   U29305 : OR2_X2 port map( A1 => n8000, A2 => n21152, Z => n8311);
   U29307 : XOR2_X1 port map( A1 => n24575, A2 => n13190, Z => n31075);
   U29315 : NOR2_X1 port map( A1 => n32981, A2 => n36454, ZN => n15033);
   U29317 : XOR2_X1 port map( A1 => n39430, A2 => n33674, Z => n8454);
   U29323 : XOR2_X1 port map( A1 => n29836, A2 => n39490, Z => n39430);
   U29324 : NAND2_X1 port map( A1 => n2866, A2 => n12081, ZN => n39431);
   U29328 : INV_X2 port map( I => n39433, ZN => n8042);
   U29329 : NAND2_X2 port map( A1 => n6601, A2 => n6599, ZN => n2792);
   U29337 : NOR2_X2 port map( A1 => n29559, A2 => n6252, ZN => n29551);
   U29342 : NOR2_X1 port map( A1 => n39435, A2 => n12527, ZN => n10992);
   U29343 : NOR2_X1 port map( A1 => n39436, A2 => n29012, ZN => n36013);
   U29345 : NOR2_X2 port map( A1 => n14833, A2 => n5450, ZN => n21449);
   U29348 : NAND2_X2 port map( A1 => n5449, A2 => n5448, ZN => n5450);
   U29352 : XOR2_X1 port map( A1 => n6596, A2 => n39437, Z => n6657);
   U29353 : XOR2_X1 port map( A1 => n25200, A2 => n37234, Z => n39437);
   U29359 : XOR2_X1 port map( A1 => n39438, A2 => n26309, Z => n13528);
   U29372 : XOR2_X1 port map( A1 => n12933, A2 => n12429, Z => n39438);
   U29376 : NAND2_X2 port map( A1 => n38881, A2 => n17960, ZN => n17959);
   U29379 : XOR2_X1 port map( A1 => n12181, A2 => n12180, Z => n12179);
   U29381 : NAND2_X2 port map( A1 => n6926, A2 => n32778, ZN => n9668);
   U29391 : OAI22_X2 port map( A1 => n39439, A2 => n36207, B1 => n36225, B2 => 
                           n16672, ZN => n31453);
   U29397 : AOI22_X2 port map( A1 => n34389, A2 => n30196, B1 => n1755, B2 => 
                           n33861, ZN => n39439);
   U29399 : XOR2_X1 port map( A1 => n382, A2 => n25252, Z => n10616);
   U29402 : OAI22_X2 port map( A1 => n24731, A2 => n11712, B1 => n24730, B2 => 
                           n39157, ZN => n382);
   U29404 : OAI21_X2 port map( A1 => n39441, A2 => n39440, B => n14331, ZN => 
                           n15953);
   U29419 : INV_X2 port map( I => n23200, ZN => n39440);
   U29426 : NAND2_X2 port map( A1 => n11183, A2 => n11185, ZN => n23814);
   U29434 : INV_X2 port map( I => n39444, ZN => n25434);
   U29437 : XNOR2_X1 port map( A1 => n25220, A2 => n39657, ZN => n39444);
   U29439 : XOR2_X1 port map( A1 => Plaintext(80), A2 => Key(80), Z => n39680);
   U29447 : XOR2_X1 port map( A1 => n10301, A2 => n38213, Z => n27601);
   U29454 : NAND2_X2 port map( A1 => n26648, A2 => n36953, ZN => n27689);
   U29455 : OAI21_X1 port map( A1 => n29358, A2 => n7376, B => n29372, ZN => 
                           n13646);
   U29467 : OAI21_X2 port map( A1 => n14311, A2 => n8089, B => n39445, ZN => 
                           n13766);
   U29468 : INV_X2 port map( I => n22133, ZN => n39445);
   U29488 : OAI22_X2 port map( A1 => n9252, A2 => n22131, B1 => n31573, B2 => 
                           n35780, ZN => n22133);
   U29497 : INV_X2 port map( I => n39446, ZN => n8197);
   U29502 : XNOR2_X1 port map( A1 => n7037, A2 => n7040, ZN => n39446);
   U29503 : XOR2_X1 port map( A1 => n9187, A2 => n14902, Z => n39447);
   U29504 : NOR2_X2 port map( A1 => n18536, A2 => n18537, ZN => n24857);
   U29510 : NOR2_X2 port map( A1 => n1420, A2 => n9668, ZN => n4531);
   U29513 : AND2_X1 port map( A1 => n39449, A2 => n26863, Z => n14732);
   U29515 : NOR2_X1 port map( A1 => n4633, A2 => n34987, ZN => n10634);
   U29521 : XOR2_X1 port map( A1 => n39450, A2 => n34092, Z => n10835);
   U29526 : XOR2_X1 port map( A1 => n33505, A2 => n15405, Z => n39450);
   U29534 : OAI21_X2 port map( A1 => n14125, A2 => n39451, B => n6295, ZN => 
                           n2696);
   U29535 : AND2_X1 port map( A1 => n5751, A2 => n14124, Z => n39451);
   U29536 : NOR2_X2 port map( A1 => n31948, A2 => n39452, ZN => n32601);
   U29542 : NOR3_X1 port map( A1 => n22792, A2 => n33925, A3 => n33544, ZN => 
                           n39452);
   U29547 : XOR2_X1 port map( A1 => n21227, A2 => n32383, Z => n32382);
   U29549 : XOR2_X1 port map( A1 => n11383, A2 => n3448, Z => n21227);
   U29550 : NOR2_X1 port map( A1 => n34286, A2 => n34285, ZN => n39453);
   U29559 : NAND2_X2 port map( A1 => n33987, A2 => n34526, ZN => n6791);
   U29563 : INV_X1 port map( I => n26290, ZN => n34009);
   U29569 : XNOR2_X1 port map( A1 => n26381, A2 => n26290, ZN => n32175);
   U29572 : NAND2_X2 port map( A1 => n4189, A2 => n25891, ZN => n26290);
   U29580 : OAI21_X1 port map( A1 => n39602, A2 => n30989, B => n33455, ZN => 
                           n26578);
   U29582 : INV_X2 port map( I => n39455, ZN => n2707);
   U29589 : XOR2_X1 port map( A1 => n21035, A2 => n35626, Z => n39456);
   U29590 : NAND3_X2 port map( A1 => n17811, A2 => n19069, A3 => n33101, ZN => 
                           n31650);
   U29591 : NAND2_X2 port map( A1 => n39457, A2 => n6463, ZN => n23707);
   U29592 : NAND2_X1 port map( A1 => n18618, A2 => n34012, ZN => n39457);
   U29597 : NAND3_X1 port map( A1 => n23172, A2 => n39418, A3 => n38752, ZN => 
                           n20176);
   U29603 : OAI21_X2 port map( A1 => n39599, A2 => n6731, B => n25637, ZN => 
                           n39458);
   U29604 : XOR2_X1 port map( A1 => n39459, A2 => n20270, Z => n20394);
   U29605 : XOR2_X1 port map( A1 => n39460, A2 => n24074, Z => n39459);
   U29609 : NAND2_X2 port map( A1 => n39461, A2 => n39338, ZN => n7);
   U29612 : NAND2_X2 port map( A1 => n27300, A2 => n4033, ZN => n39461);
   U29613 : XOR2_X1 port map( A1 => n27751, A2 => n39462, Z => n19009);
   U29614 : XOR2_X1 port map( A1 => n9013, A2 => n35464, Z => n39462);
   U29617 : NAND3_X2 port map( A1 => n4439, A2 => n13982, A3 => n23509, ZN => 
                           n11669);
   U29621 : NOR2_X2 port map( A1 => n3659, A2 => n30934, ZN => n13155);
   U29625 : INV_X2 port map( I => n39463, ZN => n37052);
   U29628 : XNOR2_X1 port map( A1 => n6924, A2 => n6922, ZN => n39463);
   U29629 : NAND2_X2 port map( A1 => n39517, A2 => n26778, ZN => n2947);
   U29636 : OAI21_X2 port map( A1 => n22683, A2 => n8339, B => n17568, ZN => 
                           n39464);
   U29638 : XOR2_X1 port map( A1 => n35218, A2 => n8402, Z => n39465);
   U29640 : NAND2_X2 port map( A1 => n39466, A2 => n9504, ZN => n12289);
   U29643 : NAND2_X1 port map( A1 => n9506, A2 => n19769, ZN => n39466);
   U29644 : XOR2_X1 port map( A1 => n24942, A2 => n5845, Z => n15531);
   U29645 : AOI21_X2 port map( A1 => n37208, A2 => n23225, B => n15074, ZN => 
                           n15073);
   U29648 : XOR2_X1 port map( A1 => n16368, A2 => n17462, Z => n9122);
   U29665 : NAND2_X2 port map( A1 => n7725, A2 => n9178, ZN => n39514);
   U29672 : OAI22_X2 port map( A1 => n19134, A2 => n32228, B1 => n11295, B2 => 
                           n23124, ZN => n14343);
   U29680 : INV_X2 port map( I => n20897, ZN => n32228);
   U29681 : XOR2_X1 port map( A1 => n11382, A2 => n32847, Z => n20897);
   U29686 : NAND2_X2 port map( A1 => n2193, A2 => n8570, ZN => n9116);
   U29687 : NOR2_X2 port map( A1 => n36507, A2 => n26372, ZN => n27389);
   U29691 : INV_X2 port map( I => n35164, ZN => n18619);
   U29692 : NAND2_X1 port map( A1 => n39467, A2 => n24395, ZN => n24181);
   U29701 : INV_X2 port map( I => n8760, ZN => n39467);
   U29703 : NAND2_X2 port map( A1 => n24716, A2 => n14534, ZN => n25226);
   U29705 : NOR3_X1 port map( A1 => n20418, A2 => n23399, A3 => n36810, ZN => 
                           n23320);
   U29706 : XOR2_X1 port map( A1 => n39809, A2 => n36190, Z => n22968);
   U29708 : NOR3_X2 port map( A1 => n840, A2 => n949, A3 => n9743, ZN => n33433
                           );
   U29710 : AOI21_X2 port map( A1 => n34720, A2 => n37477, B => n31796, ZN => 
                           n39469);
   U29713 : OR2_X2 port map( A1 => n5104, A2 => n39470, Z => n34475);
   U29714 : OAI22_X1 port map( A1 => n21519, A2 => n19397, B1 => n21520, B2 => 
                           n21521, ZN => n39470);
   U29725 : XOR2_X1 port map( A1 => n15776, A2 => n27703, Z => n27500);
   U29733 : XOR2_X1 port map( A1 => n39471, A2 => n1051, Z => Ciphertext(161));
   U29741 : AOI22_X1 port map( A1 => n30107, A2 => n12204, B1 => n18483, B2 => 
                           n16180, ZN => n39471);
   U29750 : XNOR2_X1 port map( A1 => n26356, A2 => n9151, ZN => n6477);
   U29752 : INV_X2 port map( I => n39472, ZN => n17692);
   U29754 : XOR2_X1 port map( A1 => n39474, A2 => n7180, Z => n20649);
   U29755 : XOR2_X1 port map( A1 => n28984, A2 => n7182, Z => n39474);
   U29761 : NAND2_X2 port map( A1 => n11889, A2 => n20859, ZN => n36798);
   U29763 : XOR2_X1 port map( A1 => n39475, A2 => n16601, Z => n16599);
   U29767 : XOR2_X1 port map( A1 => n33387, A2 => n14487, Z => n39475);
   U29769 : NAND3_X2 port map( A1 => n23248, A2 => n22852, A3 => n23270, ZN => 
                           n15491);
   U29772 : XOR2_X1 port map( A1 => n39476, A2 => n16679, Z => n6165);
   U29775 : XOR2_X1 port map( A1 => n2585, A2 => n34188, Z => n39476);
   U29778 : NAND2_X2 port map( A1 => n3120, A2 => n24637, ZN => n24635);
   U29796 : OAI21_X2 port map( A1 => n15496, A2 => n15497, B => n24230, ZN => 
                           n24637);
   U29811 : NAND2_X1 port map( A1 => n36474, A2 => n29124, ZN => n36473);
   U29819 : XOR2_X1 port map( A1 => n30687, A2 => n13205, Z => n36552);
   U29823 : INV_X4 port map( I => n7852, ZN => n24691);
   U29834 : INV_X2 port map( I => n30989, ZN => n39477);
   U29839 : BUF_X2 port map( I => n14379, Z => n39478);
   U29845 : INV_X2 port map( I => n39479, ZN => n39830);
   U29846 : XOR2_X1 port map( A1 => n36127, A2 => n28320, Z => n39479);
   U29847 : XOR2_X1 port map( A1 => n9085, A2 => n26480, Z => n26572);
   U29851 : AOI21_X2 port map( A1 => n8709, A2 => n8711, B => n8708, ZN => 
                           n9085);
   U29866 : NAND2_X2 port map( A1 => n32596, A2 => n39481, ZN => n18300);
   U29869 : OR2_X2 port map( A1 => n7631, A2 => n23380, Z => n30364);
   U29870 : OAI21_X2 port map( A1 => n39711, A2 => n20981, B => n4716, ZN => 
                           n14115);
   U29872 : NOR2_X2 port map( A1 => n26152, A2 => n26153, ZN => n27164);
   U29874 : XOR2_X1 port map( A1 => n31807, A2 => n27178, Z => n1859);
   U29876 : NAND2_X2 port map( A1 => n27165, A2 => n21272, ZN => n27387);
   U29879 : NAND2_X2 port map( A1 => n26445, A2 => n26446, ZN => n27165);
   U29884 : NAND2_X1 port map( A1 => n39483, A2 => n39482, ZN => n10556);
   U29885 : NAND2_X1 port map( A1 => n12661, A2 => n12660, ZN => n39483);
   U29890 : NAND2_X1 port map( A1 => n5976, A2 => n5975, ZN => n36304);
   U29892 : NAND2_X2 port map( A1 => n1222, A2 => n27197, ZN => n27354);
   U29894 : XOR2_X1 port map( A1 => n39487, A2 => n22581, Z => n1758);
   U29895 : XOR2_X1 port map( A1 => n4720, A2 => n22492, Z => n39487);
   U29897 : BUF_X2 port map( I => n2980, Z => n39488);
   U29903 : NOR3_X2 port map( A1 => n25499, A2 => n32365, A3 => n3735, ZN => 
                           n19240);
   U29912 : NAND2_X2 port map( A1 => n22327, A2 => n4108, ZN => n13163);
   U29916 : NAND2_X2 port map( A1 => n27144, A2 => n9593, ZN => n19455);
   U29927 : OAI21_X2 port map( A1 => n16708, A2 => n26684, B => n16707, ZN => 
                           n27144);
   U29942 : XOR2_X1 port map( A1 => n39631, A2 => n29092, Z => n39490);
   U29960 : NAND3_X2 port map( A1 => n13616, A2 => n13615, A3 => n22056, ZN => 
                           n22439);
   U29972 : XOR2_X1 port map( A1 => n39493, A2 => n36513, Z => Ciphertext(141))
                           ;
   U29975 : NOR2_X1 port map( A1 => n36848, A2 => n32531, ZN => n39493);
   U29978 : NOR2_X2 port map( A1 => n18304, A2 => n35253, ZN => n2057);
   U29985 : OAI21_X2 port map( A1 => n37192, A2 => n39494, B => n1223, ZN => 
                           n34890);
   U29989 : NOR2_X1 port map( A1 => n14327, A2 => n27389, ZN => n39494);
   U29995 : BUF_X2 port map( I => n18959, Z => n39495);
   U29996 : NAND2_X2 port map( A1 => n5093, A2 => n9141, ZN => n16107);
   U29997 : NAND2_X2 port map( A1 => n5498, A2 => n5496, ZN => n7432);
   U30005 : AND2_X1 port map( A1 => n28236, A2 => n39488, Z => n27990);
   U30006 : XOR2_X1 port map( A1 => n35208, A2 => n39497, Z => n32516);
   U30009 : INV_X2 port map( I => n29833, ZN => n39497);
   U30014 : OAI22_X2 port map( A1 => n28499, A2 => n27941, B1 => n4697, B2 => 
                           n28498, ZN => n29833);
   U30016 : AOI21_X1 port map( A1 => n11398, A2 => n11397, B => n1379, ZN => 
                           n30577);
   U30017 : NOR2_X1 port map( A1 => n20321, A2 => n37084, ZN => n34061);
   U30019 : AOI22_X2 port map( A1 => n15292, A2 => n18293, B1 => n11900, B2 => 
                           n8495, ZN => n4823);
   U30022 : NOR2_X2 port map( A1 => n14783, A2 => n21930, ZN => n15292);
   U30023 : XOR2_X1 port map( A1 => n11739, A2 => n24077, Z => n12798);
   U30030 : OAI21_X2 port map( A1 => n4960, A2 => n21014, B => n12746, ZN => 
                           n24077);
   U30034 : NAND3_X1 port map( A1 => n7852, A2 => n5896, A3 => n39098, ZN => 
                           n34881);
   U30035 : NAND2_X1 port map( A1 => n6539, A2 => n6540, ZN => n39498);
   U30039 : NAND2_X1 port map( A1 => n6353, A2 => n31875, ZN => n39499);
   U30041 : BUF_X2 port map( I => n14817, Z => n39500);
   U30044 : XOR2_X1 port map( A1 => n22444, A2 => n22500, Z => n22544);
   U30045 : NAND2_X2 port map( A1 => n22347, A2 => n22346, ZN => n22444);
   U30049 : XOR2_X1 port map( A1 => n22648, A2 => n22715, Z => n13961);
   U30054 : NAND2_X2 port map( A1 => n33155, A2 => n16712, ZN => n23794);
   U30056 : OAI21_X1 port map( A1 => n30145, A2 => n30134, B => n18424, ZN => 
                           n30135);
   U30058 : NAND2_X2 port map( A1 => n18588, A2 => n18241, ZN => n18424);
   U30059 : XOR2_X1 port map( A1 => n27647, A2 => n10301, Z => n27820);
   U30064 : NAND2_X2 port map( A1 => n34493, A2 => n16045, ZN => n27647);
   U30067 : NAND2_X2 port map( A1 => n30958, A2 => n12659, ZN => n35919);
   U30068 : XOR2_X1 port map( A1 => n25005, A2 => n16192, Z => n16191);
   U30071 : NAND3_X1 port map( A1 => n27334, A2 => n1218, A3 => n35115, ZN => 
                           n26846);
   U30072 : NAND2_X1 port map( A1 => n8650, A2 => n7607, ZN => n2130);
   U30078 : NAND2_X2 port map( A1 => n39509, A2 => n15834, ZN => n334);
   U30079 : INV_X2 port map( I => n39511, ZN => n4306);
   U30080 : XOR2_X1 port map( A1 => n291, A2 => n4204, Z => n39512);
   U30084 : NAND2_X1 port map( A1 => n29532, A2 => n29525, ZN => n29524);
   U30085 : NAND2_X2 port map( A1 => n36469, A2 => n10259, ZN => n29532);
   U30087 : NAND2_X2 port map( A1 => n34982, A2 => n9535, ZN => n34977);
   U30088 : NAND2_X2 port map( A1 => n3193, A2 => n18696, ZN => n28546);
   U30092 : OR3_X1 port map( A1 => n23610, A2 => n1627, A3 => n37088, Z => 
                           n35397);
   U30093 : XOR2_X1 port map( A1 => n39516, A2 => n2727, Z => n5514);
   U30095 : XOR2_X1 port map( A1 => n36915, A2 => n33007, Z => n26779);
   U30097 : XOR2_X1 port map( A1 => n20753, A2 => n22642, Z => n11377);
   U30100 : XOR2_X1 port map( A1 => n17189, A2 => n22552, Z => n22642);
   U30105 : OAI22_X2 port map( A1 => n26955, A2 => n8415, B1 => n31982, B2 => 
                           n8103, ZN => n39517);
   U30106 : NOR2_X2 port map( A1 => n20376, A2 => n19017, ZN => n20375);
   U30111 : NAND2_X2 port map( A1 => n39771, A2 => n37180, ZN => n19017);
   U30112 : INV_X2 port map( I => n39519, ZN => n36728);
   U30116 : XOR2_X1 port map( A1 => n34178, A2 => n38190, Z => n15304);
   U30122 : XOR2_X1 port map( A1 => n27645, A2 => n31233, Z => n34544);
   U30123 : XOR2_X1 port map( A1 => n19405, A2 => n12985, Z => n39520);
   U30126 : AOI21_X2 port map( A1 => n28543, A2 => n37956, B => n11474, ZN => 
                           n29067);
   U30127 : XOR2_X1 port map( A1 => n38584, A2 => n26556, Z => n26483);
   U30135 : NAND2_X2 port map( A1 => n33557, A2 => n30199, ZN => n30213);
   U30139 : XOR2_X1 port map( A1 => n39522, A2 => n19908, Z => Ciphertext(182))
                           ;
   U30143 : BUF_X2 port map( I => n16502, Z => n39523);
   U30146 : AOI22_X2 port map( A1 => n39524, A2 => n28450, B1 => n18972, B2 => 
                           n18971, ZN => n27957);
   U30147 : NOR2_X2 port map( A1 => n35830, A2 => n12543, ZN => n39524);
   U30148 : OAI21_X2 port map( A1 => n12276, A2 => n12275, B => n30048, ZN => 
                           n39525);
   U30152 : AOI22_X2 port map( A1 => n5678, A2 => n13705, B1 => n31512, B2 => 
                           n29979, ZN => n29982);
   U30154 : XOR2_X1 port map( A1 => n6325, A2 => n37194, Z => n7201);
   U30165 : XNOR2_X1 port map( A1 => n12267, A2 => n22790, ZN => n6325);
   U30169 : INV_X2 port map( I => n32981, ZN => n4573);
   U30172 : NAND2_X1 port map( A1 => n19097, A2 => n18081, ZN => n29911);
   U30175 : XOR2_X1 port map( A1 => n28999, A2 => n15565, Z => n39529);
   U30176 : OAI21_X2 port map( A1 => n39530, A2 => n32719, B => n20764, ZN => 
                           n13278);
   U30178 : XOR2_X1 port map( A1 => n26572, A2 => n26229, Z => n26577);
   U30182 : BUF_X2 port map( I => n20158, Z => n39537);
   U30183 : INV_X2 port map( I => n33323, ZN => n36867);
   U30185 : NAND3_X2 port map( A1 => n14498, A2 => n19080, A3 => n18872, ZN => 
                           n33323);
   U30186 : NAND2_X2 port map( A1 => n39539, A2 => n33392, ZN => n36301);
   U30188 : NAND2_X2 port map( A1 => n24778, A2 => n39540, ZN => n39539);
   U30189 : NAND2_X2 port map( A1 => n19593, A2 => n13300, ZN => n24778);
   U30190 : NOR2_X1 port map( A1 => n23128, A2 => n13688, ZN => n7504);
   U30201 : NAND2_X1 port map( A1 => n3725, A2 => n2944, ZN => n5107);
   U30202 : BUF_X2 port map( I => n19849, Z => n39541);
   U30204 : NOR2_X2 port map( A1 => n12509, A2 => n11240, ZN => n11434);
   U30205 : XOR2_X1 port map( A1 => n39543, A2 => n29854, Z => Ciphertext(116))
                           ;
   U30207 : NAND2_X1 port map( A1 => n19872, A2 => n30616, ZN => n39543);
   U30212 : NOR2_X1 port map( A1 => n6191, A2 => n4272, ZN => n27017);
   U30213 : XOR2_X1 port map( A1 => n5308, A2 => n25242, Z => n39544);
   U30214 : XOR2_X1 port map( A1 => n23931, A2 => n23841, Z => n23985);
   U30218 : NAND2_X2 port map( A1 => n23369, A2 => n23368, ZN => n23841);
   U30219 : XOR2_X1 port map( A1 => n233, A2 => n10309, Z => n25380);
   U30224 : INV_X1 port map( I => n31488, ZN => n39660);
   U30227 : NAND2_X2 port map( A1 => n20108, A2 => n15884, ZN => n32377);
   U30228 : INV_X2 port map( I => n4381, ZN => n25975);
   U30231 : NAND2_X2 port map( A1 => n2626, A2 => n18787, ZN => n4381);
   U30238 : XOR2_X1 port map( A1 => n14231, A2 => n19849, Z => n11899);
   U30240 : NAND3_X2 port map( A1 => n6409, A2 => n6408, A3 => n9500, ZN => 
                           n19849);
   U30242 : AOI21_X2 port map( A1 => n39545, A2 => n32977, B => n10228, ZN => 
                           n18571);
   U30243 : NAND2_X2 port map( A1 => n345, A2 => n11526, ZN => n39545);
   U30245 : AND2_X1 port map( A1 => n4272, A2 => n39546, Z => n20709);
   U30249 : XOR2_X1 port map( A1 => n39547, A2 => n27726, Z => n31442);
   U30251 : XOR2_X1 port map( A1 => n32015, A2 => n27823, Z => n39547);
   U30252 : OAI21_X2 port map( A1 => n26236, A2 => n30883, B => n14157, ZN => 
                           n26035);
   U30253 : NAND2_X2 port map( A1 => n31994, A2 => n39375, ZN => n14157);
   U30254 : NAND2_X2 port map( A1 => n7695, A2 => n8770, ZN => n5126);
   U30256 : XOR2_X1 port map( A1 => n39549, A2 => n8856, Z => n32893);
   U30263 : XOR2_X1 port map( A1 => n7358, A2 => n31541, Z => n39549);
   U30267 : XOR2_X1 port map( A1 => n25268, A2 => n25188, Z => n39550);
   U30268 : XOR2_X1 port map( A1 => Plaintext(120), A2 => Key(120), Z => n33999
                           );
   U30271 : OR2_X1 port map( A1 => n26833, A2 => n30853, Z => n32941);
   U30274 : XNOR2_X1 port map( A1 => n22736, A2 => n22714, ZN => n36195);
   U30275 : NAND2_X2 port map( A1 => n39551, A2 => n39586, ZN => n6002);
   U30277 : NAND2_X2 port map( A1 => n22101, A2 => n38830, ZN => n22098);
   U30279 : NAND2_X2 port map( A1 => n27235, A2 => n27436, ZN => n27150);
   U30281 : NOR2_X2 port map( A1 => n20492, A2 => n20493, ZN => n6435);
   U30282 : NOR2_X2 port map( A1 => n13501, A2 => n33433, ZN => n6844);
   U30289 : XOR2_X1 port map( A1 => n39552, A2 => n7664, Z => n10006);
   U30291 : XOR2_X1 port map( A1 => n27683, A2 => n27632, Z => n27782);
   U30295 : XOR2_X1 port map( A1 => n27504, A2 => n19758, Z => n27505);
   U30296 : NAND2_X2 port map( A1 => n15058, A2 => n14084, ZN => n27504);
   U30299 : XOR2_X1 port map( A1 => n39553, A2 => n16532, Z => n5603);
   U30301 : XOR2_X1 port map( A1 => n16531, A2 => n17117, Z => n39553);
   U30304 : NOR2_X1 port map( A1 => n16946, A2 => n27320, ZN => n39554);
   U30307 : XOR2_X1 port map( A1 => n39556, A2 => n30179, Z => Ciphertext(178))
                           ;
   U30311 : NAND3_X2 port map( A1 => n34903, A2 => n5422, A3 => n17168, ZN => 
                           n39556);
   U30312 : NOR2_X2 port map( A1 => n24350, A2 => n24349, ZN => n5957);
   U30313 : OAI21_X2 port map( A1 => n20022, A2 => n20021, B => n39557, ZN => 
                           n27446);
   U30318 : XOR2_X1 port map( A1 => n6196, A2 => n6930, Z => n28985);
   U30325 : NAND2_X2 port map( A1 => n11911, A2 => n9625, ZN => n6930);
   U30335 : XOR2_X1 port map( A1 => n14231, A2 => n30179, Z => n25221);
   U30339 : AOI22_X2 port map( A1 => n8296, A2 => n1122, B1 => n14266, B2 => 
                           n36228, ZN => n14231);
   U30342 : XOR2_X1 port map( A1 => n39558, A2 => n22590, Z => n36038);
   U30344 : XOR2_X1 port map( A1 => n7560, A2 => n39559, Z => n39558);
   U30345 : XOR2_X1 port map( A1 => n39560, A2 => n10365, Z => n20087);
   U30351 : XOR2_X1 port map( A1 => n28332, A2 => n28333, Z => n39560);
   U30353 : NAND2_X2 port map( A1 => n3535, A2 => n31319, ZN => n35664);
   U30355 : XOR2_X1 port map( A1 => n20213, A2 => n39561, Z => n35711);
   U30358 : NAND2_X2 port map( A1 => n15377, A2 => n15378, ZN => n20213);
   U30361 : NAND2_X2 port map( A1 => n39562, A2 => n11258, ZN => n15030);
   U30363 : XOR2_X1 port map( A1 => n39563, A2 => n518, Z => n12293);
   U30365 : XOR2_X1 port map( A1 => n26591, A2 => n26305, Z => n26210);
   U30368 : NOR2_X2 port map( A1 => n5881, A2 => n5884, ZN => n26305);
   U30369 : XOR2_X1 port map( A1 => n11350, A2 => n11349, Z => n11348);
   U30370 : INV_X4 port map( I => n19279, ZN => n32802);
   U30371 : NAND2_X2 port map( A1 => n4538, A2 => n31376, ZN => n6560);
   U30375 : AND2_X1 port map( A1 => n4386, A2 => n11415, Z => n3820);
   U30381 : NAND2_X2 port map( A1 => n9746, A2 => n36700, ZN => n14833);
   U30385 : NAND2_X1 port map( A1 => n27185, A2 => n4964, ZN => n39566);
   U30387 : XOR2_X1 port map( A1 => n27845, A2 => n16613, Z => n27763);
   U30388 : NAND2_X2 port map( A1 => n39567, A2 => n3819, ZN => n4378);
   U30389 : NOR2_X1 port map( A1 => n25813, A2 => n25936, ZN => n25937);
   U30390 : XOR2_X1 port map( A1 => n27853, A2 => n35610, Z => n27856);
   U30393 : NAND2_X2 port map( A1 => n39568, A2 => n35492, ZN => n25887);
   U30394 : NAND2_X2 port map( A1 => n19759, A2 => n8131, ZN => n5465);
   U30397 : NOR2_X2 port map( A1 => n30342, A2 => n9889, ZN => n17925);
   U30401 : INV_X2 port map( I => n39570, ZN => n9893);
   U30402 : NOR2_X1 port map( A1 => n980, A2 => n37804, ZN => n18018);
   U30404 : BUF_X2 port map( I => n23969, Z => n39575);
   U30405 : AOI22_X2 port map( A1 => n26694, A2 => n19455, B1 => n3783, B2 => 
                           n21144, ZN => n10998);
   U30406 : INV_X2 port map( I => n39577, ZN => n17314);
   U30408 : XOR2_X1 port map( A1 => n27857, A2 => n20032, Z => n39577);
   U30409 : AOI21_X1 port map( A1 => n30113, A2 => n30119, B => n39578, ZN => 
                           n30116);
   U30413 : XOR2_X1 port map( A1 => n27757, A2 => n10707, Z => n5484);
   U30415 : BUF_X2 port map( I => n12649, Z => n39579);
   U30417 : XOR2_X1 port map( A1 => n9119, A2 => n7623, Z => n9118);
   U30418 : OAI22_X1 port map( A1 => n28364, A2 => n1193, B1 => n28365, B2 => 
                           n33460, ZN => n5150);
   U30419 : XOR2_X1 port map( A1 => n39580, A2 => n36087, Z => n15903);
   U30420 : XOR2_X1 port map( A1 => n6291, A2 => n32090, Z => n39580);
   U30423 : XOR2_X1 port map( A1 => n20987, A2 => n35317, Z => n39600);
   U30424 : NAND2_X2 port map( A1 => n17093, A2 => n16842, ZN => n39581);
   U30426 : NOR2_X1 port map( A1 => n7099, A2 => n36435, ZN => n4459);
   U30431 : AND2_X1 port map( A1 => n13686, A2 => n36355, Z => n10564);
   U30432 : BUF_X2 port map( I => n840, Z => n39584);
   U30433 : NAND2_X2 port map( A1 => n39587, A2 => n13264, ZN => n24732);
   U30435 : NAND2_X2 port map( A1 => n39589, A2 => n32408, ZN => n3967);
   U30436 : OAI22_X2 port map( A1 => n22220, A2 => n22223, B1 => n8792, B2 => 
                           n22222, ZN => n39589);
   U30437 : OAI21_X2 port map( A1 => n14082, A2 => n6592, B => n19589, ZN => 
                           n14273);
   U30440 : XOR2_X1 port map( A1 => n39590, A2 => n13654, Z => n205);
   U30441 : XOR2_X1 port map( A1 => n39591, A2 => n17000, Z => n19473);
   U30443 : XOR2_X1 port map( A1 => n14191, A2 => n15978, Z => n34611);
   U30444 : OR2_X1 port map( A1 => n22084, A2 => n2257, Z => n39592);
   U30445 : XOR2_X1 port map( A1 => n26181, A2 => n26399, Z => n6134);
   U30448 : XOR2_X1 port map( A1 => n26585, A2 => n19847, Z => n26181);
   U30451 : AOI22_X2 port map( A1 => n39593, A2 => n28641, B1 => n28640, B2 => 
                           n15447, ZN => n20452);
   U30452 : OAI22_X2 port map( A1 => n15447, A2 => n28639, B1 => n4369, B2 => 
                           n28637, ZN => n39593);
   U30461 : NOR3_X2 port map( A1 => n7086, A2 => n13444, A3 => n20041, ZN => 
                           n6914);
   U30469 : NAND2_X2 port map( A1 => n32741, A2 => n16406, ZN => n39681);
   U30471 : NAND2_X1 port map( A1 => n336, A2 => n27422, ZN => n33799);
   U30473 : NAND2_X1 port map( A1 => n23518, A2 => n23517, ZN => n19283);
   U30476 : NOR2_X2 port map( A1 => n22842, A2 => n22841, ZN => n23517);
   U30477 : NAND2_X1 port map( A1 => n18850, A2 => n8660, ZN => n23312);
   U30478 : NOR2_X2 port map( A1 => n34001, A2 => n27363, ZN => n16482);
   U30480 : NAND2_X2 port map( A1 => n18023, A2 => n18024, ZN => n27363);
   U30481 : BUF_X2 port map( I => n26729, Z => n39595);
   U30482 : NAND2_X2 port map( A1 => n6282, A2 => n2349, ZN => n33539);
   U30483 : INV_X1 port map( I => n22552, ZN => n39630);
   U30484 : XOR2_X1 port map( A1 => n26509, A2 => n26587, Z => n39596);
   U30486 : OAI21_X1 port map( A1 => n26864, A2 => n26952, B => n39737, ZN => 
                           n32176);
   U30493 : INV_X2 port map( I => n39597, ZN => n27200);
   U30494 : NOR2_X2 port map( A1 => n17072, A2 => n7424, ZN => n39597);
   U30496 : BUF_X2 port map( I => n1230, Z => n39598);
   U30501 : NOR2_X1 port map( A1 => n11415, A2 => n4356, ZN => n33276);
   U30503 : NAND2_X1 port map( A1 => n22939, A2 => n10247, ZN => n39601);
   U30504 : NAND2_X1 port map( A1 => n29946, A2 => n11861, ZN => n29841);
   U30507 : XOR2_X1 port map( A1 => n25183, A2 => n39604, Z => n34911);
   U30508 : XOR2_X1 port map( A1 => n39320, A2 => n37109, Z => n39604);
   U30509 : XOR2_X1 port map( A1 => n27805, A2 => n13568, Z => n13608);
   U30516 : NAND2_X2 port map( A1 => n17893, A2 => n17891, ZN => n12846);
   U30517 : AOI21_X2 port map( A1 => n34143, A2 => n24605, B => n33392, ZN => 
                           n24607);
   U30518 : NOR2_X2 port map( A1 => n39606, A2 => n21852, ZN => n21856);
   U30519 : OAI21_X2 port map( A1 => n1355, A2 => n693, B => n6234, ZN => 
                           n39606);
   U30521 : BUF_X2 port map( I => n17861, Z => n39607);
   U30524 : INV_X2 port map( I => n39608, ZN => n34160);
   U30525 : XOR2_X1 port map( A1 => n1556, A2 => n17445, Z => n39609);
   U30528 : NOR2_X2 port map( A1 => n11469, A2 => n39610, ZN => n35793);
   U30532 : INV_X2 port map( I => n28491, ZN => n39610);
   U30533 : NAND2_X2 port map( A1 => n18910, A2 => n16619, ZN => n28491);
   U30538 : XOR2_X1 port map( A1 => n36961, A2 => n26474, Z => n39612);
   U30541 : XOR2_X1 port map( A1 => n39613, A2 => n12556, Z => n4752);
   U30543 : XOR2_X1 port map( A1 => n8952, A2 => n18577, Z => n39614);
   U30545 : XOR2_X1 port map( A1 => n26503, A2 => n39615, Z => n412);
   U30546 : XOR2_X1 port map( A1 => n26504, A2 => n36333, Z => n39615);
   U30551 : AOI22_X2 port map( A1 => n39617, A2 => n9543, B1 => n23042, B2 => 
                           n22833, ZN => n7024);
   U30554 : INV_X2 port map( I => n13485, ZN => n39617);
   U30555 : NAND2_X2 port map( A1 => n38329, A2 => n33431, ZN => n13485);
   U30556 : NAND2_X2 port map( A1 => n32, A2 => n3913, ZN => n3907);
   U30557 : NAND2_X2 port map( A1 => n8699, A2 => n8294, ZN => n10221);
   U30564 : NOR2_X2 port map( A1 => n4173, A2 => n4172, ZN => n39624);
   U30567 : OAI21_X2 port map( A1 => n21713, A2 => n19542, B => n21652, ZN => 
                           n39619);
   U30568 : XOR2_X1 port map( A1 => n24560, A2 => n24563, Z => n39621);
   U30571 : OAI22_X2 port map( A1 => n39546, A2 => n27221, B1 => n38488, B2 => 
                           n39424, ZN => n27297);
   U30575 : XOR2_X1 port map( A1 => n382, A2 => n25215, Z => n8920);
   U30578 : NAND2_X2 port map( A1 => n13386, A2 => n19682, ZN => n24342);
   U30584 : XOR2_X1 port map( A1 => n11451, A2 => n33809, Z => n11449);
   U30589 : NAND2_X2 port map( A1 => n39623, A2 => n7565, ZN => n6944);
   U30593 : NAND3_X1 port map( A1 => n24205, A2 => n37264, A3 => n24206, ZN => 
                           n39623);
   U30594 : NAND2_X2 port map( A1 => n39624, A2 => n34461, ZN => n35500);
   U30596 : NOR2_X2 port map( A1 => n30825, A2 => n37139, ZN => n3993);
   U30606 : OAI21_X2 port map( A1 => n2058, A2 => n7036, B => n35647, ZN => 
                           n5634);
   U30607 : NAND2_X2 port map( A1 => n6786, A2 => n6790, ZN => n28758);
   U30608 : AOI22_X2 port map( A1 => n23011, A2 => n5702, B1 => n4931, B2 => 
                           n1318, ZN => n16416);
   U30611 : XOR2_X1 port map( A1 => n9923, A2 => n17494, Z => n17698);
   U30613 : NAND2_X1 port map( A1 => n8027, A2 => n39629, ZN => n33667);
   U30614 : NAND2_X1 port map( A1 => n33786, A2 => n32366, ZN => n39629);
   U30616 : INV_X2 port map( I => n23970, ZN => n15336);
   U30617 : AND2_X1 port map( A1 => n33738, A2 => n2153, Z => n21991);
   U30618 : XOR2_X1 port map( A1 => n22464, A2 => n11974, Z => n15671);
   U30621 : NAND2_X2 port map( A1 => n38282, A2 => n12029, ZN => n31049);
   U30622 : OR2_X1 port map( A1 => n11764, A2 => n11763, Z => n39633);
   U30625 : XOR2_X1 port map( A1 => n10767, A2 => n39634, Z => n34223);
   U30626 : OAI21_X2 port map( A1 => n35819, A2 => n35820, B => n39635, ZN => 
                           n27914);
   U30630 : NAND2_X2 port map( A1 => n28133, A2 => n28229, ZN => n39635);
   U30632 : XOR2_X1 port map( A1 => n12183, A2 => n36952, Z => n7273);
   U30633 : XOR2_X1 port map( A1 => n9943, A2 => n14062, Z => n5891);
   U30634 : INV_X2 port map( I => n39638, ZN => n11636);
   U30637 : INV_X2 port map( I => n39639, ZN => n693);
   U30638 : XNOR2_X1 port map( A1 => Plaintext(36), A2 => Key(36), ZN => n39639
                           );
   U30639 : NAND2_X1 port map( A1 => n39642, A2 => n39640, ZN => n26640);
   U30644 : NAND2_X1 port map( A1 => n39641, A2 => n26764, ZN => n39640);
   U30653 : INV_X1 port map( I => n26763, ZN => n39641);
   U30658 : NAND2_X1 port map( A1 => n13393, A2 => n26763, ZN => n39642);
   U30659 : OAI22_X2 port map( A1 => n19893, A2 => n8082, B1 => n16067, B2 => 
                           n28390, ZN => n39643);
   U30660 : XOR2_X1 port map( A1 => n39644, A2 => n16091, Z => n287);
   U30663 : XOR2_X1 port map( A1 => n37256, A2 => n35249, Z => n39644);
   U30665 : AOI22_X2 port map( A1 => n2434, A2 => n12080, B1 => n2435, B2 => 
                           n8749, ZN => n31476);
   U30667 : XOR2_X1 port map( A1 => Key(37), A2 => Plaintext(37), Z => n35161);
   U30668 : OAI21_X2 port map( A1 => n39645, A2 => n15739, B => n33045, ZN => 
                           n6089);
   U30670 : NOR2_X2 port map( A1 => n31283, A2 => n921, ZN => n3699);
   U30673 : NAND2_X2 port map( A1 => n31205, A2 => n26023, ZN => n25771);
   U30677 : NAND3_X1 port map( A1 => n9553, A2 => n3511, A3 => n17197, ZN => 
                           n33805);
   U30679 : INV_X2 port map( I => n32153, ZN => n33599);
   U30680 : XOR2_X1 port map( A1 => n30458, A2 => n30963, Z => n32153);
   U30681 : OAI21_X2 port map( A1 => n451, A2 => n450, B => n38172, ZN => n5344
                           );
   U30683 : NAND2_X2 port map( A1 => n20959, A2 => n39649, ZN => n13917);
   U30684 : AOI22_X2 port map( A1 => n15193, A2 => n20155, B1 => n16871, B2 => 
                           n39258, ZN => n39649);
   U30686 : NAND2_X1 port map( A1 => n30844, A2 => n38197, ZN => n39821);
   U30687 : NAND2_X2 port map( A1 => n38206, A2 => n18042, ZN => n18908);
   U30688 : XOR2_X1 port map( A1 => n34894, A2 => n4305, Z => n31370);
   U30691 : AOI22_X1 port map( A1 => n29577, A2 => n20437, B1 => n31899, B2 => 
                           n29575, ZN => n17113);
   U30692 : NOR2_X2 port map( A1 => n1222, A2 => n27197, ZN => n3783);
   U30694 : XOR2_X1 port map( A1 => n19024, A2 => n39652, Z => n39651);
   U30700 : INV_X2 port map( I => n26498, ZN => n39652);
   U30701 : AOI22_X2 port map( A1 => n35274, A2 => n20357, B1 => n3833, B2 => 
                           n19778, ZN => n36886);
   U30702 : NAND2_X2 port map( A1 => n22304, A2 => n3835, ZN => n35274);
   U30705 : NAND2_X2 port map( A1 => n6228, A2 => n37215, ZN => n6727);
   U30706 : INV_X2 port map( I => n39653, ZN => n39814);
   U30707 : XOR2_X1 port map( A1 => n10275, A2 => n10278, Z => n39653);
   U30708 : INV_X1 port map( I => n27581, ZN => n19396);
   U30711 : XOR2_X1 port map( A1 => n27581, A2 => n27669, Z => n27552);
   U30712 : XOR2_X1 port map( A1 => n6757, A2 => n17455, Z => n21098);
   U30714 : NAND2_X2 port map( A1 => n25596, A2 => n35821, ZN => n6757);
   U30716 : XOR2_X1 port map( A1 => n27661, A2 => n27662, Z => n27840);
   U30717 : NOR2_X1 port map( A1 => n17121, A2 => n30194, ZN => n17120);
   U30721 : XOR2_X1 port map( A1 => n15592, A2 => n39655, Z => n30966);
   U30722 : XOR2_X1 port map( A1 => n5407, A2 => n25219, Z => n39657);
   U30725 : NOR2_X2 port map( A1 => n21738, A2 => n19335, ZN => n22295);
   U30726 : OAI21_X2 port map( A1 => n2057, A2 => n20989, B => n24382, ZN => 
                           n16184);
   U30728 : NOR2_X2 port map( A1 => n33834, A2 => n18407, ZN => n9412);
   U30729 : OR2_X2 port map( A1 => n8653, A2 => n8517, Z => n21899);
   U30731 : AOI21_X2 port map( A1 => n22288, A2 => n1687, B => n1328, ZN => 
                           n5556);
   U30732 : XNOR2_X1 port map( A1 => n31151, A2 => n33166, ZN => n39663);
   U30733 : OR2_X1 port map( A1 => n33347, A2 => n19410, Z => n27934);
   U30737 : AND2_X2 port map( A1 => n17424, A2 => n17425, Z => n29461);
   U30739 : OR2_X1 port map( A1 => n32899, A2 => n4880, Z => n31786);
   U30741 : BUF_X2 port map( I => n13285, Z => n39666);
   U30743 : XOR2_X1 port map( A1 => n26318, A2 => n26317, Z => n39667);
   U30746 : XOR2_X1 port map( A1 => n26491, A2 => n2545, Z => n32954);
   U30747 : OR2_X1 port map( A1 => n35431, A2 => n21802, Z => n39668);
   U30752 : OR2_X1 port map( A1 => n1230, A2 => n14962, Z => n26865);
   U30753 : NOR2_X2 port map( A1 => n3562, A2 => n21869, ZN => n21867);
   U30754 : NAND2_X2 port map( A1 => n12529, A2 => n34340, ZN => n5383);
   U30756 : INV_X2 port map( I => n39669, ZN => n34116);
   U30759 : NOR2_X2 port map( A1 => n14037, A2 => n18303, ZN => n39669);
   U30761 : NAND2_X2 port map( A1 => n12252, A2 => n155, ZN => n26359);
   U30765 : INV_X2 port map( I => n27233, ZN => n39671);
   U30770 : BUF_X2 port map( I => n21683, Z => n39672);
   U30771 : XOR2_X1 port map( A1 => n2512, A2 => n23841, Z => n23866);
   U30776 : NOR2_X2 port map( A1 => n13537, A2 => n39673, ZN => n13536);
   U30781 : INV_X1 port map( I => n39674, ZN => n39673);
   U30785 : NAND2_X1 port map( A1 => n10414, A2 => n37051, ZN => n39674);
   U30786 : XOR2_X1 port map( A1 => n26435, A2 => n39675, Z => n26201);
   U30790 : XOR2_X1 port map( A1 => n34469, A2 => n20600, Z => n39675);
   U30797 : AOI21_X2 port map( A1 => n33753, A2 => n39248, B => n39676, ZN => 
                           n14504);
   U30799 : INV_X2 port map( I => n18661, ZN => n39676);
   U30800 : BUF_X2 port map( I => n8219, Z => n39678);
   U30802 : XOR2_X1 port map( A1 => n39679, A2 => n26385, Z => n18390);
   U30803 : XOR2_X1 port map( A1 => n9984, A2 => n26176, Z => n39679);
   U30806 : INV_X1 port map( I => n39488, ZN => n2302);
   U30807 : XOR2_X1 port map( A1 => n2134, A2 => n31794, Z => n2980);
   U30811 : XOR2_X1 port map( A1 => n31162, A2 => n13934, Z => n29347);
   U30813 : XOR2_X1 port map( A1 => n29142, A2 => n19866, Z => n16091);
   U30814 : OAI21_X2 port map( A1 => n36517, A2 => n17447, B => n8788, ZN => 
                           n12885);
   U30817 : XOR2_X1 port map( A1 => n5316, A2 => n5315, Z => n6145);
   U30819 : XOR2_X1 port map( A1 => n27805, A2 => n12507, Z => n19989);
   U30820 : NOR2_X1 port map( A1 => n32204, A2 => n19163, ZN => n34287);
   U30821 : XOR2_X1 port map( A1 => n11290, A2 => n11288, Z => n11481);
   U30822 : NOR3_X2 port map( A1 => n19549, A2 => n39656, A3 => n16305, ZN => 
                           n7315);
   U30823 : AND2_X2 port map( A1 => n29968, A2 => n18896, Z => n29973);
   U30827 : XOR2_X1 port map( A1 => n12884, A2 => n39683, Z => n3770);
   U30828 : XOR2_X1 port map( A1 => n27753, A2 => n37195, Z => n39683);
   U30831 : XOR2_X1 port map( A1 => n3081, A2 => n3632, Z => n18806);
   U30832 : XOR2_X1 port map( A1 => n22639, A2 => n22640, Z => n34289);
   U30836 : NOR2_X2 port map( A1 => n6348, A2 => n39684, ZN => n6347);
   U30837 : OAI22_X2 port map( A1 => n21560, A2 => n19397, B1 => n21477, B2 => 
                           n8597, ZN => n39684);
   U30839 : NOR2_X2 port map( A1 => n11759, A2 => n36800, ZN => n24673);
   U30841 : NAND2_X2 port map( A1 => n21796, A2 => n7047, ZN => n31202);
   U30844 : NOR2_X1 port map( A1 => n24156, A2 => n37267, ZN => n24303);
   U30852 : NAND3_X2 port map( A1 => n28452, A2 => n35793, A3 => n4523, ZN => 
                           n29121);
   U30860 : XOR2_X1 port map( A1 => n15336, A2 => n31775, Z => n13736);
   U30861 : NAND2_X1 port map( A1 => n31812, A2 => n3978, ZN => n39721);
   U30864 : OAI21_X2 port map( A1 => n37981, A2 => n28639, B => n39355, ZN => 
                           n30757);
   U30869 : AOI21_X1 port map( A1 => n6323, A2 => n29479, B => n29478, ZN => 
                           n6322);
   U30870 : XOR2_X1 port map( A1 => n36544, A2 => n9989, Z => n26183);
   U30871 : OAI22_X2 port map( A1 => n20296, A2 => n1253, B1 => n20295, B2 => 
                           n25448, ZN => n39687);
   U30872 : NAND2_X2 port map( A1 => n20979, A2 => n10896, ZN => n29644);
   U30873 : XOR2_X1 port map( A1 => n5026, A2 => n39688, Z => n6596);
   U30874 : XOR2_X1 port map( A1 => n6598, A2 => n518, Z => n39688);
   U30875 : AND2_X1 port map( A1 => n19605, A2 => n28132, Z => n28223);
   U30876 : BUF_X2 port map( I => n29659, Z => n39689);
   U30877 : NAND2_X1 port map( A1 => n35686, A2 => n24874, ZN => n9211);
   U30878 : XOR2_X1 port map( A1 => n38154, A2 => n20454, Z => n10117);
   U30879 : NAND2_X1 port map( A1 => n6946, A2 => n21995, ZN => n6949);
   U30880 : AOI22_X2 port map( A1 => n20121, A2 => n25688, B1 => n25393, B2 => 
                           n25689, ZN => n39690);
   U30881 : XOR2_X1 port map( A1 => n34469, A2 => n20213, Z => n26569);
   U30882 : INV_X2 port map( I => n19443, ZN => n39691);
   U30883 : NAND2_X1 port map( A1 => n28017, A2 => n39692, ZN => n31799);
   U30884 : XNOR2_X1 port map( A1 => n23955, A2 => n37842, ZN => n39728);
   U30885 : OR2_X1 port map( A1 => n17692, A2 => n34013, Z => n23023);
   U30886 : NAND3_X1 port map( A1 => n22917, A2 => n23163, A3 => n36095, ZN => 
                           n11877);
   U30887 : NAND2_X1 port map( A1 => n9165, A2 => n22250, ZN => n9711);
   U30888 : NAND2_X2 port map( A1 => n7759, A2 => n9495, ZN => n9165);
   U30889 : XOR2_X1 port map( A1 => n39693, A2 => n22648, Z => n487);
   U30890 : XOR2_X1 port map( A1 => n291, A2 => n32309, Z => n39694);
   U30891 : XOR2_X1 port map( A1 => n39695, A2 => n30063, Z => Ciphertext(144))
                           ;
   U30892 : NAND2_X2 port map( A1 => n39697, A2 => n11507, ZN => n11541);
   U30893 : BUF_X2 port map( I => n6196, Z => n39698);
   U30894 : XOR2_X1 port map( A1 => n28969, A2 => n17250, Z => n10136);
   U30895 : XOR2_X1 port map( A1 => n38147, A2 => n29104, Z => n28969);
   U30896 : INV_X2 port map( I => n36380, ZN => n39699);
   U30897 : AOI21_X1 port map( A1 => n21873, A2 => n21874, B => n21872, ZN => 
                           n21879);
   U30898 : AOI21_X2 port map( A1 => n39700, A2 => n37183, B => n1546, ZN => 
                           n7097);
   U30899 : OAI22_X2 port map( A1 => n27085, A2 => n14261, B1 => n33979, B2 => 
                           n38211, ZN => n11590);
   U30900 : NAND2_X2 port map( A1 => n39701, A2 => n29948, ZN => n29979);
   U30901 : NAND2_X1 port map( A1 => n13085, A2 => n1904, ZN => n39701);
   U30902 : AOI22_X2 port map( A1 => n21020, A2 => n156, B1 => n39702, B2 => 
                           n9514, ZN => n3904);
   U30903 : OR2_X1 port map( A1 => n22796, A2 => n35213, Z => n23030);
   U30904 : XOR2_X1 port map( A1 => n130, A2 => n12205, Z => n22796);
   U30905 : NOR2_X2 port map( A1 => n23389, A2 => n4525, ZN => n9639);
   U30906 : BUF_X2 port map( I => n24300, Z => n39703);
   U30907 : BUF_X2 port map( I => n8430, Z => n39704);
   U30908 : XOR2_X1 port map( A1 => n26457, A2 => n4918, Z => n35923);
   U30909 : AOI22_X2 port map( A1 => n21766, A2 => n16945, B1 => n9759, B2 => 
                           n21499, ZN => n39705);
   U30910 : XNOR2_X1 port map( A1 => n22620, A2 => n22731, ZN => n22429);
   U30911 : OAI21_X2 port map( A1 => n5085, A2 => n37001, B => n39707, ZN => 
                           n11443);
   U30912 : XOR2_X1 port map( A1 => n39708, A2 => n7553, Z => n10737);
   U30913 : XOR2_X1 port map( A1 => n291, A2 => n12838, Z => n39708);
   U30914 : BUF_X2 port map( I => n18081, Z => n39709);
   U30915 : XOR2_X1 port map( A1 => n39710, A2 => n10920, Z => n36373);
   U30916 : BUF_X2 port map( I => n34644, Z => n39711);
   U30917 : XOR2_X1 port map( A1 => n33601, A2 => n29033, Z => n18288);
   U30918 : NAND2_X2 port map( A1 => n31486, A2 => n39768, ZN => n29747);
   U30919 : NAND2_X2 port map( A1 => n39715, A2 => n31904, ZN => n8375);
   U30920 : NAND2_X1 port map( A1 => n25305, A2 => n1535, ZN => n39715);
   U30921 : XOR2_X1 port map( A1 => n10380, A2 => n33789, Z => n10379);
   U30922 : XOR2_X1 port map( A1 => n16607, A2 => n16605, Z => n17313);
   U30923 : XOR2_X1 port map( A1 => n8755, A2 => n29293, Z => n29307);
   U30924 : NAND2_X1 port map( A1 => n4880, A2 => n10559, ZN => n34374);
   U30925 : XOR2_X1 port map( A1 => n27598, A2 => n39717, Z => n27603);
   U30926 : XOR2_X1 port map( A1 => n27597, A2 => n27596, Z => n39717);
   U30927 : XOR2_X1 port map( A1 => n22541, A2 => n39718, Z => n36812);
   U30928 : XOR2_X1 port map( A1 => n31504, A2 => n39630, Z => n39718);
   U30929 : XOR2_X1 port map( A1 => n33452, A2 => n23988, Z => n24043);
   U30930 : NOR2_X2 port map( A1 => n23016, A2 => n23015, ZN => n23988);
   U30931 : XOR2_X1 port map( A1 => n25145, A2 => n39720, Z => n39719);
   U30932 : OAI21_X1 port map( A1 => n15028, A2 => n14529, B => n31534, ZN => 
                           n15027);
   U30933 : NOR2_X2 port map( A1 => n32061, A2 => n23458, ZN => n23297);
   U30934 : NAND2_X2 port map( A1 => n39721, A2 => n4741, ZN => n9757);
   U30935 : NAND2_X2 port map( A1 => n39722, A2 => n15710, ZN => n8728);
   U30936 : BUF_X2 port map( I => n33509, Z => n39723);
   U30937 : XOR2_X1 port map( A1 => n4302, A2 => n25085, Z => n4305);
   U30938 : XOR2_X1 port map( A1 => n39726, A2 => n29091, Z => n29199);
   U30939 : XOR2_X1 port map( A1 => n7936, A2 => n6675, Z => n39726);
   U30940 : OAI21_X2 port map( A1 => n34682, A2 => n13270, B => n35258, ZN => 
                           n33255);
   U30941 : XOR2_X1 port map( A1 => n36000, A2 => n39727, Z => n8760);
   U30942 : XOR2_X1 port map( A1 => n23836, A2 => n39728, Z => n39727);
   U30943 : NAND2_X2 port map( A1 => n35926, A2 => n20825, ZN => n12793);
   U30944 : NAND3_X2 port map( A1 => n32159, A2 => n9330, A3 => n8013, ZN => 
                           n8660);
   U30945 : AOI21_X2 port map( A1 => n37106, A2 => n13495, B => n24630, ZN => 
                           n11082);
   U30946 : XOR2_X1 port map( A1 => n23947, A2 => n24006, Z => n15904);
   U30947 : XOR2_X1 port map( A1 => n27818, A2 => n31996, Z => n27884);
   U30948 : XOR2_X1 port map( A1 => n8920, A2 => n21252, Z => n8922);
   U30949 : NAND3_X2 port map( A1 => n4938, A2 => n24389, A3 => n24388, ZN => 
                           n19359);
   U30950 : AOI21_X1 port map( A1 => n32196, A2 => n31340, B => n26215, ZN => 
                           n16814);
   U30951 : NAND2_X2 port map( A1 => n12365, A2 => n14349, ZN => n17976);
   U30952 : NAND2_X1 port map( A1 => n39732, A2 => n21756, ZN => n13521);
   U30953 : INV_X2 port map( I => n39733, ZN => n39827);
   U30954 : XOR2_X1 port map( A1 => n19727, A2 => n9707, Z => n39733);
   U30955 : AOI21_X2 port map( A1 => n39735, A2 => n13030, B => n24727, ZN => 
                           n25186);
   U30956 : XOR2_X1 port map( A1 => n11416, A2 => n34181, Z => n11415);
   U30957 : BUF_X2 port map( I => n30284, Z => n39737);
   U30958 : NAND2_X2 port map( A1 => n39738, A2 => n7179, ZN => n16238);
   U30959 : AND2_X1 port map( A1 => n28339, A2 => n28400, Z => n13401);
   U30960 : NAND2_X2 port map( A1 => n33585, A2 => n33138, ZN => n23426);
   U30961 : NAND3_X2 port map( A1 => n39740, A2 => n30391, A3 => n28863, ZN => 
                           n29687);
   U30962 : XOR2_X1 port map( A1 => n39741, A2 => n27701, Z => n6644);
   U30963 : XOR2_X1 port map( A1 => n10057, A2 => n19612, Z => n39741);
   U30964 : XOR2_X1 port map( A1 => n29088, A2 => n12707, Z => n6635);
   U30965 : NAND2_X2 port map( A1 => n35776, A2 => n33686, ZN => n12707);
   U30966 : XOR2_X1 port map( A1 => n38041, A2 => n13147, Z => n39743);
   U30967 : NAND2_X2 port map( A1 => n36186, A2 => n36082, ZN => n30282);
   U30968 : NAND2_X2 port map( A1 => n4143, A2 => n121, ZN => n15559);
   U30969 : XOR2_X1 port map( A1 => n30819, A2 => n17328, Z => n39744);
   U30970 : BUF_X2 port map( I => n29996, Z => n39745);
   U30971 : XNOR2_X1 port map( A1 => n17398, A2 => n6142, ZN => n39783);
   U30972 : NAND3_X1 port map( A1 => n27934, A2 => n32977, A3 => n28118, ZN => 
                           n28347);
   U30973 : OAI21_X2 port map( A1 => n22036, A2 => n22037, B => n20388, ZN => 
                           n22509);
   U30974 : NAND2_X2 port map( A1 => n13241, A2 => n39746, ZN => n5061);
   U30975 : NOR2_X2 port map( A1 => n39747, A2 => n22091, ZN => n22014);
   U30976 : NOR3_X1 port map( A1 => n9685, A2 => n1678, A3 => n22204, ZN => 
                           n39747);
   U30977 : AOI22_X2 port map( A1 => n25364, A2 => n33114, B1 => n25366, B2 => 
                           n2576, ZN => n39748);
   U30978 : AND2_X1 port map( A1 => n16095, A2 => n33304, Z => n39749);
   U30979 : NAND2_X2 port map( A1 => n1116, A2 => n32868, ZN => n3451);
   U30980 : NAND2_X2 port map( A1 => n21565, A2 => n13472, ZN => n2166);
   U30981 : XOR2_X1 port map( A1 => n39750, A2 => n11284, Z => n17533);
   U30982 : XOR2_X1 port map( A1 => n39751, A2 => n9196, Z => n7741);
   U30983 : XOR2_X1 port map( A1 => n9195, A2 => n27795, Z => n39751);
   U30984 : OR3_X1 port map( A1 => n14369, A2 => n6106, A3 => n21301, Z => 
                           n25604);
   U30985 : BUF_X2 port map( I => n20267, Z => n39752);
   U30986 : XOR2_X1 port map( A1 => n35654, A2 => n2443, Z => n2714);
   U30987 : INV_X2 port map( I => n39753, ZN => n19016);
   U30988 : XOR2_X1 port map( A1 => Plaintext(44), A2 => Key(44), Z => n39753);
   U30989 : OAI21_X2 port map( A1 => n39754, A2 => n12405, B => n26794, ZN => 
                           n27304);
   U30990 : NOR2_X2 port map( A1 => n3041, A2 => n37589, ZN => n14429);
   U30991 : OAI21_X2 port map( A1 => n39755, A2 => n9170, B => n27893, ZN => 
                           n28704);
   U30992 : AOI21_X2 port map( A1 => n9168, A2 => n37015, B => n28419, ZN => 
                           n39755);
   U30993 : OAI21_X2 port map( A1 => n12352, A2 => n12214, B => n39757, ZN => 
                           n17884);
   U30994 : AOI22_X2 port map( A1 => n12213, A2 => n27306, B1 => n27585, B2 => 
                           n26791, ZN => n39757);
   U30995 : INV_X2 port map( I => n39759, ZN => n3452);
   U30996 : XNOR2_X1 port map( A1 => n22596, A2 => n22607, ZN => n39759);
   U30997 : OAI22_X1 port map( A1 => n1021, A2 => n2830, B1 => n15575, B2 => 
                           n17624, ZN => n2833);
   U30998 : INV_X2 port map( I => n23912, ZN => n39760);
   U30999 : INV_X2 port map( I => n28590, ZN => n39761);
   U31000 : INV_X2 port map( I => n5859, ZN => n31375);
   U31001 : NAND3_X2 port map( A1 => n5858, A2 => n5857, A3 => n12578, ZN => 
                           n5859);
   U31002 : XOR2_X1 port map( A1 => n39762, A2 => n1809, Z => n1805);
   U31003 : XOR2_X1 port map( A1 => n31012, A2 => n1807, Z => n39762);
   U31004 : XOR2_X1 port map( A1 => n17623, A2 => n39763, Z => n14953);
   U31005 : XOR2_X1 port map( A1 => n5208, A2 => n25115, Z => n39763);
   U31006 : XOR2_X1 port map( A1 => n39764, A2 => n22511, Z => n5340);
   U31007 : INV_X2 port map( I => n20335, ZN => n39764);
   U31008 : OAI22_X2 port map( A1 => n18392, A2 => n12260, B1 => n12257, B2 => 
                           n14451, ZN => n13409);
   U31009 : XOR2_X1 port map( A1 => n3290, A2 => n31125, Z => n755);
   U31010 : XOR2_X1 port map( A1 => n26397, A2 => n13064, Z => n39766);
   U31011 : XOR2_X1 port map( A1 => n28918, A2 => n28919, Z => n29903);
   U31012 : INV_X2 port map( I => n21644, ZN => n21909);
   U31013 : NAND2_X2 port map( A1 => n23608, A2 => n1637, ZN => n3744);
   U31014 : OAI21_X2 port map( A1 => n19869, A2 => n18850, B => n32013, ZN => 
                           n23608);
   U31015 : XOR2_X1 port map( A1 => n22640, A2 => n39767, Z => n35343);
   U31016 : XOR2_X1 port map( A1 => n12393, A2 => n35081, Z => n39767);
   U31017 : XOR2_X1 port map( A1 => n23902, A2 => n18849, Z => n6564);
   U31018 : NAND2_X1 port map( A1 => n29194, A2 => n29815, ZN => n39768);
   U31019 : NOR2_X1 port map( A1 => n19041, A2 => n29973, ZN => n29963);
   U31020 : INV_X2 port map( I => n10959, ZN => n11861);
   U31021 : INV_X1 port map( I => n26458, ZN => n26318);
   U31022 : XOR2_X1 port map( A1 => n26458, A2 => n17760, Z => n17759);
   U31023 : XOR2_X1 port map( A1 => n26365, A2 => n5031, Z => n26458);
   U31024 : INV_X2 port map( I => n19728, ZN => n19575);
   U31025 : NAND2_X2 port map( A1 => n39770, A2 => n23466, ZN => n2319);
   U31026 : OR2_X1 port map( A1 => n21546, A2 => n21871, Z => n11918);
   U31027 : XOR2_X1 port map( A1 => n4561, A2 => n4562, Z => n4564);
   U31028 : XOR2_X1 port map( A1 => n39772, A2 => n19616, Z => Ciphertext(85));
   U31029 : NAND2_X2 port map( A1 => n9884, A2 => n11001, ZN => n29683);
   U31030 : AOI22_X2 port map( A1 => n16367, A2 => n33349, B1 => n32616, B2 => 
                           n23556, ZN => n11529);
   U31031 : NAND2_X2 port map( A1 => n39773, A2 => n35159, ZN => n26161);
   U31032 : XOR2_X1 port map( A1 => n12818, A2 => n39774, Z => n4086);
   U31033 : XOR2_X1 port map( A1 => n7055, A2 => n27739, Z => n39774);
   U31034 : XOR2_X1 port map( A1 => n39775, A2 => n34136, Z => n35435);
   U31035 : NAND2_X2 port map( A1 => n37104, A2 => n33561, ZN => n13854);
   U31036 : INV_X2 port map( I => n1414, ZN => n4284);
   U31037 : XOR2_X1 port map( A1 => n39776, A2 => n8747, Z => n7459);
   U31038 : XOR2_X1 port map( A1 => n2283, A2 => n31909, Z => n39776);
   U31039 : OAI21_X2 port map( A1 => n2915, A2 => n12449, B => n12448, ZN => 
                           n6177);
   U31040 : NAND2_X2 port map( A1 => n24342, A2 => n24341, ZN => n30464);
   U31041 : XOR2_X1 port map( A1 => n18310, A2 => n16905, Z => n34518);
   U31042 : XOR2_X1 port map( A1 => n31401, A2 => n24941, Z => n39778);
   U31043 : XOR2_X1 port map( A1 => n22677, A2 => n22622, Z => n22592);
   U31044 : XOR2_X1 port map( A1 => n23971, A2 => n23974, Z => n11118);
   U31045 : XOR2_X1 port map( A1 => n18300, A2 => n23783, Z => n23971);
   U31046 : XOR2_X1 port map( A1 => n6369, A2 => n39779, Z => n19680);
   U31047 : XOR2_X1 port map( A1 => n22372, A2 => n6368, Z => n39779);
   U31048 : INV_X2 port map( I => n257, ZN => n8264);
   U31049 : NAND2_X2 port map( A1 => n15223, A2 => n16430, ZN => n257);
   U31050 : XOR2_X1 port map( A1 => n17651, A2 => n22383, Z => n8856);
   U31051 : OAI21_X2 port map( A1 => n37179, A2 => n3699, B => n2121, ZN => 
                           n9250);
   U31052 : XOR2_X1 port map( A1 => n25145, A2 => n25143, Z => n13260);
   U31053 : XOR2_X1 port map( A1 => n25097, A2 => n25211, Z => n25145);
   U31054 : NAND2_X1 port map( A1 => n34957, A2 => n26929, ZN => n26635);
   U31055 : NOR2_X2 port map( A1 => n39477, A2 => n31546, ZN => n26929);
   U31056 : XOR2_X1 port map( A1 => n27474, A2 => n15726, Z => n39780);
   U31057 : NOR2_X2 port map( A1 => n840, A2 => n11003, ZN => n31917);
   U31058 : AND3_X1 port map( A1 => n22326, A2 => n39489, A3 => n4108, Z => 
                           n36085);
   U31059 : NOR2_X1 port map( A1 => n21687, A2 => n21688, ZN => n21691);
   U31060 : INV_X2 port map( I => n9964, ZN => n21687);
   U31061 : XOR2_X1 port map( A1 => Plaintext(38), A2 => Key(38), Z => n9964);
   U31062 : XOR2_X1 port map( A1 => n39783, A2 => n9430, Z => n36113);
   U31063 : XOR2_X1 port map( A1 => n8473, A2 => n31591, Z => n8472);
   U31064 : NAND2_X2 port map( A1 => n16657, A2 => n16658, ZN => n8473);
   U31065 : NAND2_X2 port map( A1 => n39784, A2 => n33730, ZN => n7506);
   U31066 : NAND2_X2 port map( A1 => n2974, A2 => n2977, ZN => n39784);
   U31067 : NAND2_X2 port map( A1 => n39785, A2 => n10657, ZN => n22119);
   U31068 : XOR2_X1 port map( A1 => n22731, A2 => n31562, Z => n17413);
   U31069 : NOR2_X2 port map( A1 => n8503, A2 => n8504, ZN => n31562);
   U31070 : XOR2_X1 port map( A1 => n10520, A2 => n30094, Z => n642);
   U31071 : XOR2_X1 port map( A1 => n39790, A2 => n17834, Z => n17838);
   U31072 : XOR2_X1 port map( A1 => n18600, A2 => n25250, Z => n39790);
   U31073 : XOR2_X1 port map( A1 => n39791, A2 => n14505, Z => n779);
   U31074 : XOR2_X1 port map( A1 => n1324, A2 => n39792, Z => n39791);
   U31075 : INV_X2 port map( I => n8552, ZN => n39792);
   U31076 : NOR3_X2 port map( A1 => n16845, A2 => n14432, A3 => n29640, ZN => 
                           n19318);
   U31077 : XOR2_X1 port map( A1 => n32646, A2 => n1664, Z => n9511);
   U31078 : NOR2_X2 port map( A1 => n31966, A2 => n28109, ZN => n39794);
   U31079 : INV_X1 port map( I => n28240, ZN => n39795);
   U31080 : BUF_X2 port map( I => n7728, Z => n39797);
   U31081 : XOR2_X1 port map( A1 => n5279, A2 => n37197, Z => n12283);
   U31082 : XOR2_X1 port map( A1 => n22741, A2 => n1324, Z => n5279);
   U31083 : NOR2_X2 port map( A1 => n7391, A2 => n19813, ZN => n15635);
   U31084 : INV_X2 port map( I => n39799, ZN => n7391);
   U31085 : NOR2_X2 port map( A1 => n733, A2 => n33948, ZN => n39799);
   U31086 : OR2_X1 port map( A1 => n35757, A2 => n7459, Z => n8819);
   U31087 : XOR2_X1 port map( A1 => n35542, A2 => n14608, Z => n35757);
   U31088 : NAND2_X2 port map( A1 => n10152, A2 => n20313, ZN => n24162);
   U31089 : OAI22_X1 port map( A1 => n2866, A2 => n39392, B1 => n19544, B2 => 
                           n29059, ZN => n15492);
   U31090 : NOR2_X2 port map( A1 => n7789, A2 => n30240, ZN => n2866);
   U31091 : NAND2_X2 port map( A1 => n20875, A2 => n39802, ZN => n26089);
   U31092 : OAI21_X2 port map( A1 => n10532, A2 => n17282, B => n7236, ZN => 
                           n39802);
   U31093 : OR2_X1 port map( A1 => n35216, A2 => n32775, Z => n18207);
   U31094 : NAND2_X2 port map( A1 => n4083, A2 => n35551, ZN => n16672);
   U31095 : OAI21_X2 port map( A1 => n24187, A2 => n13167, B => n10659, ZN => 
                           n36664);
   U31096 : AOI22_X2 port map( A1 => n1133, A2 => n7885, B1 => n7886, B2 => 
                           n23504, ZN => n7884);
   U31097 : NAND2_X1 port map( A1 => n27269, A2 => n35990, ZN => n20377);
   U31098 : XOR2_X1 port map( A1 => n39807, A2 => n33695, Z => n20974);
   U31099 : XOR2_X1 port map( A1 => n34489, A2 => n26513, Z => n39807);
   U31100 : OAI22_X2 port map( A1 => n39808, A2 => n34790, B1 => n8342, B2 => 
                           n21995, ZN => n6893);
   U31101 : XOR2_X1 port map( A1 => n17569, A2 => n38216, Z => n39809);
   U31102 : INV_X2 port map( I => n7828, ZN => n21239);
   U31103 : INV_X2 port map( I => n17564, ZN => n23190);
   U31104 : INV_X1 port map( I => n38851, ZN => n22964);
   U31105 : INV_X2 port map( I => n22853, ZN => n14817);
   U31106 : OR2_X1 port map( A1 => n4600, A2 => n31611, Z => n39813);
   U31107 : AND2_X1 port map( A1 => n18907, A2 => n18402, Z => n39818);
   U31108 : BUF_X2 port map( I => n19223, Z => n14082);
   U31109 : INV_X2 port map( I => n9751, ZN => n36708);
   U31110 : XNOR2_X1 port map( A1 => n30910, A2 => n13260, ZN => n39820);
   U31111 : BUF_X2 port map( I => n6145, Z => n5314);
   U31112 : OAI22_X2 port map( A1 => n16073, A2 => n34436, B1 => n16072, B2 => 
                           n35160, ZN => n35207);
   U31113 : AOI22_X2 port map( A1 => n26097, A2 => n39351, B1 => n32748, B2 => 
                           n32747, ZN => n35238);
   U31114 : XNOR2_X1 port map( A1 => n15077, A2 => n15453, ZN => n39823);
   U31115 : INV_X2 port map( I => n28125, ZN => n10836);
   U31116 : OAI21_X2 port map( A1 => n5160, A2 => n5158, B => n31932, ZN => 
                           n6067);
   U31117 : INV_X2 port map( I => n13927, ZN => n18061);
   U31118 : INV_X2 port map( I => n3845, ZN => n31888);
   U31119 : INV_X2 port map( I => n34325, ZN => n777);
   U31120 : INV_X2 port map( I => n16803, ZN => n967);
   U31121 : XNOR2_X1 port map( A1 => n2996, A2 => n32092, ZN => n39828);
   U31122 : INV_X2 port map( I => n29184, ZN => n35551);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Top is

   port( clk : in std_logic;  Plaintext, Key : in std_logic_vector (191 downto 
         0);  Ciphertext : out std_logic_vector (191 downto 0));

end SPEEDY_Top;

architecture SYN_Behavioral of SPEEDY_Top is

   component DFFRNQ_X1
      port( D, CLK, RN : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSNQ_X1
      port( D, CLK, SN : in std_logic;  Q : out std_logic);
   end component;
   
   component SPEEDY_Rounds7_0
      port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : 
            out std_logic_vector (191 downto 0));
   end component;
   
   signal reg_in_191_port, reg_in_190_port, reg_in_189_port, reg_in_188_port, 
      reg_in_187_port, reg_in_186_port, reg_in_185_port, reg_in_184_port, 
      reg_in_183_port, reg_in_182_port, reg_in_181_port, reg_in_180_port, 
      reg_in_179_port, reg_in_178_port, reg_in_177_port, reg_in_176_port, 
      reg_in_175_port, reg_in_174_port, reg_in_173_port, reg_in_172_port, 
      reg_in_171_port, reg_in_170_port, reg_in_169_port, reg_in_168_port, 
      reg_in_167_port, reg_in_166_port, reg_in_165_port, reg_in_164_port, 
      reg_in_163_port, reg_in_162_port, reg_in_161_port, reg_in_160_port, 
      reg_in_159_port, reg_in_158_port, reg_in_157_port, reg_in_156_port, 
      reg_in_155_port, reg_in_154_port, reg_in_153_port, reg_in_152_port, 
      reg_in_151_port, reg_in_150_port, reg_in_149_port, reg_in_148_port, 
      reg_in_147_port, reg_in_146_port, reg_in_145_port, reg_in_144_port, 
      reg_in_143_port, reg_in_142_port, reg_in_141_port, reg_in_140_port, 
      reg_in_139_port, reg_in_138_port, reg_in_137_port, reg_in_136_port, 
      reg_in_135_port, reg_in_134_port, reg_in_133_port, reg_in_132_port, 
      reg_in_131_port, reg_in_130_port, reg_in_129_port, reg_in_128_port, 
      reg_in_127_port, reg_in_126_port, reg_in_125_port, reg_in_124_port, 
      reg_in_123_port, reg_in_122_port, reg_in_121_port, reg_in_120_port, 
      reg_in_119_port, reg_in_118_port, reg_in_117_port, reg_in_116_port, 
      reg_in_115_port, reg_in_114_port, reg_in_113_port, reg_in_112_port, 
      reg_in_111_port, reg_in_110_port, reg_in_109_port, reg_in_108_port, 
      reg_in_107_port, reg_in_106_port, reg_in_105_port, reg_in_104_port, 
      reg_in_103_port, reg_in_102_port, reg_in_101_port, reg_in_100_port, 
      reg_in_99_port, reg_in_98_port, reg_in_97_port, reg_in_96_port, 
      reg_in_95_port, reg_in_94_port, reg_in_93_port, reg_in_92_port, 
      reg_in_91_port, reg_in_90_port, reg_in_89_port, reg_in_88_port, 
      reg_in_87_port, reg_in_86_port, reg_in_85_port, reg_in_84_port, 
      reg_in_83_port, reg_in_82_port, reg_in_81_port, reg_in_80_port, 
      reg_in_79_port, reg_in_78_port, reg_in_77_port, reg_in_76_port, 
      reg_in_75_port, reg_in_74_port, reg_in_73_port, reg_in_72_port, 
      reg_in_71_port, reg_in_70_port, reg_in_69_port, reg_in_68_port, 
      reg_in_67_port, reg_in_66_port, reg_in_65_port, reg_in_64_port, 
      reg_in_63_port, reg_in_62_port, reg_in_61_port, reg_in_60_port, 
      reg_in_59_port, reg_in_58_port, reg_in_57_port, reg_in_56_port, 
      reg_in_55_port, reg_in_54_port, reg_in_53_port, reg_in_52_port, 
      reg_in_51_port, reg_in_50_port, reg_in_49_port, reg_in_48_port, 
      reg_in_47_port, reg_in_46_port, reg_in_45_port, reg_in_44_port, 
      reg_in_43_port, reg_in_42_port, reg_in_41_port, reg_in_40_port, 
      reg_in_39_port, reg_in_38_port, reg_in_37_port, reg_in_36_port, 
      reg_in_35_port, reg_in_34_port, reg_in_33_port, reg_in_32_port, 
      reg_in_31_port, reg_in_30_port, reg_in_29_port, reg_in_28_port, 
      reg_in_27_port, reg_in_26_port, reg_in_25_port, reg_in_24_port, 
      reg_in_23_port, reg_in_22_port, reg_in_21_port, reg_in_20_port, 
      reg_in_19_port, reg_in_18_port, reg_in_17_port, reg_in_16_port, 
      reg_in_15_port, reg_in_14_port, reg_in_13_port, reg_in_12_port, 
      reg_in_11_port, reg_in_10_port, reg_in_9_port, reg_in_8_port, 
      reg_in_7_port, reg_in_6_port, reg_in_5_port, reg_in_4_port, reg_in_3_port
      , reg_in_2_port, reg_in_1_port, reg_in_0_port, reg_key_191_port, 
      reg_key_190_port, reg_key_189_port, reg_key_188_port, reg_key_187_port, 
      reg_key_186_port, reg_key_185_port, reg_key_184_port, reg_key_183_port, 
      reg_key_182_port, reg_key_181_port, reg_key_180_port, reg_key_179_port, 
      reg_key_178_port, reg_key_177_port, reg_key_176_port, reg_key_175_port, 
      reg_key_174_port, reg_key_173_port, reg_key_172_port, reg_key_171_port, 
      reg_key_170_port, reg_key_169_port, reg_key_168_port, reg_key_167_port, 
      reg_key_166_port, reg_key_165_port, reg_key_164_port, reg_key_163_port, 
      reg_key_162_port, reg_key_161_port, reg_key_160_port, reg_key_159_port, 
      reg_key_158_port, reg_key_157_port, reg_key_156_port, reg_key_155_port, 
      reg_key_154_port, reg_key_153_port, reg_key_152_port, reg_key_151_port, 
      reg_key_150_port, reg_key_149_port, reg_key_148_port, reg_key_147_port, 
      reg_key_146_port, reg_key_145_port, reg_key_144_port, reg_key_143_port, 
      reg_key_142_port, reg_key_141_port, reg_key_140_port, reg_key_139_port, 
      reg_key_138_port, reg_key_137_port, reg_key_136_port, reg_key_135_port, 
      reg_key_134_port, reg_key_133_port, reg_key_132_port, reg_key_131_port, 
      reg_key_130_port, reg_key_129_port, reg_key_128_port, reg_key_127_port, 
      reg_key_126_port, reg_key_125_port, reg_key_124_port, reg_key_123_port, 
      reg_key_122_port, reg_key_121_port, reg_key_120_port, reg_key_119_port, 
      reg_key_118_port, reg_key_117_port, reg_key_116_port, reg_key_115_port, 
      reg_key_114_port, reg_key_113_port, reg_key_112_port, reg_key_111_port, 
      reg_key_110_port, reg_key_109_port, reg_key_108_port, reg_key_107_port, 
      reg_key_106_port, reg_key_105_port, reg_key_104_port, reg_key_103_port, 
      reg_key_102_port, reg_key_101_port, reg_key_100_port, reg_key_99_port, 
      reg_key_98_port, reg_key_97_port, reg_key_96_port, reg_key_95_port, 
      reg_key_94_port, reg_key_93_port, reg_key_92_port, reg_key_91_port, 
      reg_key_90_port, reg_key_89_port, reg_key_88_port, reg_key_87_port, 
      reg_key_86_port, reg_key_85_port, reg_key_84_port, reg_key_83_port, 
      reg_key_82_port, reg_key_81_port, reg_key_80_port, reg_key_79_port, 
      reg_key_78_port, reg_key_77_port, reg_key_76_port, reg_key_75_port, 
      reg_key_74_port, reg_key_73_port, reg_key_72_port, reg_key_71_port, 
      reg_key_70_port, reg_key_69_port, reg_key_68_port, reg_key_67_port, 
      reg_key_66_port, reg_key_65_port, reg_key_64_port, reg_key_63_port, 
      reg_key_62_port, reg_key_61_port, reg_key_60_port, reg_key_59_port, 
      reg_key_58_port, reg_key_57_port, reg_key_56_port, reg_key_55_port, 
      reg_key_54_port, reg_key_53_port, reg_key_52_port, reg_key_51_port, 
      reg_key_50_port, reg_key_49_port, reg_key_48_port, reg_key_47_port, 
      reg_key_46_port, reg_key_45_port, reg_key_44_port, reg_key_43_port, 
      reg_key_42_port, reg_key_41_port, reg_key_40_port, reg_key_39_port, 
      reg_key_38_port, reg_key_37_port, reg_key_36_port, reg_key_35_port, 
      reg_key_34_port, reg_key_33_port, reg_key_32_port, reg_key_31_port, 
      reg_key_30_port, reg_key_29_port, reg_key_28_port, reg_key_27_port, 
      reg_key_26_port, reg_key_25_port, reg_key_24_port, reg_key_23_port, 
      reg_key_22_port, reg_key_21_port, reg_key_20_port, reg_key_19_port, 
      reg_key_18_port, reg_key_17_port, reg_key_16_port, reg_key_15_port, 
      reg_key_14_port, reg_key_13_port, reg_key_12_port, reg_key_11_port, 
      reg_key_10_port, reg_key_9_port, reg_key_8_port, reg_key_7_port, 
      reg_key_6_port, reg_key_5_port, reg_key_4_port, reg_key_3_port, 
      reg_key_2_port, reg_key_1_port, reg_key_0_port, reg_out_191_port, 
      reg_out_190_port, reg_out_189_port, reg_out_188_port, reg_out_187_port, 
      reg_out_186_port, reg_out_185_port, reg_out_184_port, reg_out_183_port, 
      reg_out_182_port, reg_out_181_port, reg_out_180_port, reg_out_179_port, 
      reg_out_178_port, reg_out_177_port, reg_out_176_port, reg_out_175_port, 
      reg_out_174_port, reg_out_173_port, reg_out_172_port, reg_out_171_port, 
      reg_out_170_port, reg_out_169_port, reg_out_168_port, reg_out_167_port, 
      reg_out_166_port, reg_out_165_port, reg_out_164_port, reg_out_163_port, 
      reg_out_162_port, reg_out_161_port, reg_out_160_port, reg_out_159_port, 
      reg_out_158_port, reg_out_157_port, reg_out_156_port, reg_out_155_port, 
      reg_out_154_port, reg_out_153_port, reg_out_152_port, reg_out_151_port, 
      reg_out_150_port, reg_out_149_port, reg_out_148_port, reg_out_147_port, 
      reg_out_146_port, reg_out_145_port, reg_out_144_port, reg_out_143_port, 
      reg_out_142_port, reg_out_141_port, reg_out_140_port, reg_out_139_port, 
      reg_out_138_port, reg_out_137_port, reg_out_136_port, reg_out_135_port, 
      reg_out_134_port, reg_out_133_port, reg_out_132_port, reg_out_131_port, 
      reg_out_130_port, reg_out_129_port, reg_out_128_port, reg_out_127_port, 
      reg_out_126_port, reg_out_125_port, reg_out_124_port, reg_out_123_port, 
      reg_out_122_port, reg_out_121_port, reg_out_120_port, reg_out_119_port, 
      reg_out_118_port, reg_out_117_port, reg_out_116_port, reg_out_115_port, 
      reg_out_114_port, reg_out_113_port, reg_out_112_port, reg_out_111_port, 
      reg_out_110_port, reg_out_109_port, reg_out_108_port, reg_out_107_port, 
      reg_out_106_port, reg_out_105_port, reg_out_104_port, reg_out_103_port, 
      reg_out_102_port, reg_out_101_port, reg_out_100_port, reg_out_99_port, 
      reg_out_98_port, reg_out_97_port, reg_out_96_port, reg_out_95_port, 
      reg_out_94_port, reg_out_93_port, reg_out_92_port, reg_out_91_port, 
      reg_out_90_port, reg_out_89_port, reg_out_88_port, reg_out_87_port, 
      reg_out_86_port, reg_out_85_port, reg_out_84_port, reg_out_83_port, 
      reg_out_82_port, reg_out_81_port, reg_out_80_port, reg_out_79_port, 
      reg_out_78_port, reg_out_77_port, reg_out_76_port, reg_out_75_port, 
      reg_out_74_port, reg_out_73_port, reg_out_72_port, reg_out_71_port, 
      reg_out_70_port, reg_out_69_port, reg_out_68_port, reg_out_67_port, 
      reg_out_66_port, reg_out_65_port, reg_out_64_port, reg_out_63_port, 
      reg_out_62_port, reg_out_61_port, reg_out_60_port, reg_out_59_port, 
      reg_out_58_port, reg_out_57_port, reg_out_56_port, reg_out_55_port, 
      reg_out_54_port, reg_out_53_port, reg_out_52_port, reg_out_51_port, 
      reg_out_50_port, reg_out_49_port, reg_out_48_port, reg_out_47_port, 
      reg_out_46_port, reg_out_45_port, reg_out_44_port, reg_out_43_port, 
      reg_out_42_port, reg_out_41_port, reg_out_40_port, reg_out_39_port, 
      reg_out_38_port, reg_out_37_port, reg_out_36_port, reg_out_35_port, 
      reg_out_34_port, reg_out_33_port, reg_out_32_port, reg_out_31_port, 
      reg_out_30_port, reg_out_29_port, reg_out_28_port, reg_out_27_port, 
      reg_out_26_port, reg_out_25_port, reg_out_24_port, reg_out_23_port, 
      reg_out_22_port, reg_out_21_port, reg_out_20_port, reg_out_19_port, 
      reg_out_18_port, reg_out_17_port, reg_out_16_port, reg_out_15_port, 
      reg_out_14_port, reg_out_13_port, reg_out_12_port, reg_out_11_port, 
      reg_out_10_port, reg_out_9_port, reg_out_8_port, reg_out_7_port, 
      reg_out_6_port, reg_out_5_port, reg_out_4_port, reg_out_3_port, 
      reg_out_2_port, reg_out_1_port, reg_out_0_port, n2, n3, n5, n6, n7, n8, 
      n12, n13, n14, n16, n17, n18, n19, n20, n23, n25, n26, n28, n30, n32, n35
      , n36, n37, n38, n39, n41, n42, n43, n44, n45, n46, n47, n48, n49, n51, 
      n52, n53, n54, n56, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71
      , n72, n74, n75, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, 
      n90, n91, n92, n93, n94, n97, n99, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n113, n114, n116, n119, n120, n122, n123, n124, n127, 
      n128, n129, n130, n135, n136, n139, n140, n141, n142, n143, n145, n146, 
      n148, n149, n150, n151, n152, n156, n157, n158, n159, n162, n164, n167, 
      n168, n169, n171, n173, n174, n176, n177, n178, n179, n180, n182, n184, 
      n185, n188, n189, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
      n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, 
      n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n345, n346, 
      n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, 
      n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
      n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
      n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
      n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, 
      n407, n408, n409, n413, n415, n416, n417, n418, n419, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n469, n470, n471, n472, n473, 
      n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, 
      n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, 
      n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n526, n527, n528, n529, n530, n532, n533, n534, n535, n536, 
      n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, 
      n549, n550, n551, n552, n553, n555, n556, n557, n558, n559, n560, n561, 
      n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, 
      n574, n575, n577, n578, n579, n580, n581, n582, n583, n584, n586, n587, 
      n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
      n600, n601, n602, n603, n604, n605, n606, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, 
      n625, n626, n627, n628, n629, n630, n631, n632, n633, n635, n636, n637, 
      n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, 
      n650, n651, n652, n653, n654, n655, n656 : std_logic;

begin
   
   reg_in_regx190x : DFFSNQ_X1 port map( D => Plaintext(190), CLK => clk, SN =>
                           n575, Q => reg_in_190_port);
   reg_in_regx189x : DFFSNQ_X1 port map( D => Plaintext(189), CLK => clk, SN =>
                           n574, Q => reg_in_189_port);
   reg_in_regx188x : DFFSNQ_X1 port map( D => Plaintext(188), CLK => clk, SN =>
                           n573, Q => reg_in_188_port);
   reg_in_regx187x : DFFSNQ_X1 port map( D => Plaintext(187), CLK => clk, SN =>
                           n572, Q => reg_in_187_port);
   reg_in_regx186x : DFFSNQ_X1 port map( D => Plaintext(186), CLK => clk, SN =>
                           n571, Q => reg_in_186_port);
   reg_in_regx185x : DFFSNQ_X1 port map( D => Plaintext(185), CLK => clk, SN =>
                           n570, Q => reg_in_185_port);
   reg_in_regx184x : DFFSNQ_X1 port map( D => Plaintext(184), CLK => clk, SN =>
                           n569, Q => reg_in_184_port);
   reg_in_regx183x : DFFSNQ_X1 port map( D => Plaintext(183), CLK => clk, SN =>
                           n568, Q => reg_in_183_port);
   reg_in_regx182x : DFFSNQ_X1 port map( D => Plaintext(182), CLK => clk, SN =>
                           n567, Q => reg_in_182_port);
   reg_in_regx181x : DFFSNQ_X1 port map( D => Plaintext(181), CLK => clk, SN =>
                           n566, Q => reg_in_181_port);
   reg_in_regx180x : DFFSNQ_X1 port map( D => Plaintext(180), CLK => clk, SN =>
                           n565, Q => reg_in_180_port);
   reg_in_regx179x : DFFSNQ_X1 port map( D => Plaintext(179), CLK => clk, SN =>
                           n564, Q => reg_in_179_port);
   reg_in_regx178x : DFFSNQ_X1 port map( D => Plaintext(178), CLK => clk, SN =>
                           n563, Q => reg_in_178_port);
   reg_in_regx177x : DFFSNQ_X1 port map( D => Plaintext(177), CLK => clk, SN =>
                           n562, Q => reg_in_177_port);
   reg_in_regx176x : DFFSNQ_X1 port map( D => Plaintext(176), CLK => clk, SN =>
                           n561, Q => reg_in_176_port);
   reg_in_regx175x : DFFSNQ_X1 port map( D => Plaintext(175), CLK => clk, SN =>
                           n560, Q => reg_in_175_port);
   reg_in_regx174x : DFFSNQ_X1 port map( D => Plaintext(174), CLK => clk, SN =>
                           n559, Q => reg_in_174_port);
   reg_in_regx173x : DFFSNQ_X1 port map( D => Plaintext(173), CLK => clk, SN =>
                           n558, Q => reg_in_173_port);
   reg_in_regx172x : DFFSNQ_X1 port map( D => Plaintext(172), CLK => clk, SN =>
                           n557, Q => reg_in_172_port);
   reg_in_regx171x : DFFSNQ_X1 port map( D => Plaintext(171), CLK => clk, SN =>
                           n556, Q => reg_in_171_port);
   reg_in_regx170x : DFFSNQ_X1 port map( D => Plaintext(170), CLK => clk, SN =>
                           n555, Q => reg_in_170_port);
   reg_in_regx168x : DFFSNQ_X1 port map( D => Plaintext(168), CLK => clk, SN =>
                           n553, Q => reg_in_168_port);
   reg_in_regx167x : DFFSNQ_X1 port map( D => Plaintext(167), CLK => clk, SN =>
                           n552, Q => reg_in_167_port);
   reg_in_regx166x : DFFSNQ_X1 port map( D => Plaintext(166), CLK => clk, SN =>
                           n551, Q => reg_in_166_port);
   reg_in_regx165x : DFFSNQ_X1 port map( D => Plaintext(165), CLK => clk, SN =>
                           n550, Q => reg_in_165_port);
   reg_in_regx164x : DFFSNQ_X1 port map( D => Plaintext(164), CLK => clk, SN =>
                           n549, Q => reg_in_164_port);
   reg_in_regx163x : DFFSNQ_X1 port map( D => Plaintext(163), CLK => clk, SN =>
                           n548, Q => reg_in_163_port);
   reg_in_regx162x : DFFSNQ_X1 port map( D => Plaintext(162), CLK => clk, SN =>
                           n547, Q => reg_in_162_port);
   reg_in_regx161x : DFFSNQ_X1 port map( D => Plaintext(161), CLK => clk, SN =>
                           n546, Q => reg_in_161_port);
   reg_in_regx160x : DFFSNQ_X1 port map( D => Plaintext(160), CLK => clk, SN =>
                           n545, Q => reg_in_160_port);
   reg_in_regx159x : DFFSNQ_X1 port map( D => Plaintext(159), CLK => clk, SN =>
                           n544, Q => reg_in_159_port);
   reg_in_regx158x : DFFSNQ_X1 port map( D => Plaintext(158), CLK => clk, SN =>
                           n543, Q => reg_in_158_port);
   reg_in_regx157x : DFFSNQ_X1 port map( D => Plaintext(157), CLK => clk, SN =>
                           n542, Q => reg_in_157_port);
   reg_in_regx156x : DFFSNQ_X1 port map( D => Plaintext(156), CLK => clk, SN =>
                           n541, Q => reg_in_156_port);
   reg_in_regx155x : DFFSNQ_X1 port map( D => Plaintext(155), CLK => clk, SN =>
                           n540, Q => reg_in_155_port);
   reg_in_regx154x : DFFSNQ_X1 port map( D => Plaintext(154), CLK => clk, SN =>
                           n539, Q => reg_in_154_port);
   reg_in_regx153x : DFFSNQ_X1 port map( D => Plaintext(153), CLK => clk, SN =>
                           n538, Q => reg_in_153_port);
   reg_in_regx152x : DFFSNQ_X1 port map( D => Plaintext(152), CLK => clk, SN =>
                           n537, Q => reg_in_152_port);
   reg_in_regx151x : DFFSNQ_X1 port map( D => Plaintext(151), CLK => clk, SN =>
                           n536, Q => reg_in_151_port);
   reg_in_regx150x : DFFSNQ_X1 port map( D => Plaintext(150), CLK => clk, SN =>
                           n535, Q => reg_in_150_port);
   reg_in_regx149x : DFFSNQ_X1 port map( D => Plaintext(149), CLK => clk, SN =>
                           n534, Q => reg_in_149_port);
   reg_in_regx148x : DFFSNQ_X1 port map( D => Plaintext(148), CLK => clk, SN =>
                           n533, Q => reg_in_148_port);
   reg_in_regx147x : DFFSNQ_X1 port map( D => Plaintext(147), CLK => clk, SN =>
                           n532, Q => reg_in_147_port);
   reg_in_regx145x : DFFSNQ_X1 port map( D => Plaintext(145), CLK => clk, SN =>
                           n530, Q => reg_in_145_port);
   reg_in_regx144x : DFFSNQ_X1 port map( D => Plaintext(144), CLK => clk, SN =>
                           n529, Q => reg_in_144_port);
   reg_in_regx143x : DFFSNQ_X1 port map( D => Plaintext(143), CLK => clk, SN =>
                           n528, Q => reg_in_143_port);
   reg_in_regx142x : DFFSNQ_X1 port map( D => Plaintext(142), CLK => clk, SN =>
                           n527, Q => reg_in_142_port);
   reg_in_regx141x : DFFSNQ_X1 port map( D => Plaintext(141), CLK => clk, SN =>
                           n526, Q => reg_in_141_port);
   reg_in_regx139x : DFFSNQ_X1 port map( D => Plaintext(139), CLK => clk, SN =>
                           n524, Q => reg_in_139_port);
   reg_in_regx138x : DFFSNQ_X1 port map( D => Plaintext(138), CLK => clk, SN =>
                           n523, Q => reg_in_138_port);
   reg_in_regx137x : DFFSNQ_X1 port map( D => Plaintext(137), CLK => clk, SN =>
                           n522, Q => reg_in_137_port);
   reg_in_regx136x : DFFSNQ_X1 port map( D => Plaintext(136), CLK => clk, SN =>
                           n521, Q => reg_in_136_port);
   reg_in_regx135x : DFFSNQ_X1 port map( D => Plaintext(135), CLK => clk, SN =>
                           n520, Q => reg_in_135_port);
   reg_in_regx134x : DFFSNQ_X1 port map( D => Plaintext(134), CLK => clk, SN =>
                           n519, Q => reg_in_134_port);
   reg_in_regx133x : DFFSNQ_X1 port map( D => Plaintext(133), CLK => clk, SN =>
                           n518, Q => reg_in_133_port);
   reg_in_regx132x : DFFSNQ_X1 port map( D => Plaintext(132), CLK => clk, SN =>
                           n517, Q => reg_in_132_port);
   reg_in_regx131x : DFFSNQ_X1 port map( D => Plaintext(131), CLK => clk, SN =>
                           n516, Q => reg_in_131_port);
   reg_in_regx130x : DFFSNQ_X1 port map( D => Plaintext(130), CLK => clk, SN =>
                           n515, Q => reg_in_130_port);
   reg_in_regx129x : DFFSNQ_X1 port map( D => Plaintext(129), CLK => clk, SN =>
                           n514, Q => reg_in_129_port);
   reg_in_regx128x : DFFSNQ_X1 port map( D => Plaintext(128), CLK => clk, SN =>
                           n513, Q => reg_in_128_port);
   reg_in_regx127x : DFFSNQ_X1 port map( D => Plaintext(127), CLK => clk, SN =>
                           n512, Q => reg_in_127_port);
   reg_in_regx126x : DFFSNQ_X1 port map( D => Plaintext(126), CLK => clk, SN =>
                           n511, Q => reg_in_126_port);
   reg_in_regx124x : DFFSNQ_X1 port map( D => Plaintext(124), CLK => clk, SN =>
                           n509, Q => reg_in_124_port);
   reg_in_regx123x : DFFSNQ_X1 port map( D => Plaintext(123), CLK => clk, SN =>
                           n508, Q => reg_in_123_port);
   reg_in_regx122x : DFFSNQ_X1 port map( D => Plaintext(122), CLK => clk, SN =>
                           n507, Q => reg_in_122_port);
   reg_in_regx121x : DFFSNQ_X1 port map( D => Plaintext(121), CLK => clk, SN =>
                           n506, Q => reg_in_121_port);
   reg_in_regx120x : DFFSNQ_X1 port map( D => Plaintext(120), CLK => clk, SN =>
                           n505, Q => reg_in_120_port);
   reg_in_regx119x : DFFSNQ_X1 port map( D => Plaintext(119), CLK => clk, SN =>
                           n504, Q => reg_in_119_port);
   reg_in_regx118x : DFFSNQ_X1 port map( D => Plaintext(118), CLK => clk, SN =>
                           n503, Q => reg_in_118_port);
   reg_in_regx117x : DFFSNQ_X1 port map( D => Plaintext(117), CLK => clk, SN =>
                           n502, Q => reg_in_117_port);
   reg_in_regx116x : DFFSNQ_X1 port map( D => Plaintext(116), CLK => clk, SN =>
                           n501, Q => reg_in_116_port);
   reg_in_regx115x : DFFSNQ_X1 port map( D => Plaintext(115), CLK => clk, SN =>
                           n500, Q => reg_in_115_port);
   reg_in_regx114x : DFFSNQ_X1 port map( D => Plaintext(114), CLK => clk, SN =>
                           n499, Q => reg_in_114_port);
   reg_in_regx113x : DFFSNQ_X1 port map( D => Plaintext(113), CLK => clk, SN =>
                           n498, Q => reg_in_113_port);
   reg_in_regx112x : DFFSNQ_X1 port map( D => Plaintext(112), CLK => clk, SN =>
                           n497, Q => reg_in_112_port);
   reg_in_regx111x : DFFSNQ_X1 port map( D => Plaintext(111), CLK => clk, SN =>
                           n496, Q => reg_in_111_port);
   reg_in_regx110x : DFFSNQ_X1 port map( D => Plaintext(110), CLK => clk, SN =>
                           n495, Q => reg_in_110_port);
   reg_in_regx109x : DFFSNQ_X1 port map( D => Plaintext(109), CLK => clk, SN =>
                           n494, Q => reg_in_109_port);
   reg_in_regx108x : DFFSNQ_X1 port map( D => Plaintext(108), CLK => clk, SN =>
                           n493, Q => reg_in_108_port);
   reg_in_regx107x : DFFSNQ_X1 port map( D => Plaintext(107), CLK => clk, SN =>
                           n492, Q => reg_in_107_port);
   reg_in_regx106x : DFFSNQ_X1 port map( D => Plaintext(106), CLK => clk, SN =>
                           n491, Q => reg_in_106_port);
   reg_in_regx105x : DFFSNQ_X1 port map( D => Plaintext(105), CLK => clk, SN =>
                           n490, Q => reg_in_105_port);
   reg_in_regx104x : DFFSNQ_X1 port map( D => Plaintext(104), CLK => clk, SN =>
                           n489, Q => reg_in_104_port);
   reg_in_regx103x : DFFSNQ_X1 port map( D => Plaintext(103), CLK => clk, SN =>
                           n488, Q => reg_in_103_port);
   reg_in_regx102x : DFFSNQ_X1 port map( D => Plaintext(102), CLK => clk, SN =>
                           n487, Q => reg_in_102_port);
   reg_in_regx101x : DFFSNQ_X1 port map( D => Plaintext(101), CLK => clk, SN =>
                           n486, Q => reg_in_101_port);
   reg_in_regx100x : DFFSNQ_X1 port map( D => Plaintext(100), CLK => clk, SN =>
                           n485, Q => reg_in_100_port);
   reg_in_regx99x : DFFSNQ_X1 port map( D => Plaintext(99), CLK => clk, SN => 
                           n484, Q => reg_in_99_port);
   reg_in_regx98x : DFFSNQ_X1 port map( D => Plaintext(98), CLK => clk, SN => 
                           n483, Q => reg_in_98_port);
   reg_in_regx97x : DFFSNQ_X1 port map( D => Plaintext(97), CLK => clk, SN => 
                           n482, Q => reg_in_97_port);
   reg_in_regx96x : DFFSNQ_X1 port map( D => Plaintext(96), CLK => clk, SN => 
                           n481, Q => reg_in_96_port);
   reg_in_regx95x : DFFSNQ_X1 port map( D => Plaintext(95), CLK => clk, SN => 
                           n480, Q => reg_in_95_port);
   reg_in_regx94x : DFFSNQ_X1 port map( D => Plaintext(94), CLK => clk, SN => 
                           n479, Q => reg_in_94_port);
   reg_in_regx93x : DFFSNQ_X1 port map( D => Plaintext(93), CLK => clk, SN => 
                           n478, Q => reg_in_93_port);
   reg_in_regx92x : DFFSNQ_X1 port map( D => Plaintext(92), CLK => clk, SN => 
                           n477, Q => reg_in_92_port);
   reg_in_regx91x : DFFSNQ_X1 port map( D => Plaintext(91), CLK => clk, SN => 
                           n476, Q => reg_in_91_port);
   reg_in_regx90x : DFFSNQ_X1 port map( D => Plaintext(90), CLK => clk, SN => 
                           n475, Q => reg_in_90_port);
   reg_in_regx89x : DFFSNQ_X1 port map( D => Plaintext(89), CLK => clk, SN => 
                           n474, Q => reg_in_89_port);
   reg_in_regx88x : DFFSNQ_X1 port map( D => Plaintext(88), CLK => clk, SN => 
                           n473, Q => reg_in_88_port);
   reg_in_regx87x : DFFSNQ_X1 port map( D => Plaintext(87), CLK => clk, SN => 
                           n472, Q => reg_in_87_port);
   reg_in_regx86x : DFFSNQ_X1 port map( D => Plaintext(86), CLK => clk, SN => 
                           n471, Q => reg_in_86_port);
   reg_in_regx85x : DFFSNQ_X1 port map( D => Plaintext(85), CLK => clk, SN => 
                           n470, Q => reg_in_85_port);
   reg_in_regx84x : DFFSNQ_X1 port map( D => Plaintext(84), CLK => clk, SN => 
                           n469, Q => reg_in_84_port);
   reg_in_regx82x : DFFSNQ_X1 port map( D => Plaintext(82), CLK => clk, SN => 
                           n467, Q => reg_in_82_port);
   reg_in_regx81x : DFFSNQ_X1 port map( D => Plaintext(81), CLK => clk, SN => 
                           n466, Q => reg_in_81_port);
   reg_in_regx80x : DFFSNQ_X1 port map( D => Plaintext(80), CLK => clk, SN => 
                           n465, Q => reg_in_80_port);
   reg_in_regx79x : DFFSNQ_X1 port map( D => Plaintext(79), CLK => clk, SN => 
                           n464, Q => reg_in_79_port);
   reg_in_regx78x : DFFSNQ_X1 port map( D => Plaintext(78), CLK => clk, SN => 
                           n463, Q => reg_in_78_port);
   reg_in_regx77x : DFFSNQ_X1 port map( D => Plaintext(77), CLK => clk, SN => 
                           n462, Q => reg_in_77_port);
   reg_in_regx76x : DFFSNQ_X1 port map( D => Plaintext(76), CLK => clk, SN => 
                           n461, Q => reg_in_76_port);
   reg_in_regx75x : DFFSNQ_X1 port map( D => Plaintext(75), CLK => clk, SN => 
                           n460, Q => reg_in_75_port);
   reg_in_regx74x : DFFSNQ_X1 port map( D => Plaintext(74), CLK => clk, SN => 
                           n459, Q => reg_in_74_port);
   reg_in_regx73x : DFFSNQ_X1 port map( D => Plaintext(73), CLK => clk, SN => 
                           n458, Q => reg_in_73_port);
   reg_in_regx72x : DFFSNQ_X1 port map( D => Plaintext(72), CLK => clk, SN => 
                           n457, Q => reg_in_72_port);
   reg_in_regx71x : DFFSNQ_X1 port map( D => Plaintext(71), CLK => clk, SN => 
                           n456, Q => reg_in_71_port);
   reg_in_regx70x : DFFSNQ_X1 port map( D => Plaintext(70), CLK => clk, SN => 
                           n455, Q => reg_in_70_port);
   reg_in_regx69x : DFFSNQ_X1 port map( D => Plaintext(69), CLK => clk, SN => 
                           n454, Q => reg_in_69_port);
   reg_in_regx68x : DFFSNQ_X1 port map( D => Plaintext(68), CLK => clk, SN => 
                           n453, Q => reg_in_68_port);
   reg_in_regx67x : DFFSNQ_X1 port map( D => Plaintext(67), CLK => clk, SN => 
                           n452, Q => reg_in_67_port);
   reg_in_regx66x : DFFSNQ_X1 port map( D => Plaintext(66), CLK => clk, SN => 
                           n451, Q => reg_in_66_port);
   reg_in_regx65x : DFFSNQ_X1 port map( D => Plaintext(65), CLK => clk, SN => 
                           n450, Q => reg_in_65_port);
   reg_in_regx64x : DFFSNQ_X1 port map( D => Plaintext(64), CLK => clk, SN => 
                           n449, Q => reg_in_64_port);
   reg_in_regx63x : DFFSNQ_X1 port map( D => Plaintext(63), CLK => clk, SN => 
                           n448, Q => reg_in_63_port);
   reg_in_regx62x : DFFSNQ_X1 port map( D => Plaintext(62), CLK => clk, SN => 
                           n447, Q => reg_in_62_port);
   reg_in_regx61x : DFFSNQ_X1 port map( D => Plaintext(61), CLK => clk, SN => 
                           n446, Q => reg_in_61_port);
   reg_in_regx60x : DFFSNQ_X1 port map( D => Plaintext(60), CLK => clk, SN => 
                           n445, Q => reg_in_60_port);
   reg_in_regx58x : DFFSNQ_X1 port map( D => Plaintext(58), CLK => clk, SN => 
                           n443, Q => reg_in_58_port);
   reg_in_regx57x : DFFSNQ_X1 port map( D => Plaintext(57), CLK => clk, SN => 
                           n442, Q => reg_in_57_port);
   reg_in_regx56x : DFFSNQ_X1 port map( D => Plaintext(56), CLK => clk, SN => 
                           n441, Q => reg_in_56_port);
   reg_in_regx55x : DFFSNQ_X1 port map( D => Plaintext(55), CLK => clk, SN => 
                           n440, Q => reg_in_55_port);
   reg_in_regx54x : DFFSNQ_X1 port map( D => Plaintext(54), CLK => clk, SN => 
                           n439, Q => reg_in_54_port);
   reg_in_regx53x : DFFSNQ_X1 port map( D => Plaintext(53), CLK => clk, SN => 
                           n438, Q => reg_in_53_port);
   reg_in_regx52x : DFFSNQ_X1 port map( D => Plaintext(52), CLK => clk, SN => 
                           n437, Q => reg_in_52_port);
   reg_in_regx51x : DFFSNQ_X1 port map( D => Plaintext(51), CLK => clk, SN => 
                           n436, Q => reg_in_51_port);
   reg_in_regx50x : DFFSNQ_X1 port map( D => Plaintext(50), CLK => clk, SN => 
                           n435, Q => reg_in_50_port);
   reg_in_regx49x : DFFSNQ_X1 port map( D => Plaintext(49), CLK => clk, SN => 
                           n434, Q => reg_in_49_port);
   reg_in_regx48x : DFFSNQ_X1 port map( D => Plaintext(48), CLK => clk, SN => 
                           n433, Q => reg_in_48_port);
   reg_in_regx47x : DFFSNQ_X1 port map( D => Plaintext(47), CLK => clk, SN => 
                           n432, Q => reg_in_47_port);
   reg_in_regx46x : DFFSNQ_X1 port map( D => Plaintext(46), CLK => clk, SN => 
                           n431, Q => reg_in_46_port);
   reg_in_regx45x : DFFSNQ_X1 port map( D => Plaintext(45), CLK => clk, SN => 
                           n430, Q => reg_in_45_port);
   reg_in_regx44x : DFFSNQ_X1 port map( D => Plaintext(44), CLK => clk, SN => 
                           n429, Q => reg_in_44_port);
   reg_in_regx43x : DFFSNQ_X1 port map( D => Plaintext(43), CLK => clk, SN => 
                           n428, Q => reg_in_43_port);
   reg_in_regx42x : DFFSNQ_X1 port map( D => Plaintext(42), CLK => clk, SN => 
                           n427, Q => reg_in_42_port);
   reg_in_regx41x : DFFSNQ_X1 port map( D => Plaintext(41), CLK => clk, SN => 
                           n426, Q => reg_in_41_port);
   reg_in_regx40x : DFFSNQ_X1 port map( D => Plaintext(40), CLK => clk, SN => 
                           n425, Q => reg_in_40_port);
   reg_in_regx39x : DFFSNQ_X1 port map( D => Plaintext(39), CLK => clk, SN => 
                           n424, Q => reg_in_39_port);
   reg_in_regx38x : DFFSNQ_X1 port map( D => Plaintext(38), CLK => clk, SN => 
                           n423, Q => reg_in_38_port);
   reg_in_regx37x : DFFSNQ_X1 port map( D => Plaintext(37), CLK => clk, SN => 
                           n422, Q => reg_in_37_port);
   reg_in_regx36x : DFFSNQ_X1 port map( D => Plaintext(36), CLK => clk, SN => 
                           n421, Q => reg_in_36_port);
   reg_in_regx34x : DFFSNQ_X1 port map( D => Plaintext(34), CLK => clk, SN => 
                           n419, Q => reg_in_34_port);
   reg_in_regx33x : DFFSNQ_X1 port map( D => Plaintext(33), CLK => clk, SN => 
                           n418, Q => reg_in_33_port);
   reg_in_regx32x : DFFSNQ_X1 port map( D => Plaintext(32), CLK => clk, SN => 
                           n417, Q => reg_in_32_port);
   reg_in_regx31x : DFFSNQ_X1 port map( D => Plaintext(31), CLK => clk, SN => 
                           n416, Q => reg_in_31_port);
   reg_in_regx30x : DFFSNQ_X1 port map( D => Plaintext(30), CLK => clk, SN => 
                           n415, Q => reg_in_30_port);
   reg_in_regx28x : DFFSNQ_X1 port map( D => Plaintext(28), CLK => clk, SN => 
                           n413, Q => reg_in_28_port);
   reg_in_regx24x : DFFSNQ_X1 port map( D => Plaintext(24), CLK => clk, SN => 
                           n409, Q => reg_in_24_port);
   reg_in_regx23x : DFFSNQ_X1 port map( D => Plaintext(23), CLK => clk, SN => 
                           n408, Q => reg_in_23_port);
   reg_in_regx22x : DFFSNQ_X1 port map( D => Plaintext(22), CLK => clk, SN => 
                           n407, Q => reg_in_22_port);
   reg_in_regx21x : DFFSNQ_X1 port map( D => Plaintext(21), CLK => clk, SN => 
                           n406, Q => reg_in_21_port);
   reg_in_regx20x : DFFSNQ_X1 port map( D => Plaintext(20), CLK => clk, SN => 
                           n405, Q => reg_in_20_port);
   reg_in_regx19x : DFFSNQ_X1 port map( D => Plaintext(19), CLK => clk, SN => 
                           n404, Q => reg_in_19_port);
   reg_in_regx18x : DFFSNQ_X1 port map( D => Plaintext(18), CLK => clk, SN => 
                           n403, Q => reg_in_18_port);
   reg_in_regx17x : DFFSNQ_X1 port map( D => Plaintext(17), CLK => clk, SN => 
                           n402, Q => reg_in_17_port);
   reg_in_regx16x : DFFSNQ_X1 port map( D => Plaintext(16), CLK => clk, SN => 
                           n401, Q => reg_in_16_port);
   reg_in_regx15x : DFFSNQ_X1 port map( D => Plaintext(15), CLK => clk, SN => 
                           n400, Q => reg_in_15_port);
   reg_in_regx14x : DFFSNQ_X1 port map( D => Plaintext(14), CLK => clk, SN => 
                           n399, Q => reg_in_14_port);
   reg_in_regx13x : DFFSNQ_X1 port map( D => Plaintext(13), CLK => clk, SN => 
                           n398, Q => reg_in_13_port);
   reg_in_regx12x : DFFSNQ_X1 port map( D => Plaintext(12), CLK => clk, SN => 
                           n397, Q => reg_in_12_port);
   reg_in_regx11x : DFFSNQ_X1 port map( D => Plaintext(11), CLK => clk, SN => 
                           n396, Q => reg_in_11_port);
   reg_in_regx10x : DFFSNQ_X1 port map( D => Plaintext(10), CLK => clk, SN => 
                           n395, Q => reg_in_10_port);
   reg_in_regx9x : DFFSNQ_X1 port map( D => Plaintext(9), CLK => clk, SN => 
                           n394, Q => reg_in_9_port);
   reg_in_regx8x : DFFSNQ_X1 port map( D => Plaintext(8), CLK => clk, SN => 
                           n393, Q => reg_in_8_port);
   reg_in_regx7x : DFFSNQ_X1 port map( D => Plaintext(7), CLK => clk, SN => 
                           n392, Q => reg_in_7_port);
   reg_in_regx6x : DFFSNQ_X1 port map( D => Plaintext(6), CLK => clk, SN => 
                           n391, Q => reg_in_6_port);
   reg_in_regx5x : DFFSNQ_X1 port map( D => Plaintext(5), CLK => clk, SN => 
                           n390, Q => reg_in_5_port);
   reg_in_regx4x : DFFSNQ_X1 port map( D => Plaintext(4), CLK => clk, SN => 
                           n389, Q => reg_in_4_port);
   reg_in_regx3x : DFFSNQ_X1 port map( D => Plaintext(3), CLK => clk, SN => 
                           n388, Q => reg_in_3_port);
   reg_in_regx2x : DFFSNQ_X1 port map( D => Plaintext(2), CLK => clk, SN => 
                           n387, Q => reg_in_2_port);
   reg_in_regx1x : DFFSNQ_X1 port map( D => Plaintext(1), CLK => clk, SN => 
                           n386, Q => reg_in_1_port);
   reg_in_regx0x : DFFSNQ_X1 port map( D => Plaintext(0), CLK => clk, SN => 
                           n385, Q => reg_in_0_port);
   reg_key_regx191x : DFFSNQ_X1 port map( D => Key(191), CLK => clk, SN => n384
                           , Q => reg_key_191_port);
   reg_key_regx190x : DFFSNQ_X1 port map( D => Key(190), CLK => clk, SN => n383
                           , Q => reg_key_190_port);
   reg_key_regx189x : DFFSNQ_X1 port map( D => Key(189), CLK => clk, SN => n382
                           , Q => reg_key_189_port);
   reg_key_regx188x : DFFSNQ_X1 port map( D => Key(188), CLK => clk, SN => n381
                           , Q => reg_key_188_port);
   reg_key_regx187x : DFFSNQ_X1 port map( D => Key(187), CLK => clk, SN => n380
                           , Q => reg_key_187_port);
   reg_key_regx186x : DFFSNQ_X1 port map( D => Key(186), CLK => clk, SN => n379
                           , Q => reg_key_186_port);
   reg_key_regx185x : DFFSNQ_X1 port map( D => Key(185), CLK => clk, SN => n378
                           , Q => reg_key_185_port);
   reg_key_regx184x : DFFSNQ_X1 port map( D => Key(184), CLK => clk, SN => n377
                           , Q => reg_key_184_port);
   reg_key_regx183x : DFFSNQ_X1 port map( D => Key(183), CLK => clk, SN => n376
                           , Q => reg_key_183_port);
   reg_key_regx182x : DFFSNQ_X1 port map( D => Key(182), CLK => clk, SN => n375
                           , Q => reg_key_182_port);
   reg_key_regx181x : DFFSNQ_X1 port map( D => Key(181), CLK => clk, SN => n374
                           , Q => reg_key_181_port);
   reg_key_regx180x : DFFSNQ_X1 port map( D => Key(180), CLK => clk, SN => n373
                           , Q => reg_key_180_port);
   reg_key_regx179x : DFFSNQ_X1 port map( D => Key(179), CLK => clk, SN => n372
                           , Q => reg_key_179_port);
   reg_key_regx178x : DFFSNQ_X1 port map( D => Key(178), CLK => clk, SN => n371
                           , Q => reg_key_178_port);
   reg_key_regx177x : DFFSNQ_X1 port map( D => Key(177), CLK => clk, SN => n370
                           , Q => reg_key_177_port);
   reg_key_regx176x : DFFSNQ_X1 port map( D => Key(176), CLK => clk, SN => n369
                           , Q => reg_key_176_port);
   reg_key_regx175x : DFFSNQ_X1 port map( D => Key(175), CLK => clk, SN => n368
                           , Q => reg_key_175_port);
   reg_key_regx174x : DFFSNQ_X1 port map( D => Key(174), CLK => clk, SN => n367
                           , Q => reg_key_174_port);
   reg_key_regx173x : DFFSNQ_X1 port map( D => Key(173), CLK => clk, SN => n366
                           , Q => reg_key_173_port);
   reg_key_regx172x : DFFSNQ_X1 port map( D => Key(172), CLK => clk, SN => n365
                           , Q => reg_key_172_port);
   reg_key_regx171x : DFFSNQ_X1 port map( D => Key(171), CLK => clk, SN => n364
                           , Q => reg_key_171_port);
   reg_key_regx170x : DFFSNQ_X1 port map( D => Key(170), CLK => clk, SN => n363
                           , Q => reg_key_170_port);
   reg_key_regx169x : DFFSNQ_X1 port map( D => Key(169), CLK => clk, SN => n362
                           , Q => reg_key_169_port);
   reg_key_regx168x : DFFSNQ_X1 port map( D => Key(168), CLK => clk, SN => n361
                           , Q => reg_key_168_port);
   reg_key_regx167x : DFFSNQ_X1 port map( D => Key(167), CLK => clk, SN => n360
                           , Q => reg_key_167_port);
   reg_key_regx166x : DFFSNQ_X1 port map( D => Key(166), CLK => clk, SN => n359
                           , Q => reg_key_166_port);
   reg_key_regx165x : DFFSNQ_X1 port map( D => Key(165), CLK => clk, SN => n358
                           , Q => reg_key_165_port);
   reg_key_regx164x : DFFSNQ_X1 port map( D => Key(164), CLK => clk, SN => n357
                           , Q => reg_key_164_port);
   reg_key_regx163x : DFFSNQ_X1 port map( D => Key(163), CLK => clk, SN => n356
                           , Q => reg_key_163_port);
   reg_key_regx162x : DFFSNQ_X1 port map( D => Key(162), CLK => clk, SN => n355
                           , Q => reg_key_162_port);
   reg_key_regx161x : DFFSNQ_X1 port map( D => Key(161), CLK => clk, SN => n354
                           , Q => reg_key_161_port);
   reg_key_regx160x : DFFSNQ_X1 port map( D => Key(160), CLK => clk, SN => n353
                           , Q => reg_key_160_port);
   reg_key_regx159x : DFFSNQ_X1 port map( D => Key(159), CLK => clk, SN => n352
                           , Q => reg_key_159_port);
   reg_key_regx158x : DFFSNQ_X1 port map( D => Key(158), CLK => clk, SN => n351
                           , Q => reg_key_158_port);
   reg_key_regx157x : DFFSNQ_X1 port map( D => Key(157), CLK => clk, SN => n350
                           , Q => reg_key_157_port);
   reg_key_regx156x : DFFSNQ_X1 port map( D => Key(156), CLK => clk, SN => n349
                           , Q => reg_key_156_port);
   reg_key_regx155x : DFFSNQ_X1 port map( D => Key(155), CLK => clk, SN => n348
                           , Q => reg_key_155_port);
   reg_key_regx154x : DFFSNQ_X1 port map( D => Key(154), CLK => clk, SN => n347
                           , Q => reg_key_154_port);
   reg_key_regx153x : DFFSNQ_X1 port map( D => Key(153), CLK => clk, SN => n346
                           , Q => reg_key_153_port);
   reg_key_regx152x : DFFSNQ_X1 port map( D => Key(152), CLK => clk, SN => n345
                           , Q => reg_key_152_port);
   reg_key_regx150x : DFFSNQ_X1 port map( D => Key(150), CLK => clk, SN => n343
                           , Q => reg_key_150_port);
   reg_key_regx149x : DFFSNQ_X1 port map( D => Key(149), CLK => clk, SN => n342
                           , Q => reg_key_149_port);
   reg_key_regx148x : DFFSNQ_X1 port map( D => Key(148), CLK => clk, SN => n341
                           , Q => reg_key_148_port);
   reg_key_regx147x : DFFSNQ_X1 port map( D => Key(147), CLK => clk, SN => n340
                           , Q => reg_key_147_port);
   reg_key_regx146x : DFFSNQ_X1 port map( D => Key(146), CLK => clk, SN => n339
                           , Q => reg_key_146_port);
   reg_key_regx145x : DFFSNQ_X1 port map( D => Key(145), CLK => clk, SN => n338
                           , Q => reg_key_145_port);
   reg_key_regx144x : DFFSNQ_X1 port map( D => Key(144), CLK => clk, SN => n337
                           , Q => reg_key_144_port);
   reg_key_regx143x : DFFSNQ_X1 port map( D => Key(143), CLK => clk, SN => n336
                           , Q => reg_key_143_port);
   reg_key_regx142x : DFFSNQ_X1 port map( D => Key(142), CLK => clk, SN => n335
                           , Q => reg_key_142_port);
   reg_key_regx141x : DFFSNQ_X1 port map( D => Key(141), CLK => clk, SN => n334
                           , Q => reg_key_141_port);
   reg_key_regx140x : DFFSNQ_X1 port map( D => Key(140), CLK => clk, SN => n333
                           , Q => reg_key_140_port);
   reg_key_regx139x : DFFSNQ_X1 port map( D => Key(139), CLK => clk, SN => n332
                           , Q => reg_key_139_port);
   reg_key_regx138x : DFFSNQ_X1 port map( D => Key(138), CLK => clk, SN => n331
                           , Q => reg_key_138_port);
   reg_key_regx137x : DFFSNQ_X1 port map( D => Key(137), CLK => clk, SN => n330
                           , Q => reg_key_137_port);
   reg_key_regx136x : DFFSNQ_X1 port map( D => Key(136), CLK => clk, SN => n329
                           , Q => reg_key_136_port);
   reg_key_regx135x : DFFSNQ_X1 port map( D => Key(135), CLK => clk, SN => n328
                           , Q => reg_key_135_port);
   reg_key_regx134x : DFFSNQ_X1 port map( D => Key(134), CLK => clk, SN => n327
                           , Q => reg_key_134_port);
   reg_key_regx133x : DFFSNQ_X1 port map( D => Key(133), CLK => clk, SN => n326
                           , Q => reg_key_133_port);
   reg_key_regx132x : DFFSNQ_X1 port map( D => Key(132), CLK => clk, SN => n325
                           , Q => reg_key_132_port);
   reg_key_regx131x : DFFSNQ_X1 port map( D => Key(131), CLK => clk, SN => n324
                           , Q => reg_key_131_port);
   reg_key_regx130x : DFFSNQ_X1 port map( D => Key(130), CLK => clk, SN => n323
                           , Q => reg_key_130_port);
   reg_key_regx129x : DFFSNQ_X1 port map( D => Key(129), CLK => clk, SN => n322
                           , Q => reg_key_129_port);
   reg_key_regx128x : DFFSNQ_X1 port map( D => Key(128), CLK => clk, SN => n321
                           , Q => reg_key_128_port);
   reg_key_regx127x : DFFSNQ_X1 port map( D => Key(127), CLK => clk, SN => n320
                           , Q => reg_key_127_port);
   reg_key_regx126x : DFFSNQ_X1 port map( D => Key(126), CLK => clk, SN => n319
                           , Q => reg_key_126_port);
   reg_key_regx125x : DFFSNQ_X1 port map( D => Key(125), CLK => clk, SN => n318
                           , Q => reg_key_125_port);
   reg_key_regx124x : DFFSNQ_X1 port map( D => Key(124), CLK => clk, SN => n317
                           , Q => reg_key_124_port);
   reg_key_regx123x : DFFSNQ_X1 port map( D => Key(123), CLK => clk, SN => n316
                           , Q => reg_key_123_port);
   reg_key_regx122x : DFFSNQ_X1 port map( D => Key(122), CLK => clk, SN => n315
                           , Q => reg_key_122_port);
   reg_key_regx121x : DFFSNQ_X1 port map( D => Key(121), CLK => clk, SN => n314
                           , Q => reg_key_121_port);
   reg_key_regx120x : DFFSNQ_X1 port map( D => Key(120), CLK => clk, SN => n313
                           , Q => reg_key_120_port);
   reg_key_regx119x : DFFSNQ_X1 port map( D => Key(119), CLK => clk, SN => n312
                           , Q => reg_key_119_port);
   reg_key_regx118x : DFFSNQ_X1 port map( D => Key(118), CLK => clk, SN => n311
                           , Q => reg_key_118_port);
   reg_key_regx117x : DFFSNQ_X1 port map( D => Key(117), CLK => clk, SN => n310
                           , Q => reg_key_117_port);
   reg_key_regx116x : DFFSNQ_X1 port map( D => Key(116), CLK => clk, SN => n309
                           , Q => reg_key_116_port);
   reg_key_regx115x : DFFSNQ_X1 port map( D => Key(115), CLK => clk, SN => n308
                           , Q => reg_key_115_port);
   reg_key_regx114x : DFFSNQ_X1 port map( D => Key(114), CLK => clk, SN => n307
                           , Q => reg_key_114_port);
   reg_key_regx113x : DFFSNQ_X1 port map( D => Key(113), CLK => clk, SN => n306
                           , Q => reg_key_113_port);
   reg_key_regx112x : DFFSNQ_X1 port map( D => Key(112), CLK => clk, SN => n305
                           , Q => reg_key_112_port);
   reg_key_regx111x : DFFSNQ_X1 port map( D => Key(111), CLK => clk, SN => n304
                           , Q => reg_key_111_port);
   reg_key_regx110x : DFFSNQ_X1 port map( D => Key(110), CLK => clk, SN => n303
                           , Q => reg_key_110_port);
   reg_key_regx109x : DFFSNQ_X1 port map( D => Key(109), CLK => clk, SN => n302
                           , Q => reg_key_109_port);
   reg_key_regx108x : DFFSNQ_X1 port map( D => Key(108), CLK => clk, SN => n301
                           , Q => reg_key_108_port);
   reg_key_regx107x : DFFSNQ_X1 port map( D => Key(107), CLK => clk, SN => n300
                           , Q => reg_key_107_port);
   reg_key_regx106x : DFFSNQ_X1 port map( D => Key(106), CLK => clk, SN => n299
                           , Q => reg_key_106_port);
   reg_key_regx105x : DFFSNQ_X1 port map( D => Key(105), CLK => clk, SN => n298
                           , Q => reg_key_105_port);
   reg_key_regx104x : DFFSNQ_X1 port map( D => Key(104), CLK => clk, SN => n297
                           , Q => reg_key_104_port);
   reg_key_regx103x : DFFSNQ_X1 port map( D => Key(103), CLK => clk, SN => n296
                           , Q => reg_key_103_port);
   reg_key_regx102x : DFFSNQ_X1 port map( D => Key(102), CLK => clk, SN => n295
                           , Q => reg_key_102_port);
   reg_key_regx101x : DFFSNQ_X1 port map( D => Key(101), CLK => clk, SN => n294
                           , Q => reg_key_101_port);
   reg_key_regx100x : DFFSNQ_X1 port map( D => Key(100), CLK => clk, SN => n293
                           , Q => reg_key_100_port);
   reg_key_regx99x : DFFSNQ_X1 port map( D => Key(99), CLK => clk, SN => n292, 
                           Q => reg_key_99_port);
   reg_key_regx98x : DFFSNQ_X1 port map( D => Key(98), CLK => clk, SN => n291, 
                           Q => reg_key_98_port);
   reg_key_regx97x : DFFSNQ_X1 port map( D => Key(97), CLK => clk, SN => n290, 
                           Q => reg_key_97_port);
   reg_key_regx96x : DFFSNQ_X1 port map( D => Key(96), CLK => clk, SN => n289, 
                           Q => reg_key_96_port);
   reg_key_regx95x : DFFSNQ_X1 port map( D => Key(95), CLK => clk, SN => n288, 
                           Q => reg_key_95_port);
   reg_key_regx94x : DFFSNQ_X1 port map( D => Key(94), CLK => clk, SN => n287, 
                           Q => reg_key_94_port);
   reg_key_regx93x : DFFSNQ_X1 port map( D => Key(93), CLK => clk, SN => n286, 
                           Q => reg_key_93_port);
   reg_key_regx92x : DFFSNQ_X1 port map( D => Key(92), CLK => clk, SN => n285, 
                           Q => reg_key_92_port);
   reg_key_regx91x : DFFSNQ_X1 port map( D => Key(91), CLK => clk, SN => n284, 
                           Q => reg_key_91_port);
   reg_key_regx90x : DFFSNQ_X1 port map( D => Key(90), CLK => clk, SN => n283, 
                           Q => reg_key_90_port);
   reg_key_regx89x : DFFSNQ_X1 port map( D => Key(89), CLK => clk, SN => n282, 
                           Q => reg_key_89_port);
   reg_key_regx88x : DFFSNQ_X1 port map( D => Key(88), CLK => clk, SN => n281, 
                           Q => reg_key_88_port);
   reg_key_regx87x : DFFSNQ_X1 port map( D => Key(87), CLK => clk, SN => n280, 
                           Q => reg_key_87_port);
   reg_key_regx86x : DFFSNQ_X1 port map( D => Key(86), CLK => clk, SN => n279, 
                           Q => reg_key_86_port);
   reg_key_regx85x : DFFSNQ_X1 port map( D => Key(85), CLK => clk, SN => n278, 
                           Q => reg_key_85_port);
   reg_key_regx84x : DFFSNQ_X1 port map( D => Key(84), CLK => clk, SN => n277, 
                           Q => reg_key_84_port);
   reg_key_regx83x : DFFSNQ_X1 port map( D => Key(83), CLK => clk, SN => n276, 
                           Q => reg_key_83_port);
   reg_key_regx82x : DFFSNQ_X1 port map( D => Key(82), CLK => clk, SN => n275, 
                           Q => reg_key_82_port);
   reg_key_regx81x : DFFSNQ_X1 port map( D => Key(81), CLK => clk, SN => n274, 
                           Q => reg_key_81_port);
   reg_key_regx80x : DFFSNQ_X1 port map( D => Key(80), CLK => clk, SN => n273, 
                           Q => reg_key_80_port);
   reg_key_regx79x : DFFSNQ_X1 port map( D => Key(79), CLK => clk, SN => n272, 
                           Q => reg_key_79_port);
   reg_key_regx78x : DFFSNQ_X1 port map( D => Key(78), CLK => clk, SN => n271, 
                           Q => reg_key_78_port);
   reg_key_regx77x : DFFSNQ_X1 port map( D => Key(77), CLK => clk, SN => n270, 
                           Q => reg_key_77_port);
   reg_key_regx76x : DFFSNQ_X1 port map( D => Key(76), CLK => clk, SN => n269, 
                           Q => reg_key_76_port);
   reg_key_regx75x : DFFSNQ_X1 port map( D => Key(75), CLK => clk, SN => n268, 
                           Q => reg_key_75_port);
   reg_key_regx74x : DFFSNQ_X1 port map( D => Key(74), CLK => clk, SN => n267, 
                           Q => reg_key_74_port);
   reg_key_regx73x : DFFSNQ_X1 port map( D => Key(73), CLK => clk, SN => n266, 
                           Q => reg_key_73_port);
   reg_key_regx72x : DFFSNQ_X1 port map( D => Key(72), CLK => clk, SN => n265, 
                           Q => reg_key_72_port);
   reg_key_regx71x : DFFSNQ_X1 port map( D => Key(71), CLK => clk, SN => n264, 
                           Q => reg_key_71_port);
   reg_key_regx70x : DFFSNQ_X1 port map( D => Key(70), CLK => clk, SN => n263, 
                           Q => reg_key_70_port);
   reg_key_regx69x : DFFSNQ_X1 port map( D => Key(69), CLK => clk, SN => n262, 
                           Q => reg_key_69_port);
   reg_key_regx68x : DFFSNQ_X1 port map( D => Key(68), CLK => clk, SN => n261, 
                           Q => reg_key_68_port);
   reg_key_regx67x : DFFSNQ_X1 port map( D => Key(67), CLK => clk, SN => n260, 
                           Q => reg_key_67_port);
   reg_key_regx66x : DFFSNQ_X1 port map( D => Key(66), CLK => clk, SN => n259, 
                           Q => reg_key_66_port);
   reg_key_regx65x : DFFSNQ_X1 port map( D => Key(65), CLK => clk, SN => n258, 
                           Q => reg_key_65_port);
   reg_key_regx64x : DFFSNQ_X1 port map( D => Key(64), CLK => clk, SN => n257, 
                           Q => reg_key_64_port);
   reg_key_regx63x : DFFSNQ_X1 port map( D => Key(63), CLK => clk, SN => n256, 
                           Q => reg_key_63_port);
   reg_key_regx62x : DFFSNQ_X1 port map( D => Key(62), CLK => clk, SN => n255, 
                           Q => reg_key_62_port);
   reg_key_regx61x : DFFSNQ_X1 port map( D => Key(61), CLK => clk, SN => n254, 
                           Q => reg_key_61_port);
   reg_key_regx60x : DFFSNQ_X1 port map( D => Key(60), CLK => clk, SN => n253, 
                           Q => reg_key_60_port);
   reg_key_regx59x : DFFSNQ_X1 port map( D => Key(59), CLK => clk, SN => n252, 
                           Q => reg_key_59_port);
   reg_key_regx58x : DFFSNQ_X1 port map( D => Key(58), CLK => clk, SN => n251, 
                           Q => reg_key_58_port);
   reg_key_regx57x : DFFSNQ_X1 port map( D => Key(57), CLK => clk, SN => n250, 
                           Q => reg_key_57_port);
   reg_key_regx56x : DFFSNQ_X1 port map( D => Key(56), CLK => clk, SN => n249, 
                           Q => reg_key_56_port);
   reg_key_regx55x : DFFSNQ_X1 port map( D => Key(55), CLK => clk, SN => n248, 
                           Q => reg_key_55_port);
   reg_key_regx54x : DFFSNQ_X1 port map( D => Key(54), CLK => clk, SN => n247, 
                           Q => reg_key_54_port);
   reg_key_regx53x : DFFSNQ_X1 port map( D => Key(53), CLK => clk, SN => n246, 
                           Q => reg_key_53_port);
   reg_key_regx52x : DFFSNQ_X1 port map( D => Key(52), CLK => clk, SN => n245, 
                           Q => reg_key_52_port);
   reg_key_regx51x : DFFSNQ_X1 port map( D => Key(51), CLK => clk, SN => n244, 
                           Q => reg_key_51_port);
   reg_key_regx50x : DFFSNQ_X1 port map( D => Key(50), CLK => clk, SN => n243, 
                           Q => reg_key_50_port);
   reg_key_regx49x : DFFSNQ_X1 port map( D => Key(49), CLK => clk, SN => n242, 
                           Q => reg_key_49_port);
   reg_key_regx48x : DFFSNQ_X1 port map( D => Key(48), CLK => clk, SN => n241, 
                           Q => reg_key_48_port);
   reg_key_regx47x : DFFSNQ_X1 port map( D => Key(47), CLK => clk, SN => n240, 
                           Q => reg_key_47_port);
   reg_key_regx46x : DFFSNQ_X1 port map( D => Key(46), CLK => clk, SN => n239, 
                           Q => reg_key_46_port);
   reg_key_regx45x : DFFSNQ_X1 port map( D => Key(45), CLK => clk, SN => n238, 
                           Q => reg_key_45_port);
   reg_key_regx44x : DFFSNQ_X1 port map( D => Key(44), CLK => clk, SN => n237, 
                           Q => reg_key_44_port);
   reg_key_regx43x : DFFSNQ_X1 port map( D => Key(43), CLK => clk, SN => n236, 
                           Q => reg_key_43_port);
   reg_key_regx42x : DFFSNQ_X1 port map( D => Key(42), CLK => clk, SN => n235, 
                           Q => reg_key_42_port);
   reg_key_regx41x : DFFSNQ_X1 port map( D => Key(41), CLK => clk, SN => n234, 
                           Q => reg_key_41_port);
   reg_key_regx40x : DFFSNQ_X1 port map( D => Key(40), CLK => clk, SN => n233, 
                           Q => reg_key_40_port);
   reg_key_regx39x : DFFSNQ_X1 port map( D => Key(39), CLK => clk, SN => n232, 
                           Q => reg_key_39_port);
   reg_key_regx38x : DFFSNQ_X1 port map( D => Key(38), CLK => clk, SN => n231, 
                           Q => reg_key_38_port);
   reg_key_regx36x : DFFSNQ_X1 port map( D => Key(36), CLK => clk, SN => n229, 
                           Q => reg_key_36_port);
   reg_key_regx35x : DFFSNQ_X1 port map( D => Key(35), CLK => clk, SN => n228, 
                           Q => reg_key_35_port);
   reg_key_regx34x : DFFSNQ_X1 port map( D => Key(34), CLK => clk, SN => n227, 
                           Q => reg_key_34_port);
   reg_key_regx33x : DFFSNQ_X1 port map( D => Key(33), CLK => clk, SN => n226, 
                           Q => reg_key_33_port);
   reg_key_regx32x : DFFSNQ_X1 port map( D => Key(32), CLK => clk, SN => n225, 
                           Q => reg_key_32_port);
   reg_key_regx31x : DFFSNQ_X1 port map( D => Key(31), CLK => clk, SN => n224, 
                           Q => reg_key_31_port);
   reg_key_regx30x : DFFSNQ_X1 port map( D => Key(30), CLK => clk, SN => n223, 
                           Q => reg_key_30_port);
   reg_key_regx29x : DFFSNQ_X1 port map( D => Key(29), CLK => clk, SN => n222, 
                           Q => reg_key_29_port);
   reg_key_regx28x : DFFSNQ_X1 port map( D => Key(28), CLK => clk, SN => n221, 
                           Q => reg_key_28_port);
   reg_key_regx27x : DFFSNQ_X1 port map( D => Key(27), CLK => clk, SN => n220, 
                           Q => reg_key_27_port);
   reg_key_regx26x : DFFSNQ_X1 port map( D => Key(26), CLK => clk, SN => n219, 
                           Q => reg_key_26_port);
   reg_key_regx25x : DFFSNQ_X1 port map( D => Key(25), CLK => clk, SN => n218, 
                           Q => reg_key_25_port);
   reg_key_regx24x : DFFSNQ_X1 port map( D => Key(24), CLK => clk, SN => n217, 
                           Q => reg_key_24_port);
   reg_key_regx23x : DFFSNQ_X1 port map( D => Key(23), CLK => clk, SN => n216, 
                           Q => reg_key_23_port);
   reg_key_regx22x : DFFSNQ_X1 port map( D => Key(22), CLK => clk, SN => n215, 
                           Q => reg_key_22_port);
   reg_key_regx21x : DFFSNQ_X1 port map( D => Key(21), CLK => clk, SN => n214, 
                           Q => reg_key_21_port);
   reg_key_regx20x : DFFSNQ_X1 port map( D => Key(20), CLK => clk, SN => n213, 
                           Q => reg_key_20_port);
   reg_key_regx19x : DFFSNQ_X1 port map( D => Key(19), CLK => clk, SN => n212, 
                           Q => reg_key_19_port);
   reg_key_regx18x : DFFSNQ_X1 port map( D => Key(18), CLK => clk, SN => n211, 
                           Q => reg_key_18_port);
   reg_key_regx17x : DFFSNQ_X1 port map( D => Key(17), CLK => clk, SN => n210, 
                           Q => reg_key_17_port);
   reg_key_regx16x : DFFSNQ_X1 port map( D => Key(16), CLK => clk, SN => n209, 
                           Q => reg_key_16_port);
   reg_key_regx15x : DFFSNQ_X1 port map( D => Key(15), CLK => clk, SN => n208, 
                           Q => reg_key_15_port);
   reg_key_regx14x : DFFSNQ_X1 port map( D => Key(14), CLK => clk, SN => n207, 
                           Q => reg_key_14_port);
   reg_key_regx13x : DFFSNQ_X1 port map( D => Key(13), CLK => clk, SN => n206, 
                           Q => reg_key_13_port);
   reg_key_regx12x : DFFSNQ_X1 port map( D => Key(12), CLK => clk, SN => n205, 
                           Q => reg_key_12_port);
   reg_key_regx11x : DFFSNQ_X1 port map( D => Key(11), CLK => clk, SN => n204, 
                           Q => reg_key_11_port);
   reg_key_regx10x : DFFSNQ_X1 port map( D => Key(10), CLK => clk, SN => n203, 
                           Q => reg_key_10_port);
   reg_key_regx9x : DFFSNQ_X1 port map( D => Key(9), CLK => clk, SN => n202, Q 
                           => reg_key_9_port);
   reg_key_regx8x : DFFSNQ_X1 port map( D => Key(8), CLK => clk, SN => n201, Q 
                           => reg_key_8_port);
   reg_key_regx7x : DFFSNQ_X1 port map( D => Key(7), CLK => clk, SN => n200, Q 
                           => reg_key_7_port);
   reg_key_regx6x : DFFSNQ_X1 port map( D => Key(6), CLK => clk, SN => n199, Q 
                           => reg_key_6_port);
   reg_key_regx5x : DFFSNQ_X1 port map( D => Key(5), CLK => clk, SN => n198, Q 
                           => reg_key_5_port);
   reg_key_regx4x : DFFSNQ_X1 port map( D => Key(4), CLK => clk, SN => n197, Q 
                           => reg_key_4_port);
   reg_key_regx3x : DFFSNQ_X1 port map( D => Key(3), CLK => clk, SN => n196, Q 
                           => reg_key_3_port);
   reg_key_regx2x : DFFSNQ_X1 port map( D => Key(2), CLK => clk, SN => n195, Q 
                           => reg_key_2_port);
   reg_key_regx1x : DFFSNQ_X1 port map( D => Key(1), CLK => clk, SN => n194, Q 
                           => reg_key_1_port);
   reg_key_regx0x : DFFSNQ_X1 port map( D => Key(0), CLK => clk, SN => n193, Q 
                           => reg_key_0_port);
   Ciphertext_regx191x : DFFSNQ_X1 port map( D => reg_out_191_port, CLK => clk,
                           SN => n192, Q => Ciphertext(191));
   Ciphertext_regx188x : DFFSNQ_X1 port map( D => reg_out_188_port, CLK => clk,
                           SN => n189, Q => Ciphertext(188));
   Ciphertext_regx187x : DFFSNQ_X1 port map( D => reg_out_187_port, CLK => clk,
                           SN => n188, Q => Ciphertext(187));
   Ciphertext_regx184x : DFFSNQ_X1 port map( D => reg_out_184_port, CLK => clk,
                           SN => n185, Q => Ciphertext(184));
   Ciphertext_regx183x : DFFSNQ_X1 port map( D => reg_out_183_port, CLK => clk,
                           SN => n184, Q => Ciphertext(183));
   Ciphertext_regx181x : DFFSNQ_X1 port map( D => reg_out_181_port, CLK => clk,
                           SN => n182, Q => Ciphertext(181));
   Ciphertext_regx179x : DFFSNQ_X1 port map( D => reg_out_179_port, CLK => clk,
                           SN => n180, Q => Ciphertext(179));
   Ciphertext_regx178x : DFFSNQ_X1 port map( D => reg_out_178_port, CLK => clk,
                           SN => n179, Q => Ciphertext(178));
   Ciphertext_regx177x : DFFSNQ_X1 port map( D => reg_out_177_port, CLK => clk,
                           SN => n178, Q => Ciphertext(177));
   Ciphertext_regx176x : DFFSNQ_X1 port map( D => reg_out_176_port, CLK => clk,
                           SN => n177, Q => Ciphertext(176));
   Ciphertext_regx175x : DFFSNQ_X1 port map( D => reg_out_175_port, CLK => clk,
                           SN => n176, Q => Ciphertext(175));
   Ciphertext_regx173x : DFFSNQ_X1 port map( D => reg_out_173_port, CLK => clk,
                           SN => n174, Q => Ciphertext(173));
   Ciphertext_regx172x : DFFSNQ_X1 port map( D => reg_out_172_port, CLK => clk,
                           SN => n173, Q => Ciphertext(172));
   Ciphertext_regx170x : DFFSNQ_X1 port map( D => reg_out_170_port, CLK => clk,
                           SN => n171, Q => Ciphertext(170));
   Ciphertext_regx168x : DFFSNQ_X1 port map( D => reg_out_168_port, CLK => clk,
                           SN => n169, Q => Ciphertext(168));
   Ciphertext_regx167x : DFFSNQ_X1 port map( D => reg_out_167_port, CLK => clk,
                           SN => n168, Q => Ciphertext(167));
   Ciphertext_regx166x : DFFSNQ_X1 port map( D => reg_out_166_port, CLK => clk,
                           SN => n167, Q => Ciphertext(166));
   Ciphertext_regx163x : DFFSNQ_X1 port map( D => reg_out_163_port, CLK => clk,
                           SN => n164, Q => Ciphertext(163));
   Ciphertext_regx161x : DFFSNQ_X1 port map( D => reg_out_161_port, CLK => clk,
                           SN => n162, Q => Ciphertext(161));
   Ciphertext_regx158x : DFFSNQ_X1 port map( D => reg_out_158_port, CLK => clk,
                           SN => n159, Q => Ciphertext(158));
   Ciphertext_regx157x : DFFSNQ_X1 port map( D => reg_out_157_port, CLK => clk,
                           SN => n158, Q => Ciphertext(157));
   Ciphertext_regx156x : DFFSNQ_X1 port map( D => reg_out_156_port, CLK => clk,
                           SN => n157, Q => Ciphertext(156));
   Ciphertext_regx155x : DFFSNQ_X1 port map( D => reg_out_155_port, CLK => clk,
                           SN => n156, Q => Ciphertext(155));
   Ciphertext_regx151x : DFFSNQ_X1 port map( D => reg_out_151_port, CLK => clk,
                           SN => n152, Q => Ciphertext(151));
   Ciphertext_regx150x : DFFSNQ_X1 port map( D => reg_out_150_port, CLK => clk,
                           SN => n151, Q => Ciphertext(150));
   Ciphertext_regx149x : DFFSNQ_X1 port map( D => reg_out_149_port, CLK => clk,
                           SN => n150, Q => Ciphertext(149));
   Ciphertext_regx148x : DFFSNQ_X1 port map( D => reg_out_148_port, CLK => clk,
                           SN => n149, Q => Ciphertext(148));
   Ciphertext_regx147x : DFFSNQ_X1 port map( D => reg_out_147_port, CLK => clk,
                           SN => n148, Q => Ciphertext(147));
   Ciphertext_regx145x : DFFSNQ_X1 port map( D => reg_out_145_port, CLK => clk,
                           SN => n146, Q => Ciphertext(145));
   Ciphertext_regx144x : DFFSNQ_X1 port map( D => reg_out_144_port, CLK => clk,
                           SN => n145, Q => Ciphertext(144));
   Ciphertext_regx142x : DFFSNQ_X1 port map( D => reg_out_142_port, CLK => clk,
                           SN => n143, Q => Ciphertext(142));
   Ciphertext_regx141x : DFFSNQ_X1 port map( D => reg_out_141_port, CLK => clk,
                           SN => n142, Q => Ciphertext(141));
   Ciphertext_regx140x : DFFSNQ_X1 port map( D => reg_out_140_port, CLK => clk,
                           SN => n141, Q => Ciphertext(140));
   Ciphertext_regx139x : DFFSNQ_X1 port map( D => reg_out_139_port, CLK => clk,
                           SN => n140, Q => Ciphertext(139));
   Ciphertext_regx138x : DFFSNQ_X1 port map( D => reg_out_138_port, CLK => clk,
                           SN => n139, Q => Ciphertext(138));
   Ciphertext_regx135x : DFFSNQ_X1 port map( D => reg_out_135_port, CLK => clk,
                           SN => n136, Q => Ciphertext(135));
   Ciphertext_regx134x : DFFSNQ_X1 port map( D => reg_out_134_port, CLK => clk,
                           SN => n135, Q => Ciphertext(134));
   Ciphertext_regx129x : DFFSNQ_X1 port map( D => reg_out_129_port, CLK => clk,
                           SN => n130, Q => Ciphertext(129));
   Ciphertext_regx128x : DFFSNQ_X1 port map( D => reg_out_128_port, CLK => clk,
                           SN => n129, Q => Ciphertext(128));
   Ciphertext_regx127x : DFFSNQ_X1 port map( D => reg_out_127_port, CLK => clk,
                           SN => n128, Q => Ciphertext(127));
   Ciphertext_regx126x : DFFSNQ_X1 port map( D => reg_out_126_port, CLK => clk,
                           SN => n127, Q => Ciphertext(126));
   Ciphertext_regx123x : DFFSNQ_X1 port map( D => reg_out_123_port, CLK => clk,
                           SN => n124, Q => Ciphertext(123));
   Ciphertext_regx122x : DFFSNQ_X1 port map( D => reg_out_122_port, CLK => clk,
                           SN => n123, Q => Ciphertext(122));
   Ciphertext_regx121x : DFFSNQ_X1 port map( D => reg_out_121_port, CLK => clk,
                           SN => n122, Q => Ciphertext(121));
   Ciphertext_regx119x : DFFSNQ_X1 port map( D => reg_out_119_port, CLK => clk,
                           SN => n120, Q => Ciphertext(119));
   Ciphertext_regx118x : DFFSNQ_X1 port map( D => reg_out_118_port, CLK => clk,
                           SN => n119, Q => Ciphertext(118));
   Ciphertext_regx115x : DFFSNQ_X1 port map( D => reg_out_115_port, CLK => clk,
                           SN => n116, Q => Ciphertext(115));
   Ciphertext_regx113x : DFFSNQ_X1 port map( D => reg_out_113_port, CLK => clk,
                           SN => n114, Q => Ciphertext(113));
   Ciphertext_regx112x : DFFSNQ_X1 port map( D => reg_out_112_port, CLK => clk,
                           SN => n113, Q => Ciphertext(112));
   Ciphertext_regx110x : DFFSNQ_X1 port map( D => reg_out_110_port, CLK => clk,
                           SN => n111, Q => Ciphertext(110));
   Ciphertext_regx109x : DFFSNQ_X1 port map( D => reg_out_109_port, CLK => clk,
                           SN => n110, Q => Ciphertext(109));
   Ciphertext_regx108x : DFFSNQ_X1 port map( D => reg_out_108_port, CLK => clk,
                           SN => n109, Q => Ciphertext(108));
   Ciphertext_regx107x : DFFSNQ_X1 port map( D => reg_out_107_port, CLK => clk,
                           SN => n108, Q => Ciphertext(107));
   Ciphertext_regx106x : DFFSNQ_X1 port map( D => reg_out_106_port, CLK => clk,
                           SN => n107, Q => Ciphertext(106));
   Ciphertext_regx105x : DFFSNQ_X1 port map( D => reg_out_105_port, CLK => clk,
                           SN => n106, Q => Ciphertext(105));
   Ciphertext_regx104x : DFFSNQ_X1 port map( D => reg_out_104_port, CLK => clk,
                           SN => n105, Q => Ciphertext(104));
   Ciphertext_regx103x : DFFSNQ_X1 port map( D => reg_out_103_port, CLK => clk,
                           SN => n104, Q => Ciphertext(103));
   Ciphertext_regx102x : DFFSNQ_X1 port map( D => reg_out_102_port, CLK => clk,
                           SN => n103, Q => Ciphertext(102));
   Ciphertext_regx98x : DFFSNQ_X1 port map( D => reg_out_98_port, CLK => clk, 
                           SN => n99, Q => Ciphertext(98));
   Ciphertext_regx96x : DFFSNQ_X1 port map( D => reg_out_96_port, CLK => clk, 
                           SN => n97, Q => Ciphertext(96));
   Ciphertext_regx93x : DFFSNQ_X1 port map( D => reg_out_93_port, CLK => clk, 
                           SN => n94, Q => Ciphertext(93));
   Ciphertext_regx92x : DFFSNQ_X1 port map( D => reg_out_92_port, CLK => clk, 
                           SN => n93, Q => Ciphertext(92));
   Ciphertext_regx91x : DFFSNQ_X1 port map( D => reg_out_91_port, CLK => clk, 
                           SN => n92, Q => Ciphertext(91));
   Ciphertext_regx90x : DFFSNQ_X1 port map( D => reg_out_90_port, CLK => clk, 
                           SN => n91, Q => Ciphertext(90));
   Ciphertext_regx89x : DFFSNQ_X1 port map( D => reg_out_89_port, CLK => clk, 
                           SN => n90, Q => Ciphertext(89));
   Ciphertext_regx86x : DFFSNQ_X1 port map( D => reg_out_86_port, CLK => clk, 
                           SN => n87, Q => Ciphertext(86));
   Ciphertext_regx85x : DFFSNQ_X1 port map( D => reg_out_85_port, CLK => clk, 
                           SN => n86, Q => Ciphertext(85));
   Ciphertext_regx84x : DFFSNQ_X1 port map( D => reg_out_84_port, CLK => clk, 
                           SN => n85, Q => Ciphertext(84));
   Ciphertext_regx83x : DFFSNQ_X1 port map( D => reg_out_83_port, CLK => clk, 
                           SN => n84, Q => Ciphertext(83));
   Ciphertext_regx82x : DFFSNQ_X1 port map( D => reg_out_82_port, CLK => clk, 
                           SN => n83, Q => Ciphertext(82));
   Ciphertext_regx81x : DFFSNQ_X1 port map( D => reg_out_81_port, CLK => clk, 
                           SN => n82, Q => Ciphertext(81));
   Ciphertext_regx80x : DFFSNQ_X1 port map( D => reg_out_80_port, CLK => clk, 
                           SN => n81, Q => Ciphertext(80));
   Ciphertext_regx79x : DFFSNQ_X1 port map( D => reg_out_79_port, CLK => clk, 
                           SN => n80, Q => Ciphertext(79));
   Ciphertext_regx78x : DFFSNQ_X1 port map( D => reg_out_78_port, CLK => clk, 
                           SN => n79, Q => Ciphertext(78));
   Ciphertext_regx77x : DFFSNQ_X1 port map( D => reg_out_77_port, CLK => clk, 
                           SN => n78, Q => Ciphertext(77));
   Ciphertext_regx76x : DFFSNQ_X1 port map( D => reg_out_76_port, CLK => clk, 
                           SN => n77, Q => Ciphertext(76));
   Ciphertext_regx74x : DFFSNQ_X1 port map( D => reg_out_74_port, CLK => clk, 
                           SN => n75, Q => Ciphertext(74));
   Ciphertext_regx73x : DFFSNQ_X1 port map( D => reg_out_73_port, CLK => clk, 
                           SN => n74, Q => Ciphertext(73));
   Ciphertext_regx71x : DFFSNQ_X1 port map( D => reg_out_71_port, CLK => clk, 
                           SN => n72, Q => Ciphertext(71));
   Ciphertext_regx70x : DFFSNQ_X1 port map( D => reg_out_70_port, CLK => clk, 
                           SN => n71, Q => Ciphertext(70));
   Ciphertext_regx69x : DFFSNQ_X1 port map( D => reg_out_69_port, CLK => clk, 
                           SN => n70, Q => Ciphertext(69));
   Ciphertext_regx68x : DFFSNQ_X1 port map( D => reg_out_68_port, CLK => clk, 
                           SN => n69, Q => Ciphertext(68));
   Ciphertext_regx67x : DFFSNQ_X1 port map( D => reg_out_67_port, CLK => clk, 
                           SN => n68, Q => Ciphertext(67));
   Ciphertext_regx66x : DFFSNQ_X1 port map( D => reg_out_66_port, CLK => clk, 
                           SN => n67, Q => Ciphertext(66));
   Ciphertext_regx65x : DFFSNQ_X1 port map( D => reg_out_65_port, CLK => clk, 
                           SN => n66, Q => Ciphertext(65));
   Ciphertext_regx64x : DFFSNQ_X1 port map( D => reg_out_64_port, CLK => clk, 
                           SN => n65, Q => Ciphertext(64));
   Ciphertext_regx63x : DFFSNQ_X1 port map( D => reg_out_63_port, CLK => clk, 
                           SN => n64, Q => Ciphertext(63));
   Ciphertext_regx62x : DFFSNQ_X1 port map( D => reg_out_62_port, CLK => clk, 
                           SN => n63, Q => Ciphertext(62));
   Ciphertext_regx61x : DFFSNQ_X1 port map( D => reg_out_61_port, CLK => clk, 
                           SN => n62, Q => Ciphertext(61));
   Ciphertext_regx60x : DFFSNQ_X1 port map( D => reg_out_60_port, CLK => clk, 
                           SN => n61, Q => Ciphertext(60));
   Ciphertext_regx55x : DFFSNQ_X1 port map( D => reg_out_55_port, CLK => clk, 
                           SN => n56, Q => Ciphertext(55));
   Ciphertext_regx53x : DFFSNQ_X1 port map( D => reg_out_53_port, CLK => clk, 
                           SN => n54, Q => Ciphertext(53));
   Ciphertext_regx52x : DFFSNQ_X1 port map( D => reg_out_52_port, CLK => clk, 
                           SN => n53, Q => Ciphertext(52));
   Ciphertext_regx51x : DFFSNQ_X1 port map( D => reg_out_51_port, CLK => clk, 
                           SN => n52, Q => Ciphertext(51));
   Ciphertext_regx50x : DFFSNQ_X1 port map( D => reg_out_50_port, CLK => clk, 
                           SN => n51, Q => Ciphertext(50));
   Ciphertext_regx48x : DFFSNQ_X1 port map( D => reg_out_48_port, CLK => clk, 
                           SN => n49, Q => Ciphertext(48));
   Ciphertext_regx47x : DFFSNQ_X1 port map( D => reg_out_47_port, CLK => clk, 
                           SN => n48, Q => Ciphertext(47));
   Ciphertext_regx46x : DFFSNQ_X1 port map( D => reg_out_46_port, CLK => clk, 
                           SN => n47, Q => Ciphertext(46));
   Ciphertext_regx45x : DFFSNQ_X1 port map( D => reg_out_45_port, CLK => clk, 
                           SN => n46, Q => Ciphertext(45));
   Ciphertext_regx44x : DFFSNQ_X1 port map( D => reg_out_44_port, CLK => clk, 
                           SN => n45, Q => Ciphertext(44));
   Ciphertext_regx43x : DFFSNQ_X1 port map( D => reg_out_43_port, CLK => clk, 
                           SN => n44, Q => Ciphertext(43));
   Ciphertext_regx42x : DFFSNQ_X1 port map( D => reg_out_42_port, CLK => clk, 
                           SN => n43, Q => Ciphertext(42));
   Ciphertext_regx41x : DFFSNQ_X1 port map( D => reg_out_41_port, CLK => clk, 
                           SN => n42, Q => Ciphertext(41));
   Ciphertext_regx40x : DFFSNQ_X1 port map( D => reg_out_40_port, CLK => clk, 
                           SN => n41, Q => Ciphertext(40));
   Ciphertext_regx38x : DFFSNQ_X1 port map( D => reg_out_38_port, CLK => clk, 
                           SN => n39, Q => Ciphertext(38));
   Ciphertext_regx37x : DFFSNQ_X1 port map( D => reg_out_37_port, CLK => clk, 
                           SN => n38, Q => Ciphertext(37));
   Ciphertext_regx36x : DFFSNQ_X1 port map( D => reg_out_36_port, CLK => clk, 
                           SN => n37, Q => Ciphertext(36));
   Ciphertext_regx35x : DFFSNQ_X1 port map( D => reg_out_35_port, CLK => clk, 
                           SN => n36, Q => Ciphertext(35));
   Ciphertext_regx34x : DFFSNQ_X1 port map( D => reg_out_34_port, CLK => clk, 
                           SN => n35, Q => Ciphertext(34));
   Ciphertext_regx31x : DFFSNQ_X1 port map( D => reg_out_31_port, CLK => clk, 
                           SN => n32, Q => Ciphertext(31));
   Ciphertext_regx29x : DFFSNQ_X1 port map( D => reg_out_29_port, CLK => clk, 
                           SN => n30, Q => Ciphertext(29));
   Ciphertext_regx27x : DFFSNQ_X1 port map( D => reg_out_27_port, CLK => clk, 
                           SN => n28, Q => Ciphertext(27));
   Ciphertext_regx25x : DFFSNQ_X1 port map( D => reg_out_25_port, CLK => clk, 
                           SN => n26, Q => Ciphertext(25));
   Ciphertext_regx24x : DFFSNQ_X1 port map( D => reg_out_24_port, CLK => clk, 
                           SN => n25, Q => Ciphertext(24));
   Ciphertext_regx22x : DFFSNQ_X1 port map( D => reg_out_22_port, CLK => clk, 
                           SN => n23, Q => Ciphertext(22));
   Ciphertext_regx19x : DFFSNQ_X1 port map( D => reg_out_19_port, CLK => clk, 
                           SN => n20, Q => Ciphertext(19));
   Ciphertext_regx18x : DFFSNQ_X1 port map( D => reg_out_18_port, CLK => clk, 
                           SN => n19, Q => Ciphertext(18));
   Ciphertext_regx17x : DFFSNQ_X1 port map( D => reg_out_17_port, CLK => clk, 
                           SN => n18, Q => Ciphertext(17));
   Ciphertext_regx16x : DFFSNQ_X1 port map( D => reg_out_16_port, CLK => clk, 
                           SN => n17, Q => Ciphertext(16));
   Ciphertext_regx15x : DFFSNQ_X1 port map( D => reg_out_15_port, CLK => clk, 
                           SN => n16, Q => Ciphertext(15));
   Ciphertext_regx13x : DFFSNQ_X1 port map( D => reg_out_13_port, CLK => clk, 
                           SN => n14, Q => Ciphertext(13));
   Ciphertext_regx12x : DFFSNQ_X1 port map( D => reg_out_12_port, CLK => clk, 
                           SN => n13, Q => Ciphertext(12));
   Ciphertext_regx11x : DFFSNQ_X1 port map( D => reg_out_11_port, CLK => clk, 
                           SN => n12, Q => Ciphertext(11));
   Ciphertext_regx7x : DFFSNQ_X1 port map( D => reg_out_7_port, CLK => clk, SN 
                           => n8, Q => Ciphertext(7));
   Ciphertext_regx6x : DFFSNQ_X1 port map( D => reg_out_6_port, CLK => clk, SN 
                           => n7, Q => Ciphertext(6));
   Ciphertext_regx5x : DFFSNQ_X1 port map( D => reg_out_5_port, CLK => clk, SN 
                           => n6, Q => Ciphertext(5));
   Ciphertext_regx4x : DFFSNQ_X1 port map( D => reg_out_4_port, CLK => clk, SN 
                           => n5, Q => Ciphertext(4));
   Ciphertext_regx2x : DFFSNQ_X1 port map( D => reg_out_2_port, CLK => clk, SN 
                           => n3, Q => Ciphertext(2));
   Ciphertext_regx1x : DFFSNQ_X1 port map( D => reg_out_1_port, CLK => clk, SN 
                           => n2, Q => Ciphertext(1));
   n2 <= '1';
   n3 <= '1';
   n5 <= '1';
   n6 <= '1';
   n7 <= '1';
   n8 <= '1';
   n12 <= '1';
   n13 <= '1';
   n14 <= '1';
   n16 <= '1';
   n17 <= '1';
   n18 <= '1';
   n19 <= '1';
   n20 <= '1';
   n23 <= '1';
   n25 <= '1';
   n26 <= '1';
   n28 <= '1';
   n30 <= '1';
   n32 <= '1';
   n35 <= '1';
   n36 <= '1';
   n37 <= '1';
   n38 <= '1';
   n39 <= '1';
   n41 <= '1';
   n42 <= '1';
   n43 <= '1';
   n44 <= '1';
   n45 <= '1';
   n46 <= '1';
   n47 <= '1';
   n48 <= '1';
   n49 <= '1';
   n51 <= '1';
   n52 <= '1';
   n53 <= '1';
   n54 <= '1';
   n56 <= '1';
   n61 <= '1';
   n62 <= '1';
   n63 <= '1';
   n64 <= '1';
   n65 <= '1';
   n66 <= '1';
   n67 <= '1';
   n68 <= '1';
   n69 <= '1';
   n70 <= '1';
   n71 <= '1';
   n72 <= '1';
   n74 <= '1';
   n75 <= '1';
   n77 <= '1';
   n78 <= '1';
   n79 <= '1';
   n80 <= '1';
   n81 <= '1';
   n82 <= '1';
   n83 <= '1';
   n84 <= '1';
   n85 <= '1';
   n86 <= '1';
   n87 <= '1';
   n90 <= '1';
   n91 <= '1';
   n92 <= '1';
   n93 <= '1';
   n94 <= '1';
   n97 <= '1';
   n99 <= '1';
   n103 <= '1';
   n104 <= '1';
   n105 <= '1';
   n106 <= '1';
   n107 <= '1';
   n108 <= '1';
   n109 <= '1';
   n110 <= '1';
   n111 <= '1';
   n113 <= '1';
   n114 <= '1';
   n116 <= '1';
   n119 <= '1';
   n120 <= '1';
   n122 <= '1';
   n123 <= '1';
   n124 <= '1';
   n127 <= '1';
   n128 <= '1';
   n129 <= '1';
   n130 <= '1';
   n135 <= '1';
   n136 <= '1';
   n139 <= '1';
   n140 <= '1';
   n141 <= '1';
   n142 <= '1';
   n143 <= '1';
   n145 <= '1';
   n146 <= '1';
   n148 <= '1';
   n149 <= '1';
   n150 <= '1';
   n151 <= '1';
   n152 <= '1';
   n156 <= '1';
   n157 <= '1';
   n158 <= '1';
   n159 <= '1';
   n162 <= '1';
   n164 <= '1';
   n167 <= '1';
   n168 <= '1';
   n169 <= '1';
   n171 <= '1';
   n173 <= '1';
   n174 <= '1';
   n176 <= '1';
   n177 <= '1';
   n178 <= '1';
   n179 <= '1';
   n180 <= '1';
   n182 <= '1';
   n184 <= '1';
   n185 <= '1';
   n188 <= '1';
   n189 <= '1';
   n192 <= '1';
   n193 <= '1';
   n194 <= '1';
   n195 <= '1';
   n196 <= '1';
   n197 <= '1';
   n198 <= '1';
   n199 <= '1';
   n200 <= '1';
   n201 <= '1';
   n202 <= '1';
   n203 <= '1';
   n204 <= '1';
   n205 <= '1';
   n206 <= '1';
   n207 <= '1';
   n208 <= '1';
   n209 <= '1';
   n210 <= '1';
   n211 <= '1';
   n212 <= '1';
   n213 <= '1';
   n214 <= '1';
   n215 <= '1';
   n216 <= '1';
   n217 <= '1';
   n218 <= '1';
   n219 <= '1';
   n220 <= '1';
   n221 <= '1';
   n222 <= '1';
   n223 <= '1';
   n224 <= '1';
   n225 <= '1';
   n226 <= '1';
   n227 <= '1';
   n228 <= '1';
   n229 <= '1';
   n231 <= '1';
   n232 <= '1';
   n233 <= '1';
   n234 <= '1';
   n235 <= '1';
   n236 <= '1';
   n237 <= '1';
   n238 <= '1';
   n239 <= '1';
   n240 <= '1';
   n241 <= '1';
   n242 <= '1';
   n243 <= '1';
   n244 <= '1';
   n245 <= '1';
   n246 <= '1';
   n247 <= '1';
   n248 <= '1';
   n249 <= '1';
   n250 <= '1';
   n251 <= '1';
   n252 <= '1';
   n253 <= '1';
   n254 <= '1';
   n255 <= '1';
   n256 <= '1';
   n257 <= '1';
   n258 <= '1';
   n259 <= '1';
   n260 <= '1';
   n261 <= '1';
   n262 <= '1';
   n263 <= '1';
   n264 <= '1';
   n265 <= '1';
   n266 <= '1';
   n267 <= '1';
   n268 <= '1';
   n269 <= '1';
   n270 <= '1';
   n271 <= '1';
   n272 <= '1';
   n273 <= '1';
   n274 <= '1';
   n275 <= '1';
   n276 <= '1';
   n277 <= '1';
   n278 <= '1';
   n279 <= '1';
   n280 <= '1';
   n281 <= '1';
   n282 <= '1';
   n283 <= '1';
   n284 <= '1';
   n285 <= '1';
   n286 <= '1';
   n287 <= '1';
   n288 <= '1';
   n289 <= '1';
   n290 <= '1';
   n291 <= '1';
   n292 <= '1';
   n293 <= '1';
   n294 <= '1';
   n295 <= '1';
   n296 <= '1';
   n297 <= '1';
   n298 <= '1';
   n299 <= '1';
   n300 <= '1';
   n301 <= '1';
   n302 <= '1';
   n303 <= '1';
   n304 <= '1';
   n305 <= '1';
   n306 <= '1';
   n307 <= '1';
   n308 <= '1';
   n309 <= '1';
   n310 <= '1';
   n311 <= '1';
   n312 <= '1';
   n313 <= '1';
   n314 <= '1';
   n315 <= '1';
   n316 <= '1';
   n317 <= '1';
   n318 <= '1';
   n319 <= '1';
   n320 <= '1';
   n321 <= '1';
   n322 <= '1';
   n323 <= '1';
   n324 <= '1';
   n325 <= '1';
   n326 <= '1';
   n327 <= '1';
   n328 <= '1';
   n329 <= '1';
   n330 <= '1';
   n331 <= '1';
   n332 <= '1';
   n333 <= '1';
   n334 <= '1';
   n335 <= '1';
   n336 <= '1';
   n337 <= '1';
   n338 <= '1';
   n339 <= '1';
   n340 <= '1';
   n341 <= '1';
   n342 <= '1';
   n343 <= '1';
   n345 <= '1';
   n346 <= '1';
   n347 <= '1';
   n348 <= '1';
   n349 <= '1';
   n350 <= '1';
   n351 <= '1';
   n352 <= '1';
   n353 <= '1';
   n354 <= '1';
   n355 <= '1';
   n356 <= '1';
   n357 <= '1';
   n358 <= '1';
   n359 <= '1';
   n360 <= '1';
   n361 <= '1';
   n362 <= '1';
   n363 <= '1';
   n364 <= '1';
   n365 <= '1';
   n366 <= '1';
   n367 <= '1';
   n368 <= '1';
   n369 <= '1';
   n370 <= '1';
   n371 <= '1';
   n372 <= '1';
   n373 <= '1';
   n374 <= '1';
   n375 <= '1';
   n376 <= '1';
   n377 <= '1';
   n378 <= '1';
   n379 <= '1';
   n380 <= '1';
   n381 <= '1';
   n382 <= '1';
   n383 <= '1';
   n384 <= '1';
   n385 <= '1';
   n386 <= '1';
   n387 <= '1';
   n388 <= '1';
   n389 <= '1';
   n390 <= '1';
   n391 <= '1';
   n392 <= '1';
   n393 <= '1';
   n394 <= '1';
   n395 <= '1';
   n396 <= '1';
   n397 <= '1';
   n398 <= '1';
   n399 <= '1';
   n400 <= '1';
   n401 <= '1';
   n402 <= '1';
   n403 <= '1';
   n404 <= '1';
   n405 <= '1';
   n406 <= '1';
   n407 <= '1';
   n408 <= '1';
   n409 <= '1';
   n413 <= '1';
   n415 <= '1';
   n416 <= '1';
   n417 <= '1';
   n418 <= '1';
   n419 <= '1';
   n421 <= '1';
   n422 <= '1';
   n423 <= '1';
   n424 <= '1';
   n425 <= '1';
   n426 <= '1';
   n427 <= '1';
   n428 <= '1';
   n429 <= '1';
   n430 <= '1';
   n431 <= '1';
   n432 <= '1';
   n433 <= '1';
   n434 <= '1';
   n435 <= '1';
   n436 <= '1';
   n437 <= '1';
   n438 <= '1';
   n439 <= '1';
   n440 <= '1';
   n441 <= '1';
   n442 <= '1';
   n443 <= '1';
   n445 <= '1';
   n446 <= '1';
   n447 <= '1';
   n448 <= '1';
   n449 <= '1';
   n450 <= '1';
   n451 <= '1';
   n452 <= '1';
   n453 <= '1';
   n454 <= '1';
   n455 <= '1';
   n456 <= '1';
   n457 <= '1';
   n458 <= '1';
   n459 <= '1';
   n460 <= '1';
   n461 <= '1';
   n462 <= '1';
   n463 <= '1';
   n464 <= '1';
   n465 <= '1';
   n466 <= '1';
   n467 <= '1';
   n469 <= '1';
   n470 <= '1';
   n471 <= '1';
   n472 <= '1';
   n473 <= '1';
   n474 <= '1';
   n475 <= '1';
   n476 <= '1';
   n477 <= '1';
   n478 <= '1';
   n479 <= '1';
   n480 <= '1';
   n481 <= '1';
   n482 <= '1';
   n483 <= '1';
   n484 <= '1';
   n485 <= '1';
   n486 <= '1';
   n487 <= '1';
   n488 <= '1';
   n489 <= '1';
   n490 <= '1';
   n491 <= '1';
   n492 <= '1';
   n493 <= '1';
   n494 <= '1';
   n495 <= '1';
   n496 <= '1';
   n497 <= '1';
   n498 <= '1';
   n499 <= '1';
   n500 <= '1';
   n501 <= '1';
   n502 <= '1';
   n503 <= '1';
   n504 <= '1';
   n505 <= '1';
   n506 <= '1';
   n507 <= '1';
   n508 <= '1';
   n509 <= '1';
   n511 <= '1';
   n512 <= '1';
   n513 <= '1';
   n514 <= '1';
   n515 <= '1';
   n516 <= '1';
   n517 <= '1';
   n518 <= '1';
   n519 <= '1';
   n520 <= '1';
   n521 <= '1';
   n522 <= '1';
   n523 <= '1';
   n524 <= '1';
   n526 <= '1';
   n527 <= '1';
   n528 <= '1';
   n529 <= '1';
   n530 <= '1';
   n532 <= '1';
   n533 <= '1';
   n534 <= '1';
   n535 <= '1';
   n536 <= '1';
   n537 <= '1';
   n538 <= '1';
   n539 <= '1';
   n540 <= '1';
   n541 <= '1';
   n542 <= '1';
   n543 <= '1';
   n544 <= '1';
   n545 <= '1';
   n546 <= '1';
   n547 <= '1';
   n548 <= '1';
   n549 <= '1';
   n550 <= '1';
   n551 <= '1';
   n552 <= '1';
   n553 <= '1';
   n555 <= '1';
   n556 <= '1';
   n557 <= '1';
   n558 <= '1';
   n559 <= '1';
   n560 <= '1';
   n561 <= '1';
   n562 <= '1';
   n563 <= '1';
   n564 <= '1';
   n565 <= '1';
   n566 <= '1';
   n567 <= '1';
   n568 <= '1';
   n569 <= '1';
   n570 <= '1';
   n571 <= '1';
   n572 <= '1';
   n573 <= '1';
   n574 <= '1';
   n575 <= '1';
   Ciphertext_regx160x : DFFRNQ_X1 port map( D => reg_out_160_port, CLK => clk,
                           RN => n616, Q => Ciphertext(160));
   Ciphertext_regx159x : DFFRNQ_X1 port map( D => reg_out_159_port, CLK => clk,
                           RN => n615, Q => Ciphertext(159));
   Ciphertext_regx10x : DFFRNQ_X1 port map( D => reg_out_10_port, CLK => clk, 
                           RN => n614, Q => Ciphertext(10));
   reg_in_regx125x : DFFRNQ_X1 port map( D => Plaintext(125), CLK => clk, RN =>
                           n613, Q => reg_in_125_port);
   Ciphertext_regx132x : DFFRNQ_X1 port map( D => reg_out_132_port, CLK => clk,
                           RN => n612, Q => Ciphertext(132));
   Ciphertext_regx49x : DFFRNQ_X1 port map( D => reg_out_49_port, CLK => clk, 
                           RN => n611, Q => Ciphertext(49));
   Ciphertext_regx33x : DFFRNQ_X1 port map( D => reg_out_33_port, CLK => clk, 
                           RN => n610, Q => Ciphertext(33));
   Ciphertext_regx3x : DFFRNQ_X1 port map( D => reg_out_3_port, CLK => clk, RN 
                           => n609, Q => Ciphertext(3));
   Ciphertext_regx185x : DFFRNQ_X1 port map( D => reg_out_185_port, CLK => clk,
                           RN => n608, Q => Ciphertext(185));
   reg_in_regx25x : DFFRNQ_X1 port map( D => Plaintext(25), CLK => clk, RN => 
                           n606, Q => reg_in_25_port);
   Ciphertext_regx99x : DFFRNQ_X1 port map( D => reg_out_99_port, CLK => clk, 
                           RN => n605, Q => Ciphertext(99));
   Ciphertext_regx116x : DFFRNQ_X1 port map( D => reg_out_116_port, CLK => clk,
                           RN => n604, Q => Ciphertext(116));
   Ciphertext_regx32x : DFFRNQ_X1 port map( D => reg_out_32_port, CLK => clk, 
                           RN => n603, Q => Ciphertext(32));
   Ciphertext_regx125x : DFFRNQ_X1 port map( D => reg_out_125_port, CLK => clk,
                           RN => n602, Q => Ciphertext(125));
   Ciphertext_regx94x : DFFRNQ_X1 port map( D => reg_out_94_port, CLK => clk, 
                           RN => n601, Q => Ciphertext(94));
   Ciphertext_regx143x : DFFRNQ_X1 port map( D => reg_out_143_port, CLK => clk,
                           RN => n600, Q => Ciphertext(143));
   Ciphertext_regx75x : DFFRNQ_X1 port map( D => reg_out_75_port, CLK => clk, 
                           RN => n599, Q => Ciphertext(75));
   Ciphertext_regx114x : DFFRNQ_X1 port map( D => reg_out_114_port, CLK => clk,
                           RN => n598, Q => Ciphertext(114));
   Ciphertext_regx186x : DFFRNQ_X1 port map( D => reg_out_186_port, CLK => clk,
                           RN => n597, Q => Ciphertext(186));
   Ciphertext_regx21x : DFFRNQ_X1 port map( D => reg_out_21_port, CLK => clk, 
                           RN => n596, Q => Ciphertext(21));
   Ciphertext_regx154x : DFFRNQ_X1 port map( D => reg_out_154_port, CLK => clk,
                           RN => n595, Q => Ciphertext(154));
   Ciphertext_regx14x : DFFRNQ_X1 port map( D => reg_out_14_port, CLK => clk, 
                           RN => n594, Q => Ciphertext(14));
   reg_in_regx140x : DFFRNQ_X1 port map( D => Plaintext(140), CLK => clk, RN =>
                           n593, Q => reg_in_140_port);
   Ciphertext_regx20x : DFFRNQ_X1 port map( D => reg_out_20_port, CLK => clk, 
                           RN => n592, Q => Ciphertext(20));
   reg_in_regx35x : DFFRNQ_X1 port map( D => Plaintext(35), CLK => clk, RN => 
                           n591, Q => reg_in_35_port);
   Ciphertext_regx124x : DFFRNQ_X1 port map( D => reg_out_124_port, CLK => clk,
                           RN => n590, Q => Ciphertext(124));
   Ciphertext_regx136x : DFFRNQ_X1 port map( D => reg_out_136_port, CLK => clk,
                           RN => n589, Q => Ciphertext(136));
   Ciphertext_regx9x : DFFRNQ_X1 port map( D => reg_out_9_port, CLK => clk, RN 
                           => n588, Q => Ciphertext(9));
   Ciphertext_regx28x : DFFRNQ_X1 port map( D => reg_out_28_port, CLK => clk, 
                           RN => n587, Q => Ciphertext(28));
   Ciphertext_regx23x : DFFRNQ_X1 port map( D => reg_out_23_port, CLK => clk, 
                           RN => n586, Q => Ciphertext(23));
   Ciphertext_regx111x : DFFRNQ_X1 port map( D => reg_out_111_port, CLK => clk,
                           RN => n584, Q => Ciphertext(111));
   Ciphertext_regx30x : DFFRNQ_X1 port map( D => reg_out_30_port, CLK => clk, 
                           RN => n583, Q => Ciphertext(30));
   Ciphertext_regx101x : DFFRNQ_X1 port map( D => reg_out_101_port, CLK => clk,
                           RN => n582, Q => Ciphertext(101));
   Ciphertext_regx87x : DFFRNQ_X1 port map( D => reg_out_87_port, CLK => clk, 
                           RN => n581, Q => Ciphertext(87));
   reg_in_regx169x : DFFRNQ_X1 port map( D => Plaintext(169), CLK => clk, RN =>
                           n580, Q => reg_in_169_port);
   Ciphertext_regx117x : DFFRNQ_X1 port map( D => reg_out_117_port, CLK => clk,
                           RN => n579, Q => Ciphertext(117));
   Ciphertext_regx133x : DFFRNQ_X1 port map( D => reg_out_133_port, CLK => clk,
                           RN => n578, Q => Ciphertext(133));
   Ciphertext_regx146x : DFFRNQ_X1 port map( D => reg_out_146_port, CLK => clk,
                           RN => n577, Q => Ciphertext(146));
   n577 <= '1';
   n578 <= '1';
   n579 <= '1';
   n580 <= '1';
   n581 <= '1';
   n582 <= '1';
   n583 <= '1';
   n584 <= '1';
   n586 <= '1';
   n587 <= '1';
   n588 <= '1';
   n589 <= '1';
   n590 <= '1';
   n591 <= '1';
   n592 <= '1';
   n593 <= '1';
   n594 <= '1';
   n595 <= '1';
   n596 <= '1';
   n597 <= '1';
   n598 <= '1';
   n599 <= '1';
   n600 <= '1';
   n601 <= '1';
   n602 <= '1';
   n603 <= '1';
   n604 <= '1';
   n605 <= '1';
   n606 <= '1';
   n608 <= '1';
   n609 <= '1';
   n610 <= '1';
   n611 <= '1';
   n612 <= '1';
   n613 <= '1';
   n614 <= '1';
   n615 <= '1';
   n616 <= '1';
   Ciphertext_regx88x : DFFSNQ_X1 port map( D => reg_out_88_port, CLK => clk, 
                           SN => n644, Q => Ciphertext(88));
   Ciphertext_regx72x : DFFRNQ_X1 port map( D => reg_out_72_port, CLK => clk, 
                           RN => n643, Q => Ciphertext(72));
   Ciphertext_regx100x : DFFRNQ_X1 port map( D => reg_out_100_port, CLK => clk,
                           RN => n642, Q => Ciphertext(100));
   Ciphertext_regx130x : DFFRNQ_X1 port map( D => reg_out_130_port, CLK => clk,
                           RN => n641, Q => Ciphertext(130));
   Ciphertext_regx59x : DFFRNQ_X1 port map( D => reg_out_59_port, CLK => clk, 
                           RN => n640, Q => Ciphertext(59));
   Ciphertext_regx0x : DFFRNQ_X1 port map( D => reg_out_0_port, CLK => clk, RN 
                           => n639, Q => Ciphertext(0));
   Ciphertext_regx58x : DFFRNQ_X1 port map( D => reg_out_58_port, CLK => clk, 
                           RN => n638, Q => Ciphertext(58));
   Ciphertext_regx26x : DFFRNQ_X1 port map( D => reg_out_26_port, CLK => clk, 
                           RN => n637, Q => Ciphertext(26));
   Ciphertext_regx131x : DFFRNQ_X1 port map( D => reg_out_131_port, CLK => clk,
                           RN => n636, Q => Ciphertext(131));
   Ciphertext_regx189x : DFFRNQ_X1 port map( D => reg_out_189_port, CLK => clk,
                           RN => n635, Q => Ciphertext(189));
   Ciphertext_regx56x : DFFRNQ_X1 port map( D => reg_out_56_port, CLK => clk, 
                           RN => n633, Q => Ciphertext(56));
   Ciphertext_regx54x : DFFRNQ_X1 port map( D => reg_out_54_port, CLK => clk, 
                           RN => n632, Q => Ciphertext(54));
   Ciphertext_regx153x : DFFRNQ_X1 port map( D => reg_out_153_port, CLK => clk,
                           RN => n631, Q => Ciphertext(153));
   Ciphertext_regx174x : DFFRNQ_X1 port map( D => reg_out_174_port, CLK => clk,
                           RN => n630, Q => Ciphertext(174));
   reg_in_regx146x : DFFRNQ_X1 port map( D => Plaintext(146), CLK => clk, RN =>
                           n629, Q => reg_in_146_port);
   Ciphertext_regx171x : DFFRNQ_X1 port map( D => reg_out_171_port, CLK => clk,
                           RN => n628, Q => Ciphertext(171));
   Ciphertext_regx180x : DFFRNQ_X1 port map( D => reg_out_180_port, CLK => clk,
                           RN => n627, Q => Ciphertext(180));
   reg_key_regx37x : DFFRNQ_X1 port map( D => Key(37), CLK => clk, RN => n626, 
                           Q => reg_key_37_port);
   Ciphertext_regx182x : DFFRNQ_X1 port map( D => reg_out_182_port, CLK => clk,
                           RN => n625, Q => Ciphertext(182));
   reg_in_regx83x : DFFRNQ_X1 port map( D => Plaintext(83), CLK => clk, RN => 
                           n624, Q => reg_in_83_port);
   Ciphertext_regx152x : DFFRNQ_X1 port map( D => reg_out_152_port, CLK => clk,
                           RN => n623, Q => Ciphertext(152));
   Ciphertext_regx120x : DFFRNQ_X1 port map( D => reg_out_120_port, CLK => clk,
                           RN => n622, Q => Ciphertext(120));
   Ciphertext_regx137x : DFFRNQ_X1 port map( D => reg_out_137_port, CLK => clk,
                           RN => n621, Q => Ciphertext(137));
   reg_in_regx191x : DFFSNQ_X1 port map( D => Plaintext(191), CLK => clk, SN =>
                           n620, Q => reg_in_191_port);
   Ciphertext_regx190x : DFFRNQ_X1 port map( D => reg_out_190_port, CLK => clk,
                           RN => n619, Q => Ciphertext(190));
   Ciphertext_regx97x : DFFRNQ_X1 port map( D => reg_out_97_port, CLK => clk, 
                           RN => n618, Q => Ciphertext(97));
   reg_in_regx59x : DFFRNQ_X1 port map( D => Plaintext(59), CLK => clk, RN => 
                           n617, Q => reg_in_59_port);
   n617 <= '1';
   n618 <= '1';
   n619 <= '1';
   n620 <= '1';
   n621 <= '1';
   n622 <= '1';
   n623 <= '1';
   n624 <= '1';
   n625 <= '1';
   n626 <= '1';
   n627 <= '1';
   n628 <= '1';
   n629 <= '1';
   n630 <= '1';
   n631 <= '1';
   n632 <= '1';
   n633 <= '1';
   n635 <= '1';
   n636 <= '1';
   n637 <= '1';
   n638 <= '1';
   n639 <= '1';
   n640 <= '1';
   n641 <= '1';
   n642 <= '1';
   n643 <= '1';
   n644 <= '1';
   SPEEDY_instance : SPEEDY_Rounds7_0 port map( Plaintext(191) => 
                           reg_in_191_port, Plaintext(190) => reg_in_190_port, 
                           Plaintext(189) => reg_in_189_port, Plaintext(188) =>
                           reg_in_188_port, Plaintext(187) => reg_in_187_port, 
                           Plaintext(186) => reg_in_186_port, Plaintext(185) =>
                           reg_in_185_port, Plaintext(184) => reg_in_184_port, 
                           Plaintext(183) => reg_in_183_port, Plaintext(182) =>
                           reg_in_182_port, Plaintext(181) => reg_in_181_port, 
                           Plaintext(180) => reg_in_180_port, Plaintext(179) =>
                           reg_in_179_port, Plaintext(178) => reg_in_178_port, 
                           Plaintext(177) => reg_in_177_port, Plaintext(176) =>
                           reg_in_176_port, Plaintext(175) => reg_in_175_port, 
                           Plaintext(174) => reg_in_174_port, Plaintext(173) =>
                           reg_in_173_port, Plaintext(172) => reg_in_172_port, 
                           Plaintext(171) => reg_in_171_port, Plaintext(170) =>
                           reg_in_170_port, Plaintext(169) => reg_in_169_port, 
                           Plaintext(168) => reg_in_168_port, Plaintext(167) =>
                           reg_in_167_port, Plaintext(166) => reg_in_166_port, 
                           Plaintext(165) => reg_in_165_port, Plaintext(164) =>
                           reg_in_164_port, Plaintext(163) => reg_in_163_port, 
                           Plaintext(162) => reg_in_162_port, Plaintext(161) =>
                           reg_in_161_port, Plaintext(160) => reg_in_160_port, 
                           Plaintext(159) => reg_in_159_port, Plaintext(158) =>
                           reg_in_158_port, Plaintext(157) => reg_in_157_port, 
                           Plaintext(156) => reg_in_156_port, Plaintext(155) =>
                           reg_in_155_port, Plaintext(154) => reg_in_154_port, 
                           Plaintext(153) => reg_in_153_port, Plaintext(152) =>
                           reg_in_152_port, Plaintext(151) => reg_in_151_port, 
                           Plaintext(150) => reg_in_150_port, Plaintext(149) =>
                           reg_in_149_port, Plaintext(148) => reg_in_148_port, 
                           Plaintext(147) => reg_in_147_port, Plaintext(146) =>
                           reg_in_146_port, Plaintext(145) => reg_in_145_port, 
                           Plaintext(144) => reg_in_144_port, Plaintext(143) =>
                           reg_in_143_port, Plaintext(142) => reg_in_142_port, 
                           Plaintext(141) => reg_in_141_port, Plaintext(140) =>
                           reg_in_140_port, Plaintext(139) => reg_in_139_port, 
                           Plaintext(138) => reg_in_138_port, Plaintext(137) =>
                           reg_in_137_port, Plaintext(136) => reg_in_136_port, 
                           Plaintext(135) => reg_in_135_port, Plaintext(134) =>
                           reg_in_134_port, Plaintext(133) => reg_in_133_port, 
                           Plaintext(132) => reg_in_132_port, Plaintext(131) =>
                           reg_in_131_port, Plaintext(130) => reg_in_130_port, 
                           Plaintext(129) => reg_in_129_port, Plaintext(128) =>
                           reg_in_128_port, Plaintext(127) => reg_in_127_port, 
                           Plaintext(126) => reg_in_126_port, Plaintext(125) =>
                           reg_in_125_port, Plaintext(124) => reg_in_124_port, 
                           Plaintext(123) => reg_in_123_port, Plaintext(122) =>
                           reg_in_122_port, Plaintext(121) => reg_in_121_port, 
                           Plaintext(120) => reg_in_120_port, Plaintext(119) =>
                           reg_in_119_port, Plaintext(118) => reg_in_118_port, 
                           Plaintext(117) => reg_in_117_port, Plaintext(116) =>
                           reg_in_116_port, Plaintext(115) => reg_in_115_port, 
                           Plaintext(114) => reg_in_114_port, Plaintext(113) =>
                           reg_in_113_port, Plaintext(112) => reg_in_112_port, 
                           Plaintext(111) => reg_in_111_port, Plaintext(110) =>
                           reg_in_110_port, Plaintext(109) => reg_in_109_port, 
                           Plaintext(108) => reg_in_108_port, Plaintext(107) =>
                           reg_in_107_port, Plaintext(106) => reg_in_106_port, 
                           Plaintext(105) => reg_in_105_port, Plaintext(104) =>
                           reg_in_104_port, Plaintext(103) => reg_in_103_port, 
                           Plaintext(102) => reg_in_102_port, Plaintext(101) =>
                           reg_in_101_port, Plaintext(100) => reg_in_100_port, 
                           Plaintext(99) => reg_in_99_port, Plaintext(98) => 
                           reg_in_98_port, Plaintext(97) => reg_in_97_port, 
                           Plaintext(96) => reg_in_96_port, Plaintext(95) => 
                           reg_in_95_port, Plaintext(94) => reg_in_94_port, 
                           Plaintext(93) => reg_in_93_port, Plaintext(92) => 
                           reg_in_92_port, Plaintext(91) => reg_in_91_port, 
                           Plaintext(90) => reg_in_90_port, Plaintext(89) => 
                           reg_in_89_port, Plaintext(88) => reg_in_88_port, 
                           Plaintext(87) => reg_in_87_port, Plaintext(86) => 
                           reg_in_86_port, Plaintext(85) => reg_in_85_port, 
                           Plaintext(84) => reg_in_84_port, Plaintext(83) => 
                           reg_in_83_port, Plaintext(82) => reg_in_82_port, 
                           Plaintext(81) => reg_in_81_port, Plaintext(80) => 
                           reg_in_80_port, Plaintext(79) => reg_in_79_port, 
                           Plaintext(78) => reg_in_78_port, Plaintext(77) => 
                           reg_in_77_port, Plaintext(76) => reg_in_76_port, 
                           Plaintext(75) => reg_in_75_port, Plaintext(74) => 
                           reg_in_74_port, Plaintext(73) => reg_in_73_port, 
                           Plaintext(72) => reg_in_72_port, Plaintext(71) => 
                           reg_in_71_port, Plaintext(70) => reg_in_70_port, 
                           Plaintext(69) => reg_in_69_port, Plaintext(68) => 
                           reg_in_68_port, Plaintext(67) => reg_in_67_port, 
                           Plaintext(66) => reg_in_66_port, Plaintext(65) => 
                           reg_in_65_port, Plaintext(64) => reg_in_64_port, 
                           Plaintext(63) => reg_in_63_port, Plaintext(62) => 
                           reg_in_62_port, Plaintext(61) => reg_in_61_port, 
                           Plaintext(60) => reg_in_60_port, Plaintext(59) => 
                           reg_in_59_port, Plaintext(58) => reg_in_58_port, 
                           Plaintext(57) => reg_in_57_port, Plaintext(56) => 
                           reg_in_56_port, Plaintext(55) => reg_in_55_port, 
                           Plaintext(54) => reg_in_54_port, Plaintext(53) => 
                           reg_in_53_port, Plaintext(52) => reg_in_52_port, 
                           Plaintext(51) => reg_in_51_port, Plaintext(50) => 
                           reg_in_50_port, Plaintext(49) => reg_in_49_port, 
                           Plaintext(48) => reg_in_48_port, Plaintext(47) => 
                           reg_in_47_port, Plaintext(46) => reg_in_46_port, 
                           Plaintext(45) => reg_in_45_port, Plaintext(44) => 
                           reg_in_44_port, Plaintext(43) => reg_in_43_port, 
                           Plaintext(42) => reg_in_42_port, Plaintext(41) => 
                           reg_in_41_port, Plaintext(40) => reg_in_40_port, 
                           Plaintext(39) => reg_in_39_port, Plaintext(38) => 
                           reg_in_38_port, Plaintext(37) => reg_in_37_port, 
                           Plaintext(36) => reg_in_36_port, Plaintext(35) => 
                           reg_in_35_port, Plaintext(34) => reg_in_34_port, 
                           Plaintext(33) => reg_in_33_port, Plaintext(32) => 
                           reg_in_32_port, Plaintext(31) => reg_in_31_port, 
                           Plaintext(30) => reg_in_30_port, Plaintext(29) => 
                           reg_in_29_port, Plaintext(28) => reg_in_28_port, 
                           Plaintext(27) => reg_in_27_port, Plaintext(26) => 
                           reg_in_26_port, Plaintext(25) => reg_in_25_port, 
                           Plaintext(24) => reg_in_24_port, Plaintext(23) => 
                           reg_in_23_port, Plaintext(22) => reg_in_22_port, 
                           Plaintext(21) => reg_in_21_port, Plaintext(20) => 
                           reg_in_20_port, Plaintext(19) => reg_in_19_port, 
                           Plaintext(18) => reg_in_18_port, Plaintext(17) => 
                           reg_in_17_port, Plaintext(16) => reg_in_16_port, 
                           Plaintext(15) => reg_in_15_port, Plaintext(14) => 
                           reg_in_14_port, Plaintext(13) => reg_in_13_port, 
                           Plaintext(12) => reg_in_12_port, Plaintext(11) => 
                           reg_in_11_port, Plaintext(10) => reg_in_10_port, 
                           Plaintext(9) => reg_in_9_port, Plaintext(8) => 
                           reg_in_8_port, Plaintext(7) => reg_in_7_port, 
                           Plaintext(6) => reg_in_6_port, Plaintext(5) => 
                           reg_in_5_port, Plaintext(4) => reg_in_4_port, 
                           Plaintext(3) => reg_in_3_port, Plaintext(2) => 
                           reg_in_2_port, Plaintext(1) => reg_in_1_port, 
                           Plaintext(0) => reg_in_0_port, Key(191) => 
                           reg_key_191_port, Key(190) => reg_key_190_port, 
                           Key(189) => reg_key_189_port, Key(188) => 
                           reg_key_188_port, Key(187) => reg_key_187_port, 
                           Key(186) => reg_key_186_port, Key(185) => 
                           reg_key_185_port, Key(184) => reg_key_184_port, 
                           Key(183) => reg_key_183_port, Key(182) => 
                           reg_key_182_port, Key(181) => reg_key_181_port, 
                           Key(180) => reg_key_180_port, Key(179) => 
                           reg_key_179_port, Key(178) => reg_key_178_port, 
                           Key(177) => reg_key_177_port, Key(176) => 
                           reg_key_176_port, Key(175) => reg_key_175_port, 
                           Key(174) => reg_key_174_port, Key(173) => 
                           reg_key_173_port, Key(172) => reg_key_172_port, 
                           Key(171) => reg_key_171_port, Key(170) => 
                           reg_key_170_port, Key(169) => reg_key_169_port, 
                           Key(168) => reg_key_168_port, Key(167) => 
                           reg_key_167_port, Key(166) => reg_key_166_port, 
                           Key(165) => reg_key_165_port, Key(164) => 
                           reg_key_164_port, Key(163) => reg_key_163_port, 
                           Key(162) => reg_key_162_port, Key(161) => 
                           reg_key_161_port, Key(160) => reg_key_160_port, 
                           Key(159) => reg_key_159_port, Key(158) => 
                           reg_key_158_port, Key(157) => reg_key_157_port, 
                           Key(156) => reg_key_156_port, Key(155) => 
                           reg_key_155_port, Key(154) => reg_key_154_port, 
                           Key(153) => reg_key_153_port, Key(152) => 
                           reg_key_152_port, Key(151) => reg_key_151_port, 
                           Key(150) => reg_key_150_port, Key(149) => 
                           reg_key_149_port, Key(148) => reg_key_148_port, 
                           Key(147) => reg_key_147_port, Key(146) => 
                           reg_key_146_port, Key(145) => reg_key_145_port, 
                           Key(144) => reg_key_144_port, Key(143) => 
                           reg_key_143_port, Key(142) => reg_key_142_port, 
                           Key(141) => reg_key_141_port, Key(140) => 
                           reg_key_140_port, Key(139) => reg_key_139_port, 
                           Key(138) => reg_key_138_port, Key(137) => 
                           reg_key_137_port, Key(136) => reg_key_136_port, 
                           Key(135) => reg_key_135_port, Key(134) => 
                           reg_key_134_port, Key(133) => reg_key_133_port, 
                           Key(132) => reg_key_132_port, Key(131) => 
                           reg_key_131_port, Key(130) => reg_key_130_port, 
                           Key(129) => reg_key_129_port, Key(128) => 
                           reg_key_128_port, Key(127) => reg_key_127_port, 
                           Key(126) => reg_key_126_port, Key(125) => 
                           reg_key_125_port, Key(124) => reg_key_124_port, 
                           Key(123) => reg_key_123_port, Key(122) => 
                           reg_key_122_port, Key(121) => reg_key_121_port, 
                           Key(120) => reg_key_120_port, Key(119) => 
                           reg_key_119_port, Key(118) => reg_key_118_port, 
                           Key(117) => reg_key_117_port, Key(116) => 
                           reg_key_116_port, Key(115) => reg_key_115_port, 
                           Key(114) => reg_key_114_port, Key(113) => 
                           reg_key_113_port, Key(112) => reg_key_112_port, 
                           Key(111) => reg_key_111_port, Key(110) => 
                           reg_key_110_port, Key(109) => reg_key_109_port, 
                           Key(108) => reg_key_108_port, Key(107) => 
                           reg_key_107_port, Key(106) => reg_key_106_port, 
                           Key(105) => reg_key_105_port, Key(104) => 
                           reg_key_104_port, Key(103) => reg_key_103_port, 
                           Key(102) => reg_key_102_port, Key(101) => 
                           reg_key_101_port, Key(100) => reg_key_100_port, 
                           Key(99) => reg_key_99_port, Key(98) => 
                           reg_key_98_port, Key(97) => reg_key_97_port, Key(96)
                           => reg_key_96_port, Key(95) => reg_key_95_port, 
                           Key(94) => reg_key_94_port, Key(93) => 
                           reg_key_93_port, Key(92) => reg_key_92_port, Key(91)
                           => reg_key_91_port, Key(90) => reg_key_90_port, 
                           Key(89) => reg_key_89_port, Key(88) => 
                           reg_key_88_port, Key(87) => reg_key_87_port, Key(86)
                           => reg_key_86_port, Key(85) => reg_key_85_port, 
                           Key(84) => reg_key_84_port, Key(83) => 
                           reg_key_83_port, Key(82) => reg_key_82_port, Key(81)
                           => reg_key_81_port, Key(80) => reg_key_80_port, 
                           Key(79) => reg_key_79_port, Key(78) => 
                           reg_key_78_port, Key(77) => reg_key_77_port, Key(76)
                           => reg_key_76_port, Key(75) => reg_key_75_port, 
                           Key(74) => reg_key_74_port, Key(73) => 
                           reg_key_73_port, Key(72) => reg_key_72_port, Key(71)
                           => reg_key_71_port, Key(70) => reg_key_70_port, 
                           Key(69) => reg_key_69_port, Key(68) => 
                           reg_key_68_port, Key(67) => reg_key_67_port, Key(66)
                           => reg_key_66_port, Key(65) => reg_key_65_port, 
                           Key(64) => reg_key_64_port, Key(63) => 
                           reg_key_63_port, Key(62) => reg_key_62_port, Key(61)
                           => reg_key_61_port, Key(60) => reg_key_60_port, 
                           Key(59) => reg_key_59_port, Key(58) => 
                           reg_key_58_port, Key(57) => reg_key_57_port, Key(56)
                           => reg_key_56_port, Key(55) => reg_key_55_port, 
                           Key(54) => reg_key_54_port, Key(53) => 
                           reg_key_53_port, Key(52) => reg_key_52_port, Key(51)
                           => reg_key_51_port, Key(50) => reg_key_50_port, 
                           Key(49) => reg_key_49_port, Key(48) => 
                           reg_key_48_port, Key(47) => reg_key_47_port, Key(46)
                           => reg_key_46_port, Key(45) => reg_key_45_port, 
                           Key(44) => reg_key_44_port, Key(43) => 
                           reg_key_43_port, Key(42) => reg_key_42_port, Key(41)
                           => reg_key_41_port, Key(40) => reg_key_40_port, 
                           Key(39) => reg_key_39_port, Key(38) => 
                           reg_key_38_port, Key(37) => reg_key_37_port, Key(36)
                           => reg_key_36_port, Key(35) => reg_key_35_port, 
                           Key(34) => reg_key_34_port, Key(33) => 
                           reg_key_33_port, Key(32) => reg_key_32_port, Key(31)
                           => reg_key_31_port, Key(30) => reg_key_30_port, 
                           Key(29) => reg_key_29_port, Key(28) => 
                           reg_key_28_port, Key(27) => reg_key_27_port, Key(26)
                           => reg_key_26_port, Key(25) => reg_key_25_port, 
                           Key(24) => reg_key_24_port, Key(23) => 
                           reg_key_23_port, Key(22) => reg_key_22_port, Key(21)
                           => reg_key_21_port, Key(20) => reg_key_20_port, 
                           Key(19) => reg_key_19_port, Key(18) => 
                           reg_key_18_port, Key(17) => reg_key_17_port, Key(16)
                           => reg_key_16_port, Key(15) => reg_key_15_port, 
                           Key(14) => reg_key_14_port, Key(13) => 
                           reg_key_13_port, Key(12) => reg_key_12_port, Key(11)
                           => reg_key_11_port, Key(10) => reg_key_10_port, 
                           Key(9) => reg_key_9_port, Key(8) => reg_key_8_port, 
                           Key(7) => reg_key_7_port, Key(6) => reg_key_6_port, 
                           Key(5) => reg_key_5_port, Key(4) => reg_key_4_port, 
                           Key(3) => reg_key_3_port, Key(2) => reg_key_2_port, 
                           Key(1) => reg_key_1_port, Key(0) => reg_key_0_port, 
                           Ciphertext(191) => reg_out_191_port, Ciphertext(190)
                           => reg_out_190_port, Ciphertext(189) => 
                           reg_out_189_port, Ciphertext(188) => 
                           reg_out_188_port, Ciphertext(187) => 
                           reg_out_187_port, Ciphertext(186) => 
                           reg_out_186_port, Ciphertext(185) => 
                           reg_out_185_port, Ciphertext(184) => 
                           reg_out_184_port, Ciphertext(183) => 
                           reg_out_183_port, Ciphertext(182) => 
                           reg_out_182_port, Ciphertext(181) => 
                           reg_out_181_port, Ciphertext(180) => 
                           reg_out_180_port, Ciphertext(179) => 
                           reg_out_179_port, Ciphertext(178) => 
                           reg_out_178_port, Ciphertext(177) => 
                           reg_out_177_port, Ciphertext(176) => 
                           reg_out_176_port, Ciphertext(175) => 
                           reg_out_175_port, Ciphertext(174) => 
                           reg_out_174_port, Ciphertext(173) => 
                           reg_out_173_port, Ciphertext(172) => 
                           reg_out_172_port, Ciphertext(171) => 
                           reg_out_171_port, Ciphertext(170) => 
                           reg_out_170_port, Ciphertext(169) => 
                           reg_out_169_port, Ciphertext(168) => 
                           reg_out_168_port, Ciphertext(167) => 
                           reg_out_167_port, Ciphertext(166) => 
                           reg_out_166_port, Ciphertext(165) => 
                           reg_out_165_port, Ciphertext(164) => 
                           reg_out_164_port, Ciphertext(163) => 
                           reg_out_163_port, Ciphertext(162) => 
                           reg_out_162_port, Ciphertext(161) => 
                           reg_out_161_port, Ciphertext(160) => 
                           reg_out_160_port, Ciphertext(159) => 
                           reg_out_159_port, Ciphertext(158) => 
                           reg_out_158_port, Ciphertext(157) => 
                           reg_out_157_port, Ciphertext(156) => 
                           reg_out_156_port, Ciphertext(155) => 
                           reg_out_155_port, Ciphertext(154) => 
                           reg_out_154_port, Ciphertext(153) => 
                           reg_out_153_port, Ciphertext(152) => 
                           reg_out_152_port, Ciphertext(151) => 
                           reg_out_151_port, Ciphertext(150) => 
                           reg_out_150_port, Ciphertext(149) => 
                           reg_out_149_port, Ciphertext(148) => 
                           reg_out_148_port, Ciphertext(147) => 
                           reg_out_147_port, Ciphertext(146) => 
                           reg_out_146_port, Ciphertext(145) => 
                           reg_out_145_port, Ciphertext(144) => 
                           reg_out_144_port, Ciphertext(143) => 
                           reg_out_143_port, Ciphertext(142) => 
                           reg_out_142_port, Ciphertext(141) => 
                           reg_out_141_port, Ciphertext(140) => 
                           reg_out_140_port, Ciphertext(139) => 
                           reg_out_139_port, Ciphertext(138) => 
                           reg_out_138_port, Ciphertext(137) => 
                           reg_out_137_port, Ciphertext(136) => 
                           reg_out_136_port, Ciphertext(135) => 
                           reg_out_135_port, Ciphertext(134) => 
                           reg_out_134_port, Ciphertext(133) => 
                           reg_out_133_port, Ciphertext(132) => 
                           reg_out_132_port, Ciphertext(131) => 
                           reg_out_131_port, Ciphertext(130) => 
                           reg_out_130_port, Ciphertext(129) => 
                           reg_out_129_port, Ciphertext(128) => 
                           reg_out_128_port, Ciphertext(127) => 
                           reg_out_127_port, Ciphertext(126) => 
                           reg_out_126_port, Ciphertext(125) => 
                           reg_out_125_port, Ciphertext(124) => 
                           reg_out_124_port, Ciphertext(123) => 
                           reg_out_123_port, Ciphertext(122) => 
                           reg_out_122_port, Ciphertext(121) => 
                           reg_out_121_port, Ciphertext(120) => 
                           reg_out_120_port, Ciphertext(119) => 
                           reg_out_119_port, Ciphertext(118) => 
                           reg_out_118_port, Ciphertext(117) => 
                           reg_out_117_port, Ciphertext(116) => 
                           reg_out_116_port, Ciphertext(115) => 
                           reg_out_115_port, Ciphertext(114) => 
                           reg_out_114_port, Ciphertext(113) => 
                           reg_out_113_port, Ciphertext(112) => 
                           reg_out_112_port, Ciphertext(111) => 
                           reg_out_111_port, Ciphertext(110) => 
                           reg_out_110_port, Ciphertext(109) => 
                           reg_out_109_port, Ciphertext(108) => 
                           reg_out_108_port, Ciphertext(107) => 
                           reg_out_107_port, Ciphertext(106) => 
                           reg_out_106_port, Ciphertext(105) => 
                           reg_out_105_port, Ciphertext(104) => 
                           reg_out_104_port, Ciphertext(103) => 
                           reg_out_103_port, Ciphertext(102) => 
                           reg_out_102_port, Ciphertext(101) => 
                           reg_out_101_port, Ciphertext(100) => 
                           reg_out_100_port, Ciphertext(99) => reg_out_99_port,
                           Ciphertext(98) => reg_out_98_port, Ciphertext(97) =>
                           reg_out_97_port, Ciphertext(96) => reg_out_96_port, 
                           Ciphertext(95) => reg_out_95_port, Ciphertext(94) =>
                           reg_out_94_port, Ciphertext(93) => reg_out_93_port, 
                           Ciphertext(92) => reg_out_92_port, Ciphertext(91) =>
                           reg_out_91_port, Ciphertext(90) => reg_out_90_port, 
                           Ciphertext(89) => reg_out_89_port, Ciphertext(88) =>
                           reg_out_88_port, Ciphertext(87) => reg_out_87_port, 
                           Ciphertext(86) => reg_out_86_port, Ciphertext(85) =>
                           reg_out_85_port, Ciphertext(84) => reg_out_84_port, 
                           Ciphertext(83) => reg_out_83_port, Ciphertext(82) =>
                           reg_out_82_port, Ciphertext(81) => reg_out_81_port, 
                           Ciphertext(80) => reg_out_80_port, Ciphertext(79) =>
                           reg_out_79_port, Ciphertext(78) => reg_out_78_port, 
                           Ciphertext(77) => reg_out_77_port, Ciphertext(76) =>
                           reg_out_76_port, Ciphertext(75) => reg_out_75_port, 
                           Ciphertext(74) => reg_out_74_port, Ciphertext(73) =>
                           reg_out_73_port, Ciphertext(72) => reg_out_72_port, 
                           Ciphertext(71) => reg_out_71_port, Ciphertext(70) =>
                           reg_out_70_port, Ciphertext(69) => reg_out_69_port, 
                           Ciphertext(68) => reg_out_68_port, Ciphertext(67) =>
                           reg_out_67_port, Ciphertext(66) => reg_out_66_port, 
                           Ciphertext(65) => reg_out_65_port, Ciphertext(64) =>
                           reg_out_64_port, Ciphertext(63) => reg_out_63_port, 
                           Ciphertext(62) => reg_out_62_port, Ciphertext(61) =>
                           reg_out_61_port, Ciphertext(60) => reg_out_60_port, 
                           Ciphertext(59) => reg_out_59_port, Ciphertext(58) =>
                           reg_out_58_port, Ciphertext(57) => reg_out_57_port, 
                           Ciphertext(56) => reg_out_56_port, Ciphertext(55) =>
                           reg_out_55_port, Ciphertext(54) => reg_out_54_port, 
                           Ciphertext(53) => reg_out_53_port, Ciphertext(52) =>
                           reg_out_52_port, Ciphertext(51) => reg_out_51_port, 
                           Ciphertext(50) => reg_out_50_port, Ciphertext(49) =>
                           reg_out_49_port, Ciphertext(48) => reg_out_48_port, 
                           Ciphertext(47) => reg_out_47_port, Ciphertext(46) =>
                           reg_out_46_port, Ciphertext(45) => reg_out_45_port, 
                           Ciphertext(44) => reg_out_44_port, Ciphertext(43) =>
                           reg_out_43_port, Ciphertext(42) => reg_out_42_port, 
                           Ciphertext(41) => reg_out_41_port, Ciphertext(40) =>
                           reg_out_40_port, Ciphertext(39) => reg_out_39_port, 
                           Ciphertext(38) => reg_out_38_port, Ciphertext(37) =>
                           reg_out_37_port, Ciphertext(36) => reg_out_36_port, 
                           Ciphertext(35) => reg_out_35_port, Ciphertext(34) =>
                           reg_out_34_port, Ciphertext(33) => reg_out_33_port, 
                           Ciphertext(32) => reg_out_32_port, Ciphertext(31) =>
                           reg_out_31_port, Ciphertext(30) => reg_out_30_port, 
                           Ciphertext(29) => reg_out_29_port, Ciphertext(28) =>
                           reg_out_28_port, Ciphertext(27) => reg_out_27_port, 
                           Ciphertext(26) => reg_out_26_port, Ciphertext(25) =>
                           reg_out_25_port, Ciphertext(24) => reg_out_24_port, 
                           Ciphertext(23) => reg_out_23_port, Ciphertext(22) =>
                           reg_out_22_port, Ciphertext(21) => reg_out_21_port, 
                           Ciphertext(20) => reg_out_20_port, Ciphertext(19) =>
                           reg_out_19_port, Ciphertext(18) => reg_out_18_port, 
                           Ciphertext(17) => reg_out_17_port, Ciphertext(16) =>
                           reg_out_16_port, Ciphertext(15) => reg_out_15_port, 
                           Ciphertext(14) => reg_out_14_port, Ciphertext(13) =>
                           reg_out_13_port, Ciphertext(12) => reg_out_12_port, 
                           Ciphertext(11) => reg_out_11_port, Ciphertext(10) =>
                           reg_out_10_port, Ciphertext(9) => reg_out_9_port, 
                           Ciphertext(8) => reg_out_8_port, Ciphertext(7) => 
                           reg_out_7_port, Ciphertext(6) => reg_out_6_port, 
                           Ciphertext(5) => reg_out_5_port, Ciphertext(4) => 
                           reg_out_4_port, Ciphertext(3) => reg_out_3_port, 
                           Ciphertext(2) => reg_out_2_port, Ciphertext(1) => 
                           reg_out_1_port, Ciphertext(0) => reg_out_0_port);
   Ciphertext_regx164x : DFFRNQ_X1 port map( D => reg_out_164_port, CLK => clk,
                           RN => n656, Q => Ciphertext(164));
   Ciphertext_regx162x : DFFRNQ_X1 port map( D => reg_out_162_port, CLK => clk,
                           RN => n655, Q => Ciphertext(162));
   reg_in_regx29x : DFFSNQ_X1 port map( D => Plaintext(29), CLK => clk, SN => 
                           n654, Q => reg_in_29_port);
   reg_in_regx26x : DFFRNQ_X1 port map( D => Plaintext(26), CLK => clk, RN => 
                           n653, Q => reg_in_26_port);
   reg_key_regx151x : DFFRNQ_X1 port map( D => Key(151), CLK => clk, RN => n652
                           , Q => reg_key_151_port);
   Ciphertext_regx8x : DFFRNQ_X1 port map( D => reg_out_8_port, CLK => clk, RN 
                           => n651, Q => Ciphertext(8));
   Ciphertext_regx95x : DFFRNQ_X1 port map( D => reg_out_95_port, CLK => clk, 
                           RN => n650, Q => Ciphertext(95));
   Ciphertext_regx165x : DFFSNQ_X1 port map( D => reg_out_165_port, CLK => clk,
                           SN => n649, Q => Ciphertext(165));
   Ciphertext_regx169x : DFFRNQ_X1 port map( D => reg_out_169_port, CLK => clk,
                           RN => n648, Q => Ciphertext(169));
   Ciphertext_regx39x : DFFSNQ_X1 port map( D => reg_out_39_port, CLK => clk, 
                           SN => n647, Q => Ciphertext(39));
   reg_in_regx27x : DFFRNQ_X1 port map( D => Plaintext(27), CLK => clk, RN => 
                           n646, Q => reg_in_27_port);
   Ciphertext_regx57x : DFFRNQ_X1 port map( D => reg_out_57_port, CLK => clk, 
                           RN => n645, Q => Ciphertext(57));
   n645 <= '1';
   n646 <= '1';
   n647 <= '1';
   n648 <= '1';
   n649 <= '1';
   n650 <= '1';
   n651 <= '1';
   n652 <= '1';
   n653 <= '1';
   n654 <= '1';
   n655 <= '1';
   n656 <= '1';

end SYN_Behavioral;
