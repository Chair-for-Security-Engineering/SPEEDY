module SPEEDY_Rounds5_0 ( Ciphertext, Key, Plaintext );
  input [191:0] Ciphertext;
  input [191:0] Key;
  output [191:0] Plaintext;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n16, n17, n18,
         n19, n22, n23, n24, n25, n27, n28, n30, n31, n32, n35, n36, n38, n39,
         n40, n41, n42, n45, n46, n47, n48, n49, n50, n51, n52, n54, n55, n56,
         n57, n58, n60, n63, n64, n65, n67, n68, n69, n70, n71, n73, n74, n75,
         n76, n77, n82, n83, n86, n87, n89, n90, n91, n92, n93, n94, n95, n99,
         n100, n101, n102, n104, n106, n108, n110, n112, n113, n114, n115,
         n118, n119, n120, n121, n122, n125, n126, n127, n128, n129, n131,
         n132, n134, n135, n136, n137, n139, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n154, n155, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n169, n170, n171, n172,
         n173, n174, n175, n177, n180, n181, n183, n184, n185, n186, n188,
         n190, n191, n192, n193, n194, n195, n197, n198, n199, n200, n201,
         n204, n205, n206, n208, n209, n210, n211, n212, n216, n218, n219,
         n220, n222, n223, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n239, n240, n241, n242, n244, n245,
         n246, n247, n248, n250, n251, n252, n254, n255, n256, n257, n258,
         n259, n260, n261, n263, n264, n265, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n286, n287, n288, n289, n291, n293, n294, n295, n296, n297,
         n299, n300, n301, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n331, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n352, n353, n354, n355, n356, n357, n358, n362, n368, n369, n370,
         n372, n373, n374, n375, n376, n377, n381, n382, n383, n386, n388,
         n389, n390, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n405, n412, n413, n414, n417, n418, n419, n420, n423, n424, n426,
         n427, n430, n431, n432, n435, n438, n441, n442, n444, n445, n447,
         n452, n453, n454, n457, n458, n459, n460, n461, n462, n463, n467,
         n469, n471, n473, n480, n481, n483, n484, n485, n486, n487, n488,
         n489, n498, n505, n506, n507, n508, n509, n510, n511, n514, n515,
         n516, n517, n518, n522, n523, n525, n539, n540, n543, n544, n547,
         n548, n551, n555, n556, n557, n559, n560, n562, n563, n566, n567,
         n569, n574, n575, n576, n580, n581, n584, n585, n587, n588, n590,
         n591, n592, n593, n594, n596, n597, n598, n601, n602, n603, n604,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n742, n743,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n793, n794, n795, n796, n797, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n823, n824, n825,
         n826, n828, n829, n833, n834, n835, n836, n837, n838, n840, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n865,
         n866, n867, n868, n869, n870, n871, n872, n874, n875, n876, n877,
         n878, n879, n881, n882, n883, n884, n885, n886, n888, n889, n891,
         n892, n893, n894, n895, n896, n897, n899, n900, n901, n902, n903,
         n904, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n932, n933, n934, n935, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n966, n967, n968, n969, n970, n971, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1048,
         n1049, n1050, n1051, n1052, n1053, n1055, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1128, n1129, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1170, n1171, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1215, n1216, n1217, n1219, n1221, n1223, n1224,
         n1226, n1227, n1228, n1229, n1230, n1232, n1233, n1234, n1235, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1254, n1255, n1256, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1347,
         n1348, n1349, n1350, n1351, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1450, n1451, n1452,
         n1453, n1454, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1471, n1472, n1473, n1474,
         n1475, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1532, n1533, n1534, n1535, n1536, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1640, n1641, n1642, n1643, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1661, n1662, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1725, n1726, n1727, n1729, n1730, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1830, n1831, n1832, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1870, n1871,
         n1872, n1873, n1874, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1887, n1888, n1889, n1890, n1891, n1892, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2042, n2043, n2044, n2045, n2046, n2049, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2076, n2077, n2080, n2081, n2082, n2083, n2084, n2086, n2087, n2088,
         n2089, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2123, n2125, n2126, n2129, n2130, n2131, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2141, n2143, n2144, n2149, n2150,
         n2151, n2153, n2154, n2155, n2156, n2158, n2159, n2162, n2163, n2164,
         n2166, n2167, n2168, n2169, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2185, n2188, n2189, n2192, n2193,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2203, n2204, n2205,
         n2206, n2207, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2234, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2761, n2762, n2763, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2830, n2831, n2832, n2833, n2834, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2881, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2905, n2906, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2918, n2919, n2920, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3070, n3071, n3072, n3073, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3167, n3168, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3354,
         n3355, n3356, n3358, n3359, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3397,
         n3398, n3399, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3478, n3479, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3569, n3570, n3571, n3572, n3573, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3931, n3932, n3933, n3935,
         n3936, n3937, n3938, n3940, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3962, n3963, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4102, n4103, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4330, n4331, n4332, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4420, n4421, n4422, n4423, n4424, n4425, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4748, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4785, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4803, n4804, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4893,
         n4894, n4895, n4896, n4897, n4898, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4995, n4996, n4997, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5037, n5038, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5075,
         n5076, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5086, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5186, n5187, n5188, n5189, n5190, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5512, n5513, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5829, n5830, n5831, n5832, n5833,
         n5835, n5836, n5837, n5838, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5903, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6028, n6029, n6030, n6031, n6032, n6033, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6076,
         n6077, n6078, n6079, n6080, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6123, n6125, n6126, n6127, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6235, n6236, n6237, n6238, n6239, n6240, n6242, n6243, n6244, n6245,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6389,
         n6390, n6391, n6392, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6614, n6615, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6858, n6859, n6860, n6861, n6862, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6965, n6966, n6967, n6968, n6969, n6970, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7024,
         n7025, n7026, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7440, n7441, n7442, n7443, n7444, n7445, n7447, n7449, n7450, n7451,
         n7452, n7454, n7455, n7456, n7458, n7459, n7460, n7461, n7462, n7464,
         n7465, n7466, n7467, n7468, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7544, n7545, n7546, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7571, n7572,
         n7573, n7574, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7632, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8075, n8076, n8077, n8078, n8079, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8366, n8367, n8368, n8369, n8370, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8421, n8422, n8423,
         n8424, n8425, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8633, n8634, n8635, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9120, n9121, n9122,
         n9123, n9124, n9125, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10402, n10403, n10404, n10405, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10630, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11132, n11133, n11134, n11135, n11136, n11137, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11764, n11765, n11766,
         n11767, n11768, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11788, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14159, n14160, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16051,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17101, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18360, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19175, n19176, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19256, n19257, n19258, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20143, n20144, n20145, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20220, n20221, n20222, n20223, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20303, n20304, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20989, n20990, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21299, n21300, n21301, n21302, n21303, n21304,
         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
         n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
         n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,
         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
         n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
         n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360,
         n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,
         n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
         n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
         n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
         n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
         n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408,
         n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21687, n21688, n21689, n21690, n21691, n21692, n21693,
         n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701,
         n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
         n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717,
         n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
         n21726, n21727, n21728, n21729, n21730, n21731, n21733, n21734,
         n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742,
         n21743, n21744, n21746, n21748, n21749, n21750, n21751, n21752,
         n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
         n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768,
         n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
         n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
         n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792,
         n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800,
         n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
         n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
         n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
         n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840,
         n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
         n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
         n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864,
         n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872,
         n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
         n21881, n21882, n21883, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
         n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
         n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
         n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
         n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
         n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
         n21947, n21948, n21949, n21950, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
         n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
         n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
         n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22093,
         n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101,
         n22102, n22103, n22104, n22106, n22107, n22108, n22109, n22110,
         n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118,
         n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22127,
         n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
         n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
         n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,
         n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160,
         n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
         n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176,
         n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,
         n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192,
         n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,
         n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,
         n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
         n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224,
         n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,
         n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
         n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248,
         n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,
         n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
         n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
         n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280,
         n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
         n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296,
         n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304,
         n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,
         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
         n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
         n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
         n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
         n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
         n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368,
         n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
         n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
         n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,
         n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
         n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
         n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
         n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424,
         n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,
         n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440,
         n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448,
         n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,
         n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464,
         n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
         n22473, n22474, n22475, n22476, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22682, n22683, n22684,
         n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692,
         n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22701,
         n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709,
         n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717,
         n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725,
         n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733,
         n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741,
         n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749,
         n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757,
         n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765,
         n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773,
         n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781,
         n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789,
         n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22798,
         n22799, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
         n22808, n22810, n22811, n22812, n22813, n22814, n22815, n22816,
         n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,
         n22825, n22826, n22827, n22828, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22967, n22968, n22969, n22970,
         n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978,
         n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986,
         n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994,
         n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002,
         n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010,
         n23011, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23097, n23098, n23099, n23100,
         n23101, n23102, n23103, n23104, n23105, n23107, n23108, n23109,
         n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117,
         n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125,
         n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133,
         n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141,
         n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149,
         n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157,
         n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165,
         n23166, n23167, n23169, n23170, n23171, n23172, n23173, n23174,
         n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182,
         n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190,
         n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198,
         n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206,
         n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214,
         n23215, n23216, n23217, n23218, n23219, n23220, n23222, n23223,
         n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232,
         n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240,
         n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248,
         n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256,
         n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264,
         n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272,
         n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280,
         n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288,
         n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,
         n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304,
         n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312,
         n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320,
         n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328,
         n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336,
         n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344,
         n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352,
         n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360,
         n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368,
         n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376,
         n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384,
         n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392,
         n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400,
         n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408,
         n23409, n23410, n23411, n23412, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23520, n23521, n23522,
         n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530,
         n23531, n23533, n23535, n23536, n23537, n23538, n23539, n23540,
         n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548,
         n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556,
         n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564,
         n23565, n23566, n23568, n23569, n23570, n23571, n23572, n23573,
         n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581,
         n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589,
         n23590, n23591, n23592, n23593, n23594, n23595, n23597, n23598,
         n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606,
         n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614,
         n23615, n23616, n23617, n23618, n23619, n23621, n23622, n23623,
         n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631,
         n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639,
         n23640, n23641, n23642, n23643, n23644, n23645, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23710, n23711, n23712, n23713, n23714,
         n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722,
         n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730,
         n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738,
         n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746,
         n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754,
         n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762,
         n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770,
         n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778,
         n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786,
         n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794,
         n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802,
         n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810,
         n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818,
         n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826,
         n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834,
         n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842,
         n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850,
         n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858,
         n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866,
         n23867, n23868, n23869, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23975, n23976, n23977, n23978, n23979, n23980,
         n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988,
         n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996,
         n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004,
         n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012,
         n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020,
         n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028,
         n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036,
         n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044,
         n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052,
         n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060,
         n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068,
         n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076,
         n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084,
         n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092,
         n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100,
         n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108,
         n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116,
         n24117, n24118, n24119, n24120, n24121, n24123, n24124, n24126,
         n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134,
         n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142,
         n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150,
         n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158,
         n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166,
         n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174,
         n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182,
         n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190,
         n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198,
         n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206,
         n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214,
         n24215, n24216, n24217, n24218, n24220, n24221, n24222, n24223,
         n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231,
         n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239,
         n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247,
         n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255,
         n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263,
         n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271,
         n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279,
         n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287,
         n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295,
         n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303,
         n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311,
         n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319,
         n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327,
         n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
         n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343,
         n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351,
         n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359,
         n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367,
         n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375,
         n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383,
         n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391,
         n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399,
         n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
         n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415,
         n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423,
         n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431,
         n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439,
         n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447,
         n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455,
         n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463,
         n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471,
         n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479,
         n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487,
         n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496,
         n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504,
         n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512,
         n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520,
         n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528,
         n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536,
         n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544,
         n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552,
         n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560,
         n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568,
         n24569, n24570, n24571, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24878, n24879, n24880, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24990, n24991, n24992, n24993, n24994, n24995, n24996,
         n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004,
         n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012,
         n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020,
         n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028,
         n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036,
         n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044,
         n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052,
         n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060,
         n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068,
         n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076,
         n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084,
         n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093,
         n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101,
         n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109,
         n25110, n25111, n25113, n25114, n25115, n25116, n25117, n25118,
         n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126,
         n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134,
         n25135, n25136, n25137, n25138, n25139, n25141, n25142, n25143,
         n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151,
         n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159,
         n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167,
         n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175,
         n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183,
         n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191,
         n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199,
         n25200, n25201, n25202, n25203, n25204, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
         n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
         n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
         n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
         n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
         n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
         n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
         n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
         n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
         n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
         n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434,
         n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
         n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450,
         n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458,
         n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
         n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947,
         n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
         n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
         n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
         n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
         n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26021, n26023, n26024, n26025, n26026, n26027, n26028,
         n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036,
         n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044,
         n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26053,
         n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061,
         n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069,
         n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077,
         n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085,
         n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093,
         n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101,
         n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109,
         n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117,
         n26118, n26119, n26120, n26121, n26122, n26123, n26125, n26126,
         n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134,
         n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142,
         n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150,
         n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158,
         n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166,
         n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174,
         n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182,
         n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190,
         n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198,
         n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206,
         n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214,
         n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222,
         n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230,
         n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238,
         n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246,
         n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254,
         n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262,
         n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270,
         n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278,
         n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286,
         n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294,
         n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302,
         n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310,
         n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319,
         n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327,
         n26328, n26329, n26331, n26332, n26333, n26334, n26335, n26336,
         n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
         n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352,
         n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
         n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368,
         n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376,
         n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384,
         n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,
         n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400,
         n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408,
         n26409, n26410, n26411, n26412, n26413, n26414, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
         n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
         n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
         n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
         n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634,
         n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
         n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
         n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
         n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
         n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
         n26675, n26676, n26677, n26678, n26679, n26680, n26683, n26684,
         n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692,
         n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700,
         n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708,
         n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716,
         n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724,
         n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732,
         n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740,
         n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748,
         n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756,
         n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764,
         n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772,
         n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780,
         n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788,
         n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796,
         n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804,
         n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812,
         n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820,
         n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828,
         n26829, n26830, n26831, n26832, n26833, n26835, n26836, n26837,
         n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845,
         n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853,
         n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861,
         n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
         n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877,
         n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885,
         n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893,
         n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901,
         n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910,
         n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918,
         n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926,
         n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934,
         n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942,
         n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950,
         n26951, n26953, n26954, n26955, n26956, n26957, n26958, n26959,
         n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967,
         n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975,
         n26976, n26977, n26979, n26980, n26981, n26982, n26983, n26984,
         n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,
         n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000,
         n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,
         n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016,
         n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024,
         n27025, n27026, n27027, n27028, n27029, n27030, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27048, n27049, n27050,
         n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
         n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066,
         n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074,
         n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
         n27083, n27084, n27085, n27087, n27088, n27089, n27090, n27091,
         n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099,
         n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
         n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115,
         n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123,
         n27124, n27126, n27127, n27128, n27129, n27130, n27131, n27132,
         n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140,
         n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148,
         n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156,
         n27157, n27158, n27160, n27161, n27162, n27163, n27164, n27165,
         n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173,
         n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181,
         n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189,
         n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197,
         n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206,
         n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214,
         n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222,
         n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230,
         n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238,
         n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246,
         n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254,
         n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262,
         n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270,
         n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278,
         n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286,
         n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294,
         n27295, n27297, n27298, n27299, n27300, n27301, n27302, n27303,
         n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311,
         n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319,
         n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327,
         n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335,
         n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343,
         n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351,
         n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359,
         n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367,
         n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375,
         n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383,
         n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391,
         n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399,
         n27400, n27401, n27403, n27404, n27405, n27406, n27407, n27408,
         n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416,
         n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424,
         n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432,
         n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440,
         n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448,
         n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456,
         n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,
         n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472,
         n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480,
         n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27530,
         n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
         n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
         n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554,
         n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
         n27563, n27564, n27566, n27567, n27568, n27569, n27570, n27571,
         n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579,
         n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587,
         n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
         n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603,
         n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611,
         n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619,
         n27620, n27621, n27623, n27624, n27625, n27626, n27627, n27628,
         n27629, n27631, n27632, n27633, n27634, n27635, n27636, n27637,
         n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645,
         n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653,
         n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661,
         n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669,
         n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677,
         n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685,
         n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693,
         n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701,
         n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709,
         n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717,
         n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725,
         n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733,
         n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741,
         n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749,
         n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757,
         n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765,
         n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773,
         n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781,
         n27782, n27783, n27784, n27786, n27787, n27788, n27789, n27790,
         n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798,
         n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806,
         n27807, n27808, n27809, n27810, n27811, n27812, n27814, n27815,
         n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823,
         n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831,
         n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839,
         n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847,
         n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855,
         n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863,
         n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871,
         n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879,
         n27880, n27881, n27882, n27883, n27885, n27886, n27887, n27888,
         n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896,
         n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904,
         n27905, n27906, n27907, n27908, n27909, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27961, n27962,
         n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970,
         n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978,
         n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986,
         n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994,
         n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002,
         n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010,
         n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018,
         n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026,
         n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034,
         n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042,
         n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050,
         n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058,
         n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066,
         n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074,
         n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082,
         n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090,
         n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
         n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
         n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114,
         n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122,
         n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130,
         n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138,
         n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146,
         n28147, n28148, n28149, n28150, n28152, n28153, n28155, n28156,
         n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164,
         n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172,
         n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180,
         n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188,
         n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196,
         n28197, n28198, n28200, n28201, n28202, n28203, n28204, n28205,
         n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213,
         n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221,
         n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229,
         n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237,
         n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245,
         n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253,
         n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261,
         n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269,
         n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277,
         n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285,
         n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293,
         n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301,
         n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309,
         n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317,
         n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325,
         n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333,
         n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341,
         n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349,
         n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357,
         n28358, n28359, n28360, n28361, n28362, n28364, n28365, n28366,
         n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374,
         n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382,
         n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390,
         n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398,
         n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406,
         n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414,
         n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422,
         n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430,
         n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
         n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446,
         n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454,
         n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462,
         n28463, n28464, n28465, n28466, n28469, n28470, n28471, n28472,
         n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480,
         n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530,
         n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538,
         n28539, n28540, n28541, n28543, n28544, n28545, n28546, n28547,
         n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
         n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564,
         n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572,
         n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581,
         n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589,
         n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597,
         n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605,
         n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613,
         n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621,
         n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629,
         n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637,
         n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645,
         n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28654,
         n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662,
         n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670,
         n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678,
         n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686,
         n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694,
         n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702,
         n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710,
         n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718,
         n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726,
         n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734,
         n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742,
         n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750,
         n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758,
         n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766,
         n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774,
         n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782,
         n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790,
         n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798,
         n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806,
         n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814,
         n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822,
         n28823, n28824, n28825, n28826, n28827, n28828, n28830, n28831,
         n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839,
         n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847,
         n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855,
         n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863,
         n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871,
         n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879,
         n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887,
         n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895,
         n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903,
         n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911,
         n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919,
         n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927,
         n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935,
         n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943,
         n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951,
         n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959,
         n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967,
         n28968, n28970, n28971, n28972, n28973, n28974, n28975, n28976,
         n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984,
         n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992,
         n28993, n28994, n28995, n28996, n28997, n28998, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29025, n29026,
         n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034,
         n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042,
         n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050,
         n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058,
         n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066,
         n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074,
         n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082,
         n29083, n29084, n29085, n29086, n29087, n29089, n29090, n29091,
         n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099,
         n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
         n29108, n29110, n29111, n29112, n29114, n29115, n29116, n29117,
         n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125,
         n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133,
         n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141,
         n29142, n29143, n29145, n29146, n29147, n29148, n29149, n29150,
         n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158,
         n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166,
         n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174,
         n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182,
         n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190,
         n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198,
         n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206,
         n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214,
         n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222,
         n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230,
         n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238,
         n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246,
         n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254,
         n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262,
         n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270,
         n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278,
         n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286,
         n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294,
         n29295, n29296, n29298, n29299, n29300, n29301, n29302, n29303,
         n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311,
         n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319,
         n29320, n29321, n29323, n29324, n29325, n29326, n29327, n29328,
         n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336,
         n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344,
         n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352,
         n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360,
         n29361, n29362, n29363, n29364, n29365, n29366, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
         n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394,
         n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402,
         n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410,
         n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418,
         n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426,
         n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435,
         n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443,
         n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451,
         n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459,
         n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
         n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475,
         n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483,
         n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491,
         n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499,
         n29500, n29501, n29502, n29504, n29505, n29506, n29507, n29508,
         n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516,
         n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524,
         n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532,
         n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540,
         n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548,
         n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556,
         n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564,
         n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572,
         n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580,
         n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588,
         n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596,
         n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604,
         n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612,
         n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620,
         n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628,
         n29629, n29630, n29631, n29632, n29634, n29635, n29636, n29637,
         n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645,
         n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653,
         n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661,
         n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669,
         n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677,
         n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685,
         n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693,
         n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701,
         n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709,
         n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717,
         n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725,
         n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733,
         n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741,
         n29742, n29743, n29745, n29746, n29747, n29748, n29749, n29750,
         n29751, n29753, n29754, n29755, n29756, n29757, n29758, n29759,
         n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767,
         n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775,
         n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783,
         n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791,
         n29792, n29794, n29795, n29796, n29797, n29798, n29799, n29800,
         n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808,
         n29809, n29810, n29811, n29812, n29813, n29814, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30080, n30081, n30082,
         n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090,
         n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098,
         n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106,
         n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114,
         n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122,
         n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130,
         n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138,
         n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146,
         n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154,
         n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162,
         n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170,
         n30171, n30172, n30173, n30174, n30175, n30177, n30178, n30179,
         n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
         n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195,
         n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203,
         n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211,
         n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219,
         n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
         n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235,
         n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243,
         n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251,
         n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
         n30260, n30261, n30262, n30263, n30265, n30266, n30267, n30268,
         n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276,
         n30279, n30280, n30281, n30282, n30283, n30285, n30286, n30287,
         n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295,
         n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303,
         n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311,
         n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319,
         n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327,
         n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335,
         n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343,
         n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351,
         n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359,
         n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367,
         n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375,
         n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383,
         n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391,
         n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399,
         n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407,
         n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415,
         n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423,
         n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431,
         n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439,
         n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447,
         n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455,
         n30456, n30458, n30459, n30460, n30461, n30462, n30463, n30464,
         n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30615, n30616, n30617, n30618,
         n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626,
         n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634,
         n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642,
         n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650,
         n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658,
         n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666,
         n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674,
         n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682,
         n30683, n30684, n30685, n30686, n30687, n30688, n30690, n30691,
         n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699,
         n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707,
         n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715,
         n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723,
         n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731,
         n30732, n30733, n30734, n30735, n30736, n30737, n30740, n30741,
         n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749,
         n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757,
         n30758, n30759, n30760, n30761, n30762, n30763, n30764, n30765,
         n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773,
         n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781,
         n30782, n30783, n30784, n30785, n30787, n30788, n30789, n30790,
         n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798,
         n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806,
         n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814,
         n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822,
         n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830,
         n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838,
         n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846,
         n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854,
         n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862,
         n30863, n30864, n30865, n30866, n30868, n30869, n30870, n30872,
         n30873, n30876, n30877, n30878, n30879, n30880, n30881, n30882,
         n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890,
         n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898,
         n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906,
         n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914,
         n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922,
         n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930,
         n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938,
         n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947,
         n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955,
         n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963,
         n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30972,
         n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980,
         n30981, n30982, n30983, n30985, n30986, n30987, n30988, n30989,
         n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997,
         n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005,
         n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013,
         n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021,
         n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029,
         n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037,
         n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045,
         n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053,
         n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061,
         n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069,
         n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078,
         n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086,
         n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094,
         n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102,
         n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110,
         n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118,
         n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126,
         n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134,
         n31135, n31136, n31137, n31139, n31140, n31141, n31142, n31143,
         n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151,
         n31152, n31153, n31155, n31156, n31157, n31158, n31159, n31160,
         n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168,
         n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176,
         n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184,
         n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192,
         n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200,
         n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208,
         n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216,
         n31217, n31218, n31219, n31220, n31221, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31271, n31272, n31273, n31274,
         n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282,
         n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290,
         n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298,
         n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306,
         n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314,
         n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322,
         n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330,
         n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338,
         n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346,
         n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354,
         n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362,
         n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370,
         n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378,
         n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31387,
         n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31396,
         n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404,
         n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412,
         n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420,
         n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428,
         n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436,
         n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444,
         n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452,
         n31453, n31454, n31455, n31456, n31457, n31460, n31461, n31462,
         n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470,
         n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478,
         n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486,
         n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494,
         n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502,
         n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510,
         n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518,
         n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526,
         n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534,
         n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542,
         n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550,
         n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558,
         n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566,
         n31567, n31568, n31569, n31571, n31572, n31573, n31574, n31575,
         n31576, n31577, n31578, n31580, n31581, n31582, n31583, n31584,
         n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592,
         n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600,
         n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608,
         n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616,
         n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624,
         n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632,
         n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640,
         n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648,
         n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656,
         n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664,
         n31665, n31666, n31667, n31668, n31669, n31670, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31775, n31776, n31777, n31778,
         n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786,
         n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794,
         n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802,
         n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810,
         n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818,
         n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826,
         n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834,
         n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842,
         n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850,
         n31851, n31852, n31853, n31855, n31856, n31857, n31858, n31859,
         n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867,
         n31868, n31870, n31872, n31873, n31874, n31875, n31876, n31877,
         n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885,
         n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893,
         n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901,
         n31902, n31904, n31906, n31907, n31908, n31909, n31910, n31911,
         n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919,
         n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927,
         n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935,
         n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943,
         n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951,
         n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959,
         n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967,
         n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975,
         n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983,
         n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991,
         n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999,
         n32000, n32001, n32002, n32003, n32004, n32006, n32007, n32008,
         n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016,
         n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024,
         n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032,
         n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32065, n32066,
         n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074,
         n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082,
         n32083, n32084, n32086, n32087, n32088, n32089, n32090, n32091,
         n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099,
         n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107,
         n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115,
         n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123,
         n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131,
         n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139,
         n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147,
         n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155,
         n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163,
         n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171,
         n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32180,
         n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188,
         n32189, n32190, n32191, n32193, n32194, n32195, n32196, n32197,
         n32198, n32199, n32200, n32201, n32202, n32203, n32204, n32205,
         n32206, n32207, n32208, n32209, n32210, n32211, n32212, n32213,
         n32214, n32215, n32216, n32217, n32219, n32220, n32221, n32222,
         n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230,
         n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238,
         n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246,
         n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254,
         n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262,
         n32263, n32264, n32265, n32267, n32268, n32269, n32270, n32271,
         n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279,
         n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287,
         n32288, n32289, n32290, n32291, n32292, n32293, n32294, n32295,
         n32296, n32297, n32298, n32299, n32300, n32301, n32302, n32303,
         n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311,
         n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319,
         n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327,
         n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335,
         n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343,
         n32344, n32345, n32346, n32347, n32348, n32349, n32350, n32351,
         n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359,
         n32360, n32361, n32362, n32363, n32364, n32365, n32366, n32367,
         n32368, n32369, n32370, n32371, n32372, n32373, n32374, n32375,
         n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383,
         n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391,
         n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399,
         n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407,
         n32408, n32409, n32410, n32411, n32412, n32413, n32414, n32415,
         n32416, n32417, n32418, n32419, n32420, n32421, n32422, n32423,
         n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431,
         n32432, n32433, n32434, n32436, n32437, n32438, n32439, n32440,
         n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448,
         n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456,
         n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464,
         n32465, n32466, n32469, n32470, n32471, n32472, n32473, n32474,
         n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482,
         n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490,
         n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498,
         n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506,
         n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514,
         n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522,
         n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530,
         n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32540,
         n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548,
         n32549, n32550, n32551, n32552, n32553, n32554, n32555, n32556,
         n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564,
         n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572,
         n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580,
         n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588,
         n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596,
         n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604,
         n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612,
         n32613, n32614, n32615, n32616, n32617, n32618, n32620, n32621,
         n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629,
         n32630, n32631, n32632, n32633, n32634, n32635, n32636, n32637,
         n32638, n32639, n32640, n32641, n32642, n32643, n32644, n32645,
         n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653,
         n32654, n32655, n32656, n32657, n32658, n32659, n32660, n32661,
         n32662, n32663, n32664, n32665, n32666, n32667, n32668, n32669,
         n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677,
         n32678, n32679, n32680, n32681, n32682, n32683, n32684, n32685,
         n32686, n32687, n32688, n32689, n32690, n32691, n32692, n32693,
         n32694, n32695, n32696, n32697, n32698, n32699, n32700, n32701,
         n32702, n32703, n32704, n32705, n32706, n32707, n32708, n32709,
         n32710, n32711, n32712, n32713, n32714, n32715, n32716, n32717,
         n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725,
         n32726, n32727, n32728, n32729, n32730, n32731, n32732, n32733,
         n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741,
         n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749,
         n32750, n32751, n32752, n32753, n32754, n32755, n32756, n32757,
         n32758, n32759, n32760, n32761, n32762, n32763, n32764, n32765,
         n32766, n32767, n32768, n32769, n32770, n32771, n32772, n32773,
         n32774, n32775, n32776, n32777, n32778, n32779, n32780, n32781,
         n32782, n32783, n32784, n32785, n32786, n32787, n32788, n32789,
         n32790, n32791, n32792, n32793, n32794, n32795, n32796, n32797,
         n32798, n32799, n32800, n32801, n32802, n32803, n32804, n32805,
         n32806, n32807, n32808, n32809, n32810, n32811, n32812, n32813,
         n32814, n32815, n32816, n32817, n32818, n32819, n32820, n32821,
         n32822, n32823, n32824, n32825, n32826, n32827, n32828, n32829,
         n32830, n32831, n32832, n32833, n32834, n32835, n32836, n32837,
         n32838, n32839, n32840, n32841, n32842, n32843, n32844, n32845,
         n32846, n32847, n32848, n32849, n32850, n32851, n32852, n32853,
         n32854, n32855, n32856, n32857, n32858, n32859, n32860, n32861,
         n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869,
         n32870, n32871, n32873, n32874, n32875, n32876, n32877, n32878,
         n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886,
         n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894,
         n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902,
         n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910,
         n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918,
         n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926,
         n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934,
         n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942,
         n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950,
         n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958,
         n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966,
         n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974,
         n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982,
         n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990,
         n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999,
         n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007,
         n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015,
         n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023,
         n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031,
         n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039,
         n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047,
         n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055,
         n33056, n33057, n33058, n33059, n33060, n33061, n33062, n33063,
         n33064, n33065, n33066, n33067, n33068, n33070, n33071, n33072,
         n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080,
         n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088,
         n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096,
         n33097, n33098, n33099, n33100, n33101, n33102, n33103, n33104,
         n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112,
         n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120,
         n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128,
         n33129, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33154,
         n33155, n33157, n33158, n33159, n33160, n33162, n33163, n33164,
         n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172,
         n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180,
         n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188,
         n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196,
         n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204,
         n33205, n33206, n33207, n33208, n33209, n33210, n33211, n33212,
         n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220,
         n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228,
         n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236,
         n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244,
         n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252,
         n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260,
         n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268,
         n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276,
         n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284,
         n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292,
         n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300,
         n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308,
         n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316,
         n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324,
         n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332,
         n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340,
         n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348,
         n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356,
         n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364,
         n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372,
         n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380,
         n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388,
         n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396,
         n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404,
         n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412,
         n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420,
         n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428,
         n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33437,
         n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445,
         n33446, n33447, n33448, n33449, n33450, n33451, n33452, n33453,
         n33454, n33455, n33456, n33457, n33458, n33459, n33460, n33461,
         n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469,
         n33470, n33471, n33472, n33473, n33474, n33475, n33476, n33477,
         n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485,
         n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493,
         n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501,
         n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509,
         n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517,
         n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525,
         n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533,
         n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541,
         n33542, n33543, n33544, n33545, n33546, n33547, n33548, n33549,
         n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557,
         n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565,
         n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573,
         n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581,
         n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589,
         n33590, n33591, n33592, n33593, n33594, n33595, n33596, n33597,
         n33598, n33599, n33600, n33601, n33602, n33603, n33604, n33605,
         n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613,
         n33614, n33615, n33616, n33617, n33618, n33619, n33620, n33621,
         n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629,
         n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637,
         n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645,
         n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33653,
         n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661,
         n33662, n33663, n33664, n33666, n33667, n33668, n33669, n33670,
         n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678,
         n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
         n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694,
         n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702,
         n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710,
         n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718,
         n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726,
         n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734,
         n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
         n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750,
         n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758,
         n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766,
         n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774,
         n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782,
         n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790,
         n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798,
         n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806,
         n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814,
         n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822,
         n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830,
         n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838,
         n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846,
         n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
         n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862,
         n33863, n33864, n33865, n33866, n33867, n33868, n33870, n33871,
         n33872, n33873, n33874, n33875, n33876, n33877, n33878, n33879,
         n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887,
         n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895,
         n33896, n33897, n33898, n33899, n33900, n33901, n33902, n33903,
         n33904, n33905, n33906, n33907, n33908, n33909, n33910, n33911,
         n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919,
         n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927,
         n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935,
         n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943,
         n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951,
         n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959,
         n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967,
         n33968, n33969, n33970, n33971, n33973, n33974, n33975, n33976,
         n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984,
         n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992,
         n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000,
         n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008,
         n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016,
         n34017, n34018, n34019, n34020, n34021, n34022, n34025, n34026,
         n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034,
         n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042,
         n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050,
         n34051, n34052, n34053, n34054, n34055, n34056, n34057, n34058,
         n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066,
         n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074,
         n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082,
         n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090,
         n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098,
         n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106,
         n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114,
         n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122,
         n34123, n34124, n34125, n34126, n34127, n34128, n34129, n34130,
         n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138,
         n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146,
         n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154,
         n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162,
         n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170,
         n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178,
         n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186,
         n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194,
         n34195, n34196, n34197, n34198, n34199, n34200, n34201, n34202,
         n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210,
         n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218,
         n34219, n34220, n34221, n34222, n34224, n34225, n34226, n34227,
         n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235,
         n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243,
         n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251,
         n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259,
         n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267,
         n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275,
         n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283,
         n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291,
         n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299,
         n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307,
         n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315,
         n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323,
         n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331,
         n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339,
         n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347,
         n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34356,
         n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364,
         n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372,
         n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380,
         n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388,
         n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396,
         n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404,
         n34405, n34406, n34407, n34409, n34410, n34411, n34412, n34413,
         n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421,
         n34422, n34423, n34424, n34425, n34426, n34427, n34428, n34429,
         n34430, n34431, n34432, n34433, n34434, n34435, n34436, n34437,
         n34438, n34439, n34440, n34441, n34442, n34443, n34444, n34445,
         n34446, n34447, n34448, n34449, n34450, n34451, n34452, n34453,
         n34454, n34455, n34456, n34457, n34458, n34460, n34461, n34462,
         n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470,
         n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478,
         n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486,
         n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494,
         n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502,
         n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510,
         n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518,
         n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526,
         n34527, n34528, n34529, n34530, n34531, n34533, n34534, n34535,
         n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543,
         n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551,
         n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559,
         n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567,
         n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575,
         n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583,
         n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591,
         n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599,
         n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607,
         n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615,
         n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623,
         n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631,
         n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639,
         n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647,
         n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655,
         n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663,
         n34664, n34665, n34666, n34667, n34668, n34669, n34670, n34671,
         n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679,
         n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687,
         n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695,
         n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703,
         n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711,
         n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719,
         n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727,
         n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735,
         n34736, n34737, n34739, n34740, n34741, n34742, n34743, n34744,
         n34745, n34746, n34747, n34748, n34749, n34750, n34751, n34752,
         n34753, n34754, n34755, n34756, n34757, n34758, n34759, n34760,
         n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768,
         n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776,
         n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784,
         n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792,
         n34793, n34794, n34795, n34796, n34797, n34798, n34799, n34800,
         n34801, n34802, n34803, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34823, n34824, n34825, n34826,
         n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834,
         n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842,
         n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850,
         n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858,
         n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866,
         n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874,
         n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882,
         n34883, n34884, n34885, n34886, n34887, n34888, n34889, n34890,
         n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898,
         n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906,
         n34907, n34908, n34909, n34910, n34911, n34912, n34913, n34914,
         n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922,
         n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930,
         n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938,
         n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946,
         n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954,
         n34955, n34956, n34957, n34958, n34959, n34960, n34961, n34962,
         n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970,
         n34971, n34972, n34973, n34974, n34976, n34977, n34978, n34979,
         n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987,
         n34989, n34991, n34992, n34993, n34994, n34995, n34996, n34997,
         n34998, n34999, n35000, n35001, n35002, n35003, n35004, n35005,
         n35006, n35007, n35008, n35009, n35010, n35011, n35012, n35013,
         n35014, n35015, n35016, n35017, n35018, n35019, n35020, n35021,
         n35022, n35023, n35024, n35025, n35026, n35027, n35028, n35029,
         n35030, n35031, n35032, n35033, n35034, n35035, n35036, n35037,
         n35038, n35039, n35040, n35041, n35042, n35043, n35044, n35045,
         n35046, n35047, n35048, n35049, n35050, n35051, n35052, n35054,
         n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062,
         n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070,
         n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078,
         n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086,
         n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094,
         n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102,
         n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110,
         n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118,
         n35119, n35120, n35121, n35122, n35124, n35125, n35126, n35127,
         n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135,
         n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143,
         n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151,
         n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159,
         n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167,
         n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175,
         n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35184,
         n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192,
         n35193, n35194, n35195, n35196, n35197, n35199, n35200, n35201,
         n35202, n35203, n35204, n35206, n35207, n35208, n35209, n35210,
         n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218,
         n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226,
         n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234,
         n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242,
         n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250,
         n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258,
         n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266,
         n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274,
         n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282,
         n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290,
         n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298,
         n35299, n35300, n35301, n35302, n35304, n35305, n35306, n35307,
         n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315,
         n35316, n35317, n35318, n35320, n35321, n35322, n35323, n35324,
         n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332,
         n35333, n35334, n35335, n35336, n35337, n35338, n35339, n35340,
         n35341, n35342, n35343, n35344, n35345, n35346, n35347, n35348,
         n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356,
         n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35364,
         n35365, n35366, n35367, n35368, n35369, n35370, n35371, n35372,
         n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380,
         n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388,
         n35389, n35390, n35391, n35392, n35393, n35394, n35395, n35396,
         n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404,
         n35405, n35406, n35407, n35408, n35409, n35410, n35411, n35412,
         n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420,
         n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428,
         n35429, n35430, n35431, n35432, n35433, n35434, n35436, n35437,
         n35438, n35439, n35440, n35441, n35443, n35444, n35445, n35446,
         n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456,
         n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464,
         n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472,
         n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480,
         n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488,
         n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496,
         n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504,
         n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514,
         n35515, n35517, n35518, n35519, n35520, n35521, n35522, n35523,
         n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531,
         n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539,
         n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547,
         n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555,
         n35556, n35557, n35559, n35560, n35561, n35562, n35564, n35565,
         n35566, n35567, n35568, n35569, n35570, n35571, n35572, n35573,
         n35574, n35575, n35576, n35577, n35578, n35579, n35580, n35581,
         n35582, n35583, n35584, n35585, n35586, n35587, n35588, n35589,
         n35590, n35591, n35592, n35593, n35594, n35595, n35596, n35597,
         n35598, n35599, n35600, n35601, n35602, n35603, n35604, n35605,
         n35606, n35607, n35608, n35609, n35610, n35611, n35612, n35613,
         n35614, n35615, n35616, n35617, n35618, n35619, n35620, n35621,
         n35622, n35623, n35624, n35625, n35626, n35627, n35628, n35629,
         n35630, n35631, n35632, n35633, n35634, n35635, n35636, n35637,
         n35638, n35639, n35640, n35641, n35642, n35643, n35644, n35645,
         n35646, n35647, n35648, n35649, n35650, n35651, n35652, n35653,
         n35654, n35655, n35656, n35657, n35658, n35659, n35660, n35661,
         n35662, n35663, n35664, n35665, n35666, n35667, n35668, n35669,
         n35670, n35671, n35672, n35673, n35674, n35675, n35676, n35677,
         n35678, n35679, n35680, n35681, n35682, n35683, n35684, n35685,
         n35686, n35687, n35688, n35689, n35690, n35691, n35692, n35693,
         n35694, n35695, n35696, n35697, n35698, n35699, n35700, n35701,
         n35702, n35703, n35704, n35705, n35706, n35707, n35708, n35709,
         n35710, n35711, n35712, n35713, n35714, n35715, n35716, n35717,
         n35718, n35719, n35720, n35721, n35722, n35723, n35724, n35725,
         n35726, n35727, n35728, n35729, n35730, n35731, n35732, n35733,
         n35734, n35735, n35736, n35738, n35739, n35740, n35741, n35742,
         n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750,
         n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759,
         n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767,
         n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775,
         n35777, n35778, n35779, n35780, n35781, n35782, n35783, n35784,
         n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792,
         n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800,
         n35801, n35802, n35803, n35804, n35805, n35806, n35807, n35808,
         n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816,
         n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824,
         n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832,
         n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840,
         n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848,
         n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856,
         n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864,
         n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35888, n35889, n35890,
         n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898,
         n35899, n35900, n35901, n35902, n35903, n35905, n35906, n35907,
         n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915,
         n35916, n35917, n35918, n35920, n35921, n35922, n35923, n35924,
         n35925, n35927, n35928, n35929, n35930, n35931, n35932, n35933,
         n35934, n35935, n35936, n35937, n35938, n35939, n35940, n35941,
         n35942, n35943, n35944, n35945, n35946, n35947, n35948, n35949,
         n35950, n35951, n35952, n35953, n35954, n35955, n35956, n35957,
         n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965,
         n35966, n35967, n35968, n35969, n35970, n35971, n35972, n35973,
         n35974, n35975, n35976, n35977, n35978, n35979, n35980, n35981,
         n35982, n35983, n35984, n35985, n35986, n35988, n35989, n35990,
         n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998,
         n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006,
         n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014,
         n36015, n36016, n36017, n36018, n36019, n36021, n36022, n36023,
         n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031,
         n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039,
         n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047,
         n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055,
         n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063,
         n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071,
         n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079,
         n36080, n36081, n36082, n36084, n36085, n36086, n36087, n36088,
         n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096,
         n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104,
         n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112,
         n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120,
         n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128,
         n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136,
         n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144,
         n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152,
         n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160,
         n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168,
         n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176,
         n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184,
         n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192,
         n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200,
         n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208,
         n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216,
         n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224,
         n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232,
         n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240,
         n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248,
         n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256,
         n36257, n36259, n36260, n36261, n36262, n36263, n36265, n36266,
         n36267, n36268, n36269, n36270, n36271, n36272, n36274, n36275,
         n36277, n36278, n36279, n36280, n36281, n36282, n36283, n36284,
         n36285, n36286, n36287, n36289, n36290, n36291, n36292, n36293,
         n36294, n36295, n36296, n36297, n36298, n36299, n36300, n36301,
         n36302, n36303, n36304, n36305, n36306, n36307, n36308, n36309,
         n36310, n36311, n36312, n36313, n36314, n36315, n36316, n36317,
         n36318, n36319, n36320, n36321, n36322, n36323, n36324, n36325,
         n36326, n36327, n36328, n36329, n36330, n36331, n36332, n36333,
         n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36341,
         n36342, n36343, n36344, n36345, n36346, n36347, n36348, n36349,
         n36350, n36351, n36352, n36353, n36354, n36355, n36356, n36357,
         n36358, n36359, n36360, n36361, n36362, n36363, n36364, n36365,
         n36366, n36367, n36368, n36369, n36370, n36371, n36372, n36373,
         n36374, n36375, n36376, n36377, n36378, n36379, n36380, n36381,
         n36382, n36383, n36384, n36385, n36386, n36387, n36388, n36389,
         n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397,
         n36398, n36399, n36400, n36401, n36402, n36403, n36404, n36405,
         n36406, n36407, n36408, n36409, n36410, n36411, n36412, n36413,
         n36414, n36415, n36416, n36417, n36418, n36419, n36420, n36421,
         n36422, n36423, n36424, n36425, n36426, n36427, n36428, n36429,
         n36430, n36431, n36432, n36433, n36434, n36435, n36436, n36437,
         n36438, n36439, n36440, n36441, n36442, n36443, n36444, n36445,
         n36446, n36447, n36448, n36449, n36450, n36451, n36453, n36454,
         n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462,
         n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470,
         n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478,
         n36479, n36480, n36481, n36482, n36483, n36484, n36486, n36487,
         n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495,
         n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503,
         n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511,
         n36512, n36513, n36514, n36515, n36516, n36517, n36518, n36519,
         n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527,
         n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535,
         n36536, n36537, n36538, n36539, n36540, n36541, n36542, n36543,
         n36544, n36545, n36546, n36547, n36548, n36549, n36550, n36551,
         n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559,
         n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567,
         n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575,
         n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583,
         n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591,
         n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599,
         n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607,
         n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615,
         n36616, n36617, n36618, n36619, n36620, n36621, n36622, n36623,
         n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631,
         n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639,
         n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647,
         n36648, n36649, n36650, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36703, n36704, n36705, n36706,
         n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714,
         n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722,
         n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730,
         n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738,
         n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746,
         n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754,
         n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762,
         n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770,
         n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778,
         n36779, n36780, n36781, n36782, n36783, n36784, n36786, n36787,
         n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795,
         n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803,
         n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811,
         n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819,
         n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828,
         n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36836,
         n36837, n36838, n36839, n36840, n36841, n36842, n36843, n36844,
         n36845, n36846, n36847, n36849, n36850, n36851, n36852, n36853,
         n36854, n36855, n36856, n36857, n36858, n36859, n36860, n36861,
         n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869,
         n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877,
         n36878, n36879, n36880, n36881, n36882, n36883, n36884, n36885,
         n36886, n36887, n36888, n36889, n36890, n36891, n36892, n36893,
         n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901,
         n36902, n36903, n36904, n36905, n36906, n36907, n36908, n36909,
         n36910, n36911, n36912, n36913, n36914, n36915, n36916, n36917,
         n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925,
         n36926, n36927, n36928, n36929, n36930, n36931, n36932, n36933,
         n36934, n36935, n36936, n36937, n36938, n36939, n36940, n36941,
         n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949,
         n36950, n36951, n36952, n36953, n36954, n36955, n36956, n36957,
         n36958, n36959, n36960, n36961, n36962, n36963, n36964, n36965,
         n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973,
         n36974, n36975, n36976, n36977, n36978, n36979, n36980, n36981,
         n36982, n36983, n36984, n36985, n36986, n36987, n36988, n36989,
         n36990, n36991, n36992, n36993, n36994, n36995, n36996, n36997,
         n36998, n36999, n37000, n37001, n37002, n37003, n37004, n37005,
         n37006, n37007, n37008, n37009, n37010, n37011, n37012, n37013,
         n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021,
         n37022, n37023, n37024, n37025, n37026, n37027, n37028, n37029,
         n37030, n37031, n37032, n37033, n37034, n37035, n37036, n37037,
         n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045,
         n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053,
         n37054, n37055, n37056, n37057, n37058, n37059, n37060, n37061,
         n37062, n37063, n37064, n37065, n37066, n37067, n37068, n37069,
         n37070, n37071, n37072, n37073, n37074, n37075, n37076, n37077,
         n37078, n37079, n37080, n37081, n37082, n37083, n37084, n37085,
         n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093,
         n37094, n37095, n37096, n37097, n37098, n37099, n37100, n37101,
         n37102, n37103, n37104, n37105, n37106, n37107, n37108, n37109,
         n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117,
         n37118, n37119, n37120, n37121, n37122, n37123, n37124, n37125,
         n37126, n37127, n37128, n37129, n37130, n37131, n37132, n37133,
         n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141,
         n37142, n37143, n37144, n37145, n37146, n37147, n37148, n37149,
         n37150, n37151, n37152, n37153, n37154, n37155, n37156, n37157,
         n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165,
         n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173,
         n37174, n37175, n37176, n37177, n37178, n37179, n37180, n37181,
         n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189,
         n37190, n37191, n37192, n37193, n37194, n37195, n37196, n37197,
         n37198, n37199, n37200, n37201, n37202, n37203, n37204, n37205,
         n37206, n37207, n37208, n37209, n37210, n37211, n37212, n37213,
         n37214, n37215, n37216, n37217, n37219, n37220, n37221, n37222,
         n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230,
         n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238,
         n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246,
         n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254,
         n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262,
         n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270,
         n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278,
         n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287,
         n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295,
         n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303,
         n37304, n37305, n37306, n37307, n37308, n37309, n37310, n37311,
         n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319,
         n37320, n37321, n37323, n37324, n37325, n37326, n37327, n37328,
         n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336,
         n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344,
         n37345, n37346, n37347, n37348, n37349, n37350, n37351, n37352,
         n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360,
         n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368,
         n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376,
         n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384,
         n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392,
         n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400,
         n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408,
         n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416,
         n37417, n37418, n37419, n37420, n37421, n37422, n37423, n37424,
         n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432,
         n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440,
         n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448,
         n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456,
         n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464,
         n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472,
         n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480,
         n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488,
         n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496,
         n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504,
         n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512,
         n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520,
         n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528,
         n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536,
         n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544,
         n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552,
         n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560,
         n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568,
         n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576,
         n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584,
         n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592,
         n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600,
         n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608,
         n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616,
         n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624,
         n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632,
         n37633, n37634, n37635, n37636, n37637, n37638, n37639, n37640,
         n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648,
         n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656,
         n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664,
         n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672,
         n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680,
         n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688,
         n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696,
         n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37744, n37745, n37746,
         n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754,
         n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762,
         n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770,
         n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778,
         n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786,
         n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794,
         n37795, n37796, n37797, n37798, n37799, n37800, n37801, n37802,
         n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810,
         n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818,
         n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826,
         n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834,
         n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843,
         n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851,
         n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859,
         n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867,
         n37868, n37869, n37870, n37871, n37872, n37873, n37875, n37876,
         n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885,
         n37886, n37887, n37888, n37890, n37891, n37892, n37893, n37894,
         n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902,
         n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910,
         n37911, n37912, n37913, n37914, n37916, n37917, n37918, n37919,
         n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927,
         n37928, n37929, n37930, n37931, n37932, n37933, n37934, n37935,
         n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943,
         n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951,
         n37952, n37953, n37954, n37955, n37956, n37957, n37958, n37959,
         n37960, n37961, n37962, n37963, n37964, n37965, n37966, n37967,
         n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975,
         n37976, n37977, n37978, n37979, n37980, n37981, n37982, n37983,
         n37984, n37985, n37986, n37987, n37988, n37989, n37990, n37991,
         n37992, n37993, n37994, n37995, n37996, n37997, n37998, n37999,
         n38000, n38001, n38002, n38003, n38004, n38005, n38006, n38007,
         n38008, n38009, n38010, n38011, n38012, n38013, n38014, n38015,
         n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023,
         n38024, n38025, n38026, n38027, n38028, n38029, n38030, n38031,
         n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039,
         n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047,
         n38048, n38049, n38050, n38051, n38052, n38053, n38054, n38055,
         n38056, n38057, n38058, n38059, n38060, n38061, n38062, n38063,
         n38064, n38065, n38066, n38067, n38068, n38069, n38070, n38071,
         n38072, n38073, n38074, n38075, n38076, n38077, n38078, n38079,
         n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087,
         n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095,
         n38096, n38097, n38098, n38099, n38100, n38101, n38102, n38103,
         n38104, n38105, n38106, n38107, n38108, n38109, n38110, n38111,
         n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119,
         n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38127,
         n38128, n38129, n38130, n38131, n38132, n38133, n38134, n38135,
         n38136, n38137, n38138, n38139, n38140, n38141, n38142, n38143,
         n38144, n38145, n38146, n38147, n38148, n38149, n38150, n38151,
         n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159,
         n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167,
         n38168, n38169, n38170, n38171, n38173, n38174, n38175, n38176,
         n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184,
         n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192,
         n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200,
         n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208,
         n38209, n38210, n38211, n38212, n38213, n38214, n38215, n38216,
         n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224,
         n38225, n38226, n38227, n38228, n38231, n38232, n38233, n38234,
         n38235, n38236, n38237, n38239, n38240, n38241, n38242, n38243,
         n38244, n38245, n38246, n38247, n38248, n38249, n38250, n38251,
         n38252, n38253, n38254, n38255, n38256, n38257, n38258, n38259,
         n38260, n38261, n38262, n38263, n38264, n38265, n38266, n38267,
         n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275,
         n38276, n38277, n38278, n38279, n38280, n38281, n38282, n38283,
         n38284, n38285, n38286, n38287, n38288, n38289, n38290, n38291,
         n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299,
         n38300, n38301, n38302, n38303, n38304, n38305, n38306, n38307,
         n38308, n38309, n38310, n38311, n38312, n38313, n38314, n38315,
         n38316, n38317, n38318, n38319, n38320, n38321, n38322, n38323,
         n38324, n38325, n38326, n38327, n38328, n38329, n38330, n38331,
         n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339,
         n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347,
         n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355,
         n38356, n38357, n38358, n38359, n38360, n38361, n38362, n38363,
         n38364, n38365, n38366, n38367, n38368, n38369, n38370, n38371,
         n38372, n38373, n38374, n38375, n38376, n38377, n38378, n38379,
         n38380, n38381, n38382, n38383, n38384, n38385, n38386, n38387,
         n38388, n38389, n38390, n38391, n38392, n38393, n38394, n38395,
         n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38404,
         n38405, n38406, n38407, n38408, n38409, n38410, n38412, n38413,
         n38414, n38415, n38416, n38417, n38418, n38419, n38420, n38421,
         n38422, n38423, n38424, n38425, n38426, n38427, n38428, n38429,
         n38430, n38431, n38432, n38434, n38435, n38436, n38438, n38439,
         n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447,
         n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455,
         n38456, n38457, n38458, n38459, n38460, n38461, n38462, n38463,
         n38464, n38465, n38467, n38468, n38469, n38470, n38471, n38472,
         n38473, n38474, n38475, n38476, n38477, n38478, n38479, n38480,
         n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488,
         n38489, n38490, n38491, n38492, n38493, n38494, n38495, n38496,
         n38497, n38498, n38499, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38528, n38529, n38530,
         n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538,
         n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546,
         n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38555,
         n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563,
         n38564, n38565, n38566, n38567, n38568, n38569, n38570, n38571,
         n38572, n38573, n38574, n38575, n38576, n38577, n38578, n38579,
         n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587,
         n38588, n38589, n38590, n38591, n38592, n38593, n38594, n38595,
         n38596, n38597, n38598, n38599, n38600, n38601, n38602, n38603,
         n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611,
         n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619,
         n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627,
         n38628, n38629, n38630, n38631, n38632, n38633, n38635, n38636,
         n38637, n38638, n38639, n38640, n38641, n38642, n38643, n38644,
         n38645, n38646, n38647, n38648, n38649, n38650, n38651, n38652,
         n38653, n38654, n38655, n38656, n38657, n38658, n38659, n38660,
         n38661, n38662, n38663, n38664, n38665, n38666, n38667, n38668,
         n38669, n38670, n38672, n38673, n38674, n38675, n38676, n38677,
         n38678, n38679, n38680, n38681, n38682, n38683, n38684, n38685,
         n38686, n38687, n38688, n38689, n38690, n38691, n38692, n38693,
         n38694, n38695, n38696, n38697, n38698, n38699, n38700, n38701,
         n38702, n38703, n38704, n38706, n38707, n38708, n38710, n38711,
         n38712, n38713, n38714, n38715, n38716, n38717, n38718, n38719,
         n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727,
         n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38736,
         n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744,
         n38745, n38746, n38747, n38749, n38750, n38751, n38752, n38753,
         n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
         n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769,
         n38770, n38772, n38773, n38774, n38775, n38776, n38777, n38778,
         n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786,
         n38787, n38788, n38789, n38790, n38791, n38793, n38794, n38795,
         n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803,
         n38804, n38805, n38806, n38807, n38808, n38809, n38810, n38811,
         n38812, n38813, n38814, n38815, n38816, n38817, n38818, n38819,
         n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827,
         n38828, n38830, n38831, n38832, n38833, n38834, n38835, n38836,
         n38837, n38838, n38839, n38840, n38841, n38842, n38843, n38844,
         n38845, n38846, n38847, n38848, n38849, n38850, n38851, n38852,
         n38853, n38854, n38855, n38856, n38857, n38858, n38859, n38860,
         n38861, n38862, n38863, n38864, n38865, n38866, n38867, n38868,
         n38869, n38870, n38871, n38872, n38873, n38874, n38875, n38876,
         n38877, n38878, n38879, n38880, n38881, n38882, n38883, n38884,
         n38885, n38886, n38887, n38888, n38889, n38890, n38891, n38892,
         n38893, n38894, n38895, n38896, n38897, n38898, n38899, n38900,
         n38901, n38902, n38903, n38904, n38905, n38906, n38907, n38908,
         n38909, n38910, n38911, n38912, n38913, n38914, n38915, n38916,
         n38917, n38918, n38919, n38920, n38921, n38922, n38923, n38924,
         n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932,
         n38933, n38934, n38935, n38936, n38937, n38938, n38939, n38940,
         n38941, n38942, n38943, n38944, n38946, n38947, n38949, n38950,
         n38951, n38952, n38953, n38954, n38955, n38957, n38958, n38959,
         n38960, n38961, n38962, n38963, n38964, n38965, n38966, n38967,
         n38968, n38969, n38970, n38971, n38972, n38973, n38974, n38975,
         n38976, n38977, n38978, n38979, n38980, n38981, n38982, n38983,
         n38984, n38985, n38986, n38987, n38988, n38989, n38990, n38991,
         n38992, n38993, n38994, n38995, n38996, n38997, n38998, n38999,
         n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007,
         n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015,
         n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023,
         n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031,
         n39032, n39033, n39034, n39035, n39036, n39037, n39038, n39039,
         n39040, n39041, n39042, n39043, n39044, n39045, n39046, n39047,
         n39048, n39049, n39050, n39051, n39052, n39053, n39054, n39055,
         n39056, n39057, n39058, n39059, n39060, n39062, n39063, n39064,
         n39065, n39066, n39067, n39068, n39069, n39070, n39071, n39072,
         n39073, n39074, n39076, n39077, n39078, n39079, n39081, n39082,
         n39083, n39084, n39085, n39086, n39087, n39088, n39089, n39090,
         n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098,
         n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106,
         n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114,
         n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122,
         n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130,
         n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138,
         n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146,
         n39147, n39148, n39150, n39151, n39152, n39153, n39154, n39155,
         n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39163,
         n39164, n39165, n39166, n39167, n39168, n39169, n39170, n39171,
         n39172, n39173, n39174, n39175, n39176, n39177, n39178, n39179,
         n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187,
         n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195,
         n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203,
         n39204, n39205, n39206, n39207, n39208, n39210, n39211, n39212,
         n39213, n39214, n39215, n39216, n39217, n39218, n39219, n39220,
         n39221, n39222, n39223, n39224, n39225, n39226, n39227, n39228,
         n39229, n39230, n39231, n39232, n39233, n39234, n39235, n39236,
         n39237, n39238, n39239, n39240, n39242, n39243, n39244, n39245,
         n39246, n39247, n39249, n39250, n39251, n39252, n39253, n39254,
         n39255, n39256, n39257, n39258, n39259, n39260, n39261, n39262,
         n39263, n39264, n39265, n39266, n39267, n39268, n39269, n39270,
         n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278,
         n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286,
         n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294,
         n39295, n39296, n39298, n39299, n39300, n39301, n39302, n39303,
         n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311,
         n39312, n39313, n39314, n39316, n39317, n39318, n39319, n39320,
         n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328,
         n39329, n39330, n39331, n39332, n39333, n39334, n39335, n39336,
         n39337, n39338, n39339, n39340, n39341, n39342, n39343, n39344,
         n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352,
         n39353, n39354, n39355, n39356, n39358, n39359, n39360, n39361,
         n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369,
         n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377,
         n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39386,
         n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394,
         n39395, n39396, n39397, n39399, n39400, n39401, n39402, n39403,
         n39405, n39406, n39407, n39408, n39409, n39410, n39411, n39412,
         n39413, n39414, n39415, n39416, n39417, n39418, n39419, n39420,
         n39421, n39422, n39423, n39424, n39425, n39426, n39427, n39428,
         n39429, n39430, n39431, n39432, n39434, n39436, n39437, n39438,
         n39439, n39441, n39442, n39443, n39444, n39445, n39446, n39447,
         n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455,
         n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463,
         n39464, n39465, n39466, n39467, n39468, n39469, n39470, n39471,
         n39472, n39473, n39474, n39475, n39476, n39477, n39478, n39479,
         n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488,
         n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496,
         n39497, n39498, n39499, n39500, n39501, n39502, n39503, n39504,
         n39505, n39506, n39507, n39508, n39509, n39510, n39511, n39512,
         n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520,
         n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528,
         n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536,
         n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544,
         n39545, n39546, n39547, n39548, n39549, n39551, n39552, n39553,
         n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561,
         n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569,
         n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577,
         n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585,
         n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593,
         n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601,
         n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609,
         n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617,
         n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625,
         n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39636,
         n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644,
         n39645, n39646, n39647, n39648, n39649, n39650, n39651, n39652,
         n39653, n39654, n39655, n39656, n39657, n39658, n39660, n39661,
         n39662, n39663, n39664, n39665, n39666, n39667, n39668, n39669,
         n39670, n39671, n39672, n39673, n39674, n39675, n39676, n39677,
         n39678, n39679, n39680, n39681, n39682, n39683, n39684, n39685,
         n39686, n39687, n39688, n39689, n39690, n39691, n39692, n39693,
         n39694, n39695, n39696, n39697, n39698, n39699, n39700, n39701,
         n39702, n39703, n39704, n39705, n39706, n39707, n39708, n39709,
         n39710, n39711, n39712, n39713, n39714, n39715, n39716, n39717,
         n39718, n39719, n39720, n39721, n39722, n39723, n39724, n39725,
         n39726, n39727, n39728, n39730, n39731, n39732, n39733, n39734,
         n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742,
         n39743, n39744, n39746, n39747, n39748, n39749, n39750, n39751,
         n39752, n39753, n39754, n39755, n39756, n39757, n39758, n39759,
         n39760, n39761, n39762, n39763, n39764, n39765, n39766, n39767,
         n39768, n39769, n39770, n39771, n39772, n39774, n39775, n39776,
         n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784,
         n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792,
         n39793, n39794, n39795, n39796, n39797, n39799, n39800, n39801,
         n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809,
         n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
         n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825,
         n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833,
         n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841,
         n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849,
         n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857,
         n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865,
         n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873,
         n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881,
         n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
         n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897,
         n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905,
         n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913,
         n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921,
         n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929,
         n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937,
         n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39946,
         n39947, n39948, n39949, n39950, n39951, n39952, n39953, n39954,
         n39955, n39956, n39957, n39958, n39959, n39960, n39961, n39962,
         n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970,
         n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978,
         n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986,
         n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994,
         n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002,
         n40003, n40004, n40005, n40006, n40007, n40008, n40009, n40010,
         n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018,
         n40019, n40020, n40021, n40022, n40023, n40024, n40025, n40026,
         n40027, n40028, n40029, n40030, n40031, n40032, n40033, n40034,
         n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042,
         n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050,
         n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058,
         n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066,
         n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074,
         n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082,
         n40083, n40084, n40085, n40087, n40088, n40089, n40090, n40091,
         n40092, n40093, n40094, n40095, n40096, n40097, n40098, n40099,
         n40100, n40101, n40102, n40103, n40104, n40105, n40106, n40107,
         n40108, n40110, n40111, n40112, n40113, n40114, n40115, n40116,
         n40118, n40119, n40120, n40121, n40122, n40123, n40124, n40125,
         n40126, n40127, n40128, n40129, n40130, n40131, n40132, n40133,
         n40134, n40136, n40137, n40138, n40139, n40140, n40141, n40142,
         n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40151,
         n40153, n40154, n40155, n40156, n40157, n40158, n40159, n40160,
         n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168,
         n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176,
         n40177, n40178, n40179, n40180, n40181, n40182, n40184, n40185,
         n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
         n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201,
         n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209,
         n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217,
         n40218, n40219, n40221, n40222, n40223, n40224, n40225, n40226,
         n40227, n40228, n40229, n40230, n40231, n40232, n40233, n40234,
         n40235, n40236, n40237, n40238, n40239, n40240, n40241, n40242,
         n40243, n40244, n40245, n40246, n40247, n40248, n40249, n40250,
         n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258,
         n40259, n40261, n40262, n40263, n40264, n40265, n40266, n40267,
         n40268, n40269, n40271, n40272, n40273, n40274, n40275, n40276,
         n40277, n40278, n40279, n40280, n40281, n40282, n40283, n40284,
         n40285, n40286, n40287, n40288, n40289, n40290, n40291, n40292,
         n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300,
         n40301, n40302, n40303, n40304, n40305, n40306, n40307, n40308,
         n40309, n40310, n40311, n40312, n40313, n40314, n40315, n40316,
         n40317, n40318, n40319, n40320, n40321, n40322, n40323, n40324,
         n40325, n40326, n40327, n40328, n40329, n40330, n40331, n40332,
         n40333, n40334, n40335, n40336, n40337, n40338, n40339, n40340,
         n40341, n40342, n40343, n40344, n40345, n40346, n40347, n40348,
         n40349, n40350, n40351, n40352, n40353, n40354, n40355, n40356,
         n40357, n40358, n40359, n40360, n40361, n40362, n40363, n40364,
         n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372,
         n40373, n40374, n40375, n40376, n40377, n40378, n40379, n40380,
         n40381, n40382, n40383, n40384, n40385, n40386, n40387, n40388,
         n40389, n40390, n40391, n40392, n40393, n40394, n40395, n40396,
         n40397, n40398, n40399, n40400, n40401, n40402, n40403, n40404,
         n40405, n40406, n40407, n40408, n40409, n40410, n40411, n40412,
         n40413, n40414, n40415, n40416, n40417, n40418, n40419, n40420,
         n40421, n40422, n40423, n40424, n40425, n40426, n40427, n40428,
         n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436,
         n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444,
         n40445, n40446, n40447, n40448, n40449, n40450, n40451, n40452,
         n40453, n40454, n40455, n40456, n40457, n40458, n40459, n40460,
         n40461, n40462, n40463, n40464, n40465, n40466, n40467, n40468,
         n40469, n40470, n40471, n40472, n40473, n40474, n40475, n40476,
         n40477, n40478, n40479, n40480, n40481, n40482, n40483, n40484,
         n40485, n40486, n40487, n40488, n40489, n40490, n40491, n40492,
         n40493, n40494, n40496, n40497, n40498, n40499, n40500, n40501,
         n40502, n40503, n40504, n40505, n40506, n40507, n40508, n40509,
         n40510, n40511, n40512, n40513, n40514, n40515, n40517, n40518,
         n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526,
         n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534,
         n40535, n40536, n40537, n40538, n40539, n40540, n40541, n40542,
         n40543, n40544, n40545, n40546, n40547, n40548, n40549, n40550,
         n40551, n40552, n40553, n40555, n40556, n40557, n40558, n40559,
         n40560, n40561, n40562, n40563, n40564, n40565, n40566, n40567,
         n40569, n40570, n40571, n40572, n40573, n40574, n40575, n40576,
         n40577, n40578, n40579, n40580, n40581, n40582, n40583, n40584,
         n40585, n40586, n40587, n40588, n40589, n40590, n40591, n40592,
         n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600,
         n40601, n40602, n40603, n40605, n40606, n40607, n40608, n40609,
         n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617,
         n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625,
         n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633,
         n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641,
         n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649,
         n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657,
         n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665,
         n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673,
         n40674, n40675, n40676, n40677, n40678, n40679, n40681, n40682,
         n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690,
         n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698,
         n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706,
         n40707, n40708, n40709, n40712, n40713, n40714, n40715, n40716,
         n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724,
         n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732,
         n40733, n40734, n40735, n40736, n40737, n40738, n40739, n40740,
         n40741, n40742, n40744, n40745, n40746, n40747, n40748, n40749,
         n40750, n40751, n40752, n40753, n40754, n40755, n40756, n40757,
         n40758, n40759, n40760, n40761, n40762, n40763, n40764, n40765,
         n40766, n40767, n40768, n40769, n40770, n40771, n40772, n40773,
         n40774, n40775, n40776, n40777, n40778, n40779, n40780, n40781,
         n40782, n40783, n40784, n40785, n40786, n40787, n40788, n40789,
         n40790, n40791, n40792, n40793, n40794, n40795, n40796, n40797,
         n40798, n40799, n40800, n40801, n40802, n40803, n40804, n40805,
         n40806, n40807, n40808, n40809, n40810, n40811, n40812, n40813,
         n40814, n40815, n40816, n40817, n40818, n40819, n40820, n40821,
         n40822, n40823, n40824, n40825, n40826, n40827, n40828, n40830,
         n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40838,
         n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846,
         n40847, n40848, n40849, n40850, n40851, n40852, n40853, n40854,
         n40855, n40856, n40857, n40858, n40859, n40860, n40861, n40862,
         n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870,
         n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878,
         n40879, n40880, n40881, n40882, n40883, n40884, n40885, n40886,
         n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894,
         n40895, n40896, n40897, n40898, n40899, n40900, n40901, n40902,
         n40903, n40904, n40905, n40906, n40907, n40908, n40909, n40910,
         n40911, n40912, n40913, n40914, n40915, n40916, n40917, n40918,
         n40919, n40920, n40921, n40922, n40923, n40924, n40925, n40926,
         n40927, n40928, n40929, n40930, n40931, n40932, n40933, n40934,
         n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942,
         n40943, n40944, n40945, n40946, n40947, n40948, n40949, n40950,
         n40951, n40952, n40953, n40954, n40955, n40956, n40957, n40958,
         n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966,
         n40967, n40968, n40969, n40970, n40971, n40972, n40974, n40975,
         n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983,
         n40984, n40985, n40986, n40988, n40989, n40990, n40991, n40992,
         n40993, n40994, n40995, n40996, n40997, n40998, n40999, n41000,
         n41001, n41002, n41003, n41004, n41006, n41007, n41008, n41009,
         n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41018,
         n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026,
         n41027, n41028, n41029, n41030, n41031, n41032, n41033, n41034,
         n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042,
         n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050,
         n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058,
         n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066,
         n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074,
         n41075, n41076, n41077, n41078, n41079, n41080, n41081, n41082,
         n41083, n41084, n41085, n41086, n41087, n41088, n41089, n41090,
         n41091, n41092, n41093, n41094, n41095, n41096, n41097, n41098,
         n41099, n41100, n41101, n41102, n41103, n41104, n41105, n41106,
         n41107, n41108, n41109, n41110, n41111, n41112, n41113, n41114,
         n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122,
         n41123, n41124, n41125, n41126, n41127, n41129, n41130, n41131,
         n41132, n41134, n41135, n41136, n41137, n41138, n41139, n41140,
         n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148,
         n41149, n41150, n41152, n41153, n41154, n41155, n41156, n41157,
         n41158, n41159, n41160, n41161, n41162, n41163, n41164, n41165,
         n41166, n41167, n41168, n41169, n41170, n41171, n41172, n41173,
         n41174, n41175, n41176, n41177, n41178, n41179, n41180, n41181,
         n41182, n41183, n41184, n41185, n41186, n41187, n41188, n41189,
         n41190, n41191, n41192, n41193, n41194, n41195, n41196, n41197,
         n41198, n41199, n41200, n41201, n41202, n41203, n41204, n41205,
         n41206, n41207, n41208, n41209, n41210, n41211, n41212, n41213,
         n41214, n41215, n41216, n41217, n41218, n41219, n41220, n41221,
         n41222, n41223, n41224, n41225, n41226, n41227, n41228, n41229,
         n41230, n41231, n41232, n41233, n41234, n41235, n41236, n41237,
         n41238, n41239, n41240, n41241, n41242, n41243, n41244, n41245,
         n41246, n41247, n41248, n41249, n41250, n41251, n41252, n41253,
         n41254, n41256, n41257, n41258, n41259, n41260, n41261, n41262,
         n41263, n41264, n41265, n41266, n41267, n41268, n41269, n41270,
         n41271, n41272, n41273, n41274, n41275, n41276, n41277, n41278,
         n41279, n41280, n41281, n41282, n41283, n41284, n41285, n41286,
         n41287, n41288, n41289, n41290, n41291, n41292, n41293, n41294,
         n41295, n41296, n41297, n41298, n41299, n41300, n41301, n41302,
         n41303, n41304, n41305, n41306, n41307, n41308, n41309, n41310,
         n41311, n41312, n41313, n41314, n41315, n41316, n41317, n41318,
         n41319, n41320, n41321, n41322, n41323, n41324, n41325, n41326,
         n41327, n41328, n41329, n41330, n41331, n41332, n41333, n41334,
         n41335, n41336, n41337, n41338, n41339, n41340, n41341, n41342,
         n41343, n41344, n41345, n41346, n41347, n41348, n41349, n41350,
         n41351, n41352, n41353, n41354, n41355, n41356, n41357, n41358,
         n41359, n41360, n41361, n41362, n41363, n41364, n41365, n41366,
         n41367, n41368, n41370, n41371, n41372, n41373, n41374, n41375,
         n41376, n41377, n41378, n41379, n41380, n41381, n41382, n41383,
         n41384, n41385, n41386, n41387, n41388, n41389, n41390, n41391,
         n41392, n41393, n41394, n41395, n41396, n41397, n41398, n41399,
         n41400, n41401, n41402, n41403, n41404, n41405, n41406, n41407,
         n41408, n41409, n41410, n41411, n41412, n41413, n41414, n41415,
         n41416, n41417, n41418, n41419, n41420, n41421, n41422, n41423,
         n41424, n41425, n41426, n41427, n41428, n41429, n41430, n41431,
         n41432, n41433, n41434, n41435, n41436, n41437, n41438, n41439,
         n41440, n41441, n41442, n41443, n41444, n41445, n41446, n41447,
         n41448, n41449, n41450, n41451, n41452, n41453, n41454, n41455,
         n41456, n41457, n41458, n41459, n41460, n41461, n41462, n41463,
         n41464, n41465, n41466, n41467, n41468, n41469, n41470, n41471,
         n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479,
         n41480, n41481, n41482, n41483, n41484, n41485, n41486, n41487,
         n41488, n41489, n41490, n41491, n41492, n41493, n41494, n41495,
         n41496, n41497, n41498, n41499, n41500, n41501, n41502, n41503,
         n41504, n41505, n41506, n41507, n41508, n41509, n41510, n41511,
         n41512, n41513, n41514, n41515, n41516, n41517, n41518, n41519,
         n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527,
         n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535,
         n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543,
         n41544, n41545, n41546, n41547, n41548, n41550, n41551, n41552,
         n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560,
         n41561, n41562, n41563, n41564, n41565, n41566, n41567, n41568,
         n41569, n41570, n41571, n41572, n41573, n41574, n41575, n41576,
         n41577, n41578, n41579, n41580, n41581, n41582, n41583, n41584,
         n41585, n41586, n41587, n41588, n41589, n41590, n41591, n41592,
         n41593, n41594, n41595, n41596, n41597, n41598, n41599, n41600,
         n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608,
         n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616,
         n41617, n41618, n41619, n41620, n41621, n41622, n41623, n41624,
         n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632,
         n41633, n41634, n41635, n41636, n41637, n41638, n41639, n41640,
         n41641, n41642, n41643, n41644, n41645, n41646, n41647, n41648,
         n41649, n41650, n41651, n41652, n41653, n41654, n41655, n41656,
         n41657, n41658, n41659, n41660, n41661, n41662, n41663, n41664,
         n41665, n41666, n41667, n41668, n41669, n41670, n41671, n41672,
         n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680,
         n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688,
         n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696,
         n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704,
         n41705, n41706, n41707, n41708, n41709, n41710, n41711, n41712,
         n41713, n41714, n41716, n41717, n41718, n41719, n41720, n41721,
         n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729,
         n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737,
         n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745,
         n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753,
         n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761,
         n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769,
         n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777,
         n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785,
         n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793,
         n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801,
         n41802, n41803, n41804, n41805, n41806, n41808, n41809, n41810,
         n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818,
         n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826,
         n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834,
         n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842,
         n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850,
         n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858,
         n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866,
         n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874,
         n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882,
         n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891,
         n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899,
         n41900, n41901, n41902, n41903, n41904, n41905, n41906, n41907,
         n41908, n41909, n41910, n41911, n41912, n41913, n41914, n41915,
         n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923,
         n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931,
         n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939,
         n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947,
         n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955,
         n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963,
         n41964, n41966, n41967, n41968, n41969, n41970, n41971, n41972,
         n41973, n41974, n41975, n41976, n41977, n41978, n41979, n41980,
         n41981, n41982, n41983, n41984, n41985, n41986, n41987, n41988,
         n41989, n41990, n41991, n41992, n41993, n41994, n41995, n41996,
         n41997, n41998, n41999, n42000, n42001, n42002, n42003, n42004,
         n42005, n42006, n42007, n42008, n42009, n42010, n42011, n42012,
         n42013, n42014, n42015, n42016, n42017, n42018, n42019, n42020,
         n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028,
         n42029, n42030, n42031, n42032, n42033, n42034, n42035, n42036,
         n42037, n42038, n42039, n42040, n42041, n42042, n42043, n42044,
         n42045, n42046, n42047, n42048, n42049, n42050, n42051, n42052,
         n42053, n42054, n42055, n42056, n42057, n42058, n42059, n42060,
         n42061, n42062, n42063, n42064, n42065, n42066, n42067, n42068,
         n42069, n42070, n42071, n42072, n42073, n42074, n42075, n42076,
         n42077, n42078, n42079, n42080, n42081, n42082, n42083, n42084,
         n42085, n42086, n42087, n42088, n42089, n42090, n42091, n42092,
         n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100,
         n42101, n42102, n42103, n42104, n42105, n42106, n42107, n42109,
         n42110, n42111, n42112, n42113, n42114, n42115, n42116, n42117,
         n42118, n42119, n42120, n42121, n42122, n42123, n42124, n42125,
         n42126, n42127, n42128, n42129, n42130, n42131, n42132, n42133,
         n42134, n42135, n42136, n42138, n42139, n42140, n42141, n42142,
         n42143, n42144, n42145, n42146, n42147, n42148, n42149, n42150,
         n42151, n42152, n42153, n42154, n42155, n42156, n42157, n42158,
         n42159, n42160, n42161, n42162, n42163, n42164, n42165, n42166,
         n42167, n42168, n42169, n42170, n42171, n42172, n42173, n42174,
         n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182,
         n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190,
         n42191, n42192, n42193, n42194, n42195, n42196, n42197, n42198,
         n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206,
         n42207, n42208, n42209, n42210, n42211, n42212, n42213, n42214,
         n42215, n42216, n42217, n42218, n42219, n42220, n42221, n42222,
         n42223, n42224, n42225, n42226, n42227, n42228, n42229, n42230,
         n42231, n42232, n42233, n42234, n42235, n42236, n42237, n42238,
         n42239, n42240, n42241, n42242, n42243, n42244, n42245, n42246,
         n42247, n42248, n42250, n42251, n42253, n42254, n42255, n42256,
         n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264,
         n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272,
         n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280,
         n42281, n42282, n42283, n42284, n42285, n42286, n42287, n42289,
         n42290, n42291, n42292, n42293, n42294, n42295, n42296, n42297,
         n42298, n42299, n42300, n42301, n42302, n42303, n42304, n42305,
         n42306, n42307, n42308, n42309, n42310, n42311, n42312, n42313,
         n42314, n42315, n42316, n42317, n42318, n42319, n42320, n42321,
         n42322, n42323, n42324, n42326, n42327, n42328, n42329, n42330,
         n42331, n42332, n42333, n42334, n42335, n42336, n42337, n42338,
         n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346,
         n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354,
         n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362,
         n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370,
         n42371, n42372, n42373, n42374, n42375, n42376, n42377, n42378,
         n42379, n42380, n42381, n42382, n42383, n42384, n42385, n42386,
         n42387, n42388, n42389, n42390, n42391, n42392, n42393, n42394,
         n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402,
         n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410,
         n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418,
         n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426,
         n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434,
         n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442,
         n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450,
         n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458,
         n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466,
         n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474,
         n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482,
         n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490,
         n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498,
         n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506,
         n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514,
         n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522,
         n42523, n42524, n42525, n42526, n42527, n42528, n42529, n42530,
         n42531, n42532, n42533, n42534, n42535, n42537, n42538, n42539,
         n42540, n42541, n42542, n42543, n42544, n42545, n42546, n42547,
         n42548, n42549, n42550, n42551, n42552, n42553, n42554, n42555,
         n42556, n42557, n42558, n42559, n42560, n42561, n42562, n42563,
         n42564, n42565, n42566, n42567, n42568, n42569, n42570, n42571,
         n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579,
         n42580, n42581, n42582, n42583, n42584, n42585, n42587, n42588,
         n42589, n42590, n42591, n42592, n42593, n42594, n42595, n42596,
         n42597, n42598, n42599, n42600, n42602, n42603, n42604, n42605,
         n42606, n42607, n42608, n42609, n42610, n42611, n42612, n42613,
         n42614, n42615, n42616, n42617, n42618, n42619, n42620, n42621,
         n42622, n42623, n42624, n42625, n42626, n42628, n42629, n42630,
         n42631, n42632, n42633, n42634, n42635, n42636, n42637, n42638,
         n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646,
         n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654,
         n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662,
         n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670,
         n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678,
         n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686,
         n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694,
         n42695, n42696, n42697, n42698, n42699, n42700, n42701, n42702,
         n42703, n42704, n42705, n42706, n42707, n42708, n42709, n42710,
         n42711, n42712, n42713, n42714, n42715, n42716, n42717, n42718,
         n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726,
         n42727, n42728, n42729, n42730, n42731, n42732, n42733, n42734,
         n42735, n42736, n42737, n42738, n42739, n42740, n42741, n42742,
         n42743, n42744, n42745, n42746, n42748, n42749, n42750, n42751,
         n42752, n42753, n42754, n42755, n42756, n42757, n42758, n42759,
         n42760, n42761, n42762, n42763, n42764, n42765, n42766, n42767,
         n42768, n42769, n42770, n42771, n42772, n42773, n42774, n42775,
         n42776, n42777, n42778, n42779, n42780, n42781, n42782, n42783,
         n42784, n42785, n42786, n42787, n42788, n42789, n42790, n42791,
         n42792, n42793, n42794, n42795, n42796, n42797, n42798, n42799,
         n42800, n42801, n42802, n42803, n42804, n42805, n42807, n42808,
         n42809, n42810, n42811, n42812, n42813, n42814, n42815, n42816,
         n42817, n42818, n42819, n42820, n42821, n42822, n42823, n42824,
         n42825, n42826, n42827, n42828, n42829, n42830, n42831, n42832,
         n42833, n42834, n42835, n42836, n42837, n42839, n42840, n42841,
         n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849,
         n42850, n42851, n42852, n42853, n42854, n42855, n42856, n42857,
         n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865,
         n42866, n42867, n42868, n42869, n42870, n42871, n42872, n42873,
         n42874, n42875, n42876, n42877, n42878, n42879, n42880, n42881,
         n42882, n42883, n42884, n42885, n42886, n42887, n42888, n42889,
         n42890, n42891, n42892, n42893, n42894, n42895, n42896, n42897,
         n42898, n42899, n42900, n42901, n42902, n42903, n42904, n42905,
         n42906, n42907, n42908, n42909, n42910, n42911, n42912, n42913,
         n42914, n42915, n42916, n42917, n42918, n42919, n42920, n42921,
         n42922, n42923, n42924, n42925, n42926, n42927, n42928, n42930,
         n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938,
         n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946,
         n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42955,
         n42956, n42957, n42958, n42959, n42960, n42961, n42962, n42963,
         n42964, n42965, n42966, n42967, n42968, n42969, n42970, n42971,
         n42972, n42973, n42974, n42975, n42976, n42977, n42978, n42979,
         n42980, n42981, n42982, n42983, n42984, n42985, n42986, n42987,
         n42988, n42989, n42990, n42991, n42992, n42993, n42994, n42995,
         n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003,
         n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011,
         n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019,
         n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027,
         n43028, n43029, n43030, n43031, n43032, n43033, n43034, n43035,
         n43036, n43037, n43038, n43039, n43040, n43041, n43042, n43043,
         n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051,
         n43052, n43053, n43054, n43055, n43056, n43057, n43058, n43059,
         n43060, n43061, n43062, n43063, n43064, n43065, n43066, n43067,
         n43068, n43069, n43070, n43071, n43072, n43073, n43074, n43075,
         n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083,
         n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091,
         n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099,
         n43100, n43101, n43102, n43103, n43104, n43105, n43106, n43107,
         n43108, n43109, n43110, n43111, n43112, n43113, n43114, n43115,
         n43116, n43117, n43118, n43119, n43120, n43121, n43122, n43123,
         n43124, n43125, n43126, n43127, n43128, n43129, n43130, n43131,
         n43132, n43133, n43134, n43135, n43136, n43137, n43138, n43139,
         n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147,
         n43148, n43149, n43150, n43151, n43152, n43153, n43154, n43155,
         n43156, n43157, n43158, n43159, n43160, n43161, n43162, n43163,
         n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171,
         n43172, n43173, n43174, n43175, n43176, n43177, n43178, n43179,
         n43180, n43181, n43182, n43183, n43184, n43185, n43186, n43187,
         n43188, n43189, n43190, n43191, n43192, n43193, n43194, n43195,
         n43196, n43197, n43198, n43199, n43200, n43201, n43202, n43203,
         n43204, n43205, n43206, n43207, n43208, n43209, n43210, n43211,
         n43212, n43213, n43214, n43215, n43216, n43217, n43218, n43219,
         n43220, n43221, n43222, n43223, n43224, n43225, n43226, n43227,
         n43228, n43229, n43230, n43231, n43232, n43233, n43234, n43235,
         n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243,
         n43244, n43245, n43246, n43247, n43248, n43249, n43250, n43251,
         n43252, n43253, n43254, n43255, n43256, n43257, n43258, n43259,
         n43260, n43261, n43262, n43263, n43264, n43265, n43266, n43267,
         n43268, n43269, n43270, n43271, n43272, n43273, n43274, n43275,
         n43276, n43277, n43278, n43279, n43280, n43281, n43282, n43283,
         n43284, n43285, n43286, n43287, n43288, n43289, n43290, n43291,
         n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299,
         n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307,
         n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315,
         n43316, n43317, n43318, n43319, n43320, n43321, n43322, n43323,
         n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331,
         n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339,
         n43340, n43341, n43342, n43343, n43344, n43345, n43346, n43347,
         n43348, n43349, n43350, n43351, n43352, n43353, n43354, n43355,
         n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363,
         n43364, n43365, n43366, n43368, n43369, n43370, n43371, n43372,
         n43373, n43374, n43375, n43376, n43377, n43378, n43379, n43380,
         n43381, n43382, n43383, n43384, n43385, n43386, n43387, n43388,
         n43389, n43390, n43391, n43392, n43393, n43394, n43395, n43396,
         n43398, n43399, n43400, n43401, n43402, n43403, n43404, n43405,
         n43406, n43407, n43408, n43409, n43410, n43411, n43412, n43413,
         n43414, n43415, n43416, n43417, n43419, n43420, n43421, n43422,
         n43423, n43424, n43425, n43426, n43427, n43428, n43429, n43430,
         n43431, n43432, n43433, n43434, n43435, n43436, n43437, n43438,
         n43440, n43442, n43443, n43444, n43445, n43446, n43447, n43448,
         n43449, n43450, n43451, n43452, n43453, n43454, n43455, n43456,
         n43457, n43458, n43459, n43460, n43461, n43462, n43463, n43464,
         n43465, n43466, n43467, n43468, n43469, n43470, n43471, n43472,
         n43473, n43474, n43475, n43476, n43477, n43478, n43479, n43480,
         n43481, n43482, n43483, n43484, n43485, n43486, n43487, n43488,
         n43489, n43490, n43491, n43492, n43493, n43494, n43495, n43496,
         n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505,
         n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513,
         n43514, n43515, n43516, n43517, n43518, n43519, n43520, n43521,
         n43522, n43523, n43524, n43525, n43526, n43527, n43528, n43529,
         n43530, n43531, n43532, n43533, n43534, n43536, n43537, n43538,
         n43539, n43540, n43541, n43542, n43543, n43544, n43545, n43546,
         n43547, n43548, n43549, n43550, n43551, n43552, n43553, n43554,
         n43555, n43556, n43557, n43558, n43559, n43560, n43561, n43562,
         n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570,
         n43571, n43572, n43573, n43574, n43575, n43577, n43578, n43579,
         n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587,
         n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595,
         n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603,
         n43604, n43605, n43606, n43607, n43608, n43609, n43610, n43611,
         n43612, n43613, n43614, n43615, n43616, n43617, n43618, n43619,
         n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627,
         n43628, n43629, n43630, n43631, n43632, n43633, n43634, n43635,
         n43636, n43637, n43638, n43639, n43640, n43641, n43642, n43643,
         n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651,
         n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659,
         n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667,
         n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675,
         n43676, n43677, n43678, n43679, n43680, n43681, n43682, n43683,
         n43684, n43685, n43686, n43687, n43688, n43689, n43690, n43691,
         n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699,
         n43700, n43701, n43702, n43703, n43704, n43705, n43706, n43707,
         n43708, n43709, n43710, n43711, n43712, n43713, n43714, n43715,
         n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723,
         n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731,
         n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739,
         n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747,
         n43748, n43749, n43750, n43751, n43752, n43753, n43754, n43755,
         n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763,
         n43764, n43765, n43766, n43767, n43768, n43769, n43770, n43771,
         n43772, n43773, n43774, n43775, n43776, n43777, n43778, n43779,
         n43780, n43781, n43782, n43783, n43784, n43785, n43786, n43787,
         n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795,
         n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803,
         n43804, n43805, n43806, n43807, n43808, n43809, n43810, n43811,
         n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819,
         n43820, n43821, n43822, n43823, n43824, n43825, n43826, n43827,
         n43828, n43829, n43830, n43831, n43832, n43833, n43834, n43835,
         n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843,
         n43844, n43845, n43846, n43848, n43849, n43850, n43851, n43852,
         n43853, n43854, n43855, n43856, n43857, n43858, n43859, n43860,
         n43861, n43862, n43863, n43864, n43865, n43866, n43867, n43868,
         n43869, n43870, n43871, n43872, n43873, n43874, n43875, n43876,
         n43877, n43878, n43879, n43880, n43881, n43882, n43883, n43884,
         n43885, n43886, n43887, n43888, n43889, n43890, n43891, n43892,
         n43893, n43894, n43895, n43896, n43897, n43898, n43899, n43900,
         n43901, n43902, n43903, n43904, n43905, n43906, n43907, n43908,
         n43909, n43910, n43911, n43912, n43913, n43914, n43915, n43916,
         n43917, n43918, n43919, n43920, n43921, n43922, n43923, n43924,
         n43925, n43926, n43927, n43928, n43929, n43930, n43931, n43932,
         n43933, n43934, n43935, n43936, n43937, n43938, n43939, n43940,
         n43941, n43942, n43943, n43944, n43945, n43946, n43947, n43948,
         n43949, n43950, n43951, n43952, n43953, n43954, n43955, n43956,
         n43957, n43958, n43959, n43960, n43961, n43962, n43963, n43964,
         n43965, n43966, n43967, n43968, n43969, n43970, n43971, n43972,
         n43973, n43974, n43975, n43976, n43977, n43978, n43979, n43980,
         n43981, n43982, n43983, n43984, n43985, n43986, n43987, n43988,
         n43989, n43990, n43991, n43992, n43993, n43994, n43995, n43996,
         n43997, n43998, n43999, n44000, n44001, n44002, n44003, n44004,
         n44005, n44006, n44007, n44008, n44009, n44010, n44011, n44012,
         n44013, n44014, n44015, n44016, n44017, n44018, n44019, n44020,
         n44021, n44022, n44023, n44024, n44025, n44026, n44027, n44028,
         n44029, n44030, n44031, n44032, n44033, n44034, n44035, n44036,
         n44037, n44038, n44039, n44040, n44041, n44042, n44043, n44044,
         n44045, n44046, n44047, n44048, n44049, n44050, n44051, n44052,
         n44053, n44054, n44055, n44056, n44057, n44058, n44059, n44060,
         n44061, n44062, n44063, n44064, n44065, n44066, n44067, n44068,
         n44069, n44070, n44071, n44072, n44073, n44074, n44075, n44076,
         n44077, n44078, n44079, n44080, n44081, n44082, n44083, n44084,
         n44085, n44086, n44087, n44088, n44089, n44090, n44091, n44092,
         n44093, n44094, n44095, n44096, n44097, n44098, n44099, n44100,
         n44101, n44102, n44103, n44104, n44105, n44106, n44107, n44108,
         n44109, n44110, n44111, n44112, n44113, n44114, n44115, n44116,
         n44117, n44118, n44119, n44120, n44121, n44122, n44124, n44125,
         n44126, n44127, n44128, n44129, n44130, n44131, n44132, n44133,
         n44134, n44135, n44136, n44137, n44138, n44139, n44140, n44141,
         n44142, n44143, n44144, n44145, n44146, n44147, n44148, n44149,
         n44150, n44151, n44152, n44153, n44154, n44155, n44156, n44157,
         n44158, n44159, n44160, n44161, n44162, n44163, n44164, n44165,
         n44166, n44167, n44168, n44169, n44170, n44171, n44172, n44173,
         n44174, n44175, n44176, n44177, n44178, n44179, n44180, n44181,
         n44182, n44183, n44184, n44185, n44186, n44187, n44188, n44189,
         n44190, n44191, n44192, n44193, n44194, n44195, n44196, n44197,
         n44198, n44199, n44200, n44201, n44202, n44203, n44204, n44205,
         n44206, n44207, n44208, n44209, n44210, n44211, n44213, n44214,
         n44215, n44216, n44217, n44218, n44219, n44220, n44221, n44222,
         n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230,
         n44231, n44232, n44233, n44234, n44235, n44236, n44237, n44238,
         n44239, n44240, n44241, n44242, n44243, n44244, n44245, n44246,
         n44248, n44249, n44250, n44251, n44252, n44253, n44254, n44255,
         n44256, n44257, n44258, n44259, n44260, n44261, n44262, n44263,
         n44264, n44265, n44266, n44267, n44268, n44269, n44270, n44271,
         n44272, n44273, n44274, n44275, n44276, n44277, n44278, n44279,
         n44280, n44281, n44282, n44283, n44284, n44285, n44286, n44287,
         n44288, n44289, n44290, n44291, n44292, n44293, n44294, n44295,
         n44296, n44297, n44298, n44299, n44300, n44301, n44302, n44303,
         n44304, n44305, n44306, n44307, n44308, n44309, n44310, n44311,
         n44312, n44313, n44314, n44315, n44316, n44317, n44318, n44319,
         n44320, n44321, n44322, n44323, n44324, n44325, n44326, n44327,
         n44328, n44329, n44330, n44331, n44332, n44333, n44334, n44335,
         n44336, n44337, n44338, n44339, n44340, n44341, n44342, n44343,
         n44344, n44345, n44346, n44347, n44348, n44349, n44350, n44351,
         n44353, n44354, n44355, n44356, n44357, n44358, n44359, n44360,
         n44361, n44362, n44363, n44364, n44365, n44366, n44367, n44368,
         n44369, n44370, n44371, n44372, n44373, n44374, n44375, n44376,
         n44377, n44378, n44379, n44380, n44381, n44382, n44383, n44384,
         n44385, n44386, n44387, n44388, n44389, n44390, n44391, n44392,
         n44393, n44394, n44395, n44396, n44397, n44398, n44399, n44400,
         n44401, n44402, n44403, n44404, n44405, n44406, n44407, n44408,
         n44409, n44410, n44411, n44412, n44413, n44414, n44415, n44416,
         n44417, n44418, n44419, n44420, n44421, n44422, n44423, n44424,
         n44425, n44426, n44427, n44428, n44429, n44430, n44431, n44432,
         n44433, n44434, n44435, n44436, n44437, n44438, n44439, n44440,
         n44441, n44442, n44443, n44444, n44445, n44446, n44447, n44448,
         n44449, n44450, n44451, n44452, n44453, n44454, n44455, n44456,
         n44457, n44458, n44459, n44460, n44461, n44462, n44463, n44464,
         n44465, n44466, n44467, n44468, n44469, n44470, n44471, n44472,
         n44473, n44474, n44475, n44476, n44477, n44478, n44479, n44480,
         n44481, n44482, n44483, n44484, n44485, n44486, n44487, n44488,
         n44489, n44490, n44491, n44493, n44494, n44495, n44496, n44497,
         n44498, n44499, n44500, n44501, n44502, n44503, n44504, n44505,
         n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513,
         n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44521,
         n44522, n44523, n44524, n44525, n44526, n44527, n44528, n44529,
         n44530, n44531, n44532, n44533, n44534, n44535, n44536, n44537,
         n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545,
         n44546, n44547, n44548, n44549, n44550, n44551, n44552, n44553,
         n44554, n44555, n44556, n44557, n44558, n44559, n44560, n44561,
         n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569,
         n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577,
         n44578, n44579, n44580, n44581, n44582, n44583, n44584, n44585,
         n44586, n44587, n44588, n44589, n44590, n44591, n44592, n44593,
         n44594, n44595, n44596, n44597, n44598, n44599, n44600, n44601,
         n44602, n44603, n44604, n44605, n44606, n44607, n44608, n44609,
         n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617,
         n44618, n44619, n44620, n44621, n44622, n44623, n44624, n44625,
         n44626, n44627, n44628, n44629, n44630, n44631, n44632, n44633,
         n44634, n44635, n44636, n44637, n44638, n44640, n44641, n44642,
         n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650,
         n44651, n44652, n44653, n44654, n44655, n44657, n44658, n44659,
         n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667,
         n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675,
         n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683,
         n44684, n44685, n44686, n44687, n44688, n44689, n44690, n44691,
         n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699,
         n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707,
         n44708, n44709, n44710, n44711, n44712, n44713, n44714, n44715,
         n44716, n44717, n44718, n44720, n44721, n44722, n44723, n44724,
         n44725, n44726, n44727, n44728, n44729, n44730, n44731, n44732,
         n44733, n44734, n44735, n44736, n44737, n44738, n44739, n44740,
         n44741, n44742, n44743, n44744, n44745, n44746, n44747, n44748,
         n44750, n44751, n44752, n44753, n44754, n44755, n44756, n44757,
         n44758, n44759, n44760, n44761, n44762, n44763, n44764, n44765,
         n44766, n44767, n44768, n44769, n44770, n44771, n44772, n44773,
         n44774, n44775, n44776, n44777, n44778, n44779, n44780, n44781,
         n44782, n44783, n44784, n44785, n44786, n44787, n44788, n44789,
         n44790, n44791, n44792, n44793, n44794, n44795, n44796, n44797,
         n44798, n44799, n44800, n44801, n44802, n44803, n44804, n44805,
         n44806, n44807, n44808, n44809, n44810, n44811, n44812, n44813,
         n44814, n44815, n44816, n44817, n44818, n44819, n44820, n44821,
         n44822, n44823, n44825, n44826, n44827, n44828, n44829, n44830,
         n44831, n44832, n44833, n44835, n44836, n44837, n44838, n44839,
         n44840, n44841, n44842, n44843, n44844, n44845, n44846, n44847,
         n44848, n44850, n44851, n44852, n44853, n44854, n44855, n44856,
         n44857, n44858, n44859, n44860, n44861, n44862, n44863, n44864,
         n44865, n44866, n44867, n44868, n44869, n44870, n44871, n44872,
         n44873, n44874, n44875, n44876, n44877, n44878, n44879, n44880,
         n44881, n44882, n44883, n44884, n44885, n44886, n44887, n44888,
         n44889, n44890, n44891, n44892, n44893, n44894, n44895, n44896,
         n44897, n44898, n44900, n44901, n44902, n44903, n44904, n44905,
         n44906, n44907, n44908, n44909, n44910, n44911, n44912, n44913,
         n44914, n44915, n44916, n44917, n44918, n44919, n44920, n44921,
         n44922, n44923, n44924, n44925, n44926, n44927, n44928, n44929,
         n44930, n44931, n44932, n44933, n44934, n44935, n44936, n44937,
         n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946,
         n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954,
         n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962,
         n44963, n44964, n44965, n44966, n44967, n44968, n44969, n44970,
         n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978,
         n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986,
         n44987, n44988, n44989, n44990, n44991, n44992, n44993, n44994,
         n44995, n44996, n44997, n44998, n44999, n45000, n45001, n45002,
         n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010,
         n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018,
         n45019, n45020, n45021, n45022, n45024, n45025, n45026, n45027,
         n45028, n45029, n45030, n45031, n45032, n45034, n45035, n45036,
         n45037, n45038, n45039, n45040, n45041, n45042, n45043, n45044,
         n45045, n45046, n45047, n45048, n45049, n45050, n45051, n45052,
         n45053, n45054, n45055, n45056, n45057, n45058, n45059, n45060,
         n45061, n45062, n45063, n45064, n45065, n45066, n45067, n45068,
         n45069, n45070, n45071, n45072, n45073, n45075, n45076, n45077,
         n45078, n45079, n45080, n45081, n45082, n45083, n45084, n45085,
         n45086, n45087, n45088, n45089, n45090, n45091, n45092, n45093,
         n45094, n45095, n45096, n45097, n45098, n45099, n45100, n45101,
         n45102, n45103, n45104, n45105, n45106, n45107, n45108, n45109,
         n45110, n45111, n45112, n45113, n45114, n45115, n45116, n45117,
         n45118, n45119, n45120, n45121, n45122, n45123, n45124, n45125,
         n45126, n45127, n45128, n45129, n45130, n45131, n45132, n45133,
         n45134, n45135, n45136, n45137, n45138, n45139, n45140, n45141,
         n45142, n45143, n45144, n45145, n45146, n45147, n45148, n45149,
         n45150, n45151, n45152, n45153, n45156, n45157, n45158, n45159,
         n45160, n45161, n45162, n45163, n45164, n45165, n45166, n45167,
         n45168, n45169, n45170, n45171, n45172, n45173, n45174, n45175,
         n45176, n45177, n45178, n45179, n45180, n45181, n45182, n45183,
         n45184, n45185, n45186, n45187, n45188, n45189, n45190, n45191,
         n45192, n45193, n45194, n45195, n45196, n45197, n45198, n45199,
         n45200, n45201, n45202, n45203, n45204, n45205, n45206, n45207,
         n45208, n45209, n45210, n45211, n45212, n45213, n45214, n45215,
         n45216, n45217, n45218, n45219, n45220, n45221, n45222, n45223,
         n45224, n45225, n45226, n45227, n45228, n45229, n45230, n45231,
         n45232, n45233, n45234, n45235, n45236, n45237, n45238, n45239,
         n45240, n45241, n45242, n45243, n45244, n45245, n45246, n45247,
         n45248, n45249, n45250, n45251, n45252, n45253, n45254, n45255,
         n45256, n45257, n45258, n45259, n45260, n45261, n45262, n45263,
         n45264, n45265, n45266, n45267, n45268, n45269, n45270, n45271,
         n45272, n45273, n45274, n45275, n45276, n45277, n45278, n45279,
         n45280, n45281, n45282, n45283, n45284, n45285, n45286, n45287,
         n45288, n45289, n45290, n45291, n45293, n45294, n45295, n45296,
         n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304,
         n45305, n45306, n45307, n45308, n45309, n45310, n45311, n45312,
         n45313, n45314, n45315, n45316, n45317, n45318, n45319, n45320,
         n45321, n45322, n45323, n45324, n45325, n45326, n45327, n45328,
         n45329, n45330, n45331, n45332, n45333, n45334, n45335, n45336,
         n45337, n45338, n45339, n45340, n45341, n45342, n45343, n45344,
         n45345, n45346, n45347, n45348, n45349, n45350, n45351, n45352,
         n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360,
         n45361, n45362, n45363, n45365, n45366, n45367, n45368, n45369,
         n45370, n45371, n45372, n45373, n45374, n45375, n45376, n45377,
         n45378, n45379, n45380, n45381, n45382, n45383, n45384, n45385,
         n45386, n45387, n45388, n45389, n45390, n45391, n45392, n45393,
         n45394, n45395, n45396, n45397, n45398, n45399, n45400, n45401,
         n45402, n45403, n45404, n45405, n45406, n45407, n45408, n45409,
         n45410, n45411, n45412, n45413, n45414, n45415, n45416, n45417,
         n45418, n45419, n45420, n45421, n45422, n45423, n45424, n45425,
         n45426, n45427, n45428, n45429, n45430, n45431, n45432, n45433,
         n45434, n45435, n45436, n45437, n45438, n45439, n45440, n45441,
         n45442, n45443, n45444, n45445, n45446, n45447, n45448, n45449,
         n45450, n45451, n45452, n45453, n45454, n45455, n45456, n45457,
         n45458, n45459, n45460, n45461, n45462, n45463, n45464, n45465,
         n45466, n45467, n45468, n45469, n45470, n45471, n45472, n45473,
         n45474, n45475, n45476, n45477, n45478, n45479, n45480, n45481,
         n45482, n45483, n45484, n45485, n45486, n45487, n45488, n45489,
         n45490, n45491, n45492, n45493, n45494, n45495, n45496, n45497,
         n45498, n45499, n45500, n45501, n45502, n45503, n45504, n45505,
         n45506, n45507, n45509, n45510, n45511, n45512, n45513, n45514,
         n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522,
         n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530,
         n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538,
         n45539, n45540, n45541, n45542, n45543, n45544, n45545, n45546,
         n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554,
         n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562,
         n45563, n45564, n45565, n45566, n45567, n45568, n45569, n45570,
         n45571, n45572, n45573, n45574, n45575, n45576, n45577, n45578,
         n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586,
         n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594,
         n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602,
         n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610,
         n45611, n45612, n45613, n45614, n45615, n45616, n45617, n45618,
         n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626,
         n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634,
         n45635, n45636, n45637, n45638, n45639, n45640, n45641, n45642,
         n45643, n45644, n45645, n45646, n45647, n45648, n45649, n45650,
         n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658,
         n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666,
         n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674,
         n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682,
         n45683, n45684, n45685, n45686, n45687, n45688, n45689, n45690,
         n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698,
         n45700, n45701, n45702, n45703, n45704, n45706, n45707, n45708,
         n45709, n45710, n45711, n45712, n45713, n45714, n45715, n45716,
         n45717, n45718, n45719, n45720, n45722, n45723, n45724, n45725,
         n45726, n45727, n45728, n45729, n45730, n45731, n45732, n45733,
         n45734, n45735, n45736, n45737, n45739, n45740, n45741, n45742,
         n45743, n45744, n45745, n45746, n45747, n45748, n45749, n45750,
         n45751, n45752, n45753, n45754, n45755, n45756, n45757, n45758,
         n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766,
         n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774,
         n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782,
         n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790,
         n45791, n45792, n45793, n45794, n45795, n45796, n45797, n45798,
         n45799, n45800, n45801, n45802, n45804, n45805, n45806, n45807,
         n45808, n45809, n45810, n45811, n45812, n45813, n45814, n45815,
         n45816, n45817, n45818, n45819, n45820, n45821, n45822, n45823,
         n45824, n45825, n45826, n45827, n45828, n45829, n45830, n45831,
         n45832, n45833, n45834, n45835, n45836, n45837, n45838, n45839,
         n45840, n45841, n45842, n45843, n45844, n45845, n45847, n45848,
         n45849, n45850, n45851, n45852, n45853, n45854, n45855, n45856,
         n45857, n45858, n45859, n45860, n45861, n45862, n45863, n45864,
         n45865, n45866, n45868, n45869, n45870, n45871, n45872, n45873,
         n45874, n45875, n45876, n45877, n45878, n45880, n45881, n45882,
         n45883, n45884, n45886, n45887, n45888, n45889, n45890, n45891,
         n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899,
         n45900, n45901, n45902, n45904, n45905, n45906, n45907, n45908,
         n45909, n45910, n45911, n45912, n45913, n45914, n45915, n45916,
         n45917, n45918, n45919, n45920, n45921, n45922, n45923, n45924,
         n45925, n45926, n45927, n45928, n45929, n45930, n45931, n45932,
         n45933, n45934, n45935, n45936, n45937, n45938, n45939, n45940,
         n45941, n45942, n45943, n45944, n45945, n45946, n45947, n45948,
         n45949, n45950, n45951, n45952, n45953, n45954, n45955, n45956,
         n45957, n45958, n45959, n45960, n45961, n45962, n45963, n45964,
         n45965, n45966, n45967, n45968, n45969, n45970, n45971, n45972,
         n45973, n45974, n45975, n45976, n45977, n45978, n45979, n45980,
         n45981, n45982, n45983, n45984, n45985, n45986, n45987, n45988,
         n45989, n45990, n45991, n45992, n45993, n45994, n45995, n45996,
         n45997, n45998, n45999, n46000, n46001, n46002, n46003, n46004,
         n46005, n46006, n46007, n46008, n46009, n46010, n46011, n46012,
         n46013, n46014, n46015, n46016, n46017, n46018, n46020, n46021,
         n46022, n46023, n46024, n46025, n46026, n46027, n46028, n46029,
         n46030, n46031, n46032, n46033, n46034, n46035, n46036, n46037,
         n46038, n46039, n46040, n46041, n46042, n46043, n46044, n46045,
         n46046, n46047, n46048, n46049, n46050, n46051, n46052, n46053,
         n46054, n46055, n46056, n46057, n46058, n46059, n46060, n46061,
         n46062, n46063, n46064, n46065, n46066, n46067, n46068, n46069,
         n46070, n46071, n46072, n46073, n46074, n46075, n46076, n46077,
         n46078, n46079, n46080, n46081, n46082, n46083, n46084, n46085,
         n46086, n46087, n46089, n46090, n46091, n46092, n46093, n46094,
         n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102,
         n46103, n46104, n46105, n46106, n46107, n46108, n46109, n46110,
         n46111, n46112, n46113, n46114, n46115, n46116, n46117, n46118,
         n46119, n46120, n46121, n46122, n46123, n46124, n46125, n46126,
         n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46134,
         n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142,
         n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150,
         n46151, n46152, n46153, n46154, n46155, n46156, n46157, n46158,
         n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166,
         n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174,
         n46175, n46176, n46177, n46178, n46179, n46180, n46181, n46182,
         n46183, n46184, n46186, n46187, n46188, n46189, n46190, n46191,
         n46192, n46193, n46194, n46195, n46196, n46197, n46198, n46199,
         n46200, n46201, n46202, n46203, n46204, n46205, n46206, n46207,
         n46208, n46209, n46210, n46211, n46213, n46214, n46215, n46216,
         n46217, n46218, n46219, n46220, n46221, n46222, n46223, n46224,
         n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232,
         n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240,
         n46241, n46242, n46243, n46244, n46245, n46246, n46247, n46248,
         n46249, n46250, n46251, n46252, n46253, n46254, n46255, n46256,
         n46257, n46258, n46259, n46260, n46261, n46262, n46263, n46264,
         n46265, n46266, n46267, n46268, n46269, n46270, n46271, n46272,
         n46273, n46274, n46275, n46276, n46277, n46278, n46279, n46280,
         n46281, n46282, n46283, n46284, n46285, n46286, n46287, n46288,
         n46289, n46290, n46291, n46292, n46293, n46294, n46295, n46296,
         n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304,
         n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312,
         n46313, n46314, n46315, n46316, n46317, n46318, n46319, n46320,
         n46321, n46322, n46324, n46325, n46326, n46327, n46328, n46329,
         n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339,
         n46340, n46341, n46342, n46343, n46344, n46345, n46346, n46347,
         n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355,
         n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363,
         n46364, n46365, n46366, n46367, n46368, n46369, n46370, n46371,
         n46372, n46373, n46374, n46376, n46377, n46378, n46379, n46380,
         n46381, n46382, n46383, n46384, n46385, n46386, n46387, n46388,
         n46389, n46390, n46392, n46393, n46394, n46395, n46396, n46397,
         n46398, n46399, n46400, n46401, n46402, n46403, n46404, n46405,
         n46406, n46407, n46408, n46409, n46410, n46411, n46412, n46413,
         n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421,
         n46422, n46423, n46424, n46425, n46426, n46427, n46428, n46429,
         n46430, n46431, n46432, n46433, n46434, n46435, n46436, n46437,
         n46438, n46439, n46440, n46441, n46442, n46443, n46444, n46445,
         n46446, n46447, n46448, n46449, n46450, n46451, n46453, n46454,
         n46455, n46456, n46457, n46458, n46459, n46460, n46461, n46462,
         n46463, n46464, n46465, n46466, n46467, n46468, n46469, n46470,
         n46471, n46472, n46473, n46474, n46475, n46476, n46477, n46478,
         n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486,
         n46487, n46488, n46489, n46490, n46491, n46492, n46493, n46494,
         n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502,
         n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510,
         n46511, n46512, n46513, n46514, n46515, n46516, n46517, n46518,
         n46519, n46520, n46521, n46522, n46523, n46524, n46525, n46526,
         n46527, n46529, n46530, n46532, n46533, n46534, n46535, n46536,
         n46537, n46538, n46539, n46540, n46541, n46542, n46543, n46544,
         n46546, n46547, n46548, n46549, n46550, n46551, n46552, n46553,
         n46554, n46555, n46557, n46558, n46559, n46560, n46561, n46562,
         n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570,
         n46571, n46572, n46573, n46574, n46575, n46576, n46577, n46578,
         n46579, n46580, n46581, n46582, n46583, n46584, n46585, n46586,
         n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594,
         n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602,
         n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610,
         n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618,
         n46619, n46620, n46621, n46622, n46623, n46624, n46625, n46626,
         n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634,
         n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642,
         n46643, n46644, n46645, n46646, n46647, n46648, n46649, n46650,
         n46651, n46652, n46653, n46654, n46655, n46656, n46657, n46658,
         n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666,
         n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674,
         n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682,
         n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690,
         n46691, n46692, n46693, n46694, n46695, n46696, n46697, n46698,
         n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706,
         n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714,
         n46715, n46716, n46717, n46718, n46719, n46720, n46721, n46722,
         n46723, n46724, n46725, n46726, n46727, n46728, n46729, n46730,
         n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738,
         n46739, n46740, n46741, n46742, n46743, n46744, n46746, n46747,
         n46748, n46749, n46750, n46751, n46752, n46753, n46754, n46755,
         n46756, n46757, n46760, n46761, n46762, n46763, n46764, n46766,
         n46767, n46768, n46769, n46770, n46772, n46773, n46774, n46775,
         n46776, n46777, n46778, n46779, n46780, n46781, n46782, n46783,
         n46784, n46785, n46786, n46787, n46788, n46789, n46790, n46791,
         n46792, n46793, n46794, n46795, n46796, n46797, n46798, n46799,
         n46800, n46801, n46802, n46803, n46804, n46805, n46806, n46807,
         n46808, n46809, n46810, n46811, n46812, n46813, n46814, n46815,
         n46816, n46817, n46818, n46819, n46820, n46821, n46822, n46823,
         n46824, n46825, n46826, n46827, n46828, n46829, n46830, n46831,
         n46832, n46833, n46834, n46835, n46836, n46837, n46838, n46839,
         n46840, n46841, n46842, n46843, n46844, n46845, n46846, n46847,
         n46848, n46849, n46850, n46851, n46852, n46853, n46854, n46855,
         n46856, n46857, n46858, n46859, n46860, n46861, n46862, n46863,
         n46864, n46865, n46866, n46867, n46868, n46869, n46870, n46871,
         n46872, n46873, n46874, n46875, n46876, n46877, n46878, n46879,
         n46880, n46881, n46882, n46883, n46884, n46885, n46886, n46887,
         n46888, n46889, n46890, n46891, n46892, n46893, n46894, n46895,
         n46896, n46897, n46898, n46899, n46900, n46901, n46902, n46903,
         n46904, n46905, n46906, n46907, n46908, n46909, n46910, n46911,
         n46912, n46913, n46915, n46916, n46917, n46918, n46919, n46920,
         n46921, n46922, n46923, n46924, n46925, n46926, n46927, n46929,
         n46930, n46931, n46932, n46933, n46934, n46935, n46936, n46938,
         n46939, n46940, n46941, n46942, n46943, n46944, n46945, n46946,
         n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954,
         n46956, n46957, n46958, n46959, n46960, n46961, n46962, n46963,
         n46964, n46965, n46966, n46967, n46968, n46969, n46970, n46971,
         n46972, n46973, n46974, n46975, n46976, n46977, n46978, n46979,
         n46980, n46981, n46982, n46983, n46984, n46985, n46986, n46987,
         n46988, n46989, n46990, n46991, n46992, n46993, n46994, n46995,
         n46996, n46997, n46998, n46999, n47000, n47001, n47002, n47003,
         n47004, n47005, n47006, n47007, n47008, n47009, n47010, n47011,
         n47012, n47013, n47014, n47015, n47016, n47017, n47018, n47019,
         n47020, n47021, n47022, n47023, n47024, n47025, n47026, n47027,
         n47028, n47029, n47030, n47031, n47032, n47033, n47034, n47035,
         n47036, n47037, n47038, n47040, n47041, n47042, n47043, n47044,
         n47045, n47046, n47047, n47048, n47049, n47050, n47051, n47052,
         n47053, n47054, n47055, n47056, n47057, n47058, n47059, n47060,
         n47061, n47062, n47063, n47064, n47065, n47066, n47067, n47068,
         n47069, n47070, n47071, n47072, n47073, n47074, n47075, n47076,
         n47077, n47078, n47079, n47080, n47081, n47082, n47083, n47084,
         n47085, n47086, n47087, n47088, n47089, n47090, n47091, n47092,
         n47093, n47094, n47095, n47096, n47097, n47098, n47099, n47100,
         n47101, n47102, n47103, n47104, n47105, n47106, n47107, n47108,
         n47109, n47110, n47111, n47112, n47113, n47114, n47115, n47116,
         n47117, n47118, n47119, n47120, n47121, n47122, n47123, n47124,
         n47125, n47126, n47127, n47128, n47129, n47130, n47131, n47132,
         n47133, n47134, n47135, n47136, n47137, n47138, n47139, n47140,
         n47141, n47142, n47143, n47144, n47145, n47146, n47147, n47148,
         n47149, n47150, n47151, n47152, n47153, n47154, n47155, n47156,
         n47157, n47158, n47159, n47160, n47161, n47162, n47163, n47164,
         n47165, n47166, n47167, n47168, n47169, n47170, n47171, n47172,
         n47173, n47174, n47175, n47176, n47177, n47178, n47179, n47180,
         n47181, n47182, n47183, n47184, n47185, n47186, n47187, n47188,
         n47189, n47190, n47191, n47192, n47193, n47194, n47195, n47196,
         n47198, n47199, n47200, n47201, n47202, n47203, n47204, n47205,
         n47206, n47207, n47208, n47209, n47210, n47211, n47212, n47213,
         n47214, n47215, n47216, n47217, n47218, n47219, n47220, n47221,
         n47222, n47223, n47224, n47225, n47226, n47227, n47228, n47229,
         n47230, n47231, n47232, n47233, n47234, n47236, n47237, n47238,
         n47239, n47240, n47241, n47242, n47243, n47244, n47245, n47246,
         n47247, n47248, n47249, n47250, n47251, n47252, n47253, n47254,
         n47255, n47256, n47257, n47258, n47259, n47260, n47261, n47262,
         n47263, n47264, n47265, n47266, n47267, n47268, n47269, n47270,
         n47271, n47272, n47273, n47274, n47275, n47276, n47277, n47278,
         n47279, n47280, n47281, n47282, n47283, n47284, n47285, n47286,
         n47287, n47288, n47289, n47290, n47291, n47292, n47293, n47294,
         n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302,
         n47304, n47305, n47306, n47307, n47308, n47309, n47310, n47311,
         n47312, n47313, n47314, n47315, n47316, n47317, n47318, n47319,
         n47320, n47321, n47322, n47323, n47324, n47325, n47326, n47327,
         n47328, n47329, n47330, n47331, n47332, n47333, n47334, n47335,
         n47336, n47337, n47338, n47339, n47340, n47341, n47342, n47343,
         n47344, n47345, n47346, n47347, n47348, n47349, n47350, n47351,
         n47352, n47353, n47354, n47355, n47356, n47357, n47358, n47359,
         n47360, n47361, n47362, n47363, n47364, n47365, n47366, n47367,
         n47368, n47369, n47370, n47371, n47372, n47373, n47374, n47375,
         n47376, n47377, n47378, n47379, n47380, n47381, n47382, n47383,
         n47384, n47385, n47386, n47387, n47388, n47389, n47390, n47391,
         n47392, n47393, n47394, n47395, n47396, n47397, n47398, n47399,
         n47400, n47401, n47402, n47403, n47404, n47405, n47406, n47407,
         n47408, n47409, n47410, n47411, n47412, n47413, n47414, n47415,
         n47416, n47417, n47418, n47419, n47420, n47421, n47422, n47423,
         n47424, n47425, n47426, n47427, n47429, n47430, n47431, n47432,
         n47433, n47434, n47435, n47436, n47437, n47438, n47439, n47440,
         n47441, n47442, n47443, n47444, n47445, n47446, n47448, n47449,
         n47450, n47451, n47452, n47453, n47454, n47455, n47456, n47457,
         n47458, n47459, n47461, n47462, n47463, n47464, n47465, n47466,
         n47467, n47468, n47469, n47471, n47472, n47473, n47474, n47475,
         n47476, n47477, n47478, n47479, n47480, n47481, n47482, n47483,
         n47484, n47485, n47486, n47487, n47488, n47489, n47490, n47491,
         n47492, n47493, n47494, n47495, n47496, n47497, n47498, n47499,
         n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507,
         n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515,
         n47516, n47517, n47518, n47519, n47520, n47521, n47522, n47523,
         n47524, n47525, n47526, n47527, n47528, n47530, n47532, n47533,
         n47534, n47535, n47536, n47537, n47538, n47539, n47540, n47541,
         n47542, n47543, n47544, n47545, n47546, n47547, n47548, n47549,
         n47550, n47551, n47552, n47553, n47554, n47555, n47556, n47557,
         n47558, n47559, n47560, n47561, n47563, n47564, n47565, n47566,
         n47567, n47568, n47569, n47570, n47571, n47572, n47573, n47574,
         n47575, n47576, n47577, n47578, n47579, n47580, n47581, n47582,
         n47583, n47584, n47586, n47587, n47588, n47589, n47590, n47591,
         n47592, n47593, n47594, n47595, n47596, n47598, n47599, n47600,
         n47601, n47602, n47603, n47604, n47605, n47606, n47607, n47608,
         n47609, n47610, n47612, n47613, n47614, n47615, n47616, n47617,
         n47618, n47619, n47620, n47621, n47622, n47623, n47624, n47625,
         n47626, n47627, n47628, n47629, n47630, n47631, n47632, n47633,
         n47634, n47635, n47636, n47637, n47638, n47639, n47640, n47641,
         n47642, n47643, n47644, n47645, n47646, n47647, n47648, n47649,
         n47650, n47651, n47652, n47653, n47654, n47655, n47656, n47657,
         n47658, n47659, n47660, n47661, n47662, n47663, n47664, n47665,
         n47666, n47667, n47668, n47669, n47670, n47671, n47672, n47673,
         n47674, n47675, n47676, n47677, n47678, n47679, n47680, n47681,
         n47682, n47683, n47684, n47685, n47686, n47687, n47688, n47689,
         n47690, n47691, n47692, n47693, n47694, n47695, n47696, n47697,
         n47698, n47699, n47700, n47701, n47702, n47703, n47704, n47705,
         n47706, n47707, n47708, n47710, n47711, n47712, n47713, n47714,
         n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722,
         n47723, n47724, n47725, n47727, n47728, n47729, n47730, n47731,
         n47732, n47733, n47734, n47735, n47736, n47737, n47738, n47739,
         n47740, n47741, n47742, n47743, n47744, n47745, n47746, n47747,
         n47748, n47749, n47750, n47751, n47752, n47753, n47754, n47755,
         n47756, n47757, n47758, n47759, n47760, n47761, n47762, n47763,
         n47764, n47765, n47766, n47767, n47768, n47769, n47770, n47771,
         n47772, n47773, n47774, n47775, n47776, n47777, n47778, n47779,
         n47780, n47781, n47782, n47783, n47784, n47785, n47786, n47787,
         n47788, n47789, n47790, n47791, n47792, n47793, n47794, n47795,
         n47796, n47797, n47798, n47799, n47800, n47801, n47802, n47803,
         n47804, n47805, n47806, n47807, n47808, n47809, n47810, n47811,
         n47812, n47813, n47814, n47816, n47817, n47818, n47819, n47820,
         n47821, n47822, n47823, n47824, n47825, n47826, n47827, n47828,
         n47831, n47832, n47833, n47834, n47835, n47836, n47837, n47838,
         n47839, n47840, n47841, n47842, n47843, n47844, n47845, n47846,
         n47847, n47848, n47849, n47850, n47851, n47852, n47853, n47854,
         n47855, n47856, n47857, n47858, n47859, n47860, n47861, n47862,
         n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870,
         n47871, n47872, n47873, n47874, n47875, n47876, n47877, n47878,
         n47879, n47880, n47881, n47882, n47883, n47884, n47885, n47886,
         n47887, n47888, n47889, n47890, n47891, n47892, n47893, n47894,
         n47895, n47896, n47897, n47898, n47899, n47900, n47901, n47902,
         n47903, n47905, n47906, n47907, n47908, n47909, n47910, n47911,
         n47912, n47913, n47914, n47915, n47916, n47917, n47918, n47919,
         n47920, n47921, n47922, n47923, n47924, n47925, n47926, n47927,
         n47928, n47930, n47931, n47932, n47934, n47935, n47936, n47937,
         n47938, n47939, n47940, n47941, n47942, n47943, n47944, n47945,
         n47946, n47947, n47948, n47949, n47950, n47951, n47952, n47953,
         n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962,
         n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970,
         n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978,
         n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986,
         n47987, n47988, n47989, n47990, n47991, n47992, n47994, n47995,
         n47996, n47997, n47998, n47999, n48000, n48001, n48002, n48003,
         n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011,
         n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019,
         n48020, n48021, n48022, n48023, n48024, n48025, n48026, n48027,
         n48028, n48029, n48030, n48031, n48032, n48033, n48034, n48035,
         n48036, n48037, n48038, n48039, n48040, n48041, n48042, n48043,
         n48044, n48045, n48046, n48047, n48048, n48049, n48050, n48051,
         n48052, n48053, n48054, n48055, n48056, n48058, n48059, n48060,
         n48061, n48062, n48063, n48064, n48065, n48066, n48067, n48068,
         n48069, n48070, n48071, n48072, n48073, n48074, n48075, n48076,
         n48077, n48078, n48079, n48080, n48081, n48082, n48083, n48084,
         n48085, n48086, n48087, n48088, n48089, n48090, n48091, n48093,
         n48094, n48095, n48096, n48097, n48098, n48099, n48100, n48101,
         n48102, n48103, n48104, n48105, n48106, n48107, n48108, n48110,
         n48111, n48112, n48113, n48114, n48115, n48116, n48117, n48118,
         n48119, n48120, n48121, n48122, n48123, n48124, n48125, n48126,
         n48127, n48128, n48129, n48130, n48131, n48132, n48133, n48134,
         n48135, n48136, n48137, n48138, n48139, n48140, n48141, n48142,
         n48143, n48144, n48145, n48146, n48147, n48148, n48149, n48150,
         n48151, n48152, n48153, n48154, n48155, n48156, n48157, n48158,
         n48159, n48160, n48161, n48162, n48163, n48164, n48165, n48166,
         n48167, n48168, n48169, n48170, n48171, n48172, n48173, n48174,
         n48175, n48176, n48177, n48178, n48179, n48180, n48181, n48182,
         n48183, n48184, n48185, n48186, n48187, n48188, n48189, n48190,
         n48191, n48192, n48193, n48194, n48195, n48196, n48197, n48198,
         n48199, n48200, n48201, n48203, n48204, n48205, n48206, n48207,
         n48208, n48209, n48210, n48211, n48212, n48213, n48214, n48215,
         n48216, n48217, n48218, n48219, n48220, n48221, n48222, n48223,
         n48224, n48225, n48226, n48227, n48228, n48229, n48230, n48231,
         n48232, n48233, n48234, n48236, n48237, n48238, n48239, n48240,
         n48241, n48242, n48243, n48244, n48246, n48247, n48248, n48249,
         n48250, n48251, n48252, n48253, n48254, n48255, n48256, n48257,
         n48258, n48259, n48260, n48261, n48262, n48263, n48264, n48265,
         n48266, n48267, n48268, n48269, n48270, n48271, n48272, n48273,
         n48274, n48275, n48276, n48277, n48278, n48279, n48280, n48281,
         n48282, n48283, n48284, n48285, n48286, n48287, n48288, n48289,
         n48290, n48291, n48292, n48293, n48294, n48295, n48296, n48297,
         n48298, n48299, n48300, n48301, n48302, n48303, n48304, n48305,
         n48306, n48307, n48308, n48309, n48310, n48311, n48312, n48313,
         n48314, n48315, n48316, n48317, n48318, n48319, n48320, n48321,
         n48322, n48323, n48324, n48325, n48326, n48327, n48328, n48329,
         n48330, n48331, n48332, n48333, n48334, n48335, n48336, n48337,
         n48338, n48339, n48340, n48341, n48342, n48343, n48344, n48345,
         n48346, n48347, n48348, n48349, n48350, n48351, n48352, n48353,
         n48354, n48355, n48356, n48357, n48358, n48359, n48360, n48361,
         n48362, n48363, n48364, n48365, n48366, n48367, n48368, n48369,
         n48370, n48371, n48372, n48373, n48374, n48375, n48376, n48377,
         n48378, n48379, n48380, n48381, n48382, n48386, n48387, n48388,
         n48389, n48390, n48391, n48392, n48393, n48394, n48395, n48396,
         n48397, n48398, n48399, n48400, n48401, n48402, n48403, n48404,
         n48405, n48406, n48407, n48408, n48409, n48410, n48411, n48412,
         n48413, n48414, n48415, n48416, n48417, n48418, n48419, n48420,
         n48421, n48422, n48423, n48424, n48425, n48426, n48427, n48428,
         n48429, n48430, n48431, n48432, n48433, n48434, n48435, n48436,
         n48437, n48438, n48439, n48441, n48442, n48443, n48444, n48445,
         n48446, n48447, n48448, n48449, n48450, n48451, n48452, n48453,
         n48454, n48455, n48456, n48457, n48458, n48459, n48460, n48461,
         n48462, n48463, n48464, n48465, n48466, n48467, n48468, n48469,
         n48470, n48471, n48472, n48473, n48474, n48475, n48476, n48477,
         n48478, n48479, n48480, n48481, n48482, n48483, n48484, n48485,
         n48486, n48487, n48488, n48489, n48490, n48491, n48492, n48493,
         n48494, n48495, n48496, n48497, n48498, n48499, n48500, n48501,
         n48502, n48503, n48504, n48505, n48506, n48507, n48508, n48509,
         n48510, n48512, n48513, n48514, n48515, n48516, n48517, n48518,
         n48519, n48520, n48521, n48522, n48523, n48524, n48525, n48526,
         n48527, n48528, n48529, n48530, n48531, n48532, n48533, n48534,
         n48535, n48536, n48537, n48538, n48539, n48540, n48541, n48542,
         n48543, n48544, n48545, n48546, n48547, n48548, n48549, n48550,
         n48551, n48552, n48553, n48554, n48555, n48556, n48557, n48558,
         n48559, n48560, n48561, n48562, n48563, n48564, n48565, n48566,
         n48567, n48568, n48569, n48570, n48571, n48572, n48573, n48574,
         n48575, n48576, n48577, n48578, n48579, n48580, n48581, n48582,
         n48583, n48584, n48585, n48586, n48587, n48588, n48589, n48590,
         n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598,
         n48599, n48600, n48602, n48603, n48604, n48605, n48606, n48607,
         n48608, n48609, n48610, n48611, n48612, n48613, n48614, n48615,
         n48616, n48617, n48618, n48620, n48621, n48622, n48623, n48624,
         n48625, n48626, n48627, n48628, n48629, n48630, n48631, n48632,
         n48633, n48635, n48636, n48638, n48639, n48640, n48641, n48642,
         n48643, n48644, n48646, n48647, n48648, n48649, n48650, n48651,
         n48652, n48653, n48654, n48655, n48656, n48657, n48658, n48659,
         n48661, n48662, n48663, n48664, n48665, n48666, n48667, n48668,
         n48669, n48670, n48671, n48672, n48674, n48675, n48676, n48677,
         n48678, n48679, n48682, n48683, n48684, n48685, n48686, n48687,
         n48688, n48689, n48690, n48691, n48692, n48694, n48695, n48696,
         n48697, n48698, n48699, n48700, n48701, n48702, n48703, n48704,
         n48705, n48706, n48707, n48708, n48709, n48710, n48711, n48712,
         n48713, n48714, n48715, n48716, n48717, n48718, n48719, n48720,
         n48721, n48722, n48723, n48724, n48725, n48726, n48727, n48728,
         n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736,
         n48737, n48738, n48739, n48740, n48741, n48742, n48743, n48744,
         n48745, n48747, n48748, n48749, n48750, n48751, n48752, n48753,
         n48754, n48755, n48756, n48757, n48759, n48760, n48762, n48763,
         n48764, n48765, n48766, n48767, n48768, n48769, n48770, n48771,
         n48772, n48773, n48774, n48775, n48776, n48777, n48778, n48779,
         n48780, n48781, n48782, n48783, n48784, n48785, n48786, n48787,
         n48788, n48789, n48790, n48791, n48792, n48793, n48794, n48795,
         n48796, n48797, n48798, n48799, n48800, n48801, n48802, n48803,
         n48804, n48805, n48806, n48807, n48808, n48809, n48810, n48811,
         n48812, n48813, n48814, n48815, n48816, n48817, n48818, n48819,
         n48820, n48821, n48823, n48824, n48825, n48826, n48827, n48828,
         n48829, n48830, n48831, n48832, n48833, n48834, n48835, n48836,
         n48837, n48838, n48839, n48840, n48841, n48842, n48843, n48844,
         n48845, n48846, n48847, n48848, n48849, n48850, n48851, n48852,
         n48853, n48854, n48855, n48856, n48857, n48858, n48859, n48860,
         n48861, n48862, n48863, n48864, n48865, n48866, n48867, n48868,
         n48869, n48870, n48871, n48872, n48873, n48874, n48875, n48876,
         n48877, n48878, n48879, n48880, n48881, n48882, n48883, n48884,
         n48885, n48886, n48887, n48888, n48889, n48890, n48891, n48892,
         n48893, n48894, n48895, n48896, n48897, n48898, n48899, n48900,
         n48901, n48902, n48903, n48904, n48905, n48906, n48907, n48908,
         n48909, n48910, n48911, n48912, n48913, n48914, n48915, n48916,
         n48917, n48918, n48919, n48920, n48921, n48922, n48923, n48924,
         n48925, n48926, n48927, n48928, n48929, n48930, n48931, n48932,
         n48933, n48934, n48935, n48936, n48937, n48938, n48939, n48940,
         n48941, n48942, n48943, n48944, n48945, n48946, n48947, n48948,
         n48949, n48950, n48951, n48952, n48953, n48954, n48955, n48956,
         n48957, n48958, n48959, n48960, n48961, n48962, n48963, n48964,
         n48965, n48966, n48967, n48968, n48969, n48970, n48971, n48972,
         n48973, n48974, n48975, n48976, n48977, n48978, n48979, n48980,
         n48981, n48982, n48983, n48984, n48985, n48986, n48987, n48988,
         n48989, n48990, n48991, n48992, n48993, n48994, n48995, n48996,
         n48997, n48998, n48999, n49000, n49001, n49002, n49003, n49004,
         n49005, n49006, n49007, n49008, n49009, n49010, n49011, n49012,
         n49013, n49014, n49015, n49016, n49017, n49018, n49019, n49020,
         n49021, n49022, n49023, n49024, n49025, n49026, n49027, n49029,
         n49030, n49031, n49032, n49034, n49035, n49036, n49037, n49038,
         n49039, n49040, n49041, n49042, n49043, n49044, n49045, n49046,
         n49047, n49048, n49049, n49050, n49051, n49052, n49053, n49054,
         n49055, n49056, n49057, n49058, n49059, n49060, n49061, n49062,
         n49063, n49065, n49066, n49067, n49068, n49069, n49070, n49071,
         n49072, n49073, n49074, n49075, n49076, n49077, n49078, n49079,
         n49080, n49081, n49082, n49083, n49084, n49085, n49086, n49087,
         n49088, n49089, n49090, n49091, n49092, n49093, n49094, n49095,
         n49096, n49097, n49098, n49099, n49100, n49101, n49102, n49103,
         n49104, n49105, n49106, n49107, n49108, n49109, n49110, n49111,
         n49112, n49113, n49114, n49115, n49116, n49117, n49118, n49119,
         n49120, n49122, n49123, n49124, n49125, n49126, n49127, n49128,
         n49129, n49130, n49131, n49132, n49133, n49134, n49135, n49136,
         n49137, n49138, n49139, n49140, n49141, n49142, n49143, n49144,
         n49145, n49146, n49147, n49148, n49149, n49150, n49151, n49152,
         n49153, n49154, n49155, n49156, n49157, n49158, n49159, n49160,
         n49161, n49162, n49163, n49164, n49165, n49166, n49167, n49168,
         n49169, n49170, n49171, n49172, n49173, n49174, n49175, n49176,
         n49177, n49178, n49179, n49180, n49181, n49182, n49183, n49184,
         n49185, n49186, n49187, n49188, n49189, n49190, n49191, n49192,
         n49193, n49194, n49195, n49196, n49197, n49198, n49199, n49200,
         n49201, n49202, n49203, n49204, n49205, n49207, n49208, n49209,
         n49210, n49211, n49212, n49213, n49214, n49215, n49216, n49217,
         n49218, n49220, n49221, n49222, n49223, n49224, n49225, n49226,
         n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49235,
         n49236, n49237, n49238, n49240, n49241, n49242, n49243, n49244,
         n49245, n49246, n49247, n49248, n49249, n49250, n49251, n49252,
         n49253, n49254, n49255, n49256, n49257, n49258, n49259, n49260,
         n49261, n49262, n49263, n49264, n49265, n49266, n49267, n49268,
         n49269, n49270, n49271, n49272, n49273, n49274, n49275, n49276,
         n49277, n49278, n49279, n49280, n49281, n49282, n49283, n49284,
         n49285, n49286, n49287, n49288, n49289, n49290, n49291, n49292,
         n49293, n49294, n49295, n49296, n49297, n49298, n49299, n49300,
         n49301, n49302, n49303, n49304, n49305, n49306, n49307, n49308,
         n49309, n49310, n49311, n49312, n49313, n49314, n49315, n49316,
         n49317, n49318, n49319, n49320, n49321, n49322, n49323, n49324,
         n49325, n49326, n49327, n49328, n49329, n49330, n49331, n49332,
         n49333, n49334, n49335, n49336, n49337, n49338, n49339, n49340,
         n49341, n49342, n49343, n49344, n49345, n49346, n49347, n49348,
         n49349, n49350, n49351, n49352, n49353, n49354, n49356, n49357,
         n49358, n49359, n49360, n49361, n49362, n49363, n49364, n49365,
         n49366, n49367, n49368, n49369, n49370, n49371, n49372, n49373,
         n49374, n49375, n49376, n49377, n49378, n49379, n49380, n49381,
         n49382, n49383, n49384, n49385, n49386, n49387, n49389, n49390,
         n49391, n49392, n49393, n49394, n49395, n49396, n49397, n49398,
         n49399, n49400, n49402, n49403, n49404, n49405, n49406, n49407,
         n49408, n49409, n49410, n49411, n49412, n49413, n49414, n49415,
         n49416, n49417, n49418, n49419, n49420, n49421, n49422, n49423,
         n49424, n49425, n49426, n49427, n49428, n49429, n49430, n49431,
         n49432, n49433, n49434, n49435, n49436, n49437, n49439, n49440,
         n49441, n49442, n49443, n49444, n49445, n49446, n49448, n49449,
         n49450, n49451, n49452, n49453, n49454, n49455, n49456, n49457,
         n49458, n49459, n49460, n49461, n49462, n49463, n49464, n49465,
         n49466, n49467, n49468, n49469, n49470, n49471, n49472, n49473,
         n49474, n49475, n49476, n49477, n49478, n49479, n49480, n49481,
         n49482, n49483, n49484, n49485, n49486, n49487, n49488, n49489,
         n49490, n49491, n49492, n49493, n49494, n49495, n49496, n49497,
         n49498, n49499, n49500, n49501, n49502, n49503, n49504, n49505,
         n49506, n49507, n49508, n49509, n49510, n49511, n49512, n49514,
         n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522,
         n49523, n49524, n49525, n49526, n49528, n49529, n49530, n49531,
         n49532, n49533, n49534, n49536, n49537, n49538, n49539, n49540,
         n49541, n49542, n49543, n49544, n49545, n49546, n49547, n49548,
         n49549, n49551, n49552, n49553, n49554, n49555, n49556, n49557,
         n49558, n49559, n49560, n49561, n49562, n49563, n49564, n49565,
         n49566, n49567, n49568, n49569, n49570, n49571, n49572, n49573,
         n49574, n49575, n49576, n49577, n49578, n49579, n49580, n49581,
         n49582, n49583, n49584, n49585, n49586, n49587, n49588, n49589,
         n49590, n49591, n49592, n49593, n49594, n49595, n49596, n49597,
         n49598, n49599, n49600, n49601, n49602, n49603, n49604, n49605,
         n49606, n49607, n49608, n49609, n49610, n49611, n49612, n49613,
         n49614, n49615, n49616, n49617, n49618, n49619, n49620, n49621,
         n49622, n49623, n49624, n49625, n49626, n49627, n49628, n49629,
         n49630, n49631, n49632, n49633, n49634, n49635, n49636, n49637,
         n49638, n49639, n49640, n49641, n49642, n49643, n49644, n49645,
         n49646, n49647, n49648, n49649, n49650, n49651, n49652, n49653,
         n49654, n49655, n49656, n49657, n49658, n49659, n49660, n49661,
         n49662, n49663, n49664, n49665, n49666, n49667, n49668, n49669,
         n49671, n49672, n49673, n49674, n49675, n49676, n49677, n49678,
         n49679, n49680, n49681, n49682, n49683, n49684, n49685, n49686,
         n49687, n49688, n49689, n49690, n49691, n49692, n49693, n49694,
         n49695, n49696, n49698, n49699, n49700, n49701, n49702, n49703,
         n49704, n49705, n49706, n49707, n49708, n49709, n49710, n49711,
         n49712, n49713, n49714, n49715, n49716, n49717, n49718, n49719,
         n49720, n49721, n49722, n49723, n49724, n49725, n49726, n49727,
         n49728, n49729, n49730, n49731, n49732, n49733, n49734, n49735,
         n49736, n49737, n49738, n49739, n49740, n49742, n49743, n49744,
         n49745, n49746, n49747, n49748, n49749, n49750, n49751, n49752,
         n49753, n49754, n49755, n49756, n49757, n49758, n49759, n49760,
         n49761, n49762, n49763, n49764, n49765, n49766, n49767, n49768,
         n49769, n49770, n49771, n49772, n49773, n49774, n49775, n49776,
         n49777, n49778, n49779, n49780, n49781, n49782, n49783, n49784,
         n49785, n49786, n49787, n49788, n49789, n49790, n49791, n49792,
         n49793, n49794, n49795, n49796, n49797, n49798, n49799, n49800,
         n49801, n49802, n49803, n49804, n49805, n49806, n49807, n49808,
         n49809, n49810, n49811, n49812, n49813, n49814, n49815, n49816,
         n49817, n49818, n49819, n49820, n49821, n49822, n49823, n49824,
         n49825, n49826, n49827, n49828, n49829, n49830, n49831, n49832,
         n49833, n49834, n49835, n49836, n49837, n49839, n49840, n49841,
         n49842, n49843, n49844, n49845, n49846, n49847, n49848, n49849,
         n49850, n49851, n49852, n49853, n49854, n49855, n49856, n49857,
         n49858, n49859, n49860, n49861, n49862, n49863, n49864, n49865,
         n49866, n49867, n49868, n49869, n49870, n49871, n49872, n49873,
         n49874, n49875, n49876, n49877, n49878, n49879, n49880, n49881,
         n49882, n49883, n49884, n49885, n49886, n49887, n49888, n49889,
         n49890, n49891, n49892, n49893, n49894, n49895, n49896, n49897,
         n49898, n49899, n49900, n49901, n49902, n49903, n49904, n49905,
         n49906, n49907, n49908, n49909, n49910, n49911, n49912, n49913,
         n49914, n49915, n49916, n49917, n49918, n49919, n49920, n49923,
         n49924, n49925, n49926, n49927, n49928, n49929, n49930, n49931,
         n49932, n49933, n49934, n49935, n49936, n49937, n49938, n49939,
         n49940, n49941, n49942, n49944, n49945, n49946, n49947, n49948,
         n49949, n49950, n49951, n49952, n49953, n49954, n49955, n49956,
         n49957, n49958, n49959, n49960, n49961, n49962, n49963, n49964,
         n49965, n49966, n49967, n49968, n49969, n49970, n49971, n49972,
         n49973, n49975, n49976, n49977, n49978, n49979, n49980, n49981,
         n49982, n49983, n49984, n49985, n49986, n49987, n49988, n49989,
         n49990, n49991, n49992, n49993, n49994, n49995, n49996, n49997,
         n49998, n49999, n50000, n50001, n50002, n50003, n50005, n50006,
         n50007, n50008, n50009, n50010, n50011, n50012, n50013, n50014,
         n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022,
         n50023, n50024, n50025, n50026, n50027, n50028, n50029, n50030,
         n50031, n50032, n50033, n50034, n50035, n50036, n50037, n50038,
         n50039, n50040, n50041, n50042, n50043, n50044, n50045, n50047,
         n50048, n50049, n50050, n50051, n50052, n50053, n50054, n50055,
         n50056, n50057, n50058, n50059, n50060, n50061, n50062, n50063,
         n50064, n50065, n50066, n50067, n50068, n50069, n50070, n50071,
         n50072, n50073, n50074, n50075, n50076, n50077, n50078, n50079,
         n50080, n50081, n50082, n50083, n50084, n50085, n50086, n50087,
         n50088, n50089, n50090, n50091, n50092, n50093, n50094, n50095,
         n50096, n50097, n50098, n50099, n50100, n50101, n50102, n50103,
         n50104, n50105, n50106, n50107, n50110, n50111, n50112, n50113,
         n50114, n50115, n50116, n50118, n50119, n50120, n50121, n50122,
         n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130,
         n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138,
         n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146,
         n50147, n50148, n50149, n50150, n50151, n50152, n50153, n50154,
         n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162,
         n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170,
         n50172, n50173, n50175, n50176, n50177, n50178, n50179, n50180,
         n50181, n50182, n50183, n50184, n50185, n50186, n50187, n50188,
         n50189, n50191, n50192, n50193, n50194, n50195, n50196, n50197,
         n50198, n50199, n50200, n50201, n50202, n50203, n50204, n50205,
         n50206, n50207, n50208, n50209, n50210, n50211, n50212, n50213,
         n50214, n50215, n50216, n50217, n50218, n50219, n50220, n50222,
         n50223, n50224, n50225, n50226, n50227, n50228, n50229, n50230,
         n50231, n50232, n50233, n50234, n50235, n50236, n50237, n50238,
         n50239, n50240, n50241, n50242, n50243, n50244, n50245, n50246,
         n50247, n50248, n50249, n50250, n50251, n50252, n50253, n50254,
         n50255, n50256, n50257, n50258, n50259, n50260, n50261, n50262,
         n50263, n50264, n50265, n50266, n50267, n50268, n50269, n50270,
         n50271, n50272, n50273, n50274, n50275, n50276, n50277, n50278,
         n50279, n50280, n50281, n50282, n50283, n50284, n50285, n50286,
         n50287, n50288, n50289, n50290, n50291, n50292, n50293, n50294,
         n50295, n50296, n50297, n50299, n50300, n50301, n50302, n50303,
         n50304, n50305, n50306, n50307, n50308, n50309, n50310, n50311,
         n50312, n50313, n50314, n50315, n50316, n50317, n50318, n50319,
         n50320, n50321, n50322, n50323, n50324, n50325, n50326, n50327,
         n50328, n50329, n50330, n50331, n50332, n50333, n50334, n50335,
         n50336, n50337, n50338, n50339, n50340, n50341, n50342, n50343,
         n50344, n50345, n50346, n50347, n50348, n50349, n50350, n50351,
         n50352, n50353, n50354, n50355, n50356, n50357, n50358, n50359,
         n50360, n50361, n50362, n50363, n50364, n50365, n50366, n50367,
         n50368, n50369, n50370, n50371, n50372, n50373, n50374, n50375,
         n50376, n50377, n50378, n50379, n50380, n50381, n50382, n50383,
         n50384, n50385, n50386, n50387, n50388, n50389, n50390, n50391,
         n50392, n50393, n50394, n50395, n50396, n50397, n50398, n50399,
         n50400, n50401, n50402, n50403, n50404, n50405, n50406, n50407,
         n50408, n50409, n50410, n50411, n50412, n50413, n50414, n50415,
         n50416, n50417, n50418, n50419, n50420, n50421, n50422, n50423,
         n50424, n50425, n50426, n50427, n50428, n50429, n50430, n50431,
         n50433, n50434, n50435, n50436, n50437, n50438, n50439, n50440,
         n50441, n50442, n50443, n50444, n50445, n50446, n50447, n50448,
         n50449, n50450, n50451, n50452, n50453, n50454, n50455, n50456,
         n50457, n50458, n50459, n50460, n50461, n50462, n50463, n50465,
         n50466, n50467, n50468, n50469, n50470, n50471, n50472, n50473,
         n50474, n50475, n50476, n50477, n50478, n50479, n50480, n50481,
         n50482, n50483, n50484, n50485, n50486, n50487, n50488, n50489,
         n50490, n50491, n50492, n50493, n50494, n50495, n50496, n50497,
         n50500, n50501, n50502, n50503, n50504, n50505, n50506, n50507,
         n50508, n50509, n50510, n50511, n50512, n50513, n50514, n50515,
         n50516, n50517, n50518, n50519, n50520, n50521, n50522, n50523,
         n50524, n50525, n50526, n50527, n50528, n50529, n50530, n50531,
         n50532, n50533, n50534, n50535, n50536, n50537, n50538, n50539,
         n50540, n50541, n50542, n50543, n50544, n50545, n50546, n50547,
         n50548, n50549, n50550, n50551, n50552, n50553, n50554, n50555,
         n50556, n50557, n50558, n50559, n50560, n50561, n50562, n50563,
         n50564, n50565, n50566, n50567, n50568, n50570, n50571, n50572,
         n50573, n50574, n50575, n50576, n50577, n50578, n50579, n50580,
         n50581, n50582, n50583, n50584, n50585, n50586, n50587, n50588,
         n50589, n50590, n50591, n50592, n50593, n50594, n50595, n50596,
         n50597, n50598, n50599, n50600, n50601, n50602, n50603, n50604,
         n50605, n50606, n50607, n50608, n50609, n50610, n50611, n50612,
         n50613, n50614, n50615, n50616, n50617, n50618, n50619, n50620,
         n50621, n50622, n50623, n50624, n50625, n50626, n50627, n50628,
         n50629, n50630, n50631, n50632, n50633, n50634, n50635, n50636,
         n50637, n50638, n50639, n50640, n50641, n50642, n50643, n50644,
         n50645, n50646, n50647, n50648, n50649, n50650, n50651, n50652,
         n50653, n50654, n50655, n50656, n50657, n50658, n50659, n50660,
         n50661, n50662, n50663, n50664, n50665, n50666, n50667, n50668,
         n50669, n50670, n50671, n50672, n50673, n50674, n50675, n50676,
         n50677, n50678, n50679, n50680, n50681, n50682, n50683, n50684,
         n50685, n50686, n50687, n50688, n50689, n50690, n50691, n50692,
         n50693, n50694, n50695, n50696, n50697, n50698, n50699, n50700,
         n50701, n50702, n50703, n50704, n50705, n50706, n50707, n50708,
         n50709, n50710, n50711, n50712, n50713, n50714, n50715, n50716,
         n50717, n50718, n50719, n50720, n50721, n50722, n50723, n50724,
         n50725, n50726, n50727, n50728, n50729, n50730, n50731, n50732,
         n50733, n50734, n50735, n50736, n50737, n50738, n50739, n50740,
         n50741, n50742, n50743, n50744, n50745, n50746, n50747, n50748,
         n50749, n50750, n50751, n50752, n50753, n50754, n50755, n50756,
         n50757, n50758, n50759, n50761, n50762, n50763, n50764, n50765,
         n50766, n50767, n50768, n50769, n50770, n50771, n50772, n50773,
         n50774, n50775, n50776, n50777, n50778, n50779, n50780, n50781,
         n50782, n50783, n50784, n50785, n50786, n50787, n50788, n50790,
         n50791, n50792, n50793, n50794, n50795, n50797, n50798, n50799,
         n50800, n50801, n50802, n50803, n50804, n50805, n50806, n50807,
         n50808, n50809, n50810, n50811, n50812, n50813, n50814, n50815,
         n50816, n50817, n50819, n50820, n50821, n50822, n50823, n50824,
         n50825, n50826, n50827, n50828, n50829, n50830, n50831, n50832,
         n50833, n50834, n50835, n50836, n50837, n50839, n50840, n50841,
         n50842, n50843, n50844, n50845, n50846, n50847, n50848, n50849,
         n50850, n50851, n50852, n50853, n50854, n50855, n50856, n50857,
         n50858, n50859, n50860, n50861, n50862, n50863, n50864, n50865,
         n50866, n50867, n50868, n50869, n50870, n50871, n50872, n50873,
         n50874, n50875, n50876, n50877, n50878, n50879, n50880, n50881,
         n50882, n50883, n50884, n50885, n50886, n50887, n50888, n50889,
         n50890, n50892, n50893, n50894, n50895, n50896, n50897, n50898,
         n50899, n50900, n50901, n50902, n50903, n50904, n50906, n50907,
         n50908, n50909, n50910, n50911, n50912, n50913, n50914, n50915,
         n50916, n50917, n50918, n50919, n50920, n50921, n50922, n50923,
         n50924, n50925, n50926, n50927, n50928, n50929, n50930, n50931,
         n50932, n50933, n50934, n50935, n50936, n50937, n50938, n50939,
         n50940, n50941, n50942, n50943, n50944, n50945, n50946, n50947,
         n50948, n50949, n50950, n50951, n50952, n50953, n50954, n50955,
         n50956, n50957, n50958, n50959, n50960, n50961, n50962, n50963,
         n50964, n50965, n50966, n50967, n50976, n50977, n50980, n50981,
         n50982, n50983, n50984, n50986, n50987, n50990, n50991, n50992,
         n50997, n51001, n51004, n51006, n51009, n51012, n51013, n51014,
         n51015, n51016, n51017, n51018, n51019, n51021, n51022, n51023,
         n51025, n51026, n51029, n51031, n51032, n51033, n51034, n51039,
         n51046, n51047, n51048, n51049, n51050, n51052, n51056, n51057,
         n51058, n51062, n51063, n51064, n51066, n51067, n51068, n51072,
         n51077, n51080, n51081, n51085, n51086, n51087, n51088, n51090,
         n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51099,
         n51100, n51101, n51102, n51103, n51105, n51106, n51107, n51108,
         n51109, n51110, n51111, n51112, n51113, n51114, n51115, n51116,
         n51117, n51118, n51119, n51120, n51121, n51122, n51123, n51124,
         n51125, n51126, n51127, n51128, n51129, n51130, n51132, n51133,
         n51134, n51135, n51136, n51137, n51138, n51139, n51140, n51141,
         n51142, n51143, n51144, n51145, n51146, n51147, n51148, n51149,
         n51150, n51151, n51152, n51153, n51154, n51155, n51156, n51157,
         n51158, n51159, n51160, n51161, n51162, n51163, n51164, n51165,
         n51166, n51167, n51168, n51169, n51170, n51171, n51172, n51173,
         n51174, n51175, n51176, n51177, n51178, n51179, n51180, n51181,
         n51182, n51183, n51185, n51186, n51187, n51189, n51190, n51191,
         n51192, n51193, n51194, n51196, n51197, n51198, n51199, n51200,
         n51201, n51202, n51203, n51204, n51205, n51206, n51207, n51208,
         n51209, n51210, n51211, n51212, n51213, n51214, n51215, n51216,
         n51217, n51218, n51219, n51220, n51222, n51223, n51224, n51225,
         n51226, n51227, n51228, n51229, n51230, n51231, n51232, n51233,
         n51234, n51235, n51236, n51237, n51238, n51239, n51240, n51241,
         n51242, n51243, n51244, n51245, n51246, n51247, n51248, n51249,
         n51250, n51251, n51252, n51253, n51254, n51255, n51256, n51257,
         n51258, n51259, n51261, n51262, n51263, n51264, n51265, n51266,
         n51267, n51269, n51270, n51271, n51272, n51273, n51274, n51276,
         n51277, n51278, n51279, n51281, n51282, n51283, n51284, n51285,
         n51286, n51287, n51289, n51290, n51291, n51292, n51294, n51295,
         n51296, n51297, n51298, n51299, n51300, n51301, n51302, n51303,
         n51304, n51305, n51306, n51307, n51308, n51309, n51310, n51312,
         n51313, n51314, n51315, n51316, n51317, n51318, n51320, n51321,
         n51322, n51323, n51324, n51325, n51326, n51327, n51328, n51329,
         n51330, n51331, n51332, n51333, n51334, n51335, n51336, n51337,
         n51338, n51339, n51340, n51341, n51342, n51343, n51344, n51346,
         n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354,
         n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362,
         n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370,
         n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378,
         n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386,
         n51388, n51389, n51390, n51391, n51392, n51393, n51394, n51395,
         n51396, n51397, n51398, n51399, n51400, n51401, n51402, n51403,
         n51404, n51406, n51407, n51408, n51409, n51410, n51411, n51413,
         n51414, n51415, n51416, n51417, n51418, n51419, n51420, n51421,
         n51422, n51423, n51424, n51425, n51426, n51427, n51429, n51430,
         n51431, n51432, n51433, n51434, n51435, n51436, n51437, n51438,
         n51439, n51440, n51441, n51442, n51444, n51445, n51446, n51447,
         n51448, n51449, n51450, n51451, n51452, n51453, n51454, n51455,
         n51456, n51458, n51459, n51460, n51461, n51462, n51463, n51464,
         n51465, n51467, n51468, n51469, n51470, n51471, n51472, n51473,
         n51474, n51478, n51479, n51480, n51481, n51482, n51483, n51484,
         n51485, n51486, n51487, n51488, n51489, n51490, n51491, n51492,
         n51493, n51494, n51495, n51496, n51497, n51498, n51500, n51501,
         n51502, n51503, n51504, n51507, n51508, n51509, n51510, n51511,
         n51512, n51513, n51514, n51515, n51516, n51517, n51518, n51519,
         n51520, n51521, n51522, n51523, n51524, n51525, n51526, n51529,
         n51530, n51531, n51532, n51533, n51534, n51535, n51536, n51537,
         n51538, n51539, n51540, n51541, n51542, n51543, n51544, n51545,
         n51546, n51547, n51548, n51549, n51550, n51551, n51552, n51553,
         n51554, n51556, n51557, n51558, n51559, n51560, n51562, n51564,
         n51565, n51566, n51567, n51568, n51569, n51570, n51571, n51572,
         n51573, n51574, n51575, n51576, n51577, n51578, n51579, n51580,
         n51581, n51582, n51583, n51584, n51585, n51586, n51587, n51588,
         n51589, n51590, n51591, n51592, n51593, n51594, n51595, n51596,
         n51597, n51598, n51599, n51601, n51602, n51603, n51605, n51606,
         n51607, n51608, n51609, n51610, n51611, n51612, n51613, n51614,
         n51616, n51617, n51618, n51619, n51620, n51621, n51622, n51623,
         n51624, n51625, n51626, n51627, n51628, n51629, n51630, n51631,
         n51632, n51633, n51634, n51635, n51636, n51637, n51638, n51639,
         n51640, n51641, n51642, n51643, n51644, n51645, n51646, n51647,
         n51648, n51649, n51650, n51652, n51653, n51654, n51655, n51656,
         n51657, n51658, n51659, n51660, n51661, n51662, n51663, n51664,
         n51665, n51666, n51667, n51668, n51669, n51670, n51671, n51672,
         n51673, n51674, n51675, n51676, n51677, n51678, n51679, n51680,
         n51681, n51682, n51683, n51684, n51685, n51686, n51687, n51688,
         n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696,
         n51697, n51698, n51699, n51700, n51702, n51703, n51704, n51705,
         n51706, n51708, n51709, n51710, n51711, n51712, n51713, n51714,
         n51715, n51716, n51717, n51719, n51720, n51721, n51722, n51723,
         n51724, n51725, n51726, n51727, n51728, n51729, n51730, n51731,
         n51732, n51733, n51734, n51735, n51736, n51737, n51738, n51739,
         n51740, n51742, n51743, n51744, n51746, n51747, n51748, n51749,
         n51750, n51751, n51752, n51753, n51754, n51755, n51756, n51757,
         n51758, n51760, n51761, n51762, n51763, n51764, n51765, n51766,
         n51767, n51768, n51769, n51770, n51771, n51772, n51773, n51774,
         n51775, n51776, n51777, n51778, n51779, n51780, n51781, n51782,
         n51783, n51784, n51785, n51786, n51787, n51788, n51789, n51790,
         n51791, n51792, n51793, n51794, n51795, n51796, n51797, n51798,
         n51799, n51800, n51801, n51802, n51803, n51804, n51805, n51806,
         n51807, n51808, n51809, n51810, n51811, n51812, n51813, n51814,
         n51815, n51816, n51817, n51818, n51819, n51820, n51821, n51822,
         n51823, n51824, n51825, n51826, n51827, n51828, n51829, n51830,
         n51831, n51832, n51833, n51834, n51835, n51836, n51837, n51838,
         n51839, n51840, n51841, n51842, n51843, n51844, n51845, n51846,
         n51847, n51848, n51849, n51850, n51851, n51852, n51853, n51854,
         n51855, n51856, n51857, n51858, n51859, n51860, n51861, n51862,
         n51863, n51864, n51865, n51866, n51867, n51868, n51869, n51870,
         n51871, n51872, n51873, n51874, n51875, n51876, n51877, n51878,
         n51879, n51880, n51881, n51882, n51883, n51884, n51885, n51886,
         n51887, n51888, n51889, n51890, n51891, n51892, n51893, n51894,
         n51895, n51896, n51897, n51898, n51899, n51900, n51901, n51902,
         n51903, n51904, n51905, n51906, n51907, n51908, n51909, n51910,
         n51911, n51912, n51913, n51914, n51915, n51916, n51917, n51918,
         n51919, n51920, n51921, n51922, n51923, n51924, n51925, n51926,
         n51927, n51928, n51929, n51930, n51931, n51932, n51933, n51934,
         n51935, n51936, n51937, n51938, n51939, n51940, n51941, n51942,
         n51943, n51944, n51945, n51946, n51947, n51948, n51949, n51950,
         n51951, n51952, n51953, n51954, n51955, n51956, n51957, n51958,
         n51959, n51960, n51961, n51962, n51963, n51964, n51965, n51966,
         n51967, n51968, n51969, n51970, n51971, n51972, n51973, n51974,
         n51975, n51976, n51977, n51978, n51979, n51980, n51981, n51982,
         n51983, n51984, n51985, n51986, n51987, n51988, n51989, n51990,
         n51991, n51992, n51993, n51994, n51995, n51996, n51997, n51998,
         n51999, n52000, n52001, n52002, n52003, n52004, n52005, n52006,
         n52007, n52008, n52009, n52010, n52011, n52012, n52013, n52014,
         n52015, n52016, n52017, n52018, n52019, n52020, n52021, n52022,
         n52023, n52024, n52025, n52026, n52027, n52028, n52029, n52030,
         n52031, n52032, n52033, n52034, n52035, n52036, n52037, n52038,
         n52039, n52040, n52041, n52042, n52043, n52044, n52045, n52046,
         n52047, n52048, n52049, n52050, n52051, n52052, n52053, n52054,
         n52055, n52056, n52057, n52058, n52059, n52060, n52061, n52062,
         n52063, n52064, n52065, n52066, n52067, n52068, n52069, n52070,
         n52071, n52072, n52073, n52074, n52075, n52076, n52077, n52078,
         n52079, n52080, n52081, n52082, n52083, n52084, n52085, n52086,
         n52087, n52088, n52089, n52090, n52091, n52092, n52093, n52094,
         n52095, n52096, n52097, n52098, n52099, n52100, n52101, n52102,
         n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110,
         n52111, n52112, n52113, n52114, n52115, n52116, n52117, n52118,
         n52119, n52120, n52121, n52122, n52123, n52124, n52125, n52126,
         n52127, n52128, n52129, n52130, n52131, n52132, n52133, n52134,
         n52135, n52136, n52137, n52138, n52139, n52140, n52141, n52142,
         n52143, n52144, n52145, n52146, n52147, n52148, n52149, n52150,
         n52151, n52152, n52153, n52154, n52155, n52156, n52157, n52158,
         n52159, n52160, n52161, n52162, n52163, n52164, n52165, n52166,
         n52167, n52168, n52169, n52170, n52171, n52172, n52173, n52174,
         n52175, n52176, n52177, n52178, n52179, n52180, n52181, n52182,
         n52183, n52184, n52185, n52186, n52187, n52188, n52189, n52190,
         n52191, n52192, n52193, n52194, n52195, n52196, n52197, n52198,
         n52199, n52200, n52201, n52202, n52203, n52204, n52205, n52206,
         n52207, n52208, n52209, n52210, n52211, n52212, n52213, n52214,
         n52215, n52216, n52217, n52218, n52219, n52220, n52221, n52222,
         n52223, n52224, n52225, n52226, n52227, n52228, n52229, n52230,
         n52231, n52232, n52233, n52234, n52235, n52236, n52237, n52238,
         n52239, n52240, n52241, n52242, n52243, n52244, n52245, n52246,
         n52247, n52248, n52249, n52250, n52251, n52252, n52253, n52254,
         n52255, n52256, n52257, n52258, n52259, n52260, n52261, n52262,
         n52263, n52264, n52265, n52266, n52267, n52268, n52269, n52270,
         n52271, n52272, n52273, n52274, n52275, n52276, n52277, n52278,
         n52279, n52280, n52281, n52282, n52283, n52284, n52285, n52286,
         n52287, n52288, n52289, n52290, n52291, n52292, n52293, n52294,
         n52295, n52296, n52297, n52298, n52299, n52300, n52301, n52302,
         n52303, n52304, n52305, n52306, n52307, n52308, n52309, n52310,
         n52311, n52312, n52313, n52314, n52315, n52316, n52317, n52318,
         n52319, n52320, n52321, n52322, n52323, n52324, n52325, n52326,
         n52327, n52328, n52329, n52330, n52331, n52332, n52333, n52334,
         n52335, n52336, n52337, n52338, n52339, n52340, n52341, n52342,
         n52343, n52344, n52345, n52346, n52347, n52348, n52349, n52350,
         n52351, n52352, n52353, n52354, n52355, n52356, n52357, n52358,
         n52359, n52360, n52361, n52362, n52363, n52364, n52365, n52366,
         n52367, n52368, n52369, n52370, n52371, n52372, n52373, n52374,
         n52375, n52376, n52377, n52378, n52379, n52380, n52381, n52382,
         n52383, n52384, n52385, n52386, n52387, n52388, n52389, n52390,
         n52391, n52392, n52393, n52394, n52395, n52396, n52397, n52398,
         n52399, n52400, n52401, n52402, n52403, n52404, n52405, n52406,
         n52407, n52408, n52409, n52410, n52411, n52412, n52413, n52414,
         n52415, n52416, n52417, n52418, n52419, n52420, n52421, n52422,
         n52423, n52424, n52425, n52426, n52427, n52428, n52429, n52430,
         n52431, n52432, n52433, n52434;

  AND2_X1 U1 ( .A1(n50731), .A2(n50700), .ZN(n44630) );
  OR2_X1 U2 ( .A1(n48912), .A2(n48853), .ZN(n48918) );
  BUF_X1 U8 ( .A(n50854), .Z(n601) );
  AND2_X1 U9 ( .A1(n1716), .A2(n1717), .ZN(n47991) );
  NOR2_X1 U14 ( .A1(n47326), .A2(n50390), .ZN(n139) );
  OR2_X1 U15 ( .A1(n50372), .A2(n667), .ZN(n134) );
  AND2_X1 U16 ( .A1(n45802), .A2(n46746), .ZN(n86) );
  AND2_X1 U17 ( .A1(n46743), .A2(n1760), .ZN(n46751) );
  AND2_X1 U25 ( .A1(n7577), .A2(n49231), .ZN(n145) );
  AND2_X1 U32 ( .A1(n5895), .A2(n5892), .ZN(n42122) );
  AND2_X1 U34 ( .A1(n36095), .A2(n7241), .ZN(n7237) );
  NAND4_X1 U35 ( .A1(n40844), .A2(n40843), .A3(n40842), .A4(n40841), .ZN(
        n42643) );
  AND2_X1 U37 ( .A1(n40476), .A2(n41268), .ZN(n58) );
  OR2_X1 U38 ( .A1(n39707), .A2(n39706), .ZN(n55) );
  INV_X1 U39 ( .A(n38814), .ZN(n40637) );
  NOR2_X1 U40 ( .A1(n51633), .A2(n186), .ZN(n185) );
  OR2_X1 U41 ( .A1(n38810), .A2(n41792), .ZN(n41799) );
  AND3_X1 U43 ( .A1(n41645), .A2(n41650), .A3(n41647), .ZN(n226) );
  OR2_X1 U44 ( .A1(n6859), .A2(n38416), .ZN(n246) );
  INV_X1 U48 ( .A(n40792), .ZN(n40777) );
  INV_X1 U49 ( .A(n40558), .ZN(n40564) );
  AND3_X1 U51 ( .A1(n1335), .A2(n241), .A3(n36784), .ZN(n8644) );
  AND2_X1 U52 ( .A1(n68), .A2(n37219), .ZN(n38263) );
  AOI22_X1 U53 ( .A1(n3027), .A2(n34797), .B1(n34799), .B2(n34798), .ZN(n2) );
  OR2_X1 U54 ( .A1(n36640), .A2(n36629), .ZN(n38072) );
  OR2_X1 U55 ( .A1(n38196), .A2(n6869), .ZN(n263) );
  OR2_X1 U56 ( .A1(n35736), .A2(n36410), .ZN(n289) );
  NOR2_X1 U58 ( .A1(n38949), .A2(n39210), .ZN(n38943) );
  NAND2_X1 U59 ( .A1(n35888), .A2(n38341), .ZN(n14) );
  NAND2_X1 U61 ( .A1(n39273), .A2(n5262), .ZN(n39270) );
  OR2_X1 U63 ( .A1(n38565), .A2(n36105), .ZN(n38570) );
  AND2_X1 U64 ( .A1(n38200), .A2(n35151), .ZN(n38567) );
  BUF_X1 U69 ( .A(n32678), .Z(n35028) );
  INV_X1 U71 ( .A(n38635), .ZN(n197) );
  INV_X1 U73 ( .A(n37023), .ZN(n165) );
  XNOR2_X1 U74 ( .A(n50983), .B(n31187), .ZN(n82) );
  BUF_X1 U75 ( .A(n35104), .Z(n35471) );
  XNOR2_X1 U76 ( .A(n2155), .B(n36869), .ZN(n35372) );
  NAND4_X1 U81 ( .A1(n30524), .A2(n30523), .A3(n30522), .A4(n30521), .ZN(
        n32860) );
  AOI21_X1 U82 ( .B1(n33116), .B2(n33115), .A(n33114), .ZN(n33893) );
  AND4_X1 U83 ( .A1(n30909), .A2(n30596), .A3(n30595), .A4(n30594), .ZN(n30615) );
  AND2_X1 U84 ( .A1(n32992), .A2(n32993), .ZN(n200) );
  AND3_X1 U85 ( .A1(n30970), .A2(n1099), .A3(n1098), .ZN(n30972) );
  OR2_X1 U86 ( .A1(n29587), .A2(n31111), .ZN(n1129) );
  OR2_X1 U87 ( .A1(n30935), .A2(n30082), .ZN(n30080) );
  OR2_X1 U88 ( .A1(n29840), .A2(n169), .ZN(n31272) );
  AND2_X1 U89 ( .A1(n31934), .A2(n31338), .ZN(n19) );
  AND2_X1 U90 ( .A1(n31221), .A2(n32209), .ZN(n31224) );
  INV_X1 U91 ( .A(n706), .ZN(n31640) );
  OR2_X1 U92 ( .A1(n31512), .A2(n30925), .ZN(n29648) );
  AND2_X1 U93 ( .A1(n32212), .A2(n32210), .ZN(n31221) );
  NOR2_X1 U94 ( .A1(n29618), .A2(n29622), .ZN(n28164) );
  NOR2_X1 U97 ( .A1(n51744), .A2(n31338), .ZN(n31347) );
  AND2_X1 U100 ( .A1(n32916), .A2(n32909), .ZN(n158) );
  INV_X1 U101 ( .A(n29622), .ZN(n32990) );
  OR2_X1 U102 ( .A1(n31873), .A2(n31870), .ZN(n31028) );
  INV_X1 U103 ( .A(n31748), .ZN(n31740) );
  AND2_X1 U106 ( .A1(n29857), .A2(n29856), .ZN(n70) );
  AND2_X1 U108 ( .A1(n29545), .A2(n29557), .ZN(n27048) );
  OR2_X1 U109 ( .A1(n30784), .A2(n160), .ZN(n6789) );
  NOR2_X1 U110 ( .A1(n29131), .A2(n159), .ZN(n29136) );
  AND2_X1 U111 ( .A1(n29132), .A2(n30181), .ZN(n159) );
  AOI21_X1 U112 ( .B1(n28555), .B2(n2110), .A(n51748), .ZN(n195) );
  AND2_X1 U113 ( .A1(n29306), .A2(n29291), .ZN(n29311) );
  AND2_X1 U114 ( .A1(n28517), .A2(n2328), .ZN(n30446) );
  AND2_X1 U115 ( .A1(n27881), .A2(n29346), .ZN(n1059) );
  INV_X1 U117 ( .A(n29495), .ZN(n257) );
  INV_X1 U119 ( .A(n30783), .ZN(n161) );
  AND2_X1 U121 ( .A1(n30461), .A2(n427), .ZN(n2328) );
  OR2_X1 U122 ( .A1(n28841), .A2(n30461), .ZN(n29735) );
  AND2_X1 U123 ( .A1(n27680), .A2(n27686), .ZN(n27579) );
  AND2_X1 U124 ( .A1(n28449), .A2(n29749), .ZN(n28841) );
  AND2_X1 U126 ( .A1(n28523), .A2(n28521), .ZN(n28991) );
  AND2_X1 U128 ( .A1(n27119), .A2(n27987), .ZN(n177) );
  AND2_X1 U135 ( .A1(n28874), .A2(n29029), .ZN(n29045) );
  BUF_X1 U138 ( .A(n27633), .Z(n597) );
  BUF_X1 U141 ( .A(n23651), .Z(n25669) );
  OAI21_X2 U142 ( .B1(n24018), .B2(n24017), .A(n24016), .ZN(n26377) );
  AND3_X1 U143 ( .A1(n20553), .A2(n7718), .A3(n20554), .ZN(n27197) );
  AND2_X1 U146 ( .A1(n20282), .A2(n20281), .ZN(n20288) );
  AND2_X1 U147 ( .A1(n22144), .A2(n19560), .ZN(n19563) );
  AOI21_X1 U150 ( .B1(n22183), .B2(n22180), .A(n22179), .ZN(n22181) );
  AND2_X1 U151 ( .A1(n3876), .A2(n23171), .ZN(n22548) );
  OR2_X1 U152 ( .A1(n24124), .A2(n24123), .ZN(n119) );
  OR2_X1 U153 ( .A1(n23708), .A2(n5415), .ZN(n171) );
  OR2_X1 U159 ( .A1(n23531), .A2(n50990), .ZN(n4882) );
  INV_X1 U164 ( .A(n22506), .ZN(n288) );
  AOI22_X1 U165 ( .A1(n20652), .A2(n15834), .B1(n15833), .B2(n15832), .ZN(
        n15839) );
  INV_X1 U166 ( .A(n19950), .ZN(n21423) );
  OAI21_X1 U167 ( .B1(n18893), .B2(n21528), .A(n301), .ZN(n3458) );
  INV_X1 U168 ( .A(n20131), .ZN(n20130) );
  OR2_X1 U169 ( .A1(n15630), .A2(n19891), .ZN(n19896) );
  AOI21_X1 U170 ( .B1(n21544), .B2(n20624), .A(n6929), .ZN(n18494) );
  NAND2_X1 U171 ( .A1(n19391), .A2(n19392), .ZN(n76) );
  OR2_X1 U172 ( .A1(n20052), .A2(n20062), .ZN(n19135) );
  BUF_X1 U176 ( .A(n19860), .Z(n585) );
  BUF_X1 U177 ( .A(n1417), .Z(n18344) );
  NOR2_X1 U179 ( .A1(n5058), .A2(n17018), .ZN(n20119) );
  AND2_X1 U181 ( .A1(n17577), .A2(n17576), .ZN(n19389) );
  BUF_X1 U183 ( .A(n18865), .Z(n498) );
  OR2_X1 U184 ( .A1(n15400), .A2(n17873), .ZN(n2222) );
  OAI211_X1 U186 ( .C1(n15249), .C2(n15248), .A(n15247), .B(n15246), .ZN(
        n16416) );
  NOR2_X1 U188 ( .A1(n14831), .A2(n15448), .ZN(n128) );
  NOR2_X1 U189 ( .A1(n15030), .A2(n69), .ZN(n11806) );
  INV_X1 U190 ( .A(n13801), .ZN(n69) );
  OR2_X1 U191 ( .A1(n11820), .A2(n13102), .ZN(n12820) );
  OR2_X1 U192 ( .A1(n12894), .A2(n12893), .ZN(n64) );
  AND3_X1 U193 ( .A1(n7734), .A2(n14816), .A3(n14815), .ZN(n5257) );
  OR2_X1 U195 ( .A1(n15357), .A2(n15380), .ZN(n205) );
  BUF_X1 U197 ( .A(Key[175]), .Z(n4529) );
  BUF_X1 U198 ( .A(Key[157]), .Z(n4712) );
  BUF_X1 U199 ( .A(Key[65]), .Z(n4645) );
  CLKBUF_X1 U200 ( .A(Key[166]), .Z(n4471) );
  BUF_X1 U201 ( .A(Key[121]), .Z(n45736) );
  BUF_X1 U202 ( .A(Key[104]), .Z(n49323) );
  BUF_X1 U203 ( .A(Key[21]), .Z(n45883) );
  INV_X1 U204 ( .A(n14033), .ZN(n47) );
  BUF_X1 U205 ( .A(Key[136]), .Z(n1341) );
  BUF_X1 U207 ( .A(Key[106]), .Z(n4585) );
  NAND4_X2 U212 ( .A1(n10753), .A2(n10752), .A3(n10751), .A4(n10750), .ZN(
        n14006) );
  AND2_X1 U215 ( .A1(n8901), .A2(n12678), .ZN(n32) );
  OAI211_X1 U216 ( .C1(n9750), .C2(n9749), .A(n9748), .B(n875), .ZN(n3418) );
  INV_X1 U217 ( .A(n9423), .ZN(n12251) );
  OAI21_X1 U219 ( .B1(n10939), .B2(n12314), .A(n12309), .ZN(n8) );
  AND2_X1 U221 ( .A1(n10302), .A2(n12303), .ZN(n9758) );
  BUF_X1 U222 ( .A(n11932), .Z(n2156) );
  CLKBUF_X1 U223 ( .A(n11899), .Z(n510) );
  BUF_X1 U225 ( .A(n9207), .Z(n12631) );
  INV_X1 U228 ( .A(n11932), .ZN(n12709) );
  AND2_X1 U229 ( .A1(n9001), .A2(n10722), .ZN(n12292) );
  OR2_X1 U231 ( .A1(n11884), .A2(n11501), .ZN(n8901) );
  BUF_X1 U232 ( .A(n12496), .Z(n642) );
  BUF_X1 U233 ( .A(n9204), .Z(n10465) );
  BUF_X1 U236 ( .A(n12453), .Z(n592) );
  XNOR2_X2 U246 ( .A(n26540), .B(n28274), .ZN(n27235) );
  AND2_X2 U247 ( .A1(n7288), .A2(n20774), .ZN(n22623) );
  OR2_X1 U249 ( .A1(n19761), .A2(n22979), .ZN(n19038) );
  NOR2_X1 U250 ( .A1(n32725), .A2(n1085), .ZN(n32715) );
  XNOR2_X1 U254 ( .A(n42535), .B(n42534), .ZN(n43742) );
  AND2_X1 U256 ( .A1(n46279), .A2(n23), .ZN(n49008) );
  AOI22_X1 U258 ( .A1(n27011), .A2(n27010), .B1(n27755), .B2(n27743), .ZN(
        n27021) );
  AND2_X1 U259 ( .A1(n51346), .A2(n47573), .ZN(n47519) );
  NOR2_X1 U269 ( .A1(n36777), .A2(n36776), .ZN(n36786) );
  OR2_X1 U271 ( .A1(n39201), .A2(n38943), .ZN(n247) );
  OR2_X1 U272 ( .A1(n30449), .A2(n29734), .ZN(n28526) );
  INV_X1 U274 ( .A(n49037), .ZN(n23) );
  NOR2_X1 U276 ( .A1(n49377), .A2(n51729), .ZN(n49349) );
  INV_X1 U278 ( .A(n49574), .ZN(n43407) );
  OR2_X1 U279 ( .A1(n52151), .A2(n40822), .ZN(n40839) );
  INV_X1 U283 ( .A(n50299), .ZN(n49953) );
  OR2_X1 U285 ( .A1(n42105), .A2(n41797), .ZN(n38814) );
  OR2_X1 U287 ( .A1(n50465), .A2(n544), .ZN(n50435) );
  AND2_X1 U288 ( .A1(n51344), .A2(n2092), .ZN(n45190) );
  OR2_X1 U289 ( .A1(n49308), .A2(n49309), .ZN(n49311) );
  OR2_X1 U291 ( .A1(n49217), .A2(n132), .ZN(n131) );
  OR2_X1 U294 ( .A1(n38409), .A2(n38410), .ZN(n38412) );
  INV_X1 U300 ( .A(n46632), .ZN(n44423) );
  OR2_X1 U301 ( .A1(n46632), .A2(n44864), .ZN(n5309) );
  AND2_X1 U303 ( .A1(n50188), .A2(n50233), .ZN(n93) );
  OR2_X1 U308 ( .A1(n26937), .A2(n27668), .ZN(n26871) );
  INV_X1 U310 ( .A(n20343), .ZN(n50) );
  AND2_X1 U313 ( .A1(n29426), .A2(n26905), .ZN(n29429) );
  AND2_X2 U321 ( .A1(n2086), .A2(n36571), .ZN(n36565) );
  AND2_X1 U322 ( .A1(n174), .A2(n47934), .ZN(n173) );
  INV_X1 U323 ( .A(n20752), .ZN(n20739) );
  OR2_X1 U326 ( .A1(n36045), .A2(n36052), .ZN(n36050) );
  AND2_X1 U328 ( .A1(n13797), .A2(n13804), .ZN(n15030) );
  AND2_X1 U329 ( .A1(n9279), .A2(n11590), .ZN(n11247) );
  XNOR2_X1 U331 ( .A(n5612), .B(n8087), .ZN(n35104) );
  OR2_X1 U332 ( .A1(n15257), .A2(n15259), .ZN(n15266) );
  NAND2_X1 U335 ( .A1(n51049), .A2(n3243), .ZN(n21520) );
  OR2_X1 U336 ( .A1(n19170), .A2(n20428), .ZN(n20420) );
  NOR2_X1 U339 ( .A1(n14545), .A2(n14550), .ZN(n13362) );
  XNOR2_X1 U340 ( .A(n26414), .B(n26413), .ZN(n83) );
  NAND4_X2 U341 ( .A1(n31736), .A2(n31738), .A3(n31735), .A4(n31737), .ZN(
        n34604) );
  NAND3_X1 U350 ( .A1(n35948), .A2(n38504), .A3(n35574), .ZN(n35585) );
  INV_X1 U356 ( .A(n41025), .ZN(n40422) );
  AND2_X1 U357 ( .A1(n41025), .A2(n41034), .ZN(n35185) );
  NAND2_X1 U359 ( .A1(n986), .A2(n48464), .ZN(n985) );
  NAND2_X1 U360 ( .A1(n5324), .A2(n397), .ZN(n8613) );
  NAND3_X1 U363 ( .A1(n46814), .A2(n46767), .A3(n4), .ZN(n47085) );
  XNOR2_X2 U365 ( .A(n34407), .B(n5), .ZN(n36052) );
  XNOR2_X1 U366 ( .A(n34394), .B(n34395), .ZN(n5) );
  AND2_X1 U368 ( .A1(n21142), .A2(n21141), .ZN(n6) );
  NAND2_X1 U379 ( .A1(n10952), .A2(n7), .ZN(n9661) );
  INV_X1 U380 ( .A(n8), .ZN(n7) );
  NOR2_X1 U381 ( .A1(n9772), .A2(n10938), .ZN(n10952) );
  AOI21_X1 U383 ( .B1(n11433), .B2(n9), .A(n14103), .ZN(n6491) );
  NAND4_X2 U384 ( .A1(n22451), .A2(n22450), .A3(n22449), .A4(n22448), .ZN(
        n25755) );
  NAND3_X1 U385 ( .A1(n28637), .A2(n28641), .A3(n28636), .ZN(n28648) );
  XNOR2_X2 U387 ( .A(n28431), .B(n25320), .ZN(n27445) );
  NAND4_X2 U388 ( .A1(n23325), .A2(n23324), .A3(n23326), .A4(n23327), .ZN(
        n28431) );
  NAND2_X1 U389 ( .A1(n10), .A2(n9436), .ZN(n5510) );
  NAND2_X1 U390 ( .A1(n5512), .A2(n12133), .ZN(n10) );
  NAND4_X2 U393 ( .A1(n28612), .A2(n28613), .A3(n32594), .A4(n28611), .ZN(
        n36672) );
  NAND2_X1 U400 ( .A1(n14), .A2(n12), .ZN(n35892) );
  NAND2_X1 U401 ( .A1(n13), .A2(n35407), .ZN(n12) );
  OAI22_X1 U402 ( .A1(n6615), .A2(n38339), .B1(n38335), .B2(n38337), .ZN(n13)
         );
  XNOR2_X1 U404 ( .A(n16), .B(n35373), .ZN(n35406) );
  XNOR2_X1 U405 ( .A(n35369), .B(n35370), .ZN(n16) );
  INV_X1 U407 ( .A(n17), .ZN(n13194) );
  OAI21_X1 U408 ( .B1(n13947), .B2(n13193), .A(n13192), .ZN(n17) );
  OR2_X2 U414 ( .A1(n18), .A2(n8289), .ZN(n30037) );
  NAND3_X1 U415 ( .A1(n2674), .A2(n2670), .A3(n2672), .ZN(n18) );
  NAND2_X1 U416 ( .A1(n31339), .A2(n19), .ZN(n31343) );
  NAND2_X1 U417 ( .A1(n31931), .A2(n31346), .ZN(n31339) );
  NAND2_X1 U420 ( .A1(n7954), .A2(n36121), .ZN(n36131) );
  AND2_X2 U421 ( .A1(n10945), .A2(n9057), .ZN(n10939) );
  NAND2_X1 U424 ( .A1(n31910), .A2(n31075), .ZN(n32850) );
  AND4_X2 U425 ( .A1(n3743), .A2(n28855), .A3(n28856), .A4(n3744), .ZN(n31075)
         );
  NAND4_X1 U426 ( .A1(n9369), .A2(n51138), .A3(n11353), .A4(n10687), .ZN(
        n12092) );
  NOR2_X2 U432 ( .A1(n6226), .A2(n19510), .ZN(n598) );
  NAND2_X1 U434 ( .A1(n25836), .A2(n8744), .ZN(n26329) );
  NAND2_X1 U435 ( .A1(n42618), .A2(n48971), .ZN(n42807) );
  NAND3_X1 U442 ( .A1(n3197), .A2(n20065), .A3(n6022), .ZN(n3196) );
  NAND3_X1 U443 ( .A1(n18501), .A2(n18502), .A3(n18500), .ZN(n18503) );
  NAND2_X1 U445 ( .A1(n22), .A2(n11771), .ZN(n4963) );
  OAI211_X1 U446 ( .C1(n11767), .C2(n11768), .A(n12886), .B(n11766), .ZN(n22)
         );
  NAND2_X1 U449 ( .A1(n40185), .A2(n41193), .ZN(n40186) );
  NAND2_X1 U450 ( .A1(n2896), .A2(n38627), .ZN(n2895) );
  NAND2_X1 U451 ( .A1(n20082), .A2(n16218), .ZN(n20072) );
  NAND4_X2 U460 ( .A1(n19941), .A2(n24), .A3(n19940), .A4(n19939), .ZN(n24030)
         );
  NAND4_X1 U461 ( .A1(n19936), .A2(n19937), .A3(n19935), .A4(n19938), .ZN(n24)
         );
  AND2_X1 U464 ( .A1(n14318), .A2(n51064), .ZN(n25) );
  NAND2_X1 U469 ( .A1(n8908), .A2(n8909), .ZN(n11082) );
  NAND2_X1 U470 ( .A1(n30147), .A2(n28600), .ZN(n5706) );
  NAND3_X1 U471 ( .A1(n28535), .A2(n28534), .A3(n29030), .ZN(n269) );
  NAND3_X1 U475 ( .A1(n31240), .A2(n24365), .A3(n24366), .ZN(n6117) );
  NAND2_X1 U476 ( .A1(n5496), .A2(n32410), .ZN(n32413) );
  NAND3_X1 U482 ( .A1(n3539), .A2(n3540), .A3(n27), .ZN(n49809) );
  XNOR2_X2 U486 ( .A(n18822), .B(n2263), .ZN(n18823) );
  NAND3_X1 U490 ( .A1(n12582), .A2(n14955), .A3(n12581), .ZN(n12588) );
  OAI21_X1 U495 ( .B1(n2899), .B2(n4259), .A(n42809), .ZN(n30) );
  OR2_X2 U496 ( .A1(n45228), .A2(n45227), .ZN(n45711) );
  AND3_X1 U500 ( .A1(n31194), .A2(n31990), .A3(n7897), .ZN(n31999) );
  XNOR2_X1 U501 ( .A(n31), .B(n47627), .ZN(Plaintext[11]) );
  NAND4_X1 U502 ( .A1(n47626), .A2(n47624), .A3(n47625), .A4(n47623), .ZN(n31)
         );
  NAND2_X1 U503 ( .A1(n11881), .A2(n32), .ZN(n11883) );
  OAI211_X1 U506 ( .C1(n28469), .C2(n32172), .A(n51628), .B(n51629), .ZN(
        n28470) );
  XNOR2_X1 U515 ( .A(n36), .B(n50532), .ZN(Plaintext[159]) );
  NAND3_X1 U516 ( .A1(n7468), .A2(n50531), .A3(n7467), .ZN(n36) );
  NAND3_X1 U522 ( .A1(n36132), .A2(n38589), .A3(n52104), .ZN(n37582) );
  NAND2_X1 U524 ( .A1(n38), .A2(n22828), .ZN(n22839) );
  OAI22_X1 U525 ( .A1(n22824), .A2(n22825), .B1(n22827), .B2(n22826), .ZN(n38)
         );
  NAND2_X1 U530 ( .A1(n3882), .A2(n11663), .ZN(n7184) );
  XNOR2_X2 U534 ( .A(n39), .B(n33668), .ZN(n38142) );
  XNOR2_X1 U535 ( .A(n33539), .B(n31842), .ZN(n39) );
  NAND2_X1 U536 ( .A1(n40), .A2(n20422), .ZN(n19330) );
  XNOR2_X2 U537 ( .A(n291), .B(n17817), .ZN(n20422) );
  INV_X1 U538 ( .A(n17838), .ZN(n40) );
  INV_X1 U539 ( .A(n5073), .ZN(n39585) );
  AND3_X2 U544 ( .A1(n12320), .A2(n8561), .A3(n8415), .ZN(n14709) );
  XNOR2_X1 U545 ( .A(n41), .B(n17189), .ZN(n17193) );
  XNOR2_X1 U546 ( .A(n17187), .B(n17188), .ZN(n41) );
  NAND3_X1 U547 ( .A1(n37460), .A2(n40585), .A3(n40775), .ZN(n5421) );
  NAND2_X1 U548 ( .A1(n727), .A2(n30452), .ZN(n1926) );
  AND4_X2 U553 ( .A1(n29476), .A2(n29477), .A3(n29475), .A4(n3388), .ZN(n31067) );
  NAND3_X1 U554 ( .A1(n51158), .A2(n42), .A3(n7321), .ZN(n146) );
  INV_X1 U556 ( .A(n32852), .ZN(n30495) );
  NAND2_X1 U557 ( .A1(n32843), .A2(n32386), .ZN(n32852) );
  NAND2_X1 U561 ( .A1(n3308), .A2(n24343), .ZN(n28291) );
  INV_X2 U562 ( .A(n29677), .ZN(n32509) );
  NAND3_X1 U564 ( .A1(n24335), .A2(n457), .A3(n24334), .ZN(n24341) );
  NAND2_X1 U565 ( .A1(n24332), .A2(n23531), .ZN(n24334) );
  NAND3_X1 U573 ( .A1(n13289), .A2(n13288), .A3(n46), .ZN(n13294) );
  NAND3_X1 U574 ( .A1(n13308), .A2(n14034), .A3(n47), .ZN(n46) );
  OR3_X1 U575 ( .A1(n36233), .A2(n35457), .A3(n37591), .ZN(n33784) );
  AND3_X1 U578 ( .A1(n48), .A2(n47887), .A3(n47888), .ZN(n4031) );
  AOI22_X1 U579 ( .A1(n47865), .A2(n47883), .B1(n47866), .B2(n47867), .ZN(n48)
         );
  NAND3_X1 U583 ( .A1(n3826), .A2(n5057), .A3(n28862), .ZN(n28509) );
  NAND2_X1 U586 ( .A1(n51), .A2(n49), .ZN(n18058) );
  NAND2_X1 U587 ( .A1(n20430), .A2(n50), .ZN(n49) );
  NAND2_X1 U588 ( .A1(n52), .A2(n20343), .ZN(n51) );
  NAND2_X1 U589 ( .A1(n20425), .A2(n20345), .ZN(n52) );
  OR2_X2 U590 ( .A1(n17838), .A2(n20422), .ZN(n20354) );
  XNOR2_X2 U593 ( .A(n5777), .B(n3524), .ZN(n36807) );
  XNOR2_X2 U596 ( .A(n23390), .B(n23391), .ZN(n2774) );
  XNOR2_X1 U597 ( .A(n54), .B(n48091), .ZN(Plaintext[41]) );
  NAND4_X1 U598 ( .A1(n48090), .A2(n48087), .A3(n48089), .A4(n48088), .ZN(n54)
         );
  NAND2_X1 U603 ( .A1(n7704), .A2(n40651), .ZN(n7414) );
  AND2_X1 U604 ( .A1(n12266), .A2(n10741), .ZN(n12242) );
  NAND2_X1 U606 ( .A1(n26455), .A2(n3160), .ZN(n28194) );
  NAND2_X1 U607 ( .A1(n39705), .A2(n55), .ZN(n41076) );
  NAND2_X1 U612 ( .A1(n56), .A2(n37975), .ZN(n4034) );
  NAND2_X1 U613 ( .A1(n1144), .A2(n36082), .ZN(n56) );
  NAND2_X1 U615 ( .A1(n40723), .A2(n674), .ZN(n1561) );
  NAND2_X1 U616 ( .A1(n41328), .A2(n41332), .ZN(n674) );
  NAND3_X1 U617 ( .A1(n31141), .A2(n8677), .A3(n29989), .ZN(n8676) );
  OAI22_X1 U621 ( .A1(n287), .A2(n32178), .B1(n32181), .B2(n32180), .ZN(n32191) );
  NAND4_X2 U623 ( .A1(n19557), .A2(n19556), .A3(n3271), .A4(n19558), .ZN(
        n26044) );
  NAND2_X1 U627 ( .A1(n18086), .A2(n1517), .ZN(n1516) );
  NAND2_X1 U631 ( .A1(n57), .A2(n10314), .ZN(n10315) );
  NAND2_X1 U632 ( .A1(n818), .A2(n10312), .ZN(n57) );
  NAND3_X1 U634 ( .A1(n867), .A2(n14739), .A3(n866), .ZN(n14749) );
  NAND3_X1 U638 ( .A1(n41728), .A2(n41730), .A3(n58), .ZN(n40475) );
  NAND2_X1 U639 ( .A1(n22503), .A2(n22502), .ZN(n5459) );
  NAND2_X1 U640 ( .A1(n12694), .A2(n12710), .ZN(n12701) );
  OR2_X1 U642 ( .A1(n12695), .A2(n12690), .ZN(n12694) );
  NAND3_X1 U645 ( .A1(n20387), .A2(n18002), .A3(n19370), .ZN(n19377) );
  NAND2_X1 U646 ( .A1(n51130), .A2(n19370), .ZN(n20387) );
  XNOR2_X1 U648 ( .A(n15846), .B(n60), .ZN(n15848) );
  XNOR2_X1 U649 ( .A(n15844), .B(n7115), .ZN(n60) );
  NAND3_X1 U650 ( .A1(n3084), .A2(n5188), .A3(n14964), .ZN(n3083) );
  OR2_X1 U651 ( .A1(n14950), .A2(n14962), .ZN(n14936) );
  NAND2_X1 U655 ( .A1(n9808), .A2(n10214), .ZN(n9809) );
  AND4_X2 U659 ( .A1(n17010), .A2(n17009), .A3(n17011), .A4(n21086), .ZN(n7350) );
  AOI21_X1 U660 ( .B1(n15902), .B2(n20232), .A(n51624), .ZN(n15920) );
  NAND2_X1 U663 ( .A1(n507), .A2(n40121), .ZN(n40194) );
  NAND2_X1 U666 ( .A1(n8625), .A2(n39381), .ZN(n37037) );
  NAND2_X1 U667 ( .A1(n26818), .A2(n27575), .ZN(n4156) );
  INV_X1 U668 ( .A(n36572), .ZN(n36481) );
  AND2_X1 U669 ( .A1(n36572), .A2(n63), .ZN(n36018) );
  NAND3_X1 U674 ( .A1(n12672), .A2(n11870), .A3(n7354), .ZN(n12450) );
  NAND2_X1 U678 ( .A1(n65), .A2(n64), .ZN(n12895) );
  OAI22_X1 U679 ( .A1(n12891), .A2(n483), .B1(n13441), .B2(n4383), .ZN(n65) );
  XNOR2_X2 U680 ( .A(n6448), .B(n6447), .ZN(n27690) );
  INV_X2 U685 ( .A(n47435), .ZN(n48730) );
  OR2_X2 U686 ( .A1(n46410), .A2(n46409), .ZN(n47435) );
  OR2_X2 U689 ( .A1(n6721), .A2(n20658), .ZN(n18846) );
  NAND2_X1 U690 ( .A1(n35732), .A2(n34628), .ZN(n6638) );
  NAND2_X1 U691 ( .A1(n40261), .A2(n42749), .ZN(n42142) );
  XNOR2_X1 U697 ( .A(n17321), .B(n18540), .ZN(n15851) );
  NAND4_X2 U698 ( .A1(n13810), .A2(n13809), .A3(n13808), .A4(n13807), .ZN(
        n17321) );
  NAND4_X2 U701 ( .A1(n67), .A2(n39658), .A3(n39656), .A4(n39657), .ZN(n43155)
         );
  NAND2_X1 U702 ( .A1(n39655), .A2(n40154), .ZN(n67) );
  NAND3_X1 U703 ( .A1(n31706), .A2(n31700), .A3(n26349), .ZN(n32122) );
  AND2_X1 U704 ( .A1(n32923), .A2(n28824), .ZN(n212) );
  NAND2_X1 U709 ( .A1(n46766), .A2(n46767), .ZN(n46769) );
  NAND3_X1 U710 ( .A1(n3690), .A2(n20923), .A3(n20922), .ZN(n20924) );
  NAND2_X1 U711 ( .A1(n48505), .A2(n46474), .ZN(n46313) );
  OR2_X1 U713 ( .A1(n35923), .A2(n37745), .ZN(n37500) );
  XNOR2_X2 U719 ( .A(n32748), .B(n32747), .ZN(n38565) );
  AND3_X2 U720 ( .A1(n29858), .A2(n7943), .A3(n70), .ZN(n32345) );
  INV_X1 U721 ( .A(n7414), .ZN(n41441) );
  NAND2_X1 U722 ( .A1(n71), .A2(n40643), .ZN(n36390) );
  NAND2_X1 U723 ( .A1(n39767), .A2(n7414), .ZN(n71) );
  OAI22_X1 U727 ( .A1(n27796), .A2(n27795), .B1(n27797), .B2(n28618), .ZN(
        n3007) );
  OAI21_X1 U730 ( .B1(n29379), .B2(n30575), .A(n73), .ZN(n29380) );
  NAND3_X1 U731 ( .A1(n31034), .A2(n6107), .A3(n31827), .ZN(n73) );
  XNOR2_X1 U733 ( .A(n6856), .B(n6858), .ZN(n74) );
  NAND3_X1 U734 ( .A1(n29448), .A2(n29446), .A3(n29447), .ZN(n29449) );
  OR3_X1 U736 ( .A1(n40591), .A2(n431), .A3(n40768), .ZN(n7861) );
  NAND2_X1 U737 ( .A1(n4047), .A2(n22409), .ZN(n22414) );
  NAND2_X1 U738 ( .A1(n7316), .A2(n7315), .ZN(n7314) );
  NAND4_X2 U742 ( .A1(n6891), .A2(n6890), .A3(n29689), .A4(n6893), .ZN(n35482)
         );
  NAND2_X1 U749 ( .A1(n22861), .A2(n22856), .ZN(n22865) );
  NAND2_X1 U751 ( .A1(n6639), .A2(n7059), .ZN(n7057) );
  NAND3_X1 U752 ( .A1(n49532), .A2(n49533), .A3(n49531), .ZN(n49546) );
  INV_X1 U754 ( .A(n11647), .ZN(n10013) );
  NAND2_X1 U755 ( .A1(n9305), .A2(n10572), .ZN(n11647) );
  NAND2_X1 U756 ( .A1(n13301), .A2(n4634), .ZN(n13302) );
  NAND2_X1 U760 ( .A1(n77), .A2(n76), .ZN(n2832) );
  INV_X1 U761 ( .A(n19390), .ZN(n77) );
  NOR2_X1 U764 ( .A1(n20448), .A2(n21480), .ZN(n20817) );
  AND3_X2 U769 ( .A1(n43473), .A2(n43472), .A3(n43471), .ZN(n43490) );
  OR2_X2 U771 ( .A1(n2831), .A2(n19394), .ZN(n23020) );
  NAND3_X1 U772 ( .A1(n3969), .A2(n19329), .A3(n3970), .ZN(n19334) );
  NAND2_X2 U775 ( .A1(n51094), .A2(n42990), .ZN(n49725) );
  OR2_X2 U781 ( .A1(n1465), .A2(n3071), .ZN(n42136) );
  OR2_X2 U782 ( .A1(n29325), .A2(n52216), .ZN(n29315) );
  INV_X1 U783 ( .A(n34698), .ZN(n34699) );
  NAND2_X1 U785 ( .A1(n26416), .A2(n28915), .ZN(n28571) );
  NAND2_X1 U786 ( .A1(n981), .A2(n27069), .ZN(n2669) );
  NAND3_X1 U788 ( .A1(n45889), .A2(n45890), .A3(n45888), .ZN(n45891) );
  BUF_X2 U797 ( .A(n18535), .Z(n461) );
  NAND2_X1 U799 ( .A1(n20161), .A2(n23409), .ZN(n22046) );
  XNOR2_X1 U801 ( .A(n36832), .B(n82), .ZN(n1892) );
  XNOR2_X2 U803 ( .A(n26412), .B(n83), .ZN(n28923) );
  NOR2_X1 U807 ( .A1(n21144), .A2(n21755), .ZN(n21730) );
  NAND2_X2 U809 ( .A1(n6304), .A2(n6306), .ZN(n34400) );
  NAND2_X1 U810 ( .A1(n19075), .A2(n19076), .ZN(n20131) );
  OAI211_X1 U813 ( .C1(n46731), .C2(n45799), .A(n45801), .B(n86), .ZN(n45806)
         );
  NAND2_X1 U816 ( .A1(n52120), .A2(n40943), .ZN(n41553) );
  NAND2_X1 U818 ( .A1(n21439), .A2(n21427), .ZN(n19950) );
  NAND3_X1 U819 ( .A1(n14795), .A2(n14139), .A3(n14788), .ZN(n5139) );
  XNOR2_X1 U820 ( .A(n87), .B(n48719), .ZN(Plaintext[65]) );
  NAND2_X1 U822 ( .A1(n14600), .A2(n14601), .ZN(n13317) );
  NAND2_X1 U823 ( .A1(n10391), .A2(n11400), .ZN(n9607) );
  INV_X1 U824 ( .A(n30043), .ZN(n1158) );
  NAND2_X1 U825 ( .A1(n29602), .A2(n31340), .ZN(n30043) );
  NAND2_X1 U826 ( .A1(n19348), .A2(n20506), .ZN(n19349) );
  OAI21_X1 U827 ( .B1(n12271), .B2(n8994), .A(n11335), .ZN(n8993) );
  NAND2_X1 U828 ( .A1(n11346), .A2(n8994), .ZN(n11335) );
  NAND2_X1 U831 ( .A1(n39271), .A2(n39284), .ZN(n39275) );
  NAND2_X1 U835 ( .A1(n2151), .A2(n14950), .ZN(n15286) );
  NAND3_X1 U837 ( .A1(n2613), .A2(n49611), .A3(n49602), .ZN(n6009) );
  NAND4_X2 U839 ( .A1(n19041), .A2(n19040), .A3(n19042), .A4(n19043), .ZN(
        n25548) );
  NAND3_X2 U842 ( .A1(n1358), .A2(n40347), .A3(n40345), .ZN(n1357) );
  NAND4_X2 U844 ( .A1(n3884), .A2(n7782), .A3(n26748), .A4(n26749), .ZN(n31684) );
  NAND3_X1 U848 ( .A1(n273), .A2(n4581), .A3(n47582), .ZN(n272) );
  XNOR2_X2 U851 ( .A(n3710), .B(n14508), .ZN(n19250) );
  NOR2_X1 U854 ( .A1(n89), .A2(n22106), .ZN(n22112) );
  OAI22_X1 U855 ( .A1(n22104), .A2(n22103), .B1(n6103), .B2(n22102), .ZN(n89)
         );
  AND2_X2 U857 ( .A1(n39014), .A2(n39007), .ZN(n39259) );
  AND2_X2 U858 ( .A1(n2166), .A2(n590), .ZN(n20015) );
  XNOR2_X1 U862 ( .A(n26123), .B(n90), .ZN(n26128) );
  XNOR2_X1 U863 ( .A(n26520), .B(n26122), .ZN(n90) );
  NAND2_X1 U864 ( .A1(n50299), .A2(n51300), .ZN(n50301) );
  NAND2_X1 U867 ( .A1(n1941), .A2(n20592), .ZN(n1940) );
  XNOR2_X2 U873 ( .A(n34150), .B(n34149), .ZN(n36557) );
  NAND4_X1 U874 ( .A1(n91), .A2(n21882), .A3(n21883), .A4(n21881), .ZN(n21893)
         );
  NAND4_X1 U878 ( .A1(n20179), .A2(n20180), .A3(n20182), .A4(n20181), .ZN(n92)
         );
  XNOR2_X1 U879 ( .A(n35085), .B(n35224), .ZN(n7611) );
  NAND3_X1 U882 ( .A1(n41009), .A2(n40801), .A3(n38763), .ZN(n8264) );
  NAND2_X1 U883 ( .A1(n30709), .A2(n29855), .ZN(n28799) );
  NAND2_X1 U887 ( .A1(n50232), .A2(n93), .ZN(n50168) );
  NAND2_X1 U890 ( .A1(n525), .A2(n36272), .ZN(n3163) );
  NAND2_X1 U891 ( .A1(n27736), .A2(n27730), .ZN(n27726) );
  INV_X1 U898 ( .A(n47085), .ZN(n6565) );
  NAND2_X1 U899 ( .A1(n34528), .A2(n2788), .ZN(n37617) );
  NAND3_X1 U901 ( .A1(n5753), .A2(n32494), .A3(n5751), .ZN(n32801) );
  NAND3_X2 U902 ( .A1(n38296), .A2(n38295), .A3(n38294), .ZN(n40869) );
  OAI21_X1 U905 ( .B1(n39744), .B2(n5747), .A(n7662), .ZN(n39750) );
  AND3_X1 U906 ( .A1(n29483), .A2(n29502), .A3(n29484), .ZN(n95) );
  NAND3_X1 U911 ( .A1(n4794), .A2(n13351), .A3(n51152), .ZN(n13360) );
  NAND2_X1 U917 ( .A1(n8200), .A2(n39941), .ZN(n39961) );
  NAND2_X1 U918 ( .A1(n19797), .A2(n5388), .ZN(n3604) );
  NAND2_X1 U919 ( .A1(n18888), .A2(n19795), .ZN(n5388) );
  INV_X1 U922 ( .A(n10686), .ZN(n12383) );
  NAND2_X1 U923 ( .A1(n26661), .A2(n28701), .ZN(n29303) );
  NAND2_X1 U927 ( .A1(n51340), .A2(n47599), .ZN(n47618) );
  NAND3_X1 U928 ( .A1(n28896), .A2(n28897), .A3(n28898), .ZN(n28899) );
  OR2_X2 U931 ( .A1(n1170), .A2(n99), .ZN(n26378) );
  NAND4_X1 U932 ( .A1(n5035), .A2(n5034), .A3(n23031), .A4(n23030), .ZN(n99)
         );
  NAND2_X1 U933 ( .A1(n100), .A2(n50520), .ZN(n7468) );
  NAND3_X1 U937 ( .A1(n30637), .A2(n30636), .A3(n2496), .ZN(n4135) );
  NAND3_X1 U939 ( .A1(n3407), .A2(n26079), .A3(n26080), .ZN(n26082) );
  XNOR2_X1 U940 ( .A(n101), .B(n44638), .ZN(Plaintext[169]) );
  NAND4_X1 U941 ( .A1(n44637), .A2(n44635), .A3(n44636), .A4(n44634), .ZN(n101) );
  NAND3_X1 U942 ( .A1(n29973), .A2(n26347), .A3(n32138), .ZN(n26351) );
  NAND2_X1 U944 ( .A1(n7222), .A2(n22189), .ZN(n20563) );
  NAND2_X1 U946 ( .A1(n1092), .A2(n16039), .ZN(n13034) );
  NAND3_X1 U947 ( .A1(n2928), .A2(n26088), .A3(n26087), .ZN(n26203) );
  NAND2_X1 U948 ( .A1(n102), .A2(n29139), .ZN(n27087) );
  NAND3_X1 U951 ( .A1(n18330), .A2(n18342), .A3(n18074), .ZN(n18329) );
  AND2_X2 U952 ( .A1(n3073), .A2(n18331), .ZN(n18330) );
  NAND2_X1 U953 ( .A1(n1031), .A2(n45960), .ZN(n1339) );
  NAND2_X1 U956 ( .A1(n790), .A2(n4540), .ZN(n806) );
  INV_X2 U973 ( .A(n15324), .ZN(n15435) );
  AOI21_X1 U976 ( .B1(n32816), .B2(n32823), .A(n106), .ZN(n8749) );
  NAND3_X1 U977 ( .A1(n32814), .A2(n8536), .A3(n51630), .ZN(n106) );
  NAND2_X1 U983 ( .A1(n19538), .A2(n19539), .ZN(n19541) );
  NAND2_X1 U987 ( .A1(n45958), .A2(n49677), .ZN(n50025) );
  XNOR2_X2 U989 ( .A(n16707), .B(n16475), .ZN(n20157) );
  NAND3_X2 U990 ( .A1(n4285), .A2(n9882), .A3(n9880), .ZN(n13930) );
  NAND2_X1 U991 ( .A1(n110), .A2(n108), .ZN(n47471) );
  NAND3_X1 U992 ( .A1(n6604), .A2(n8448), .A3(n6831), .ZN(n108) );
  NAND2_X1 U993 ( .A1(n47469), .A2(n47617), .ZN(n110) );
  NAND2_X1 U994 ( .A1(n32335), .A2(n2091), .ZN(n32699) );
  NAND2_X1 U995 ( .A1(n32684), .A2(n32691), .ZN(n32335) );
  NAND3_X1 U996 ( .A1(n47771), .A2(n47786), .A3(n47755), .ZN(n45007) );
  NAND3_X1 U1003 ( .A1(n45523), .A2(n45533), .A3(n113), .ZN(n112) );
  INV_X1 U1004 ( .A(n45816), .ZN(n113) );
  XNOR2_X1 U1006 ( .A(n114), .B(n41963), .ZN(n41967) );
  XNOR2_X1 U1007 ( .A(n41964), .B(n42962), .ZN(n114) );
  NAND3_X1 U1008 ( .A1(n2963), .A2(n24146), .A3(n4025), .ZN(n7076) );
  NAND4_X2 U1009 ( .A1(n8745), .A2(n31571), .A3(n31572), .A4(n115), .ZN(n36855) );
  NAND3_X1 U1010 ( .A1(n1890), .A2(n31568), .A3(n31569), .ZN(n115) );
  XNOR2_X2 U1011 ( .A(n26611), .B(n25778), .ZN(n27479) );
  NOR2_X2 U1012 ( .A1(n23517), .A2(n23516), .ZN(n26611) );
  AOI22_X1 U1013 ( .A1(n15835), .A2(n20657), .B1(n15836), .B2(n20655), .ZN(
        n15838) );
  NOR2_X1 U1014 ( .A1(n9952), .A2(n10555), .ZN(n9829) );
  NOR2_X1 U1021 ( .A1(n24126), .A2(n118), .ZN(n4148) );
  NAND2_X1 U1022 ( .A1(n190), .A2(n119), .ZN(n118) );
  INV_X1 U1023 ( .A(n120), .ZN(n5675) );
  OAI21_X1 U1024 ( .B1(n3290), .B2(n41491), .A(n36287), .ZN(n120) );
  NAND3_X1 U1026 ( .A1(n21768), .A2(n21766), .A3(n819), .ZN(n21790) );
  NAND2_X1 U1027 ( .A1(n4314), .A2(n4315), .ZN(n21768) );
  NAND2_X2 U1028 ( .A1(n1700), .A2(n1699), .ZN(n36930) );
  NAND3_X1 U1032 ( .A1(n35900), .A2(n38640), .A3(n37682), .ZN(n35903) );
  NAND2_X1 U1033 ( .A1(n51736), .A2(n39225), .ZN(n39233) );
  NAND3_X1 U1034 ( .A1(n121), .A2(n37913), .A3(n37914), .ZN(n8553) );
  NAND2_X1 U1035 ( .A1(n4675), .A2(n4674), .ZN(n121) );
  NAND2_X1 U1036 ( .A1(n1874), .A2(n39906), .ZN(n39902) );
  NAND3_X1 U1038 ( .A1(n48939), .A2(n48940), .A3(n48938), .ZN(n48948) );
  NAND3_X2 U1042 ( .A1(n901), .A2(n30467), .A3(n30465), .ZN(n900) );
  NOR2_X1 U1043 ( .A1(n48952), .A2(n48950), .ZN(n48934) );
  NAND2_X1 U1044 ( .A1(n52137), .A2(n48944), .ZN(n48952) );
  NAND2_X1 U1047 ( .A1(n745), .A2(n51489), .ZN(n29754) );
  NAND2_X1 U1049 ( .A1(n51103), .A2(n32214), .ZN(n32199) );
  OAI211_X2 U1055 ( .C1(n18297), .C2(n18298), .A(n18296), .B(n18295), .ZN(
        n22121) );
  OAI211_X1 U1056 ( .C1(n46957), .C2(n46956), .A(n126), .B(n125), .ZN(n46959)
         );
  NAND2_X1 U1057 ( .A1(n46954), .A2(n3198), .ZN(n125) );
  AOI21_X1 U1058 ( .B1(n46954), .B2(n46953), .A(n51478), .ZN(n126) );
  NAND2_X1 U1059 ( .A1(n44109), .A2(n46830), .ZN(n46772) );
  NAND3_X2 U1061 ( .A1(n23544), .A2(n6917), .A3(n23543), .ZN(n26435) );
  NAND4_X2 U1062 ( .A1(n5803), .A2(n11911), .A3(n127), .A4(n8665), .ZN(n15440)
         );
  NOR2_X1 U1064 ( .A1(n129), .A2(n128), .ZN(n13911) );
  NAND2_X1 U1066 ( .A1(n1657), .A2(n23044), .ZN(n22087) );
  NAND2_X1 U1067 ( .A1(n10475), .A2(n12589), .ZN(n10477) );
  INV_X1 U1068 ( .A(n32119), .ZN(n31705) );
  NAND2_X1 U1069 ( .A1(n32119), .A2(n32130), .ZN(n5305) );
  NAND2_X1 U1073 ( .A1(n3951), .A2(n30549), .ZN(n28724) );
  NAND3_X1 U1074 ( .A1(n36401), .A2(n37647), .A3(n36410), .ZN(n35726) );
  OR2_X2 U1079 ( .A1(n42177), .A2(n44640), .ZN(n45533) );
  NAND3_X2 U1081 ( .A1(n4084), .A2(n31951), .A3(n4085), .ZN(n36792) );
  BUF_X1 U1082 ( .A(n37158), .Z(n37927) );
  BUF_X1 U1083 ( .A(n19214), .Z(n2180) );
  NAND2_X1 U1090 ( .A1(n27852), .A2(n29478), .ZN(n26667) );
  INV_X2 U1091 ( .A(n11740), .ZN(n14482) );
  NAND3_X1 U1092 ( .A1(n38720), .A2(n39300), .A3(n39293), .ZN(n39312) );
  NAND3_X1 U1093 ( .A1(n50545), .A2(n50544), .A3(n50549), .ZN(n50547) );
  XNOR2_X2 U1095 ( .A(n43909), .B(n44198), .ZN(n2051) );
  NAND3_X1 U1101 ( .A1(n46980), .A2(n46981), .A3(n134), .ZN(n46988) );
  NAND2_X1 U1109 ( .A1(n41150), .A2(n135), .ZN(n39839) );
  NAND4_X2 U1111 ( .A1(n32148), .A2(n32147), .A3(n32145), .A4(n32146), .ZN(
        n41150) );
  NAND2_X1 U1112 ( .A1(n30855), .A2(n30856), .ZN(n706) );
  XNOR2_X2 U1113 ( .A(n31620), .B(n31619), .ZN(n38057) );
  NOR2_X2 U1115 ( .A1(n17418), .A2(n17420), .ZN(n24206) );
  NAND3_X1 U1116 ( .A1(n47546), .A2(n47545), .A3(n51346), .ZN(n47549) );
  XNOR2_X2 U1117 ( .A(n136), .B(n8512), .ZN(n19396) );
  XNOR2_X1 U1118 ( .A(n10658), .B(n10657), .ZN(n136) );
  XNOR2_X1 U1124 ( .A(n137), .B(n50503), .ZN(Plaintext[157]) );
  NAND4_X1 U1125 ( .A1(n7471), .A2(n7472), .A3(n7473), .A4(n2446), .ZN(n137)
         );
  NOR2_X1 U1126 ( .A1(n139), .A2(n51636), .ZN(n46170) );
  NAND2_X1 U1128 ( .A1(n46811), .A2(n46822), .ZN(n46784) );
  AOI21_X1 U1132 ( .B1(n41132), .B2(n141), .A(n41131), .ZN(n41140) );
  NAND3_X1 U1133 ( .A1(n44421), .A2(n44424), .A3(n3449), .ZN(n141) );
  NAND4_X2 U1138 ( .A1(n6362), .A2(n143), .A3(n142), .A4(n26680), .ZN(n31815)
         );
  NAND2_X1 U1139 ( .A1(n26672), .A2(n26671), .ZN(n142) );
  NAND2_X1 U1140 ( .A1(n26673), .A2(n29495), .ZN(n143) );
  NAND3_X1 U1146 ( .A1(n6629), .A2(n21655), .A3(n20659), .ZN(n6628) );
  NAND3_X1 U1147 ( .A1(n14954), .A2(n14952), .A3(n14953), .ZN(n14964) );
  NAND3_X1 U1148 ( .A1(n39169), .A2(n38667), .A3(n7729), .ZN(n38658) );
  BUF_X2 U1149 ( .A(n10881), .Z(n13525) );
  OR2_X2 U1151 ( .A1(n25479), .A2(n29182), .ZN(n29270) );
  XNOR2_X1 U1152 ( .A(n144), .B(n32265), .ZN(n33213) );
  XNOR2_X1 U1153 ( .A(n32223), .B(n32224), .ZN(n144) );
  NAND3_X1 U1155 ( .A1(n30598), .A2(n30599), .A3(n30597), .ZN(n30600) );
  INV_X1 U1157 ( .A(n49691), .ZN(n49692) );
  NAND2_X1 U1158 ( .A1(n2668), .A2(n145), .ZN(n49691) );
  NAND3_X2 U1159 ( .A1(n148), .A2(n37744), .A3(n147), .ZN(n41770) );
  NAND2_X1 U1160 ( .A1(n37738), .A2(n37737), .ZN(n147) );
  XNOR2_X2 U1162 ( .A(n32337), .B(n5045), .ZN(n6826) );
  NAND2_X2 U1163 ( .A1(n17018), .A2(n20157), .ZN(n20124) );
  NAND3_X2 U1164 ( .A1(n149), .A2(n30615), .A3(n30613), .ZN(n37113) );
  NAND2_X1 U1167 ( .A1(n30604), .A2(n30603), .ZN(n151) );
  XNOR2_X2 U1170 ( .A(n3924), .B(n33324), .ZN(n37759) );
  NAND2_X1 U1173 ( .A1(n10858), .A2(n14123), .ZN(n14128) );
  NAND2_X1 U1177 ( .A1(n7984), .A2(n1901), .ZN(n1900) );
  INV_X1 U1181 ( .A(n155), .ZN(n154) );
  OAI21_X1 U1182 ( .B1(n11088), .B2(n11087), .A(n11085), .ZN(n155) );
  NAND3_X1 U1187 ( .A1(n709), .A2(n32487), .A3(n32486), .ZN(n157) );
  AND2_X2 U1189 ( .A1(n30758), .A2(n24351), .ZN(n6048) );
  NAND2_X1 U1190 ( .A1(n28823), .A2(n158), .ZN(n32923) );
  NAND2_X1 U1195 ( .A1(n161), .A2(n30785), .ZN(n160) );
  AOI21_X1 U1197 ( .B1(n11008), .B2(n10199), .A(n9748), .ZN(n9037) );
  AND2_X2 U1200 ( .A1(n754), .A2(n23950), .ZN(n23963) );
  XNOR2_X2 U1201 ( .A(n26367), .B(n26366), .ZN(n28926) );
  NAND2_X1 U1203 ( .A1(n21297), .A2(n21296), .ZN(n162) );
  NAND3_X1 U1205 ( .A1(n49703), .A2(n164), .A3(n163), .ZN(n6906) );
  INV_X1 U1206 ( .A(n44748), .ZN(n163) );
  INV_X1 U1207 ( .A(n44747), .ZN(n164) );
  NAND2_X1 U1209 ( .A1(n166), .A2(n2083), .ZN(n22484) );
  NAND2_X1 U1210 ( .A1(n22476), .A2(n22480), .ZN(n166) );
  OR2_X2 U1212 ( .A1(n19806), .A2(n19801), .ZN(n21300) );
  NAND2_X1 U1213 ( .A1(n31269), .A2(n31490), .ZN(n169) );
  NAND2_X1 U1214 ( .A1(n5913), .A2(n31489), .ZN(n29840) );
  NAND2_X1 U1215 ( .A1(n23707), .A2(n171), .ZN(n170) );
  OR2_X1 U1217 ( .A1(n29622), .A2(n29616), .ZN(n30506) );
  NAND2_X1 U1219 ( .A1(n47926), .A2(n47927), .ZN(n172) );
  NAND2_X1 U1220 ( .A1(n47960), .A2(n52056), .ZN(n174) );
  NAND3_X1 U1221 ( .A1(n47672), .A2(n47670), .A3(n47671), .ZN(n47678) );
  NAND2_X1 U1223 ( .A1(n6619), .A2(n50675), .ZN(n6618) );
  NOR2_X1 U1224 ( .A1(n51631), .A2(n175), .ZN(n3114) );
  NAND2_X1 U1227 ( .A1(n27129), .A2(n177), .ZN(n28584) );
  NAND2_X1 U1230 ( .A1(n1070), .A2(n5073), .ZN(n1069) );
  NAND3_X1 U1232 ( .A1(n20710), .A2(n20709), .A3(n51626), .ZN(n20719) );
  XNOR2_X1 U1234 ( .A(n180), .B(n50817), .ZN(Plaintext[178]) );
  NAND4_X1 U1235 ( .A1(n50816), .A2(n50813), .A3(n50815), .A4(n50814), .ZN(
        n180) );
  NOR2_X1 U1236 ( .A1(n28857), .A2(n28784), .ZN(n28786) );
  NAND4_X1 U1237 ( .A1(n5390), .A2(n29060), .A3(n745), .A4(n28783), .ZN(n28857) );
  NAND2_X1 U1238 ( .A1(n181), .A2(n9432), .ZN(n5513) );
  NAND2_X1 U1239 ( .A1(n11418), .A2(n9431), .ZN(n181) );
  NAND2_X1 U1246 ( .A1(n31205), .A2(n32491), .ZN(n27647) );
  NAND3_X2 U1248 ( .A1(n1996), .A2(n21088), .A3(n1995), .ZN(n24905) );
  NAND2_X1 U1249 ( .A1(n28177), .A2(n28187), .ZN(n29719) );
  XNOR2_X2 U1250 ( .A(n2596), .B(n28367), .ZN(n28187) );
  AND2_X2 U1253 ( .A1(n28867), .A2(n2707), .ZN(n28952) );
  NAND3_X1 U1254 ( .A1(n22277), .A2(n23551), .A3(n23562), .ZN(n22278) );
  OAI211_X1 U1258 ( .C1(n20424), .C2(n20425), .A(n20432), .B(n20423), .ZN(
        n20440) );
  NAND4_X1 U1265 ( .A1(n183), .A2(n9554), .A3(n9552), .A4(n9553), .ZN(n9556)
         );
  NAND2_X1 U1266 ( .A1(n11128), .A2(n9547), .ZN(n183) );
  NAND3_X1 U1267 ( .A1(n7511), .A2(n21914), .A3(n21916), .ZN(n21917) );
  AND3_X2 U1268 ( .A1(n46365), .A2(n46364), .A3(n46366), .ZN(n47442) );
  NAND3_X1 U1269 ( .A1(n184), .A2(n37538), .A3(n3165), .ZN(n37540) );
  NAND2_X1 U1270 ( .A1(n3163), .A2(n37396), .ZN(n184) );
  NAND2_X1 U1271 ( .A1(n12590), .A2(n11920), .ZN(n9540) );
  NAND2_X1 U1275 ( .A1(n40681), .A2(n185), .ZN(n40699) );
  NAND2_X1 U1276 ( .A1(n40678), .A2(n40679), .ZN(n186) );
  NAND3_X1 U1278 ( .A1(n6985), .A2(n49595), .A3(n49574), .ZN(n45728) );
  BUF_X2 U1283 ( .A(n42604), .Z(n46276) );
  NAND3_X1 U1285 ( .A1(n40767), .A2(n40785), .A3(n40598), .ZN(n7105) );
  XNOR2_X1 U1286 ( .A(n188), .B(n45737), .ZN(Plaintext[121]) );
  NAND4_X1 U1287 ( .A1(n45732), .A2(n45733), .A3(n45734), .A4(n45735), .ZN(
        n188) );
  NAND4_X1 U1288 ( .A1(n24121), .A2(n4726), .A3(n24413), .A4(n24120), .ZN(n190) );
  NAND3_X1 U1295 ( .A1(n29735), .A2(n29734), .A3(n29733), .ZN(n191) );
  XNOR2_X1 U1296 ( .A(n192), .B(n28362), .ZN(n28366) );
  XNOR2_X1 U1297 ( .A(n28355), .B(n28356), .ZN(n192) );
  XNOR2_X1 U1300 ( .A(n4522), .B(n42955), .ZN(n193) );
  XNOR2_X2 U1301 ( .A(n35059), .B(n35609), .ZN(n33470) );
  NAND3_X2 U1302 ( .A1(n32515), .A2(n5121), .A3(n5159), .ZN(n35609) );
  NAND4_X1 U1305 ( .A1(n27118), .A2(n195), .A3(n24876), .A4(n194), .ZN(n4598)
         );
  NAND2_X1 U1306 ( .A1(n24859), .A2(n28545), .ZN(n194) );
  NAND2_X1 U1307 ( .A1(n197), .A2(n38630), .ZN(n38640) );
  XNOR2_X2 U1308 ( .A(n35269), .B(n35268), .ZN(n38630) );
  NAND2_X1 U1309 ( .A1(n198), .A2(n20247), .ZN(n20248) );
  NAND2_X1 U1310 ( .A1(n20245), .A2(n21629), .ZN(n198) );
  OR3_X1 U1314 ( .A1(n23518), .A2(n23129), .A3(n51001), .ZN(n24067) );
  XNOR2_X1 U1316 ( .A(n199), .B(n18652), .ZN(n7270) );
  XNOR2_X1 U1317 ( .A(n2290), .B(n18660), .ZN(n199) );
  NAND3_X2 U1318 ( .A1(n32994), .A2(n32995), .A3(n200), .ZN(n35537) );
  NAND3_X1 U1319 ( .A1(n48220), .A2(n2119), .A3(n48200), .ZN(n45000) );
  NAND4_X2 U1321 ( .A1(n201), .A2(n41808), .A3(n41805), .A4(n41806), .ZN(
        n45327) );
  NAND2_X1 U1323 ( .A1(n28025), .A2(n30305), .ZN(n28028) );
  NAND3_X1 U1325 ( .A1(n20464), .A2(n20465), .A3(n20463), .ZN(n8589) );
  NAND2_X1 U1328 ( .A1(n4819), .A2(n13927), .ZN(n17786) );
  AND2_X2 U1332 ( .A1(n27090), .A2(n27089), .ZN(n29677) );
  NAND2_X1 U1333 ( .A1(n13924), .A2(n204), .ZN(n13926) );
  NAND2_X1 U1334 ( .A1(n7735), .A2(n205), .ZN(n204) );
  NOR2_X2 U1339 ( .A1(n24025), .A2(n22101), .ZN(n23675) );
  NAND4_X1 U1340 ( .A1(n206), .A2(n11524), .A3(n11522), .A4(n11523), .ZN(
        n13914) );
  OAI21_X1 U1341 ( .B1(n11519), .B2(n11520), .A(n11567), .ZN(n206) );
  NAND3_X2 U1343 ( .A1(n8590), .A2(n20486), .A3(n8588), .ZN(n22479) );
  NAND4_X2 U1349 ( .A1(n33888), .A2(n33886), .A3(n33887), .A4(n33885), .ZN(
        n3526) );
  NAND2_X2 U1361 ( .A1(n19118), .A2(n21270), .ZN(n19122) );
  NAND3_X2 U1362 ( .A1(n208), .A2(n840), .A3(n37428), .ZN(n40768) );
  NAND2_X1 U1363 ( .A1(n4571), .A2(n38111), .ZN(n208) );
  OAI211_X1 U1364 ( .C1(n44850), .C2(n46760), .A(n209), .B(n46757), .ZN(n46761) );
  NAND2_X1 U1365 ( .A1(n46754), .A2(n44850), .ZN(n209) );
  XNOR2_X1 U1366 ( .A(n210), .B(n35788), .ZN(n35529) );
  XNOR2_X1 U1367 ( .A(n35515), .B(n35514), .ZN(n210) );
  NAND2_X1 U1368 ( .A1(n36157), .A2(n37432), .ZN(n36164) );
  AOI21_X1 U1370 ( .B1(n14764), .B2(n15237), .A(n15242), .ZN(n211) );
  INV_X1 U1374 ( .A(n32895), .ZN(n6269) );
  NAND2_X1 U1375 ( .A1(n6270), .A2(n32895), .ZN(n32919) );
  NAND3_X2 U1376 ( .A1(n28776), .A2(n28777), .A3(n28778), .ZN(n32895) );
  BUF_X2 U1377 ( .A(n11144), .Z(n15233) );
  XNOR2_X2 U1380 ( .A(Key[15]), .B(Ciphertext[86]), .ZN(n9895) );
  XNOR2_X1 U1384 ( .A(n17847), .B(n17730), .ZN(n16292) );
  NAND2_X1 U1390 ( .A1(n19891), .A2(n15630), .ZN(n18932) );
  NAND4_X1 U1393 ( .A1(n33066), .A2(n33065), .A3(n35713), .A4(n33064), .ZN(
        n216) );
  NAND4_X2 U1394 ( .A1(n22841), .A2(n22839), .A3(n22838), .A4(n22840), .ZN(
        n25947) );
  NAND3_X1 U1396 ( .A1(n11445), .A2(n6409), .A3(n51674), .ZN(n6406) );
  NAND3_X1 U1397 ( .A1(n40388), .A2(n40385), .A3(n51012), .ZN(n38620) );
  INV_X1 U1398 ( .A(n41143), .ZN(n218) );
  NAND3_X1 U1400 ( .A1(n36519), .A2(n36518), .A3(n36517), .ZN(n36520) );
  NAND2_X1 U1401 ( .A1(n37990), .A2(n37975), .ZN(n36519) );
  NAND2_X1 U1402 ( .A1(n2754), .A2(n47151), .ZN(n2708) );
  NAND2_X1 U1403 ( .A1(n47159), .A2(n47154), .ZN(n2754) );
  XNOR2_X1 U1404 ( .A(n34724), .B(n219), .ZN(n33135) );
  XNOR2_X1 U1405 ( .A(n33129), .B(n33128), .ZN(n219) );
  NAND2_X1 U1406 ( .A1(n13275), .A2(n220), .ZN(n13280) );
  AOI21_X1 U1407 ( .B1(n14763), .B2(n15199), .A(n2013), .ZN(n220) );
  NAND3_X1 U1410 ( .A1(n46344), .A2(n46274), .A3(n46354), .ZN(n46275) );
  XNOR2_X2 U1413 ( .A(n24425), .B(n24424), .ZN(n1484) );
  INV_X1 U1418 ( .A(n39288), .ZN(n222) );
  INV_X2 U1420 ( .A(n49021), .ZN(n49019) );
  NOR2_X1 U1423 ( .A1(n3997), .A2(n7786), .ZN(n265) );
  NAND3_X1 U1424 ( .A1(n3790), .A2(n30999), .A3(n29840), .ZN(n3788) );
  NAND2_X1 U1425 ( .A1(n36458), .A2(n36454), .ZN(n36462) );
  XNOR2_X2 U1426 ( .A(n34344), .B(n3926), .ZN(n36454) );
  OAI211_X1 U1428 ( .C1(n51165), .C2(n223), .A(n1095), .B(n50500), .ZN(n7471)
         );
  NAND2_X1 U1429 ( .A1(n50496), .A2(n50521), .ZN(n223) );
  OAI21_X1 U1431 ( .B1(n41979), .B2(n41975), .A(n225), .ZN(n40614) );
  NAND2_X1 U1432 ( .A1(n41981), .A2(n226), .ZN(n225) );
  NAND2_X1 U1434 ( .A1(n30161), .A2(n227), .ZN(n30317) );
  BUF_X2 U1436 ( .A(n5454), .Z(n2155) );
  NAND2_X1 U1441 ( .A1(n21480), .A2(n21494), .ZN(n20828) );
  NAND3_X1 U1444 ( .A1(n19903), .A2(n19902), .A3(n22764), .ZN(n19910) );
  NAND2_X1 U1445 ( .A1(n10184), .A2(n2093), .ZN(n10544) );
  NAND2_X1 U1446 ( .A1(n49819), .A2(n6689), .ZN(n49821) );
  NAND2_X1 U1448 ( .A1(n31804), .A2(n31805), .ZN(n7200) );
  NAND2_X1 U1450 ( .A1(n228), .A2(n32505), .ZN(n32515) );
  NOR2_X1 U1451 ( .A1(n32502), .A2(n3358), .ZN(n228) );
  NAND3_X1 U1455 ( .A1(n32389), .A2(n28914), .A3(n1140), .ZN(n28940) );
  NAND2_X1 U1459 ( .A1(n41974), .A2(n41973), .ZN(n41976) );
  XNOR2_X1 U1460 ( .A(n229), .B(n19923), .ZN(n20541) );
  XNOR2_X1 U1461 ( .A(n19628), .B(n1384), .ZN(n229) );
  XNOR2_X2 U1466 ( .A(n2578), .B(n19258), .ZN(n19891) );
  NAND3_X1 U1468 ( .A1(n13417), .A2(n10651), .A3(n10650), .ZN(n14353) );
  NAND3_X1 U1471 ( .A1(n230), .A2(n22559), .A3(n22998), .ZN(n22560) );
  NAND2_X1 U1472 ( .A1(n3691), .A2(n22557), .ZN(n230) );
  AND4_X2 U1473 ( .A1(n38308), .A2(n38307), .A3(n38306), .A4(n38309), .ZN(
        n40526) );
  OAI22_X1 U1474 ( .A1(n1574), .A2(n26974), .B1(n398), .B2(n26975), .ZN(n1572)
         );
  XNOR2_X1 U1476 ( .A(n231), .B(n25129), .ZN(n7429) );
  XNOR2_X1 U1477 ( .A(n25139), .B(n25138), .ZN(n231) );
  NAND2_X1 U1486 ( .A1(n41940), .A2(n233), .ZN(n35993) );
  NAND2_X1 U1488 ( .A1(n50027), .A2(n49650), .ZN(n49660) );
  NAND2_X1 U1490 ( .A1(n234), .A2(n4091), .ZN(n6223) );
  OAI211_X1 U1491 ( .C1(n36241), .C2(n37748), .A(n35924), .B(n37764), .ZN(n234) );
  NAND3_X1 U1492 ( .A1(n11971), .A2(n10340), .A3(n10339), .ZN(n10342) );
  NAND2_X1 U1494 ( .A1(n31783), .A2(n31782), .ZN(n31785) );
  NOR2_X1 U1496 ( .A1(n236), .A2(n235), .ZN(n7056) );
  NOR2_X1 U1497 ( .A1(n48688), .A2(n48682), .ZN(n235) );
  INV_X1 U1498 ( .A(n48684), .ZN(n236) );
  OAI211_X1 U1506 ( .C1(n30160), .C2(n30177), .A(n29139), .B(n237), .ZN(n4082)
         );
  NAND3_X1 U1511 ( .A1(n27642), .A2(n27640), .A3(n27641), .ZN(n8275) );
  NAND2_X1 U1512 ( .A1(n239), .A2(n38676), .ZN(n38240) );
  OAI21_X1 U1513 ( .B1(n38245), .B2(n38237), .A(n39167), .ZN(n239) );
  AND3_X2 U1516 ( .A1(n19548), .A2(n19547), .A3(n19546), .ZN(n20903) );
  BUF_X2 U1519 ( .A(n17287), .Z(n21270) );
  NAND2_X1 U1520 ( .A1(n420), .A2(n37924), .ZN(n39169) );
  OR2_X2 U1522 ( .A1(n38251), .A2(n38250), .ZN(n40874) );
  BUF_X2 U1523 ( .A(n18804), .Z(n2225) );
  NAND4_X1 U1525 ( .A1(n50730), .A2(n240), .A3(n7745), .A4(n7744), .ZN(n7742)
         );
  INV_X1 U1526 ( .A(n7748), .ZN(n240) );
  OAI21_X1 U1527 ( .B1(n36782), .B2(n8462), .A(n2571), .ZN(n241) );
  NAND4_X2 U1536 ( .A1(n35912), .A2(n35913), .A3(n35911), .A4(n35910), .ZN(
        n1491) );
  NAND4_X1 U1537 ( .A1(n244), .A2(n43431), .A3(n43422), .A4(n43423), .ZN(n5684) );
  NAND2_X1 U1538 ( .A1(n43430), .A2(n45945), .ZN(n244) );
  NAND3_X1 U1539 ( .A1(n48469), .A2(n48457), .A3(n46411), .ZN(n42509) );
  XNOR2_X2 U1540 ( .A(n43366), .B(n245), .ZN(n49137) );
  XNOR2_X1 U1541 ( .A(n43361), .B(n43362), .ZN(n245) );
  NAND3_X1 U1543 ( .A1(n29254), .A2(n29119), .A3(n29259), .ZN(n25632) );
  NAND2_X1 U1549 ( .A1(n3589), .A2(n19837), .ZN(n19527) );
  NAND3_X1 U1551 ( .A1(n6883), .A2(n6887), .A3(n246), .ZN(n6882) );
  NAND4_X2 U1553 ( .A1(n20912), .A2(n20913), .A3(n20914), .A4(n20911), .ZN(
        n28370) );
  NAND2_X1 U1555 ( .A1(n38944), .A2(n39201), .ZN(n248) );
  NAND2_X2 U1557 ( .A1(n35439), .A2(n35438), .ZN(n44027) );
  NAND4_X2 U1560 ( .A1(n23265), .A2(n23264), .A3(n23263), .A4(n23262), .ZN(
        n6656) );
  NAND3_X1 U1562 ( .A1(n38644), .A2(n4139), .A3(n38643), .ZN(n38645) );
  NAND2_X1 U1564 ( .A1(n12253), .A2(n11345), .ZN(n9423) );
  NAND2_X1 U1565 ( .A1(n4479), .A2(n250), .ZN(n24007) );
  NAND3_X1 U1567 ( .A1(n252), .A2(n37640), .A3(n251), .ZN(n35199) );
  NAND2_X1 U1568 ( .A1(n37649), .A2(n34632), .ZN(n251) );
  NAND2_X1 U1569 ( .A1(n36403), .A2(n5590), .ZN(n252) );
  NAND3_X2 U1570 ( .A1(n30897), .A2(n4489), .A3(n30896), .ZN(n34841) );
  AND2_X2 U1576 ( .A1(n4246), .A2(n36015), .ZN(n36558) );
  BUF_X1 U1577 ( .A(n18780), .Z(n2162) );
  AND3_X2 U1582 ( .A1(n8816), .A2(n8815), .A3(n8814), .ZN(n13590) );
  OR2_X2 U1586 ( .A1(n30500), .A2(n30499), .ZN(n35075) );
  NAND2_X1 U1591 ( .A1(n256), .A2(n255), .ZN(n27866) );
  NAND2_X1 U1592 ( .A1(n27864), .A2(n29495), .ZN(n255) );
  NAND2_X1 U1593 ( .A1(n27865), .A2(n257), .ZN(n256) );
  NAND2_X1 U1597 ( .A1(n29988), .A2(n2366), .ZN(n259) );
  XNOR2_X1 U1602 ( .A(n35825), .B(n260), .ZN(n34584) );
  XNOR2_X1 U1603 ( .A(n34454), .B(n34037), .ZN(n260) );
  NAND3_X1 U1605 ( .A1(n1427), .A2(n32404), .A3(n714), .ZN(n32072) );
  XNOR2_X1 U1607 ( .A(n261), .B(n35562), .ZN(n35564) );
  XNOR2_X1 U1608 ( .A(n35559), .B(n35560), .ZN(n261) );
  NAND3_X1 U1609 ( .A1(n14226), .A2(n14227), .A3(n16221), .ZN(n13224) );
  NAND2_X1 U1610 ( .A1(n32346), .A2(n32437), .ZN(n32349) );
  AND2_X2 U1613 ( .A1(n17740), .A2(n21473), .ZN(n20316) );
  NAND2_X1 U1617 ( .A1(n264), .A2(n263), .ZN(n36107) );
  NAND2_X1 U1618 ( .A1(n688), .A2(n38196), .ZN(n264) );
  AOI21_X2 U1621 ( .B1(n20382), .B2(n3411), .A(n20381), .ZN(n22085) );
  NAND4_X2 U1622 ( .A1(n32362), .A2(n32363), .A3(n32364), .A4(n32361), .ZN(
        n37261) );
  NAND3_X1 U1624 ( .A1(n26773), .A2(n6290), .A3(n26810), .ZN(n4097) );
  NAND3_X1 U1625 ( .A1(n39502), .A2(n40665), .A3(n685), .ZN(n36180) );
  NAND2_X1 U1635 ( .A1(n43462), .A2(n49722), .ZN(n45993) );
  NAND2_X1 U1636 ( .A1(n49717), .A2(n49725), .ZN(n43462) );
  NAND2_X2 U1638 ( .A1(n3442), .A2(n21059), .ZN(n26147) );
  XNOR2_X1 U1639 ( .A(n15019), .B(n51417), .ZN(n15026) );
  AND2_X2 U1642 ( .A1(n11359), .A2(n12113), .ZN(n12111) );
  NAND3_X1 U1646 ( .A1(n21171), .A2(n21188), .A3(n5271), .ZN(n5274) );
  NAND2_X1 U1647 ( .A1(n10932), .A2(n10219), .ZN(n10135) );
  NAND3_X2 U1651 ( .A1(n2941), .A2(n2942), .A3(n31102), .ZN(n35105) );
  NAND2_X1 U1655 ( .A1(n5272), .A2(n21181), .ZN(n267) );
  INV_X1 U1656 ( .A(n268), .ZN(n35886) );
  OAI21_X1 U1657 ( .B1(n36462), .B2(n36448), .A(n36598), .ZN(n268) );
  NAND2_X1 U1658 ( .A1(n50265), .A2(n47058), .ZN(n47333) );
  NAND3_X1 U1659 ( .A1(n16870), .A2(n2869), .A3(n16871), .ZN(n17005) );
  NAND3_X1 U1660 ( .A1(n28541), .A2(n28540), .A3(n269), .ZN(n28543) );
  NAND2_X1 U1670 ( .A1(n3604), .A2(n19713), .ZN(n18886) );
  INV_X1 U1674 ( .A(n22179), .ZN(n22178) );
  NAND2_X1 U1675 ( .A1(n21700), .A2(n21714), .ZN(n22179) );
  AND3_X2 U1678 ( .A1(n2558), .A2(n2561), .A3(n2562), .ZN(n22186) );
  INV_X1 U1679 ( .A(n46398), .ZN(n46394) );
  NAND2_X1 U1680 ( .A1(n46483), .A2(n46503), .ZN(n46398) );
  INV_X1 U1687 ( .A(n38367), .ZN(n270) );
  NAND2_X1 U1691 ( .A1(n2684), .A2(n2459), .ZN(n271) );
  NAND2_X2 U1692 ( .A1(n7392), .A2(n7574), .ZN(n31624) );
  XNOR2_X1 U1694 ( .A(n272), .B(n47584), .ZN(Plaintext[5]) );
  AND2_X1 U1695 ( .A1(n47583), .A2(n47568), .ZN(n273) );
  NAND4_X2 U1696 ( .A1(n21159), .A2(n21160), .A3(n21161), .A4(n22273), .ZN(
        n27232) );
  XNOR2_X1 U1699 ( .A(n275), .B(n50795), .ZN(Plaintext[177]) );
  NAND4_X1 U1700 ( .A1(n50794), .A2(n50791), .A3(n50793), .A4(n50792), .ZN(
        n275) );
  NAND4_X2 U1702 ( .A1(n9416), .A2(n9415), .A3(n9414), .A4(n9413), .ZN(n11315)
         );
  NAND3_X1 U1707 ( .A1(n21779), .A2(n24452), .A3(n21778), .ZN(n21785) );
  NAND2_X1 U1710 ( .A1(n36490), .A2(n35315), .ZN(n36472) );
  BUF_X1 U1715 ( .A(n9218), .Z(n12055) );
  NAND2_X1 U1718 ( .A1(n276), .A2(n15046), .ZN(n10407) );
  NAND2_X1 U1719 ( .A1(n13480), .A2(n277), .ZN(n276) );
  OR2_X2 U1720 ( .A1(n18014), .A2(n5336), .ZN(n19398) );
  OAI211_X1 U1723 ( .C1(n8764), .C2(n50549), .A(n50568), .B(n50567), .ZN(
        n50571) );
  NAND2_X1 U1729 ( .A1(n29886), .A2(n30734), .ZN(n30743) );
  NAND3_X2 U1731 ( .A1(n7497), .A2(n3773), .A3(n7496), .ZN(n3772) );
  AND4_X2 U1735 ( .A1(n44697), .A2(n44699), .A3(n44700), .A4(n44698), .ZN(
        n47962) );
  NAND3_X1 U1736 ( .A1(n17613), .A2(n2478), .A3(n50991), .ZN(n22152) );
  AND3_X2 U1742 ( .A1(n27406), .A2(n1120), .A3(n1123), .ZN(n32787) );
  NAND3_X1 U1744 ( .A1(n30847), .A2(n31820), .A3(n6107), .ZN(n30851) );
  NAND2_X1 U1746 ( .A1(n3393), .A2(n30080), .ZN(n30090) );
  XNOR2_X2 U1747 ( .A(n278), .B(n41850), .ZN(n45393) );
  NAND2_X1 U1748 ( .A1(n43671), .A2(n4308), .ZN(n278) );
  NAND2_X1 U1749 ( .A1(n30824), .A2(n31301), .ZN(n30825) );
  NOR2_X1 U1751 ( .A1(n16797), .A2(n18291), .ZN(n15089) );
  NAND2_X1 U1752 ( .A1(n633), .A2(n17522), .ZN(n18291) );
  NAND2_X1 U1753 ( .A1(n12068), .A2(n9207), .ZN(n12073) );
  NAND2_X2 U1757 ( .A1(n4356), .A2(n4355), .ZN(n40330) );
  INV_X2 U1762 ( .A(n900), .ZN(n31904) );
  NOR2_X2 U1763 ( .A1(n4345), .A2(n13061), .ZN(n15254) );
  INV_X1 U1768 ( .A(n49646), .ZN(n49666) );
  NAND2_X1 U1769 ( .A1(n52212), .A2(n51733), .ZN(n49646) );
  NAND2_X1 U1770 ( .A1(n279), .A2(n48646), .ZN(n48629) );
  OAI22_X1 U1771 ( .A1(n48625), .A2(n48616), .B1(n48617), .B2(n48618), .ZN(
        n279) );
  XNOR2_X1 U1773 ( .A(n18421), .B(n18420), .ZN(n280) );
  AND2_X2 U1774 ( .A1(n49209), .A2(n45970), .ZN(n49203) );
  NAND2_X1 U1776 ( .A1(n26891), .A2(n27618), .ZN(n24571) );
  BUF_X2 U1778 ( .A(n45370), .Z(n48227) );
  NAND3_X2 U1779 ( .A1(n5778), .A2(n32086), .A3(n32084), .ZN(n5777) );
  OR2_X2 U1784 ( .A1(n13229), .A2(n13237), .ZN(n13221) );
  XNOR2_X2 U1785 ( .A(n282), .B(n33428), .ZN(n37774) );
  AND4_X2 U1789 ( .A1(n2001), .A2(n43092), .A3(n2002), .A4(n43093), .ZN(n49569) );
  NAND3_X2 U1791 ( .A1(n41713), .A2(n283), .A3(n51634), .ZN(n46113) );
  NAND2_X1 U1792 ( .A1(n41701), .A2(n41700), .ZN(n283) );
  AOI22_X1 U1795 ( .A1(n1712), .A2(n22697), .B1(n21778), .B2(n22287), .ZN(
        n1710) );
  OAI21_X1 U1797 ( .B1(n11100), .B2(n8944), .A(n286), .ZN(n8956) );
  NAND2_X1 U1798 ( .A1(n8944), .A2(n8942), .ZN(n286) );
  NAND2_X1 U1799 ( .A1(n8389), .A2(n32177), .ZN(n287) );
  NOR2_X2 U1802 ( .A1(n21200), .A2(n6078), .ZN(n21208) );
  NAND2_X1 U1804 ( .A1(n8155), .A2(n5966), .ZN(n3320) );
  NAND3_X1 U1805 ( .A1(n46651), .A2(n46846), .A3(n46676), .ZN(n46650) );
  NAND2_X1 U1807 ( .A1(n288), .A2(n22509), .ZN(n21070) );
  NAND2_X1 U1809 ( .A1(n11881), .A2(n8901), .ZN(n8907) );
  OAI21_X1 U1810 ( .B1(n11884), .B2(n12680), .A(n12462), .ZN(n11881) );
  NAND2_X1 U1812 ( .A1(n31803), .A2(n52047), .ZN(n31789) );
  BUF_X2 U1813 ( .A(n19214), .Z(n2181) );
  INV_X2 U1814 ( .A(n22748), .ZN(n23054) );
  OR2_X2 U1815 ( .A1(n33879), .A2(n33878), .ZN(n43669) );
  NAND2_X1 U1819 ( .A1(n12178), .A2(n12170), .ZN(n3615) );
  NAND2_X1 U1820 ( .A1(n52132), .A2(n11322), .ZN(n12170) );
  NAND3_X1 U1821 ( .A1(n36002), .A2(n37649), .A3(n289), .ZN(n6647) );
  XNOR2_X1 U1824 ( .A(n17819), .B(n17818), .ZN(n291) );
  NAND2_X1 U1829 ( .A1(n293), .A2(n30789), .ZN(n3503) );
  OAI22_X1 U1830 ( .A1(n27564), .A2(n30794), .B1(n29907), .B2(n29899), .ZN(
        n293) );
  NAND4_X2 U1832 ( .A1(n37995), .A2(n37993), .A3(n37992), .A4(n37994), .ZN(
        n40909) );
  NAND3_X1 U1835 ( .A1(n294), .A2(n12072), .A3(n9208), .ZN(n12078) );
  NAND2_X1 U1836 ( .A1(n1167), .A2(n12067), .ZN(n294) );
  NAND2_X1 U1837 ( .A1(n16490), .A2(n19535), .ZN(n19055) );
  NAND2_X1 U1841 ( .A1(n17310), .A2(n17413), .ZN(n21239) );
  AND2_X2 U1842 ( .A1(n7340), .A2(n51760), .ZN(n12557) );
  NAND2_X1 U1843 ( .A1(n295), .A2(n39728), .ZN(n39736) );
  OAI211_X1 U1844 ( .C1(n41040), .C2(n41286), .A(n41031), .B(n40430), .ZN(n295) );
  NAND3_X1 U1846 ( .A1(n3938), .A2(n24296), .A3(n24295), .ZN(n3937) );
  NAND3_X1 U1847 ( .A1(n41633), .A2(n41635), .A3(n41634), .ZN(n1207) );
  NAND2_X1 U1848 ( .A1(n48722), .A2(n995), .ZN(n48726) );
  NAND2_X1 U1849 ( .A1(n1150), .A2(n32138), .ZN(n32139) );
  XNOR2_X1 U1850 ( .A(n296), .B(n45363), .ZN(n45369) );
  XNOR2_X1 U1851 ( .A(n45361), .B(n45362), .ZN(n296) );
  NAND2_X1 U1852 ( .A1(n10111), .A2(n10112), .ZN(n10113) );
  NAND3_X1 U1853 ( .A1(n14019), .A2(n14022), .A3(n14020), .ZN(n2006) );
  NOR2_X2 U1857 ( .A1(n32251), .A2(n31778), .ZN(n31238) );
  OR2_X2 U1859 ( .A1(n401), .A2(n30393), .ZN(n30696) );
  OAI22_X1 U1862 ( .A1(n10935), .A2(n10934), .B1(n10933), .B2(n10932), .ZN(
        n297) );
  NAND2_X1 U1864 ( .A1(n21312), .A2(n21313), .ZN(n21317) );
  OR2_X2 U1865 ( .A1(n21252), .A2(n3885), .ZN(n19475) );
  NAND3_X1 U1869 ( .A1(n37942), .A2(n39270), .A3(n39016), .ZN(n36775) );
  NAND2_X1 U1873 ( .A1(n300), .A2(n299), .ZN(n5456) );
  NAND2_X1 U1874 ( .A1(n17065), .A2(n51403), .ZN(n299) );
  NAND2_X1 U1875 ( .A1(n16567), .A2(n19071), .ZN(n300) );
  NAND2_X1 U1878 ( .A1(n21528), .A2(n51625), .ZN(n301) );
  NAND3_X1 U1881 ( .A1(n303), .A2(n1993), .A3(n20286), .ZN(n20287) );
  NAND2_X1 U1882 ( .A1(n1992), .A2(n24242), .ZN(n303) );
  NAND2_X1 U1891 ( .A1(n52132), .A2(n10413), .ZN(n12175) );
  BUF_X1 U1898 ( .A(n11558), .Z(n15385) );
  OAI22_X1 U1901 ( .A1(n18846), .A2(n1704), .B1(n18847), .B2(n20660), .ZN(
        n15833) );
  NAND2_X1 U1902 ( .A1(n17584), .A2(n20515), .ZN(n18081) );
  AND2_X1 U1905 ( .A1(n6627), .A2(n15837), .ZN(n6625) );
  INV_X1 U1906 ( .A(n22188), .ZN(n7119) );
  NAND2_X1 U1907 ( .A1(n452), .A2(n23409), .ZN(n23425) );
  INV_X1 U1908 ( .A(n26565), .ZN(n1026) );
  INV_X1 U1910 ( .A(n23810), .ZN(n23814) );
  NAND4_X1 U1912 ( .A1(n21943), .A2(n21941), .A3(n21940), .A4(n21942), .ZN(
        n24655) );
  XNOR2_X1 U1915 ( .A(n26015), .B(n26014), .ZN(n1023) );
  INV_X1 U1917 ( .A(n30265), .ZN(n29235) );
  XNOR2_X1 U1918 ( .A(n24916), .B(n24923), .ZN(n1500) );
  OR2_X1 U1919 ( .A1(n30710), .A2(n30706), .ZN(n1153) );
  NAND2_X1 U1922 ( .A1(n51111), .A2(n27695), .ZN(n29549) );
  NAND2_X1 U1923 ( .A1(n51514), .A2(n29159), .ZN(n7532) );
  AND2_X1 U1925 ( .A1(n31816), .A2(n30576), .ZN(n2028) );
  OR2_X1 U1926 ( .A1(n29736), .A2(n29749), .ZN(n30449) );
  NOR2_X1 U1927 ( .A1(n30647), .A2(n51086), .ZN(n30652) );
  INV_X1 U1928 ( .A(n31546), .ZN(n31169) );
  AND2_X1 U1929 ( .A1(n32883), .A2(n719), .ZN(n5498) );
  NAND2_X1 U1932 ( .A1(n37499), .A2(n37757), .ZN(n34914) );
  NAND2_X1 U1934 ( .A1(n38164), .A2(n38593), .ZN(n37448) );
  INV_X1 U1935 ( .A(n5711), .ZN(n37980) );
  OR2_X1 U1937 ( .A1(n37765), .A2(n36248), .ZN(n37753) );
  AND2_X1 U1940 ( .A1(n40876), .A2(n678), .ZN(n38356) );
  AND2_X1 U1941 ( .A1(n41645), .A2(n41103), .ZN(n41638) );
  INV_X1 U1945 ( .A(n41691), .ZN(n41695) );
  OR2_X1 U1946 ( .A1(n51853), .A2(n40963), .ZN(n41372) );
  AOI21_X1 U1947 ( .B1(n41646), .B2(n41094), .A(n1706), .ZN(n1705) );
  OR2_X1 U1948 ( .A1(n540), .A2(n664), .ZN(n1586) );
  INV_X1 U1950 ( .A(n46899), .ZN(n46903) );
  INV_X1 U1951 ( .A(n44665), .ZN(n660) );
  NOR2_X1 U1952 ( .A1(n49237), .A2(n656), .ZN(n1251) );
  OAI21_X1 U1953 ( .B1(n49178), .B2(n49177), .A(n49176), .ZN(n49179) );
  INV_X1 U1954 ( .A(n5668), .ZN(n45937) );
  OR2_X1 U1958 ( .A1(n12106), .A2(n9639), .ZN(n304) );
  OR2_X1 U1960 ( .A1(n12711), .A2(n1781), .ZN(n306) );
  AND3_X1 U1961 ( .A1(n9999), .A2(n9998), .A3(n807), .ZN(n307) );
  AND3_X1 U1962 ( .A1(n10001), .A2(n10577), .A3(n1280), .ZN(n308) );
  XOR2_X1 U1963 ( .A(n33768), .B(n17685), .Z(n309) );
  XOR2_X1 U1965 ( .A(n45040), .B(n45039), .Z(n310) );
  AND3_X1 U1966 ( .A1(n13057), .A2(n14791), .A3(n11055), .ZN(n311) );
  AND3_X1 U1967 ( .A1(n14038), .A2(n14026), .A3(n14027), .ZN(n312) );
  OR2_X1 U1968 ( .A1(n13334), .A2(n14197), .ZN(n313) );
  INV_X1 U1969 ( .A(n22403), .ZN(n23230) );
  AND2_X1 U1970 ( .A1(n39716), .A2(n6870), .ZN(n314) );
  BUF_X1 U1971 ( .A(n48413), .Z(n506) );
  AND2_X1 U1972 ( .A1(n48515), .A2(n48514), .ZN(n315) );
  INV_X1 U1973 ( .A(n16546), .ZN(n18356) );
  AND3_X1 U1975 ( .A1(n3342), .A2(n20322), .A3(n20840), .ZN(n316) );
  XNOR2_X2 U1976 ( .A(n18466), .B(n17965), .ZN(n18704) );
  OR2_X1 U1977 ( .A1(n20266), .A2(n1704), .ZN(n317) );
  AND2_X1 U1978 ( .A1(n21401), .A2(n21399), .ZN(n318) );
  OR2_X1 U1981 ( .A1(n21222), .A2(n1456), .ZN(n319) );
  BUF_X2 U1982 ( .A(n24029), .Z(n354) );
  NAND4_X2 U1985 ( .A1(n15839), .A2(n6626), .A3(n6625), .A4(n15838), .ZN(
        n23821) );
  NAND2_X1 U1986 ( .A1(n22832), .A2(n22826), .ZN(n320) );
  OR2_X1 U1987 ( .A1(n22562), .A2(n22982), .ZN(n321) );
  XOR2_X1 U1988 ( .A(n3110), .B(n2541), .Z(n322) );
  NAND4_X2 U1989 ( .A1(n1954), .A2(n1955), .A3(n1956), .A4(n1958), .ZN(n26390)
         );
  BUF_X2 U1992 ( .A(n27281), .Z(n28974) );
  AND2_X1 U1993 ( .A1(n24248), .A2(n20285), .ZN(n323) );
  AND2_X1 U1995 ( .A1(n4971), .A2(n23110), .ZN(n324) );
  OR2_X1 U1997 ( .A1(n29989), .A2(n31425), .ZN(n325) );
  OR2_X1 U1999 ( .A1(n27760), .A2(n27745), .ZN(n326) );
  INV_X2 U2000 ( .A(n31067), .ZN(n3099) );
  AND3_X1 U2003 ( .A1(n31487), .A2(n30102), .A3(n1738), .ZN(n327) );
  XOR2_X1 U2004 ( .A(n34889), .B(n34157), .Z(n328) );
  XNOR2_X1 U2005 ( .A(n33112), .B(n33111), .ZN(n329) );
  BUF_X2 U2008 ( .A(n33981), .Z(n2168) );
  AND2_X1 U2009 ( .A1(n3490), .A2(n3489), .ZN(n331) );
  AND4_X2 U2012 ( .A1(n35740), .A2(n35739), .A3(n35738), .A4(n6646), .ZN(
        n39906) );
  AND2_X1 U2017 ( .A1(n41702), .A2(n41694), .ZN(n333) );
  AND3_X1 U2019 ( .A1(n38618), .A2(n33178), .A3(n1100), .ZN(n334) );
  XOR2_X1 U2021 ( .A(n44932), .B(n43759), .Z(n335) );
  BUF_X1 U2022 ( .A(n42181), .Z(n44828) );
  AND2_X1 U2028 ( .A1(n48309), .A2(n912), .ZN(n336) );
  OR2_X1 U2029 ( .A1(n49265), .A2(n49263), .ZN(n337) );
  AND2_X1 U2030 ( .A1(n49521), .A2(n49487), .ZN(n338) );
  AND2_X1 U2031 ( .A1(n1176), .A2(n1175), .ZN(n339) );
  NAND3_X2 U2032 ( .A1(n45249), .A2(n45248), .A3(n45247), .ZN(n45739) );
  AND2_X1 U2034 ( .A1(n47435), .A2(n47442), .ZN(n340) );
  AND3_X1 U2036 ( .A1(n50136), .A2(n50097), .A3(n50088), .ZN(n341) );
  OR2_X1 U2037 ( .A1(n50469), .A2(n50468), .ZN(n342) );
  AND3_X1 U2038 ( .A1(n45845), .A2(n46692), .A3(n52169), .ZN(n343) );
  OR2_X1 U2039 ( .A1(n50871), .A2(n1441), .ZN(n344) );
  AND3_X1 U2040 ( .A1(n47791), .A2(n47789), .A3(n52118), .ZN(n345) );
  NAND4_X1 U2045 ( .A1(n49179), .A2(n8020), .A3(n49180), .A4(n49173), .ZN(
        n49375) );
  XNOR2_X1 U2048 ( .A(n9253), .B(Key[138]), .ZN(n12612) );
  NAND4_X1 U2050 ( .A1(n8957), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(n15102)
         );
  BUF_X1 U2053 ( .A(n17170), .Z(n355) );
  BUF_X2 U2054 ( .A(n17170), .Z(n356) );
  XNOR2_X1 U2055 ( .A(n16064), .B(n18134), .ZN(n17170) );
  NAND2_X2 U2056 ( .A1(n47376), .A2(n47377), .ZN(n50235) );
  OR2_X2 U2057 ( .A1(n46358), .A2(n46267), .ZN(n46277) );
  XNOR2_X1 U2060 ( .A(Key[21]), .B(Ciphertext[32]), .ZN(n11136) );
  XNOR2_X1 U2062 ( .A(n17979), .B(n17978), .ZN(n21391) );
  XNOR2_X1 U2065 ( .A(n44937), .B(n45314), .ZN(n46042) );
  NAND4_X1 U2070 ( .A1(n7293), .A2(n26984), .A3(n2295), .A4(n7292), .ZN(n31940) );
  NAND4_X1 U2077 ( .A1(n13835), .A2(n13836), .A3(n13834), .A4(n13833), .ZN(
        n18431) );
  XNOR2_X1 U2080 ( .A(n28423), .B(n8368), .ZN(n28301) );
  OAI21_X1 U2083 ( .B1(n41140), .B2(n41139), .A(n5309), .ZN(n47868) );
  XNOR2_X1 U2086 ( .A(n6599), .B(n16969), .ZN(n18261) );
  NAND4_X1 U2088 ( .A1(n26715), .A2(n26714), .A3(n26716), .A4(n26713), .ZN(
        n34544) );
  XNOR2_X1 U2091 ( .A(n25491), .B(n25490), .ZN(n27783) );
  NAND2_X1 U2096 ( .A1(n8180), .A2(n30730), .ZN(n31545) );
  XNOR2_X1 U2100 ( .A(n25875), .B(n25874), .ZN(n28638) );
  NOR2_X1 U2101 ( .A1(n16892), .A2(n18847), .ZN(n1990) );
  NOR2_X2 U2103 ( .A1(n7684), .A2(n51025), .ZN(n50352) );
  NAND4_X1 U2105 ( .A1(n27947), .A2(n27949), .A3(n27948), .A4(n27950), .ZN(
        n31748) );
  BUF_X1 U2107 ( .A(n46996), .Z(n388) );
  BUF_X1 U2108 ( .A(n46996), .Z(n389) );
  XNOR2_X1 U2110 ( .A(n25567), .B(n25568), .ZN(n28659) );
  NAND4_X1 U2113 ( .A1(n30190), .A2(n30302), .A3(n30319), .A4(n30189), .ZN(
        n31567) );
  XNOR2_X1 U2118 ( .A(n28430), .B(n25589), .ZN(n7877) );
  NAND2_X2 U2120 ( .A1(n1103), .A2(n44274), .ZN(n48051) );
  OR2_X1 U2121 ( .A1(n6775), .A2(n6779), .ZN(n397) );
  XNOR2_X1 U2123 ( .A(n26219), .B(n26218), .ZN(n29533) );
  BUF_X1 U2126 ( .A(n29930), .Z(n401) );
  XNOR2_X1 U2128 ( .A(n24015), .B(n24014), .ZN(n29930) );
  NOR2_X2 U2131 ( .A1(n30568), .A2(n30567), .ZN(n32859) );
  BUF_X1 U2134 ( .A(n45793), .Z(n405) );
  XNOR2_X1 U2136 ( .A(n41366), .B(n41365), .ZN(n45793) );
  XNOR2_X1 U2137 ( .A(n42856), .B(n42857), .ZN(n49695) );
  BUF_X2 U2146 ( .A(n23208), .Z(n413) );
  NAND4_X1 U2147 ( .A1(n6316), .A2(n6314), .A3(n6315), .A4(n18325), .ZN(n23208) );
  NOR2_X1 U2149 ( .A1(n46684), .A2(n46683), .ZN(n47528) );
  AND2_X2 U2150 ( .A1(n27858), .A2(n51110), .ZN(n2294) );
  NAND2_X2 U2153 ( .A1(n8362), .A2(n8363), .ZN(n24026) );
  NAND3_X2 U2154 ( .A1(n3972), .A2(n5144), .A3(n2374), .ZN(n23924) );
  XNOR2_X2 U2155 ( .A(n36764), .B(n37325), .ZN(n35283) );
  BUF_X1 U2157 ( .A(n22403), .Z(n417) );
  BUF_X1 U2158 ( .A(n22403), .Z(n418) );
  OAI211_X1 U2159 ( .C1(n20027), .C2(n18379), .A(n7582), .B(n7579), .ZN(n22403) );
  BUF_X2 U2161 ( .A(n39181), .Z(n420) );
  XNOR2_X1 U2162 ( .A(n37076), .B(n37075), .ZN(n39181) );
  XNOR2_X1 U2168 ( .A(n46136), .B(n46135), .ZN(n50382) );
  NAND2_X1 U2169 ( .A1(n31904), .A2(n32830), .ZN(n8536) );
  AND4_X2 U2170 ( .A1(n5841), .A2(n30373), .A3(n5840), .A4(n30372), .ZN(n32830) );
  BUF_X2 U2171 ( .A(n45192), .Z(n50906) );
  NAND4_X1 U2175 ( .A1(n37459), .A2(n37458), .A3(n37457), .A4(n37456), .ZN(
        n40792) );
  XNOR2_X1 U2177 ( .A(n28406), .B(n28405), .ZN(n30442) );
  XNOR2_X1 U2180 ( .A(n44061), .B(n5379), .ZN(n45122) );
  NAND2_X2 U2182 ( .A1(n30972), .A2(n30973), .ZN(n37081) );
  NAND4_X2 U2184 ( .A1(n38932), .A2(n38935), .A3(n38934), .A4(n38933), .ZN(
        n43170) );
  NAND4_X2 U2186 ( .A1(n1607), .A2(n1606), .A3(n24163), .A4(n24162), .ZN(
        n26175) );
  BUF_X2 U2187 ( .A(n21698), .Z(n21712) );
  NAND4_X2 U2189 ( .A1(n20293), .A2(n18277), .A3(n18276), .A4(n18278), .ZN(
        n26119) );
  XNOR2_X1 U2191 ( .A(n26037), .B(n26038), .ZN(n29442) );
  NAND2_X1 U2194 ( .A1(n4806), .A2(n40062), .ZN(n40781) );
  XNOR2_X1 U2197 ( .A(n27220), .B(n27219), .ZN(n29718) );
  XNOR2_X1 U2201 ( .A(n8487), .B(Key[59]), .ZN(n12145) );
  NAND4_X2 U2202 ( .A1(n14557), .A2(n14555), .A3(n14556), .A4(n14554), .ZN(
        n16464) );
  XNOR2_X1 U2205 ( .A(n43894), .B(n43895), .ZN(n50338) );
  BUF_X2 U2206 ( .A(n23304), .Z(n441) );
  NAND4_X1 U2207 ( .A1(n5535), .A2(n5537), .A3(n5534), .A4(n21518), .ZN(n23304) );
  OAI21_X2 U2208 ( .B1(n43673), .B2(n43672), .A(n43671), .ZN(n45258) );
  XNOR2_X1 U2210 ( .A(n8931), .B(Key[53]), .ZN(n12542) );
  XNOR2_X1 U2215 ( .A(n25124), .B(n24022), .ZN(n7558) );
  NAND4_X1 U2220 ( .A1(n48226), .A2(n48225), .A3(n48223), .A4(n48224), .ZN(
        n48391) );
  BUF_X1 U2221 ( .A(n27663), .Z(n447) );
  XNOR2_X1 U2223 ( .A(n5387), .B(n5386), .ZN(n27663) );
  BUF_X1 U2229 ( .A(n11636), .Z(n453) );
  BUF_X2 U2230 ( .A(n11636), .Z(n454) );
  XNOR2_X1 U2231 ( .A(n9095), .B(Key[62]), .ZN(n11636) );
  XNOR2_X1 U2234 ( .A(n34502), .B(n34501), .ZN(n34529) );
  NAND4_X1 U2238 ( .A1(n20690), .A2(n6919), .A3(n20691), .A4(n20689), .ZN(
        n24333) );
  AND3_X2 U2240 ( .A1(n5404), .A2(n5401), .A3(n5398), .ZN(n46059) );
  XNOR2_X1 U2242 ( .A(n34108), .B(n34107), .ZN(n36575) );
  XNOR2_X1 U2245 ( .A(n35483), .B(n35683), .ZN(n36881) );
  XNOR2_X1 U2248 ( .A(n17902), .B(n16980), .ZN(n18535) );
  BUF_X2 U2249 ( .A(n22188), .Z(n463) );
  AND2_X2 U2252 ( .A1(n50031), .A2(n50032), .ZN(n50145) );
  BUF_X1 U2258 ( .A(n39028), .Z(n467) );
  NAND4_X1 U2262 ( .A1(n10975), .A2(n10974), .A3(n10973), .A4(n10972), .ZN(
        n14029) );
  BUF_X2 U2264 ( .A(n26228), .Z(n471) );
  XNOR2_X1 U2265 ( .A(n7350), .B(n7254), .ZN(n26228) );
  XNOR2_X1 U2272 ( .A(n33842), .B(n33841), .ZN(n38972) );
  XNOR2_X1 U2275 ( .A(Key[134]), .B(Ciphertext[7]), .ZN(n11409) );
  XNOR2_X2 U2279 ( .A(n33488), .B(n33487), .ZN(n38495) );
  NOR2_X2 U2280 ( .A1(n13740), .A2(n13739), .ZN(n17158) );
  AND3_X2 U2281 ( .A1(n6855), .A2(n28034), .A3(n6854), .ZN(n29618) );
  OAI211_X1 U2286 ( .C1(n36281), .C2(n36280), .A(n36279), .B(n36278), .ZN(
        n42054) );
  OR2_X1 U2290 ( .A1(n12324), .A2(n9667), .ZN(n12328) );
  NAND3_X2 U2292 ( .A1(n46564), .A2(n46563), .A3(n46562), .ZN(n47617) );
  BUF_X2 U2294 ( .A(n12890), .Z(n483) );
  NAND3_X1 U2295 ( .A1(n9967), .A2(n9966), .A3(n6041), .ZN(n12890) );
  NAND4_X1 U2299 ( .A1(n2005), .A2(n14040), .A3(n312), .A4(n14039), .ZN(n16470) );
  AND3_X2 U2302 ( .A1(n38989), .A2(n7207), .A3(n38990), .ZN(n41692) );
  BUF_X2 U2303 ( .A(n30426), .Z(n486) );
  XNOR2_X1 U2305 ( .A(n5984), .B(n27464), .ZN(n30426) );
  BUF_X2 U2306 ( .A(n28264), .Z(n488) );
  XNOR2_X1 U2307 ( .A(n23290), .B(n27232), .ZN(n28264) );
  XNOR2_X1 U2310 ( .A(n1110), .B(n17372), .ZN(n19336) );
  INV_X1 U2315 ( .A(n5713), .ZN(n25860) );
  XNOR2_X1 U2316 ( .A(n24655), .B(n25501), .ZN(n5713) );
  AND4_X2 U2317 ( .A1(n7398), .A2(n36334), .A3(n36332), .A4(n7397), .ZN(n39768) );
  OR2_X2 U2318 ( .A1(n40367), .A2(n5127), .ZN(n42962) );
  NOR2_X1 U2321 ( .A1(n7047), .A2(n46830), .ZN(n46824) );
  NAND3_X2 U2322 ( .A1(n8106), .A2(n12762), .A3(n8105), .ZN(n16923) );
  NAND4_X1 U2324 ( .A1(n33284), .A2(n334), .A3(n33282), .A4(n33283), .ZN(
        n46121) );
  XNOR2_X1 U2330 ( .A(n26448), .B(n28238), .ZN(n26607) );
  BUF_X1 U2338 ( .A(n47026), .Z(n505) );
  NAND2_X1 U2345 ( .A1(n4070), .A2(n4367), .ZN(n507) );
  BUF_X2 U2347 ( .A(n22061), .Z(n23182) );
  XNOR2_X1 U2355 ( .A(n18146), .B(n18145), .ZN(n21303) );
  XNOR2_X2 U2356 ( .A(n5517), .B(n23939), .ZN(n27632) );
  XNOR2_X2 U2357 ( .A(n24226), .B(n24225), .ZN(n27558) );
  XNOR2_X1 U2358 ( .A(Key[175]), .B(Ciphertext[54]), .ZN(n11899) );
  NAND4_X2 U2362 ( .A1(n20899), .A2(n20900), .A3(n20898), .A4(n20897), .ZN(
        n25240) );
  AND4_X2 U2366 ( .A1(n5908), .A2(n11800), .A3(n5906), .A4(n5903), .ZN(n19186)
         );
  BUF_X2 U2367 ( .A(n30345), .Z(n514) );
  XNOR2_X1 U2368 ( .A(n28321), .B(n28320), .ZN(n30345) );
  BUF_X2 U2369 ( .A(n11433), .Z(n14455) );
  BUF_X2 U2370 ( .A(n43757), .Z(n516) );
  BUF_X1 U2371 ( .A(n37135), .Z(n517) );
  XNOR2_X1 U2372 ( .A(n34514), .B(n34163), .ZN(n37135) );
  BUF_X1 U2376 ( .A(n49369), .Z(n522) );
  BUF_X2 U2377 ( .A(n49369), .Z(n523) );
  NOR2_X1 U2378 ( .A1(n49281), .A2(n49280), .ZN(n49369) );
  AND4_X2 U2387 ( .A1(n29130), .A2(n29129), .A3(n29128), .A4(n29127), .ZN(
        n32066) );
  XNOR2_X1 U2399 ( .A(n1254), .B(n42254), .ZN(n46245) );
  BUF_X2 U2403 ( .A(n17134), .Z(n543) );
  NAND2_X1 U2404 ( .A1(n50286), .A2(n8763), .ZN(n544) );
  OR2_X2 U2406 ( .A1(n4206), .A2(n7344), .ZN(n46137) );
  BUF_X1 U2407 ( .A(n10419), .Z(n548) );
  XNOR2_X1 U2409 ( .A(n8680), .B(Key[12]), .ZN(n10419) );
  XNOR2_X1 U2411 ( .A(n36753), .B(n36754), .ZN(n39272) );
  BUF_X1 U2417 ( .A(n16373), .Z(n556) );
  XNOR2_X1 U2419 ( .A(n17646), .B(n5996), .ZN(n16373) );
  XNOR2_X2 U2420 ( .A(n2713), .B(n15618), .ZN(n19636) );
  XNOR2_X2 U2424 ( .A(n8833), .B(Key[98]), .ZN(n10143) );
  XNOR2_X2 U2433 ( .A(n23805), .B(n23804), .ZN(n27602) );
  XNOR2_X2 U2434 ( .A(n23579), .B(n27295), .ZN(n26239) );
  NAND2_X2 U2442 ( .A1(n1196), .A2(n7586), .ZN(n41276) );
  AND2_X1 U2443 ( .A1(n1716), .A2(n1717), .ZN(n567) );
  XNOR2_X1 U2447 ( .A(n41968), .B(n43354), .ZN(n44972) );
  NAND4_X2 U2451 ( .A1(n39848), .A2(n39845), .A3(n39846), .A4(n39847), .ZN(
        n44164) );
  NAND4_X1 U2452 ( .A1(n2709), .A2(n2710), .A3(n49971), .A4(n49970), .ZN(
        n50115) );
  XNOR2_X2 U2456 ( .A(n8966), .B(Key[105]), .ZN(n12700) );
  BUF_X2 U2458 ( .A(n16938), .Z(n576) );
  XNOR2_X1 U2459 ( .A(n17973), .B(n16559), .ZN(n16938) );
  XNOR2_X1 U2461 ( .A(n25444), .B(n27501), .ZN(n28127) );
  XNOR2_X1 U2464 ( .A(n8819), .B(Key[103]), .ZN(n11028) );
  XNOR2_X1 U2466 ( .A(n3467), .B(n17896), .ZN(n21392) );
  OAI21_X1 U2469 ( .B1(n10133), .B2(n10970), .A(n10132), .ZN(n13131) );
  XNOR2_X1 U2473 ( .A(n42901), .B(n42900), .ZN(n45922) );
  XNOR2_X1 U2478 ( .A(n3508), .B(n15962), .ZN(n17526) );
  XNOR2_X1 U2480 ( .A(n8898), .B(Key[72]), .ZN(n12453) );
  XNOR2_X2 U2481 ( .A(n3392), .B(Key[112]), .ZN(n10148) );
  XNOR2_X1 U2482 ( .A(n18615), .B(n18194), .ZN(n18820) );
  BUF_X2 U2483 ( .A(n28410), .Z(n593) );
  XNOR2_X1 U2486 ( .A(n6582), .B(n33928), .ZN(n5711) );
  XNOR2_X2 U2489 ( .A(n16518), .B(n16519), .ZN(n20147) );
  NOR2_X1 U2494 ( .A1(n43416), .A2(n647), .ZN(n4072) );
  NOR2_X1 U2495 ( .A1(n49906), .A2(n47423), .ZN(n1820) );
  OR2_X1 U2499 ( .A1(n48140), .A2(n46542), .ZN(n48116) );
  INV_X2 U2500 ( .A(n47945), .ZN(n47990) );
  INV_X1 U2501 ( .A(n48975), .ZN(n46954) );
  INV_X1 U2502 ( .A(n50128), .ZN(n50097) );
  NOR2_X1 U2503 ( .A1(n49580), .A2(n49606), .ZN(n49592) );
  INV_X2 U2504 ( .A(n2859), .ZN(n49442) );
  OR2_X1 U2507 ( .A1(n544), .A2(n50452), .ZN(n50473) );
  INV_X1 U2508 ( .A(n51298), .ZN(n50934) );
  OR2_X1 U2511 ( .A1(n50679), .A2(n50708), .ZN(n50700) );
  INV_X1 U2516 ( .A(n48734), .ZN(n995) );
  NAND2_X1 U2517 ( .A1(n47554), .A2(n47547), .ZN(n47527) );
  NAND2_X1 U2521 ( .A1(n48417), .A2(n46511), .ZN(n46337) );
  NOR2_X1 U2522 ( .A1(n46449), .A2(n7275), .ZN(n5429) );
  INV_X1 U2523 ( .A(n49659), .ZN(n1488) );
  CLKBUF_X1 U2524 ( .A(n45597), .Z(n48482) );
  INV_X1 U2526 ( .A(n46917), .ZN(n603) );
  INV_X1 U2529 ( .A(n7275), .ZN(n883) );
  NAND2_X1 U2530 ( .A1(n7216), .A2(n51326), .ZN(n49982) );
  INV_X1 U2531 ( .A(n50338), .ZN(n47271) );
  OR2_X1 U2537 ( .A1(n665), .A2(n48481), .ZN(n48485) );
  INV_X1 U2538 ( .A(n46635), .ZN(n47909) );
  INV_X1 U2542 ( .A(n48491), .ZN(n604) );
  INV_X1 U2545 ( .A(n50382), .ZN(n50034) );
  XNOR2_X1 U2559 ( .A(n1628), .B(n672), .ZN(n1627) );
  XNOR2_X1 U2560 ( .A(n45116), .B(n44944), .ZN(n43757) );
  XNOR2_X1 U2561 ( .A(n43950), .B(n2185), .ZN(n44878) );
  BUF_X1 U2562 ( .A(n40998), .Z(n44962) );
  BUF_X1 U2564 ( .A(n42380), .Z(n43915) );
  NAND4_X1 U2566 ( .A1(n39608), .A2(n39607), .A3(n39606), .A4(n39605), .ZN(
        n42590) );
  BUF_X2 U2567 ( .A(n44031), .Z(n608) );
  AND4_X1 U2568 ( .A1(n815), .A2(n40772), .A3(n40588), .A4(n40589), .ZN(n40603) );
  AND2_X1 U2571 ( .A1(n51348), .A2(n41057), .ZN(n2016) );
  INV_X1 U2572 ( .A(n39767), .ZN(n40652) );
  INV_X1 U2573 ( .A(n40903), .ZN(n40274) );
  NOR2_X1 U2575 ( .A1(n677), .A2(n40377), .ZN(n1822) );
  INV_X1 U2577 ( .A(n40800), .ZN(n609) );
  INV_X1 U2578 ( .A(n43323), .ZN(n40801) );
  AND2_X1 U2580 ( .A1(n41480), .A2(n42062), .ZN(n1333) );
  INV_X1 U2582 ( .A(n41049), .ZN(n610) );
  AND3_X1 U2588 ( .A1(n40063), .A2(n40060), .A3(n40061), .ZN(n4806) );
  NOR2_X1 U2589 ( .A1(n37369), .A2(n37370), .ZN(n40062) );
  OR2_X1 U2591 ( .A1(n35452), .A2(n694), .ZN(n983) );
  INV_X1 U2593 ( .A(n38056), .ZN(n611) );
  INV_X1 U2595 ( .A(n37488), .ZN(n37442) );
  INV_X1 U2598 ( .A(n37730), .ZN(n612) );
  INV_X1 U2600 ( .A(n37809), .ZN(n39474) );
  NAND2_X1 U2601 ( .A1(n3708), .A2(n38664), .ZN(n39182) );
  BUF_X1 U2603 ( .A(n37900), .Z(n39430) );
  AND2_X1 U2606 ( .A1(n36616), .A2(n698), .ZN(n34929) );
  INV_X1 U2607 ( .A(n38291), .ZN(n613) );
  INV_X1 U2608 ( .A(n37983), .ZN(n37987) );
  INV_X1 U2611 ( .A(n34210), .ZN(n614) );
  INV_X1 U2612 ( .A(n36632), .ZN(n36313) );
  INV_X1 U2617 ( .A(n37753), .ZN(n615) );
  CLKBUF_X1 U2623 ( .A(n51418), .Z(n37544) );
  INV_X1 U2624 ( .A(n38722), .ZN(n616) );
  CLKBUF_X1 U2625 ( .A(n2176), .Z(n2177) );
  INV_X1 U2627 ( .A(n37439), .ZN(n617) );
  XNOR2_X1 U2628 ( .A(n6142), .B(n35807), .ZN(n34911) );
  XNOR2_X1 U2631 ( .A(n32626), .B(n702), .ZN(n36874) );
  XNOR2_X1 U2632 ( .A(n34121), .B(n6555), .ZN(n35247) );
  CLKBUF_X1 U2633 ( .A(n34121), .Z(n35595) );
  BUF_X1 U2635 ( .A(n33419), .Z(n37045) );
  BUF_X1 U2638 ( .A(n31967), .Z(n35070) );
  OAI211_X1 U2640 ( .C1(n30643), .C2(n724), .A(n920), .B(n30646), .ZN(n921) );
  NOR2_X1 U2642 ( .A1(n31999), .A2(n707), .ZN(n1870) );
  AND2_X1 U2647 ( .A1(n31484), .A2(n31273), .ZN(n3767) );
  INV_X2 U2648 ( .A(n31544), .ZN(n32665) );
  INV_X2 U2651 ( .A(n32841), .ZN(n32389) );
  OR2_X1 U2652 ( .A1(n32420), .A2(n726), .ZN(n31394) );
  AND2_X1 U2653 ( .A1(n32420), .A2(n726), .ZN(n32428) );
  INV_X1 U2655 ( .A(n31425), .ZN(n620) );
  AND2_X1 U2659 ( .A1(n723), .A2(n1385), .ZN(n32057) );
  INV_X1 U2660 ( .A(n30102), .ZN(n621) );
  INV_X1 U2663 ( .A(n32252), .ZN(n622) );
  INV_X1 U2669 ( .A(n32107), .ZN(n624) );
  AND3_X1 U2671 ( .A1(n30723), .A2(n30712), .A3(n731), .ZN(n29850) );
  AND2_X1 U2673 ( .A1(n30773), .A2(n26842), .ZN(n26840) );
  NOR2_X1 U2674 ( .A1(n735), .A2(n30202), .ZN(n1871) );
  AND2_X1 U2677 ( .A1(n26842), .A2(n30768), .ZN(n1898) );
  BUF_X1 U2679 ( .A(n26779), .Z(n27760) );
  AND3_X1 U2682 ( .A1(n29545), .A2(n29550), .A3(n743), .ZN(n26753) );
  INV_X1 U2683 ( .A(n29718), .ZN(n28189) );
  INV_X1 U2687 ( .A(n27132), .ZN(n27119) );
  OR2_X1 U2688 ( .A1(n29447), .A2(n2213), .ZN(n27828) );
  INV_X1 U2692 ( .A(n24354), .ZN(n30768) );
  BUF_X1 U2694 ( .A(n24570), .Z(n26891) );
  AND2_X1 U2695 ( .A1(n6403), .A2(n30431), .ZN(n29692) );
  INV_X1 U2698 ( .A(n30269), .ZN(n625) );
  INV_X1 U2700 ( .A(n746), .ZN(n1693) );
  OR2_X1 U2701 ( .A1(n29439), .A2(n747), .ZN(n27840) );
  AND2_X1 U2704 ( .A1(n24984), .A2(n6730), .ZN(n27951) );
  INV_X1 U2705 ( .A(n30244), .ZN(n626) );
  XNOR2_X1 U2707 ( .A(n6141), .B(n25393), .ZN(n29347) );
  INV_X1 U2710 ( .A(n447), .ZN(n27070) );
  INV_X1 U2711 ( .A(n5228), .ZN(n28641) );
  XNOR2_X1 U2715 ( .A(n26156), .B(n26157), .ZN(n27695) );
  INV_X1 U2716 ( .A(n29568), .ZN(n29542) );
  XNOR2_X1 U2720 ( .A(n1376), .B(n26233), .ZN(n29507) );
  XNOR2_X1 U2721 ( .A(n6644), .B(n6643), .ZN(n30256) );
  XNOR2_X1 U2722 ( .A(n25020), .B(n25021), .ZN(n27918) );
  XNOR2_X1 U2723 ( .A(n24263), .B(n26292), .ZN(n27372) );
  BUF_X1 U2724 ( .A(n24976), .Z(n28292) );
  BUF_X1 U2725 ( .A(n22762), .Z(n27502) );
  OR2_X1 U2726 ( .A1(n1710), .A2(n758), .ZN(n2004) );
  NAND4_X1 U2728 ( .A1(n23969), .A2(n23968), .A3(n23967), .A4(n23966), .ZN(
        n27501) );
  AOI22_X1 U2730 ( .A1(n23341), .A2(n22264), .B1(n21148), .B2(n21145), .ZN(
        n20869) );
  AND2_X1 U2732 ( .A1(n24157), .A2(n23833), .ZN(n24148) );
  INV_X1 U2733 ( .A(n24157), .ZN(n24159) );
  AND2_X1 U2734 ( .A1(n21060), .A2(n50977), .ZN(n1198) );
  AND2_X1 U2735 ( .A1(n23546), .A2(n17074), .ZN(n22272) );
  AND2_X1 U2736 ( .A1(n24246), .A2(n6744), .ZN(n1495) );
  NOR2_X1 U2737 ( .A1(n51355), .A2(n23207), .ZN(n23231) );
  INV_X1 U2738 ( .A(n23254), .ZN(n628) );
  AND3_X1 U2742 ( .A1(n23411), .A2(n452), .A3(n23409), .ZN(n1177) );
  INV_X1 U2745 ( .A(n25064), .ZN(n25057) );
  INV_X1 U2747 ( .A(n24247), .ZN(n6744) );
  BUF_X1 U2757 ( .A(n23229), .Z(n2102) );
  INV_X1 U2758 ( .A(n23827), .ZN(n630) );
  NOR2_X1 U2760 ( .A1(n17311), .A2(n770), .ZN(n2045) );
  NOR2_X1 U2762 ( .A1(n5083), .A2(n16986), .ZN(n19860) );
  BUF_X1 U2766 ( .A(n16994), .Z(n20215) );
  AND2_X1 U2768 ( .A1(n18063), .A2(n1715), .ZN(n1714) );
  BUF_X1 U2770 ( .A(n17856), .Z(n20426) );
  INV_X1 U2774 ( .A(n21391), .ZN(n21397) );
  OR2_X2 U2776 ( .A1(n21354), .A2(n21605), .ZN(n20768) );
  CLKBUF_X1 U2777 ( .A(n17405), .Z(n21213) );
  NAND2_X1 U2778 ( .A1(n17484), .A2(n17576), .ZN(n18015) );
  XNOR2_X1 U2780 ( .A(n16531), .B(n16530), .ZN(n18357) );
  INV_X1 U2784 ( .A(n777), .ZN(n631) );
  INV_X1 U2787 ( .A(n17584), .ZN(n632) );
  INV_X1 U2791 ( .A(n20359), .ZN(n20435) );
  INV_X1 U2793 ( .A(n20488), .ZN(n634) );
  XNOR2_X1 U2794 ( .A(n1294), .B(n17675), .ZN(n19359) );
  XNOR2_X1 U2797 ( .A(n18146), .B(n16289), .ZN(n21251) );
  XNOR2_X1 U2798 ( .A(n8513), .B(n8512), .ZN(n16986) );
  BUF_X1 U2799 ( .A(n17887), .Z(n18409) );
  BUF_X2 U2800 ( .A(n18592), .Z(n635) );
  INV_X1 U2802 ( .A(n15018), .ZN(n636) );
  BUF_X2 U2803 ( .A(n18522), .Z(n637) );
  AND2_X1 U2807 ( .A1(n12204), .A2(n784), .ZN(n13574) );
  INV_X1 U2808 ( .A(n15437), .ZN(n15343) );
  AND2_X1 U2809 ( .A1(n13206), .A2(n2173), .ZN(n1579) );
  AND2_X1 U2810 ( .A1(n51657), .A2(n2173), .ZN(n1580) );
  NAND2_X1 U2821 ( .A1(n14411), .A2(n14393), .ZN(n14394) );
  INV_X1 U2824 ( .A(n2173), .ZN(n638) );
  INV_X2 U2825 ( .A(n13856), .ZN(n13853) );
  INV_X1 U2826 ( .A(n15163), .ZN(n15173) );
  INV_X1 U2833 ( .A(n14294), .ZN(n13588) );
  INV_X1 U2835 ( .A(n14228), .ZN(n639) );
  INV_X1 U2836 ( .A(n14106), .ZN(n640) );
  INV_X1 U2837 ( .A(n14712), .ZN(n14704) );
  BUF_X1 U2838 ( .A(n14643), .Z(n2114) );
  OR2_X2 U2840 ( .A1(n11536), .A2(n13914), .ZN(n11853) );
  INV_X1 U2842 ( .A(n13089), .ZN(n641) );
  OAI21_X1 U2845 ( .B1(n1999), .B2(n789), .A(n10457), .ZN(n10458) );
  AND2_X1 U2850 ( .A1(n11123), .A2(n802), .ZN(n1868) );
  BUF_X1 U2851 ( .A(n9022), .Z(n10272) );
  NOR2_X1 U2855 ( .A1(n9188), .A2(n796), .ZN(n1848) );
  OR2_X1 U2859 ( .A1(n12651), .A2(n796), .ZN(n10455) );
  NAND2_X1 U2860 ( .A1(n10037), .A2(n9465), .ZN(n10555) );
  NAND2_X1 U2864 ( .A1(n803), .A2(n10037), .ZN(n10539) );
  CLKBUF_X1 U2866 ( .A(n25898), .Z(n2602) );
  INV_X1 U2868 ( .A(n10147), .ZN(n9807) );
  CLKBUF_X1 U2871 ( .A(n8916), .Z(n12515) );
  CLKBUF_X1 U2873 ( .A(n8790), .Z(n10267) );
  OR2_X1 U2874 ( .A1(n804), .A2(n12301), .ZN(n9763) );
  CLKBUF_X1 U2875 ( .A(n42630), .Z(n2599) );
  BUF_X1 U2876 ( .A(n9459), .Z(n10540) );
  BUF_X1 U2877 ( .A(n12651), .Z(n2227) );
  BUF_X1 U2880 ( .A(n8880), .Z(n12720) );
  CLKBUF_X1 U2884 ( .A(n9148), .Z(n9491) );
  BUF_X1 U2885 ( .A(Key[92]), .Z(n4624) );
  CLKBUF_X1 U2887 ( .A(Key[124]), .Z(n4518) );
  BUF_X1 U2889 ( .A(Key[110]), .Z(n49429) );
  CLKBUF_X2 U2891 ( .A(Key[77]), .Z(n48843) );
  CLKBUF_X1 U2892 ( .A(Key[38]), .Z(n3336) );
  CLKBUF_X1 U2893 ( .A(Key[78]), .Z(n1336) );
  CLKBUF_X1 U2894 ( .A(Key[23]), .Z(n4636) );
  BUF_X1 U2895 ( .A(Key[182]), .Z(n4909) );
  BUF_X1 U2896 ( .A(Key[14]), .Z(n4723) );
  CLKBUF_X1 U2898 ( .A(Key[189]), .Z(n2117) );
  BUF_X1 U2899 ( .A(Key[32]), .Z(n4121) );
  BUF_X1 U2900 ( .A(Key[158]), .Z(n4641) );
  BUF_X1 U2903 ( .A(Key[176]), .Z(n4746) );
  CLKBUF_X1 U2905 ( .A(Key[74]), .Z(n4650) );
  BUF_X1 U2907 ( .A(Key[177]), .Z(n4565) );
  BUF_X1 U2910 ( .A(Key[84]), .Z(n4752) );
  BUF_X1 U2912 ( .A(Key[80]), .Z(n4939) );
  CLKBUF_X1 U2913 ( .A(Key[152]), .Z(n4076) );
  BUF_X1 U2917 ( .A(Key[35]), .Z(n4837) );
  BUF_X1 U2918 ( .A(Key[174]), .Z(n4325) );
  BUF_X1 U2919 ( .A(Key[155]), .Z(n4487) );
  BUF_X1 U2920 ( .A(Key[185]), .Z(n4890) );
  BUF_X1 U2921 ( .A(Key[95]), .Z(n4884) );
  BUF_X1 U2922 ( .A(Key[119]), .Z(n4879) );
  BUF_X1 U2924 ( .A(Key[83]), .Z(n4653) );
  BUF_X1 U2925 ( .A(Key[59]), .Z(n4826) );
  CLKBUF_X1 U2926 ( .A(Key[101]), .Z(n1313) );
  BUF_X1 U2927 ( .A(Key[41]), .Z(n4537) );
  CLKBUF_X1 U2928 ( .A(Key[93]), .Z(n4423) );
  BUF_X1 U2929 ( .A(Key[105]), .Z(n4868) );
  BUF_X1 U2931 ( .A(Key[45]), .Z(n4501) );
  BUF_X1 U2932 ( .A(Key[81]), .Z(n4883) );
  CLKBUF_X1 U2933 ( .A(Key[17]), .Z(n33221) );
  BUF_X1 U2934 ( .A(Key[29]), .Z(n4720) );
  BUF_X1 U2935 ( .A(Key[51]), .Z(n4637) );
  BUF_X1 U2936 ( .A(Key[135]), .Z(n4605) );
  BUF_X1 U2937 ( .A(Key[123]), .Z(n4157) );
  BUF_X1 U2938 ( .A(Key[125]), .Z(n3481) );
  BUF_X1 U2939 ( .A(Key[5]), .Z(n4535) );
  BUF_X1 U2941 ( .A(Key[39]), .Z(n4937) );
  BUF_X1 U2942 ( .A(Key[151]), .Z(n4788) );
  CLKBUF_X1 U2943 ( .A(Key[109]), .Z(n2230) );
  BUF_X1 U2944 ( .A(Key[191]), .Z(n4668) );
  BUF_X1 U2945 ( .A(Key[148]), .Z(n4676) );
  BUF_X1 U2946 ( .A(Key[100]), .Z(n49109) );
  BUF_X1 U2947 ( .A(Key[76]), .Z(n48814) );
  BUF_X1 U2948 ( .A(Key[52]), .Z(n4827) );
  BUF_X1 U2950 ( .A(Key[22]), .Z(n4628) );
  BUF_X1 U2953 ( .A(Key[10]), .Z(n4835) );
  BUF_X1 U2954 ( .A(Key[130]), .Z(n4733) );
  BUF_X1 U2955 ( .A(Key[19]), .Z(n4429) );
  BUF_X1 U2956 ( .A(Key[183]), .Z(n4940) );
  BUF_X1 U2957 ( .A(Key[7]), .Z(n47268) );
  CLKBUF_X1 U2959 ( .A(Key[28]), .Z(n4502) );
  BUF_X1 U2960 ( .A(Key[103]), .Z(n4895) );
  BUF_X1 U2961 ( .A(Key[112]), .Z(n4803) );
  BUF_X1 U2962 ( .A(Key[4]), .Z(n4237) );
  BUF_X1 U2963 ( .A(Key[172]), .Z(n4864) );
  BUF_X1 U2964 ( .A(Key[64]), .Z(n4737) );
  BUF_X1 U2965 ( .A(Key[137]), .Z(n49937) );
  CLKBUF_X1 U2967 ( .A(Key[145]), .Z(n4897) );
  CLKBUF_X1 U2968 ( .A(Key[143]), .Z(n4286) );
  BUF_X1 U2969 ( .A(Key[107]), .Z(n4177) );
  BUF_X1 U2970 ( .A(Key[184]), .Z(n4526) );
  BUF_X1 U2971 ( .A(Key[89]), .Z(n4874) );
  BUF_X1 U2972 ( .A(Key[149]), .Z(n4618) );
  BUF_X1 U2973 ( .A(Key[13]), .Z(n4908) );
  BUF_X1 U2975 ( .A(Key[169]), .Z(n4838) );
  BUF_X1 U2977 ( .A(Key[49]), .Z(n4916) );
  CLKBUF_X1 U2978 ( .A(Key[66]), .Z(n4490) );
  CLKBUF_X1 U2979 ( .A(Key[109]), .Z(n2231) );
  CLKBUF_X1 U2980 ( .A(Key[94]), .Z(n4275) );
  CLKBUF_X1 U2981 ( .A(Key[54]), .Z(n2947) );
  BUF_X1 U2983 ( .A(Key[179]), .Z(n4627) );
  CLKBUF_X1 U2984 ( .A(Key[82]), .Z(n4026) );
  BUF_X1 U2985 ( .A(Key[61]), .Z(n4691) );
  XNOR2_X1 U2986 ( .A(n4213), .B(Key[93]), .ZN(n43368) );
  BUF_X1 U2987 ( .A(Key[25]), .Z(n4836) );
  BUF_X1 U2988 ( .A(Key[181]), .Z(n4667) );
  BUF_X1 U2990 ( .A(Key[1]), .Z(n4926) );
  BUF_X1 U2991 ( .A(Key[139]), .Z(n4655) );
  BUF_X1 U2993 ( .A(Key[99]), .Z(n4554) );
  BUF_X1 U2995 ( .A(Key[186]), .Z(n4415) );
  BUF_X1 U2998 ( .A(Key[108]), .Z(n49414) );
  BUF_X1 U2999 ( .A(Key[132]), .Z(n42769) );
  CLKBUF_X1 U3000 ( .A(Key[150]), .Z(n4296) );
  BUF_X1 U3001 ( .A(Key[90]), .Z(n4639) );
  BUF_X1 U3002 ( .A(Key[96]), .Z(n4597) );
  BUF_X1 U3003 ( .A(Key[43]), .Z(n4869) );
  BUF_X1 U3005 ( .A(Key[138]), .Z(n4880) );
  BUF_X1 U3007 ( .A(Key[72]), .Z(n4536) );
  BUF_X1 U3008 ( .A(Key[102]), .Z(n4665) );
  BUF_X1 U3011 ( .A(Key[126]), .Z(n4705) );
  BUF_X1 U3012 ( .A(Key[127]), .Z(n49790) );
  BUF_X1 U3013 ( .A(Key[8]), .Z(n4647) );
  BUF_X1 U3014 ( .A(Key[120]), .Z(n4755) );
  BUF_X1 U3015 ( .A(Key[63]), .Z(n4666) );
  BUF_X1 U3017 ( .A(Key[68]), .Z(n4558) );
  CLKBUF_X1 U3018 ( .A(Key[159]), .Z(n3367) );
  BUF_X1 U3022 ( .A(Key[164]), .Z(n4800) );
  BUF_X1 U3023 ( .A(Key[97]), .Z(n4865) );
  BUF_X1 U3024 ( .A(Key[79]), .Z(n4824) );
  BUF_X1 U3025 ( .A(Key[144]), .Z(n4651) );
  BUF_X1 U3026 ( .A(Key[87]), .Z(n4885) );
  BUF_X1 U3027 ( .A(Key[44]), .Z(n4589) );
  BUF_X1 U3028 ( .A(Key[58]), .Z(n4654) );
  BUF_X1 U3029 ( .A(Key[187]), .Z(n4934) );
  CLKBUF_X1 U3030 ( .A(Key[117]), .Z(n4213) );
  BUF_X1 U3031 ( .A(Key[73]), .Z(n4923) );
  CLKBUF_X1 U3033 ( .A(Key[15]), .Z(n4587) );
  INV_X1 U3034 ( .A(n9926), .ZN(n643) );
  BUF_X1 U3036 ( .A(Key[168]), .Z(n4706) );
  BUF_X1 U3038 ( .A(Key[46]), .Z(n4048) );
  BUF_X1 U3039 ( .A(Key[16]), .Z(n47679) );
  CLKBUF_X1 U3041 ( .A(Key[190]), .Z(n4599) );
  NOR2_X1 U3042 ( .A1(n1736), .A2(n1583), .ZN(n1734) );
  AND4_X1 U3043 ( .A1(n48812), .A2(n5391), .A3(n4923), .A4(n5392), .ZN(n1729)
         );
  AND2_X1 U3044 ( .A1(n48342), .A2(n48343), .ZN(n1750) );
  OAI21_X1 U3045 ( .B1(n50651), .B2(n1468), .A(n50679), .ZN(n50660) );
  AND3_X1 U3046 ( .A1(n49508), .A2(n338), .A3(n4572), .ZN(n1636) );
  NOR3_X1 U3047 ( .A1(n1584), .A2(n2034), .A3(n52090), .ZN(n1583) );
  AND3_X1 U3048 ( .A1(n50823), .A2(n1445), .A3(n1444), .ZN(n1443) );
  OR2_X1 U3049 ( .A1(n1735), .A2(n45743), .ZN(n48812) );
  AND3_X1 U3050 ( .A1(n342), .A2(n50467), .A3(n1189), .ZN(n1312) );
  OAI21_X1 U3052 ( .B1(n49350), .B2(n51308), .A(n49367), .ZN(n49288) );
  INV_X1 U3053 ( .A(n50475), .ZN(n1311) );
  OAI21_X1 U3054 ( .B1(n52434), .B2(n1585), .A(n48821), .ZN(n48826) );
  OR2_X1 U3055 ( .A1(n43416), .A2(n1976), .ZN(n45734) );
  AND3_X1 U3056 ( .A1(n45984), .A2(n45982), .A3(n45981), .ZN(n3299) );
  INV_X1 U3057 ( .A(n50227), .ZN(n50191) );
  AND2_X1 U3058 ( .A1(n45753), .A2(n45754), .ZN(n1737) );
  AOI21_X1 U3059 ( .B1(n994), .B2(n48759), .A(n340), .ZN(n47438) );
  OR2_X1 U3063 ( .A1(n47728), .A2(n1994), .ZN(n47742) );
  NOR2_X1 U3064 ( .A1(n50906), .A2(n51298), .ZN(n1757) );
  INV_X1 U3065 ( .A(n47592), .ZN(n1187) );
  OR2_X1 U3067 ( .A1(n46934), .A2(n46933), .ZN(n49036) );
  AND2_X1 U3068 ( .A1(n50955), .A2(n50929), .ZN(n1756) );
  NOR2_X1 U3070 ( .A1(n49508), .A2(n49529), .ZN(n7209) );
  OR2_X1 U3071 ( .A1(n50949), .A2(n47391), .ZN(n50909) );
  AND2_X1 U3072 ( .A1(n47589), .A2(n8449), .ZN(n47622) );
  OR2_X1 U3073 ( .A1(n51400), .A2(n47586), .ZN(n47588) );
  OR2_X1 U3074 ( .A1(n562), .A2(n8508), .ZN(n50088) );
  INV_X1 U3076 ( .A(n48847), .ZN(n48846) );
  AND2_X1 U3077 ( .A1(n50681), .A2(n50734), .ZN(n50718) );
  AND2_X1 U3078 ( .A1(n6665), .A2(n50533), .ZN(n50539) );
  INV_X1 U3079 ( .A(n47620), .ZN(n47592) );
  OR2_X1 U3081 ( .A1(n50451), .A2(n4692), .ZN(n50440) );
  INV_X1 U3082 ( .A(n50700), .ZN(n50675) );
  OR2_X1 U3083 ( .A1(n47674), .A2(n47686), .ZN(n1089) );
  AND2_X1 U3084 ( .A1(n47528), .A2(n51289), .ZN(n47541) );
  NOR2_X1 U3085 ( .A1(n3782), .A2(n48908), .ZN(n48915) );
  AND2_X1 U3087 ( .A1(n49534), .A2(n2193), .ZN(n4984) );
  INV_X1 U3088 ( .A(n49491), .ZN(n45021) );
  AND4_X1 U3089 ( .A1(n1467), .A2(n50716), .A3(n50681), .A4(n51367), .ZN(n1468) );
  OR2_X1 U3091 ( .A1(n48834), .A2(n48808), .ZN(n1735) );
  INV_X1 U3092 ( .A(n47743), .ZN(n645) );
  INV_X1 U3093 ( .A(n48116), .ZN(n646) );
  OR2_X1 U3094 ( .A1(n50435), .A2(n50357), .ZN(n50411) );
  NOR2_X1 U3095 ( .A1(n567), .A2(n47989), .ZN(n47996) );
  AND2_X1 U3096 ( .A1(n47824), .A2(n47873), .ZN(n47866) );
  INV_X1 U3097 ( .A(n49534), .ZN(n49508) );
  INV_X1 U3099 ( .A(n49285), .ZN(n49350) );
  OR2_X1 U3100 ( .A1(n45739), .A2(n45711), .ZN(n48831) );
  AND2_X1 U3101 ( .A1(n48888), .A2(n48919), .ZN(n48898) );
  INV_X1 U3102 ( .A(n48853), .ZN(n48913) );
  AND2_X1 U3104 ( .A1(n48853), .A2(n51689), .ZN(n48847) );
  OR2_X1 U3105 ( .A1(n48944), .A2(n48935), .ZN(n48971) );
  NOR2_X1 U3106 ( .A1(n2034), .A2(n45739), .ZN(n48805) );
  NOR2_X1 U3107 ( .A1(n51291), .A2(n655), .ZN(n48695) );
  BUF_X1 U3108 ( .A(n45739), .Z(n45752) );
  INV_X1 U3109 ( .A(n49119), .ZN(n1155) );
  INV_X1 U3110 ( .A(n49592), .ZN(n647) );
  INV_X1 U3111 ( .A(n51687), .ZN(n3782) );
  INV_X1 U3114 ( .A(n48792), .ZN(n2033) );
  NOR2_X1 U3116 ( .A1(n49070), .A2(n44772), .ZN(n49066) );
  BUF_X1 U3117 ( .A(n42192), .Z(n47873) );
  OR2_X1 U3118 ( .A1(n50542), .A2(n50550), .ZN(n50495) );
  AND2_X1 U3119 ( .A1(n50486), .A2(n50465), .ZN(n1190) );
  INV_X1 U3120 ( .A(n47991), .ZN(n648) );
  INV_X1 U3122 ( .A(n42192), .ZN(n1420) );
  INV_X1 U3123 ( .A(n42192), .ZN(n47842) );
  NOR2_X1 U3124 ( .A1(n372), .A2(n47857), .ZN(n47824) );
  INV_X1 U3127 ( .A(n50681), .ZN(n649) );
  NOR2_X1 U3129 ( .A1(n47987), .A2(n47945), .ZN(n47928) );
  AND2_X1 U3130 ( .A1(n1945), .A2(n315), .ZN(n48565) );
  INV_X1 U3131 ( .A(n50727), .ZN(n50734) );
  OAI211_X1 U3132 ( .C1(n45594), .C2(n40180), .A(n40179), .B(n1634), .ZN(
        n42192) );
  INV_X1 U3134 ( .A(n48652), .ZN(n48640) );
  INV_X1 U3135 ( .A(n49569), .ZN(n49598) );
  BUF_X1 U3137 ( .A(n42810), .Z(n48973) );
  INV_X1 U3138 ( .A(n48051), .ZN(n650) );
  INV_X1 U3140 ( .A(n47841), .ZN(n651) );
  NOR2_X1 U3141 ( .A1(n47891), .A2(n1718), .ZN(n1717) );
  INV_X1 U3143 ( .A(n50552), .ZN(n1151) );
  INV_X1 U3146 ( .A(n50780), .ZN(n50808) );
  OR2_X1 U3147 ( .A1(n46173), .A2(n49916), .ZN(n49928) );
  AND4_X1 U3148 ( .A1(n46601), .A2(n46600), .A3(n3304), .A4(n7680), .ZN(n7678)
         );
  CLKBUF_X1 U3149 ( .A(n45872), .Z(n47721) );
  INV_X1 U3150 ( .A(n49932), .ZN(n652) );
  OAI211_X1 U3154 ( .C1(n46898), .C2(n46897), .A(n46896), .B(n46895), .ZN(
        n50854) );
  INV_X1 U3155 ( .A(n1718), .ZN(n1392) );
  OAI21_X1 U3156 ( .B1(n40178), .B2(n48443), .A(n40177), .ZN(n1634) );
  INV_X1 U3157 ( .A(n44705), .ZN(n1722) );
  INV_X1 U3158 ( .A(n49037), .ZN(n6389) );
  AND3_X1 U3162 ( .A1(n47351), .A2(n47350), .A3(n1009), .ZN(n47365) );
  AND3_X1 U3166 ( .A1(n44272), .A2(n44271), .A3(n44273), .ZN(n1103) );
  OAI21_X2 U3167 ( .B1(n50395), .B2(n50394), .A(n50393), .ZN(n50433) );
  INV_X1 U3169 ( .A(n49899), .ZN(n654) );
  AND4_X1 U3170 ( .A1(n5851), .A2(n43686), .A3(n5852), .A4(n43689), .ZN(n5848)
         );
  INV_X1 U3171 ( .A(n48698), .ZN(n655) );
  NOR2_X1 U3173 ( .A1(n47082), .A2(n47083), .ZN(n47084) );
  AND2_X1 U3175 ( .A1(n1588), .A2(n45144), .ZN(n6588) );
  INV_X1 U3176 ( .A(n46521), .ZN(n2017) );
  AOI21_X1 U3177 ( .B1(n2427), .B2(n5163), .A(n5162), .ZN(n6958) );
  OR2_X1 U3178 ( .A1(n882), .A2(n881), .ZN(n46418) );
  AND3_X1 U3179 ( .A1(n49181), .A2(n2875), .A3(n2874), .ZN(n8020) );
  AND2_X1 U3180 ( .A1(n44575), .A2(n47112), .ZN(n1199) );
  AND2_X1 U3181 ( .A1(n44645), .A2(n42176), .ZN(n1718) );
  AND2_X1 U3182 ( .A1(n1474), .A2(n1473), .ZN(n1623) );
  INV_X1 U3184 ( .A(n2040), .ZN(n1664) );
  AND3_X1 U3185 ( .A1(n916), .A2(n41917), .A3(n41916), .ZN(n914) );
  OR2_X1 U3187 ( .A1(n47908), .A2(n46635), .ZN(n2039) );
  OAI21_X1 U3190 ( .B1(n43087), .B2(n43088), .A(n43086), .ZN(n2001) );
  NOR2_X1 U3192 ( .A1(n46337), .A2(n48166), .ZN(n46518) );
  NOR2_X1 U3195 ( .A1(n7176), .A2(n7175), .ZN(n49971) );
  AND2_X1 U3196 ( .A1(n5844), .A2(n45525), .ZN(n1720) );
  AND2_X1 U3197 ( .A1(n46725), .A2(n46721), .ZN(n1588) );
  OR2_X1 U3198 ( .A1(n45066), .A2(n46854), .ZN(n46852) );
  AND2_X1 U3199 ( .A1(n45031), .A2(n51359), .ZN(n1508) );
  AOI21_X1 U3200 ( .B1(n1478), .B2(n5506), .A(n1475), .ZN(n1474) );
  OAI21_X1 U3201 ( .B1(n46033), .B2(n7724), .A(n43091), .ZN(n2002) );
  OR2_X1 U3202 ( .A1(n48550), .A2(n48551), .ZN(n1340) );
  AND2_X1 U3203 ( .A1(n4809), .A2(n4808), .ZN(n44699) );
  AND3_X1 U3204 ( .A1(n337), .A2(n46207), .A3(n46200), .ZN(n1602) );
  AND2_X1 U3205 ( .A1(n5429), .A2(n48457), .ZN(n1972) );
  OR2_X1 U3206 ( .A1(n43444), .A2(n45961), .ZN(n43445) );
  AND2_X1 U3207 ( .A1(n45790), .A2(n46589), .ZN(n46584) );
  NAND2_X1 U3208 ( .A1(n50366), .A2(n44595), .ZN(n50372) );
  AND4_X1 U3209 ( .A1(n49977), .A2(n47354), .A3(n49972), .A4(n49990), .ZN(
        n1475) );
  OR2_X1 U3210 ( .A1(n2119), .A2(n48208), .ZN(n1101) );
  AND2_X1 U3212 ( .A1(n47151), .A2(n2178), .ZN(n47000) );
  NOR2_X1 U3213 ( .A1(n8569), .A2(n46444), .ZN(n48457) );
  OR2_X1 U3215 ( .A1(n46434), .A2(n51732), .ZN(n45618) );
  AND2_X1 U3216 ( .A1(n49651), .A2(n1806), .ZN(n45961) );
  OR2_X1 U3217 ( .A1(n47069), .A2(n46772), .ZN(n46814) );
  AND2_X1 U3218 ( .A1(n42365), .A2(n46204), .ZN(n6942) );
  NOR2_X1 U3221 ( .A1(n1943), .A2(n48165), .ZN(n48169) );
  BUF_X1 U3222 ( .A(n45773), .Z(n46654) );
  AND2_X1 U3223 ( .A1(n46693), .A2(n46614), .ZN(n1507) );
  AND2_X1 U3224 ( .A1(n48179), .A2(n48165), .ZN(n1752) );
  OR2_X1 U3225 ( .A1(n49150), .A2(n49148), .ZN(n1161) );
  OR2_X1 U3226 ( .A1(n46731), .A2(n46735), .ZN(n46555) );
  NOR2_X1 U3228 ( .A1(n45757), .A2(n1655), .ZN(n44867) );
  INV_X1 U3230 ( .A(n7777), .ZN(n47153) );
  OR2_X1 U3231 ( .A1(n40175), .A2(n6674), .ZN(n1643) );
  NOR2_X1 U3232 ( .A1(n49972), .A2(n49990), .ZN(n43178) );
  AND2_X1 U3233 ( .A1(n46714), .A2(n46572), .ZN(n46574) );
  INV_X1 U3234 ( .A(n40175), .ZN(n1645) );
  AND2_X1 U3235 ( .A1(n42177), .A2(n44640), .ZN(n45521) );
  AND2_X1 U3239 ( .A1(n49978), .A2(n49980), .ZN(n1010) );
  NOR2_X1 U3240 ( .A1(n1654), .A2(n46637), .ZN(n46628) );
  AND3_X1 U3241 ( .A1(n2726), .A2(n49663), .A3(n51733), .ZN(n1806) );
  INV_X1 U3242 ( .A(n3610), .ZN(n50361) );
  AND2_X1 U3244 ( .A1(n44583), .A2(n50270), .ZN(n50262) );
  NOR2_X1 U3245 ( .A1(n48474), .A2(n48491), .ZN(n48254) );
  OR2_X1 U3246 ( .A1(n47044), .A2(n5237), .ZN(n50279) );
  BUF_X1 U3247 ( .A(n41470), .Z(n46589) );
  NAND2_X1 U3248 ( .A1(n47128), .A2(n45772), .ZN(n46859) );
  AND2_X1 U3249 ( .A1(n47309), .A2(n50390), .ZN(n47019) );
  OR2_X1 U3251 ( .A1(n50001), .A2(n50010), .ZN(n1811) );
  OR2_X1 U3252 ( .A1(n45551), .A2(n44992), .ZN(n48208) );
  AND2_X1 U3253 ( .A1(n46908), .A2(n51513), .ZN(n46917) );
  AOI21_X1 U3258 ( .B1(n1586), .B2(n49177), .A(n44784), .ZN(n45211) );
  INV_X1 U3259 ( .A(n46395), .ZN(n991) );
  AND2_X1 U3260 ( .A1(n46744), .A2(n46747), .ZN(n46735) );
  INV_X1 U3261 ( .A(n49688), .ZN(n656) );
  BUF_X1 U3262 ( .A(n45628), .Z(n48524) );
  AND2_X1 U3263 ( .A1(n46498), .A2(n46487), .ZN(n46387) );
  CLKBUF_X1 U3264 ( .A(n43688), .Z(n46998) );
  BUF_X1 U3266 ( .A(n39812), .Z(n48268) );
  INV_X1 U3269 ( .A(n43688), .ZN(n47151) );
  BUF_X1 U3270 ( .A(n42177), .Z(n45819) );
  INV_X1 U3271 ( .A(n44786), .ZN(n49177) );
  OR2_X1 U3272 ( .A1(n45848), .A2(n46904), .ZN(n46609) );
  AND2_X1 U3276 ( .A1(n49629), .A2(n49983), .ZN(n49973) );
  AND2_X1 U3278 ( .A1(n47126), .A2(n46649), .ZN(n46863) );
  CLKBUF_X1 U3281 ( .A(n42703), .Z(n46228) );
  NAND2_X1 U3282 ( .A1(n48481), .A2(n44678), .ZN(n48474) );
  OR2_X1 U3283 ( .A1(n46572), .A2(n405), .ZN(n46701) );
  INV_X1 U3285 ( .A(n46342), .ZN(n657) );
  INV_X1 U3288 ( .A(n47333), .ZN(n658) );
  NOR2_X1 U3290 ( .A1(n48201), .A2(n48213), .ZN(n44263) );
  INV_X1 U3293 ( .A(n46918), .ZN(n659) );
  OR2_X1 U3295 ( .A1(n44673), .A2(n48479), .ZN(n48251) );
  OR2_X1 U3296 ( .A1(n45848), .A2(n51359), .ZN(n46606) );
  CLKBUF_X1 U3297 ( .A(n52136), .Z(n46489) );
  NOR2_X1 U3298 ( .A1(n46498), .A2(n988), .ZN(n46403) );
  AND2_X1 U3299 ( .A1(n50325), .A2(n50010), .ZN(n47369) );
  NOR2_X1 U3301 ( .A1(n2742), .A2(n48416), .ZN(n6194) );
  NAND2_X1 U3302 ( .A1(n44409), .A2(n48479), .ZN(n48491) );
  XNOR2_X1 U3307 ( .A(n810), .B(n42282), .ZN(n44786) );
  CLKBUF_X1 U3308 ( .A(n42508), .Z(n48449) );
  INV_X1 U3310 ( .A(n39813), .ZN(n48259) );
  XNOR2_X1 U3311 ( .A(n43843), .B(n43844), .ZN(n47026) );
  XNOR2_X1 U3312 ( .A(n43964), .B(n43963), .ZN(n47341) );
  AND2_X1 U3313 ( .A1(n44118), .A2(n50280), .ZN(n50259) );
  XNOR2_X1 U3314 ( .A(n43982), .B(n43983), .ZN(n47044) );
  XNOR2_X1 U3315 ( .A(n1466), .B(n43659), .ZN(n43688) );
  XNOR2_X1 U3316 ( .A(n7696), .B(n42882), .ZN(n49231) );
  INV_X1 U3317 ( .A(n46828), .ZN(n661) );
  INV_X1 U3318 ( .A(n988), .ZN(n46487) );
  BUF_X1 U3319 ( .A(n43432), .Z(n49208) );
  BUF_X1 U3322 ( .A(n43278), .Z(n49656) );
  XNOR2_X1 U3325 ( .A(n4750), .B(n2303), .ZN(n46899) );
  INV_X1 U3328 ( .A(n46510), .ZN(n48404) );
  CLKBUF_X1 U3329 ( .A(n42081), .Z(n45818) );
  XNOR2_X1 U3331 ( .A(n43829), .B(n43828), .ZN(n50350) );
  INV_X1 U3333 ( .A(n45209), .ZN(n664) );
  XNOR2_X1 U3334 ( .A(n43630), .B(n43629), .ZN(n46996) );
  INV_X1 U3335 ( .A(n44678), .ZN(n665) );
  XNOR2_X1 U3336 ( .A(n42364), .B(n42363), .ZN(n46196) );
  INV_X1 U3338 ( .A(n46197), .ZN(n666) );
  XNOR2_X1 U3341 ( .A(n1174), .B(n42766), .ZN(n988) );
  XNOR2_X1 U3342 ( .A(n41787), .B(n44479), .ZN(n6717) );
  XNOR2_X1 U3343 ( .A(n42916), .B(n42348), .ZN(n1599) );
  XNOR2_X1 U3344 ( .A(n43534), .B(n43193), .ZN(n1033) );
  INV_X1 U3345 ( .A(n47096), .ZN(n669) );
  XNOR2_X1 U3346 ( .A(n1598), .B(n42666), .ZN(n44022) );
  XNOR2_X1 U3347 ( .A(n45432), .B(n43194), .ZN(n1035) );
  XNOR2_X1 U3349 ( .A(n44512), .B(n45389), .ZN(n42666) );
  XNOR2_X1 U3351 ( .A(n2103), .B(n42351), .ZN(n1598) );
  XNOR2_X1 U3353 ( .A(n1836), .B(n51408), .ZN(n45042) );
  BUF_X1 U3354 ( .A(n43027), .Z(n45059) );
  INV_X1 U3355 ( .A(n7608), .ZN(n43079) );
  XNOR2_X1 U3356 ( .A(n43920), .B(n50987), .ZN(n42786) );
  XNOR2_X1 U3357 ( .A(n7608), .B(n6031), .ZN(n43504) );
  INV_X1 U3358 ( .A(n42560), .ZN(n45041) );
  BUF_X1 U3360 ( .A(n44031), .Z(n2228) );
  NAND4_X1 U3363 ( .A1(n41456), .A2(n41455), .A3(n41454), .A4(n41453), .ZN(
        n42980) );
  XNOR2_X1 U3365 ( .A(n42560), .B(n310), .ZN(n1836) );
  NAND4_X1 U3372 ( .A1(n39897), .A2(n8755), .A3(n39896), .A4(n39898), .ZN(
        n42979) );
  AND4_X2 U3374 ( .A1(n6840), .A2(n37821), .A3(n7423), .A4(n37820), .ZN(n42560) );
  NAND3_X1 U3375 ( .A1(n41108), .A2(n6543), .A3(n6542), .ZN(n44951) );
  AND3_X1 U3378 ( .A1(n35009), .A2(n40508), .A3(n35007), .ZN(n3389) );
  AND2_X1 U3380 ( .A1(n1147), .A2(n1146), .ZN(n43671) );
  AND4_X1 U3381 ( .A1(n39994), .A2(n39993), .A3(n39992), .A4(n39991), .ZN(
        n44154) );
  NAND4_X1 U3382 ( .A1(n37615), .A2(n37614), .A3(n37613), .A4(n41020), .ZN(
        n42659) );
  AND3_X1 U3384 ( .A1(n39557), .A2(n39556), .A3(n39558), .ZN(n7122) );
  NAND4_X2 U3389 ( .A1(n1399), .A2(n1401), .A3(n41739), .A4(n41262), .ZN(
        n46138) );
  NAND4_X2 U3390 ( .A1(n39108), .A2(n39106), .A3(n39107), .A4(n39109), .ZN(
        n44373) );
  NOR2_X1 U3392 ( .A1(n41145), .A2(n2356), .ZN(n6549) );
  INV_X1 U3393 ( .A(n43928), .ZN(n672) );
  NAND3_X1 U3395 ( .A1(n40364), .A2(n40363), .A3(n40362), .ZN(n46143) );
  AND3_X1 U3396 ( .A1(n8197), .A2(n8196), .A3(n8195), .ZN(n4918) );
  AND2_X1 U3397 ( .A1(n37872), .A2(n37873), .ZN(n1216) );
  AND3_X1 U3399 ( .A1(n35725), .A2(n4068), .A3(n35723), .ZN(n5033) );
  AND2_X1 U3400 ( .A1(n2789), .A2(n1014), .ZN(n42089) );
  OR2_X1 U3401 ( .A1(n37845), .A2(n37844), .ZN(n39663) );
  AND4_X1 U3402 ( .A1(n40427), .A2(n40426), .A3(n40425), .A4(n40424), .ZN(
        n40434) );
  AND4_X1 U3403 ( .A1(n40144), .A2(n7153), .A3(n7155), .A4(n40145), .ZN(n4814)
         );
  AOI21_X1 U3405 ( .B1(n1388), .B2(n40396), .A(n39740), .ZN(n1102) );
  AND2_X1 U3407 ( .A1(n40405), .A2(n40395), .ZN(n1403) );
  AND3_X1 U3408 ( .A1(n38602), .A2(n38608), .A3(n38601), .ZN(n3463) );
  AND2_X1 U3409 ( .A1(n41738), .A2(n1400), .ZN(n1399) );
  AND4_X1 U3412 ( .A1(n5597), .A2(n5596), .A3(n40538), .A4(n40532), .ZN(n5595)
         );
  AND2_X1 U3413 ( .A1(n39162), .A2(n39163), .ZN(n1301) );
  AND3_X1 U3415 ( .A1(n36656), .A2(n36657), .A3(n36655), .ZN(n36661) );
  NOR3_X1 U3416 ( .A1(n7462), .A2(n40122), .A3(n2324), .ZN(n7461) );
  OAI21_X1 U3418 ( .B1(n1382), .B2(n40436), .A(n1380), .ZN(n39994) );
  OR2_X1 U3419 ( .A1(n38376), .A2(n38377), .ZN(n1388) );
  AOI22_X1 U3420 ( .A1(n34325), .A2(n40327), .B1(n39853), .B2(n40336), .ZN(
        n34327) );
  AND2_X1 U3421 ( .A1(n38373), .A2(n38372), .ZN(n1391) );
  AND3_X1 U3422 ( .A1(n39705), .A2(n38867), .A3(n3095), .ZN(n38884) );
  INV_X1 U3424 ( .A(n1705), .ZN(n41108) );
  AND2_X1 U3425 ( .A1(n40008), .A2(n1613), .ZN(n6887) );
  NOR2_X1 U3426 ( .A1(n40396), .A2(n40447), .ZN(n40462) );
  OR2_X1 U3427 ( .A1(n39788), .A2(n51377), .ZN(n38447) );
  OR2_X1 U3428 ( .A1(n42104), .A2(n38817), .ZN(n41789) );
  AND2_X1 U3430 ( .A1(n41735), .A2(n41736), .ZN(n1402) );
  AND2_X1 U3431 ( .A1(n3029), .A2(n6040), .ZN(n38932) );
  AND4_X1 U3432 ( .A1(n5421), .A2(n7861), .A3(n1126), .A4(n1125), .ZN(n3982)
         );
  AND2_X1 U3433 ( .A1(n40346), .A2(n40344), .ZN(n1358) );
  AND2_X1 U3434 ( .A1(n40968), .A2(n41372), .ZN(n41385) );
  AND3_X1 U3435 ( .A1(n7860), .A2(n1884), .A3(n1883), .ZN(n5422) );
  INV_X1 U3436 ( .A(n38850), .ZN(n38849) );
  AOI22_X1 U3437 ( .A1(n41900), .A2(n38606), .B1(n41327), .B2(n4876), .ZN(
        n38610) );
  OR2_X1 U3438 ( .A1(n42015), .A2(n41581), .ZN(n1067) );
  NOR2_X1 U3439 ( .A1(n40686), .A2(n40689), .ZN(n39682) );
  OR2_X1 U3440 ( .A1(n37865), .A2(n7117), .ZN(n38850) );
  INV_X1 U3441 ( .A(n1822), .ZN(n41148) );
  OR2_X1 U3442 ( .A1(n40590), .A2(n40776), .ZN(n1884) );
  INV_X1 U3443 ( .A(n41262), .ZN(n41731) );
  INV_X1 U3444 ( .A(n41339), .ZN(n40359) );
  OR2_X1 U3445 ( .A1(n38805), .A2(n43665), .ZN(n38808) );
  AND2_X1 U3446 ( .A1(n38352), .A2(n38353), .ZN(n1165) );
  OR2_X1 U3447 ( .A1(n4116), .A2(n39830), .ZN(n4115) );
  AOI22_X1 U3448 ( .A1(n41345), .A2(n41346), .B1(n41344), .B2(n41343), .ZN(
        n1408) );
  NOR2_X1 U3449 ( .A1(n40459), .A2(n39979), .ZN(n1382) );
  AND2_X1 U3450 ( .A1(n41511), .A2(n41581), .ZN(n41513) );
  OR2_X1 U3452 ( .A1(n40899), .A2(n2224), .ZN(n1070) );
  NAND2_X1 U3453 ( .A1(n930), .A2(n41797), .ZN(n932) );
  OR2_X1 U3454 ( .A1(n41348), .A2(n41352), .ZN(n41339) );
  NOR2_X1 U3455 ( .A1(n39912), .A2(n1874), .ZN(n39566) );
  INV_X1 U3457 ( .A(n42441), .ZN(n1334) );
  NOR2_X1 U3458 ( .A1(n40617), .A2(n41647), .ZN(n41978) );
  AND2_X1 U3460 ( .A1(n40388), .A2(n1931), .ZN(n40379) );
  INV_X1 U3463 ( .A(n42441), .ZN(n42042) );
  OR2_X1 U3464 ( .A1(n51853), .A2(n40972), .ZN(n40916) );
  INV_X1 U3465 ( .A(n42111), .ZN(n42112) );
  OR2_X1 U3466 ( .A1(n40377), .A2(n39834), .ZN(n39831) );
  NOR2_X1 U3468 ( .A1(n41638), .A2(n41646), .ZN(n1706) );
  AND2_X1 U3469 ( .A1(n42138), .A2(n42156), .ZN(n41751) );
  AND2_X1 U3470 ( .A1(n40868), .A2(n1984), .ZN(n40864) );
  AND3_X1 U3471 ( .A1(n41588), .A2(n41997), .A3(n42006), .ZN(n1133) );
  OR2_X1 U3473 ( .A1(n41144), .A2(n52083), .ZN(n1100) );
  OR2_X2 U3476 ( .A1(n6775), .A2(n6779), .ZN(n41039) );
  NOR2_X1 U3477 ( .A1(n42008), .A2(n41587), .ZN(n41512) );
  INV_X1 U3479 ( .A(n40500), .ZN(n41064) );
  OR2_X1 U3480 ( .A1(n38448), .A2(n51377), .ZN(n39785) );
  AND2_X1 U3481 ( .A1(n41348), .A2(n40740), .ZN(n41344) );
  INV_X1 U3482 ( .A(n1464), .ZN(n42442) );
  AND2_X1 U3483 ( .A1(n39738), .A2(n40450), .ZN(n1178) );
  AND2_X1 U3485 ( .A1(n39614), .A2(n41004), .ZN(n1261) );
  AND2_X1 U3489 ( .A1(n41211), .A2(n41212), .ZN(n8752) );
  AND2_X1 U3490 ( .A1(n41319), .A2(n41323), .ZN(n1562) );
  INV_X1 U3492 ( .A(n41111), .ZN(n41112) );
  NOR2_X1 U3493 ( .A1(n40295), .A2(n42062), .ZN(n1464) );
  INV_X1 U3495 ( .A(n42062), .ZN(n41481) );
  AND2_X1 U3497 ( .A1(n5318), .A2(n41323), .ZN(n41330) );
  OR2_X2 U3499 ( .A1(n8236), .A2(n6968), .ZN(n41902) );
  NOR2_X1 U3500 ( .A1(n41319), .A2(n40730), .ZN(n40373) );
  INV_X1 U3501 ( .A(n38810), .ZN(n42106) );
  NOR2_X1 U3502 ( .A1(n51684), .A2(n51950), .ZN(n930) );
  AND2_X1 U3503 ( .A1(n38810), .A2(n51950), .ZN(n40636) );
  INV_X1 U3504 ( .A(n40778), .ZN(n40775) );
  INV_X1 U3505 ( .A(n40943), .ZN(n41535) );
  AND2_X1 U3506 ( .A1(n38428), .A2(n39101), .ZN(n6884) );
  INV_X1 U3508 ( .A(n39674), .ZN(n40685) );
  OR2_X1 U3510 ( .A1(n41690), .A2(n5475), .ZN(n41698) );
  AND2_X1 U3513 ( .A1(n39097), .A2(n39103), .ZN(n1611) );
  OR2_X1 U3514 ( .A1(n35431), .A2(n35430), .ZN(n1614) );
  INV_X1 U3515 ( .A(n40240), .ZN(n676) );
  AND2_X1 U3516 ( .A1(n38810), .A2(n43666), .ZN(n42110) );
  NOR2_X1 U3518 ( .A1(n40250), .A2(n41938), .ZN(n42202) );
  INV_X1 U3519 ( .A(n41149), .ZN(n1931) );
  OR2_X2 U3520 ( .A1(n897), .A2(n5142), .ZN(n41702) );
  AND3_X1 U3523 ( .A1(n1741), .A2(n1740), .A3(n36526), .ZN(n36649) );
  AND2_X1 U3524 ( .A1(n41796), .A2(n43666), .ZN(n38817) );
  INV_X1 U3525 ( .A(n40525), .ZN(n678) );
  NAND4_X2 U3527 ( .A1(n5555), .A2(n5554), .A3(n5553), .A4(n39314), .ZN(n41670) );
  AND2_X1 U3528 ( .A1(n35182), .A2(n35181), .ZN(n7586) );
  NOR2_X1 U3529 ( .A1(n40869), .A2(n1984), .ZN(n40860) );
  INV_X1 U3530 ( .A(n42061), .ZN(n679) );
  INV_X1 U3531 ( .A(n40447), .ZN(n6851) );
  INV_X1 U3532 ( .A(n41975), .ZN(n6940) );
  INV_X1 U3533 ( .A(n42205), .ZN(n680) );
  INV_X1 U3534 ( .A(n40388), .ZN(n41143) );
  INV_X1 U3536 ( .A(n43666), .ZN(n40632) );
  INV_X1 U3538 ( .A(n39673), .ZN(n40676) );
  INV_X1 U3540 ( .A(n42138), .ZN(n42131) );
  INV_X1 U3541 ( .A(n40768), .ZN(n681) );
  INV_X1 U3542 ( .A(n52083), .ZN(n682) );
  INV_X1 U3543 ( .A(n41587), .ZN(n683) );
  NAND2_X1 U3546 ( .A1(n8355), .A2(n36418), .ZN(n39944) );
  INV_X1 U3549 ( .A(n39752), .ZN(n684) );
  AND3_X1 U3552 ( .A1(n34697), .A2(n34695), .A3(n34696), .ZN(n6766) );
  INV_X1 U3553 ( .A(n41796), .ZN(n41791) );
  AND2_X1 U3555 ( .A1(n36217), .A2(n36218), .ZN(n1949) );
  NAND4_X2 U3556 ( .A1(n37196), .A2(n37197), .A3(n4992), .A4(n4991), .ZN(
        n40453) );
  INV_X1 U3558 ( .A(n42054), .ZN(n686) );
  INV_X1 U3560 ( .A(n40526), .ZN(n1984) );
  AND2_X1 U3562 ( .A1(n31359), .A2(n7930), .ZN(n2948) );
  AND3_X1 U3564 ( .A1(n4887), .A2(n37936), .A3(n37935), .ZN(n1119) );
  NAND4_X2 U3565 ( .A1(n33275), .A2(n7976), .A3(n33277), .A4(n33276), .ZN(
        n40388) );
  AND4_X1 U3567 ( .A1(n1013), .A2(n38121), .A3(n38120), .A4(n1012), .ZN(n38129) );
  NOR2_X1 U3569 ( .A1(n36447), .A2(n36446), .ZN(n36509) );
  AND3_X1 U3570 ( .A1(n36419), .A2(n36417), .A3(n36416), .ZN(n8355) );
  INV_X1 U3571 ( .A(n42136), .ZN(n687) );
  AND4_X1 U3573 ( .A1(n36892), .A2(n36891), .A3(n36890), .A4(n36889), .ZN(
        n36893) );
  AND4_X1 U3574 ( .A1(n36346), .A2(n36333), .A3(n36347), .A4(n7396), .ZN(n7398) );
  AOI22_X1 U3576 ( .A1(n36538), .A2(n36537), .B1(n36536), .B2(n36535), .ZN(
        n36650) );
  AND3_X1 U3579 ( .A1(n38326), .A2(n37193), .A3(n4760), .ZN(n4992) );
  AND3_X1 U3580 ( .A1(n36409), .A2(n6263), .A3(n36408), .ZN(n36418) );
  AND3_X1 U3581 ( .A1(n1525), .A2(n34916), .A3(n1524), .ZN(n1530) );
  AND2_X1 U3584 ( .A1(n38256), .A2(n38628), .ZN(n37677) );
  AND4_X1 U3585 ( .A1(n36245), .A2(n5940), .A3(n37513), .A4(n36253), .ZN(n5939) );
  AND3_X1 U3587 ( .A1(n37567), .A2(n37565), .A3(n37566), .ZN(n1094) );
  AOI22_X1 U3588 ( .A1(n38331), .A2(n38332), .B1(n38333), .B2(n2714), .ZN(
        n38350) );
  AND2_X1 U3590 ( .A1(n1044), .A2(n36216), .ZN(n36213) );
  AND2_X1 U3591 ( .A1(n37444), .A2(n37445), .ZN(n852) );
  AND3_X1 U3592 ( .A1(n37641), .A2(n37642), .A3(n4352), .ZN(n37651) );
  AND3_X1 U3593 ( .A1(n35692), .A2(n35691), .A3(n35690), .ZN(n35698) );
  OAI211_X1 U3594 ( .C1(n36530), .C2(n5405), .A(n3068), .B(n36522), .ZN(n1742)
         );
  NOR2_X1 U3595 ( .A1(n34690), .A2(n39353), .ZN(n34696) );
  AND2_X1 U3597 ( .A1(n37429), .A2(n37427), .ZN(n840) );
  AND2_X1 U3598 ( .A1(n39312), .A2(n39313), .ZN(n5554) );
  OR2_X1 U3599 ( .A1(n38572), .A2(n1764), .ZN(n8577) );
  AND2_X1 U3600 ( .A1(n39488), .A2(n39471), .ZN(n39485) );
  AND3_X1 U3601 ( .A1(n35916), .A2(n35915), .A3(n37497), .ZN(n6222) );
  AND2_X1 U3602 ( .A1(n37512), .A2(n37513), .ZN(n5637) );
  AND3_X1 U3603 ( .A1(n37768), .A2(n37509), .A3(n37508), .ZN(n37514) );
  OR2_X1 U3604 ( .A1(n36037), .A2(n1914), .ZN(n34094) );
  OAI21_X1 U3605 ( .B1(n36590), .B2(n1692), .A(n1691), .ZN(n35874) );
  AND2_X1 U3606 ( .A1(n8459), .A2(n38328), .ZN(n37197) );
  AOI22_X1 U3607 ( .A1(n38260), .A2(n38261), .B1(n38263), .B2(n38262), .ZN(
        n38267) );
  AOI22_X1 U3608 ( .A1(n36142), .A2(n2245), .B1(n38545), .B2(n2719), .ZN(
        n31360) );
  INV_X1 U3609 ( .A(n38570), .ZN(n688) );
  INV_X1 U3610 ( .A(n37916), .ZN(n37917) );
  OR2_X1 U3611 ( .A1(n37766), .A2(n1569), .ZN(n1528) );
  INV_X1 U3612 ( .A(n38339), .ZN(n1605) );
  AND3_X1 U3613 ( .A1(n36188), .A2(n37778), .A3(n36186), .ZN(n34690) );
  AND2_X1 U3614 ( .A1(n36589), .A2(n36045), .ZN(n1692) );
  INV_X1 U3618 ( .A(n35942), .ZN(n39351) );
  INV_X1 U3619 ( .A(n34938), .ZN(n34947) );
  INV_X1 U3620 ( .A(n38467), .ZN(n38119) );
  AND2_X1 U3621 ( .A1(n37980), .A2(n37983), .ZN(n36535) );
  AND2_X1 U3622 ( .A1(n37804), .A2(n39472), .ZN(n39484) );
  AOI21_X1 U3624 ( .B1(n1005), .B2(n37594), .A(n1004), .ZN(n1003) );
  NOR2_X1 U3625 ( .A1(n38056), .A2(n36338), .ZN(n38131) );
  AND2_X1 U3626 ( .A1(n39335), .A2(n36199), .ZN(n39353) );
  INV_X1 U3628 ( .A(n37884), .ZN(n39401) );
  NOR2_X1 U3629 ( .A1(n1950), .A2(n38484), .ZN(n6318) );
  NOR2_X1 U3630 ( .A1(n34963), .A2(n1360), .ZN(n34186) );
  AND2_X1 U3631 ( .A1(n39208), .A2(n39426), .ZN(n902) );
  INV_X1 U3632 ( .A(n38108), .ZN(n1974) );
  INV_X1 U3633 ( .A(n39473), .ZN(n1582) );
  OR2_X1 U3634 ( .A1(n37517), .A2(n38493), .ZN(n33558) );
  AND2_X1 U3635 ( .A1(n34676), .A2(n37557), .ZN(n37562) );
  AND2_X1 U3636 ( .A1(n38092), .A2(n36627), .ZN(n36640) );
  INV_X1 U3637 ( .A(n7916), .ZN(n2049) );
  NAND2_X1 U3638 ( .A1(n35010), .A2(n38132), .ZN(n38056) );
  INV_X1 U3639 ( .A(n35452), .ZN(n37594) );
  AND2_X1 U3642 ( .A1(n33174), .A2(n34210), .ZN(n38029) );
  BUF_X1 U3647 ( .A(n34210), .Z(n35156) );
  AND2_X1 U3649 ( .A1(n38731), .A2(n38313), .ZN(n8077) );
  AND2_X1 U3652 ( .A1(n52054), .A2(n37774), .ZN(n1469) );
  INV_X1 U3653 ( .A(n1006), .ZN(n36231) );
  AND2_X1 U3654 ( .A1(n39245), .A2(n38701), .ZN(n4257) );
  OR2_X1 U3655 ( .A1(n36225), .A2(n1006), .ZN(n1005) );
  OR2_X1 U3656 ( .A1(n52191), .A2(n38483), .ZN(n38108) );
  INV_X1 U3658 ( .A(n37757), .ZN(n1569) );
  INV_X1 U3660 ( .A(n37762), .ZN(n1570) );
  NOR2_X1 U3663 ( .A1(n39464), .A2(n39438), .ZN(n1843) );
  INV_X1 U3664 ( .A(n2089), .ZN(n39347) );
  AND2_X1 U3666 ( .A1(n37762), .A2(n33370), .ZN(n3529) );
  OR2_X1 U3668 ( .A1(n38635), .A2(n38630), .ZN(n37688) );
  CLKBUF_X1 U3670 ( .A(n35927), .Z(n37538) );
  XNOR2_X1 U3671 ( .A(n35980), .B(n37596), .ZN(n37595) );
  AND2_X1 U3673 ( .A1(n35890), .A2(n38329), .ZN(n38345) );
  AND2_X1 U3674 ( .A1(n36047), .A2(n36590), .ZN(n36581) );
  INV_X1 U3676 ( .A(n38702), .ZN(n38700) );
  CLKBUF_X1 U3677 ( .A(n33562), .Z(n38492) );
  OR2_X1 U3678 ( .A1(n38593), .A2(n36122), .ZN(n37568) );
  NOR2_X1 U3679 ( .A1(n51334), .A2(n37646), .ZN(n37635) );
  INV_X1 U3682 ( .A(n37385), .ZN(n37387) );
  NAND2_X1 U3683 ( .A1(n35457), .A2(n35973), .ZN(n35452) );
  INV_X1 U3684 ( .A(n38566), .ZN(n689) );
  OR2_X1 U3689 ( .A1(n5482), .A2(n37667), .ZN(n35889) );
  INV_X1 U3691 ( .A(n37804), .ZN(n37806) );
  INV_X1 U3692 ( .A(n36225), .ZN(n690) );
  AND2_X1 U3693 ( .A1(n1970), .A2(n2176), .ZN(n39483) );
  INV_X1 U3694 ( .A(n36616), .ZN(n34648) );
  CLKBUF_X1 U3696 ( .A(n35531), .Z(n37438) );
  INV_X1 U3697 ( .A(n38201), .ZN(n1764) );
  OR2_X1 U3698 ( .A1(n7729), .A2(n38659), .ZN(n38666) );
  NAND2_X1 U3699 ( .A1(n38035), .A2(n38040), .ZN(n36383) );
  INV_X1 U3703 ( .A(n37747), .ZN(n691) );
  BUF_X1 U3705 ( .A(n33456), .Z(n36189) );
  OR2_X1 U3706 ( .A1(n36232), .A2(n37591), .ZN(n1006) );
  BUF_X1 U3709 ( .A(n35828), .Z(n38732) );
  INV_X1 U3713 ( .A(n37665), .ZN(n6614) );
  AND2_X1 U3714 ( .A1(n37596), .A2(n37371), .ZN(n37590) );
  BUF_X1 U3716 ( .A(n36771), .Z(n39014) );
  XNOR2_X1 U3718 ( .A(n1620), .B(n1619), .ZN(n38635) );
  INV_X1 U3719 ( .A(n37501), .ZN(n692) );
  INV_X1 U3721 ( .A(n37448), .ZN(n693) );
  AND2_X1 U3722 ( .A1(n31358), .A2(n51738), .ZN(n38545) );
  INV_X1 U3723 ( .A(n38084), .ZN(n38094) );
  OR2_X1 U3724 ( .A1(n34958), .A2(n36632), .ZN(n1360) );
  INV_X1 U3726 ( .A(n38040), .ZN(n35155) );
  XNOR2_X1 U3727 ( .A(n35249), .B(n36955), .ZN(n1619) );
  CLKBUF_X1 U3728 ( .A(n33174), .Z(n38037) );
  XNOR2_X1 U3729 ( .A(n8336), .B(n33538), .ZN(n38496) );
  INV_X1 U3730 ( .A(n37378), .ZN(n694) );
  XNOR2_X1 U3733 ( .A(n34772), .B(n34771), .ZN(n39028) );
  AND2_X1 U3734 ( .A1(n37399), .A2(n37406), .ZN(n37551) );
  INV_X1 U3735 ( .A(n36458), .ZN(n36590) );
  XNOR2_X1 U3738 ( .A(n34582), .B(n34583), .ZN(n37633) );
  INV_X1 U3740 ( .A(n34187), .ZN(n695) );
  XNOR2_X1 U3743 ( .A(n7337), .B(n32938), .ZN(n38575) );
  INV_X1 U3744 ( .A(n51474), .ZN(n1698) );
  CLKBUF_X1 U3745 ( .A(n33995), .Z(n36518) );
  INV_X1 U3746 ( .A(n34908), .ZN(n37885) );
  AND2_X1 U3747 ( .A1(n34971), .A2(n36364), .ZN(n38001) );
  BUF_X1 U3748 ( .A(n33780), .Z(n36232) );
  AND2_X1 U3749 ( .A1(n36248), .A2(n37759), .ZN(n33370) );
  INV_X1 U3752 ( .A(n36772), .ZN(n8429) );
  INV_X1 U3753 ( .A(n34189), .ZN(n5530) );
  XNOR2_X1 U3754 ( .A(n34607), .B(n34427), .ZN(n5448) );
  INV_X1 U3756 ( .A(n35215), .ZN(n696) );
  XNOR2_X1 U3759 ( .A(n35247), .B(n35248), .ZN(n36955) );
  XNOR2_X1 U3761 ( .A(n36769), .B(n1887), .ZN(n36772) );
  XNOR2_X1 U3762 ( .A(n34308), .B(n34307), .ZN(n34656) );
  INV_X1 U3763 ( .A(n36429), .ZN(n698) );
  XNOR2_X1 U3764 ( .A(n33251), .B(n35402), .ZN(n36312) );
  INV_X1 U3765 ( .A(n37969), .ZN(n699) );
  XNOR2_X1 U3767 ( .A(n35280), .B(n32855), .ZN(n38561) );
  XNOR2_X1 U3768 ( .A(n7190), .B(n33582), .ZN(n37406) );
  INV_X1 U3769 ( .A(n38464), .ZN(n38471) );
  BUF_X1 U3770 ( .A(n33778), .Z(n37593) );
  XNOR2_X1 U3771 ( .A(n31018), .B(n7447), .ZN(n36299) );
  XNOR2_X1 U3772 ( .A(n6707), .B(n6706), .ZN(n36105) );
  XNOR2_X1 U3774 ( .A(n35492), .B(n35491), .ZN(n37439) );
  XNOR2_X1 U3775 ( .A(n3365), .B(n34112), .ZN(n36015) );
  XNOR2_X1 U3776 ( .A(n34229), .B(n1489), .ZN(n34231) );
  XNOR2_X1 U3778 ( .A(n35259), .B(n35260), .ZN(n1620) );
  XNOR2_X1 U3779 ( .A(n36874), .B(n328), .ZN(n32655) );
  XNOR2_X1 U3781 ( .A(n35404), .B(n33540), .ZN(n35280) );
  INV_X1 U3783 ( .A(n33540), .ZN(n35680) );
  XNOR2_X1 U3785 ( .A(n36934), .B(n1490), .ZN(n1489) );
  INV_X1 U3786 ( .A(n35247), .ZN(n36856) );
  INV_X1 U3787 ( .A(n35748), .ZN(n34608) );
  XNOR2_X1 U3788 ( .A(n868), .B(n34156), .ZN(n33542) );
  AND3_X1 U3789 ( .A1(n6000), .A2(n7907), .A3(n31293), .ZN(n35749) );
  INV_X1 U3790 ( .A(n51472), .ZN(n1490) );
  INV_X1 U3794 ( .A(n35391), .ZN(n701) );
  XNOR2_X1 U3795 ( .A(n35047), .B(n4990), .ZN(n6603) );
  XNOR2_X1 U3796 ( .A(n37326), .B(n908), .ZN(n37327) );
  XNOR2_X1 U3797 ( .A(n34594), .B(n35075), .ZN(n33212) );
  NAND2_X1 U3800 ( .A1(n2289), .A2(n6195), .ZN(n35086) );
  INV_X1 U3802 ( .A(n36880), .ZN(n908) );
  XNOR2_X1 U3803 ( .A(n33911), .B(n37241), .ZN(n35047) );
  XNOR2_X1 U3804 ( .A(n33541), .B(n34369), .ZN(n868) );
  XNOR2_X1 U3806 ( .A(n51446), .B(n36671), .ZN(n37063) );
  INV_X1 U3807 ( .A(n35075), .ZN(n34104) );
  NAND3_X1 U3811 ( .A1(n3046), .A2(n31837), .A3(n3045), .ZN(n34620) );
  INV_X1 U3813 ( .A(n31525), .ZN(n1021) );
  AND2_X1 U3815 ( .A1(n32412), .A2(n32406), .ZN(n8250) );
  NOR2_X1 U3818 ( .A1(n31524), .A2(n31525), .ZN(n33326) );
  AND4_X1 U3819 ( .A1(n7908), .A2(n31292), .A3(n31287), .A4(n31288), .ZN(n6000) );
  XNOR2_X1 U3823 ( .A(n33806), .B(n842), .ZN(n34296) );
  NAND2_X1 U3826 ( .A1(n30992), .A2(n31500), .ZN(n8484) );
  XNOR2_X1 U3827 ( .A(n34604), .B(n34603), .ZN(n1117) );
  AND2_X1 U3828 ( .A1(n1292), .A2(n1290), .ZN(n32061) );
  BUF_X2 U3830 ( .A(n33335), .Z(n704) );
  AND3_X1 U3831 ( .A1(n28494), .A2(n28493), .A3(n28492), .ZN(n829) );
  AND3_X1 U3832 ( .A1(n29394), .A2(n5122), .A3(n6135), .ZN(n4785) );
  NAND4_X2 U3833 ( .A1(n31330), .A2(n31329), .A3(n31328), .A4(n31327), .ZN(
        n36829) );
  NAND4_X1 U3834 ( .A1(n25985), .A2(n25986), .A3(n25987), .A4(n25984), .ZN(
        n33566) );
  NAND4_X2 U3835 ( .A1(n29358), .A2(n29361), .A3(n29360), .A4(n29359), .ZN(
        n34382) );
  AND3_X1 U3838 ( .A1(n30656), .A2(n30655), .A3(n925), .ZN(n923) );
  NAND3_X1 U3840 ( .A1(n32322), .A2(n5599), .A3(n32323), .ZN(n5598) );
  NAND4_X1 U3841 ( .A1(n32651), .A2(n32650), .A3(n32653), .A4(n32652), .ZN(
        n34360) );
  AND4_X1 U3843 ( .A1(n29845), .A2(n4848), .A3(n31276), .A4(n29844), .ZN(
        n29846) );
  AND2_X1 U3844 ( .A1(n33162), .A2(n33152), .ZN(n1396) );
  NOR2_X1 U3845 ( .A1(n1870), .A2(n27152), .ZN(n27157) );
  AOI22_X1 U3846 ( .A1(n32445), .A2(n31958), .B1(n31956), .B2(n31957), .ZN(
        n1566) );
  NAND3_X1 U3847 ( .A1(n1247), .A2(n30938), .A3(n30937), .ZN(n32337) );
  AOI21_X1 U3848 ( .B1(n31254), .B2(n31253), .A(n895), .ZN(n31255) );
  AND2_X1 U3849 ( .A1(n2011), .A2(n3846), .ZN(n31168) );
  OAI21_X1 U3850 ( .B1(n1485), .B2(n31675), .A(n2094), .ZN(n29099) );
  AND2_X1 U3851 ( .A1(n26637), .A2(n6561), .ZN(n6560) );
  AND4_X1 U3852 ( .A1(n29090), .A2(n3136), .A3(n29091), .A4(n32134), .ZN(n3139) );
  AOI21_X1 U3853 ( .B1(n32127), .B2(n32126), .A(n1684), .ZN(n32140) );
  INV_X1 U3854 ( .A(n31450), .ZN(n31440) );
  AND3_X1 U3855 ( .A1(n29107), .A2(n29108), .A3(n29106), .ZN(n1699) );
  INV_X1 U3857 ( .A(n32588), .ZN(n1181) );
  NOR2_X1 U3858 ( .A1(n6421), .A2(n6420), .ZN(n6419) );
  NOR2_X1 U3859 ( .A1(n32396), .A2(n1428), .ZN(n1426) );
  AND4_X1 U3860 ( .A1(n31419), .A2(n52111), .A3(n31146), .A4(n31892), .ZN(
        n1343) );
  AND3_X1 U3861 ( .A1(n31065), .A2(n30926), .A3(n30927), .ZN(n1247) );
  OAI21_X1 U3862 ( .B1(n3240), .B2(n31626), .A(n31580), .ZN(n28727) );
  OR2_X1 U3863 ( .A1(n30516), .A2(n28607), .ZN(n30518) );
  AND2_X1 U3864 ( .A1(n6107), .A2(n30576), .ZN(n31819) );
  OAI21_X1 U3866 ( .B1(n31989), .B2(n31990), .A(n32004), .ZN(n1770) );
  NOR2_X1 U3867 ( .A1(n32124), .A2(n32130), .ZN(n872) );
  AND2_X1 U3868 ( .A1(n31815), .A2(n6107), .ZN(n3612) );
  INV_X1 U3869 ( .A(n31391), .ZN(n895) );
  INV_X1 U3872 ( .A(n30143), .ZN(n1988) );
  NOR2_X1 U3874 ( .A1(n31586), .A2(n31639), .ZN(n3240) );
  INV_X1 U3875 ( .A(n30976), .ZN(n1610) );
  INV_X1 U3876 ( .A(n30981), .ZN(n31693) );
  INV_X1 U3877 ( .A(n31265), .ZN(n30103) );
  NOR2_X1 U3879 ( .A1(n32595), .A2(n32590), .ZN(n32587) );
  OR2_X1 U3880 ( .A1(n32225), .A2(n1038), .ZN(n32227) );
  AND2_X1 U3881 ( .A1(n30647), .A2(n31302), .ZN(n920) );
  AND2_X1 U3882 ( .A1(n31454), .A2(n31538), .ZN(n31172) );
  NOR2_X1 U3883 ( .A1(n29618), .A2(n32590), .ZN(n1458) );
  AND2_X1 U3884 ( .A1(n32251), .A2(n31777), .ZN(n1072) );
  INV_X1 U3885 ( .A(n31394), .ZN(n32831) );
  INV_X1 U3886 ( .A(n31301), .ZN(n30647) );
  NAND2_X1 U3887 ( .A1(n3373), .A2(n8750), .ZN(n32815) );
  OR2_X1 U3888 ( .A1(n31876), .A2(n51743), .ZN(n31885) );
  INV_X1 U3891 ( .A(n31269), .ZN(n30110) );
  INV_X1 U3892 ( .A(n32420), .ZN(n32816) );
  AND2_X1 U3893 ( .A1(n32788), .A2(n32157), .ZN(n1115) );
  INV_X1 U3895 ( .A(n32566), .ZN(n854) );
  AND2_X1 U3896 ( .A1(n32251), .A2(n32243), .ZN(n29363) );
  NOR2_X1 U3897 ( .A1(n31683), .A2(n31684), .ZN(n30004) );
  OR2_X2 U3898 ( .A1(n1880), .A2(n30779), .ZN(n31546) );
  INV_X1 U3900 ( .A(n33036), .ZN(n705) );
  OR2_X1 U3901 ( .A1(n32507), .A2(n31986), .ZN(n31987) );
  AND2_X1 U3902 ( .A1(n32420), .A2(n31401), .ZN(n31391) );
  OR2_X1 U3903 ( .A1(n31986), .A2(n31995), .ZN(n30872) );
  AND2_X1 U3904 ( .A1(n31725), .A2(n5995), .ZN(n32151) );
  NOR2_X1 U3905 ( .A1(n30058), .A2(n31114), .ZN(n30943) );
  OR2_X1 U3908 ( .A1(n31567), .A2(n31558), .ZN(n31569) );
  OR2_X1 U3909 ( .A1(n7430), .A2(n32407), .ZN(n33159) );
  AND2_X1 U3910 ( .A1(n29622), .A2(n32595), .ZN(n1194) );
  NOR2_X1 U3911 ( .A1(n3224), .A2(n30102), .ZN(n30106) );
  NOR2_X1 U3912 ( .A1(n31510), .A2(n31513), .ZN(n1767) );
  OR2_X1 U3914 ( .A1(n50981), .A2(n32194), .ZN(n32216) );
  OR2_X1 U3916 ( .A1(n29998), .A2(n31679), .ZN(n30976) );
  OR2_X1 U3917 ( .A1(n31055), .A2(n30931), .ZN(n31511) );
  OR2_X1 U3918 ( .A1(n29837), .A2(n31496), .ZN(n30098) );
  AND2_X1 U3919 ( .A1(n31725), .A2(n32787), .ZN(n32778) );
  INV_X1 U3920 ( .A(n31989), .ZN(n707) );
  INV_X1 U3922 ( .A(n1385), .ZN(n32440) );
  OR2_X1 U3923 ( .A1(n31904), .A2(n31398), .ZN(n1269) );
  AND2_X1 U3924 ( .A1(n1037), .A2(n32252), .ZN(n32225) );
  OR2_X1 U3926 ( .A1(n32386), .A2(n31910), .ZN(n1140) );
  AOI22_X1 U3928 ( .A1(n26827), .A2(n26960), .B1(n26826), .B2(n27582), .ZN(
        n26849) );
  INV_X1 U3929 ( .A(n32491), .ZN(n709) );
  NOR2_X1 U3930 ( .A1(n31496), .A2(n31484), .ZN(n31269) );
  INV_X1 U3931 ( .A(n31781), .ZN(n710) );
  NAND4_X2 U3932 ( .A1(n3047), .A2(n28553), .A3(n28564), .A4(n2634), .ZN(
        n32684) );
  INV_X1 U3933 ( .A(n32254), .ZN(n1037) );
  AND2_X1 U3934 ( .A1(n32724), .A2(n32725), .ZN(n1168) );
  BUF_X1 U3935 ( .A(n27023), .Z(n31338) );
  INV_X1 U3936 ( .A(n30854), .ZN(n1672) );
  NOR2_X1 U3937 ( .A1(n31401), .A2(n900), .ZN(n32819) );
  AND2_X1 U3938 ( .A1(n32915), .A2(n32633), .ZN(n879) );
  AND2_X1 U3939 ( .A1(n32793), .A2(n32785), .ZN(n31726) );
  BUF_X1 U3940 ( .A(n28597), .Z(n31668) );
  BUF_X2 U3941 ( .A(n31753), .Z(n711) );
  OR2_X1 U3942 ( .A1(n1085), .A2(n32719), .ZN(n1479) );
  AND2_X1 U3943 ( .A1(n31384), .A2(n30534), .ZN(n8517) );
  OR2_X1 U3945 ( .A1(n6969), .A2(n32210), .ZN(n32197) );
  AND2_X1 U3947 ( .A1(n1038), .A2(n32252), .ZN(n32255) );
  NAND2_X2 U3948 ( .A1(n27825), .A2(n838), .ZN(n31425) );
  INV_X1 U3951 ( .A(n32386), .ZN(n713) );
  INV_X1 U3953 ( .A(n32128), .ZN(n715) );
  AND2_X1 U3954 ( .A1(n32089), .A2(n32558), .ZN(n31610) );
  AND2_X1 U3955 ( .A1(n1855), .A2(n1853), .ZN(n31286) );
  INV_X1 U3958 ( .A(n32210), .ZN(n5109) );
  AND2_X1 U3959 ( .A1(n31512), .A2(n30924), .ZN(n31510) );
  INV_X1 U3960 ( .A(n31899), .ZN(n717) );
  AND3_X1 U3962 ( .A1(n7313), .A2(n24677), .A3(n8598), .ZN(n6113) );
  AND3_X1 U3964 ( .A1(n5028), .A2(n5027), .A3(n30748), .ZN(n1086) );
  AND3_X1 U3966 ( .A1(n4117), .A2(n4360), .A3(n4359), .ZN(n27867) );
  AND2_X1 U3969 ( .A1(n8601), .A2(n24676), .ZN(n7312) );
  INV_X1 U3970 ( .A(n30534), .ZN(n720) );
  AND2_X1 U3971 ( .A1(n26790), .A2(n26791), .ZN(n29096) );
  INV_X1 U3972 ( .A(n31870), .ZN(n31800) );
  INV_X1 U3973 ( .A(n32251), .ZN(n1038) );
  NAND4_X1 U3975 ( .A1(n1323), .A2(n1322), .A3(n26932), .A4(n26931), .ZN(
        n31113) );
  INV_X1 U3978 ( .A(n6969), .ZN(n32212) );
  NAND2_X1 U3980 ( .A1(n5420), .A2(n7382), .ZN(n31850) );
  NAND2_X2 U3981 ( .A1(n1855), .A2(n29209), .ZN(n32402) );
  NOR2_X1 U3982 ( .A1(n32066), .A2(n1854), .ZN(n1853) );
  INV_X1 U3983 ( .A(n29209), .ZN(n1854) );
  INV_X1 U3984 ( .A(n31712), .ZN(n721) );
  AND3_X1 U3985 ( .A1(n5567), .A2(n27740), .A3(n27741), .ZN(n4113) );
  INV_X1 U3986 ( .A(n27725), .ZN(n5568) );
  INV_X1 U3987 ( .A(n31484), .ZN(n722) );
  AND2_X1 U3989 ( .A1(n1852), .A2(n1851), .ZN(n1855) );
  INV_X1 U3990 ( .A(n31306), .ZN(n724) );
  AND2_X1 U3991 ( .A1(n27544), .A2(n27543), .ZN(n1804) );
  AND3_X1 U3992 ( .A1(n6056), .A2(n26346), .A3(n26344), .ZN(n1154) );
  AND2_X1 U3994 ( .A1(n30468), .A2(n30466), .ZN(n901) );
  OAI211_X1 U3995 ( .C1(n24355), .C2(n30764), .A(n1674), .B(n8377), .ZN(n1679)
         );
  AND2_X1 U3996 ( .A1(n24353), .A2(n1678), .ZN(n1677) );
  AND2_X1 U3998 ( .A1(n8273), .A2(n8274), .ZN(n1163) );
  AND2_X1 U4000 ( .A1(n28961), .A2(n29796), .ZN(n28967) );
  AND4_X1 U4001 ( .A1(n30454), .A2(n30447), .A3(n28445), .A4(n28444), .ZN(
        n28454) );
  AND4_X1 U4002 ( .A1(n27405), .A2(n27404), .A3(n30743), .A4(n27403), .ZN(
        n27406) );
  AND2_X1 U4003 ( .A1(n7816), .A2(n29349), .ZN(n1050) );
  NAND4_X2 U4004 ( .A1(n6014), .A2(n6015), .A3(n27705), .A4(n6017), .ZN(n29686) );
  AND3_X1 U4006 ( .A1(n28554), .A2(n30301), .A3(n28552), .ZN(n3047) );
  NAND2_X1 U4007 ( .A1(n27399), .A2(n30376), .ZN(n1123) );
  OAI21_X1 U4009 ( .B1(n29690), .B2(n29692), .A(n1982), .ZN(n28746) );
  NAND4_X2 U4010 ( .A1(n3465), .A2(n3464), .A3(n27102), .A4(n27101), .ZN(
        n32503) );
  AND4_X1 U4011 ( .A1(n27138), .A2(n27137), .A3(n27136), .A4(n27135), .ZN(
        n27142) );
  AND3_X1 U4013 ( .A1(n29919), .A2(n27556), .A3(n26925), .ZN(n1323) );
  OR2_X1 U4015 ( .A1(n27828), .A2(n29450), .ZN(n5545) );
  OR2_X1 U4018 ( .A1(n24355), .A2(n30763), .ZN(n1674) );
  AND2_X1 U4019 ( .A1(n26928), .A2(n30766), .ZN(n1081) );
  OR2_X1 U4020 ( .A1(n30752), .A2(n30757), .ZN(n29919) );
  NOR2_X1 U4021 ( .A1(n28458), .A2(n28496), .ZN(n1166) );
  AOI21_X1 U4022 ( .B1(n6403), .B2(n30427), .A(n1983), .ZN(n28337) );
  AOI22_X1 U4023 ( .A1(n30756), .A2(n29926), .B1(n29927), .B2(n30766), .ZN(
        n29928) );
  AND2_X1 U4024 ( .A1(n27834), .A2(n27835), .ZN(n29437) );
  AND2_X1 U4025 ( .A1(n29208), .A2(n29207), .ZN(n1852) );
  OAI21_X1 U4026 ( .B1(n4405), .B2(n29352), .A(n29206), .ZN(n1851) );
  AND4_X1 U4027 ( .A1(n8435), .A2(n3740), .A3(n25733), .A4(n26659), .ZN(n843)
         );
  AND2_X1 U4028 ( .A1(n26874), .A2(n26873), .ZN(n1564) );
  AND2_X1 U4029 ( .A1(n1638), .A2(n27561), .ZN(n27562) );
  AND3_X1 U4030 ( .A1(n30385), .A2(n30386), .A3(n1905), .ZN(n30388) );
  AND2_X1 U4031 ( .A1(n28782), .A2(n28781), .ZN(n28817) );
  AOI21_X1 U4035 ( .B1(n26829), .B2(n1374), .A(n1372), .ZN(n27415) );
  AND2_X1 U4036 ( .A1(n27168), .A2(n27169), .ZN(n1803) );
  OR2_X1 U4037 ( .A1(n29139), .A2(n1771), .ZN(n26472) );
  AND2_X1 U4038 ( .A1(n1153), .A2(n5369), .ZN(n4759) );
  AND4_X1 U4039 ( .A1(n24567), .A2(n29463), .A3(n24566), .A4(n24565), .ZN(
        n8648) );
  INV_X1 U4040 ( .A(n31401), .ZN(n726) );
  AND2_X1 U4041 ( .A1(n27109), .A2(n29043), .ZN(n3464) );
  AND2_X1 U4042 ( .A1(n5564), .A2(n29220), .ZN(n1694) );
  AND2_X1 U4044 ( .A1(n30436), .A2(n1983), .ZN(n1982) );
  OAI21_X1 U4045 ( .B1(n27795), .B2(n28626), .A(n29513), .ZN(n1574) );
  NAND4_X1 U4046 ( .A1(n30177), .A2(n30159), .A3(n30178), .A4(n30181), .ZN(
        n29139) );
  OR2_X1 U4047 ( .A1(n6048), .A2(n26842), .ZN(n30764) );
  OR2_X1 U4049 ( .A1(n29439), .A2(n906), .ZN(n907) );
  AND2_X1 U4050 ( .A1(n30235), .A2(n30234), .ZN(n857) );
  INV_X1 U4051 ( .A(n26840), .ZN(n1471) );
  NOR2_X1 U4052 ( .A1(n6048), .A2(n1676), .ZN(n1675) );
  AND2_X1 U4053 ( .A1(n1839), .A2(n30771), .ZN(n26929) );
  NOR2_X1 U4054 ( .A1(n28907), .A2(n28577), .ZN(n27998) );
  OR2_X1 U4055 ( .A1(n28194), .A2(n29008), .ZN(n28937) );
  NOR2_X1 U4057 ( .A1(n29915), .A2(n29916), .ZN(n1939) );
  INV_X1 U4058 ( .A(n26956), .ZN(n1482) );
  INV_X1 U4059 ( .A(n26879), .ZN(n1563) );
  OR2_X1 U4060 ( .A1(n30688), .A2(n30692), .ZN(n29936) );
  NOR2_X1 U4061 ( .A1(n30434), .A2(n1983), .ZN(n29706) );
  AOI21_X1 U4062 ( .B1(n30783), .B2(n1373), .A(n29901), .ZN(n1372) );
  INV_X1 U4063 ( .A(n24569), .ZN(n27641) );
  AND2_X1 U4064 ( .A1(n26775), .A2(n27686), .ZN(n824) );
  INV_X1 U4065 ( .A(n26842), .ZN(n30755) );
  INV_X1 U4066 ( .A(n51746), .ZN(n1981) );
  AND2_X1 U4067 ( .A1(n28918), .A2(n29013), .ZN(n29018) );
  INV_X1 U4068 ( .A(n27828), .ZN(n1030) );
  INV_X1 U4069 ( .A(n30451), .ZN(n727) );
  AND2_X1 U4070 ( .A1(n6449), .A2(n27690), .ZN(n27686) );
  BUF_X1 U4071 ( .A(n27709), .Z(n2115) );
  NAND2_X1 U4072 ( .A1(n402), .A2(n30393), .ZN(n30389) );
  AND2_X1 U4073 ( .A1(n29202), .A2(n51109), .ZN(n1156) );
  OR2_X1 U4074 ( .A1(n29774), .A2(n29784), .ZN(n28766) );
  OR2_X1 U4075 ( .A1(n7805), .A2(n24687), .ZN(n2799) );
  NOR2_X1 U4076 ( .A1(n1983), .A2(n51746), .ZN(n29697) );
  OR2_X1 U4077 ( .A1(n30210), .A2(n29200), .ZN(n29350) );
  AND2_X1 U4078 ( .A1(n30211), .A2(n30210), .ZN(n27885) );
  INV_X1 U4079 ( .A(n29549), .ZN(n29541) );
  NOR2_X1 U4080 ( .A1(n27890), .A2(n29314), .ZN(n27805) );
  AND2_X1 U4084 ( .A1(n30768), .A2(n30769), .ZN(n30766) );
  INV_X1 U4086 ( .A(n30430), .ZN(n728) );
  INV_X1 U4087 ( .A(n30757), .ZN(n1839) );
  AND2_X1 U4088 ( .A1(n6059), .A2(n29526), .ZN(n26974) );
  AND2_X1 U4089 ( .A1(n27837), .A2(n27835), .ZN(n1547) );
  OR2_X1 U4091 ( .A1(n51746), .A2(n30426), .ZN(n30429) );
  AND2_X1 U4092 ( .A1(n30758), .A2(n29921), .ZN(n24355) );
  NAND2_X1 U4094 ( .A1(n28189), .A2(n28796), .ZN(n28982) );
  OR2_X1 U4095 ( .A1(n26722), .A2(n6602), .ZN(n27033) );
  INV_X1 U4096 ( .A(n30452), .ZN(n1927) );
  INV_X1 U4097 ( .A(n29552), .ZN(n26764) );
  AND2_X1 U4099 ( .A1(n24776), .A2(n982), .ZN(n981) );
  INV_X1 U4100 ( .A(n26977), .ZN(n29509) );
  INV_X1 U4101 ( .A(n29518), .ZN(n729) );
  NAND2_X1 U4102 ( .A1(n26039), .A2(n1023), .ZN(n6602) );
  INV_X1 U4103 ( .A(n30768), .ZN(n730) );
  INV_X1 U4104 ( .A(n1023), .ZN(n29438) );
  OR2_X1 U4105 ( .A1(n28971), .A2(n27278), .ZN(n29715) );
  INV_X1 U4107 ( .A(n7614), .ZN(n30280) );
  INV_X1 U4108 ( .A(n27158), .ZN(n28810) );
  NOR2_X1 U4111 ( .A1(n27654), .A2(n3765), .ZN(n1048) );
  BUF_X1 U4114 ( .A(n24563), .Z(n29471) );
  INV_X1 U4115 ( .A(n30724), .ZN(n731) );
  AND2_X1 U4116 ( .A1(n30771), .A2(n24354), .ZN(n30763) );
  INV_X1 U4117 ( .A(n27558), .ZN(n30758) );
  NAND2_X1 U4118 ( .A1(n1680), .A2(n29550), .ZN(n26761) );
  NAND2_X1 U4122 ( .A1(n30218), .A2(n30233), .ZN(n29248) );
  OR2_X1 U4124 ( .A1(n28659), .A2(n30233), .ZN(n30226) );
  OR2_X1 U4125 ( .A1(n29546), .A2(n29545), .ZN(n1285) );
  INV_X1 U4126 ( .A(n28738), .ZN(n29867) );
  OR2_X1 U4127 ( .A1(n5211), .A2(n30431), .ZN(n29868) );
  OR2_X1 U4129 ( .A1(n29346), .A2(n967), .ZN(n30211) );
  AND2_X1 U4132 ( .A1(n29692), .A2(n5330), .ZN(n813) );
  INV_X1 U4133 ( .A(n487), .ZN(n1983) );
  AND2_X1 U4134 ( .A1(n24354), .A2(n30769), .ZN(n29921) );
  INV_X1 U4135 ( .A(n51111), .ZN(n6339) );
  AND2_X1 U4136 ( .A1(n29439), .A2(n2213), .ZN(n1805) );
  OR2_X1 U4137 ( .A1(n30312), .A2(n30182), .ZN(n6342) );
  INV_X1 U4138 ( .A(n29901), .ZN(n29892) );
  AND2_X1 U4139 ( .A1(n29513), .A2(n29507), .ZN(n29522) );
  OR2_X1 U4140 ( .A1(n28708), .A2(n5656), .ZN(n29185) );
  NOR2_X1 U4141 ( .A1(n7052), .A2(n29190), .ZN(n29281) );
  INV_X1 U4143 ( .A(n29320), .ZN(n1817) );
  INV_X1 U4144 ( .A(n29461), .ZN(n732) );
  INV_X1 U4145 ( .A(n28615), .ZN(n27796) );
  INV_X1 U4146 ( .A(n30387), .ZN(n1906) );
  INV_X1 U4147 ( .A(n29346), .ZN(n733) );
  INV_X1 U4148 ( .A(n27093), .ZN(n967) );
  INV_X1 U4149 ( .A(n30694), .ZN(n734) );
  OR2_X1 U4150 ( .A1(n30245), .A2(n51726), .ZN(n2889) );
  INV_X1 U4151 ( .A(n29347), .ZN(n735) );
  AND2_X1 U4153 ( .A1(n27040), .A2(n26039), .ZN(n1015) );
  XNOR2_X1 U4155 ( .A(n27372), .B(n1658), .ZN(n30374) );
  INV_X1 U4157 ( .A(n27669), .ZN(n736) );
  INV_X1 U4159 ( .A(n25734), .ZN(n29309) );
  BUF_X1 U4160 ( .A(n26619), .Z(n29033) );
  INV_X1 U4161 ( .A(n30718), .ZN(n27164) );
  BUF_X1 U4163 ( .A(n25297), .Z(n28588) );
  NOR2_X1 U4164 ( .A1(n28623), .A2(n29507), .ZN(n28616) );
  BUF_X1 U4165 ( .A(n26288), .Z(n28626) );
  XNOR2_X1 U4166 ( .A(n24954), .B(n24955), .ZN(n30244) );
  XNOR2_X1 U4167 ( .A(n25835), .B(n25834), .ZN(n29488) );
  OR2_X1 U4169 ( .A1(n51116), .A2(n25479), .ZN(n28711) );
  XNOR2_X1 U4170 ( .A(n4491), .B(n8280), .ZN(n24878) );
  XNOR2_X1 U4171 ( .A(n27432), .B(n27431), .ZN(n28738) );
  INV_X1 U4173 ( .A(n30771), .ZN(n1676) );
  BUF_X1 U4175 ( .A(n25626), .Z(n29259) );
  INV_X1 U4176 ( .A(n27729), .ZN(n27623) );
  INV_X1 U4177 ( .A(n2707), .ZN(n3827) );
  INV_X1 U4178 ( .A(n27618), .ZN(n737) );
  AND2_X1 U4179 ( .A1(n30345), .A2(n7721), .ZN(n30340) );
  OR2_X1 U4182 ( .A1(n27070), .A2(n27652), .ZN(n982) );
  INV_X1 U4183 ( .A(n29550), .ZN(n27049) );
  OR2_X1 U4184 ( .A1(n25626), .A2(n25603), .ZN(n30232) );
  AND2_X1 U4185 ( .A1(n26944), .A2(n26937), .ZN(n1565) );
  OR2_X1 U4187 ( .A1(n30265), .A2(n6486), .ZN(n29221) );
  OR2_X1 U4188 ( .A1(n7721), .A2(n30345), .ZN(n28849) );
  NAND2_X1 U4189 ( .A1(n8640), .A2(n51723), .ZN(n29901) );
  INV_X1 U4190 ( .A(n2677), .ZN(n24774) );
  OR2_X1 U4192 ( .A1(n1484), .A2(n26954), .ZN(n27677) );
  XNOR2_X1 U4196 ( .A(n3232), .B(n27444), .ZN(n6403) );
  INV_X1 U4198 ( .A(n30780), .ZN(n30795) );
  XNOR2_X1 U4199 ( .A(n24746), .B(n24745), .ZN(n26937) );
  INV_X1 U4200 ( .A(n29923), .ZN(n738) );
  XNOR2_X1 U4202 ( .A(n26400), .B(n27183), .ZN(n28919) );
  INV_X1 U4203 ( .A(n30179), .ZN(n739) );
  INV_X1 U4205 ( .A(n30191), .ZN(n740) );
  INV_X1 U4207 ( .A(n29782), .ZN(n742) );
  INV_X1 U4209 ( .A(n27695), .ZN(n743) );
  XNOR2_X1 U4210 ( .A(n25194), .B(n25193), .ZN(n25198) );
  INV_X1 U4211 ( .A(n29507), .ZN(n29535) );
  XNOR2_X1 U4212 ( .A(n24983), .B(n7551), .ZN(n6730) );
  XNOR2_X1 U4213 ( .A(n26128), .B(n2316), .ZN(n26197) );
  INV_X1 U4217 ( .A(n7721), .ZN(n745) );
  XNOR2_X1 U4218 ( .A(n25895), .B(n25894), .ZN(n5228) );
  XNOR2_X1 U4219 ( .A(n1514), .B(n1515), .ZN(n1513) );
  INV_X1 U4220 ( .A(n27918), .ZN(n746) );
  INV_X1 U4221 ( .A(n29442), .ZN(n747) );
  XNOR2_X1 U4223 ( .A(n4239), .B(n21002), .ZN(n27633) );
  XNOR2_X1 U4224 ( .A(n8464), .B(n24691), .ZN(n25803) );
  XNOR2_X1 U4226 ( .A(n5518), .B(n21764), .ZN(n23939) );
  INV_X1 U4227 ( .A(n28068), .ZN(n1270) );
  XNOR2_X1 U4228 ( .A(n28295), .B(n5313), .ZN(n1515) );
  XNOR2_X1 U4229 ( .A(n24915), .B(n28248), .ZN(n1498) );
  XNOR2_X1 U4230 ( .A(n27264), .B(n27263), .ZN(n28367) );
  BUF_X1 U4231 ( .A(n27480), .Z(n27330) );
  INV_X1 U4233 ( .A(n28296), .ZN(n1514) );
  BUF_X1 U4234 ( .A(n26536), .Z(n2212) );
  XNOR2_X1 U4235 ( .A(n26274), .B(n7319), .ZN(n25935) );
  XNOR2_X1 U4236 ( .A(n27419), .B(n1027), .ZN(n27421) );
  INV_X1 U4237 ( .A(n25682), .ZN(n27196) );
  XNOR2_X1 U4239 ( .A(n51122), .B(n24793), .ZN(n23793) );
  XNOR2_X1 U4240 ( .A(n51122), .B(n24757), .ZN(n25609) );
  XNOR2_X1 U4243 ( .A(n23402), .B(n1377), .ZN(n23403) );
  XNOR2_X1 U4245 ( .A(n25047), .B(n25308), .ZN(n27234) );
  INV_X1 U4246 ( .A(n3110), .ZN(n3031) );
  AND2_X1 U4248 ( .A1(n22708), .A2(n6285), .ZN(n24455) );
  INV_X1 U4250 ( .A(n7319), .ZN(n1027) );
  XNOR2_X1 U4251 ( .A(n26093), .B(n26100), .ZN(n26046) );
  XNOR2_X1 U4252 ( .A(n25903), .B(n1377), .ZN(n22810) );
  XNOR2_X1 U4254 ( .A(n6434), .B(n24556), .ZN(n2125) );
  AND4_X2 U4256 ( .A1(n20870), .A2(n20871), .A3(n7133), .A4(n20869), .ZN(n7319) );
  XNOR2_X1 U4257 ( .A(n1377), .B(n28291), .ZN(n25896) );
  NAND4_X1 U4260 ( .A1(n21858), .A2(n21857), .A3(n21856), .A4(n21855), .ZN(
        n23772) );
  AND3_X1 U4261 ( .A1(n8213), .A2(n4230), .A3(n8216), .ZN(n3110) );
  NAND3_X1 U4264 ( .A1(n22410), .A2(n21729), .A3(n2259), .ZN(n25003) );
  XNOR2_X1 U4265 ( .A(n6434), .B(n1377), .ZN(n28119) );
  XNOR2_X1 U4267 ( .A(n27211), .B(n4564), .ZN(n28246) );
  XNOR2_X1 U4271 ( .A(n25747), .B(n24302), .ZN(n27459) );
  XNOR2_X1 U4272 ( .A(n24795), .B(n2203), .ZN(n25882) );
  XNOR2_X1 U4276 ( .A(n1377), .B(n26402), .ZN(n26409) );
  AND2_X1 U4280 ( .A1(n20537), .A2(n20533), .ZN(n1954) );
  XNOR2_X1 U4281 ( .A(n1377), .B(n27354), .ZN(n27356) );
  AND2_X1 U4282 ( .A1(n1966), .A2(n1965), .ZN(n21721) );
  NAND4_X2 U4283 ( .A1(n22280), .A2(n7831), .A3(n1412), .A4(n1413), .ZN(n28353) );
  AND3_X1 U4284 ( .A1(n22871), .A2(n22870), .A3(n22869), .ZN(n6266) );
  NAND4_X1 U4288 ( .A1(n22139), .A2(n22138), .A3(n22137), .A4(n22136), .ZN(
        n27272) );
  NAND2_X1 U4290 ( .A1(n5019), .A2(n8151), .ZN(n27211) );
  NAND3_X1 U4291 ( .A1(n3666), .A2(n3665), .A3(n17615), .ZN(n24736) );
  INV_X1 U4293 ( .A(n25946), .ZN(n1025) );
  NAND4_X1 U4295 ( .A1(n5005), .A2(n5000), .A3(n5591), .A4(n4999), .ZN(n27303)
         );
  OAI211_X1 U4296 ( .C1(n16854), .C2(n2130), .A(n16853), .B(n989), .ZN(n22762)
         );
  AND2_X1 U4299 ( .A1(n20536), .A2(n1959), .ZN(n1955) );
  AND4_X1 U4300 ( .A1(n4986), .A2(n16852), .A3(n16850), .A4(n16851), .ZN(
        n16853) );
  AND3_X1 U4301 ( .A1(n6134), .A2(n7028), .A3(n22250), .ZN(n6133) );
  AND2_X1 U4302 ( .A1(n21341), .A2(n990), .ZN(n989) );
  AND3_X1 U4303 ( .A1(n21509), .A2(n21511), .A3(n21510), .ZN(n6761) );
  INV_X1 U4304 ( .A(n20282), .ZN(n6736) );
  AND2_X1 U4305 ( .A1(n21995), .A2(n21984), .ZN(n1558) );
  AND2_X1 U4306 ( .A1(n21087), .A2(n21086), .ZN(n1996) );
  NOR2_X1 U4307 ( .A1(n21742), .A2(n17512), .ZN(n17515) );
  AND2_X1 U4309 ( .A1(n22510), .A2(n1431), .ZN(n1430) );
  NAND4_X1 U4310 ( .A1(n1493), .A2(n24251), .A3(n24252), .A4(n1492), .ZN(
        n24253) );
  NOR2_X1 U4311 ( .A1(n323), .A2(n20283), .ZN(n1993) );
  AND3_X1 U4312 ( .A1(n24342), .A2(n24340), .A3(n24341), .ZN(n3308) );
  OAI22_X1 U4313 ( .A1(n1998), .A2(n1997), .B1(n21908), .B2(n7247), .ZN(n1995)
         );
  AND3_X1 U4315 ( .A1(n22678), .A2(n22676), .A3(n22675), .ZN(n3820) );
  AND4_X1 U4316 ( .A1(n22077), .A2(n22078), .A3(n22079), .A4(n22076), .ZN(
        n22095) );
  AND4_X1 U4317 ( .A1(n20976), .A2(n23217), .A3(n20313), .A4(n20312), .ZN(
        n2096) );
  INV_X1 U4318 ( .A(n1968), .ZN(n1967) );
  INV_X1 U4319 ( .A(n24148), .ZN(n1609) );
  OAI211_X1 U4321 ( .C1(n21343), .C2(n19624), .A(n19623), .B(n19622), .ZN(
        n19626) );
  AOI22_X1 U4322 ( .A1(n22913), .A2(n22912), .B1(n22910), .B2(n22911), .ZN(
        n8000) );
  INV_X1 U4323 ( .A(n973), .ZN(n20964) );
  INV_X1 U4325 ( .A(n23754), .ZN(n23750) );
  INV_X1 U4326 ( .A(n8402), .ZN(n942) );
  OAI21_X1 U4327 ( .B1(n5539), .B2(n22255), .A(n21011), .ZN(n24016) );
  OR2_X1 U4328 ( .A1(n23253), .A2(n1777), .ZN(n1776) );
  NAND2_X1 U4329 ( .A1(n21834), .A2(n628), .ZN(n1903) );
  OR2_X1 U4330 ( .A1(n20992), .A2(n23485), .ZN(n990) );
  AND2_X1 U4331 ( .A1(n19553), .A2(n19552), .ZN(n3271) );
  OAI21_X1 U4332 ( .B1(n1411), .B2(n23232), .A(n23231), .ZN(n23233) );
  NOR2_X1 U4333 ( .A1(n23762), .A2(n23761), .ZN(n4722) );
  OR2_X1 U4334 ( .A1(n891), .A2(n1743), .ZN(n21817) );
  OAI21_X1 U4336 ( .B1(n23105), .B2(n23104), .A(n23103), .ZN(n1847) );
  OAI21_X1 U4337 ( .B1(n23964), .B2(n23965), .A(n23963), .ZN(n23966) );
  INV_X1 U4339 ( .A(n21778), .ZN(n1712) );
  OR2_X1 U4340 ( .A1(n22285), .A2(n20944), .ZN(n1958) );
  AND3_X1 U4341 ( .A1(n5802), .A2(n23396), .A3(n5801), .ZN(n5800) );
  OR2_X1 U4342 ( .A1(n5311), .A2(n22169), .ZN(n1522) );
  OAI21_X1 U4343 ( .B1(n21019), .B2(n975), .A(n974), .ZN(n973) );
  AND2_X1 U4344 ( .A1(n21886), .A2(n21887), .ZN(n2846) );
  OR2_X1 U4345 ( .A1(n22120), .A2(n22119), .ZN(n2053) );
  INV_X1 U4346 ( .A(n23456), .ZN(n1603) );
  OR2_X1 U4347 ( .A1(n23761), .A2(n24190), .ZN(n23754) );
  INV_X1 U4348 ( .A(n23351), .ZN(n23549) );
  OAI21_X1 U4350 ( .B1(n24028), .B2(n23392), .A(n24026), .ZN(n8254) );
  AND2_X1 U4351 ( .A1(n22123), .A2(n1777), .ZN(n23255) );
  OR2_X1 U4352 ( .A1(n23730), .A2(n24111), .ZN(n24097) );
  NOR2_X1 U4353 ( .A1(n22124), .A2(n8730), .ZN(n1904) );
  OR2_X1 U4354 ( .A1(n20309), .A2(n3646), .ZN(n20976) );
  OR2_X1 U4355 ( .A1(n21712), .A2(n22188), .ZN(n22183) );
  AND2_X1 U4357 ( .A1(n17074), .A2(n23547), .ZN(n904) );
  AOI21_X1 U4358 ( .B1(n22830), .B2(n22509), .A(n1145), .ZN(n22508) );
  OR2_X1 U4359 ( .A1(n23923), .A2(n23898), .ZN(n1148) );
  INV_X1 U4361 ( .A(n24242), .ZN(n1745) );
  NOR2_X1 U4362 ( .A1(n24245), .A2(n6744), .ZN(n1496) );
  AND2_X1 U4363 ( .A1(n21767), .A2(n21780), .ZN(n819) );
  INV_X1 U4364 ( .A(n23247), .ZN(n1777) );
  NOR2_X1 U4365 ( .A1(n5415), .A2(n24332), .ZN(n23705) );
  AND2_X1 U4367 ( .A1(n23569), .A2(n1648), .ZN(n7832) );
  OR2_X1 U4368 ( .A1(n23213), .A2(n413), .ZN(n18371) );
  OR2_X1 U4369 ( .A1(n23440), .A2(n23446), .ZN(n21999) );
  AND2_X1 U4370 ( .A1(n22358), .A2(n22359), .ZN(n1305) );
  XNOR2_X1 U4371 ( .A(n1657), .B(n23052), .ZN(n23055) );
  AND2_X1 U4373 ( .A1(n20005), .A2(n23392), .ZN(n24043) );
  NOR2_X1 U4374 ( .A1(n21671), .A2(n24413), .ZN(n23730) );
  AND2_X1 U4375 ( .A1(n8695), .A2(n22144), .ZN(n21018) );
  OAI21_X1 U4379 ( .B1(n24250), .B2(n24247), .A(n24239), .ZN(n1743) );
  OR2_X1 U4380 ( .A1(n24332), .A2(n23535), .ZN(n5260) );
  INV_X1 U4381 ( .A(n22491), .ZN(n22834) );
  INV_X1 U4383 ( .A(n22491), .ZN(n1145) );
  BUF_X1 U4384 ( .A(n21900), .Z(n7519) );
  AND2_X1 U4385 ( .A1(n8303), .A2(n23303), .ZN(n21864) );
  AND3_X1 U4386 ( .A1(n5625), .A2(n5624), .A3(n19115), .ZN(n2019) );
  INV_X1 U4387 ( .A(n23336), .ZN(n21145) );
  AND2_X1 U4388 ( .A1(n20876), .A2(n21820), .ZN(n24242) );
  INV_X1 U4389 ( .A(n22977), .ZN(n22557) );
  INV_X1 U4393 ( .A(n1648), .ZN(n1647) );
  INV_X1 U4395 ( .A(n23832), .ZN(n23828) );
  AND2_X1 U4397 ( .A1(n50992), .A2(n979), .ZN(n22143) );
  INV_X1 U4398 ( .A(n452), .ZN(n23407) );
  AND2_X1 U4399 ( .A1(n23020), .A2(n22856), .ZN(n1273) );
  OR2_X1 U4400 ( .A1(n23664), .A2(n24026), .ZN(n23670) );
  AND2_X1 U4401 ( .A1(n23306), .A2(n23316), .ZN(n3602) );
  NAND3_X1 U4403 ( .A1(n413), .A2(n22121), .A3(n418), .ZN(n20309) );
  INV_X1 U4404 ( .A(n21016), .ZN(n22859) );
  INV_X1 U4405 ( .A(n23554), .ZN(n752) );
  OR2_X1 U4406 ( .A1(n7303), .A2(n23513), .ZN(n24291) );
  OR2_X1 U4407 ( .A1(n25056), .A2(n25064), .ZN(n23104) );
  OR2_X1 U4409 ( .A1(n3822), .A2(n50990), .ZN(n23693) );
  INV_X1 U4411 ( .A(n22140), .ZN(n979) );
  AND2_X1 U4414 ( .A1(n23229), .A2(n22121), .ZN(n23209) );
  INV_X1 U4415 ( .A(n22875), .ZN(n23094) );
  NAND2_X1 U4416 ( .A1(n20403), .A2(n8230), .ZN(n22946) );
  AND2_X1 U4418 ( .A1(n18104), .A2(n1540), .ZN(n1539) );
  INV_X1 U4420 ( .A(n22085), .ZN(n23048) );
  NAND4_X1 U4423 ( .A1(n16832), .A2(n16829), .A3(n16830), .A4(n16831), .ZN(
        n16849) );
  INV_X1 U4425 ( .A(n23513), .ZN(n755) );
  INV_X1 U4426 ( .A(n17420), .ZN(n23590) );
  NAND4_X1 U4427 ( .A1(n6932), .A2(n6931), .A3(n1917), .A4(n1916), .ZN(n6930)
         );
  NAND2_X1 U4429 ( .A1(n20846), .A2(n5491), .ZN(n23957) );
  AND3_X1 U4430 ( .A1(n8590), .A2(n20486), .A3(n8588), .ZN(n2083) );
  AND3_X2 U4432 ( .A1(n6954), .A2(n6955), .A3(n6953), .ZN(n23489) );
  AOI21_X1 U4436 ( .B1(n19294), .B2(n21358), .A(n969), .ZN(n19299) );
  INV_X1 U4437 ( .A(n23244), .ZN(n757) );
  AND4_X1 U4438 ( .A1(n19419), .A2(n19434), .A3(n19420), .A4(n19421), .ZN(
        n5559) );
  AND2_X1 U4439 ( .A1(n5536), .A2(n5538), .ZN(n5535) );
  AND3_X1 U4440 ( .A1(n2693), .A2(n21746), .A3(n2692), .ZN(n8160) );
  INV_X1 U4441 ( .A(n24452), .ZN(n758) );
  NOR2_X1 U4444 ( .A1(n17854), .A2(n17855), .ZN(n17864) );
  OR2_X1 U4446 ( .A1(n8605), .A2(n17565), .ZN(n3640) );
  AND2_X1 U4448 ( .A1(n17042), .A2(n17041), .ZN(n1398) );
  AND3_X1 U4450 ( .A1(n20402), .A2(n20401), .A3(n20400), .ZN(n8230) );
  AND3_X1 U4452 ( .A1(n21643), .A2(n21641), .A3(n21642), .ZN(n1615) );
  AND2_X1 U4453 ( .A1(n4528), .A2(n19519), .ZN(n1916) );
  AND3_X1 U4454 ( .A1(n17461), .A2(n16393), .A3(n16394), .ZN(n5782) );
  OR2_X1 U4455 ( .A1(n18383), .A2(n16819), .ZN(n16397) );
  AND3_X1 U4457 ( .A1(n16396), .A2(n7584), .A3(n20039), .ZN(n16399) );
  MUX2_X1 U4458 ( .A(n16828), .B(n16827), .S(n17448), .Z(n16829) );
  AND4_X1 U4459 ( .A1(n16839), .A2(n16838), .A3(n16837), .A4(n16836), .ZN(
        n2130) );
  AND2_X1 U4460 ( .A1(n17555), .A2(n17562), .ZN(n980) );
  AOI22_X1 U4461 ( .A1(n20234), .A2(n20235), .B1(n8302), .B2(n20233), .ZN(
        n20236) );
  NAND4_X1 U4463 ( .A1(n5871), .A2(n5870), .A3(n5869), .A4(n18309), .ZN(n23229) );
  AND4_X1 U4464 ( .A1(n18321), .A2(n18320), .A3(n18322), .A4(n18319), .ZN(
        n18325) );
  OAI21_X1 U4466 ( .B1(n2058), .B2(n18330), .A(n18333), .ZN(n18334) );
  OR2_X1 U4467 ( .A1(n19638), .A2(n19637), .ZN(n19710) );
  NOR2_X1 U4469 ( .A1(n21479), .A2(n20446), .ZN(n20810) );
  OR2_X1 U4470 ( .A1(n17470), .A2(n2222), .ZN(n4193) );
  OAI21_X1 U4471 ( .B1(n1519), .B2(n18333), .A(n18061), .ZN(n1518) );
  AND2_X1 U4472 ( .A1(n16002), .A2(n21639), .ZN(n1451) );
  AND3_X1 U4473 ( .A1(n20845), .A2(n5492), .A3(n20844), .ZN(n5491) );
  AND3_X1 U4474 ( .A1(n8263), .A2(n8262), .A3(n20454), .ZN(n8261) );
  AND2_X1 U4475 ( .A1(n21462), .A2(n17712), .ZN(n20317) );
  AND2_X1 U4476 ( .A1(n5333), .A2(n590), .ZN(n20018) );
  AND2_X1 U4477 ( .A1(n21243), .A2(n19472), .ZN(n21257) );
  NOR2_X1 U4478 ( .A1(n19813), .A2(n21196), .ZN(n18108) );
  OR2_X1 U4479 ( .A1(n19513), .A2(n19514), .ZN(n19521) );
  OR2_X1 U4480 ( .A1(n20514), .A2(n1516), .ZN(n17622) );
  AND2_X1 U4481 ( .A1(n17427), .A2(n1714), .ZN(n1713) );
  OR2_X1 U4482 ( .A1(n17604), .A2(n17503), .ZN(n5197) );
  NOR2_X1 U4483 ( .A1(n20015), .A2(n1786), .ZN(n1785) );
  INV_X1 U4488 ( .A(n16891), .ZN(n20648) );
  AND2_X1 U4489 ( .A1(n17412), .A2(n2044), .ZN(n21237) );
  AND2_X1 U4491 ( .A1(n21592), .A2(n970), .ZN(n969) );
  INV_X1 U4492 ( .A(n18963), .ZN(n21254) );
  OR2_X1 U4493 ( .A1(n1053), .A2(n20399), .ZN(n14746) );
  NAND2_X1 U4494 ( .A1(n19114), .A2(n1406), .ZN(n1454) );
  AND2_X1 U4495 ( .A1(n21494), .A2(n20815), .ZN(n1366) );
  INV_X1 U4496 ( .A(n21479), .ZN(n759) );
  AND2_X1 U4497 ( .A1(n1856), .A2(n3971), .ZN(n1857) );
  NOR2_X1 U4498 ( .A1(n18047), .A2(n3181), .ZN(n5558) );
  INV_X1 U4500 ( .A(n1789), .ZN(n20458) );
  AND2_X1 U4501 ( .A1(n20681), .A2(n20232), .ZN(n20686) );
  INV_X1 U4502 ( .A(n18102), .ZN(n18869) );
  INV_X1 U4503 ( .A(n21474), .ZN(n21466) );
  OR4_X1 U4504 ( .A1(n17533), .A2(n5813), .A3(n17522), .A4(n2166), .ZN(n2645)
         );
  OR2_X1 U4505 ( .A1(n19687), .A2(n20220), .ZN(n1223) );
  AND2_X1 U4506 ( .A1(n21214), .A2(n21200), .ZN(n1319) );
  INV_X1 U4507 ( .A(n17311), .ZN(n2044) );
  NOR2_X1 U4509 ( .A1(n21234), .A2(n19514), .ZN(n17313) );
  INV_X1 U4510 ( .A(n20841), .ZN(n1797) );
  INV_X1 U4511 ( .A(n20497), .ZN(n21462) );
  INV_X1 U4512 ( .A(n20672), .ZN(n760) );
  AND2_X1 U4516 ( .A1(n17045), .A2(n1157), .ZN(n1671) );
  INV_X1 U4517 ( .A(n19513), .ZN(n761) );
  NOR2_X1 U4518 ( .A1(n20812), .A2(n20821), .ZN(n1369) );
  NOR2_X1 U4519 ( .A1(n20446), .A2(n1365), .ZN(n1364) );
  AND2_X1 U4520 ( .A1(n20473), .A2(n17639), .ZN(n866) );
  OR2_X1 U4521 ( .A1(n19933), .A2(n20638), .ZN(n21538) );
  NOR2_X1 U4522 ( .A1(n18287), .A2(n6952), .ZN(n1786) );
  AND2_X1 U4523 ( .A1(n18062), .A2(n1715), .ZN(n18333) );
  OR2_X1 U4525 ( .A1(n19424), .A2(n17869), .ZN(n1227) );
  INV_X1 U4526 ( .A(n17557), .ZN(n19411) );
  OR2_X1 U4527 ( .A1(n17311), .A2(n19514), .ZN(n21222) );
  NOR2_X1 U4528 ( .A1(n19276), .A2(n19965), .ZN(n1296) );
  NOR2_X1 U4530 ( .A1(n19957), .A2(n21427), .ZN(n20836) );
  NOR2_X1 U4531 ( .A1(n21407), .A2(n20779), .ZN(n949) );
  INV_X1 U4532 ( .A(n17045), .ZN(n17457) );
  INV_X1 U4533 ( .A(n1715), .ZN(n17544) );
  AND2_X1 U4534 ( .A1(n20063), .A2(n4459), .ZN(n17026) );
  INV_X1 U4535 ( .A(n18865), .ZN(n20681) );
  OR2_X1 U4536 ( .A1(n498), .A2(n20232), .ZN(n18102) );
  OR2_X1 U4537 ( .A1(n21530), .A2(n7431), .ZN(n21527) );
  CLKBUF_X1 U4540 ( .A(n19156), .Z(n21421) );
  BUF_X1 U4541 ( .A(n16834), .Z(n18062) );
  OR2_X1 U4542 ( .A1(n19016), .A2(n8441), .ZN(n19459) );
  INV_X1 U4543 ( .A(n970), .ZN(n20760) );
  INV_X1 U4545 ( .A(n16000), .ZN(n20240) );
  AND2_X1 U4546 ( .A1(n15997), .A2(n20698), .ZN(n18731) );
  INV_X1 U4548 ( .A(n632), .ZN(n1517) );
  INV_X1 U4549 ( .A(n21212), .ZN(n19822) );
  INV_X1 U4550 ( .A(n19289), .ZN(n762) );
  AND2_X1 U4551 ( .A1(n20088), .A2(n17057), .ZN(n18318) );
  OR2_X1 U4552 ( .A1(n20423), .A2(n20357), .ZN(n20362) );
  NAND2_X1 U4556 ( .A1(n2222), .A2(n51374), .ZN(n3181) );
  BUF_X1 U4557 ( .A(n16279), .Z(n19477) );
  CLKBUF_X1 U4558 ( .A(n634), .Z(n21469) );
  INV_X1 U4559 ( .A(n20811), .ZN(n763) );
  INV_X1 U4560 ( .A(n17567), .ZN(n764) );
  NOR2_X1 U4561 ( .A1(n590), .A2(n2166), .ZN(n6168) );
  AND2_X1 U4563 ( .A1(n20795), .A2(n1860), .ZN(n885) );
  NAND2_X1 U4566 ( .A1(n18356), .A2(n18346), .ZN(n19076) );
  OR2_X1 U4571 ( .A1(n19381), .A2(n20383), .ZN(n1788) );
  INV_X1 U4572 ( .A(n631), .ZN(n951) );
  NOR2_X1 U4573 ( .A1(n5192), .A2(n21584), .ZN(n21567) );
  OR2_X1 U4574 ( .A1(n20426), .A2(n20432), .ZN(n850) );
  INV_X1 U4575 ( .A(n598), .ZN(n765) );
  OR2_X1 U4576 ( .A1(n21300), .A2(n18217), .ZN(n18995) );
  INV_X1 U4577 ( .A(n17021), .ZN(n20123) );
  INV_X1 U4579 ( .A(n19156), .ZN(n5500) );
  INV_X1 U4580 ( .A(n1370), .ZN(n1365) );
  INV_X1 U4581 ( .A(n15400), .ZN(n17871) );
  OR2_X1 U4582 ( .A1(n8575), .A2(n21303), .ZN(n19793) );
  AND2_X1 U4583 ( .A1(n20266), .A2(n21664), .ZN(n21653) );
  OR2_X1 U4586 ( .A1(n17639), .A2(n20478), .ZN(n14744) );
  NOR2_X1 U4588 ( .A1(n373), .A2(n51385), .ZN(n19639) );
  INV_X1 U4589 ( .A(n21300), .ZN(n766) );
  XNOR2_X1 U4590 ( .A(n16929), .B(n16928), .ZN(n5083) );
  AND2_X1 U4591 ( .A1(n18217), .A2(n18997), .ZN(n19794) );
  AND2_X1 U4592 ( .A1(n15724), .A2(n19673), .ZN(n18234) );
  AND2_X1 U4593 ( .A1(n18377), .A2(n17047), .ZN(n18381) );
  NAND2_X1 U4594 ( .A1(n18962), .A2(n3885), .ZN(n17079) );
  XNOR2_X1 U4599 ( .A(n5667), .B(n16577), .ZN(n18865) );
  NAND2_X1 U4604 ( .A1(n16792), .A2(n17057), .ZN(n20086) );
  INV_X1 U4605 ( .A(n21460), .ZN(n767) );
  XNOR2_X1 U4611 ( .A(n18606), .B(n2265), .ZN(n19156) );
  INV_X1 U4612 ( .A(n18331), .ZN(n17545) );
  INV_X1 U4613 ( .A(n21392), .ZN(n21388) );
  INV_X1 U4615 ( .A(n21450), .ZN(n1618) );
  OR2_X1 U4616 ( .A1(n18294), .A2(n18288), .ZN(n6363) );
  AND2_X1 U4617 ( .A1(n19514), .A2(n5177), .ZN(n21235) );
  AND2_X1 U4618 ( .A1(n20441), .A2(n20821), .ZN(n20815) );
  INV_X1 U4619 ( .A(n17018), .ZN(n20155) );
  INV_X1 U4621 ( .A(n21397), .ZN(n769) );
  AND2_X1 U4622 ( .A1(n21584), .A2(n21578), .ZN(n20779) );
  NAND2_X1 U4623 ( .A1(n4081), .A2(n17018), .ZN(n19048) );
  INV_X1 U4624 ( .A(n17873), .ZN(n8378) );
  XNOR2_X1 U4627 ( .A(n5700), .B(n5699), .ZN(n20244) );
  INV_X1 U4628 ( .A(n20037), .ZN(n771) );
  INV_X1 U4629 ( .A(n8490), .ZN(n21604) );
  XNOR2_X1 U4630 ( .A(n15919), .B(n15918), .ZN(n20684) );
  CLKBUF_X1 U4631 ( .A(n16986), .Z(n19033) );
  BUF_X1 U4632 ( .A(n15725), .Z(n19679) );
  AND2_X1 U4633 ( .A1(n21303), .A2(n19796), .ZN(n3507) );
  INV_X1 U4634 ( .A(n14381), .ZN(n772) );
  XNOR2_X1 U4636 ( .A(n15534), .B(n15533), .ZN(n17584) );
  XNOR2_X1 U4637 ( .A(n4495), .B(n17660), .ZN(n20488) );
  INV_X1 U4638 ( .A(n19514), .ZN(n773) );
  INV_X1 U4639 ( .A(n21468), .ZN(n774) );
  INV_X1 U4642 ( .A(n20211), .ZN(n775) );
  XNOR2_X1 U4643 ( .A(n17238), .B(n8683), .ZN(n19016) );
  XNOR2_X1 U4644 ( .A(n18787), .B(n18788), .ZN(n21414) );
  XNOR2_X1 U4647 ( .A(n18398), .B(n3766), .ZN(n20638) );
  XNOR2_X1 U4648 ( .A(n15752), .B(n8129), .ZN(n1232) );
  XNOR2_X1 U4649 ( .A(n17801), .B(n17800), .ZN(n17838) );
  XNOR2_X1 U4650 ( .A(n18216), .B(n18215), .ZN(n19795) );
  INV_X1 U4652 ( .A(n20795), .ZN(n776) );
  XNOR2_X1 U4653 ( .A(n7642), .B(n7641), .ZN(n20472) );
  INV_X1 U4654 ( .A(n19989), .ZN(n777) );
  XNOR2_X1 U4655 ( .A(n17724), .B(n17723), .ZN(n21473) );
  INV_X1 U4656 ( .A(n17059), .ZN(n778) );
  XNOR2_X1 U4657 ( .A(n18418), .B(n16247), .ZN(n1480) );
  INV_X1 U4659 ( .A(n16360), .ZN(n1896) );
  CLKBUF_X1 U4660 ( .A(n16328), .Z(n2081) );
  XNOR2_X1 U4662 ( .A(n19235), .B(n1521), .ZN(n16454) );
  INV_X1 U4663 ( .A(n16328), .ZN(n779) );
  XNOR2_X1 U4664 ( .A(n15746), .B(n16661), .ZN(n16770) );
  XNOR2_X1 U4666 ( .A(n16201), .B(n17232), .ZN(n17134) );
  XNOR2_X1 U4668 ( .A(n15903), .B(n2200), .ZN(n16525) );
  INV_X1 U4669 ( .A(n17847), .ZN(n15746) );
  INV_X1 U4673 ( .A(n17887), .ZN(n16952) );
  XNOR2_X1 U4675 ( .A(n14698), .B(n1877), .ZN(n16071) );
  INV_X1 U4676 ( .A(n14698), .ZN(n1878) );
  AND2_X1 U4677 ( .A1(n1437), .A2(n1434), .ZN(n15896) );
  NAND4_X1 U4678 ( .A1(n15311), .A2(n15310), .A3(n15312), .A4(n15313), .ZN(
        n16186) );
  XNOR2_X1 U4680 ( .A(n4979), .B(n18438), .ZN(n17348) );
  INV_X1 U4681 ( .A(n16064), .ZN(n1877) );
  XNOR2_X1 U4682 ( .A(n18202), .B(n4800), .ZN(n18644) );
  XNOR2_X1 U4683 ( .A(n14698), .B(n309), .ZN(n17686) );
  XNOR2_X1 U4686 ( .A(n14698), .B(n1876), .ZN(n17384) );
  AND3_X1 U4689 ( .A1(n10090), .A2(n10091), .A3(n13187), .ZN(n1338) );
  XNOR2_X1 U4690 ( .A(n16470), .B(n16904), .ZN(n8212) );
  XNOR2_X1 U4691 ( .A(n17690), .B(n7191), .ZN(n5611) );
  XNOR2_X1 U4693 ( .A(n14176), .B(n16943), .ZN(n18692) );
  NAND3_X1 U4694 ( .A1(n14326), .A2(n14327), .A3(n1241), .ZN(n17822) );
  AND2_X1 U4697 ( .A1(n15428), .A2(n1831), .ZN(n1834) );
  NAND2_X1 U4700 ( .A1(n5258), .A2(n5257), .ZN(n5256) );
  NAND4_X1 U4701 ( .A1(n12011), .A2(n12010), .A3(n14336), .A4(n12012), .ZN(
        n948) );
  NAND2_X1 U4702 ( .A1(n7156), .A2(n3958), .ZN(n17947) );
  NAND4_X1 U4704 ( .A1(n14078), .A2(n14077), .A3(n14076), .A4(n14075), .ZN(
        n14508) );
  OR2_X1 U4705 ( .A1(n13185), .A2(n13780), .ZN(n3733) );
  AND4_X1 U4706 ( .A1(n13183), .A2(n13182), .A3(n13181), .A4(n13180), .ZN(
        n3732) );
  NOR2_X1 U4707 ( .A1(n10315), .A2(n1063), .ZN(n1062) );
  NAND3_X1 U4710 ( .A1(n15122), .A2(n4249), .A3(n4248), .ZN(n17258) );
  AND2_X1 U4711 ( .A1(n15290), .A2(n15288), .ZN(n1226) );
  AND3_X1 U4714 ( .A1(n4669), .A2(n15110), .A3(n15111), .ZN(n4248) );
  NAND3_X1 U4715 ( .A1(n14565), .A2(n14564), .A3(n14563), .ZN(n17643) );
  AND4_X1 U4717 ( .A1(n11866), .A2(n11859), .A3(n11867), .A4(n12880), .ZN(
        n2972) );
  OR2_X1 U4719 ( .A1(n12424), .A2(n13787), .ZN(n13185) );
  NOR2_X1 U4720 ( .A1(n12934), .A2(n12935), .ZN(n12941) );
  INV_X1 U4721 ( .A(n12416), .ZN(n12423) );
  OR2_X1 U4722 ( .A1(n14329), .A2(n14328), .ZN(n1241) );
  AOI22_X1 U4725 ( .A1(n13014), .A2(n13015), .B1(n13016), .B2(n13017), .ZN(
        n13020) );
  NAND4_X1 U4726 ( .A1(n12898), .A2(n12897), .A3(n12896), .A4(n12895), .ZN(
        n2121) );
  AND2_X1 U4727 ( .A1(n15279), .A2(n14054), .ZN(n1309) );
  AOI21_X1 U4728 ( .B1(n1439), .B2(n1436), .A(n1435), .ZN(n1434) );
  AND2_X1 U4729 ( .A1(n13468), .A2(n13469), .ZN(n1097) );
  AND3_X1 U4730 ( .A1(n12947), .A2(n12945), .A3(n1046), .ZN(n1045) );
  OR2_X1 U4731 ( .A1(n5628), .A2(n2471), .ZN(n1061) );
  OR2_X1 U4733 ( .A1(n13479), .A2(n13794), .ZN(n2023) );
  NOR2_X1 U4734 ( .A1(n1438), .A2(n13440), .ZN(n1435) );
  OR2_X1 U4735 ( .A1(n14786), .A2(n1780), .ZN(n15268) );
  INV_X1 U4737 ( .A(n4443), .ZN(n1096) );
  OAI21_X1 U4738 ( .B1(n15423), .B2(n14875), .A(n1832), .ZN(n1831) );
  AND4_X1 U4739 ( .A1(n12864), .A2(n12863), .A3(n12862), .A4(n14405), .ZN(
        n12875) );
  AND2_X1 U4740 ( .A1(n13993), .A2(n13998), .ZN(n9993) );
  AND3_X1 U4741 ( .A1(n15266), .A2(n14135), .A3(n14136), .ZN(n1961) );
  AND2_X1 U4742 ( .A1(n10638), .A2(n13005), .ZN(n2137) );
  AND2_X1 U4743 ( .A1(n1580), .A2(n13206), .ZN(n1578) );
  AND3_X1 U4744 ( .A1(n13812), .A2(n2061), .A3(n4231), .ZN(n2059) );
  AND2_X1 U4745 ( .A1(n13498), .A2(n13499), .ZN(n1066) );
  AND2_X1 U4746 ( .A1(n13497), .A2(n13496), .ZN(n3462) );
  NOR2_X1 U4747 ( .A1(n12409), .A2(n13296), .ZN(n1909) );
  AND2_X1 U4749 ( .A1(n14122), .A2(n14115), .ZN(n1631) );
  OR2_X1 U4750 ( .A1(n14771), .A2(n15207), .ZN(n14772) );
  OR2_X1 U4751 ( .A1(n14873), .A2(n3704), .ZN(n15416) );
  AOI21_X1 U4752 ( .B1(n13005), .B2(n13004), .A(n13401), .ZN(n14357) );
  OR2_X1 U4753 ( .A1(n14785), .A2(n15257), .ZN(n14786) );
  OR2_X1 U4754 ( .A1(n14133), .A2(n5208), .ZN(n1359) );
  OAI21_X1 U4755 ( .B1(n14635), .B2(n13653), .A(n11303), .ZN(n1046) );
  NOR2_X1 U4756 ( .A1(n2249), .A2(n1554), .ZN(n1553) );
  NAND2_X1 U4757 ( .A1(n14660), .A2(n14652), .ZN(n1439) );
  NOR2_X1 U4758 ( .A1(n1930), .A2(n1929), .ZN(n12828) );
  AND2_X1 U4759 ( .A1(n13441), .A2(n12041), .ZN(n1438) );
  OR2_X1 U4760 ( .A1(n13944), .A2(n638), .ZN(n13953) );
  NOR2_X1 U4761 ( .A1(n15205), .A2(n2014), .ZN(n15187) );
  NAND2_X1 U4762 ( .A1(n11753), .A2(n14657), .ZN(n1448) );
  OAI21_X1 U4763 ( .B1(n14024), .B2(n14023), .A(n14022), .ZN(n2007) );
  OR2_X1 U4765 ( .A1(n14880), .A2(n14870), .ZN(n2249) );
  AND2_X1 U4767 ( .A1(n13505), .A2(n13514), .ZN(n13503) );
  AND2_X1 U4768 ( .A1(n14331), .A2(n13417), .ZN(n13424) );
  OR2_X1 U4770 ( .A1(n6481), .A2(n640), .ZN(n14445) );
  NOR2_X1 U4771 ( .A1(n8075), .A2(n14984), .ZN(n14980) );
  NOR2_X1 U4772 ( .A1(n11762), .A2(n51656), .ZN(n1577) );
  NAND2_X1 U4776 ( .A1(n1556), .A2(n1555), .ZN(n1554) );
  OR2_X1 U4777 ( .A1(n10628), .A2(n7411), .ZN(n13005) );
  AND2_X1 U4778 ( .A1(n1556), .A2(n14880), .ZN(n13256) );
  INV_X1 U4779 ( .A(n14870), .ZN(n1206) );
  OR2_X1 U4780 ( .A1(n13509), .A2(n9358), .ZN(n963) );
  OR2_X1 U4781 ( .A1(n13530), .A2(n11841), .ZN(n960) );
  NOR2_X1 U4783 ( .A1(n11840), .A2(n13525), .ZN(n12765) );
  OR2_X1 U4784 ( .A1(n51018), .A2(n16039), .ZN(n13372) );
  OR2_X1 U4785 ( .A1(n14929), .A2(n7572), .ZN(n15077) );
  NOR3_X1 U4787 ( .A1(n15425), .A2(n2640), .A3(n14870), .ZN(n14877) );
  AND2_X1 U4788 ( .A1(n14791), .A2(n14139), .ZN(n1963) );
  INV_X1 U4789 ( .A(n13006), .ZN(n12224) );
  OR2_X1 U4790 ( .A1(n7688), .A2(n14294), .ZN(n14297) );
  AND2_X1 U4791 ( .A1(n14260), .A2(n10501), .ZN(n13696) );
  NOR2_X1 U4793 ( .A1(n15133), .A2(n15126), .ZN(n13711) );
  INV_X1 U4794 ( .A(n14117), .ZN(n2014) );
  INV_X1 U4795 ( .A(n12886), .ZN(n781) );
  INV_X1 U4796 ( .A(n2189), .ZN(n1486) );
  NAND2_X1 U4797 ( .A1(n11865), .A2(n11765), .ZN(n13204) );
  AND2_X1 U4798 ( .A1(n13174), .A2(n13780), .ZN(n1282) );
  INV_X1 U4799 ( .A(n14533), .ZN(n1283) );
  INV_X1 U4800 ( .A(n15233), .ZN(n2013) );
  NOR2_X1 U4802 ( .A1(n11853), .A2(n15365), .ZN(n15378) );
  AND2_X1 U4803 ( .A1(n13076), .A2(n3081), .ZN(n1930) );
  AND2_X1 U4804 ( .A1(n15440), .A2(n15341), .ZN(n14863) );
  INV_X1 U4807 ( .A(n13849), .ZN(n13854) );
  NOR2_X1 U4809 ( .A1(n51534), .A2(n14601), .ZN(n14612) );
  BUF_X1 U4810 ( .A(n11740), .Z(n14883) );
  AND2_X1 U4811 ( .A1(n14929), .A2(n15067), .ZN(n820) );
  NAND2_X1 U4813 ( .A1(n13514), .A2(n13526), .ZN(n12767) );
  AND2_X1 U4814 ( .A1(n15206), .A2(n15244), .ZN(n14117) );
  INV_X1 U4815 ( .A(n12787), .ZN(n13450) );
  INV_X1 U4816 ( .A(n15068), .ZN(n7572) );
  INV_X1 U4818 ( .A(n12787), .ZN(n2072) );
  AND2_X1 U4819 ( .A1(n14412), .A2(n14070), .ZN(n1111) );
  OR2_X1 U4820 ( .A1(n2062), .A2(n14345), .ZN(n2061) );
  INV_X1 U4824 ( .A(n13296), .ZN(n782) );
  INV_X1 U4825 ( .A(n13885), .ZN(n1555) );
  AND2_X1 U4827 ( .A1(n13820), .A2(n8226), .ZN(n14312) );
  AND2_X1 U4828 ( .A1(n14644), .A2(n9162), .ZN(n13653) );
  INV_X1 U4829 ( .A(n12204), .ZN(n13979) );
  OR2_X1 U4831 ( .A1(n15243), .A2(n15206), .ZN(n14115) );
  OR2_X1 U4834 ( .A1(n14155), .A2(n14149), .ZN(n2556) );
  AND2_X1 U4837 ( .A1(n9162), .A2(n12750), .ZN(n828) );
  AND2_X1 U4838 ( .A1(n14139), .A2(n14137), .ZN(n14141) );
  INV_X1 U4839 ( .A(n13439), .ZN(n12891) );
  OR2_X1 U4840 ( .A1(n14784), .A2(n15256), .ZN(n13057) );
  INV_X1 U4847 ( .A(n14287), .ZN(n784) );
  INV_X1 U4848 ( .A(n15189), .ZN(n1267) );
  AND2_X1 U4850 ( .A1(n51657), .A2(n1571), .ZN(n13941) );
  OR2_X2 U4852 ( .A1(n5832), .A2(n5831), .ZN(n14234) );
  NOR2_X1 U4856 ( .A1(n9695), .A2(n1074), .ZN(n1073) );
  INV_X1 U4857 ( .A(n11841), .ZN(n13506) );
  INV_X1 U4858 ( .A(n13102), .ZN(n1244) );
  AND4_X2 U4859 ( .A1(n2589), .A2(n2586), .A3(n2583), .A4(n2580), .ZN(n14929)
         );
  OR2_X1 U4860 ( .A1(n9720), .A2(n11737), .ZN(n11740) );
  NAND2_X1 U4861 ( .A1(n6382), .A2(n6762), .ZN(n6384) );
  AND2_X1 U4863 ( .A1(n15309), .A2(n14911), .ZN(n14914) );
  INV_X1 U4866 ( .A(n13170), .ZN(n13174) );
  NAND2_X1 U4867 ( .A1(n9616), .A2(n9615), .ZN(n14784) );
  INV_X1 U4869 ( .A(n12890), .ZN(n786) );
  NOR2_X1 U4874 ( .A1(n1571), .A2(n51656), .ZN(n11765) );
  NAND2_X1 U4876 ( .A1(n10644), .A2(n10637), .ZN(n2062) );
  OR2_X1 U4882 ( .A1(n11924), .A2(n11925), .ZN(n15341) );
  AND3_X1 U4884 ( .A1(n4450), .A2(n10035), .A3(n10034), .ZN(n13170) );
  NOR2_X1 U4885 ( .A1(n11607), .A2(n11606), .ZN(n1091) );
  NOR2_X1 U4887 ( .A1(n9561), .A2(n1849), .ZN(n9616) );
  AND3_X1 U4888 ( .A1(n9090), .A2(n9091), .A3(n9092), .ZN(n4586) );
  AND3_X1 U4890 ( .A1(n4881), .A2(n7425), .A3(n11541), .ZN(n14813) );
  AND3_X1 U4891 ( .A1(n9596), .A2(n9595), .A3(n9594), .ZN(n3565) );
  AOI21_X1 U4893 ( .B1(n9195), .B2(n9194), .A(n9193), .ZN(n9196) );
  AND3_X1 U4895 ( .A1(n3980), .A2(n9734), .A3(n9733), .ZN(n9736) );
  OAI21_X1 U4896 ( .B1(n2892), .B2(n9717), .A(n9716), .ZN(n11737) );
  INV_X1 U4899 ( .A(n13172), .ZN(n788) );
  INV_X1 U4900 ( .A(n14339), .ZN(n13412) );
  OR2_X1 U4901 ( .A1(n8457), .A2(n8456), .ZN(n1665) );
  AND4_X1 U4903 ( .A1(n3806), .A2(n3807), .A3(n3805), .A4(n3804), .ZN(n3803)
         );
  AND3_X1 U4905 ( .A1(n9501), .A2(n9502), .A3(n1078), .ZN(n9503) );
  AND3_X1 U4906 ( .A1(n5328), .A2(n10060), .A3(n13227), .ZN(n2073) );
  OAI21_X1 U4908 ( .B1(n3689), .B2(n10700), .A(n12105), .ZN(n860) );
  AND2_X1 U4909 ( .A1(n10577), .A2(n10576), .ZN(n1666) );
  AND2_X1 U4910 ( .A1(n10944), .A2(n10943), .ZN(n1790) );
  OR2_X1 U4912 ( .A1(n9949), .A2(n9950), .ZN(n12790) );
  OAI21_X1 U4913 ( .B1(n10283), .B2(n10284), .A(n1064), .ZN(n4820) );
  OAI22_X1 U4916 ( .A1(n1827), .A2(n1826), .B1(n1825), .B2(n1824), .ZN(n10171)
         );
  AND4_X1 U4917 ( .A1(n10131), .A2(n10130), .A3(n10129), .A4(n10128), .ZN(
        n10132) );
  INV_X1 U4918 ( .A(n9822), .ZN(n10012) );
  AOI22_X1 U4920 ( .A1(n12524), .A2(n10838), .B1(n10837), .B2(n10836), .ZN(
        n10839) );
  AND2_X1 U4922 ( .A1(n12712), .A2(n12435), .ZN(n1784) );
  AND3_X1 U4923 ( .A1(n9027), .A2(n9747), .A3(n3348), .ZN(n9041) );
  INV_X1 U4924 ( .A(n10170), .ZN(n1825) );
  INV_X1 U4925 ( .A(n11022), .ZN(n1827) );
  OR2_X1 U4926 ( .A1(n10157), .A2(n11031), .ZN(n833) );
  AND2_X1 U4927 ( .A1(n10046), .A2(n10556), .ZN(n1461) );
  AND2_X1 U4928 ( .A1(n10149), .A2(n10222), .ZN(n1039) );
  AOI21_X1 U4929 ( .B1(n9377), .B2(n10661), .A(n4464), .ZN(n4463) );
  NOR2_X1 U4930 ( .A1(n8838), .A2(n10223), .ZN(n1040) );
  NOR2_X1 U4932 ( .A1(n7530), .A2(n10456), .ZN(n1999) );
  AOI21_X1 U4933 ( .B1(n3649), .B2(n10281), .A(n870), .ZN(n1064) );
  NAND2_X1 U4935 ( .A1(n9997), .A2(n8410), .ZN(n11040) );
  INV_X1 U4936 ( .A(n2018), .ZN(n12719) );
  OAI21_X1 U4937 ( .B1(n3849), .B2(n3848), .A(n10173), .ZN(n9467) );
  AND2_X1 U4938 ( .A1(n7781), .A2(n11123), .ZN(n12691) );
  AND2_X1 U4939 ( .A1(n9542), .A2(n1307), .ZN(n12613) );
  OR2_X1 U4940 ( .A1(n10182), .A2(n9461), .ZN(n10046) );
  INV_X1 U4941 ( .A(n11387), .ZN(n12062) );
  OR2_X1 U4942 ( .A1(n10134), .A2(n1137), .ZN(n10927) );
  NOR2_X1 U4943 ( .A1(n9484), .A2(n10096), .ZN(n1932) );
  INV_X1 U4944 ( .A(n9585), .ZN(n6147) );
  OAI211_X1 U4945 ( .C1(n12304), .C2(n12300), .A(n9758), .B(n10951), .ZN(n1792) );
  AND2_X1 U4946 ( .A1(n12254), .A2(n12253), .ZN(n1105) );
  OR2_X1 U4947 ( .A1(n12711), .A2(n12705), .ZN(n1782) );
  INV_X1 U4949 ( .A(n9484), .ZN(n8438) );
  INV_X1 U4950 ( .A(n10186), .ZN(n10548) );
  INV_X1 U4951 ( .A(n10003), .ZN(n11025) );
  INV_X1 U4952 ( .A(n12521), .ZN(n11544) );
  OR2_X1 U4953 ( .A1(n10045), .A2(n10182), .ZN(n10042) );
  AND2_X1 U4954 ( .A1(n10580), .A2(n8639), .ZN(n11037) );
  INV_X1 U4955 ( .A(n9539), .ZN(n12590) );
  AND2_X1 U4956 ( .A1(n12292), .A2(n9014), .ZN(n9704) );
  AND2_X1 U4957 ( .A1(n11005), .A2(n876), .ZN(n875) );
  AND2_X1 U4959 ( .A1(n51139), .A2(n9538), .ZN(n11915) );
  AND2_X1 U4961 ( .A1(n9049), .A2(n9045), .ZN(n10673) );
  INV_X1 U4962 ( .A(n10455), .ZN(n789) );
  AND2_X1 U4964 ( .A1(n12166), .A2(n9235), .ZN(n12171) );
  INV_X1 U4965 ( .A(n33567), .ZN(n1876) );
  AND2_X1 U4966 ( .A1(n12635), .A2(n10465), .ZN(n12628) );
  INV_X1 U4970 ( .A(n11023), .ZN(n790) );
  AND2_X1 U4975 ( .A1(n12277), .A2(n12285), .ZN(n10723) );
  INV_X1 U4978 ( .A(n10584), .ZN(n1281) );
  AND2_X1 U4980 ( .A1(n9510), .A2(n9939), .ZN(n11648) );
  AND2_X1 U4982 ( .A1(n11345), .A2(n10734), .ZN(n12254) );
  INV_X1 U4983 ( .A(n51139), .ZN(n1307) );
  AND2_X1 U4984 ( .A1(n12291), .A2(n12277), .ZN(n10726) );
  OR2_X1 U4986 ( .A1(n10526), .A2(n10519), .ZN(n1208) );
  INV_X1 U4987 ( .A(n51762), .ZN(n876) );
  AND2_X1 U4989 ( .A1(n10831), .A2(n12518), .ZN(n12521) );
  NAND2_X1 U4992 ( .A1(n11704), .A2(n9139), .ZN(n11711) );
  INV_X1 U4993 ( .A(n11210), .ZN(n791) );
  AND2_X1 U4997 ( .A1(n9425), .A2(n9647), .ZN(n12253) );
  NAND2_X1 U4999 ( .A1(n9103), .A2(n7482), .ZN(n11460) );
  INV_X1 U5000 ( .A(n8050), .ZN(n793) );
  AND2_X1 U5001 ( .A1(n4555), .A2(n9519), .ZN(n11270) );
  INV_X1 U5005 ( .A(n10513), .ZN(n10522) );
  CLKBUF_X1 U5007 ( .A(n9605), .Z(n12132) );
  NAND2_X1 U5008 ( .A1(n9419), .A2(n10741), .ZN(n12258) );
  OR2_X1 U5009 ( .A1(n51761), .A2(n9830), .ZN(n10186) );
  AND2_X1 U5011 ( .A1(n10419), .A2(n12161), .ZN(n12178) );
  BUF_X1 U5013 ( .A(n8961), .Z(n11123) );
  CLKBUF_X1 U5015 ( .A(n9510), .Z(n10566) );
  INV_X1 U5016 ( .A(n10445), .ZN(n794) );
  BUF_X1 U5018 ( .A(n9519), .Z(n10589) );
  OR2_X1 U5019 ( .A1(n9335), .A2(n9339), .ZN(n11268) );
  CLKBUF_X1 U5020 ( .A(n9336), .Z(n9340) );
  INV_X1 U5021 ( .A(n10419), .ZN(n12169) );
  BUF_X1 U5024 ( .A(n9056), .Z(n12303) );
  BUF_X1 U5027 ( .A(n9147), .Z(n9932) );
  AND2_X1 U5028 ( .A1(n12602), .A2(n9547), .ZN(n9542) );
  AND2_X1 U5030 ( .A1(n9459), .A2(n10552), .ZN(n10174) );
  AND2_X1 U5031 ( .A1(n9417), .A2(n10742), .ZN(n12257) );
  OR2_X1 U5032 ( .A1(n9057), .A2(n12315), .ZN(n12300) );
  INV_X1 U5033 ( .A(n9830), .ZN(n10536) );
  BUF_X1 U5035 ( .A(n9004), .Z(n12277) );
  AND2_X1 U5036 ( .A1(n11932), .A2(n12700), .ZN(n10487) );
  BUF_X1 U5038 ( .A(n9365), .Z(n10687) );
  OR2_X1 U5039 ( .A1(n10959), .A2(n10127), .ZN(n10954) );
  AND2_X1 U5042 ( .A1(n10360), .A2(n9218), .ZN(n10665) );
  NOR2_X1 U5049 ( .A1(n11611), .A2(n11608), .ZN(n11591) );
  AND2_X1 U5051 ( .A1(n12542), .A2(n8945), .ZN(n11445) );
  NAND2_X1 U5053 ( .A1(n2976), .A2(n9104), .ZN(n11630) );
  INV_X1 U5055 ( .A(n9098), .ZN(n11468) );
  XNOR2_X1 U5056 ( .A(n9231), .B(Key[73]), .ZN(n9234) );
  INV_X1 U5057 ( .A(n50546), .ZN(n6031) );
  BUF_X1 U5058 ( .A(n8945), .Z(n12538) );
  INV_X1 U5059 ( .A(n12659), .ZN(n796) );
  INV_X1 U5060 ( .A(n11978), .ZN(n797) );
  BUF_X1 U5063 ( .A(n9153), .Z(n12516) );
  CLKBUF_X1 U5064 ( .A(n26297), .Z(n2606) );
  BUF_X1 U5065 ( .A(n9073), .Z(n11588) );
  BUF_X1 U5067 ( .A(n9292), .Z(n10607) );
  CLKBUF_X1 U5070 ( .A(n9103), .Z(n11619) );
  XNOR2_X1 U5071 ( .A(n8772), .B(Key[168]), .ZN(n11016) );
  CLKBUF_X1 U5072 ( .A(n9098), .Z(n11226) );
  INV_X1 U5073 ( .A(n9218), .ZN(n799) );
  CLKBUF_X1 U5074 ( .A(n9384), .Z(n12058) );
  INV_X1 U5077 ( .A(n48064), .ZN(n5016) );
  INV_X1 U5079 ( .A(n48614), .ZN(n2112) );
  XNOR2_X1 U5081 ( .A(n9403), .B(Key[50]), .ZN(n11376) );
  INV_X1 U5082 ( .A(n11899), .ZN(n800) );
  BUF_X1 U5084 ( .A(Key[147]), .Z(n4739) );
  XNOR2_X1 U5085 ( .A(Key[48]), .B(Ciphertext[77]), .ZN(n11186) );
  INV_X1 U5086 ( .A(n43368), .ZN(n801) );
  XNOR2_X2 U5087 ( .A(Key[78]), .B(Key[54]), .ZN(n29662) );
  BUF_X1 U5088 ( .A(Key[141]), .Z(n4793) );
  CLKBUF_X1 U5089 ( .A(Key[180]), .Z(n1326) );
  CLKBUF_X1 U5090 ( .A(Key[69]), .Z(n4431) );
  CLKBUF_X1 U5091 ( .A(Key[142]), .Z(n4486) );
  CLKBUF_X1 U5092 ( .A(Key[113]), .Z(n4287) );
  INV_X1 U5093 ( .A(n12690), .ZN(n802) );
  CLKBUF_X1 U5094 ( .A(Key[133]), .Z(n4782) );
  CLKBUF_X1 U5096 ( .A(Key[116]), .Z(n4817) );
  CLKBUF_X1 U5097 ( .A(Key[53]), .Z(n4781) );
  INV_X1 U5098 ( .A(n9465), .ZN(n803) );
  XNOR2_X1 U5100 ( .A(Key[88]), .B(Ciphertext[165]), .ZN(n9667) );
  XNOR2_X1 U5101 ( .A(Key[57]), .B(Ciphertext[92]), .ZN(n9926) );
  XNOR2_X1 U5102 ( .A(Key[126]), .B(Ciphertext[143]), .ZN(n10919) );
  INV_X1 U5105 ( .A(n10296), .ZN(n804) );
  CLKBUF_X1 U5106 ( .A(Key[18]), .Z(n4542) );
  INV_X1 U5107 ( .A(n8795), .ZN(n805) );
  CLKBUF_X1 U5108 ( .A(Key[98]), .Z(n2903) );
  XNOR2_X1 U5109 ( .A(Key[127]), .B(Ciphertext[102]), .ZN(n11640) );
  CLKBUF_X2 U5110 ( .A(Key[20]), .Z(n47737) );
  CLKBUF_X1 U5111 ( .A(Key[161]), .Z(n4612) );
  INV_X1 U5113 ( .A(n21837), .ZN(n1774) );
  NOR2_X1 U5114 ( .A1(n15424), .A2(n1206), .ZN(n1205) );
  NAND3_X1 U5115 ( .A1(n4540), .A2(n790), .A3(n10580), .ZN(n807) );
  NAND2_X1 U5116 ( .A1(n806), .A2(n2503), .ZN(n5643) );
  NAND2_X1 U5117 ( .A1(n806), .A2(n5645), .ZN(n5644) );
  XNOR2_X1 U5120 ( .A(n51438), .B(n637), .ZN(n18524) );
  XNOR2_X2 U5121 ( .A(n18682), .B(n18683), .ZN(n21355) );
  AND3_X1 U5123 ( .A1(n13427), .A2(n13406), .A3(n13405), .ZN(n808) );
  NAND2_X1 U5125 ( .A1(n47869), .A2(n47831), .ZN(n47875) );
  NAND2_X1 U5126 ( .A1(n29627), .A2(n2509), .ZN(n4228) );
  NAND2_X1 U5127 ( .A1(n809), .A2(n41911), .ZN(n919) );
  NAND3_X1 U5128 ( .A1(n1259), .A2(n41884), .A3(n48200), .ZN(n809) );
  XNOR2_X1 U5129 ( .A(n42953), .B(n43645), .ZN(n810) );
  NOR2_X2 U5130 ( .A1(n811), .A2(n1264), .ZN(n36500) );
  NAND3_X1 U5132 ( .A1(n5540), .A2(n639), .A3(n13219), .ZN(n14233) );
  OAI21_X1 U5133 ( .B1(n5110), .B2(n32214), .A(n32193), .ZN(n32196) );
  INV_X1 U5134 ( .A(n36082), .ZN(n36086) );
  XNOR2_X1 U5135 ( .A(n51750), .B(n25883), .ZN(n24924) );
  NAND2_X1 U5137 ( .A1(n37666), .A2(n35405), .ZN(n812) );
  NAND2_X1 U5138 ( .A1(n29873), .A2(n813), .ZN(n29694) );
  NAND2_X1 U5140 ( .A1(n12110), .A2(n11365), .ZN(n11366) );
  NAND2_X1 U5141 ( .A1(n9408), .A2(n10701), .ZN(n12110) );
  XNOR2_X1 U5143 ( .A(n15668), .B(n15669), .ZN(n15983) );
  NOR2_X1 U5145 ( .A1(n26969), .A2(n7091), .ZN(n814) );
  NAND3_X1 U5146 ( .A1(n40584), .A2(n40585), .A3(n40586), .ZN(n815) );
  NAND3_X2 U5148 ( .A1(n24360), .A2(n7007), .A3(n7006), .ZN(n32252) );
  NAND2_X1 U5150 ( .A1(n11056), .A2(n15264), .ZN(n816) );
  NAND2_X1 U5151 ( .A1(n1419), .A2(n19070), .ZN(n16804) );
  INV_X1 U5152 ( .A(n11813), .ZN(n5650) );
  XNOR2_X1 U5154 ( .A(n817), .B(n16543), .ZN(n16545) );
  XNOR2_X1 U5155 ( .A(n16538), .B(n16537), .ZN(n817) );
  NAND3_X1 U5156 ( .A1(n6177), .A2(n19310), .A3(n19352), .ZN(n6176) );
  NAND2_X1 U5157 ( .A1(n10261), .A2(n9786), .ZN(n9780) );
  NAND4_X2 U5161 ( .A1(n39089), .A2(n39087), .A3(n39088), .A4(n39086), .ZN(
        n42170) );
  NAND2_X1 U5162 ( .A1(n821), .A2(n820), .ZN(n13790) );
  NAND2_X1 U5163 ( .A1(n13789), .A2(n13788), .ZN(n821) );
  OR2_X1 U5164 ( .A1(n21122), .A2(n21780), .ZN(n22285) );
  NAND3_X1 U5165 ( .A1(n13206), .A2(n6668), .A3(n13949), .ZN(n13944) );
  NAND3_X2 U5167 ( .A1(n26697), .A2(n26696), .A3(n26695), .ZN(n31816) );
  XNOR2_X1 U5171 ( .A(n6658), .B(n25478), .ZN(n29182) );
  XNOR2_X1 U5172 ( .A(n36950), .B(n823), .ZN(n36954) );
  XNOR2_X1 U5173 ( .A(n36951), .B(n36949), .ZN(n823) );
  OAI21_X1 U5174 ( .B1(n6913), .B2(n21872), .A(n6915), .ZN(n943) );
  NOR2_X1 U5175 ( .A1(n38637), .A2(n197), .ZN(n37228) );
  NAND3_X1 U5176 ( .A1(n5141), .A2(n27716), .A3(n27717), .ZN(n855) );
  NAND3_X1 U5177 ( .A1(n4547), .A2(n39525), .A3(n39526), .ZN(n3452) );
  NAND2_X1 U5180 ( .A1(n49492), .A2(n7209), .ZN(n49483) );
  NAND3_X1 U5181 ( .A1(n46282), .A2(n45937), .A3(n46292), .ZN(n43424) );
  NAND3_X1 U5182 ( .A1(n27586), .A2(n27585), .A3(n27584), .ZN(n7925) );
  NAND2_X1 U5183 ( .A1(n27683), .A2(n824), .ZN(n27584) );
  XNOR2_X1 U5184 ( .A(n43320), .B(n825), .ZN(n43321) );
  XNOR2_X1 U5185 ( .A(n52125), .B(n43319), .ZN(n825) );
  XNOR2_X1 U5186 ( .A(n826), .B(n45027), .ZN(Plaintext[115]) );
  NAND3_X1 U5187 ( .A1(n3899), .A2(n3898), .A3(n3896), .ZN(n826) );
  NAND2_X1 U5188 ( .A1(n3254), .A2(n828), .ZN(n14634) );
  XNOR2_X1 U5189 ( .A(n322), .B(n27420), .ZN(n27334) );
  NAND2_X1 U5191 ( .A1(n23756), .A2(n24186), .ZN(n24182) );
  NAND3_X1 U5192 ( .A1(n50021), .A2(n49673), .A3(n49667), .ZN(n45958) );
  NAND2_X2 U5193 ( .A1(n829), .A2(n28495), .ZN(n34141) );
  NAND2_X1 U5196 ( .A1(n40725), .A2(n6325), .ZN(n3252) );
  NAND3_X1 U5197 ( .A1(n24184), .A2(n6718), .A3(n24183), .ZN(n24196) );
  XNOR2_X1 U5199 ( .A(n556), .B(n16466), .ZN(n16468) );
  NAND3_X1 U5200 ( .A1(n17093), .A2(n19535), .A3(n17094), .ZN(n17095) );
  NAND2_X1 U5201 ( .A1(n20122), .A2(n20124), .ZN(n17093) );
  NAND2_X1 U5202 ( .A1(n30051), .A2(n51744), .ZN(n27075) );
  NAND2_X1 U5203 ( .A1(n39942), .A2(n39938), .ZN(n39950) );
  NAND2_X1 U5204 ( .A1(n20652), .A2(n16891), .ZN(n6627) );
  NAND4_X1 U5205 ( .A1(n833), .A2(n1422), .A3(n10167), .A4(n10168), .ZN(n1421)
         );
  AND3_X1 U5206 ( .A1(n20978), .A2(n20976), .A3(n20977), .ZN(n834) );
  OAI22_X1 U5210 ( .A1(n15089), .A2(n20018), .B1(n17489), .B2(n2166), .ZN(
        n15099) );
  AOI21_X1 U5211 ( .B1(n1694), .B2(n29224), .A(n5793), .ZN(n5792) );
  XNOR2_X1 U5212 ( .A(n835), .B(n17349), .ZN(n16232) );
  XNOR2_X1 U5213 ( .A(n16525), .B(n16230), .ZN(n835) );
  NAND4_X1 U5214 ( .A1(n5708), .A2(n48856), .A3(n48857), .A4(n48858), .ZN(
        n4124) );
  OAI21_X1 U5215 ( .B1(n16220), .B2(n837), .A(n836), .ZN(n16224) );
  OR2_X1 U5217 ( .A1(n16219), .A2(n16221), .ZN(n837) );
  NAND3_X1 U5218 ( .A1(n14060), .A2(n14951), .A3(n14950), .ZN(n13724) );
  INV_X1 U5219 ( .A(n9892), .ZN(n11589) );
  NAND2_X1 U5220 ( .A1(n23590), .A2(n23066), .ZN(n23604) );
  NAND4_X1 U5223 ( .A1(n39878), .A2(n39879), .A3(n39880), .A4(n39881), .ZN(
        n40998) );
  NAND3_X1 U5224 ( .A1(n12431), .A2(n13354), .A3(n13347), .ZN(n12432) );
  NAND3_X1 U5225 ( .A1(n1881), .A2(n30765), .A3(n1882), .ZN(n1880) );
  NAND2_X1 U5228 ( .A1(n51377), .A2(n38448), .ZN(n38455) );
  NAND3_X1 U5229 ( .A1(n910), .A2(n8649), .A3(n27746), .ZN(n6111) );
  NAND3_X1 U5230 ( .A1(n732), .A2(n29455), .A3(n29469), .ZN(n27746) );
  NAND3_X1 U5232 ( .A1(n1262), .A2(n15999), .A3(n20249), .ZN(n1453) );
  NAND2_X1 U5233 ( .A1(n31380), .A2(n33014), .ZN(n3525) );
  NAND2_X1 U5234 ( .A1(n7459), .A2(n50681), .ZN(n50665) );
  NAND2_X1 U5236 ( .A1(n28970), .A2(n29718), .ZN(n29724) );
  NAND2_X1 U5239 ( .A1(n42131), .A2(n8332), .ZN(n42148) );
  NAND2_X1 U5240 ( .A1(n31263), .A2(n31262), .ZN(n35748) );
  AND2_X1 U5241 ( .A1(n42136), .A2(n41770), .ZN(n40886) );
  NAND2_X2 U5242 ( .A1(n843), .A2(n3741), .ZN(n31870) );
  AOI21_X1 U5245 ( .B1(n17518), .B2(n17517), .A(n844), .ZN(n17540) );
  NAND2_X1 U5246 ( .A1(n17519), .A2(n17520), .ZN(n844) );
  INV_X1 U5247 ( .A(n24675), .ZN(n29422) );
  INV_X1 U5248 ( .A(n21018), .ZN(n21921) );
  AOI22_X1 U5249 ( .A1(n32206), .A2(n929), .B1(n30888), .B2(n32214), .ZN(
        n29108) );
  NAND4_X2 U5250 ( .A1(n19599), .A2(n19598), .A3(n19600), .A4(n19601), .ZN(
        n25747) );
  NAND4_X1 U5252 ( .A1(n38872), .A2(n38877), .A3(n41084), .A4(n38871), .ZN(
        n845) );
  NAND2_X1 U5254 ( .A1(n29181), .A2(n6660), .ZN(n846) );
  AOI21_X1 U5256 ( .B1(n849), .B2(n18061), .A(n848), .ZN(n847) );
  NOR2_X1 U5257 ( .A1(n17430), .A2(n18061), .ZN(n848) );
  INV_X1 U5258 ( .A(n17429), .ZN(n849) );
  NAND2_X1 U5259 ( .A1(n5875), .A2(n850), .ZN(n20429) );
  NAND2_X1 U5260 ( .A1(n20522), .A2(n22717), .ZN(n851) );
  NAND2_X1 U5261 ( .A1(n8240), .A2(n29828), .ZN(n8239) );
  NAND3_X1 U5262 ( .A1(n19287), .A2(n20771), .A3(n21597), .ZN(n3284) );
  NAND3_X1 U5264 ( .A1(n12174), .A2(n548), .A3(n12171), .ZN(n9237) );
  NAND2_X2 U5266 ( .A1(n4113), .A2(n5568), .ZN(n30592) );
  NAND2_X1 U5267 ( .A1(n38204), .A2(n38572), .ZN(n35704) );
  NAND3_X1 U5268 ( .A1(n36525), .A2(n36535), .A3(n36524), .ZN(n36526) );
  NAND2_X1 U5269 ( .A1(n47778), .A2(n47763), .ZN(n47711) );
  OR2_X2 U5270 ( .A1(n36122), .A2(n35666), .ZN(n38589) );
  NAND3_X1 U5271 ( .A1(n22116), .A2(n23209), .A3(n18369), .ZN(n20304) );
  NAND4_X1 U5272 ( .A1(n13424), .A2(n13423), .A3(n14352), .A4(n13425), .ZN(
        n13426) );
  OR2_X2 U5273 ( .A1(n32943), .A2(n32944), .ZN(n33722) );
  NAND2_X1 U5274 ( .A1(n30819), .A2(n32135), .ZN(n32943) );
  NAND4_X1 U5275 ( .A1(n37433), .A2(n37447), .A3(n37434), .A4(n852), .ZN(n5308) );
  NAND3_X1 U5278 ( .A1(n853), .A2(n39371), .A3(n39372), .ZN(n39373) );
  NAND2_X1 U5279 ( .A1(n39370), .A2(n39378), .ZN(n853) );
  AOI21_X1 U5280 ( .B1(n31610), .B2(n624), .A(n32559), .ZN(n31611) );
  NAND2_X1 U5283 ( .A1(n5140), .A2(n855), .ZN(n1136) );
  NAND2_X1 U5284 ( .A1(n729), .A2(n28615), .ZN(n6058) );
  NAND2_X1 U5285 ( .A1(n34674), .A2(n37559), .ZN(n34680) );
  NAND2_X1 U5286 ( .A1(n37437), .A2(n37438), .ZN(n37480) );
  INV_X1 U5287 ( .A(n856), .ZN(n38824) );
  OAI211_X1 U5288 ( .C1(n934), .C2(n41789), .A(n38813), .B(n38814), .ZN(n856)
         );
  INV_X1 U5289 ( .A(n51474), .ZN(n3735) );
  NAND2_X1 U5291 ( .A1(n2997), .A2(n4307), .ZN(n2149) );
  INV_X1 U5292 ( .A(n28568), .ZN(n28565) );
  INV_X1 U5293 ( .A(n37562), .ZN(n37550) );
  NAND2_X1 U5296 ( .A1(n28991), .A2(n30461), .ZN(n28990) );
  NAND2_X1 U5297 ( .A1(n1011), .A2(n38119), .ZN(n1012) );
  NAND3_X1 U5298 ( .A1(n10764), .A2(n14595), .A3(n14171), .ZN(n4262) );
  NAND2_X1 U5299 ( .A1(n858), .A2(n857), .ZN(n30236) );
  NAND2_X1 U5300 ( .A1(n3594), .A2(n30232), .ZN(n858) );
  NAND2_X2 U5301 ( .A1(n859), .A2(n41336), .ZN(n44314) );
  NAND4_X2 U5302 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n860), .ZN(
        n14605) );
  NAND2_X1 U5304 ( .A1(n3416), .A2(n36400), .ZN(n861) );
  NAND2_X1 U5305 ( .A1(n29371), .A2(n29370), .ZN(n862) );
  NAND2_X1 U5307 ( .A1(n38365), .A2(n4577), .ZN(n1185) );
  NAND2_X1 U5308 ( .A1(n31238), .A2(n31244), .ZN(n31788) );
  NAND2_X1 U5309 ( .A1(n48549), .A2(n2663), .ZN(n2662) );
  NAND2_X1 U5310 ( .A1(n863), .A2(n12354), .ZN(n8798) );
  NAND2_X1 U5311 ( .A1(n9781), .A2(n51137), .ZN(n863) );
  NAND2_X1 U5312 ( .A1(n12358), .A2(n12350), .ZN(n9781) );
  INV_X1 U5313 ( .A(n22142), .ZN(n975) );
  NAND4_X2 U5314 ( .A1(n11790), .A2(n11791), .A3(n11793), .A4(n11792), .ZN(
        n18832) );
  NAND2_X1 U5315 ( .A1(n4753), .A2(n36202), .ZN(n1807) );
  AND3_X1 U5316 ( .A1(n31272), .A2(n31271), .A3(n8203), .ZN(n31278) );
  NAND2_X1 U5317 ( .A1(n21938), .A2(n865), .ZN(n20953) );
  NAND2_X1 U5318 ( .A1(n22143), .A2(n21018), .ZN(n865) );
  NAND2_X1 U5319 ( .A1(n31108), .A2(n31109), .ZN(n31128) );
  NAND4_X4 U5320 ( .A1(n11892), .A2(n13894), .A3(n13895), .A4(n13896), .ZN(
        n15437) );
  AND4_X2 U5321 ( .A1(n16685), .A2(n16683), .A3(n16682), .A4(n16686), .ZN(
        n23473) );
  NAND2_X1 U5322 ( .A1(n20432), .A2(n20428), .ZN(n18053) );
  XNOR2_X2 U5323 ( .A(n17769), .B(n18526), .ZN(n20428) );
  NAND3_X1 U5324 ( .A1(n20436), .A2(n19173), .A3(n20354), .ZN(n18051) );
  NAND2_X1 U5325 ( .A1(n19378), .A2(n20466), .ZN(n867) );
  INV_X1 U5326 ( .A(n37654), .ZN(n38720) );
  NAND4_X1 U5327 ( .A1(n41359), .A2(n41358), .A3(n1410), .A4(n41360), .ZN(
        n1409) );
  NOR2_X1 U5328 ( .A1(n18847), .A2(n317), .ZN(n18848) );
  NOR2_X1 U5329 ( .A1(n31146), .A2(n31425), .ZN(n2609) );
  NOR2_X1 U5330 ( .A1(n746), .A2(n52147), .ZN(n29241) );
  NOR2_X1 U5331 ( .A1(n27578), .A2(n1482), .ZN(n26811) );
  NOR2_X1 U5332 ( .A1(n40032), .A2(n40033), .ZN(n40664) );
  NAND2_X1 U5333 ( .A1(n10018), .A2(n11658), .ZN(n10569) );
  NAND2_X1 U5335 ( .A1(n38301), .A2(n39236), .ZN(n869) );
  NAND2_X1 U5336 ( .A1(n3827), .A2(n28860), .ZN(n28948) );
  INV_X1 U5337 ( .A(n10282), .ZN(n870) );
  NAND3_X1 U5338 ( .A1(n24238), .A2(n24237), .A3(n24239), .ZN(n24240) );
  NAND2_X1 U5340 ( .A1(n3983), .A2(n29273), .ZN(n871) );
  NOR2_X1 U5341 ( .A1(n32128), .A2(n872), .ZN(n31702) );
  NAND2_X1 U5346 ( .A1(n6060), .A2(n38811), .ZN(n4738) );
  NOR2_X1 U5347 ( .A1(n49503), .A2(n2193), .ZN(n49487) );
  NAND2_X1 U5348 ( .A1(n46449), .A2(n48465), .ZN(n46437) );
  NAND3_X1 U5350 ( .A1(n4604), .A2(n12310), .A3(n10292), .ZN(n9769) );
  NAND4_X1 U5351 ( .A1(n874), .A2(n32623), .A3(n32621), .A4(n32622), .ZN(
        n32624) );
  NAND2_X1 U5352 ( .A1(n1890), .A2(n32618), .ZN(n874) );
  NOR2_X2 U5353 ( .A1(n12065), .A2(n12064), .ZN(n14545) );
  NAND3_X1 U5354 ( .A1(n26994), .A2(n29426), .A3(n877), .ZN(n24672) );
  OR2_X1 U5355 ( .A1(n26901), .A2(n27711), .ZN(n877) );
  NAND3_X1 U5357 ( .A1(n43483), .A2(n43482), .A3(n43484), .ZN(n43485) );
  NAND2_X1 U5358 ( .A1(n51090), .A2(n20230), .ZN(n20231) );
  XNOR2_X2 U5359 ( .A(n15870), .B(n1480), .ZN(n20230) );
  NAND2_X1 U5360 ( .A1(n32894), .A2(n32899), .ZN(n32631) );
  AOI21_X1 U5361 ( .B1(n34920), .B2(n41645), .A(n41647), .ZN(n7367) );
  NAND2_X1 U5362 ( .A1(n31599), .A2(n879), .ZN(n878) );
  NAND3_X1 U5365 ( .A1(n8275), .A2(n1162), .A3(n1163), .ZN(n8272) );
  NAND3_X1 U5366 ( .A1(n7666), .A2(n32503), .A3(n32507), .ZN(n31992) );
  NAND2_X1 U5368 ( .A1(n7665), .A2(n48480), .ZN(n4787) );
  NOR2_X1 U5369 ( .A1(n45614), .A2(n7275), .ZN(n881) );
  AOI21_X1 U5370 ( .B1(n46417), .B2(n48448), .A(n883), .ZN(n882) );
  NAND4_X1 U5371 ( .A1(n884), .A2(n20373), .A3(n20374), .A4(n769), .ZN(n20382)
         );
  NAND2_X1 U5372 ( .A1(n21398), .A2(n885), .ZN(n884) );
  NAND3_X1 U5373 ( .A1(n22771), .A2(n2534), .A3(n22770), .ZN(n886) );
  NAND3_X1 U5376 ( .A1(n21868), .A2(n21867), .A3(n22251), .ZN(n939) );
  NAND2_X1 U5377 ( .A1(n8941), .A2(n12536), .ZN(n11089) );
  XNOR2_X1 U5378 ( .A(n888), .B(n34026), .ZN(n33852) );
  XNOR2_X1 U5379 ( .A(n33850), .B(n37097), .ZN(n888) );
  NAND2_X1 U5380 ( .A1(n38939), .A2(n39421), .ZN(n896) );
  NAND2_X1 U5381 ( .A1(n38951), .A2(n39423), .ZN(n39421) );
  NAND2_X1 U5382 ( .A1(n19732), .A2(n19006), .ZN(n4623) );
  NAND2_X1 U5384 ( .A1(n42109), .A2(n2529), .ZN(n889) );
  NAND2_X1 U5388 ( .A1(n40453), .A2(n40446), .ZN(n39979) );
  NAND4_X1 U5389 ( .A1(n14489), .A2(n14492), .A3(n14490), .A4(n14491), .ZN(
        n14493) );
  INV_X1 U5390 ( .A(n18047), .ZN(n984) );
  NAND2_X1 U5391 ( .A1(n5165), .A2(n21811), .ZN(n891) );
  NOR2_X1 U5392 ( .A1(n891), .A2(n1745), .ZN(n1744) );
  NAND2_X1 U5393 ( .A1(n24240), .A2(n891), .ZN(n24241) );
  NAND2_X1 U5394 ( .A1(n892), .A2(n31910), .ZN(n28945) );
  NAND2_X1 U5395 ( .A1(n30491), .A2(n32381), .ZN(n892) );
  NAND2_X1 U5396 ( .A1(n894), .A2(n893), .ZN(n30491) );
  NOR2_X1 U5397 ( .A1(n713), .A2(n32843), .ZN(n893) );
  INV_X1 U5398 ( .A(n32851), .ZN(n894) );
  NOR2_X1 U5400 ( .A1(n32424), .A2(n895), .ZN(n32427) );
  NAND2_X1 U5402 ( .A1(n896), .A2(n39204), .ZN(n899) );
  NAND2_X1 U5404 ( .A1(n32815), .A2(n900), .ZN(n32828) );
  NAND2_X1 U5405 ( .A1(n900), .A2(n31398), .ZN(n32822) );
  NOR2_X1 U5406 ( .A1(n8542), .A2(n900), .ZN(n30473) );
  NAND3_X1 U5407 ( .A1(n3011), .A2(n32831), .A3(n900), .ZN(n3010) );
  NAND2_X1 U5408 ( .A1(n39208), .A2(n39210), .ZN(n38651) );
  NAND3_X1 U5409 ( .A1(n39204), .A2(n39208), .A3(n39423), .ZN(n36889) );
  NAND2_X1 U5410 ( .A1(n39414), .A2(n902), .ZN(n39415) );
  NAND4_X1 U5411 ( .A1(n36888), .A2(n39208), .A3(n38953), .A4(n38946), .ZN(
        n36892) );
  NAND2_X1 U5413 ( .A1(n20726), .A2(n904), .ZN(n903) );
  NAND3_X1 U5414 ( .A1(n26642), .A2(n907), .A3(n27830), .ZN(n26644) );
  NAND2_X1 U5415 ( .A1(n1022), .A2(n430), .ZN(n906) );
  INV_X1 U5416 ( .A(n29439), .ZN(n26069) );
  XNOR2_X1 U5417 ( .A(n34294), .B(n908), .ZN(n33312) );
  XNOR2_X1 U5418 ( .A(n36758), .B(n909), .ZN(n36880) );
  INV_X1 U5419 ( .A(n47244), .ZN(n909) );
  MUX2_X1 U5420 ( .A(n41574), .B(n41575), .S(n41513), .Z(n41592) );
  NAND2_X1 U5422 ( .A1(n24562), .A2(n911), .ZN(n910) );
  NAND2_X1 U5423 ( .A1(n26786), .A2(n29472), .ZN(n911) );
  NAND2_X1 U5424 ( .A1(n29469), .A2(n27758), .ZN(n26786) );
  NAND2_X1 U5425 ( .A1(n913), .A2(n48487), .ZN(n44674) );
  NAND3_X1 U5426 ( .A1(n913), .A2(n48247), .A3(n48248), .ZN(n48249) );
  OAI21_X1 U5427 ( .B1(n48488), .B2(n48487), .A(n913), .ZN(n48489) );
  OAI211_X1 U5428 ( .C1(n48488), .C2(n48482), .A(n913), .B(n48474), .ZN(n45606) );
  NAND2_X1 U5429 ( .A1(n913), .A2(n48244), .ZN(n48473) );
  OR2_X1 U5430 ( .A1(n8097), .A2(n913), .ZN(n8096) );
  NAND3_X1 U5431 ( .A1(n45600), .A2(n913), .A3(n48478), .ZN(n45602) );
  OR2_X1 U5432 ( .A1(n46458), .A2(n913), .ZN(n912) );
  NAND2_X1 U5434 ( .A1(n915), .A2(n47875), .ZN(n47826) );
  NAND3_X1 U5435 ( .A1(n47873), .A2(n47824), .A3(n51469), .ZN(n915) );
  NAND2_X1 U5436 ( .A1(n41919), .A2(n45545), .ZN(n916) );
  NAND2_X1 U5437 ( .A1(n41920), .A2(n45002), .ZN(n918) );
  NAND2_X1 U5440 ( .A1(n30828), .A2(n30648), .ZN(n924) );
  NAND2_X1 U5441 ( .A1(n31298), .A2(n926), .ZN(n925) );
  NAND2_X1 U5442 ( .A1(n29650), .A2(n4936), .ZN(n926) );
  NAND2_X1 U5443 ( .A1(n928), .A2(n30834), .ZN(n927) );
  NAND2_X1 U5444 ( .A1(n30641), .A2(n30640), .ZN(n928) );
  NAND2_X1 U5445 ( .A1(n32207), .A2(n32197), .ZN(n929) );
  NAND3_X1 U5446 ( .A1(n38810), .A2(n41796), .A3(n51950), .ZN(n42111) );
  NAND2_X1 U5447 ( .A1(n41797), .A2(n41792), .ZN(n933) );
  NAND3_X1 U5448 ( .A1(n932), .A2(n41789), .A3(n41790), .ZN(n41808) );
  OAI21_X1 U5450 ( .B1(n933), .B2(n43665), .A(n43666), .ZN(n33883) );
  NAND3_X1 U5452 ( .A1(n42110), .A2(n43665), .A3(n933), .ZN(n42114) );
  NAND2_X1 U5453 ( .A1(n32487), .A2(n32485), .ZN(n32024) );
  NAND4_X1 U5454 ( .A1(n2385), .A2(n32026), .A3(n3664), .A4(n935), .ZN(n32032)
         );
  NAND2_X1 U5455 ( .A1(n32024), .A2(n32491), .ZN(n937) );
  NAND4_X1 U5456 ( .A1(n939), .A2(n946), .A3(n21870), .A4(n938), .ZN(n945) );
  NAND2_X1 U5457 ( .A1(n51858), .A2(n3602), .ZN(n938) );
  NAND2_X1 U5458 ( .A1(n8402), .A2(n23316), .ZN(n21867) );
  NAND3_X1 U5459 ( .A1(n940), .A2(n21871), .A3(n941), .ZN(n944) );
  NAND2_X1 U5460 ( .A1(n943), .A2(n942), .ZN(n940) );
  NAND2_X1 U5461 ( .A1(n23312), .A2(n21874), .ZN(n941) );
  NAND2_X1 U5462 ( .A1(n51125), .A2(n441), .ZN(n21872) );
  NAND3_X1 U5464 ( .A1(n21862), .A2(n23312), .A3(n947), .ZN(n946) );
  AND2_X1 U5465 ( .A1(n23310), .A2(n21863), .ZN(n947) );
  XNOR2_X1 U5466 ( .A(n484), .B(n18689), .ZN(n18564) );
  XNOR2_X1 U5468 ( .A(n18832), .B(n484), .ZN(n15317) );
  XNOR2_X1 U5469 ( .A(n15746), .B(n484), .ZN(n12027) );
  XNOR2_X1 U5470 ( .A(n15004), .B(n484), .ZN(n15889) );
  NAND2_X1 U5471 ( .A1(n24188), .A2(n22605), .ZN(n23761) );
  INV_X2 U5472 ( .A(n23866), .ZN(n24188) );
  AND2_X1 U5473 ( .A1(n21407), .A2(n631), .ZN(n19993) );
  OAI21_X1 U5474 ( .B1(n20780), .B2(n21557), .A(n949), .ZN(n2987) );
  OAI21_X1 U5475 ( .B1(n20782), .B2(n21580), .A(n950), .ZN(n18841) );
  NAND2_X1 U5476 ( .A1(n21407), .A2(n951), .ZN(n950) );
  NAND3_X1 U5477 ( .A1(n952), .A2(n9939), .A3(n10018), .ZN(n9319) );
  NAND2_X1 U5478 ( .A1(n11644), .A2(n11650), .ZN(n952) );
  NAND2_X1 U5479 ( .A1(n952), .A2(n10018), .ZN(n9941) );
  NAND2_X1 U5480 ( .A1(n10015), .A2(n952), .ZN(n10024) );
  NOR2_X1 U5481 ( .A1(n9952), .A2(n803), .ZN(n10043) );
  NAND2_X1 U5482 ( .A1(n954), .A2(n953), .ZN(n9959) );
  NAND2_X1 U5483 ( .A1(n10043), .A2(n9953), .ZN(n953) );
  NAND2_X1 U5484 ( .A1(n9951), .A2(n9953), .ZN(n954) );
  INV_X1 U5485 ( .A(n11841), .ZN(n955) );
  AND3_X1 U5487 ( .A1(n9359), .A2(n12936), .A3(n956), .ZN(n957) );
  NAND4_X1 U5488 ( .A1(n9357), .A2(n13505), .A3(n11841), .A4(n13514), .ZN(n956) );
  INV_X1 U5489 ( .A(n13527), .ZN(n9357) );
  NAND3_X2 U5490 ( .A1(n957), .A2(n961), .A3(n958), .ZN(n17804) );
  NAND2_X1 U5491 ( .A1(n959), .A2(n13515), .ZN(n958) );
  NAND2_X1 U5492 ( .A1(n11843), .A2(n960), .ZN(n959) );
  NAND3_X1 U5493 ( .A1(n963), .A2(n962), .A3(n13500), .ZN(n961) );
  NAND2_X1 U5494 ( .A1(n11843), .A2(n13505), .ZN(n962) );
  NAND2_X1 U5495 ( .A1(n13501), .A2(n11841), .ZN(n11843) );
  NAND2_X1 U5496 ( .A1(n36201), .A2(n36200), .ZN(n39338) );
  INV_X1 U5497 ( .A(n39338), .ZN(n964) );
  NAND2_X1 U5499 ( .A1(n51105), .A2(n29677), .ZN(n31990) );
  NAND2_X1 U5500 ( .A1(n51105), .A2(n32503), .ZN(n31994) );
  AND2_X1 U5501 ( .A1(n31995), .A2(n51105), .ZN(n32001) );
  AOI21_X1 U5503 ( .B1(n24178), .B2(n966), .A(n24180), .ZN(n24199) );
  INV_X1 U5504 ( .A(n4722), .ZN(n966) );
  NAND2_X1 U5505 ( .A1(n21354), .A2(n21605), .ZN(n970) );
  NAND2_X1 U5506 ( .A1(n20768), .A2(n970), .ZN(n19296) );
  NAND2_X1 U5507 ( .A1(n20765), .A2(n968), .ZN(n18720) );
  NAND2_X1 U5508 ( .A1(n762), .A2(n20760), .ZN(n968) );
  NAND2_X1 U5509 ( .A1(n21591), .A2(n970), .ZN(n21593) );
  AOI21_X1 U5510 ( .B1(n21607), .B2(n970), .A(n21362), .ZN(n20762) );
  MUX2_X1 U5511 ( .A(n21352), .B(n21353), .S(n20760), .Z(n21368) );
  NAND2_X1 U5512 ( .A1(n41997), .A2(n971), .ZN(n42000) );
  INV_X1 U5513 ( .A(n42006), .ZN(n971) );
  AND2_X1 U5514 ( .A1(n41997), .A2(n683), .ZN(n4944) );
  NAND2_X1 U5516 ( .A1(n46824), .A2(n51404), .ZN(n46767) );
  NAND2_X1 U5517 ( .A1(n20952), .A2(n22141), .ZN(n974) );
  NAND2_X1 U5518 ( .A1(n21931), .A2(n22154), .ZN(n21019) );
  NOR2_X1 U5519 ( .A1(n28765), .A2(n30732), .ZN(n978) );
  NAND2_X1 U5520 ( .A1(n977), .A2(n976), .ZN(n28777) );
  AOI21_X1 U5521 ( .B1(n28766), .B2(n30732), .A(n742), .ZN(n976) );
  NAND2_X1 U5522 ( .A1(n28765), .A2(n28766), .ZN(n977) );
  NAND2_X1 U5523 ( .A1(n978), .A2(n742), .ZN(n30372) );
  OAI21_X1 U5524 ( .B1(n978), .B2(n30741), .A(n30740), .ZN(n30744) );
  AND2_X1 U5525 ( .A1(n22155), .A2(n979), .ZN(n19560) );
  NOR2_X1 U5526 ( .A1(n50992), .A2(n979), .ZN(n21934) );
  NAND2_X1 U5527 ( .A1(n22154), .A2(n979), .ZN(n21928) );
  NAND3_X1 U5528 ( .A1(n20955), .A2(n20956), .A3(n979), .ZN(n20957) );
  NAND2_X1 U5529 ( .A1(n26877), .A2(n27671), .ZN(n27069) );
  NAND3_X1 U5530 ( .A1(n37381), .A2(n37380), .A3(n983), .ZN(n37383) );
  NAND2_X1 U5531 ( .A1(n17467), .A2(n984), .ZN(n2693) );
  NAND2_X1 U5532 ( .A1(n17466), .A2(n17559), .ZN(n18047) );
  NAND2_X1 U5533 ( .A1(n18039), .A2(n17873), .ZN(n17466) );
  OAI211_X1 U5534 ( .C1(n48469), .C2(n987), .A(n985), .B(n46444), .ZN(n46420)
         );
  INV_X1 U5535 ( .A(n46411), .ZN(n986) );
  INV_X1 U5536 ( .A(n48464), .ZN(n987) );
  NAND2_X1 U5537 ( .A1(n48463), .A2(n48455), .ZN(n48469) );
  AND2_X1 U5538 ( .A1(n46498), .A2(n988), .ZN(n46505) );
  INV_X1 U5540 ( .A(n45188), .ZN(n46746) );
  INV_X1 U5541 ( .A(n41723), .ZN(n45186) );
  NAND3_X1 U5543 ( .A1(n31553), .A2(n31471), .A3(n32614), .ZN(n31554) );
  NAND4_X1 U5544 ( .A1(n32617), .A2(n32614), .A3(n31471), .A4(n32616), .ZN(
        n30324) );
  NAND2_X1 U5545 ( .A1(n23486), .A2(n20994), .ZN(n21341) );
  NAND3_X2 U5546 ( .A1(n6463), .A2(n31834), .A3(n31833), .ZN(n1512) );
  NOR2_X1 U5549 ( .A1(n46396), .A2(n2656), .ZN(n46186) );
  OAI22_X1 U5550 ( .A1(n46396), .A2(n992), .B1(n45218), .B2(n991), .ZN(n45228)
         );
  NAND2_X1 U5551 ( .A1(n46387), .A2(n993), .ZN(n992) );
  INV_X1 U5552 ( .A(n991), .ZN(n993) );
  NAND2_X1 U5553 ( .A1(n653), .A2(n52179), .ZN(n46934) );
  NAND2_X1 U5554 ( .A1(n49036), .A2(n48994), .ZN(n46935) );
  NOR2_X1 U5555 ( .A1(n47435), .A2(n995), .ZN(n994) );
  NOR2_X1 U5557 ( .A1(n30570), .A2(n996), .ZN(n30589) );
  NAND2_X1 U5558 ( .A1(n999), .A2(n997), .ZN(n996) );
  NAND2_X1 U5559 ( .A1(n998), .A2(n31816), .ZN(n997) );
  INV_X1 U5560 ( .A(n30581), .ZN(n998) );
  NAND4_X2 U5563 ( .A1(n44580), .A2(n2286), .A3(n44579), .A4(n46567), .ZN(
        n50708) );
  NAND2_X1 U5564 ( .A1(n1000), .A2(n21756), .ZN(n17513) );
  NAND2_X1 U5565 ( .A1(n23336), .A2(n629), .ZN(n1000) );
  NAND2_X2 U5566 ( .A1(n8160), .A2(n21748), .ZN(n23336) );
  AOI21_X1 U5568 ( .B1(n40638), .B2(n1001), .A(n40637), .ZN(n1146) );
  NAND2_X1 U5569 ( .A1(n42112), .A2(n1001), .ZN(n42113) );
  INV_X1 U5570 ( .A(n38808), .ZN(n1001) );
  NAND2_X1 U5571 ( .A1(n1003), .A2(n33779), .ZN(n33787) );
  NOR2_X1 U5572 ( .A1(n37587), .A2(n37378), .ZN(n1004) );
  NAND2_X1 U5573 ( .A1(n50166), .A2(n1007), .ZN(n50167) );
  NOR2_X1 U5574 ( .A1(n1008), .A2(n50227), .ZN(n1007) );
  NAND2_X1 U5575 ( .A1(n51480), .A2(n50209), .ZN(n1008) );
  NAND2_X1 U5576 ( .A1(n47349), .A2(n49987), .ZN(n1009) );
  NAND2_X1 U5577 ( .A1(n49989), .A2(n1010), .ZN(n47350) );
  AND2_X2 U5578 ( .A1(n49629), .A2(n49627), .ZN(n49989) );
  NOR2_X1 U5579 ( .A1(n38108), .A2(n37420), .ZN(n1011) );
  OR2_X1 U5580 ( .A1(n38118), .A2(n38117), .ZN(n1013) );
  NAND2_X1 U5581 ( .A1(n37417), .A2(n38478), .ZN(n38118) );
  NAND2_X1 U5582 ( .A1(n40916), .A2(n676), .ZN(n1014) );
  NAND3_X1 U5583 ( .A1(n1015), .A2(n26068), .A3(n29448), .ZN(n27041) );
  NOR2_X1 U5584 ( .A1(n27830), .A2(n26039), .ZN(n26071) );
  NAND3_X1 U5585 ( .A1(n38570), .A2(n38201), .A3(n38200), .ZN(n1016) );
  NAND3_X1 U5586 ( .A1(n1016), .A2(n38196), .A3(n38562), .ZN(n38195) );
  NAND2_X1 U5587 ( .A1(n33061), .A2(n1016), .ZN(n33063) );
  XNOR2_X1 U5588 ( .A(n33502), .B(n35586), .ZN(n36691) );
  NAND2_X1 U5589 ( .A1(n1020), .A2(n1017), .ZN(n35586) );
  NAND3_X1 U5590 ( .A1(n1018), .A2(n33419), .A3(n1021), .ZN(n1017) );
  XNOR2_X1 U5591 ( .A(n33764), .B(n36691), .ZN(n32737) );
  INV_X1 U5592 ( .A(n31524), .ZN(n1018) );
  OAI21_X1 U5593 ( .B1(n31524), .B2(n31525), .A(n1019), .ZN(n1020) );
  INV_X1 U5594 ( .A(n33419), .ZN(n1019) );
  INV_X1 U5595 ( .A(n26039), .ZN(n27829) );
  NAND2_X1 U5596 ( .A1(n26723), .A2(n29446), .ZN(n27834) );
  NAND2_X1 U5597 ( .A1(n1022), .A2(n26039), .ZN(n26723) );
  INV_X1 U5598 ( .A(n1023), .ZN(n1022) );
  NAND2_X1 U5599 ( .A1(n29447), .A2(n1023), .ZN(n27025) );
  NAND2_X1 U5600 ( .A1(n27034), .A2(n1023), .ZN(n26065) );
  NAND2_X1 U5601 ( .A1(n21758), .A2(n23336), .ZN(n20865) );
  XNOR2_X1 U5602 ( .A(n7319), .B(n28370), .ZN(n28372) );
  XNOR2_X1 U5603 ( .A(n1025), .B(n7319), .ZN(n20886) );
  XNOR2_X1 U5604 ( .A(n1026), .B(n7319), .ZN(n24850) );
  XNOR2_X1 U5605 ( .A(n7319), .B(n801), .ZN(n25127) );
  XNOR2_X1 U5606 ( .A(n24922), .B(n1027), .ZN(n24923) );
  INV_X1 U5607 ( .A(n26641), .ZN(n1028) );
  NAND2_X1 U5608 ( .A1(n27834), .A2(n430), .ZN(n27032) );
  NAND4_X2 U5609 ( .A1(n5566), .A2(n26648), .A3(n1028), .A4(n1029), .ZN(n31033) );
  NAND3_X1 U5610 ( .A1(n27834), .A2(n1030), .A3(n430), .ZN(n1029) );
  NAND2_X1 U5611 ( .A1(n1031), .A2(n1488), .ZN(n1487) );
  OAI21_X1 U5612 ( .B1(n43443), .B2(n49666), .A(n43442), .ZN(n1031) );
  NAND2_X1 U5613 ( .A1(n6333), .A2(n18040), .ZN(n17557) );
  NAND2_X1 U5615 ( .A1(n45024), .A2(n51395), .ZN(n1032) );
  XNOR2_X1 U5616 ( .A(n1034), .B(n1033), .ZN(n43198) );
  XNOR2_X1 U5617 ( .A(n43195), .B(n1035), .ZN(n1034) );
  NAND2_X1 U5619 ( .A1(n1036), .A2(n34093), .ZN(n8009) );
  NAND2_X1 U5620 ( .A1(n1036), .A2(n5688), .ZN(n3555) );
  NAND2_X1 U5621 ( .A1(n32246), .A2(n32251), .ZN(n24365) );
  NAND2_X1 U5622 ( .A1(n622), .A2(n32251), .ZN(n32237) );
  NAND3_X1 U5623 ( .A1(n32256), .A2(n32257), .A3(n1038), .ZN(n32258) );
  AOI21_X1 U5624 ( .B1(n1040), .B2(n10150), .A(n1039), .ZN(n10154) );
  OAI21_X1 U5625 ( .B1(n1040), .B2(n5047), .A(n8841), .ZN(n8846) );
  NAND2_X1 U5626 ( .A1(n665), .A2(n48481), .ZN(n46458) );
  NAND2_X1 U5627 ( .A1(n1041), .A2(n48252), .ZN(n7665) );
  NAND3_X1 U5628 ( .A1(n48247), .A2(n48479), .A3(n46458), .ZN(n48252) );
  INV_X1 U5629 ( .A(n48254), .ZN(n1041) );
  NAND2_X1 U5630 ( .A1(n37590), .A2(n35980), .ZN(n37588) );
  INV_X1 U5631 ( .A(n2774), .ZN(n30792) );
  INV_X1 U5632 ( .A(n30780), .ZN(n1042) );
  NAND2_X1 U5634 ( .A1(n1043), .A2(n51722), .ZN(n27573) );
  NAND2_X1 U5635 ( .A1(n30793), .A2(n1043), .ZN(n3340) );
  OAI21_X1 U5636 ( .B1(n29906), .B2(n30790), .A(n1043), .ZN(n29912) );
  INV_X1 U5638 ( .A(n39475), .ZN(n1044) );
  OR2_X1 U5639 ( .A1(n7299), .A2(n1046), .ZN(n5584) );
  NAND3_X1 U5640 ( .A1(n10815), .A2(n11608), .A3(n11613), .ZN(n9892) );
  AND2_X1 U5641 ( .A1(n10815), .A2(n11608), .ZN(n9281) );
  NAND2_X1 U5642 ( .A1(n9892), .A2(n11610), .ZN(n9089) );
  NAND2_X1 U5644 ( .A1(n736), .A2(n1048), .ZN(n26940) );
  NAND3_X1 U5645 ( .A1(n26933), .A2(n27665), .A3(n1049), .ZN(n26876) );
  NAND2_X1 U5646 ( .A1(n621), .A2(n31490), .ZN(n5913) );
  NAND2_X1 U5647 ( .A1(n32105), .A2(n32559), .ZN(n32114) );
  INV_X2 U5649 ( .A(n47962), .ZN(n47936) );
  NAND2_X1 U5650 ( .A1(n47966), .A2(n47962), .ZN(n47987) );
  NAND2_X1 U5652 ( .A1(n23995), .A2(n23996), .ZN(n23997) );
  NAND2_X1 U5653 ( .A1(n2008), .A2(n23987), .ZN(n23995) );
  NAND2_X1 U5654 ( .A1(n10924), .A2(n10222), .ZN(n10914) );
  NAND2_X1 U5656 ( .A1(n23153), .A2(n23157), .ZN(n21962) );
  INV_X1 U5657 ( .A(n47426), .ZN(n47427) );
  NAND2_X1 U5658 ( .A1(n49933), .A2(n49923), .ZN(n47426) );
  NAND2_X1 U5659 ( .A1(n30723), .A2(n27588), .ZN(n28800) );
  NAND3_X1 U5661 ( .A1(n36523), .A2(n2916), .A3(n5712), .ZN(n1741) );
  NAND4_X2 U5662 ( .A1(n13020), .A2(n13019), .A3(n14276), .A4(n13021), .ZN(
        n18773) );
  NOR2_X1 U5663 ( .A1(n37626), .A2(n37625), .ZN(n1051) );
  NAND2_X1 U5664 ( .A1(n28560), .A2(n28147), .ZN(n30290) );
  NAND2_X1 U5665 ( .A1(n31466), .A2(n32608), .ZN(n31463) );
  AND2_X1 U5666 ( .A1(n49037), .A2(n653), .ZN(n49034) );
  NOR2_X1 U5668 ( .A1(n23483), .A2(n21975), .ZN(n23486) );
  AOI21_X1 U5672 ( .B1(n1052), .B2(n27161), .A(n27160), .ZN(n27539) );
  NAND2_X1 U5674 ( .A1(n1933), .A2(n47442), .ZN(n47437) );
  NAND2_X1 U5676 ( .A1(n20473), .A2(n1789), .ZN(n20399) );
  NAND2_X1 U5677 ( .A1(n14745), .A2(n20480), .ZN(n1053) );
  AND4_X2 U5680 ( .A1(n8507), .A2(n1938), .A3(n29929), .A4(n1937), .ZN(n1385)
         );
  XNOR2_X1 U5681 ( .A(n1055), .B(n34342), .ZN(n34344) );
  XNOR2_X1 U5682 ( .A(n34343), .B(n34341), .ZN(n1055) );
  XNOR2_X1 U5685 ( .A(n34157), .B(n36873), .ZN(n32811) );
  NAND2_X1 U5686 ( .A1(n1058), .A2(n29198), .ZN(n30622) );
  NAND2_X1 U5687 ( .A1(n27883), .A2(n29205), .ZN(n29198) );
  NOR2_X1 U5688 ( .A1(n1059), .A2(n735), .ZN(n1058) );
  NAND3_X1 U5690 ( .A1(n32097), .A2(n32569), .A3(n32096), .ZN(n32098) );
  NAND4_X4 U5692 ( .A1(n7958), .A2(n18892), .A3(n1060), .A4(n18891), .ZN(
        n23314) );
  NAND2_X1 U5693 ( .A1(n18889), .A2(n18890), .ZN(n1060) );
  NAND2_X1 U5695 ( .A1(n1065), .A2(n326), .ZN(n27748) );
  NAND2_X1 U5696 ( .A1(n27743), .A2(n732), .ZN(n1065) );
  NOR2_X1 U5697 ( .A1(n27006), .A2(n27015), .ZN(n27743) );
  NAND2_X1 U5698 ( .A1(n30434), .A2(n51746), .ZN(n8040) );
  XNOR2_X2 U5699 ( .A(n17906), .B(n3772), .ZN(n17145) );
  NAND2_X1 U5702 ( .A1(n31781), .A2(n32242), .ZN(n29372) );
  NAND2_X2 U5703 ( .A1(n24362), .A2(n24361), .ZN(n31781) );
  NAND3_X1 U5705 ( .A1(n28146), .A2(n28545), .A3(n28560), .ZN(n30301) );
  NOR4_X1 U5706 ( .A1(n31383), .A2(n51740), .A3(n33005), .A4(n31385), .ZN(
        n6421) );
  NAND3_X1 U5707 ( .A1(n41512), .A2(n42019), .A3(n1067), .ZN(n40705) );
  NAND2_X1 U5708 ( .A1(n19059), .A2(n1068), .ZN(n16493) );
  AND2_X1 U5709 ( .A1(n19545), .A2(n20156), .ZN(n1068) );
  NAND2_X1 U5710 ( .A1(n20120), .A2(n20114), .ZN(n19059) );
  NAND2_X1 U5711 ( .A1(n37734), .A2(n37733), .ZN(n37744) );
  NAND3_X1 U5712 ( .A1(n38103), .A2(n38102), .A3(n1069), .ZN(n38106) );
  OAI21_X1 U5713 ( .B1(n31424), .B2(n620), .A(n325), .ZN(n7481) );
  NAND2_X1 U5714 ( .A1(n1071), .A2(n31780), .ZN(n31787) );
  OAI21_X1 U5715 ( .B1(n32253), .B2(n31778), .A(n1072), .ZN(n1071) );
  NAND2_X1 U5717 ( .A1(n9696), .A2(n304), .ZN(n1074) );
  INV_X1 U5718 ( .A(n38972), .ZN(n1075) );
  NAND3_X1 U5719 ( .A1(n1076), .A2(n5958), .A3(n49936), .ZN(n5957) );
  NAND3_X1 U5720 ( .A1(n49920), .A2(n49919), .A3(n1077), .ZN(n1076) );
  NAND3_X1 U5722 ( .A1(n734), .A2(n28757), .A3(n29938), .ZN(n30396) );
  OR2_X1 U5723 ( .A1(n47307), .A2(n49637), .ZN(n49641) );
  NAND3_X1 U5724 ( .A1(n14770), .A2(n15189), .A3(n14771), .ZN(n1079) );
  NAND2_X1 U5725 ( .A1(n7024), .A2(n46756), .ZN(n1080) );
  NAND2_X1 U5727 ( .A1(n24350), .A2(n1081), .ZN(n24356) );
  NAND4_X2 U5728 ( .A1(n1082), .A2(n45855), .A3(n45853), .A4(n45854), .ZN(
        n47651) );
  NAND3_X1 U5729 ( .A1(n45849), .A2(n45848), .A3(n46692), .ZN(n1082) );
  OAI21_X1 U5732 ( .B1(n30170), .B2(n30169), .A(n1084), .ZN(n6083) );
  NAND2_X1 U5733 ( .A1(n30303), .A2(n6084), .ZN(n1084) );
  NOR2_X1 U5734 ( .A1(n5911), .A2(n51357), .ZN(n41009) );
  INV_X1 U5737 ( .A(n37551), .ZN(n1087) );
  INV_X1 U5738 ( .A(n47858), .ZN(n3386) );
  NAND2_X1 U5739 ( .A1(n1626), .A2(n39198), .ZN(n7890) );
  NAND2_X1 U5741 ( .A1(n39378), .A2(n51102), .ZN(n1088) );
  OAI21_X1 U5742 ( .B1(n47671), .B2(n47669), .A(n1089), .ZN(n47654) );
  INV_X1 U5743 ( .A(n11618), .ZN(n1090) );
  INV_X1 U5744 ( .A(n11723), .ZN(n1092) );
  NAND2_X1 U5745 ( .A1(n1093), .A2(n20363), .ZN(n17862) );
  OAI22_X1 U5746 ( .A1(n20430), .A2(n5875), .B1(n20347), .B2(n20360), .ZN(
        n1093) );
  NAND3_X2 U5747 ( .A1(n1094), .A2(n8539), .A3(n37542), .ZN(n41004) );
  NAND2_X1 U5748 ( .A1(n40002), .A2(n40016), .ZN(n35437) );
  OAI211_X1 U5749 ( .C1(n1605), .C2(n2714), .A(n35410), .B(n38332), .ZN(n35411) );
  NAND3_X2 U5751 ( .A1(n1097), .A2(n5764), .A3(n1096), .ZN(n17707) );
  NAND3_X1 U5752 ( .A1(n33035), .A2(n8544), .A3(n30969), .ZN(n1098) );
  NAND2_X1 U5753 ( .A1(n705), .A2(n33026), .ZN(n1099) );
  OAI22_X1 U5754 ( .A1(n48069), .A2(n48068), .B1(n650), .B2(n48070), .ZN(
        n48071) );
  NAND2_X1 U5755 ( .A1(n4031), .A2(n47889), .ZN(n4030) );
  NAND3_X1 U5756 ( .A1(n48211), .A2(n44261), .A3(n1101), .ZN(n44262) );
  NAND3_X2 U5757 ( .A1(n1389), .A2(n1102), .A3(n38378), .ZN(n44006) );
  XNOR2_X1 U5758 ( .A(n1104), .B(n44931), .ZN(n44985) );
  XNOR2_X1 U5759 ( .A(n44930), .B(n44929), .ZN(n1104) );
  XNOR2_X2 U5760 ( .A(n16459), .B(n8700), .ZN(n17018) );
  NAND3_X1 U5761 ( .A1(n27894), .A2(n27822), .A3(n29317), .ZN(n27823) );
  NAND2_X1 U5762 ( .A1(n12250), .A2(n1105), .ZN(n11337) );
  INV_X1 U5763 ( .A(n49344), .ZN(n49305) );
  NAND2_X1 U5764 ( .A1(n49375), .A2(n522), .ZN(n49344) );
  NAND2_X1 U5765 ( .A1(n1107), .A2(n1106), .ZN(n42309) );
  NAND2_X1 U5766 ( .A1(n42304), .A2(n46249), .ZN(n1106) );
  NAND2_X1 U5767 ( .A1(n49162), .A2(n42303), .ZN(n1107) );
  NAND2_X1 U5769 ( .A1(n26775), .A2(n26771), .ZN(n26813) );
  NAND4_X2 U5770 ( .A1(n22372), .A2(n7192), .A3(n22366), .A4(n1109), .ZN(
        n25501) );
  NAND4_X1 U5771 ( .A1(n22353), .A2(n22352), .A3(n22350), .A4(n22351), .ZN(
        n1109) );
  XNOR2_X1 U5772 ( .A(n15514), .B(n15513), .ZN(n1110) );
  NAND2_X1 U5774 ( .A1(n14071), .A2(n1111), .ZN(n14077) );
  NAND2_X1 U5775 ( .A1(n11296), .A2(n14397), .ZN(n14071) );
  NAND3_X1 U5776 ( .A1(n1112), .A2(n20578), .A3(n20577), .ZN(n20583) );
  NAND2_X1 U5777 ( .A1(n3286), .A2(n3288), .ZN(n1112) );
  INV_X1 U5778 ( .A(n7287), .ZN(n36533) );
  INV_X1 U5779 ( .A(n1484), .ZN(n8481) );
  XNOR2_X1 U5780 ( .A(n33235), .B(n32338), .ZN(n1113) );
  NAND3_X1 U5781 ( .A1(n4209), .A2(n5411), .A3(n13574), .ZN(n13579) );
  MUX2_X1 U5782 ( .A(n20818), .B(n20819), .S(n21492), .Z(n20834) );
  NAND2_X1 U5784 ( .A1(n1114), .A2(n8804), .ZN(n8805) );
  NAND2_X1 U5785 ( .A1(n10963), .A2(n2865), .ZN(n1114) );
  NAND2_X1 U5786 ( .A1(n31726), .A2(n1115), .ZN(n31727) );
  AND3_X1 U5787 ( .A1(n7682), .A2(n26741), .A3(n7681), .ZN(n4728) );
  INV_X1 U5788 ( .A(n50721), .ZN(n1467) );
  XNOR2_X1 U5789 ( .A(n1116), .B(n8751), .ZN(n34612) );
  XNOR2_X1 U5790 ( .A(n34610), .B(n34607), .ZN(n1116) );
  XNOR2_X1 U5791 ( .A(n1117), .B(n8087), .ZN(n34606) );
  NAND3_X1 U5792 ( .A1(n17560), .A2(n17558), .A3(n17559), .ZN(n17561) );
  NAND3_X2 U5793 ( .A1(n1119), .A2(n37934), .A3(n1118), .ZN(n41539) );
  INV_X1 U5794 ( .A(n37938), .ZN(n1118) );
  NAND2_X1 U5795 ( .A1(n1122), .A2(n1121), .ZN(n1120) );
  OAI211_X1 U5796 ( .C1(n28765), .C2(n7410), .A(n30742), .B(n27380), .ZN(n1122) );
  XNOR2_X2 U5798 ( .A(n1124), .B(n44491), .ZN(n46872) );
  XNOR2_X1 U5799 ( .A(n44480), .B(n44481), .ZN(n1124) );
  NAND2_X1 U5800 ( .A1(n37462), .A2(n40767), .ZN(n1125) );
  NAND2_X1 U5801 ( .A1(n40787), .A2(n40073), .ZN(n1126) );
  NAND2_X1 U5804 ( .A1(n1128), .A2(n9017), .ZN(n9018) );
  OAI21_X1 U5805 ( .B1(n9016), .B2(n9704), .A(n10726), .ZN(n1128) );
  NAND4_X1 U5806 ( .A1(n1129), .A2(n29585), .A3(n31125), .A4(n30066), .ZN(
        n7427) );
  OAI21_X1 U5807 ( .B1(n41590), .B2(n41589), .A(n1132), .ZN(n8673) );
  NAND2_X1 U5808 ( .A1(n41589), .A2(n1133), .ZN(n1132) );
  XNOR2_X1 U5809 ( .A(n1134), .B(n45612), .ZN(Plaintext[43]) );
  NOR2_X1 U5813 ( .A1(n19642), .A2(n1135), .ZN(n18254) );
  NAND2_X1 U5814 ( .A1(n19643), .A2(n19033), .ZN(n1135) );
  NAND2_X1 U5815 ( .A1(n1751), .A2(n1754), .ZN(n48187) );
  NAND2_X1 U5816 ( .A1(n48180), .A2(n668), .ZN(n48165) );
  NAND2_X1 U5817 ( .A1(n8686), .A2(n48498), .ZN(n8684) );
  NAND2_X1 U5818 ( .A1(n30758), .A2(n29924), .ZN(n30772) );
  OR2_X2 U5819 ( .A1(n1136), .A2(n27718), .ZN(n30912) );
  NAND2_X1 U5820 ( .A1(n14345), .A2(n14339), .ZN(n12228) );
  NAND2_X1 U5821 ( .A1(n10926), .A2(n10925), .ZN(n1137) );
  XNOR2_X1 U5825 ( .A(n8623), .B(n8622), .ZN(n1138) );
  NAND3_X2 U5828 ( .A1(n1139), .A2(n4309), .A3(n14357), .ZN(n17208) );
  NAND3_X1 U5829 ( .A1(n13010), .A2(n13009), .A3(n4311), .ZN(n1139) );
  NAND2_X1 U5832 ( .A1(n1142), .A2(n1141), .ZN(n37908) );
  NAND2_X1 U5833 ( .A1(n2507), .A2(n39428), .ZN(n1141) );
  NAND2_X1 U5834 ( .A1(n1143), .A2(n39204), .ZN(n1142) );
  NAND3_X1 U5836 ( .A1(n7393), .A2(n7394), .A3(n31550), .ZN(n7395) );
  NAND2_X1 U5837 ( .A1(n36087), .A2(n37977), .ZN(n1144) );
  NAND2_X1 U5838 ( .A1(n36080), .A2(n36353), .ZN(n36087) );
  NAND2_X1 U5839 ( .A1(n40640), .A2(n40639), .ZN(n1147) );
  NAND3_X1 U5841 ( .A1(n28146), .A2(n30289), .A3(n27111), .ZN(n30299) );
  NAND2_X1 U5843 ( .A1(n6541), .A2(n38015), .ZN(n38184) );
  OAI211_X1 U5846 ( .C1(n610), .C2(n39603), .A(n40506), .B(n1667), .ZN(n1668)
         );
  NAND3_X1 U5847 ( .A1(n51355), .A2(n413), .A3(n23223), .ZN(n22118) );
  NAND3_X1 U5849 ( .A1(n48178), .A2(n48421), .A3(n48409), .ZN(n48183) );
  AOI21_X1 U5850 ( .B1(n3096), .B2(n32137), .A(n32136), .ZN(n1150) );
  NAND2_X1 U5851 ( .A1(n1151), .A2(n50553), .ZN(n50540) );
  OAI21_X1 U5855 ( .B1(n41696), .B2(n41695), .A(n333), .ZN(n41701) );
  OAI211_X1 U5856 ( .C1(n30306), .C2(n2201), .A(n30307), .B(n1152), .ZN(n27089) );
  NAND2_X1 U5857 ( .A1(n30306), .A2(n29140), .ZN(n1152) );
  XNOR2_X1 U5858 ( .A(n43522), .B(n51444), .ZN(n41192) );
  NAND2_X1 U5859 ( .A1(n46510), .A2(n46336), .ZN(n48412) );
  XNOR2_X1 U5860 ( .A(n34275), .B(n33609), .ZN(n33610) );
  XNOR2_X2 U5861 ( .A(n34869), .B(n35331), .ZN(n34275) );
  XOR2_X1 U5862 ( .A(n25152), .B(n2209), .Z(n1278) );
  OR2_X1 U5863 ( .A1(n1789), .A2(n20468), .ZN(n19378) );
  AND2_X1 U5864 ( .A1(n2007), .A2(n2006), .ZN(n2005) );
  XNOR2_X1 U5866 ( .A(n17930), .B(n17929), .ZN(n20795) );
  NAND2_X1 U5867 ( .A1(n10832), .A2(n12521), .ZN(n11260) );
  INV_X1 U5868 ( .A(n12964), .ZN(n1317) );
  NAND3_X1 U5869 ( .A1(n32862), .A2(n32870), .A3(n32883), .ZN(n32863) );
  XNOR2_X2 U5870 ( .A(n46050), .B(n43920), .ZN(n45303) );
  NAND2_X1 U5871 ( .A1(n1155), .A2(n49070), .ZN(n49128) );
  NAND4_X2 U5872 ( .A1(n44738), .A2(n44739), .A3(n44736), .A4(n44737), .ZN(
        n49119) );
  NAND2_X1 U5873 ( .A1(n45937), .A2(n49137), .ZN(n44733) );
  NAND3_X1 U5874 ( .A1(n7134), .A2(n20866), .A3(n20867), .ZN(n7133) );
  NAND2_X1 U5875 ( .A1(n11943), .A2(n11108), .ZN(n11955) );
  NAND2_X1 U5876 ( .A1(n29198), .A2(n1156), .ZN(n29209) );
  NAND2_X1 U5877 ( .A1(n18374), .A2(n6711), .ZN(n1157) );
  NAND3_X1 U5880 ( .A1(n1158), .A2(n31346), .A3(n51744), .ZN(n30047) );
  NAND3_X1 U5881 ( .A1(n37598), .A2(n37597), .A3(n37593), .ZN(n37375) );
  INV_X1 U5882 ( .A(n30098), .ZN(n30992) );
  OAI21_X1 U5883 ( .B1(n5937), .B2(n1161), .A(n1160), .ZN(n44725) );
  NAND2_X1 U5884 ( .A1(n44724), .A2(n49150), .ZN(n1160) );
  INV_X1 U5885 ( .A(n20555), .ZN(n22641) );
  NAND2_X1 U5886 ( .A1(n17420), .A2(n22639), .ZN(n20555) );
  INV_X1 U5887 ( .A(n27511), .ZN(n1376) );
  NAND4_X1 U5888 ( .A1(n45716), .A2(n8163), .A3(n45710), .A4(n8164), .ZN(
        n45718) );
  AOI21_X1 U5889 ( .B1(n8023), .B2(n51709), .A(n5845), .ZN(n8025) );
  NAND2_X1 U5890 ( .A1(n6853), .A2(n30182), .ZN(n26468) );
  NAND2_X1 U5891 ( .A1(n41112), .A2(n41268), .ZN(n41257) );
  AND2_X2 U5892 ( .A1(n2224), .A2(n3655), .ZN(n40893) );
  NAND2_X1 U5894 ( .A1(n32396), .A2(n32407), .ZN(n31280) );
  NAND2_X1 U5895 ( .A1(n40420), .A2(n52193), .ZN(n41287) );
  OR2_X1 U5896 ( .A1(n17627), .A2(n20507), .ZN(n18077) );
  NAND3_X1 U5897 ( .A1(n23913), .A2(n6207), .A3(n23924), .ZN(n4349) );
  NAND2_X1 U5899 ( .A1(n32878), .A2(n1164), .ZN(n32880) );
  NAND2_X1 U5900 ( .A1(n705), .A2(n719), .ZN(n1164) );
  INV_X2 U5901 ( .A(n25421), .ZN(n25107) );
  NAND3_X1 U5902 ( .A1(n6786), .A2(n11354), .A3(n51138), .ZN(n10683) );
  NAND3_X1 U5903 ( .A1(n3372), .A2(n38354), .A3(n1165), .ZN(n38360) );
  NAND3_X1 U5904 ( .A1(n27130), .A2(n28894), .A3(n27129), .ZN(n28890) );
  NAND2_X1 U5906 ( .A1(n19680), .A2(n16994), .ZN(n20220) );
  NOR2_X1 U5908 ( .A1(n2531), .A2(n1166), .ZN(n5001) );
  NAND2_X1 U5909 ( .A1(n3347), .A2(n12617), .ZN(n1167) );
  NAND2_X1 U5912 ( .A1(n30772), .A2(n29917), .ZN(n3201) );
  NAND2_X1 U5914 ( .A1(n1238), .A2(n13467), .ZN(n13468) );
  XNOR2_X2 U5915 ( .A(n1171), .B(n24734), .ZN(n27668) );
  XNOR2_X1 U5916 ( .A(n24731), .B(n24730), .ZN(n1171) );
  NAND2_X1 U5919 ( .A1(n1173), .A2(n22826), .ZN(n21065) );
  OAI21_X1 U5920 ( .B1(n22830), .B2(n22832), .A(n288), .ZN(n1173) );
  NAND2_X1 U5921 ( .A1(n41900), .A2(n40724), .ZN(n5128) );
  NOR2_X1 U5922 ( .A1(n46872), .A2(n47096), .ZN(n47089) );
  AOI21_X1 U5924 ( .B1(n1201), .B2(n46570), .A(n1199), .ZN(n44580) );
  NAND3_X1 U5925 ( .A1(n20760), .A2(n20759), .A3(n21361), .ZN(n20761) );
  XNOR2_X1 U5926 ( .A(n43937), .B(n42763), .ZN(n1174) );
  OAI21_X1 U5929 ( .B1(n9862), .B2(n9793), .A(n10960), .ZN(n5328) );
  NAND3_X1 U5930 ( .A1(n49043), .A2(n49016), .A3(n51321), .ZN(n1175) );
  NAND2_X1 U5931 ( .A1(n51310), .A2(n49018), .ZN(n1176) );
  OR2_X1 U5932 ( .A1(n40917), .A2(n1633), .ZN(n40954) );
  INV_X1 U5933 ( .A(n22623), .ZN(n23637) );
  XNOR2_X1 U5934 ( .A(n43645), .B(n43646), .ZN(n7777) );
  NAND4_X1 U5935 ( .A1(n2023), .A2(n13494), .A3(n13477), .A4(n13478), .ZN(
        n2022) );
  NAND3_X1 U5938 ( .A1(n46449), .A2(n8585), .A3(n46441), .ZN(n48470) );
  NAND2_X1 U5939 ( .A1(n12045), .A2(n11387), .ZN(n10364) );
  XNOR2_X2 U5941 ( .A(n15457), .B(n15456), .ZN(n18041) );
  INV_X1 U5942 ( .A(n47588), .ZN(n47257) );
  NAND2_X1 U5943 ( .A1(n23417), .A2(n1177), .ZN(n20162) );
  NAND2_X1 U5944 ( .A1(n39990), .A2(n1178), .ZN(n4016) );
  NOR2_X1 U5945 ( .A1(n345), .A2(n1179), .ZN(n47799) );
  OAI21_X1 U5946 ( .B1(n47796), .B2(n45876), .A(n47794), .ZN(n1179) );
  NAND2_X1 U5947 ( .A1(n7474), .A2(n27040), .ZN(n27836) );
  NAND2_X1 U5948 ( .A1(n27838), .A2(n27837), .ZN(n1180) );
  NAND4_X1 U5949 ( .A1(n32586), .A2(n1182), .A3(n32587), .A4(n1181), .ZN(n7487) );
  INV_X1 U5950 ( .A(n32975), .ZN(n1182) );
  INV_X1 U5951 ( .A(n24272), .ZN(n1687) );
  NAND3_X1 U5953 ( .A1(n12397), .A2(n12396), .A3(n313), .ZN(n12398) );
  NAND2_X1 U5954 ( .A1(n39703), .A2(n39713), .ZN(n1183) );
  NAND2_X1 U5956 ( .A1(n3798), .A2(n47831), .ZN(n47825) );
  NAND2_X1 U5957 ( .A1(n3797), .A2(n47858), .ZN(n42193) );
  NAND3_X1 U5958 ( .A1(n7185), .A2(n11641), .A3(n11639), .ZN(n11642) );
  INV_X1 U5960 ( .A(n30635), .ZN(n5669) );
  NAND2_X1 U5961 ( .A1(n711), .A2(n31740), .ZN(n30635) );
  NAND2_X1 U5962 ( .A1(n1184), .A2(n13781), .ZN(n1910) );
  NAND2_X1 U5963 ( .A1(n12416), .A2(n10905), .ZN(n1184) );
  NAND2_X1 U5964 ( .A1(n13782), .A2(n12419), .ZN(n12416) );
  NAND4_X2 U5966 ( .A1(n6598), .A2(n2251), .A3(n34657), .A4(n34658), .ZN(
        n41083) );
  OAI211_X1 U5968 ( .C1(n39906), .C2(n39785), .A(n38449), .B(n39910), .ZN(
        n38453) );
  NAND3_X1 U5969 ( .A1(n30764), .A2(n30773), .A3(n30763), .ZN(n1322) );
  NAND2_X1 U5970 ( .A1(n1188), .A2(n1186), .ZN(n47603) );
  NAND2_X1 U5971 ( .A1(n47594), .A2(n1187), .ZN(n1186) );
  NAND2_X1 U5972 ( .A1(n52158), .A2(n47593), .ZN(n1188) );
  NAND2_X1 U5973 ( .A1(n50466), .A2(n1190), .ZN(n1189) );
  NAND2_X1 U5974 ( .A1(n50717), .A2(n4039), .ZN(n50720) );
  AND2_X2 U5975 ( .A1(n10959), .A2(n10127), .ZN(n10962) );
  OAI211_X1 U5978 ( .C1(n34637), .C2(n34638), .A(n34635), .B(n34636), .ZN(
        n1191) );
  NAND3_X1 U5979 ( .A1(n21564), .A2(n1192), .A3(n21563), .ZN(n20784) );
  NAND2_X1 U5980 ( .A1(n21556), .A2(n5192), .ZN(n1192) );
  NAND3_X1 U5983 ( .A1(n24103), .A2(n24104), .A3(n24109), .ZN(n1193) );
  NAND3_X1 U5984 ( .A1(n38334), .A2(n38330), .A3(n38345), .ZN(n37663) );
  AND2_X1 U5988 ( .A1(n32491), .A2(n32486), .ZN(n31203) );
  NAND3_X1 U5992 ( .A1(n38901), .A2(n38899), .A3(n41380), .ZN(n38886) );
  NAND2_X1 U5994 ( .A1(n13257), .A2(n13258), .ZN(n1195) );
  NAND3_X1 U5995 ( .A1(n10357), .A2(n10358), .A3(n10359), .ZN(n3356) );
  INV_X1 U5996 ( .A(n2699), .ZN(n5865) );
  XOR2_X1 U5997 ( .A(n27476), .B(n27475), .Z(n1239) );
  NAND4_X1 U5998 ( .A1(n48813), .A2(n48810), .A3(n48812), .A4(n48811), .ZN(
        n4301) );
  NAND4_X2 U5999 ( .A1(n42166), .A2(n42163), .A3(n42164), .A4(n42165), .ZN(
        n45421) );
  INV_X1 U6000 ( .A(n1404), .ZN(n1917) );
  NAND2_X1 U6001 ( .A1(n1197), .A2(n4051), .ZN(n4050) );
  NAND2_X1 U6002 ( .A1(n21061), .A2(n1198), .ZN(n1197) );
  NAND3_X1 U6003 ( .A1(n37985), .A2(n36351), .A3(n37977), .ZN(n7287) );
  OR2_X2 U6005 ( .A1(n12103), .A2(n12104), .ZN(n14370) );
  NAND3_X2 U6006 ( .A1(n3405), .A2(n3406), .A3(n9630), .ZN(n17125) );
  OAI21_X1 U6007 ( .B1(n44642), .B2(n44641), .A(n1720), .ZN(n1719) );
  INV_X1 U6008 ( .A(n13729), .ZN(n14032) );
  XNOR2_X1 U6009 ( .A(n1200), .B(n43258), .ZN(n43260) );
  XNOR2_X1 U6010 ( .A(n45361), .B(n43257), .ZN(n1200) );
  NAND2_X1 U6011 ( .A1(n39240), .A2(n51508), .ZN(n38702) );
  NAND2_X1 U6012 ( .A1(n5275), .A2(n47109), .ZN(n1201) );
  NAND4_X4 U6013 ( .A1(n1623), .A2(n1624), .A3(n1625), .A4(n5815), .ZN(n49606)
         );
  NAND2_X1 U6014 ( .A1(n5976), .A2(n32909), .ZN(n5975) );
  NAND2_X1 U6015 ( .A1(n32896), .A2(n32917), .ZN(n28823) );
  NAND2_X1 U6016 ( .A1(n32540), .A2(n32908), .ZN(n32896) );
  NAND2_X1 U6017 ( .A1(n12891), .A2(n12792), .ZN(n9991) );
  NAND3_X1 U6020 ( .A1(n32524), .A2(n32763), .A3(n32961), .ZN(n8389) );
  NAND2_X1 U6021 ( .A1(n41481), .A2(n42061), .ZN(n40288) );
  NAND2_X1 U6022 ( .A1(n1348), .A2(n2367), .ZN(n28756) );
  XNOR2_X1 U6023 ( .A(n35496), .B(n1203), .ZN(n33829) );
  XNOR2_X1 U6024 ( .A(n33826), .B(n33827), .ZN(n1203) );
  NAND2_X1 U6025 ( .A1(n17313), .A2(n2879), .ZN(n1481) );
  XNOR2_X2 U6026 ( .A(n36748), .B(n35105), .ZN(n35296) );
  NAND2_X1 U6027 ( .A1(n1204), .A2(n19113), .ZN(n5625) );
  NAND3_X1 U6028 ( .A1(n4791), .A2(n19111), .A3(n21223), .ZN(n1204) );
  NAND2_X1 U6029 ( .A1(n1205), .A2(n14876), .ZN(n4707) );
  NAND3_X1 U6030 ( .A1(n7795), .A2(n7796), .A3(n42993), .ZN(n7794) );
  NAND3_X1 U6033 ( .A1(n36206), .A2(n39472), .A3(n36205), .ZN(n4095) );
  OAI21_X1 U6034 ( .B1(n48431), .B2(n48443), .A(n1645), .ZN(n48446) );
  NAND2_X1 U6036 ( .A1(n21613), .A2(n21620), .ZN(n16000) );
  NAND3_X1 U6037 ( .A1(n8586), .A2(n22830), .A3(n20298), .ZN(n21066) );
  INV_X1 U6039 ( .A(n11177), .ZN(n1844) );
  NAND2_X1 U6040 ( .A1(n1209), .A2(n1208), .ZN(n10108) );
  NAND2_X1 U6041 ( .A1(n10513), .A2(n1210), .ZN(n1209) );
  INV_X1 U6042 ( .A(n10529), .ZN(n1210) );
  NAND2_X1 U6043 ( .A1(n1211), .A2(n6535), .ZN(n6533) );
  NAND2_X1 U6044 ( .A1(n6534), .A2(n40377), .ZN(n1211) );
  NAND2_X1 U6045 ( .A1(n48759), .A2(n48722), .ZN(n47452) );
  NAND2_X1 U6046 ( .A1(n1212), .A2(n48403), .ZN(n46339) );
  NAND2_X1 U6047 ( .A1(n48410), .A2(n8057), .ZN(n1212) );
  NAND3_X1 U6048 ( .A1(n47207), .A2(n47591), .A3(n47586), .ZN(n47209) );
  NAND2_X1 U6049 ( .A1(n25395), .A2(n30216), .ZN(n25394) );
  NAND2_X1 U6050 ( .A1(n3130), .A2(n3128), .ZN(n40063) );
  NAND2_X2 U6051 ( .A1(n1213), .A2(n4664), .ZN(n31466) );
  NAND3_X1 U6053 ( .A1(n30298), .A2(n30300), .A3(n30297), .ZN(n1215) );
  NAND2_X1 U6054 ( .A1(n1464), .A2(n41482), .ZN(n5673) );
  NAND2_X1 U6055 ( .A1(n47596), .A2(n47586), .ZN(n47619) );
  NAND2_X1 U6057 ( .A1(n48551), .A2(n48234), .ZN(n48538) );
  XNOR2_X2 U6059 ( .A(n37081), .B(n7787), .ZN(n34446) );
  XNOR2_X1 U6060 ( .A(n1217), .B(n25331), .ZN(n25335) );
  XNOR2_X1 U6061 ( .A(n25324), .B(n25323), .ZN(n1217) );
  NAND3_X1 U6063 ( .A1(n14657), .A2(n786), .A3(n13434), .ZN(n13993) );
  AND3_X1 U6064 ( .A1(n14649), .A2(n14646), .A3(n14648), .ZN(n1219) );
  XNOR2_X2 U6065 ( .A(n43249), .B(n8495), .ZN(n49657) );
  NAND2_X1 U6067 ( .A1(n21970), .A2(n21979), .ZN(n21978) );
  NAND2_X1 U6068 ( .A1(n1221), .A2(n7823), .ZN(n4372) );
  OAI22_X1 U6069 ( .A1(n10233), .A2(n10232), .B1(n10231), .B2(n12277), .ZN(
        n1221) );
  NAND2_X1 U6070 ( .A1(n28626), .A2(n26973), .ZN(n4075) );
  NAND2_X1 U6071 ( .A1(n2227), .A2(n796), .ZN(n10346) );
  NAND2_X1 U6073 ( .A1(n3538), .A2(n1223), .ZN(n3537) );
  NAND2_X1 U6076 ( .A1(n17471), .A2(n1227), .ZN(n17472) );
  NAND2_X1 U6077 ( .A1(n19411), .A2(n19413), .ZN(n17471) );
  NAND2_X1 U6078 ( .A1(n1229), .A2(n1228), .ZN(n4684) );
  NAND2_X1 U6079 ( .A1(n30811), .A2(n31708), .ZN(n1228) );
  NAND2_X1 U6080 ( .A1(n32122), .A2(n26350), .ZN(n1229) );
  INV_X1 U6081 ( .A(n23993), .ZN(n23991) );
  INV_X1 U6083 ( .A(n22531), .ZN(n1230) );
  NAND3_X1 U6085 ( .A1(n30419), .A2(n28793), .A3(n28971), .ZN(n28979) );
  NAND2_X1 U6086 ( .A1(n30296), .A2(n30283), .ZN(n28147) );
  OR2_X1 U6087 ( .A1(n29158), .A2(n2889), .ZN(n29160) );
  NAND3_X1 U6089 ( .A1(n37551), .A2(n37562), .A3(n37561), .ZN(n37556) );
  NAND2_X1 U6090 ( .A1(n51352), .A2(n40119), .ZN(n36094) );
  NAND3_X2 U6091 ( .A1(n4034), .A2(n36090), .A3(n36091), .ZN(n40119) );
  NAND2_X1 U6092 ( .A1(n37383), .A2(n37382), .ZN(n40060) );
  NAND2_X1 U6093 ( .A1(n39632), .A2(n41355), .ZN(n38747) );
  NAND2_X1 U6094 ( .A1(n2065), .A2(n40824), .ZN(n39514) );
  XNOR2_X2 U6095 ( .A(n1232), .B(n16576), .ZN(n20266) );
  NAND2_X1 U6096 ( .A1(n27555), .A2(n30763), .ZN(n30753) );
  AND2_X1 U6098 ( .A1(n46763), .A2(n46762), .ZN(n1233) );
  NAND2_X1 U6099 ( .A1(n3703), .A2(n32345), .ZN(n32452) );
  INV_X1 U6100 ( .A(n37468), .ZN(n37469) );
  NAND2_X1 U6101 ( .A1(n4000), .A2(n40558), .ZN(n37468) );
  NAND2_X1 U6102 ( .A1(n1234), .A2(n2444), .ZN(n6166) );
  NAND2_X1 U6103 ( .A1(n21529), .A2(n6163), .ZN(n1234) );
  NAND2_X1 U6104 ( .A1(n1235), .A2(n46863), .ZN(n46680) );
  INV_X1 U6105 ( .A(n5360), .ZN(n1235) );
  NAND2_X1 U6106 ( .A1(n47121), .A2(n46654), .ZN(n5360) );
  OAI21_X1 U6109 ( .B1(n13464), .B2(n13465), .A(n13463), .ZN(n1238) );
  OR2_X1 U6110 ( .A1(n41004), .A2(n38764), .ZN(n38759) );
  NAND3_X1 U6111 ( .A1(n49626), .A2(n49623), .A3(n43455), .ZN(n4009) );
  XNOR2_X1 U6112 ( .A(n28230), .B(n1239), .ZN(n2255) );
  XNOR2_X1 U6114 ( .A(n1240), .B(n42375), .ZN(n42379) );
  XNOR2_X1 U6115 ( .A(n44040), .B(n42788), .ZN(n1240) );
  NAND2_X1 U6116 ( .A1(n36535), .A2(n36081), .ZN(n36082) );
  OR2_X2 U6117 ( .A1(n7242), .A2(n3202), .ZN(n35237) );
  NOR2_X1 U6118 ( .A1(n1242), .A2(n341), .ZN(n50076) );
  OAI21_X1 U6119 ( .B1(n50061), .B2(n50120), .A(n50060), .ZN(n1242) );
  BUF_X1 U6120 ( .A(n41308), .Z(n46111) );
  NAND3_X2 U6121 ( .A1(n1243), .A2(n1539), .A3(n1534), .ZN(n22491) );
  NAND2_X1 U6122 ( .A1(n1244), .A2(n13088), .ZN(n12821) );
  OR2_X2 U6123 ( .A1(n9478), .A2(n9479), .ZN(n13088) );
  INV_X1 U6124 ( .A(n1929), .ZN(n13084) );
  AOI22_X1 U6125 ( .A1(n1245), .A2(n47831), .B1(n47817), .B2(n42191), .ZN(
        n42198) );
  NAND2_X1 U6126 ( .A1(n47849), .A2(n3385), .ZN(n1245) );
  NAND3_X1 U6127 ( .A1(n1246), .A2(n23573), .A3(n23574), .ZN(n23575) );
  NAND2_X1 U6129 ( .A1(n18217), .A2(n21300), .ZN(n18991) );
  NAND2_X1 U6130 ( .A1(n5389), .A2(n30346), .ZN(n29060) );
  OAI211_X1 U6132 ( .C1(n11757), .C2(n12898), .A(n1448), .B(n1447), .ZN(n4959)
         );
  AND2_X1 U6134 ( .A1(n29118), .A2(n3154), .ZN(n1429) );
  NAND3_X1 U6135 ( .A1(n45190), .A2(n46743), .A3(n46756), .ZN(n45191) );
  NOR2_X1 U6136 ( .A1(n31358), .A2(n36299), .ZN(n38213) );
  OAI21_X1 U6137 ( .B1(n47011), .B2(n50039), .A(n47020), .ZN(n8529) );
  NAND3_X1 U6138 ( .A1(n49441), .A2(n49424), .A3(n49440), .ZN(n47204) );
  NAND3_X1 U6139 ( .A1(n45681), .A2(n45930), .A3(n49275), .ZN(n45666) );
  XNOR2_X2 U6140 ( .A(n1248), .B(n37287), .ZN(n38704) );
  XNOR2_X1 U6141 ( .A(n37298), .B(n37286), .ZN(n1248) );
  NAND2_X1 U6142 ( .A1(n32895), .A2(n5111), .ZN(n32911) );
  NAND2_X1 U6143 ( .A1(n39225), .A2(n39235), .ZN(n37916) );
  OAI21_X1 U6144 ( .B1(n41555), .B2(n41556), .A(n41554), .ZN(n41557) );
  NAND2_X1 U6145 ( .A1(n3553), .A2(n21775), .ZN(n21120) );
  NAND2_X1 U6147 ( .A1(n1789), .A2(n20472), .ZN(n20475) );
  NAND2_X1 U6148 ( .A1(n1250), .A2(n1249), .ZN(n49260) );
  NAND2_X1 U6149 ( .A1(n49240), .A2(n656), .ZN(n1249) );
  NAND2_X1 U6150 ( .A1(n1252), .A2(n1251), .ZN(n1250) );
  NAND2_X1 U6154 ( .A1(n36901), .A2(n39464), .ZN(n39452) );
  NAND2_X1 U6155 ( .A1(n51478), .A2(n47481), .ZN(n1255) );
  NAND3_X1 U6156 ( .A1(n42804), .A2(n48958), .A3(n51511), .ZN(n1256) );
  NAND3_X1 U6157 ( .A1(n9144), .A2(n11199), .A3(n11711), .ZN(n9143) );
  NAND2_X1 U6158 ( .A1(n11696), .A2(n11209), .ZN(n9144) );
  NAND3_X2 U6159 ( .A1(n1258), .A2(n6650), .A3(n4185), .ZN(n22129) );
  AND2_X1 U6160 ( .A1(n8266), .A2(n19051), .ZN(n1258) );
  AOI21_X1 U6161 ( .B1(n19151), .B2(n19150), .A(n1775), .ZN(n19154) );
  INV_X1 U6163 ( .A(n20060), .ZN(n19494) );
  NAND2_X1 U6164 ( .A1(n16217), .A2(n20052), .ZN(n20060) );
  XNOR2_X1 U6165 ( .A(n4767), .B(n335), .ZN(n1466) );
  NAND3_X1 U6166 ( .A1(n47826), .A2(n47825), .A3(n4397), .ZN(n1263) );
  NAND3_X1 U6167 ( .A1(n38841), .A2(n6372), .A3(n6373), .ZN(n6371) );
  NAND3_X1 U6168 ( .A1(n26778), .A2(n26825), .A3(n26777), .ZN(n7786) );
  AND2_X1 U6169 ( .A1(n23606), .A2(n24211), .ZN(n22638) );
  INV_X1 U6170 ( .A(n44270), .ZN(n1259) );
  NOR2_X1 U6172 ( .A1(n24213), .A2(n3929), .ZN(n25464) );
  AND4_X2 U6173 ( .A1(n46926), .A2(n46923), .A3(n46925), .A4(n46924), .ZN(
        n1441) );
  NAND2_X1 U6174 ( .A1(n36242), .A2(n37763), .ZN(n35914) );
  NAND3_X1 U6175 ( .A1(n37764), .A2(n36247), .A3(n37753), .ZN(n37763) );
  NAND2_X1 U6176 ( .A1(n48411), .A2(n48408), .ZN(n45499) );
  NAND4_X4 U6177 ( .A1(n6223), .A2(n6221), .A3(n6222), .A4(n35922), .ZN(n42201) );
  NAND3_X1 U6179 ( .A1(n1260), .A2(n38757), .A3(n38758), .ZN(n38768) );
  OAI21_X1 U6180 ( .B1(n38755), .B2(n38754), .A(n1261), .ZN(n1260) );
  NAND2_X1 U6181 ( .A1(n14406), .A2(n12961), .ZN(n11294) );
  NAND2_X1 U6182 ( .A1(n14068), .A2(n12869), .ZN(n14406) );
  OAI21_X1 U6183 ( .B1(n16001), .B2(n20700), .A(n20253), .ZN(n1262) );
  NAND3_X2 U6184 ( .A1(n20599), .A2(n20598), .A3(n20597), .ZN(n26565) );
  NAND4_X1 U6185 ( .A1(n13488), .A2(n13489), .A3(n13490), .A4(n13491), .ZN(
        n2021) );
  NAND4_X1 U6186 ( .A1(n1263), .A2(n47833), .A3(n47832), .A4(n47834), .ZN(
        n47835) );
  OR2_X2 U6187 ( .A1(n26633), .A2(n26632), .ZN(n33005) );
  OAI211_X1 U6188 ( .C1(n36489), .C2(n36488), .A(n36486), .B(n36487), .ZN(
        n1264) );
  AND3_X1 U6190 ( .A1(n17064), .A2(n17061), .A3(n17062), .ZN(n1265) );
  XNOR2_X1 U6194 ( .A(n1266), .B(n45319), .ZN(n45323) );
  XNOR2_X1 U6195 ( .A(n1544), .B(n45449), .ZN(n1266) );
  NAND2_X1 U6196 ( .A1(n50276), .A2(n5617), .ZN(n44589) );
  NAND2_X1 U6198 ( .A1(n45921), .A2(n42886), .ZN(n49235) );
  XNOR2_X2 U6200 ( .A(n16749), .B(n17218), .ZN(n16973) );
  NAND2_X1 U6201 ( .A1(n30117), .A2(n31870), .ZN(n2967) );
  NAND2_X1 U6203 ( .A1(n1267), .A2(n15204), .ZN(n15236) );
  NOR2_X1 U6205 ( .A1(n13211), .A2(n13210), .ZN(n1268) );
  NAND2_X1 U6206 ( .A1(n31391), .A2(n1269), .ZN(n31392) );
  NAND2_X1 U6207 ( .A1(n5300), .A2(n402), .ZN(n29938) );
  NOR2_X1 U6209 ( .A1(n49691), .A2(n49254), .ZN(n49699) );
  NAND3_X1 U6210 ( .A1(n29011), .A2(n29008), .A3(n29007), .ZN(n29009) );
  NAND2_X1 U6211 ( .A1(n46343), .A2(n46344), .ZN(n46348) );
  NAND2_X1 U6212 ( .A1(n24668), .A2(n26734), .ZN(n24670) );
  BUF_X2 U6213 ( .A(n8988), .Z(n11341) );
  NAND2_X1 U6214 ( .A1(n2211), .A2(n11485), .ZN(n12483) );
  NAND2_X1 U6216 ( .A1(n23756), .A2(n24190), .ZN(n22601) );
  XNOR2_X1 U6217 ( .A(n18697), .B(n18831), .ZN(n15899) );
  OAI21_X1 U6220 ( .B1(n32887), .B2(n33041), .A(n32865), .ZN(n30968) );
  AND4_X2 U6221 ( .A1(n18737), .A2(n18735), .A3(n18736), .A4(n18734), .ZN(
        n24180) );
  NAND2_X1 U6222 ( .A1(n23705), .A2(n22235), .ZN(n3823) );
  NAND2_X1 U6223 ( .A1(n11697), .A2(n9500), .ZN(n9501) );
  OR2_X2 U6226 ( .A1(n739), .A2(n2201), .ZN(n30167) );
  NOR2_X1 U6227 ( .A1(n1272), .A2(n1271), .ZN(n41591) );
  NOR2_X1 U6228 ( .A1(n42000), .A2(n42020), .ZN(n1271) );
  INV_X1 U6229 ( .A(n41586), .ZN(n1272) );
  NAND2_X1 U6230 ( .A1(n22864), .A2(n1273), .ZN(n22858) );
  XNOR2_X1 U6231 ( .A(n43303), .B(n43250), .ZN(n1274) );
  XNOR2_X1 U6232 ( .A(n1275), .B(n47864), .ZN(Plaintext[28]) );
  NAND4_X1 U6233 ( .A1(n47863), .A2(n47861), .A3(n47862), .A4(n47860), .ZN(
        n1275) );
  XNOR2_X1 U6236 ( .A(n1277), .B(n41823), .ZN(n41824) );
  XNOR2_X1 U6237 ( .A(n5433), .B(n5434), .ZN(n1277) );
  NAND3_X1 U6238 ( .A1(n12454), .A2(n50997), .A3(n12464), .ZN(n11493) );
  XNOR2_X1 U6240 ( .A(n1278), .B(n25153), .ZN(n8736) );
  NAND2_X1 U6241 ( .A1(n19900), .A2(n25064), .ZN(n1279) );
  NAND2_X1 U6242 ( .A1(n11037), .A2(n1281), .ZN(n1280) );
  INV_X1 U6243 ( .A(n13188), .ZN(n10083) );
  NAND2_X1 U6244 ( .A1(n10904), .A2(n1282), .ZN(n13188) );
  AND3_X2 U6245 ( .A1(n23115), .A2(n4970), .A3(n324), .ZN(n31778) );
  INV_X1 U6246 ( .A(n14552), .ZN(n3038) );
  NAND2_X1 U6247 ( .A1(n1283), .A2(n14552), .ZN(n13352) );
  NAND4_X2 U6249 ( .A1(n50311), .A2(n50312), .A3(n50313), .A4(n50310), .ZN(
        n50485) );
  NAND2_X1 U6251 ( .A1(n1284), .A2(n47150), .ZN(n1922) );
  NAND2_X1 U6252 ( .A1(n2708), .A2(n4290), .ZN(n1284) );
  NAND3_X2 U6253 ( .A1(n1986), .A2(n1987), .A3(n32336), .ZN(n5045) );
  NAND3_X1 U6254 ( .A1(n29544), .A2(n1286), .A3(n1285), .ZN(n29548) );
  NAND2_X1 U6255 ( .A1(n8453), .A2(n29541), .ZN(n1286) );
  NAND2_X1 U6256 ( .A1(n37154), .A2(n39173), .ZN(n37157) );
  NAND2_X1 U6257 ( .A1(n5204), .A2(n24041), .ZN(n5203) );
  NAND4_X2 U6258 ( .A1(n27046), .A2(n1541), .A3(n27045), .A4(n27044), .ZN(
        n31346) );
  INV_X1 U6260 ( .A(n15376), .ZN(n1287) );
  NAND2_X1 U6261 ( .A1(n15382), .A2(n15381), .ZN(n15376) );
  NAND2_X1 U6263 ( .A1(n41265), .A2(n41113), .ZN(n39593) );
  OR2_X2 U6264 ( .A1(n6398), .A2(n31024), .ZN(n34881) );
  INV_X1 U6266 ( .A(n1741), .ZN(n1289) );
  NAND3_X1 U6267 ( .A1(n50370), .A2(n50367), .A3(n3607), .ZN(n47136) );
  NAND3_X1 U6268 ( .A1(n37800), .A2(n39473), .A3(n37801), .ZN(n37803) );
  NAND2_X1 U6269 ( .A1(n39474), .A2(n37804), .ZN(n37800) );
  NAND3_X1 U6270 ( .A1(n1291), .A2(n31955), .A3(n718), .ZN(n1290) );
  INV_X1 U6271 ( .A(n32047), .ZN(n1291) );
  NAND2_X1 U6272 ( .A1(n32043), .A2(n1293), .ZN(n1292) );
  INV_X1 U6273 ( .A(n718), .ZN(n1293) );
  XNOR2_X1 U6274 ( .A(n17674), .B(n2339), .ZN(n1294) );
  NOR2_X1 U6276 ( .A1(n47713), .A2(n1298), .ZN(n1297) );
  NAND2_X1 U6277 ( .A1(n47722), .A2(n47723), .ZN(n1298) );
  NAND2_X1 U6278 ( .A1(n47714), .A2(n47715), .ZN(n1299) );
  NOR2_X1 U6279 ( .A1(n30291), .A2(n30279), .ZN(n3870) );
  NAND2_X1 U6280 ( .A1(n32151), .A2(n32787), .ZN(n32777) );
  OR2_X1 U6282 ( .A1(n2030), .A2(n31815), .ZN(n2029) );
  NAND2_X2 U6283 ( .A1(n3835), .A2(n36435), .ZN(n41049) );
  XNOR2_X1 U6284 ( .A(n42222), .B(n51333), .ZN(n43558) );
  INV_X1 U6286 ( .A(n29531), .ZN(n26700) );
  NAND2_X1 U6287 ( .A1(n29518), .A2(n29513), .ZN(n29531) );
  NAND2_X1 U6288 ( .A1(n40683), .A2(n39673), .ZN(n38410) );
  AND4_X2 U6289 ( .A1(n36626), .A2(n36624), .A3(n36625), .A4(n36623), .ZN(
        n39673) );
  NAND2_X1 U6290 ( .A1(n1300), .A2(n12625), .ZN(n12079) );
  NAND2_X1 U6291 ( .A1(n4041), .A2(n12638), .ZN(n1300) );
  NAND2_X1 U6292 ( .A1(n8171), .A2(n8172), .ZN(n29910) );
  NAND2_X1 U6293 ( .A1(n22446), .A2(n321), .ZN(n22447) );
  NAND2_X1 U6294 ( .A1(n18989), .A2(n3604), .ZN(n7099) );
  NAND2_X1 U6295 ( .A1(n31956), .A2(n31323), .ZN(n1560) );
  INV_X1 U6296 ( .A(n17868), .ZN(n6516) );
  NAND2_X1 U6297 ( .A1(n2222), .A2(n17466), .ZN(n17868) );
  NAND2_X2 U6298 ( .A1(n4170), .A2(n3012), .ZN(n16011) );
  AND2_X1 U6299 ( .A1(n20418), .A2(n20419), .ZN(n1859) );
  NAND2_X1 U6300 ( .A1(n32210), .A2(n6969), .ZN(n32207) );
  NAND2_X1 U6302 ( .A1(n39912), .A2(n38448), .ZN(n39789) );
  XNOR2_X2 U6303 ( .A(n44370), .B(n43943), .ZN(n43363) );
  NAND3_X2 U6304 ( .A1(n39165), .A2(n1301), .A3(n39164), .ZN(n44370) );
  NAND2_X1 U6305 ( .A1(n27108), .A2(n27107), .ZN(n3465) );
  NAND2_X1 U6306 ( .A1(n6765), .A2(n26621), .ZN(n27107) );
  NAND2_X1 U6307 ( .A1(n12616), .A2(n12617), .ZN(n12623) );
  NAND3_X1 U6308 ( .A1(n12885), .A2(n13204), .A3(n1303), .ZN(n1302) );
  NAND2_X1 U6309 ( .A1(n781), .A2(n13930), .ZN(n1303) );
  NAND2_X1 U6312 ( .A1(n6761), .A2(n8394), .ZN(n25457) );
  NAND2_X1 U6314 ( .A1(n3002), .A2(n23344), .ZN(n23346) );
  NAND2_X1 U6315 ( .A1(n17469), .A2(n17559), .ZN(n17470) );
  NAND3_X1 U6317 ( .A1(n9545), .A2(n3376), .A3(n9544), .ZN(n9546) );
  AOI21_X1 U6318 ( .B1(n22904), .B2(n22918), .A(n1305), .ZN(n22361) );
  NAND2_X1 U6319 ( .A1(n49672), .A2(n49657), .ZN(n49651) );
  NAND2_X1 U6320 ( .A1(n36047), .A2(n35215), .ZN(n36457) );
  OR2_X2 U6322 ( .A1(n1306), .A2(n9556), .ZN(n15259) );
  NAND3_X1 U6324 ( .A1(n35003), .A2(n38391), .A3(n39601), .ZN(n35009) );
  NAND2_X1 U6325 ( .A1(n42042), .A2(n40295), .ZN(n42052) );
  XNOR2_X2 U6329 ( .A(n1308), .B(n42560), .ZN(n43698) );
  NAND2_X1 U6330 ( .A1(n42212), .A2(n8476), .ZN(n1308) );
  OAI21_X1 U6331 ( .B1(n36212), .B2(n36213), .A(n38971), .ZN(n36220) );
  NAND2_X1 U6332 ( .A1(n38043), .A2(n34945), .ZN(n34938) );
  NAND2_X1 U6333 ( .A1(n29740), .A2(n29741), .ZN(n29742) );
  NAND2_X1 U6334 ( .A1(n1758), .A2(n45184), .ZN(n45185) );
  NAND2_X1 U6336 ( .A1(n49689), .A2(n51095), .ZN(n44743) );
  OR2_X2 U6337 ( .A1(n1310), .A2(n7866), .ZN(n50958) );
  NAND4_X1 U6338 ( .A1(n5084), .A2(n7867), .A3(n46733), .A4(n45191), .ZN(n1310) );
  NAND3_X1 U6339 ( .A1(n13072), .A2(n13071), .A3(n14784), .ZN(n13073) );
  NAND3_X1 U6341 ( .A1(n37888), .A2(n38997), .A3(n4152), .ZN(n37891) );
  INV_X1 U6342 ( .A(n26954), .ZN(n26772) );
  INV_X1 U6343 ( .A(n38363), .ZN(n38364) );
  NAND2_X1 U6344 ( .A1(n41077), .A2(n39140), .ZN(n38363) );
  INV_X1 U6345 ( .A(n47135), .ZN(n46799) );
  NAND2_X1 U6346 ( .A1(n46989), .A2(n43798), .ZN(n47135) );
  NAND2_X1 U6348 ( .A1(n14036), .A2(n14023), .ZN(n12406) );
  NAND2_X1 U6349 ( .A1(n50367), .A2(n6811), .ZN(n46979) );
  XNOR2_X1 U6350 ( .A(n34554), .B(n34555), .ZN(n34557) );
  XNOR2_X2 U6351 ( .A(n34382), .B(n36930), .ZN(n34555) );
  NAND2_X1 U6354 ( .A1(n1317), .A2(n14400), .ZN(n12862) );
  AOI21_X1 U6356 ( .B1(n19821), .B2(n19820), .A(n1318), .ZN(n2256) );
  NAND2_X2 U6359 ( .A1(n1520), .A2(n1320), .ZN(n19235) );
  AND3_X1 U6360 ( .A1(n1912), .A2(n12414), .A3(n12408), .ZN(n1320) );
  NAND2_X1 U6361 ( .A1(n1321), .A2(n47205), .ZN(n6696) );
  NAND2_X1 U6362 ( .A1(n2694), .A2(n2833), .ZN(n1321) );
  NAND3_X1 U6363 ( .A1(n15422), .A2(n14875), .A3(n15424), .ZN(n1832) );
  NAND2_X1 U6364 ( .A1(n14880), .A2(n15425), .ZN(n15424) );
  OR2_X2 U6365 ( .A1(n2020), .A2(n2022), .ZN(n7115) );
  INV_X1 U6366 ( .A(n12605), .ZN(n12598) );
  NAND2_X1 U6367 ( .A1(n3377), .A2(n11921), .ZN(n12605) );
  NAND3_X2 U6370 ( .A1(n13157), .A2(n13158), .A3(n13159), .ZN(n18399) );
  MUX2_X1 U6371 ( .A(n36398), .B(n2141), .S(n37637), .Z(n37653) );
  XNOR2_X1 U6372 ( .A(n1324), .B(n4065), .ZN(Plaintext[85]) );
  NOR2_X1 U6373 ( .A1(n46961), .A2(n46962), .ZN(n1324) );
  NAND3_X2 U6374 ( .A1(n1530), .A2(n34915), .A3(n1527), .ZN(n41975) );
  AOI22_X1 U6375 ( .A1(n37226), .A2(n38636), .B1(n38265), .B2(n37227), .ZN(
        n37232) );
  OAI21_X1 U6379 ( .B1(n1727), .B2(n1726), .A(n45755), .ZN(n1725) );
  INV_X1 U6382 ( .A(n39775), .ZN(n39774) );
  NAND2_X1 U6383 ( .A1(n7704), .A2(n41446), .ZN(n39775) );
  XNOR2_X1 U6384 ( .A(n1327), .B(n49502), .ZN(Plaintext[116]) );
  NAND4_X1 U6385 ( .A1(n49499), .A2(n49498), .A3(n49500), .A4(n49501), .ZN(
        n1327) );
  INV_X1 U6386 ( .A(n35874), .ZN(n35873) );
  INV_X1 U6388 ( .A(n540), .ZN(n46252) );
  NOR2_X1 U6390 ( .A1(n31215), .A2(n32199), .ZN(n32208) );
  INV_X1 U6391 ( .A(n38448), .ZN(n1874) );
  OR2_X1 U6392 ( .A1(n36454), .A2(n36589), .ZN(n1691) );
  OAI211_X1 U6393 ( .C1(n49492), .C2(n49522), .A(n49491), .B(n49534), .ZN(
        n49493) );
  NAND2_X1 U6395 ( .A1(n45820), .A2(n45524), .ZN(n1328) );
  XNOR2_X1 U6396 ( .A(n1329), .B(n47802), .ZN(Plaintext[23]) );
  NAND4_X1 U6397 ( .A1(n47801), .A2(n47799), .A3(n47800), .A4(n4588), .ZN(
        n1329) );
  NAND2_X1 U6398 ( .A1(n47779), .A2(n1330), .ZN(n47784) );
  INV_X1 U6400 ( .A(n47793), .ZN(n1331) );
  NAND2_X1 U6401 ( .A1(n1334), .A2(n1333), .ZN(n1332) );
  NAND2_X1 U6403 ( .A1(n22638), .A2(n23599), .ZN(n23609) );
  NAND2_X1 U6404 ( .A1(n12363), .A2(n12364), .ZN(n12365) );
  NOR2_X1 U6407 ( .A1(n30759), .A2(n730), .ZN(n1899) );
  NAND3_X2 U6408 ( .A1(n8674), .A2(n3330), .A3(n23004), .ZN(n25124) );
  NOR2_X1 U6409 ( .A1(n38109), .A2(n38110), .ZN(n38113) );
  NAND3_X1 U6410 ( .A1(n12108), .A2(n12107), .A3(n12106), .ZN(n4778) );
  NAND2_X1 U6411 ( .A1(n12112), .A2(n11374), .ZN(n12108) );
  NAND2_X1 U6412 ( .A1(n14553), .A2(n14550), .ZN(n14535) );
  NAND3_X1 U6413 ( .A1(n24159), .A2(n23277), .A3(n23821), .ZN(n21798) );
  NAND2_X1 U6414 ( .A1(n12429), .A2(n12430), .ZN(n12433) );
  OAI21_X1 U6415 ( .B1(n39011), .B2(n37200), .A(n36770), .ZN(n1335) );
  XNOR2_X1 U6417 ( .A(n1337), .B(n32585), .ZN(n32607) );
  XNOR2_X1 U6418 ( .A(n35120), .B(n35659), .ZN(n1337) );
  NAND2_X1 U6420 ( .A1(n23638), .A2(n23622), .ZN(n5066) );
  NAND3_X1 U6421 ( .A1(n2308), .A2(n48549), .A3(n1340), .ZN(n48553) );
  NAND4_X2 U6422 ( .A1(n29383), .A2(n3657), .A3(n3656), .A4(n29384), .ZN(
        n36932) );
  NAND4_X2 U6423 ( .A1(n48560), .A2(n48559), .A3(n48558), .A4(n48557), .ZN(
        n48633) );
  NAND3_X1 U6424 ( .A1(n51257), .A2(n30399), .A3(n28758), .ZN(n29935) );
  XNOR2_X1 U6426 ( .A(n1342), .B(n25918), .ZN(n25933) );
  XNOR2_X1 U6427 ( .A(n25932), .B(n25919), .ZN(n1342) );
  NAND3_X1 U6428 ( .A1(n32699), .A2(n28596), .A3(n5217), .ZN(n31665) );
  XNOR2_X2 U6429 ( .A(n18749), .B(n18739), .ZN(n3142) );
  NOR2_X1 U6430 ( .A1(n1344), .A2(n1343), .ZN(n1549) );
  NOR2_X1 U6431 ( .A1(n31147), .A2(n31148), .ZN(n1344) );
  OAI21_X1 U6432 ( .B1(n27805), .B2(n1817), .A(n1814), .ZN(n27826) );
  OAI21_X1 U6433 ( .B1(n2060), .B2(n2059), .A(n2137), .ZN(n4088) );
  NAND2_X2 U6434 ( .A1(n1345), .A2(n1558), .ZN(n27241) );
  XNOR2_X1 U6436 ( .A(n25176), .B(n22554), .ZN(n22569) );
  XNOR2_X2 U6437 ( .A(n51009), .B(n25365), .ZN(n25176) );
  NAND2_X1 U6438 ( .A1(n17891), .A2(n3083), .ZN(n5186) );
  XNOR2_X2 U6439 ( .A(n1673), .B(n44893), .ZN(n46118) );
  NAND2_X1 U6441 ( .A1(n23986), .A2(n22426), .ZN(n22531) );
  OAI21_X1 U6442 ( .B1(n40204), .B2(n38777), .A(n1347), .ZN(n36095) );
  INV_X1 U6443 ( .A(n36094), .ZN(n1347) );
  INV_X1 U6444 ( .A(n30391), .ZN(n1348) );
  AND3_X2 U6445 ( .A1(n23863), .A2(n23862), .A3(n3532), .ZN(n3535) );
  NAND2_X1 U6446 ( .A1(n15770), .A2(n15068), .ZN(n15767) );
  NAND3_X1 U6447 ( .A1(n1349), .A2(n37762), .A3(n37764), .ZN(n37771) );
  NAND2_X1 U6448 ( .A1(n37760), .A2(n37761), .ZN(n1349) );
  NAND4_X1 U6449 ( .A1(n37785), .A2(n37776), .A3(n37784), .A4(n37777), .ZN(
        n1465) );
  NAND3_X1 U6450 ( .A1(n1511), .A2(n46604), .A3(n5022), .ZN(n1510) );
  XNOR2_X1 U6452 ( .A(n1350), .B(n28108), .ZN(n28110) );
  XNOR2_X1 U6453 ( .A(n28432), .B(n28107), .ZN(n1350) );
  NAND2_X1 U6454 ( .A1(n32397), .A2(n32398), .ZN(n32400) );
  NAND2_X1 U6455 ( .A1(n2777), .A2(n29896), .ZN(n29897) );
  NAND2_X1 U6456 ( .A1(n37585), .A2(n35452), .ZN(n37598) );
  NAND2_X1 U6457 ( .A1(n1779), .A2(n4017), .ZN(n21127) );
  AOI21_X1 U6459 ( .B1(n13292), .B2(n13293), .A(n14033), .ZN(n1351) );
  INV_X2 U6460 ( .A(n5693), .ZN(n5056) );
  OAI21_X1 U6463 ( .B1(n48971), .B2(n48931), .A(n46950), .ZN(n46952) );
  XNOR2_X1 U6466 ( .A(n1353), .B(n6146), .ZN(n5788) );
  XNOR2_X1 U6467 ( .A(n35806), .B(n35802), .ZN(n1353) );
  NAND3_X1 U6468 ( .A1(n28146), .A2(n24882), .A3(n28560), .ZN(n24884) );
  OAI211_X1 U6469 ( .C1(n49929), .C2(n47423), .A(n49933), .B(n1355), .ZN(
        n46174) );
  NAND2_X1 U6470 ( .A1(n47425), .A2(n49932), .ZN(n1355) );
  NAND2_X1 U6471 ( .A1(n1356), .A2(n49899), .ZN(n47425) );
  INV_X1 U6472 ( .A(n49889), .ZN(n1356) );
  NAND3_X1 U6473 ( .A1(n652), .A2(n49916), .A3(n7345), .ZN(n49929) );
  INV_X1 U6474 ( .A(n49889), .ZN(n7345) );
  XNOR2_X1 U6475 ( .A(n7121), .B(n1357), .ZN(n45366) );
  XNOR2_X1 U6477 ( .A(n42961), .B(n1357), .ZN(n41991) );
  XNOR2_X1 U6478 ( .A(n42534), .B(n1357), .ZN(n41882) );
  NAND4_X1 U6480 ( .A1(n14583), .A2(n1359), .A3(n5209), .A4(n15157), .ZN(n7712) );
  NAND2_X1 U6481 ( .A1(n6383), .A2(n51370), .ZN(n15157) );
  INV_X1 U6482 ( .A(n1360), .ZN(n36639) );
  INV_X1 U6483 ( .A(n34186), .ZN(n38078) );
  NAND4_X1 U6484 ( .A1(n20816), .A2(n1363), .A3(n1362), .A4(n1361), .ZN(n20835) );
  NAND3_X1 U6486 ( .A1(n1367), .A2(n763), .A3(n1369), .ZN(n1362) );
  NAND2_X1 U6487 ( .A1(n759), .A2(n1364), .ZN(n1363) );
  OAI21_X1 U6488 ( .B1(n20811), .B2(n20821), .A(n51754), .ZN(n1367) );
  INV_X1 U6490 ( .A(n21495), .ZN(n1370) );
  NAND2_X1 U6492 ( .A1(n1371), .A2(n2638), .ZN(n41145) );
  AND2_X1 U6493 ( .A1(n38624), .A2(n1371), .ZN(n4510) );
  NAND2_X1 U6494 ( .A1(n2639), .A2(n38617), .ZN(n1371) );
  INV_X1 U6495 ( .A(n30788), .ZN(n30791) );
  NAND2_X1 U6496 ( .A1(n1375), .A2(n29900), .ZN(n1373) );
  NOR2_X1 U6499 ( .A1(n2774), .A2(n1042), .ZN(n1375) );
  NAND2_X1 U6500 ( .A1(n398), .A2(n29507), .ZN(n26977) );
  XNOR2_X1 U6501 ( .A(n26119), .B(n1377), .ZN(n26121) );
  XNOR2_X1 U6502 ( .A(n44399), .B(n1378), .ZN(n45597) );
  XNOR2_X1 U6503 ( .A(n44398), .B(n1379), .ZN(n1378) );
  INV_X1 U6504 ( .A(n44397), .ZN(n1379) );
  XNOR2_X1 U6505 ( .A(n40021), .B(n42504), .ZN(n44398) );
  NAND2_X1 U6506 ( .A1(n39981), .A2(n40436), .ZN(n1380) );
  INV_X1 U6507 ( .A(n1382), .ZN(n1381) );
  NOR2_X1 U6508 ( .A1(n47786), .A2(n1383), .ZN(n47740) );
  NAND2_X1 U6509 ( .A1(n47778), .A2(n47745), .ZN(n1383) );
  XNOR2_X1 U6510 ( .A(n24533), .B(n1384), .ZN(n24536) );
  XNOR2_X1 U6511 ( .A(n1384), .B(n24275), .ZN(n24276) );
  XNOR2_X1 U6512 ( .A(n1384), .B(n24729), .ZN(n24730) );
  XNOR2_X1 U6513 ( .A(n24644), .B(n1384), .ZN(n24645) );
  XNOR2_X2 U6514 ( .A(n19627), .B(n28311), .ZN(n1384) );
  XNOR2_X2 U6515 ( .A(n5910), .B(n5909), .ZN(n36428) );
  NAND2_X1 U6517 ( .A1(n32439), .A2(n1385), .ZN(n31954) );
  NOR2_X1 U6520 ( .A1(n1385), .A2(n32438), .ZN(n32359) );
  NOR2_X1 U6521 ( .A1(n1385), .A2(n32345), .ZN(n32437) );
  NAND2_X1 U6522 ( .A1(n3703), .A2(n1385), .ZN(n3702) );
  NAND2_X1 U6523 ( .A1(n718), .A2(n1385), .ZN(n32442) );
  OAI22_X1 U6524 ( .A1(n32352), .A2(n32047), .B1(n32048), .B2(n1385), .ZN(
        n32049) );
  NAND3_X1 U6527 ( .A1(n2837), .A2(n32436), .A3(n718), .ZN(n1387) );
  INV_X1 U6529 ( .A(n40462), .ZN(n1390) );
  NAND2_X1 U6530 ( .A1(n737), .A2(n2144), .ZN(n24569) );
  NAND2_X1 U6531 ( .A1(n1716), .A2(n1392), .ZN(n47892) );
  NAND4_X1 U6532 ( .A1(n30144), .A2(n1393), .A3(n32332), .A4(n30143), .ZN(
        n30145) );
  NAND3_X1 U6533 ( .A1(n2012), .A2(n28598), .A3(n1393), .ZN(n28601) );
  NAND3_X1 U6534 ( .A1(n52301), .A2(n30140), .A3(n31668), .ZN(n1393) );
  NAND2_X1 U6537 ( .A1(n29825), .A2(n51640), .ZN(n1395) );
  NAND3_X1 U6538 ( .A1(n31587), .A2(n29827), .A3(n31632), .ZN(n1397) );
  NAND2_X1 U6539 ( .A1(n7705), .A2(n31631), .ZN(n31587) );
  NAND3_X2 U6540 ( .A1(n17043), .A2(n1398), .A3(n8411), .ZN(n23360) );
  NAND2_X1 U6541 ( .A1(n6433), .A2(n23360), .ZN(n23351) );
  AOI22_X1 U6542 ( .A1(n23549), .A2(n23550), .B1(n23551), .B2(n23563), .ZN(
        n23578) );
  NAND2_X1 U6544 ( .A1(n41732), .A2(n41733), .ZN(n1400) );
  NAND2_X1 U6545 ( .A1(n41737), .A2(n1402), .ZN(n1401) );
  NAND2_X1 U6546 ( .A1(n39599), .A2(n41110), .ZN(n41737) );
  OAI21_X1 U6547 ( .B1(n21232), .B2(n765), .A(n1405), .ZN(n1404) );
  NAND2_X1 U6548 ( .A1(n21235), .A2(n19518), .ZN(n1405) );
  INV_X1 U6549 ( .A(n21232), .ZN(n1406) );
  NAND2_X1 U6550 ( .A1(n17036), .A2(n1407), .ZN(n17035) );
  NAND2_X1 U6551 ( .A1(n21232), .A2(n761), .ZN(n1407) );
  NAND4_X2 U6552 ( .A1(n41361), .A2(n8122), .A3(n1409), .A4(n1408), .ZN(n43131) );
  NAND2_X1 U6553 ( .A1(n41353), .A2(n6471), .ZN(n1410) );
  OR3_X1 U6554 ( .A1(n23213), .A2(n23230), .A3(n413), .ZN(n23235) );
  INV_X1 U6555 ( .A(n18371), .ZN(n1411) );
  NAND3_X1 U6556 ( .A1(n23549), .A2(n22274), .A3(n7832), .ZN(n1412) );
  NAND2_X1 U6557 ( .A1(n22274), .A2(n22272), .ZN(n1413) );
  NAND2_X1 U6558 ( .A1(n23549), .A2(n7832), .ZN(n22273) );
  OR2_X1 U6559 ( .A1(n19071), .A2(n20144), .ZN(n1418) );
  NAND2_X1 U6560 ( .A1(n18356), .A2(n18357), .ZN(n20135) );
  INV_X1 U6561 ( .A(n20147), .ZN(n1414) );
  INV_X1 U6564 ( .A(n1417), .ZN(n20134) );
  INV_X1 U6566 ( .A(n20135), .ZN(n1419) );
  AND2_X1 U6568 ( .A1(n10166), .A2(n11033), .ZN(n1422) );
  NAND2_X1 U6569 ( .A1(n20021), .A2(n6952), .ZN(n1423) );
  NAND3_X1 U6570 ( .A1(n20021), .A2(n6952), .A3(n18287), .ZN(n18283) );
  NOR2_X1 U6571 ( .A1(n51208), .A2(n1423), .ZN(n17491) );
  NAND2_X1 U6572 ( .A1(n30968), .A2(n31526), .ZN(n1424) );
  NAND4_X1 U6573 ( .A1(n5497), .A2(n719), .A3(n32883), .A4(n32874), .ZN(n31526) );
  NAND2_X1 U6574 ( .A1(n1424), .A2(n32645), .ZN(n30973) );
  NAND2_X1 U6576 ( .A1(n51520), .A2(n1428), .ZN(n32395) );
  NAND3_X2 U6577 ( .A1(n1429), .A2(n3153), .A3(n29117), .ZN(n1428) );
  NAND2_X1 U6578 ( .A1(n32408), .A2(n1428), .ZN(n31947) );
  NOR2_X1 U6579 ( .A1(n1426), .A2(n714), .ZN(n1425) );
  AND2_X1 U6580 ( .A1(n1428), .A2(n32071), .ZN(n1427) );
  NAND3_X1 U6581 ( .A1(n31285), .A2(n32396), .A3(n1428), .ZN(n31288) );
  NAND3_X2 U6582 ( .A1(n22512), .A2(n22511), .A3(n1430), .ZN(n25506) );
  NAND2_X1 U6583 ( .A1(n1431), .A2(n22820), .ZN(n22821) );
  NAND3_X1 U6584 ( .A1(n8586), .A2(n22826), .A3(n22490), .ZN(n1431) );
  NAND2_X1 U6586 ( .A1(n1433), .A2(n52102), .ZN(n1432) );
  NAND2_X1 U6587 ( .A1(n2158), .A2(n30256), .ZN(n1433) );
  NAND2_X1 U6588 ( .A1(n14651), .A2(n14660), .ZN(n1436) );
  NAND2_X1 U6589 ( .A1(n14650), .A2(n1439), .ZN(n1437) );
  NAND2_X1 U6590 ( .A1(n1440), .A2(n39271), .ZN(n37943) );
  NAND3_X1 U6591 ( .A1(n39264), .A2(n2571), .A3(n2100), .ZN(n1440) );
  NAND2_X1 U6592 ( .A1(n1441), .A2(n601), .ZN(n50831) );
  NAND2_X1 U6593 ( .A1(n1441), .A2(n50837), .ZN(n50847) );
  NOR2_X1 U6594 ( .A1(n1441), .A2(n50837), .ZN(n50882) );
  NAND2_X1 U6595 ( .A1(n52097), .A2(n1441), .ZN(n50836) );
  NAND2_X1 U6596 ( .A1(n50848), .A2(n1441), .ZN(n50849) );
  XNOR2_X1 U6597 ( .A(n1442), .B(n50825), .ZN(Plaintext[180]) );
  NAND4_X1 U6598 ( .A1(n50824), .A2(n6815), .A3(n1446), .A4(n1443), .ZN(n1442)
         );
  NAND2_X1 U6599 ( .A1(n50822), .A2(n50835), .ZN(n1444) );
  NAND2_X1 U6600 ( .A1(n50872), .A2(n51312), .ZN(n1445) );
  NAND2_X1 U6601 ( .A1(n50821), .A2(n50839), .ZN(n1446) );
  NAND2_X1 U6602 ( .A1(n11752), .A2(n483), .ZN(n1447) );
  NAND2_X1 U6604 ( .A1(n21970), .A2(n23477), .ZN(n21343) );
  NAND2_X1 U6605 ( .A1(n23479), .A2(n23481), .ZN(n23477) );
  NAND2_X1 U6606 ( .A1(n8818), .A2(n10161), .ZN(n10003) );
  NAND2_X1 U6607 ( .A1(n10165), .A2(n11025), .ZN(n9822) );
  OAI21_X1 U6608 ( .B1(n316), .B2(n20836), .A(n3493), .ZN(n20846) );
  NAND2_X1 U6609 ( .A1(n24154), .A2(n1450), .ZN(n23829) );
  NAND3_X1 U6611 ( .A1(n6727), .A2(n19984), .A3(n21626), .ZN(n1452) );
  NAND2_X1 U6612 ( .A1(n10546), .A2(n9830), .ZN(n10182) );
  AND2_X1 U6613 ( .A1(n1454), .A2(n319), .ZN(n17416) );
  NAND4_X1 U6614 ( .A1(n17414), .A2(n17415), .A3(n319), .A4(n1454), .ZN(n1576)
         );
  NAND2_X1 U6618 ( .A1(n7050), .A2(n598), .ZN(n21223) );
  INV_X1 U6619 ( .A(n770), .ZN(n1456) );
  OAI21_X1 U6620 ( .B1(n1462), .B2(n10537), .A(n1459), .ZN(n1457) );
  NAND3_X1 U6621 ( .A1(n1457), .A2(n8288), .A3(n13779), .ZN(n13160) );
  OR2_X1 U6622 ( .A1(n2037), .A2(n30503), .ZN(n32980) );
  NAND2_X1 U6623 ( .A1(n712), .A2(n1458), .ZN(n30503) );
  INV_X1 U6624 ( .A(n32980), .ZN(n32985) );
  NAND2_X1 U6625 ( .A1(n5493), .A2(n20841), .ZN(n5492) );
  NOR2_X1 U6626 ( .A1(n1796), .A2(n19156), .ZN(n20841) );
  NAND3_X1 U6627 ( .A1(n10544), .A2(n1461), .A3(n1460), .ZN(n1459) );
  NAND2_X1 U6628 ( .A1(n10555), .A2(n10043), .ZN(n1460) );
  OAI21_X1 U6629 ( .B1(n10549), .B2(n10186), .A(n10042), .ZN(n1462) );
  XNOR2_X2 U6630 ( .A(n33550), .B(n1463), .ZN(n34294) );
  NAND4_X2 U6631 ( .A1(n31868), .A2(n31867), .A3(n32291), .A4(n31866), .ZN(
        n1463) );
  XNOR2_X1 U6632 ( .A(n1463), .B(n5616), .ZN(n35764) );
  XNOR2_X1 U6633 ( .A(n1463), .B(n35483), .ZN(n35276) );
  XNOR2_X1 U6634 ( .A(n1463), .B(n36759), .ZN(n36763) );
  XNOR2_X1 U6635 ( .A(n1463), .B(n34359), .ZN(n36993) );
  NOR2_X1 U6636 ( .A1(n42042), .A2(n1464), .ZN(n42047) );
  NAND2_X1 U6637 ( .A1(n3290), .A2(n1464), .ZN(n40050) );
  NAND2_X1 U6638 ( .A1(n47153), .A2(n43688), .ZN(n45159) );
  INV_X1 U6640 ( .A(n47464), .ZN(n47463) );
  NAND2_X1 U6641 ( .A1(n8450), .A2(n47620), .ZN(n47464) );
  NAND2_X2 U6642 ( .A1(n7678), .A2(n46602), .ZN(n47586) );
  NAND2_X1 U6643 ( .A1(n37778), .A2(n1469), .ZN(n36197) );
  NAND2_X1 U6644 ( .A1(n37778), .A2(n37774), .ZN(n35942) );
  NAND4_X2 U6646 ( .A1(n1679), .A2(n24356), .A3(n1677), .A4(n1471), .ZN(n32242) );
  INV_X1 U6647 ( .A(n31490), .ZN(n1472) );
  NAND3_X1 U6648 ( .A1(n722), .A2(n1472), .A3(n31489), .ZN(n31265) );
  NAND2_X1 U6649 ( .A1(n43178), .A2(n3278), .ZN(n1473) );
  NOR2_X1 U6650 ( .A1(n1477), .A2(n49980), .ZN(n47361) );
  INV_X1 U6652 ( .A(n47354), .ZN(n1477) );
  NOR2_X1 U6653 ( .A1(n49977), .A2(n47360), .ZN(n1478) );
  NAND2_X1 U6654 ( .A1(n51093), .A2(n43181), .ZN(n49977) );
  NAND2_X1 U6655 ( .A1(n47352), .A2(n47354), .ZN(n5506) );
  OR2_X2 U6656 ( .A1(n7216), .A2(n43147), .ZN(n47354) );
  NAND3_X1 U6657 ( .A1(n49972), .A2(n49990), .A3(n49978), .ZN(n47352) );
  NOR2_X1 U6658 ( .A1(n31648), .A2(n1479), .ZN(n2853) );
  OAI21_X1 U6659 ( .B1(n32465), .B2(n32716), .A(n1479), .ZN(n1936) );
  AOI21_X1 U6660 ( .B1(n32720), .B2(n1479), .A(n32729), .ZN(n32462) );
  XNOR2_X2 U6663 ( .A(n6680), .B(n33762), .ZN(n35973) );
  OAI21_X1 U6664 ( .B1(n17314), .B2(n19504), .A(n1481), .ZN(n17316) );
  NAND2_X1 U6666 ( .A1(n1483), .A2(n26774), .ZN(n26819) );
  NAND2_X1 U6667 ( .A1(n27578), .A2(n1484), .ZN(n1483) );
  AND2_X1 U6668 ( .A1(n31692), .A2(n31684), .ZN(n1485) );
  NAND2_X1 U6669 ( .A1(n2094), .A2(n31684), .ZN(n30981) );
  NAND2_X1 U6670 ( .A1(n4046), .A2(n6837), .ZN(n2094) );
  NAND3_X1 U6671 ( .A1(n1486), .A2(n14914), .A3(n14929), .ZN(n15303) );
  OAI21_X1 U6672 ( .B1(n43445), .B2(n1488), .A(n1487), .ZN(n43451) );
  NAND2_X1 U6673 ( .A1(n1085), .A2(n32719), .ZN(n32465) );
  NAND2_X1 U6674 ( .A1(n32724), .A2(n1085), .ZN(n32726) );
  NOR2_X1 U6676 ( .A1(n32732), .A2(n1085), .ZN(n29753) );
  NAND3_X1 U6677 ( .A1(n3239), .A2(n32731), .A3(n1085), .ZN(n32733) );
  XNOR2_X2 U6678 ( .A(n1491), .B(n43131), .ZN(n44893) );
  XNOR2_X1 U6679 ( .A(n1491), .B(n44240), .ZN(n40852) );
  XNOR2_X1 U6680 ( .A(n1491), .B(n42850), .ZN(n43238) );
  XNOR2_X1 U6681 ( .A(n1491), .B(n46111), .ZN(n43308) );
  NAND2_X1 U6682 ( .A1(n1495), .A2(n24248), .ZN(n1492) );
  INV_X1 U6684 ( .A(n24247), .ZN(n1497) );
  NOR2_X2 U6685 ( .A1(n23785), .A2(n21810), .ZN(n24248) );
  NAND2_X1 U6686 ( .A1(n38449), .A2(n39899), .ZN(n1604) );
  XNOR2_X1 U6687 ( .A(n6945), .B(n1500), .ZN(n1499) );
  INV_X1 U6689 ( .A(n49117), .ZN(n1501) );
  NAND2_X1 U6690 ( .A1(n49127), .A2(n1502), .ZN(n49115) );
  NOR2_X1 U6691 ( .A1(n49127), .A2(n1502), .ZN(n49122) );
  NAND2_X1 U6692 ( .A1(n49081), .A2(n1502), .ZN(n49082) );
  NAND2_X1 U6693 ( .A1(n44801), .A2(n1502), .ZN(n44802) );
  NAND2_X1 U6694 ( .A1(n49080), .A2(n1502), .ZN(n49087) );
  NOR2_X1 U6696 ( .A1(n49089), .A2(n1502), .ZN(n49067) );
  NAND2_X1 U6698 ( .A1(n40815), .A2(n39696), .ZN(n39511) );
  AND2_X1 U6699 ( .A1(n40822), .A2(n40835), .ZN(n39696) );
  NOR2_X1 U6700 ( .A1(n1504), .A2(n343), .ZN(n45037) );
  AOI21_X1 U6701 ( .B1(n1506), .B2(n1505), .A(n603), .ZN(n1504) );
  NAND2_X1 U6702 ( .A1(n46912), .A2(n46902), .ZN(n1505) );
  NAND2_X1 U6703 ( .A1(n1508), .A2(n1509), .ZN(n1506) );
  NAND2_X1 U6704 ( .A1(n659), .A2(n1507), .ZN(n1509) );
  INV_X1 U6706 ( .A(n1509), .ZN(n46915) );
  NAND2_X1 U6707 ( .A1(n45848), .A2(n51359), .ZN(n46918) );
  NAND2_X1 U6710 ( .A1(n5023), .A2(n46606), .ZN(n1511) );
  XNOR2_X1 U6712 ( .A(n1512), .B(n34620), .ZN(n31839) );
  XNOR2_X1 U6713 ( .A(n1512), .B(n32659), .ZN(n32673) );
  XNOR2_X1 U6714 ( .A(n1512), .B(n33691), .ZN(n33692) );
  XNOR2_X1 U6715 ( .A(n1512), .B(n7199), .ZN(n33314) );
  INV_X1 U6718 ( .A(n17441), .ZN(n1519) );
  NAND2_X1 U6719 ( .A1(n18064), .A2(n17440), .ZN(n17441) );
  NAND2_X1 U6721 ( .A1(n12407), .A2(n12409), .ZN(n1520) );
  XNOR2_X1 U6722 ( .A(n16011), .B(n17925), .ZN(n1521) );
  NAND2_X1 U6723 ( .A1(n675), .A2(n40139), .ZN(n2064) );
  NAND2_X1 U6724 ( .A1(n40820), .A2(n39689), .ZN(n40139) );
  NAND2_X1 U6727 ( .A1(n22902), .A2(n22901), .ZN(n1523) );
  NAND3_X1 U6728 ( .A1(n37766), .A2(n36247), .A3(n615), .ZN(n1524) );
  NAND3_X1 U6729 ( .A1(n1526), .A2(n36247), .A3(n692), .ZN(n1525) );
  INV_X1 U6730 ( .A(n37500), .ZN(n1526) );
  NAND3_X1 U6731 ( .A1(n1529), .A2(n36239), .A3(n1528), .ZN(n1527) );
  NAND2_X1 U6732 ( .A1(n34914), .A2(n691), .ZN(n1529) );
  NAND3_X1 U6733 ( .A1(n18100), .A2(n18872), .A3(n18101), .ZN(n1540) );
  NAND2_X1 U6735 ( .A1(n1532), .A2(n20672), .ZN(n1534) );
  INV_X1 U6736 ( .A(n18875), .ZN(n1532) );
  NAND3_X1 U6737 ( .A1(n5463), .A2(n18103), .A3(n18869), .ZN(n1533) );
  NAND2_X1 U6738 ( .A1(n20675), .A2(n18862), .ZN(n1535) );
  NAND2_X1 U6742 ( .A1(n1542), .A2(n27835), .ZN(n1541) );
  NAND2_X1 U6743 ( .A1(n27032), .A2(n27033), .ZN(n1542) );
  NAND3_X1 U6744 ( .A1(n45709), .A2(n48834), .A3(n1543), .ZN(n45710) );
  NAND2_X1 U6745 ( .A1(n48818), .A2(n1543), .ZN(n48820) );
  NAND2_X1 U6746 ( .A1(n48806), .A2(n45752), .ZN(n1543) );
  NAND4_X2 U6747 ( .A1(n39794), .A2(n39793), .A3(n39792), .A4(n39791), .ZN(
        n46050) );
  XNOR2_X1 U6748 ( .A(n45304), .B(n45303), .ZN(n1544) );
  NAND4_X2 U6750 ( .A1(n9284), .A2(n9285), .A3(n9283), .A4(n9282), .ZN(n11841)
         );
  INV_X1 U6752 ( .A(n23333), .ZN(n22264) );
  INV_X1 U6753 ( .A(n20376), .ZN(n20415) );
  OR2_X2 U6754 ( .A1(n776), .A2(n20376), .ZN(n21369) );
  NAND2_X1 U6755 ( .A1(n1547), .A2(n27834), .ZN(n1546) );
  NAND2_X2 U6756 ( .A1(n1548), .A2(n6300), .ZN(n31899) );
  OAI21_X1 U6757 ( .B1(n31151), .B2(n31149), .A(n31150), .ZN(n31897) );
  NAND2_X1 U6760 ( .A1(n1551), .A2(n725), .ZN(n1550) );
  NAND2_X1 U6762 ( .A1(n31897), .A2(n725), .ZN(n1552) );
  NOR2_X1 U6763 ( .A1(n1557), .A2(n1553), .ZN(n9274) );
  INV_X1 U6764 ( .A(n15412), .ZN(n1557) );
  NAND3_X1 U6765 ( .A1(n21982), .A2(n23485), .A3(n23487), .ZN(n1559) );
  XNOR2_X2 U6766 ( .A(n27241), .B(n26431), .ZN(n27289) );
  OAI21_X1 U6767 ( .B1(n32436), .B2(n32351), .A(n1560), .ZN(n31959) );
  NAND2_X1 U6768 ( .A1(n32056), .A2(n32345), .ZN(n31956) );
  NAND3_X1 U6770 ( .A1(n26829), .A2(n29908), .A3(n30789), .ZN(n2777) );
  NAND2_X1 U6771 ( .A1(n48847), .A2(n48898), .ZN(n48848) );
  NAND2_X1 U6772 ( .A1(n39628), .A2(n1561), .ZN(n39629) );
  NAND2_X1 U6773 ( .A1(n1562), .A2(n5318), .ZN(n40723) );
  AND4_X2 U6774 ( .A1(n1564), .A2(n26876), .A3(n26875), .A4(n1563), .ZN(n31484) );
  OAI21_X1 U6775 ( .B1(n722), .B2(n31490), .A(n31489), .ZN(n31491) );
  NAND3_X1 U6776 ( .A1(n2642), .A2(n1565), .A3(n27665), .ZN(n26870) );
  XNOR2_X2 U6778 ( .A(n24704), .B(n25803), .ZN(n2677) );
  AND2_X1 U6781 ( .A1(n41328), .A2(n41317), .ZN(n41326) );
  NAND3_X1 U6782 ( .A1(n46860), .A2(n46847), .A3(n46859), .ZN(n1567) );
  AND2_X1 U6783 ( .A1(n45778), .A2(n1567), .ZN(n1632) );
  NAND2_X1 U6787 ( .A1(n37762), .A2(n1569), .ZN(n4092) );
  NAND2_X1 U6788 ( .A1(n615), .A2(n37762), .ZN(n37513) );
  NAND2_X1 U6789 ( .A1(n37503), .A2(n1570), .ZN(n37504) );
  OR2_X1 U6790 ( .A1(n13930), .A2(n1571), .ZN(n13190) );
  AND2_X1 U6791 ( .A1(n13945), .A2(n1571), .ZN(n11862) );
  OAI21_X1 U6792 ( .B1(n2173), .B2(n13930), .A(n1571), .ZN(n13196) );
  NAND2_X1 U6793 ( .A1(n13949), .A2(n1571), .ZN(n12881) );
  NOR2_X1 U6794 ( .A1(n13949), .A2(n1571), .ZN(n13942) );
  NAND2_X1 U6795 ( .A1(n1575), .A2(n1572), .ZN(n7293) );
  NAND3_X1 U6796 ( .A1(n26976), .A2(n29535), .A3(n26975), .ZN(n1575) );
  NOR2_X1 U6798 ( .A1(n715), .A2(n29086), .ZN(n32129) );
  NAND4_X1 U6799 ( .A1(n32131), .A2(n3096), .A3(n32130), .A4(n715), .ZN(n32132) );
  OR2_X2 U6800 ( .A1(n1576), .A2(n17417), .ZN(n24211) );
  AOI21_X1 U6803 ( .B1(n1578), .B2(n13198), .A(n1577), .ZN(n11771) );
  NAND2_X1 U6804 ( .A1(n13198), .A2(n1579), .ZN(n1581) );
  MUX2_X1 U6805 ( .A(n1581), .B(n13199), .S(n13947), .Z(n13212) );
  NAND2_X1 U6806 ( .A1(n36213), .A2(n1582), .ZN(n38988) );
  INV_X1 U6807 ( .A(n52090), .ZN(n48829) );
  NAND3_X1 U6808 ( .A1(n52434), .A2(n48834), .A3(n1585), .ZN(n1584) );
  NAND2_X1 U6810 ( .A1(n36546), .A2(n1587), .ZN(n7990) );
  NAND3_X1 U6811 ( .A1(n7850), .A2(n36539), .A3(n2043), .ZN(n1587) );
  INV_X1 U6812 ( .A(n46568), .ZN(n1590) );
  NAND3_X1 U6813 ( .A1(n1588), .A2(n45144), .A3(n6587), .ZN(n1593) );
  NAND4_X2 U6814 ( .A1(n6589), .A2(n1589), .A3(n1591), .A4(n1593), .ZN(n47620)
         );
  NAND2_X1 U6815 ( .A1(n6586), .A2(n1590), .ZN(n1589) );
  NAND2_X1 U6816 ( .A1(n1592), .A2(n47093), .ZN(n1591) );
  NAND2_X1 U6817 ( .A1(n46566), .A2(n47095), .ZN(n1592) );
  INV_X1 U6818 ( .A(Ciphertext[171]), .ZN(n1594) );
  NAND2_X1 U6819 ( .A1(n20231), .A2(n1596), .ZN(n20233) );
  NAND2_X1 U6820 ( .A1(n1597), .A2(n51090), .ZN(n1596) );
  NAND2_X1 U6822 ( .A1(n26753), .A2(n29542), .ZN(n6337) );
  XNOR2_X2 U6823 ( .A(n26174), .B(n26173), .ZN(n29550) );
  NAND4_X2 U6825 ( .A1(n1602), .A2(n1601), .A3(n46208), .A4(n1600), .ZN(n49037) );
  NAND3_X1 U6826 ( .A1(n42365), .A2(n52079), .A3(n46204), .ZN(n1600) );
  NAND2_X1 U6827 ( .A1(n52079), .A2(n46198), .ZN(n1601) );
  OAI21_X1 U6828 ( .B1(n24248), .B2(n1603), .A(n21815), .ZN(n20282) );
  NAND3_X1 U6831 ( .A1(n24156), .A2(n24157), .A3(n24155), .ZN(n1606) );
  NAND2_X1 U6832 ( .A1(n23828), .A2(n23833), .ZN(n24155) );
  NAND2_X1 U6835 ( .A1(n1610), .A2(n31684), .ZN(n31685) );
  NAND2_X1 U6836 ( .A1(n1610), .A2(n2094), .ZN(n31686) );
  NAND2_X1 U6837 ( .A1(n29966), .A2(n1610), .ZN(n29972) );
  OAI21_X1 U6838 ( .B1(n31694), .B2(n1610), .A(n31693), .ZN(n31695) );
  NAND3_X1 U6839 ( .A1(n35433), .A2(n1612), .A3(n1611), .ZN(n1613) );
  NAND2_X1 U6840 ( .A1(n1614), .A2(n51297), .ZN(n1612) );
  NAND2_X2 U6843 ( .A1(n1615), .A2(n21644), .ZN(n24413) );
  NAND2_X1 U6844 ( .A1(n1616), .A2(n21463), .ZN(n3404) );
  NAND2_X1 U6845 ( .A1(n21449), .A2(n1617), .ZN(n1616) );
  NAND2_X1 U6846 ( .A1(n21474), .A2(n1618), .ZN(n1617) );
  NAND2_X1 U6847 ( .A1(n743), .A2(n51111), .ZN(n27053) );
  NAND4_X1 U6848 ( .A1(n27049), .A2(n743), .A3(n29545), .A4(n51111), .ZN(
        n29552) );
  NAND3_X1 U6849 ( .A1(n8093), .A2(n26752), .A3(n29552), .ZN(n8092) );
  NAND3_X1 U6850 ( .A1(n6469), .A2(n41355), .A3(n41339), .ZN(n41340) );
  NAND2_X1 U6851 ( .A1(n498), .A2(n20230), .ZN(n1621) );
  NAND3_X1 U6852 ( .A1(n18100), .A2(n8302), .A3(n498), .ZN(n16876) );
  NAND3_X1 U6853 ( .A1(n49562), .A2(n49592), .A3(n49598), .ZN(n49602) );
  NAND3_X1 U6854 ( .A1(n4009), .A2(n47360), .A3(n43186), .ZN(n1625) );
  OAI21_X1 U6855 ( .B1(n1626), .B2(n39200), .A(n37880), .ZN(n40940) );
  XNOR2_X1 U6856 ( .A(n516), .B(n1627), .ZN(n40238) );
  XNOR2_X1 U6857 ( .A(n41518), .B(n40224), .ZN(n1628) );
  NAND4_X2 U6858 ( .A1(n1631), .A2(n1629), .A3(n14121), .A4(n1630), .ZN(n16666) );
  NAND2_X1 U6859 ( .A1(n14116), .A2(n15207), .ZN(n1629) );
  NAND3_X1 U6860 ( .A1(n14119), .A2(n14761), .A3(n14118), .ZN(n1630) );
  XNOR2_X2 U6861 ( .A(n15888), .B(n15887), .ZN(n20232) );
  NAND3_X1 U6862 ( .A1(n45777), .A2(n45779), .A3(n1632), .ZN(n45782) );
  NAND2_X1 U6863 ( .A1(n40953), .A2(n41374), .ZN(n1633) );
  NAND2_X1 U6864 ( .A1(n40963), .A2(n41380), .ZN(n40917) );
  NOR2_X1 U6865 ( .A1(n1636), .A2(n1635), .ZN(n3898) );
  OAI21_X1 U6866 ( .B1(n49534), .B2(n49491), .A(n3321), .ZN(n1635) );
  NAND3_X2 U6867 ( .A1(n1841), .A2(n1637), .A3(n3662), .ZN(n32491) );
  NAND2_X1 U6868 ( .A1(n30755), .A2(n51696), .ZN(n1638) );
  NAND2_X1 U6870 ( .A1(n1898), .A2(n30773), .ZN(n1640) );
  NAND3_X1 U6871 ( .A1(n1642), .A2(n1900), .A3(n27556), .ZN(n1641) );
  NAND2_X1 U6872 ( .A1(n1899), .A2(n6048), .ZN(n1642) );
  NAND2_X1 U6873 ( .A1(n48269), .A2(n48264), .ZN(n40175) );
  AND3_X1 U6874 ( .A1(n36117), .A2(n36116), .A3(n36113), .ZN(n1646) );
  NAND2_X1 U6875 ( .A1(n34193), .A2(n38073), .ZN(n34195) );
  NAND2_X1 U6878 ( .A1(n752), .A2(n1647), .ZN(n7831) );
  NAND3_X1 U6879 ( .A1(n23553), .A2(n1648), .A3(n23570), .ZN(n23555) );
  NAND2_X1 U6880 ( .A1(n23361), .A2(n1648), .ZN(n23574) );
  AND3_X2 U6882 ( .A1(n17022), .A2(n5046), .A3(n17023), .ZN(n1648) );
  NAND2_X2 U6883 ( .A1(n1649), .A2(n45935), .ZN(n49443) );
  NOR2_X1 U6884 ( .A1(n1651), .A2(n1650), .ZN(n1649) );
  NAND2_X1 U6885 ( .A1(n45933), .A2(n45665), .ZN(n1650) );
  NAND2_X1 U6886 ( .A1(n45666), .A2(n45934), .ZN(n1651) );
  NAND2_X1 U6887 ( .A1(n45666), .A2(n45665), .ZN(n1653) );
  OR2_X2 U6888 ( .A1(n1652), .A2(n1653), .ZN(n48912) );
  INV_X1 U6890 ( .A(n46635), .ZN(n1654) );
  NAND2_X1 U6891 ( .A1(n45763), .A2(n1655), .ZN(n6742) );
  NOR2_X1 U6892 ( .A1(n45763), .A2(n46637), .ZN(n44422) );
  NAND3_X1 U6893 ( .A1(n44872), .A2(n45761), .A3(n1655), .ZN(n47908) );
  INV_X1 U6894 ( .A(n46637), .ZN(n1655) );
  INV_X1 U6895 ( .A(n23045), .ZN(n1657) );
  NOR2_X1 U6896 ( .A1(n1657), .A2(n23052), .ZN(n22932) );
  NAND3_X1 U6897 ( .A1(n23048), .A2(n23054), .A3(n1657), .ZN(n23058) );
  NAND3_X1 U6899 ( .A1(n22070), .A2(n1656), .A3(n23053), .ZN(n22079) );
  AND2_X1 U6900 ( .A1(n1657), .A2(n23048), .ZN(n1656) );
  XNOR2_X1 U6901 ( .A(n27378), .B(n27371), .ZN(n1658) );
  OAI211_X1 U6902 ( .C1(n17021), .C2(n20122), .A(n1659), .B(n20125), .ZN(n5974) );
  NAND2_X1 U6903 ( .A1(n51126), .A2(n17021), .ZN(n1659) );
  NOR2_X1 U6906 ( .A1(n4246), .A2(n1661), .ZN(n36561) );
  NOR2_X1 U6907 ( .A1(n36559), .A2(n1661), .ZN(n35320) );
  NAND2_X1 U6908 ( .A1(n36493), .A2(n36015), .ZN(n1661) );
  NAND2_X1 U6910 ( .A1(n44655), .A2(n46635), .ZN(n1662) );
  NAND4_X2 U6912 ( .A1(n1665), .A2(n2910), .A3(n11040), .A4(n1666), .ZN(n14345) );
  OAI21_X1 U6913 ( .B1(n41063), .B2(n41058), .A(n41049), .ZN(n1667) );
  NAND2_X1 U6915 ( .A1(n41049), .A2(n41058), .ZN(n40512) );
  INV_X1 U6916 ( .A(n39603), .ZN(n40505) );
  NAND2_X1 U6917 ( .A1(n1668), .A2(n39604), .ZN(n39607) );
  INV_X2 U6919 ( .A(n49511), .ZN(n49522) );
  NAND2_X1 U6920 ( .A1(n48168), .A2(n48167), .ZN(n1753) );
  NAND4_X2 U6924 ( .A1(n39491), .A2(n39490), .A3(n39489), .A4(n1669), .ZN(
        n42020) );
  NAND2_X1 U6925 ( .A1(n1670), .A2(n39488), .ZN(n1669) );
  AND2_X1 U6926 ( .A1(n39471), .A2(n39484), .ZN(n1670) );
  NAND4_X2 U6927 ( .A1(n17051), .A2(n1671), .A3(n17048), .A4(n17052), .ZN(
        n23546) );
  NAND2_X1 U6929 ( .A1(n18381), .A2(n7920), .ZN(n17045) );
  XNOR2_X1 U6930 ( .A(n45279), .B(n1673), .ZN(n45280) );
  XNOR2_X1 U6931 ( .A(n1673), .B(n45059), .ZN(n44895) );
  NAND2_X1 U6932 ( .A1(n1839), .A2(n1675), .ZN(n1678) );
  NOR2_X1 U6933 ( .A1(n26761), .A2(n29563), .ZN(n2845) );
  INV_X1 U6934 ( .A(n29545), .ZN(n1680) );
  AOI21_X1 U6935 ( .B1(n2028), .B2(n6107), .A(n1681), .ZN(n2026) );
  NAND3_X1 U6936 ( .A1(n2027), .A2(n31826), .A3(n1682), .ZN(n1681) );
  INV_X1 U6937 ( .A(n1682), .ZN(n29382) );
  INV_X1 U6938 ( .A(n31712), .ZN(n1683) );
  INV_X2 U6939 ( .A(n1685), .ZN(n31711) );
  NAND2_X1 U6940 ( .A1(n1685), .A2(n32130), .ZN(n29976) );
  NAND2_X1 U6941 ( .A1(n1685), .A2(n26203), .ZN(n29085) );
  NAND2_X1 U6942 ( .A1(n31700), .A2(n1685), .ZN(n31709) );
  NAND2_X1 U6943 ( .A1(n1683), .A2(n31711), .ZN(n32118) );
  NAND2_X1 U6944 ( .A1(n31701), .A2(n1685), .ZN(n26350) );
  AND2_X1 U6945 ( .A1(n1685), .A2(n32128), .ZN(n1684) );
  NAND3_X1 U6946 ( .A1(n20043), .A2(n16823), .A3(n20042), .ZN(n1696) );
  AND2_X1 U6947 ( .A1(n18376), .A2(n20037), .ZN(n20042) );
  XNOR2_X2 U6948 ( .A(n16329), .B(n779), .ZN(n18376) );
  NAND2_X1 U6949 ( .A1(n1688), .A2(n1687), .ZN(n1686) );
  OR3_X1 U6950 ( .A1(n24267), .A2(n24266), .A3(n24268), .ZN(n1688) );
  OAI21_X1 U6951 ( .B1(n31898), .B2(n31413), .A(n1689), .ZN(n31900) );
  OAI21_X1 U6952 ( .B1(n1690), .B2(n31424), .A(n31413), .ZN(n1689) );
  NAND2_X1 U6953 ( .A1(n29991), .A2(n29992), .ZN(n31424) );
  INV_X1 U6954 ( .A(n2609), .ZN(n1690) );
  NAND2_X1 U6955 ( .A1(n36590), .A2(n36454), .ZN(n36586) );
  NAND2_X1 U6956 ( .A1(n625), .A2(n1693), .ZN(n29220) );
  NAND2_X1 U6957 ( .A1(n41977), .A2(n41978), .ZN(n41980) );
  NAND3_X1 U6960 ( .A1(n1696), .A2(n20047), .A3(n1695), .ZN(n20048) );
  NAND3_X1 U6961 ( .A1(n20046), .A2(n5881), .A3(n20045), .ZN(n1695) );
  INV_X1 U6962 ( .A(n18376), .ZN(n7920) );
  NAND2_X1 U6963 ( .A1(n34910), .A2(n1697), .ZN(n7634) );
  NAND3_X1 U6964 ( .A1(n38999), .A2(n38998), .A3(n39393), .ZN(n1697) );
  NAND2_X1 U6965 ( .A1(n31215), .A2(n6969), .ZN(n1701) );
  NAND2_X1 U6966 ( .A1(n32215), .A2(n32211), .ZN(n31215) );
  MUX2_X1 U6968 ( .A(n32211), .B(n32210), .S(n50981), .Z(n1702) );
  NAND2_X1 U6973 ( .A1(n21664), .A2(n1704), .ZN(n21646) );
  NAND2_X1 U6974 ( .A1(n52271), .A2(n20656), .ZN(n20660) );
  AOI22_X1 U6975 ( .A1(n21653), .A2(n52186), .B1(n21654), .B2(n1704), .ZN(
        n21667) );
  NAND2_X1 U6977 ( .A1(n30106), .A2(n3767), .ZN(n30993) );
  NOR3_X1 U6979 ( .A1(n29221), .A2(n30269), .A3(n1708), .ZN(n1707) );
  INV_X1 U6980 ( .A(n5564), .ZN(n1708) );
  OR2_X1 U6981 ( .A1(n1710), .A2(n1709), .ZN(n24453) );
  NAND2_X1 U6982 ( .A1(n24452), .A2(n49387), .ZN(n1709) );
  NAND2_X1 U6983 ( .A1(n772), .A2(n1715), .ZN(n18060) );
  NAND2_X1 U6984 ( .A1(n1715), .A2(n14381), .ZN(n18059) );
  NAND3_X1 U6985 ( .A1(n17440), .A2(n17553), .A3(n1715), .ZN(n17435) );
  NAND2_X1 U6986 ( .A1(n17541), .A2(n1713), .ZN(n17430) );
  NAND2_X1 U6987 ( .A1(n44828), .A2(n1719), .ZN(n1716) );
  NAND2_X1 U6988 ( .A1(n44703), .A2(n44702), .ZN(n1721) );
  XNOR2_X1 U6989 ( .A(n7387), .B(n43352), .ZN(n41370) );
  XNOR2_X2 U6990 ( .A(n52122), .B(n44374), .ZN(n43352) );
  NAND3_X1 U6992 ( .A1(n48812), .A2(n5391), .A3(n5392), .ZN(n1726) );
  INV_X1 U6993 ( .A(n1734), .ZN(n1727) );
  NAND2_X1 U6995 ( .A1(n1733), .A2(n45755), .ZN(n1732) );
  NOR2_X1 U6996 ( .A1(n45743), .A2(n48808), .ZN(n48827) );
  OAI21_X1 U6997 ( .B1(n45742), .B2(n48834), .A(n45741), .ZN(n1736) );
  NAND2_X1 U6998 ( .A1(n31273), .A2(n30104), .ZN(n1738) );
  OR2_X1 U6999 ( .A1(n31484), .A2(n31490), .ZN(n30104) );
  NAND2_X1 U7002 ( .A1(n24243), .A2(n1744), .ZN(n23789) );
  XNOR2_X1 U7003 ( .A(n1747), .B(n48358), .ZN(Plaintext[51]) );
  NAND4_X1 U7004 ( .A1(n1748), .A2(n48355), .A3(n1750), .A4(n48357), .ZN(n1747) );
  AND2_X1 U7005 ( .A1(n1749), .A2(n48356), .ZN(n1748) );
  NAND2_X1 U7006 ( .A1(n48364), .A2(n48359), .ZN(n1749) );
  OAI21_X1 U7007 ( .B1(n1753), .B2(n1752), .A(n1755), .ZN(n1751) );
  NAND2_X1 U7008 ( .A1(n48170), .A2(n48411), .ZN(n1754) );
  INV_X1 U7009 ( .A(n48411), .ZN(n1755) );
  NAND2_X1 U7011 ( .A1(n50949), .A2(n1757), .ZN(n50932) );
  AOI21_X1 U7012 ( .B1(n47390), .B2(n1757), .A(n1756), .ZN(n47394) );
  NAND2_X1 U7014 ( .A1(n46744), .A2(n1759), .ZN(n1758) );
  INV_X1 U7015 ( .A(n46753), .ZN(n1759) );
  NAND3_X1 U7016 ( .A1(n45800), .A2(n46737), .A3(n1760), .ZN(n44857) );
  INV_X1 U7017 ( .A(n46744), .ZN(n1760) );
  NAND2_X1 U7018 ( .A1(n32042), .A2(n31323), .ZN(n1761) );
  NAND2_X1 U7019 ( .A1(n32455), .A2(n723), .ZN(n1762) );
  INV_X1 U7020 ( .A(n20432), .ZN(n1763) );
  NAND2_X1 U7021 ( .A1(n1766), .A2(n1765), .ZN(n31525) );
  NAND2_X1 U7022 ( .A1(n31514), .A2(n31513), .ZN(n1765) );
  NAND2_X1 U7023 ( .A1(n1768), .A2(n1767), .ZN(n1766) );
  NAND2_X1 U7024 ( .A1(n7183), .A2(n31511), .ZN(n1768) );
  NAND2_X1 U7025 ( .A1(n1770), .A2(n1769), .ZN(n32013) );
  OAI211_X1 U7026 ( .C1(n31988), .C2(n32509), .A(n30873), .B(n31987), .ZN(
        n1769) );
  NAND2_X1 U7027 ( .A1(n7897), .A2(n31986), .ZN(n31989) );
  NAND2_X1 U7028 ( .A1(n1772), .A2(n51023), .ZN(n9273) );
  NAND2_X1 U7029 ( .A1(n1773), .A2(n15424), .ZN(n1772) );
  INV_X1 U7030 ( .A(n15417), .ZN(n1773) );
  NAND2_X1 U7031 ( .A1(n1774), .A2(n23241), .ZN(n23251) );
  NOR2_X1 U7032 ( .A1(n22653), .A2(n1777), .ZN(n23261) );
  OAI21_X1 U7033 ( .B1(n22658), .B2(n1777), .A(n23241), .ZN(n20930) );
  NOR2_X1 U7034 ( .A1(n23247), .A2(n757), .ZN(n1775) );
  NAND2_X1 U7035 ( .A1(n21848), .A2(n1776), .ZN(n21856) );
  XNOR2_X1 U7036 ( .A(n1778), .B(n52100), .ZN(n24404) );
  XNOR2_X1 U7037 ( .A(n26274), .B(n1778), .ZN(n26276) );
  XNOR2_X1 U7038 ( .A(n24215), .B(n1778), .ZN(n24216) );
  NAND2_X1 U7040 ( .A1(n22289), .A2(n20943), .ZN(n1779) );
  NAND2_X1 U7041 ( .A1(n3553), .A2(n51694), .ZN(n22289) );
  NAND2_X1 U7042 ( .A1(n15263), .A2(n51686), .ZN(n1780) );
  NAND2_X1 U7043 ( .A1(n12441), .A2(n12710), .ZN(n1781) );
  NAND2_X1 U7044 ( .A1(n1784), .A2(n1783), .ZN(n8313) );
  INV_X1 U7045 ( .A(n12711), .ZN(n1783) );
  NAND2_X1 U7046 ( .A1(n17496), .A2(n1785), .ZN(n8159) );
  NAND2_X1 U7048 ( .A1(n1788), .A2(n1789), .ZN(n14741) );
  NAND3_X1 U7050 ( .A1(n4098), .A2(n20476), .A3(n1789), .ZN(n17635) );
  NAND3_X1 U7051 ( .A1(n12403), .A2(n7865), .A3(n13291), .ZN(n13737) );
  NAND4_X2 U7052 ( .A1(n1790), .A2(n1791), .A3(n10953), .A4(n1792), .ZN(n13291) );
  NAND3_X1 U7053 ( .A1(n10950), .A2(n10949), .A3(n12317), .ZN(n1791) );
  XNOR2_X1 U7054 ( .A(n1793), .B(n18595), .ZN(n18606) );
  XNOR2_X1 U7055 ( .A(n1794), .B(n18594), .ZN(n1793) );
  XNOR2_X1 U7056 ( .A(n1795), .B(n19266), .ZN(n1794) );
  XNOR2_X1 U7057 ( .A(n18600), .B(n18601), .ZN(n1795) );
  NAND2_X1 U7058 ( .A1(n3493), .A2(n21425), .ZN(n1796) );
  OAI22_X1 U7059 ( .A1(n1797), .A2(n21427), .B1(n21442), .B2(n19957), .ZN(
        n19158) );
  NAND2_X1 U7060 ( .A1(n1800), .A2(n1799), .ZN(n1798) );
  INV_X1 U7061 ( .A(n45204), .ZN(n1799) );
  NOR2_X1 U7062 ( .A1(n45621), .A2(n883), .ZN(n1800) );
  XNOR2_X1 U7064 ( .A(n25017), .B(n51122), .ZN(n25018) );
  NAND3_X1 U7066 ( .A1(n27545), .A2(n1804), .A3(n1803), .ZN(n27546) );
  INV_X1 U7067 ( .A(n26722), .ZN(n29441) );
  AOI21_X1 U7069 ( .B1(n29440), .B2(n29441), .A(n1805), .ZN(n29452) );
  AND2_X1 U7070 ( .A1(n2726), .A2(n49663), .ZN(n49671) );
  AND2_X1 U7071 ( .A1(n49651), .A2(n51733), .ZN(n50021) );
  INV_X1 U7073 ( .A(n19359), .ZN(n21464) );
  NOR2_X1 U7075 ( .A1(n5153), .A2(n36383), .ZN(n36379) );
  NAND2_X1 U7077 ( .A1(n1807), .A2(n33463), .ZN(n33466) );
  NOR2_X1 U7078 ( .A1(n1807), .A2(n42057), .ZN(n42058) );
  NAND2_X1 U7079 ( .A1(n1808), .A2(n50001), .ZN(n1813) );
  NAND2_X1 U7080 ( .A1(n46005), .A2(n1809), .ZN(n1808) );
  NAND2_X1 U7081 ( .A1(n47371), .A2(n6172), .ZN(n1809) );
  NAND2_X1 U7082 ( .A1(n50314), .A2(n6172), .ZN(n50001) );
  AOI21_X1 U7083 ( .B1(n1813), .B2(n1810), .A(n50325), .ZN(n46012) );
  OAI211_X1 U7084 ( .C1(n47371), .C2(n1812), .A(n1811), .B(n52224), .ZN(n1810)
         );
  INV_X1 U7085 ( .A(n50010), .ZN(n1812) );
  NAND2_X1 U7086 ( .A1(n50008), .A2(n51526), .ZN(n47371) );
  NAND2_X1 U7087 ( .A1(n1815), .A2(n1817), .ZN(n1814) );
  NAND2_X1 U7088 ( .A1(n29321), .A2(n27890), .ZN(n1815) );
  OAI21_X1 U7092 ( .B1(n49903), .B2(n49933), .A(n49932), .ZN(n1819) );
  XNOR2_X1 U7093 ( .A(n1818), .B(n49898), .ZN(Plaintext[134]) );
  NAND4_X1 U7094 ( .A1(n49897), .A2(n1821), .A3(n49896), .A4(n1819), .ZN(n1818) );
  NAND2_X1 U7095 ( .A1(n49917), .A2(n49899), .ZN(n49890) );
  NAND2_X1 U7096 ( .A1(n49917), .A2(n1820), .ZN(n1821) );
  OR3_X1 U7097 ( .A1(n41144), .A2(n1822), .A3(n682), .ZN(n5486) );
  NOR2_X1 U7100 ( .A1(n25847), .A2(n1823), .ZN(n25987) );
  NOR2_X1 U7101 ( .A1(n7200), .A2(n1823), .ZN(n5044) );
  NAND3_X1 U7102 ( .A1(n10169), .A2(n11023), .A3(n580), .ZN(n1824) );
  NAND2_X1 U7103 ( .A1(n10584), .A2(n10579), .ZN(n10169) );
  NAND2_X1 U7104 ( .A1(n11030), .A2(n10584), .ZN(n10170) );
  NAND2_X1 U7105 ( .A1(n11037), .A2(n790), .ZN(n1826) );
  XNOR2_X2 U7106 ( .A(n25601), .B(n25602), .ZN(n29260) );
  AND3_X1 U7107 ( .A1(n1828), .A2(n30234), .A3(n4775), .ZN(n25630) );
  NAND2_X1 U7108 ( .A1(n27938), .A2(n29248), .ZN(n1828) );
  NAND2_X1 U7109 ( .A1(n36521), .A2(n36522), .ZN(n2916) );
  AND2_X1 U7111 ( .A1(n24476), .A2(n24477), .ZN(n1830) );
  NAND3_X1 U7112 ( .A1(n24475), .A2(n24478), .A3(n1830), .ZN(n31301) );
  NAND2_X1 U7113 ( .A1(n29650), .A2(n31302), .ZN(n29398) );
  NAND2_X1 U7114 ( .A1(n51085), .A2(n30647), .ZN(n29650) );
  INV_X1 U7116 ( .A(n16490), .ZN(n1835) );
  NAND2_X1 U7118 ( .A1(n1839), .A2(n6048), .ZN(n6191) );
  NAND2_X1 U7119 ( .A1(n1838), .A2(n1837), .ZN(n26844) );
  NAND2_X1 U7120 ( .A1(n1839), .A2(n30768), .ZN(n1837) );
  NAND2_X1 U7121 ( .A1(n26841), .A2(n730), .ZN(n1838) );
  NAND2_X1 U7122 ( .A1(n32486), .A2(n1840), .ZN(n32021) );
  AND2_X1 U7123 ( .A1(n1841), .A2(n32019), .ZN(n1840) );
  NAND3_X1 U7124 ( .A1(n1842), .A2(n39449), .A3(n39441), .ZN(n7373) );
  NAND2_X1 U7125 ( .A1(n37722), .A2(n2465), .ZN(n1842) );
  NAND2_X1 U7126 ( .A1(n39035), .A2(n34806), .ZN(n37722) );
  NAND2_X1 U7127 ( .A1(n34806), .A2(n1843), .ZN(n39449) );
  NAND4_X1 U7129 ( .A1(n1846), .A2(n11159), .A3(n13089), .A4(n13086), .ZN(
        n1845) );
  NAND2_X1 U7130 ( .A1(n12919), .A2(n13095), .ZN(n1846) );
  NAND2_X1 U7131 ( .A1(n27688), .A2(n6092), .ZN(n27575) );
  NAND2_X1 U7132 ( .A1(n27677), .A2(n26823), .ZN(n6092) );
  NAND2_X1 U7133 ( .A1(n31497), .A2(n31269), .ZN(n31266) );
  NAND2_X1 U7134 ( .A1(n1847), .A2(n25055), .ZN(n25052) );
  NAND2_X1 U7135 ( .A1(n1847), .A2(n3728), .ZN(n25060) );
  OAI21_X1 U7136 ( .B1(n9558), .B2(n1850), .A(n9557), .ZN(n1849) );
  NAND2_X1 U7137 ( .A1(n2227), .A2(n12659), .ZN(n12657) );
  NAND2_X1 U7138 ( .A1(n2227), .A2(n1848), .ZN(n1850) );
  NAND2_X1 U7139 ( .A1(n32080), .A2(n31286), .ZN(n33157) );
  NAND2_X1 U7140 ( .A1(n20409), .A2(n21397), .ZN(n1856) );
  AND2_X1 U7141 ( .A1(n22470), .A2(n22481), .ZN(n22478) );
  NAND2_X1 U7142 ( .A1(n20410), .A2(n769), .ZN(n1858) );
  NOR2_X1 U7143 ( .A1(n1860), .A2(n581), .ZN(n1861) );
  NOR2_X1 U7145 ( .A1(n32509), .A2(n32511), .ZN(n32007) );
  NAND3_X1 U7147 ( .A1(n28561), .A2(n28557), .A3(n28563), .ZN(n1862) );
  OAI21_X1 U7148 ( .B1(n27116), .B2(n27115), .A(n27114), .ZN(n1863) );
  INV_X1 U7150 ( .A(n12651), .ZN(n10456) );
  NAND2_X1 U7151 ( .A1(n1865), .A2(n38173), .ZN(n1864) );
  NAND2_X1 U7152 ( .A1(n39836), .A2(n39834), .ZN(n39830) );
  NAND2_X1 U7153 ( .A1(n38024), .A2(n34976), .ZN(n1865) );
  AND2_X1 U7154 ( .A1(n12693), .A2(n1866), .ZN(n1867) );
  NAND2_X1 U7155 ( .A1(n7781), .A2(n1868), .ZN(n1866) );
  OAI211_X1 U7156 ( .C1(n12694), .C2(n12708), .A(n1867), .B(n12689), .ZN(n2585) );
  NAND2_X1 U7157 ( .A1(n735), .A2(n30191), .ZN(n27092) );
  XNOR2_X2 U7159 ( .A(n25335), .B(n25334), .ZN(n30191) );
  XNOR2_X2 U7160 ( .A(n33722), .B(n1872), .ZN(n34572) );
  OR2_X2 U7161 ( .A1(n5302), .A2(n5301), .ZN(n1872) );
  XNOR2_X1 U7162 ( .A(n1872), .B(n35536), .ZN(n34040) );
  XNOR2_X1 U7163 ( .A(n35345), .B(n1872), .ZN(n35346) );
  XNOR2_X1 U7164 ( .A(n37081), .B(n1872), .ZN(n37088) );
  XNOR2_X1 U7165 ( .A(n35800), .B(n1872), .ZN(n33109) );
  XNOR2_X1 U7166 ( .A(n35534), .B(n1872), .ZN(n33958) );
  NOR2_X1 U7167 ( .A1(n1873), .A2(n13735), .ZN(n13738) );
  INV_X1 U7168 ( .A(n13734), .ZN(n1873) );
  OR2_X2 U7170 ( .A1(n14752), .A2(n14751), .ZN(n22287) );
  NAND2_X1 U7174 ( .A1(n39907), .A2(n1874), .ZN(n38436) );
  INV_X2 U7175 ( .A(n3506), .ZN(n23417) );
  NOR2_X1 U7176 ( .A1(n20888), .A2(n23420), .ZN(n22045) );
  XNOR2_X1 U7177 ( .A(n52141), .B(n1878), .ZN(n17171) );
  XNOR2_X1 U7178 ( .A(n51379), .B(n1878), .ZN(n18459) );
  NAND3_X1 U7179 ( .A1(n51308), .A2(n49363), .A3(n523), .ZN(n49329) );
  MUX2_X1 U7180 ( .A(n49382), .B(n49371), .S(n51308), .Z(n49322) );
  NAND2_X1 U7181 ( .A1(n1879), .A2(n49305), .ZN(n4903) );
  NAND2_X1 U7182 ( .A1(n49294), .A2(n1879), .ZN(n49301) );
  NOR2_X1 U7184 ( .A1(n2158), .A2(n30267), .ZN(n30257) );
  NAND2_X1 U7185 ( .A1(n4476), .A2(n4475), .ZN(n1881) );
  OAI21_X1 U7186 ( .B1(n6190), .B2(n30762), .A(n30761), .ZN(n1882) );
  NAND2_X1 U7187 ( .A1(n40596), .A2(n40775), .ZN(n1883) );
  NAND2_X1 U7188 ( .A1(n39801), .A2(n6046), .ZN(n40590) );
  XNOR2_X1 U7189 ( .A(n1885), .B(n35404), .ZN(n1887) );
  XNOR2_X1 U7190 ( .A(n701), .B(n35680), .ZN(n1885) );
  XNOR2_X1 U7193 ( .A(n34796), .B(n1889), .ZN(n1888) );
  XNOR2_X1 U7194 ( .A(n34788), .B(n35278), .ZN(n1889) );
  NAND2_X1 U7195 ( .A1(n18024), .A2(n19395), .ZN(n1891) );
  NAND3_X1 U7196 ( .A1(n18024), .A2(n19395), .A3(n764), .ZN(n18027) );
  OAI211_X1 U7197 ( .C1(n19390), .C2(n19400), .A(n19389), .B(n1891), .ZN(
        n18028) );
  XNOR2_X2 U7198 ( .A(n1894), .B(n1892), .ZN(n36141) );
  XNOR2_X1 U7199 ( .A(n35474), .B(n31351), .ZN(n1894) );
  OAI21_X1 U7200 ( .B1(n13979), .B2(n13583), .A(n12198), .ZN(n12199) );
  NAND3_X1 U7201 ( .A1(n13583), .A2(n12204), .A3(n12198), .ZN(n1895) );
  NAND2_X1 U7202 ( .A1(n13577), .A2(n1895), .ZN(n12200) );
  XNOR2_X2 U7203 ( .A(n1897), .B(n1896), .ZN(n19388) );
  XNOR2_X1 U7204 ( .A(n51133), .B(n12402), .ZN(n16360) );
  XNOR2_X1 U7205 ( .A(n12879), .B(n17268), .ZN(n1897) );
  NAND2_X1 U7206 ( .A1(n3623), .A2(n32638), .ZN(n5304) );
  NAND2_X1 U7208 ( .A1(n32540), .A2(n32633), .ZN(n32912) );
  INV_X1 U7211 ( .A(n30773), .ZN(n27557) );
  INV_X1 U7212 ( .A(n30772), .ZN(n27555) );
  NAND2_X1 U7213 ( .A1(n27554), .A2(n30757), .ZN(n1901) );
  NAND2_X1 U7214 ( .A1(n1902), .A2(n47777), .ZN(n45011) );
  NAND2_X1 U7215 ( .A1(n47712), .A2(n645), .ZN(n47747) );
  INV_X1 U7216 ( .A(n1902), .ZN(n47712) );
  AOI21_X1 U7217 ( .B1(n47781), .B2(n47782), .A(n1902), .ZN(n47783) );
  OAI21_X1 U7218 ( .B1(n47755), .B2(n1902), .A(n45877), .ZN(n47756) );
  NAND2_X1 U7219 ( .A1(n47732), .A2(n1902), .ZN(n47733) );
  NAND4_X1 U7221 ( .A1(n21837), .A2(n22125), .A3(n1904), .A4(n1903), .ZN(
        n21841) );
  NAND2_X1 U7222 ( .A1(n23238), .A2(n22129), .ZN(n22124) );
  INV_X2 U7223 ( .A(n30699), .ZN(n30392) );
  NAND2_X1 U7225 ( .A1(n1906), .A2(n30392), .ZN(n1905) );
  NAND3_X1 U7226 ( .A1(n734), .A2(n30392), .A3(n30389), .ZN(n30386) );
  AND2_X1 U7227 ( .A1(n13786), .A2(n12418), .ZN(n1911) );
  NAND3_X1 U7230 ( .A1(n1910), .A2(n1911), .A3(n13185), .ZN(n1908) );
  NOR2_X1 U7231 ( .A1(n1913), .A2(n1909), .ZN(n1912) );
  NAND2_X1 U7232 ( .A1(n12413), .A2(n13288), .ZN(n1913) );
  NAND2_X1 U7233 ( .A1(n36034), .A2(n37957), .ZN(n1914) );
  NAND2_X1 U7234 ( .A1(n6219), .A2(n1915), .ZN(n37970) );
  NOR2_X1 U7235 ( .A1(n36037), .A2(n699), .ZN(n1915) );
  INV_X2 U7238 ( .A(n6930), .ZN(n23446) );
  NAND2_X1 U7240 ( .A1(n46339), .A2(n48417), .ZN(n1918) );
  NAND2_X1 U7241 ( .A1(n46334), .A2(n46333), .ZN(n1919) );
  NOR2_X1 U7242 ( .A1(n52067), .A2(n48751), .ZN(n48745) );
  NAND2_X1 U7243 ( .A1(n45744), .A2(n1920), .ZN(n8340) );
  NAND2_X1 U7244 ( .A1(n1921), .A2(n32243), .ZN(n24367) );
  NAND2_X1 U7245 ( .A1(n1921), .A2(n30839), .ZN(n30845) );
  NOR2_X1 U7246 ( .A1(n32233), .A2(n32251), .ZN(n1921) );
  NAND2_X1 U7247 ( .A1(n47160), .A2(n2752), .ZN(n1924) );
  NAND2_X1 U7250 ( .A1(n1924), .A2(n43683), .ZN(n1923) );
  INV_X1 U7251 ( .A(n36449), .ZN(n36448) );
  NAND2_X1 U7252 ( .A1(n36595), .A2(n36050), .ZN(n36449) );
  XNOR2_X2 U7253 ( .A(n34390), .B(n34389), .ZN(n36045) );
  XNOR2_X1 U7255 ( .A(n1925), .B(n46143), .ZN(n41755) );
  XNOR2_X1 U7256 ( .A(n40408), .B(n1925), .ZN(n44170) );
  XNOR2_X1 U7257 ( .A(n42459), .B(n52166), .ZN(n42469) );
  XNOR2_X1 U7258 ( .A(n42764), .B(n52166), .ZN(n44364) );
  XNOR2_X1 U7259 ( .A(n52166), .B(n43819), .ZN(n43825) );
  OAI21_X1 U7260 ( .B1(n30452), .B2(n427), .A(n1926), .ZN(n28838) );
  OAI21_X1 U7261 ( .B1(n30456), .B2(n30462), .A(n1927), .ZN(n30464) );
  NAND3_X1 U7262 ( .A1(n42050), .A2(n41487), .A3(n42048), .ZN(n41488) );
  NAND2_X1 U7264 ( .A1(n31454), .A2(n31544), .ZN(n31450) );
  NAND2_X1 U7266 ( .A1(n1928), .A2(n31712), .ZN(n29090) );
  NAND3_X1 U7267 ( .A1(n29089), .A2(n6678), .A3(n29975), .ZN(n1928) );
  NAND2_X1 U7268 ( .A1(n31711), .A2(n30814), .ZN(n29975) );
  NOR2_X1 U7269 ( .A1(n12821), .A2(n13090), .ZN(n1929) );
  NAND2_X1 U7270 ( .A1(n40379), .A2(n677), .ZN(n38615) );
  AOI21_X1 U7271 ( .B1(n38086), .B2(n695), .A(n34189), .ZN(n33271) );
  AOI22_X1 U7272 ( .A1(n9485), .A2(n1932), .B1(n9484), .B2(n10095), .ZN(n9488)
         );
  NOR2_X1 U7273 ( .A1(n1933), .A2(n48778), .ZN(n48784) );
  NAND2_X1 U7274 ( .A1(n1935), .A2(n1934), .ZN(n32466) );
  AOI22_X1 U7275 ( .A1(n32465), .A2(n32716), .B1(n32724), .B2(n32725), .ZN(
        n1934) );
  NAND2_X1 U7276 ( .A1(n1936), .A2(n32724), .ZN(n1935) );
  NAND2_X1 U7277 ( .A1(n29922), .A2(n30755), .ZN(n1937) );
  OAI21_X1 U7278 ( .B1(n1939), .B2(n26842), .A(n29917), .ZN(n1938) );
  OAI21_X1 U7279 ( .B1(n1942), .B2(n1940), .A(n23828), .ZN(n20585) );
  INV_X1 U7280 ( .A(n24157), .ZN(n1941) );
  INV_X1 U7281 ( .A(n23821), .ZN(n1942) );
  INV_X1 U7282 ( .A(n6194), .ZN(n1943) );
  AND2_X1 U7283 ( .A1(n6194), .A2(n1944), .ZN(n46335) );
  NAND2_X1 U7284 ( .A1(n51068), .A2(n48412), .ZN(n1944) );
  NAND2_X1 U7285 ( .A1(n48516), .A2(n48517), .ZN(n1945) );
  NAND3_X2 U7286 ( .A1(n315), .A2(n48564), .A3(n1945), .ZN(n48604) );
  NAND3_X1 U7287 ( .A1(n48648), .A2(n48600), .A3(n48649), .ZN(n3468) );
  XNOR2_X1 U7288 ( .A(n1946), .B(n46112), .ZN(n42587) );
  XNOR2_X1 U7289 ( .A(n44878), .B(n1946), .ZN(n44230) );
  XNOR2_X1 U7290 ( .A(n43143), .B(n1946), .ZN(n45418) );
  XNOR2_X1 U7291 ( .A(n42728), .B(n52069), .ZN(n42733) );
  XNOR2_X1 U7292 ( .A(n42224), .B(n52069), .ZN(n42414) );
  NAND2_X1 U7295 ( .A1(n14331), .A2(n14344), .ZN(n3515) );
  NAND4_X2 U7296 ( .A1(n36221), .A2(n36220), .A3(n1949), .A4(n36219), .ZN(
        n42062) );
  INV_X1 U7297 ( .A(n38477), .ZN(n1950) );
  OAI21_X1 U7298 ( .B1(n36114), .B2(n38477), .A(n1951), .ZN(n36117) );
  INV_X1 U7299 ( .A(n38484), .ZN(n1951) );
  OR2_X2 U7300 ( .A1(n6317), .A2(n35103), .ZN(n38484) );
  AND2_X1 U7301 ( .A1(n50951), .A2(n50913), .ZN(n47391) );
  NOR3_X1 U7303 ( .A1(n12657), .A2(n1953), .A3(n1952), .ZN(n9193) );
  NAND2_X1 U7304 ( .A1(n11986), .A2(n9188), .ZN(n1952) );
  INV_X1 U7305 ( .A(n10444), .ZN(n1953) );
  NAND3_X1 U7306 ( .A1(n20535), .A2(n22699), .A3(n1957), .ZN(n1956) );
  NAND2_X1 U7307 ( .A1(n51694), .A2(n3017), .ZN(n1957) );
  NAND3_X1 U7308 ( .A1(n2884), .A2(n21114), .A3(n20532), .ZN(n1959) );
  XNOR2_X1 U7309 ( .A(n14213), .B(n14212), .ZN(n1960) );
  XNOR2_X2 U7310 ( .A(n1960), .B(n15618), .ZN(n18331) );
  AND2_X1 U7311 ( .A1(n17546), .A2(n17545), .ZN(n18065) );
  NAND2_X1 U7313 ( .A1(n14140), .A2(n1963), .ZN(n1962) );
  OR2_X1 U7314 ( .A1(n30272), .A2(n30268), .ZN(n1964) );
  OAI21_X1 U7315 ( .B1(n21702), .B2(n463), .A(n22184), .ZN(n1968) );
  NAND2_X1 U7316 ( .A1(n21706), .A2(n21705), .ZN(n1965) );
  NAND3_X1 U7317 ( .A1(n21704), .A2(n21703), .A3(n1967), .ZN(n1966) );
  NAND2_X1 U7318 ( .A1(n21106), .A2(n21712), .ZN(n21703) );
  INV_X1 U7319 ( .A(n1970), .ZN(n37809) );
  XNOR2_X1 U7320 ( .A(n1969), .B(n33851), .ZN(n1970) );
  XNOR2_X1 U7321 ( .A(n33852), .B(n34102), .ZN(n1969) );
  NOR2_X1 U7322 ( .A1(n1972), .A2(n1971), .ZN(n2031) );
  OAI21_X1 U7323 ( .B1(n45208), .B2(n45207), .A(n45206), .ZN(n1971) );
  NAND4_X1 U7325 ( .A1(n1974), .A2(n38485), .A3(n38467), .A4(n38464), .ZN(
        n35441) );
  NAND2_X1 U7326 ( .A1(n13030), .A2(n13701), .ZN(n1975) );
  NAND2_X1 U7327 ( .A1(n1975), .A2(n15131), .ZN(n15129) );
  NAND4_X1 U7328 ( .A1(n13695), .A2(n1975), .A3(n5347), .A4(n13696), .ZN(
        n13707) );
  AOI22_X1 U7329 ( .A1(n13695), .A2(n1975), .B1(n2766), .B2(n15132), .ZN(n2765) );
  NAND2_X1 U7330 ( .A1(n49607), .A2(n49556), .ZN(n1976) );
  NAND2_X1 U7332 ( .A1(n6139), .A2(n6140), .ZN(n1977) );
  NAND2_X1 U7333 ( .A1(n22342), .A2(n22343), .ZN(n1978) );
  NAND2_X1 U7334 ( .A1(n1979), .A2(n23663), .ZN(n24360) );
  NAND3_X1 U7335 ( .A1(n23661), .A2(n23662), .A3(n30792), .ZN(n1979) );
  OAI211_X1 U7336 ( .C1(n28740), .C2(n1983), .A(n29861), .B(n1980), .ZN(n28741) );
  NAND2_X1 U7337 ( .A1(n29869), .A2(n28745), .ZN(n1980) );
  MUX2_X1 U7338 ( .A(n30425), .B(n29867), .S(n486), .Z(n27515) );
  NAND3_X1 U7339 ( .A1(n29700), .A2(n29863), .A3(n1983), .ZN(n6055) );
  NAND2_X1 U7342 ( .A1(n8404), .A2(n1985), .ZN(n1987) );
  NAND3_X1 U7343 ( .A1(n32331), .A2(n32332), .A3(n32704), .ZN(n1985) );
  NAND2_X1 U7344 ( .A1(n1989), .A2(n1988), .ZN(n1986) );
  OAI21_X1 U7345 ( .B1(n32704), .B2(n32327), .A(n32326), .ZN(n1989) );
  NAND2_X1 U7346 ( .A1(n1990), .A2(n21653), .ZN(n18853) );
  OAI21_X1 U7347 ( .B1(n1990), .B2(n16889), .A(n21653), .ZN(n16894) );
  OAI21_X1 U7348 ( .B1(n21819), .B2(n21823), .A(n23452), .ZN(n1992) );
  NAND2_X1 U7349 ( .A1(n24238), .A2(n24237), .ZN(n23452) );
  NAND3_X1 U7351 ( .A1(n47795), .A2(n47763), .A3(n47777), .ZN(n1994) );
  AND2_X1 U7352 ( .A1(n21908), .A2(n21907), .ZN(n1997) );
  INV_X1 U7353 ( .A(n23503), .ZN(n1998) );
  OAI21_X2 U7354 ( .B1(n14620), .B2(n14664), .A(n14619), .ZN(n2200) );
  OR2_X1 U7355 ( .A1(n49691), .A2(n2000), .ZN(n49255) );
  NAND2_X1 U7356 ( .A1(n49235), .A2(n49690), .ZN(n2000) );
  INV_X1 U7357 ( .A(n49235), .ZN(n49254) );
  AND2_X1 U7358 ( .A1(n49569), .A2(n49599), .ZN(n49564) );
  NAND2_X1 U7360 ( .A1(n2220), .A2(n19280), .ZN(n2003) );
  OAI21_X1 U7361 ( .B1(n19970), .B2(n1370), .A(n2003), .ZN(n19973) );
  NAND2_X1 U7362 ( .A1(n20337), .A2(n2003), .ZN(n20341) );
  NAND3_X1 U7363 ( .A1(n24455), .A2(n4177), .A3(n2004), .ZN(n24454) );
  NOR2_X1 U7364 ( .A1(n39906), .A2(n38448), .ZN(n38440) );
  NAND2_X1 U7366 ( .A1(n32665), .A2(n32660), .ZN(n2009) );
  NAND3_X1 U7367 ( .A1(n31454), .A2(n31538), .A3(n31546), .ZN(n32660) );
  NAND2_X1 U7368 ( .A1(n2010), .A2(n2009), .ZN(n32672) );
  NAND2_X1 U7369 ( .A1(n32661), .A2(n2011), .ZN(n2010) );
  INV_X1 U7370 ( .A(n32665), .ZN(n2011) );
  AND2_X1 U7371 ( .A1(n32694), .A2(n32332), .ZN(n2012) );
  NAND2_X1 U7372 ( .A1(n14117), .A2(n2013), .ZN(n14771) );
  NAND2_X1 U7373 ( .A1(n6588), .A2(n2015), .ZN(n45151) );
  INV_X1 U7374 ( .A(n47087), .ZN(n2015) );
  OAI21_X1 U7375 ( .B1(n41052), .B2(n41053), .A(n41051), .ZN(n41069) );
  NOR2_X1 U7377 ( .A1(n41049), .A2(n41054), .ZN(n41066) );
  NAND2_X1 U7378 ( .A1(n46521), .A2(n48416), .ZN(n46524) );
  NAND2_X1 U7379 ( .A1(n48177), .A2(n2017), .ZN(n48168) );
  AND2_X1 U7380 ( .A1(n11106), .A2(n2018), .ZN(n11117) );
  NAND2_X1 U7381 ( .A1(n5484), .A2(n10438), .ZN(n2018) );
  NOR2_X2 U7382 ( .A1(n11954), .A2(n8881), .ZN(n10438) );
  NAND2_X1 U7383 ( .A1(n757), .A2(n23254), .ZN(n21837) );
  NAND2_X2 U7384 ( .A1(n2019), .A2(n5626), .ZN(n23254) );
  NAND2_X1 U7385 ( .A1(n13495), .A2(n2021), .ZN(n2020) );
  NAND2_X1 U7387 ( .A1(n23066), .A2(n52155), .ZN(n2025) );
  NAND2_X1 U7390 ( .A1(n2025), .A2(n17420), .ZN(n23073) );
  NAND2_X1 U7391 ( .A1(n2026), .A2(n2029), .ZN(n29384) );
  NAND2_X1 U7392 ( .A1(n31043), .A2(n31816), .ZN(n2027) );
  AOI21_X1 U7394 ( .B1(n30576), .B2(n31816), .A(n31043), .ZN(n2030) );
  NAND2_X1 U7395 ( .A1(n1585), .A2(n51328), .ZN(n48828) );
  AND2_X1 U7396 ( .A1(n45739), .A2(n2031), .ZN(n45744) );
  NAND2_X1 U7397 ( .A1(n1585), .A2(n48808), .ZN(n48823) );
  NAND2_X1 U7398 ( .A1(n48834), .A2(n1585), .ZN(n45509) );
  NAND2_X1 U7399 ( .A1(n48830), .A2(n2032), .ZN(n45510) );
  AOI21_X1 U7400 ( .B1(n2034), .B2(n45739), .A(n48808), .ZN(n2032) );
  NAND2_X1 U7401 ( .A1(n45746), .A2(n1585), .ZN(n45709) );
  NAND2_X1 U7402 ( .A1(n48824), .A2(n2035), .ZN(n45516) );
  AND2_X1 U7403 ( .A1(n52434), .A2(n1585), .ZN(n2035) );
  OAI21_X1 U7404 ( .B1(n1585), .B2(n48799), .A(n48838), .ZN(n48800) );
  NOR2_X1 U7405 ( .A1(n32595), .A2(n28171), .ZN(n2036) );
  NAND2_X1 U7406 ( .A1(n32600), .A2(n2037), .ZN(n28171) );
  NAND2_X1 U7407 ( .A1(n32590), .A2(n2037), .ZN(n30513) );
  NAND2_X1 U7408 ( .A1(n32592), .A2(n32988), .ZN(n29617) );
  NAND2_X1 U7409 ( .A1(n2037), .A2(n32595), .ZN(n32989) );
  AOI21_X1 U7410 ( .B1(n712), .B2(n32990), .A(n2037), .ZN(n30519) );
  NAND3_X1 U7411 ( .A1(n52046), .A2(n32600), .A3(n32588), .ZN(n30508) );
  AND2_X1 U7412 ( .A1(n29622), .A2(n2037), .ZN(n32588) );
  NAND2_X1 U7413 ( .A1(n32975), .A2(n2036), .ZN(n30504) );
  NAND3_X1 U7415 ( .A1(n2039), .A2(n44655), .A3(n2038), .ZN(n47966) );
  NAND2_X1 U7416 ( .A1(n2040), .A2(n47909), .ZN(n2038) );
  NAND2_X1 U7417 ( .A1(n47911), .A2(n47907), .ZN(n2040) );
  NAND3_X1 U7418 ( .A1(n2042), .A2(n21758), .A3(n23338), .ZN(n21147) );
  NAND4_X1 U7419 ( .A1(n21144), .A2(n629), .A3(n21145), .A4(n21756), .ZN(n2042) );
  NAND3_X1 U7420 ( .A1(n2043), .A2(n37964), .A3(n37965), .ZN(n37967) );
  AND3_X1 U7421 ( .A1(n2043), .A2(n36539), .A3(n37964), .ZN(n37959) );
  NAND2_X1 U7422 ( .A1(n34092), .A2(n2043), .ZN(n8013) );
  AOI21_X1 U7423 ( .B1(n34663), .B2(n51077), .A(n2043), .ZN(n34664) );
  NAND3_X1 U7424 ( .A1(n34995), .A2(n2043), .A3(n34996), .ZN(n34999) );
  NAND2_X1 U7425 ( .A1(n773), .A2(n17311), .ZN(n3995) );
  NAND3_X1 U7426 ( .A1(n2044), .A2(n19518), .A3(n19504), .ZN(n21229) );
  NAND2_X1 U7427 ( .A1(n773), .A2(n2045), .ZN(n16655) );
  NAND2_X1 U7428 ( .A1(n19510), .A2(n19112), .ZN(n17311) );
  NAND2_X1 U7429 ( .A1(n11972), .A2(n789), .ZN(n11991) );
  NAND3_X1 U7430 ( .A1(n10341), .A2(n10342), .A3(n2046), .ZN(n10353) );
  NAND2_X1 U7431 ( .A1(n10455), .A2(n10451), .ZN(n2046) );
  OR2_X1 U7434 ( .A1(n34187), .A2(n34189), .ZN(n36627) );
  XNOR2_X1 U7436 ( .A(n44925), .B(n2051), .ZN(n42383) );
  XNOR2_X1 U7437 ( .A(n43914), .B(n2051), .ZN(n43534) );
  XNOR2_X1 U7438 ( .A(n2051), .B(n44546), .ZN(n42287) );
  XNOR2_X1 U7439 ( .A(n44536), .B(n2051), .ZN(n44545) );
  XNOR2_X1 U7440 ( .A(n2051), .B(n45298), .ZN(n45300) );
  NAND2_X1 U7441 ( .A1(n2056), .A2(n2052), .ZN(n26176) );
  OAI211_X1 U7442 ( .C1(n22117), .C2(n23209), .A(n2055), .B(n51355), .ZN(n2054) );
  NAND3_X1 U7443 ( .A1(n22116), .A2(n2102), .A3(n22115), .ZN(n2055) );
  NAND2_X1 U7444 ( .A1(n2057), .A2(n23231), .ZN(n2056) );
  NAND2_X1 U7445 ( .A1(n23235), .A2(n22122), .ZN(n2057) );
  NOR2_X1 U7446 ( .A1(n18332), .A2(n18331), .ZN(n2058) );
  OAI21_X1 U7447 ( .B1(n14330), .B2(n13008), .A(n13006), .ZN(n2060) );
  NAND2_X1 U7448 ( .A1(n40137), .A2(n40136), .ZN(n2063) );
  INV_X1 U7449 ( .A(n37924), .ZN(n2066) );
  INV_X1 U7450 ( .A(n37924), .ZN(n37209) );
  NAND2_X1 U7452 ( .A1(n38658), .A2(n2067), .ZN(n38661) );
  NAND2_X1 U7453 ( .A1(n39176), .A2(n700), .ZN(n2067) );
  XNOR2_X1 U7454 ( .A(n27235), .B(n26292), .ZN(n25570) );
  AND3_X1 U7455 ( .A1(n51728), .A2(n52172), .A3(n48382), .ZN(n2071) );
  OAI21_X1 U7456 ( .B1(n48376), .B2(n48306), .A(n2070), .ZN(n48307) );
  NAND3_X1 U7457 ( .A1(n51087), .A2(n48380), .A3(n2071), .ZN(n2070) );
  OR2_X2 U7458 ( .A1(n13449), .A2(n12790), .ZN(n13439) );
  NAND3_X2 U7459 ( .A1(n2073), .A2(n2074), .A3(n9797), .ZN(n14224) );
  NAND2_X1 U7460 ( .A1(n13232), .A2(n9856), .ZN(n2074) );
  NAND2_X1 U7461 ( .A1(n9796), .A2(n9795), .ZN(n13232) );
  NOR2_X1 U7462 ( .A1(n23160), .A2(n21945), .ZN(n2076) );
  INV_X1 U7463 ( .A(n22359), .ZN(n22919) );
  AND2_X1 U7464 ( .A1(n30734), .A2(n1121), .ZN(n2077) );
  NAND3_X1 U7468 ( .A1(n21966), .A2(n4619), .A3(n21965), .ZN(n26431) );
  OR2_X1 U7469 ( .A1(n21137), .A2(n21136), .ZN(n2082) );
  AND2_X1 U7470 ( .A1(n51695), .A2(n3553), .ZN(n2084) );
  OR2_X1 U7472 ( .A1(n36571), .A2(n36557), .ZN(n36488) );
  INV_X1 U7473 ( .A(n36557), .ZN(n2086) );
  NAND2_X1 U7476 ( .A1(n35939), .A2(n36196), .ZN(n2089) );
  XNOR2_X1 U7478 ( .A(n41757), .B(n41756), .ZN(n2092) );
  NAND2_X1 U7480 ( .A1(n6049), .A2(n803), .ZN(n2093) );
  AND2_X1 U7482 ( .A1(n3298), .A2(n3297), .ZN(n2097) );
  INV_X1 U7483 ( .A(n18671), .ZN(n2099) );
  INV_X1 U7484 ( .A(n16218), .ZN(n2101) );
  XNOR2_X1 U7485 ( .A(n42907), .B(n44904), .ZN(n2103) );
  INV_X1 U7487 ( .A(n12129), .ZN(n2105) );
  NAND2_X1 U7488 ( .A1(n4046), .A2(n6837), .ZN(n31683) );
  NOR2_X1 U7489 ( .A1(n26795), .A2(n30983), .ZN(n31691) );
  XNOR2_X1 U7490 ( .A(n14903), .B(n18147), .ZN(n16730) );
  XNOR2_X1 U7491 ( .A(n36680), .B(n7620), .ZN(n5262) );
  XNOR2_X1 U7492 ( .A(n16209), .B(n16210), .ZN(n19141) );
  XNOR2_X1 U7493 ( .A(n42907), .B(n44904), .ZN(n42453) );
  NAND4_X1 U7494 ( .A1(n22972), .A2(n22971), .A3(n22970), .A4(n22969), .ZN(
        n2106) );
  INV_X1 U7495 ( .A(n6944), .ZN(n2107) );
  AND2_X1 U7497 ( .A1(n21786), .A2(n20945), .ZN(n2108) );
  XNOR2_X1 U7498 ( .A(n22975), .B(n22974), .ZN(n2109) );
  AOI22_X1 U7500 ( .A1(n21636), .A2(n21637), .B1(n21635), .B2(n21634), .ZN(
        n21642) );
  OR2_X1 U7501 ( .A1(n44825), .A2(n42181), .ZN(n45532) );
  AND2_X1 U7502 ( .A1(n30283), .A2(n30296), .ZN(n2110) );
  AND2_X1 U7503 ( .A1(n28147), .A2(n28560), .ZN(n2111) );
  BUF_X1 U7505 ( .A(n18523), .Z(n2113) );
  XNOR2_X1 U7506 ( .A(n17234), .B(n18157), .ZN(n18523) );
  NAND4_X1 U7507 ( .A1(n9158), .A2(n8025), .A3(n9156), .A4(n9157), .ZN(n14643)
         );
  XNOR2_X1 U7508 ( .A(n24404), .B(n3031), .ZN(n26008) );
  INV_X1 U7510 ( .A(n11907), .ZN(n2116) );
  INV_X1 U7511 ( .A(n523), .ZN(n8021) );
  OR2_X1 U7512 ( .A1(n20210), .A2(n51006), .ZN(n2118) );
  NAND2_X1 U7513 ( .A1(n45538), .A2(n52070), .ZN(n2119) );
  AND2_X1 U7514 ( .A1(n38270), .A2(n2123), .ZN(n2120) );
  XNOR2_X1 U7517 ( .A(n18531), .B(n15956), .ZN(n2126) );
  NAND4_X1 U7520 ( .A1(n12898), .A2(n12897), .A3(n12896), .A4(n12895), .ZN(
        n18531) );
  XNOR2_X1 U7521 ( .A(n36703), .B(n34844), .ZN(n34433) );
  XNOR2_X1 U7522 ( .A(n34449), .B(n34448), .ZN(n37618) );
  XNOR2_X1 U7523 ( .A(n6434), .B(n24556), .ZN(n25821) );
  XNOR2_X1 U7524 ( .A(n15956), .B(n18531), .ZN(n16620) );
  OAI211_X1 U7525 ( .C1(n30967), .C2(n31540), .A(n30966), .B(n30965), .ZN(
        n34844) );
  NAND4_X1 U7526 ( .A1(n31049), .A2(n31047), .A3(n31046), .A4(n31048), .ZN(
        n2131) );
  XNOR2_X1 U7528 ( .A(n34413), .B(n34881), .ZN(n2133) );
  NAND4_X1 U7529 ( .A1(n31049), .A2(n31047), .A3(n31046), .A4(n31048), .ZN(
        n34413) );
  XNOR2_X1 U7530 ( .A(n34413), .B(n34881), .ZN(n5423) );
  INV_X1 U7531 ( .A(n305), .ZN(n2134) );
  INV_X1 U7532 ( .A(n305), .ZN(n2135) );
  INV_X1 U7533 ( .A(n305), .ZN(n2136) );
  AND3_X1 U7538 ( .A1(n17206), .A2(n3410), .A3(n3409), .ZN(n3408) );
  NAND3_X2 U7539 ( .A1(n46779), .A2(n6568), .A3(n46785), .ZN(n47573) );
  OR2_X1 U7541 ( .A1(n22314), .A2(n2676), .ZN(n2138) );
  NAND2_X1 U7543 ( .A1(n6825), .A2(n37739), .ZN(n2139) );
  OR2_X1 U7546 ( .A1(n16217), .A2(n20052), .ZN(n20078) );
  OAI21_X1 U7547 ( .B1(n17418), .B2(n23075), .A(n20555), .ZN(n24208) );
  AND2_X1 U7549 ( .A1(n35732), .A2(n37647), .ZN(n2141) );
  XNOR2_X1 U7554 ( .A(n28389), .B(n28388), .ZN(n30459) );
  XNOR2_X1 U7555 ( .A(n20541), .B(n20540), .ZN(n27729) );
  NAND4_X1 U7556 ( .A1(n13455), .A2(n13453), .A3(n13452), .A4(n13454), .ZN(
        n18522) );
  AOI21_X1 U7557 ( .B1(n30622), .B2(n30619), .A(n30623), .ZN(n31753) );
  XNOR2_X1 U7560 ( .A(n45420), .B(n45419), .ZN(n46510) );
  NAND4_X1 U7562 ( .A1(n30028), .A2(n30026), .A3(n30027), .A4(n30025), .ZN(
        n37112) );
  XNOR2_X1 U7565 ( .A(n1376), .B(n27512), .ZN(n30432) );
  NOR2_X1 U7568 ( .A1(n2838), .A2(n2839), .ZN(n14687) );
  NAND3_X1 U7569 ( .A1(n4094), .A2(n36043), .A3(n36041), .ZN(n2153) );
  XNOR2_X1 U7570 ( .A(n36855), .B(n35841), .ZN(n5454) );
  NAND4_X1 U7571 ( .A1(n26923), .A2(n26924), .A3(n26922), .A4(n26921), .ZN(
        n31110) );
  XNOR2_X1 U7572 ( .A(n8964), .B(Key[30]), .ZN(n11932) );
  NAND2_X2 U7574 ( .A1(n13816), .A2(n2482), .ZN(n17787) );
  XNOR2_X1 U7575 ( .A(n17691), .B(n18135), .ZN(n18592) );
  XNOR2_X1 U7576 ( .A(n44572), .B(n44571), .ZN(n46880) );
  NAND4_X1 U7579 ( .A1(n14495), .A2(n14496), .A3(n14494), .A4(n14493), .ZN(
        n18780) );
  XNOR2_X1 U7582 ( .A(n28103), .B(n28427), .ZN(n27393) );
  XNOR2_X1 U7583 ( .A(n16209), .B(n8398), .ZN(n20026) );
  XNOR2_X1 U7584 ( .A(n35325), .B(n36805), .ZN(n33981) );
  XNOR2_X1 U7585 ( .A(n8081), .B(n25429), .ZN(n28101) );
  XNOR2_X1 U7586 ( .A(n27195), .B(n22813), .ZN(n23112) );
  NAND4_X1 U7591 ( .A1(n9825), .A2(n9824), .A3(n9822), .A4(n9823), .ZN(n13945)
         );
  BUF_X1 U7592 ( .A(n22915), .Z(n2174) );
  OAI211_X1 U7593 ( .C1(n20492), .C2(n21465), .A(n17749), .B(n17748), .ZN(
        n22915) );
  XNOR2_X1 U7594 ( .A(n6345), .B(n42380), .ZN(n44925) );
  XNOR2_X1 U7595 ( .A(Key[6]), .B(n8912), .ZN(n12496) );
  INV_X1 U7597 ( .A(n41706), .ZN(n2179) );
  XNOR2_X1 U7598 ( .A(n5221), .B(n7166), .ZN(n19214) );
  XNOR2_X1 U7599 ( .A(n17326), .B(n17224), .ZN(n19119) );
  OAI211_X1 U7600 ( .C1(n36662), .C2(n36663), .A(n36661), .B(n36660), .ZN(
        n45400) );
  XNOR2_X1 U7602 ( .A(n35299), .B(n2691), .ZN(n38258) );
  BUF_X2 U7603 ( .A(n15060), .Z(n2189) );
  NAND4_X1 U7604 ( .A1(n12734), .A2(n12735), .A3(n12736), .A4(n12733), .ZN(
        n15060) );
  XNOR2_X1 U7606 ( .A(n9360), .B(Key[97]), .ZN(n12084) );
  XNOR2_X1 U7608 ( .A(n6209), .B(n2338), .ZN(n28145) );
  BUF_X1 U7609 ( .A(n45127), .Z(n2196) );
  NAND3_X1 U7610 ( .A1(n39051), .A2(n4918), .A3(n5960), .ZN(n45127) );
  XNOR2_X1 U7611 ( .A(n8696), .B(Key[131]), .ZN(n8818) );
  XNOR2_X1 U7612 ( .A(n46078), .B(n46077), .ZN(n50383) );
  XNOR2_X1 U7613 ( .A(n7429), .B(n7428), .ZN(n30180) );
  NAND4_X1 U7614 ( .A1(n30589), .A2(n30587), .A3(n30588), .A4(n30586), .ZN(
        n33709) );
  XNOR2_X1 U7615 ( .A(n22517), .B(n22516), .ZN(n30718) );
  XNOR2_X1 U7617 ( .A(n44561), .B(n43547), .ZN(n45101) );
  NAND4_X1 U7618 ( .A1(n32734), .A2(n32735), .A3(n32736), .A4(n32733), .ZN(
        n33336) );
  XNOR2_X1 U7619 ( .A(n26176), .B(n27272), .ZN(n25771) );
  INV_X1 U7620 ( .A(n33383), .ZN(n37269) );
  XNOR2_X1 U7621 ( .A(n45283), .B(n45282), .ZN(n46463) );
  XNOR2_X1 U7625 ( .A(n26508), .B(n24302), .ZN(n28312) );
  NAND4_X1 U7627 ( .A1(n18855), .A2(n18852), .A3(n18854), .A4(n18853), .ZN(
        n23755) );
  OR2_X1 U7628 ( .A1(n37759), .A2(n35923), .ZN(n37747) );
  XNOR2_X1 U7629 ( .A(Key[189]), .B(Ciphertext[56]), .ZN(n11907) );
  XNOR2_X1 U7631 ( .A(n5020), .B(n27183), .ZN(n29443) );
  XNOR2_X1 U7634 ( .A(n18539), .B(n17212), .ZN(n17913) );
  BUF_X2 U7635 ( .A(n18819), .Z(n2217) );
  XNOR2_X1 U7637 ( .A(n16923), .B(n17258), .ZN(n18819) );
  XNOR2_X1 U7640 ( .A(n7686), .B(n19212), .ZN(n21484) );
  BUF_X1 U7641 ( .A(n40272), .Z(n2223) );
  NAND4_X1 U7642 ( .A1(n37972), .A2(n37970), .A3(n37971), .A4(n37973), .ZN(
        n40272) );
  XNOR2_X1 U7643 ( .A(n15677), .B(n7079), .ZN(n18804) );
  XNOR2_X1 U7644 ( .A(Ciphertext[26]), .B(Key[171]), .ZN(n12651) );
  XNOR2_X1 U7646 ( .A(n4921), .B(n17346), .ZN(n21212) );
  INV_X1 U7647 ( .A(n10539), .ZN(n9960) );
  AND2_X1 U7648 ( .A1(n12834), .A2(n13632), .ZN(n3427) );
  NAND4_X1 U7649 ( .A1(n12872), .A2(n12871), .A3(n12870), .A4(n3512), .ZN(
        n12971) );
  XNOR2_X1 U7650 ( .A(n17963), .B(n17962), .ZN(n18825) );
  XNOR2_X1 U7651 ( .A(n18475), .B(n3013), .ZN(n17961) );
  XNOR2_X1 U7652 ( .A(n14585), .B(n6035), .ZN(n17113) );
  INV_X1 U7653 ( .A(n16158), .ZN(n6035) );
  INV_X1 U7654 ( .A(n17496), .ZN(n20025) );
  XNOR2_X1 U7655 ( .A(n16176), .B(n8220), .ZN(n16438) );
  INV_X1 U7656 ( .A(n18832), .ZN(n8220) );
  XNOR2_X1 U7658 ( .A(n636), .B(n18740), .ZN(n18741) );
  XNOR2_X1 U7659 ( .A(n17968), .B(n17967), .ZN(n17979) );
  XNOR2_X1 U7660 ( .A(n16093), .B(n15747), .ZN(n8129) );
  XNOR2_X1 U7661 ( .A(n16419), .B(n16418), .ZN(n3766) );
  INV_X1 U7662 ( .A(n51710), .ZN(n21559) );
  AND3_X1 U7664 ( .A1(n7100), .A2(n7098), .A3(n7099), .ZN(n7095) );
  AOI21_X1 U7667 ( .B1(n20097), .B2(n20086), .A(n778), .ZN(n18323) );
  AND2_X1 U7669 ( .A1(n3589), .A2(n21185), .ZN(n21171) );
  INV_X1 U7670 ( .A(n20101), .ZN(n17603) );
  INV_X1 U7671 ( .A(n21664), .ZN(n20659) );
  INV_X1 U7672 ( .A(n16489), .ZN(n5853) );
  OR2_X1 U7673 ( .A1(n23320), .A2(n23318), .ZN(n23321) );
  AND2_X1 U7674 ( .A1(n21782), .A2(n21783), .ZN(n4225) );
  XNOR2_X1 U7675 ( .A(n25740), .B(n27450), .ZN(n23841) );
  AND2_X1 U7676 ( .A1(n21330), .A2(n21331), .ZN(n3333) );
  OR2_X1 U7677 ( .A1(n29239), .A2(n29240), .ZN(n29244) );
  XNOR2_X1 U7678 ( .A(n2164), .B(n23841), .ZN(n24722) );
  XNOR2_X1 U7679 ( .A(n27480), .B(n27479), .ZN(n28068) );
  INV_X1 U7680 ( .A(n26355), .ZN(n7833) );
  OR2_X1 U7682 ( .A1(n30339), .A2(n30351), .ZN(n30342) );
  XNOR2_X1 U7683 ( .A(n34471), .B(n34726), .ZN(n35350) );
  XNOR2_X1 U7684 ( .A(n5598), .B(n35632), .ZN(n34856) );
  INV_X1 U7685 ( .A(n460), .ZN(n8321) );
  AND2_X1 U7686 ( .A1(n33044), .A2(n33045), .ZN(n3293) );
  OAI21_X1 U7688 ( .B1(n11908), .B2(n8667), .A(n8666), .ZN(n11896) );
  AND2_X1 U7690 ( .A1(n10138), .A2(n10919), .ZN(n10931) );
  NAND2_X1 U7691 ( .A1(n6049), .A2(n9465), .ZN(n10178) );
  NAND2_X1 U7692 ( .A1(n9178), .A2(n9186), .ZN(n10449) );
  INV_X1 U7693 ( .A(n12242), .ZN(n6661) );
  AND2_X1 U7694 ( .A1(n13086), .A2(n13102), .ZN(n3081) );
  INV_X1 U7695 ( .A(n12292), .ZN(n10232) );
  AND2_X1 U7696 ( .A1(n10224), .A2(n10726), .ZN(n10229) );
  INV_X1 U7697 ( .A(n9826), .ZN(n10541) );
  INV_X1 U7698 ( .A(n12383), .ZN(n7891) );
  INV_X1 U7699 ( .A(n9369), .ZN(n7895) );
  INV_X1 U7700 ( .A(n10683), .ZN(n11351) );
  INV_X1 U7701 ( .A(n10451), .ZN(n12652) );
  NOR2_X1 U7702 ( .A1(n10859), .A2(n12555), .ZN(n11575) );
  INV_X1 U7703 ( .A(n9104), .ZN(n7482) );
  AND2_X1 U7704 ( .A1(n13089), .A2(n8187), .ZN(n11157) );
  INV_X1 U7705 ( .A(n10921), .ZN(n10932) );
  INV_X1 U7707 ( .A(n10100), .ZN(n10520) );
  OR2_X1 U7708 ( .A1(n14234), .A2(n14228), .ZN(n13220) );
  AND2_X1 U7709 ( .A1(n13872), .A2(n3700), .ZN(n13892) );
  AND2_X1 U7710 ( .A1(n8981), .A2(n8979), .ZN(n4810) );
  XNOR2_X1 U7711 ( .A(n16897), .B(n42339), .ZN(n16248) );
  AND2_X1 U7712 ( .A1(n13785), .A2(n13777), .ZN(n3773) );
  NOR2_X1 U7713 ( .A1(n7498), .A2(n13772), .ZN(n7497) );
  OR2_X1 U7714 ( .A1(n13787), .A2(n13786), .ZN(n7496) );
  INV_X1 U7715 ( .A(n17280), .ZN(n8221) );
  INV_X1 U7716 ( .A(n20393), .ZN(n18000) );
  XNOR2_X1 U7717 ( .A(n51482), .B(n8034), .ZN(n17351) );
  XNOR2_X1 U7718 ( .A(n15824), .B(n8029), .ZN(n8028) );
  INV_X1 U7720 ( .A(n21525), .ZN(n20612) );
  INV_X1 U7721 ( .A(n20658), .ZN(n20657) );
  INV_X1 U7722 ( .A(n19819), .ZN(n5231) );
  INV_X1 U7723 ( .A(n20188), .ZN(n3243) );
  NOR2_X1 U7724 ( .A1(n21520), .A2(n52213), .ZN(n21531) );
  XNOR2_X1 U7726 ( .A(n15889), .B(n15890), .ZN(n16577) );
  INV_X1 U7727 ( .A(n20512), .ZN(n20506) );
  AND2_X1 U7728 ( .A1(n17579), .A2(n17580), .ZN(n3642) );
  INV_X1 U7729 ( .A(n18332), .ZN(n18336) );
  INV_X1 U7730 ( .A(n21652), .ZN(n21661) );
  XNOR2_X1 U7732 ( .A(n18561), .B(n18562), .ZN(n20326) );
  INV_X1 U7734 ( .A(n17784), .ZN(n8190) );
  AND2_X1 U7736 ( .A1(n19966), .A2(n19965), .ZN(n20451) );
  INV_X1 U7737 ( .A(n19055), .ZN(n19540) );
  INV_X1 U7738 ( .A(n20114), .ZN(n2749) );
  OR2_X1 U7739 ( .A1(n417), .A2(n23207), .ZN(n22117) );
  INV_X1 U7740 ( .A(n23207), .ZN(n6313) );
  INV_X1 U7742 ( .A(n373), .ZN(n19851) );
  AND3_X1 U7743 ( .A1(n21626), .A2(n21627), .A3(n21625), .ZN(n21644) );
  INV_X1 U7744 ( .A(n23341), .ZN(n3062) );
  OAI21_X1 U7745 ( .B1(n3598), .B2(n3600), .A(n20827), .ZN(n20832) );
  NOR2_X1 U7746 ( .A1(n20823), .A2(n20822), .ZN(n3600) );
  INV_X1 U7748 ( .A(n21200), .ZN(n19809) );
  AND2_X1 U7749 ( .A1(n21528), .A2(n20608), .ZN(n18902) );
  OAI21_X1 U7750 ( .B1(n21286), .B2(n51013), .A(n19017), .ZN(n7187) );
  OR2_X1 U7751 ( .A1(n18893), .A2(n21520), .ZN(n21518) );
  INV_X1 U7752 ( .A(n20089), .ZN(n20085) );
  AND2_X1 U7753 ( .A1(n17579), .A2(n17564), .ZN(n8605) );
  AND2_X1 U7754 ( .A1(n17561), .A2(n17556), .ZN(n8324) );
  AND2_X1 U7756 ( .A1(n17582), .A2(n16847), .ZN(n4700) );
  INV_X1 U7757 ( .A(n23207), .ZN(n23219) );
  OAI21_X1 U7758 ( .B1(n21457), .B2(n21456), .A(n21455), .ZN(n21478) );
  AND2_X1 U7759 ( .A1(n358), .A2(n21379), .ZN(n4002) );
  OR2_X1 U7760 ( .A1(n20197), .A2(n18495), .ZN(n20632) );
  INV_X1 U7761 ( .A(n22117), .ZN(n22120) );
  NOR2_X1 U7762 ( .A1(n6313), .A2(n413), .ZN(n8732) );
  NAND2_X1 U7763 ( .A1(n17608), .A2(n20105), .ZN(n6358) );
  NAND3_X1 U7764 ( .A1(n17598), .A2(n17597), .A3(n16788), .ZN(n6361) );
  INV_X1 U7765 ( .A(n17510), .ZN(n22256) );
  AOI21_X1 U7766 ( .B1(n17507), .B2(n17508), .A(n4058), .ZN(n5194) );
  INV_X1 U7767 ( .A(n21767), .ZN(n20942) );
  AOI21_X1 U7768 ( .B1(n5371), .B2(n22741), .A(n5094), .ZN(n6377) );
  AOI21_X1 U7769 ( .B1(n16800), .B2(n6949), .A(n6948), .ZN(n6953) );
  OAI21_X2 U7770 ( .B1(n18337), .B2(n17553), .A(n17552), .ZN(n22155) );
  NAND2_X2 U7771 ( .A1(n4866), .A2(n15097), .ZN(n21782) );
  INV_X1 U7772 ( .A(n5143), .ZN(n23904) );
  AND3_X1 U7773 ( .A1(n21103), .A2(n21102), .A3(n21101), .ZN(n8737) );
  OR2_X1 U7774 ( .A1(n22185), .A2(n7104), .ZN(n4807) );
  AND2_X1 U7776 ( .A1(n23469), .A2(n23468), .ZN(n6001) );
  NOR2_X1 U7777 ( .A1(n24281), .A2(n24282), .ZN(n24301) );
  INV_X1 U7778 ( .A(n23841), .ZN(n25088) );
  XNOR2_X1 U7779 ( .A(n2950), .B(n25074), .ZN(n25410) );
  INV_X1 U7780 ( .A(n25228), .ZN(n6141) );
  AND3_X1 U7781 ( .A1(n27624), .A2(n27625), .A3(n27724), .ZN(n8358) );
  AND2_X1 U7782 ( .A1(n29880), .A2(n29881), .ZN(n29887) );
  XNOR2_X1 U7783 ( .A(n28101), .B(n24968), .ZN(n25144) );
  INV_X1 U7784 ( .A(n28545), .ZN(n26500) );
  OAI211_X1 U7785 ( .C1(n28012), .C2(n28927), .A(n7146), .B(n28937), .ZN(n7145) );
  XNOR2_X1 U7786 ( .A(n25142), .B(n26397), .ZN(n27396) );
  NOR2_X1 U7787 ( .A1(n383), .A2(n459), .ZN(n29320) );
  INV_X1 U7788 ( .A(n30163), .ZN(n30159) );
  OR2_X1 U7789 ( .A1(n29172), .A2(n51473), .ZN(n30247) );
  OR2_X1 U7790 ( .A1(n30247), .A2(n29155), .ZN(n30253) );
  INV_X1 U7792 ( .A(n32830), .ZN(n7409) );
  INV_X1 U7794 ( .A(n29270), .ZN(n29186) );
  INV_X1 U7795 ( .A(n26455), .ZN(n29013) );
  OR2_X1 U7796 ( .A1(n26459), .A2(n3161), .ZN(n28014) );
  AND2_X1 U7797 ( .A1(n29007), .A2(n51115), .ZN(n3159) );
  AND2_X1 U7798 ( .A1(n29315), .A2(n29320), .ZN(n26325) );
  INV_X1 U7799 ( .A(n27808), .ZN(n27897) );
  NOR2_X1 U7800 ( .A1(n30688), .A2(n30387), .ZN(n30685) );
  OR2_X1 U7801 ( .A1(n31931), .A2(n29601), .ZN(n30048) );
  NOR2_X1 U7802 ( .A1(n31346), .A2(n30051), .ZN(n31333) );
  AND2_X1 U7805 ( .A1(n28339), .A2(n28338), .ZN(n3037) );
  INV_X1 U7806 ( .A(n31028), .ZN(n31026) );
  NOR2_X1 U7808 ( .A1(n3723), .A2(n3725), .ZN(n3720) );
  INV_X1 U7809 ( .A(n3724), .ZN(n3721) );
  INV_X1 U7810 ( .A(n32337), .ZN(n2841) );
  INV_X1 U7811 ( .A(n35810), .ZN(n33608) );
  XNOR2_X1 U7812 ( .A(n33620), .B(n8748), .ZN(n33649) );
  XNOR2_X1 U7813 ( .A(n6240), .B(n34620), .ZN(n35391) );
  XNOR2_X1 U7814 ( .A(n35282), .B(n35391), .ZN(n37329) );
  XNOR2_X1 U7815 ( .A(n34478), .B(n34477), .ZN(n34528) );
  INV_X1 U7817 ( .A(n34605), .ZN(n7544) );
  INV_X1 U7818 ( .A(n36788), .ZN(n7447) );
  AND3_X1 U7819 ( .A1(n38330), .A2(n38334), .A3(n37190), .ZN(n38346) );
  XNOR2_X1 U7820 ( .A(n35509), .B(n35510), .ZN(n34839) );
  INV_X1 U7821 ( .A(n33650), .ZN(n37399) );
  XNOR2_X1 U7822 ( .A(n5811), .B(n5810), .ZN(n5809) );
  INV_X1 U7823 ( .A(n33648), .ZN(n37543) );
  INV_X1 U7824 ( .A(n5570), .ZN(n3157) );
  OAI21_X1 U7825 ( .B1(n5571), .B2(n38321), .A(n38319), .ZN(n5570) );
  INV_X1 U7826 ( .A(n39224), .ZN(n39243) );
  INV_X1 U7827 ( .A(n37416), .ZN(n38472) );
  XNOR2_X1 U7829 ( .A(n5516), .B(n5515), .ZN(n36161) );
  XNOR2_X1 U7830 ( .A(n35806), .B(n37296), .ZN(n5515) );
  INV_X1 U7831 ( .A(n3044), .ZN(n37376) );
  NAND2_X1 U7832 ( .A1(n36306), .A2(n38547), .ZN(n36305) );
  INV_X1 U7834 ( .A(n35866), .ZN(n38292) );
  INV_X1 U7835 ( .A(n39767), .ZN(n7268) );
  AND2_X1 U7836 ( .A1(n2153), .A2(n584), .ZN(n39553) );
  NOR2_X1 U7837 ( .A1(n2153), .A2(n584), .ZN(n40196) );
  XNOR2_X1 U7838 ( .A(n34055), .B(n34054), .ZN(n37969) );
  AOI22_X1 U7839 ( .A1(n33271), .A2(n38087), .B1(n36638), .B2(n34197), .ZN(
        n33277) );
  OR2_X1 U7840 ( .A1(n40032), .A2(n51430), .ZN(n40023) );
  OAI21_X1 U7841 ( .B1(n40664), .B2(n7763), .A(n7762), .ZN(n7761) );
  AND2_X1 U7842 ( .A1(n41193), .A2(n41207), .ZN(n7762) );
  AND2_X1 U7843 ( .A1(n39067), .A2(n39066), .ZN(n4748) );
  XNOR2_X1 U7844 ( .A(n42067), .B(n43698), .ZN(n43218) );
  XNOR2_X1 U7845 ( .A(n45299), .B(n52038), .ZN(n44931) );
  AND2_X1 U7847 ( .A1(n3108), .A2(n46595), .ZN(n46703) );
  INV_X1 U7848 ( .A(n43250), .ZN(n8495) );
  INV_X1 U7849 ( .A(n46498), .ZN(n2688) );
  NOR2_X1 U7850 ( .A1(n7177), .A2(n50342), .ZN(n7176) );
  AND2_X1 U7851 ( .A1(n8987), .A2(n10742), .ZN(n8994) );
  XNOR2_X1 U7852 ( .A(Key[63]), .B(Ciphertext[38]), .ZN(n8880) );
  AND2_X1 U7853 ( .A1(n8881), .A2(n12725), .ZN(n11941) );
  OR2_X1 U7854 ( .A1(n11374), .A2(n12113), .ZN(n10699) );
  AND2_X1 U7856 ( .A1(n10234), .A2(n7081), .ZN(n7080) );
  INV_X1 U7857 ( .A(n9032), .ZN(n10246) );
  AND2_X1 U7858 ( .A1(n9744), .A2(n11016), .ZN(n10251) );
  AND2_X1 U7859 ( .A1(n15385), .A2(n15386), .ZN(n14820) );
  OR2_X1 U7861 ( .A1(n2796), .A2(n9874), .ZN(n9474) );
  OAI21_X1 U7862 ( .B1(n51761), .B2(n10178), .A(n10540), .ZN(n3848) );
  INV_X1 U7863 ( .A(n11031), .ZN(n10585) );
  AND2_X1 U7864 ( .A1(n12285), .A2(n12294), .ZN(n10716) );
  BUF_X1 U7865 ( .A(n9405), .Z(n12113) );
  INV_X1 U7866 ( .A(n11375), .ZN(n11377) );
  INV_X1 U7867 ( .A(n9184), .ZN(n7540) );
  INV_X1 U7868 ( .A(n11591), .ZN(n11599) );
  INV_X1 U7869 ( .A(n9279), .ZN(n11244) );
  OR2_X1 U7870 ( .A1(n11535), .A2(n11534), .ZN(n11536) );
  NOR2_X1 U7871 ( .A1(n10539), .A2(n9826), .ZN(n8286) );
  AND2_X1 U7872 ( .A1(n11646), .A2(n5315), .ZN(n5314) );
  OR2_X1 U7873 ( .A1(n11657), .A2(n10570), .ZN(n9321) );
  AND2_X1 U7874 ( .A1(n9317), .A2(n10572), .ZN(n9318) );
  AND2_X1 U7875 ( .A1(n12257), .A2(n12260), .ZN(n2968) );
  AND2_X1 U7876 ( .A1(n11016), .A2(n10252), .ZN(n10245) );
  INV_X1 U7877 ( .A(n10965), .ZN(n10970) );
  INV_X1 U7878 ( .A(n7942), .ZN(n11014) );
  INV_X1 U7879 ( .A(n12522), .ZN(n5268) );
  INV_X1 U7880 ( .A(n14159), .ZN(n4461) );
  AND2_X1 U7881 ( .A1(n11333), .A2(n11326), .ZN(n3617) );
  AND2_X1 U7882 ( .A1(n11331), .A2(n11332), .ZN(n3620) );
  NAND2_X1 U7883 ( .A1(n3619), .A2(n12152), .ZN(n3618) );
  AND2_X1 U7884 ( .A1(n11954), .A2(n8881), .ZN(n11958) );
  OR2_X1 U7885 ( .A1(n9322), .A2(n9323), .ZN(n8296) );
  OR2_X1 U7887 ( .A1(n12096), .A2(n12373), .ZN(n4283) );
  OR2_X1 U7890 ( .A1(n10990), .A2(n9785), .ZN(n4080) );
  NOR2_X1 U7891 ( .A1(n8024), .A2(n12498), .ZN(n10838) );
  AND4_X2 U7892 ( .A1(n9489), .A2(n9488), .A3(n9487), .A4(n9490), .ZN(n13102)
         );
  AND2_X1 U7893 ( .A1(n9964), .A2(n9965), .ZN(n6041) );
  NOR2_X1 U7894 ( .A1(n10296), .A2(n12301), .ZN(n9767) );
  AND2_X1 U7895 ( .A1(n10916), .A2(n4161), .ZN(n4160) );
  AND2_X1 U7896 ( .A1(n11403), .A2(n11410), .ZN(n12130) );
  OR2_X1 U7897 ( .A1(n13142), .A2(n12907), .ZN(n11178) );
  INV_X1 U7898 ( .A(n11178), .ZN(n12900) );
  AND2_X1 U7900 ( .A1(n2620), .A2(n13743), .ZN(n12394) );
  AND2_X1 U7901 ( .A1(n3645), .A2(n12907), .ZN(n14189) );
  AND3_X1 U7903 ( .A1(n9672), .A2(n9673), .A3(n9671), .ZN(n4410) );
  OR2_X1 U7904 ( .A1(n12101), .A2(n7895), .ZN(n7892) );
  AND2_X1 U7905 ( .A1(n2926), .A2(n7894), .ZN(n7893) );
  OR2_X1 U7906 ( .A1(n11458), .A2(n12544), .ZN(n6762) );
  NAND4_X1 U7907 ( .A1(n6250), .A2(n10857), .A3(n10856), .A4(n10855), .ZN(
        n10877) );
  OAI21_X1 U7908 ( .B1(n11575), .B2(n10861), .A(n12578), .ZN(n5620) );
  NAND4_X1 U7910 ( .A1(n9514), .A2(n9513), .A3(n11660), .A4(n9944), .ZN(n3584)
         );
  INV_X1 U7911 ( .A(n13441), .ZN(n14657) );
  OR2_X1 U7912 ( .A1(n9735), .A2(n10933), .ZN(n3980) );
  OR2_X1 U7913 ( .A1(n9835), .A2(n10527), .ZN(n10524) );
  AOI21_X1 U7914 ( .B1(n10525), .B2(n10520), .A(n10521), .ZN(n10523) );
  NOR2_X1 U7915 ( .A1(n15034), .A2(n13797), .ZN(n13475) );
  AND2_X1 U7916 ( .A1(n15034), .A2(n13801), .ZN(n15045) );
  INV_X1 U7917 ( .A(n17117), .ZN(n14848) );
  AND3_X1 U7918 ( .A1(n9528), .A2(n9526), .A3(n9527), .ZN(n4180) );
  XNOR2_X1 U7920 ( .A(n16904), .B(n17364), .ZN(n17814) );
  INV_X1 U7921 ( .A(n13888), .ZN(n14872) );
  BUF_X2 U7922 ( .A(n10877), .Z(n15167) );
  XNOR2_X1 U7923 ( .A(n18394), .B(n6933), .ZN(n18664) );
  INV_X1 U7924 ( .A(n17906), .ZN(n6933) );
  INV_X1 U7925 ( .A(n19388), .ZN(n3865) );
  INV_X1 U7926 ( .A(n18147), .ZN(n16960) );
  XNOR2_X1 U7927 ( .A(n16095), .B(n16094), .ZN(n20613) );
  XNOR2_X1 U7928 ( .A(n16382), .B(n16381), .ZN(n18380) );
  INV_X1 U7929 ( .A(n19170), .ZN(n20363) );
  INV_X1 U7930 ( .A(n6500), .ZN(n6499) );
  OAI21_X1 U7931 ( .B1(n19013), .B2(n21208), .A(n19819), .ZN(n6500) );
  INV_X1 U7933 ( .A(n16986), .ZN(n6490) );
  INV_X1 U7934 ( .A(n17113), .ZN(n15600) );
  AND2_X1 U7935 ( .A1(n7259), .A2(n51127), .ZN(n7949) );
  INV_X1 U7936 ( .A(n16788), .ZN(n7131) );
  AND2_X1 U7937 ( .A1(n16798), .A2(n2166), .ZN(n2648) );
  AND2_X1 U7938 ( .A1(n2645), .A2(n2644), .ZN(n2650) );
  OR2_X1 U7939 ( .A1(n19356), .A2(n21468), .ZN(n6177) );
  NOR2_X1 U7940 ( .A1(n767), .A2(n774), .ZN(n3366) );
  INV_X1 U7941 ( .A(n5388), .ZN(n19800) );
  INV_X1 U7942 ( .A(n19796), .ZN(n8575) );
  XNOR2_X1 U7943 ( .A(n16950), .B(n2254), .ZN(n2713) );
  AOI21_X1 U7944 ( .B1(n19407), .B2(n19408), .A(n3671), .ZN(n19409) );
  INV_X1 U7945 ( .A(n19417), .ZN(n3671) );
  AND2_X1 U7946 ( .A1(n4193), .A2(n4194), .ZN(n5560) );
  INV_X1 U7947 ( .A(n7653), .ZN(n7652) );
  AOI21_X1 U7948 ( .B1(n21254), .B2(n21255), .A(n5659), .ZN(n21259) );
  AND2_X1 U7949 ( .A1(n3885), .A2(n21253), .ZN(n5659) );
  INV_X1 U7950 ( .A(n17076), .ZN(n21245) );
  OR2_X1 U7951 ( .A1(n17997), .A2(n20474), .ZN(n8232) );
  AND2_X1 U7952 ( .A1(n20840), .A2(n5494), .ZN(n5493) );
  OR2_X1 U7953 ( .A1(n21427), .A2(n52139), .ZN(n5494) );
  OR2_X1 U7954 ( .A1(n24105), .A2(n24411), .ZN(n23521) );
  INV_X1 U7955 ( .A(n5294), .ZN(n5292) );
  XNOR2_X1 U7956 ( .A(n8356), .B(n16418), .ZN(n4974) );
  INV_X1 U7957 ( .A(n19330), .ZN(n20430) );
  AND2_X1 U7958 ( .A1(n18863), .A2(n18873), .ZN(n8302) );
  OR2_X1 U7959 ( .A1(n21391), .A2(n6395), .ZN(n21382) );
  AND2_X1 U7960 ( .A1(n19349), .A2(n19350), .ZN(n7677) );
  AOI22_X1 U7961 ( .A1(n19343), .A2(n17619), .B1(n20506), .B2(n19342), .ZN(
        n4988) );
  INV_X1 U7963 ( .A(n23068), .ZN(n23075) );
  OAI21_X1 U7964 ( .B1(n20055), .B2(n17027), .A(n3379), .ZN(n3191) );
  AND2_X1 U7965 ( .A1(n19135), .A2(n20075), .ZN(n3379) );
  INV_X1 U7966 ( .A(n16216), .ZN(n3195) );
  AND2_X1 U7967 ( .A1(n19500), .A2(n2391), .ZN(n6023) );
  AND3_X1 U7968 ( .A1(n17095), .A2(n20112), .A3(n17097), .ZN(n6845) );
  AOI22_X1 U7969 ( .A1(n20740), .A2(n21542), .B1(n20741), .B2(n20748), .ZN(
        n20756) );
  OAI21_X1 U7970 ( .B1(n19322), .B2(n5875), .A(n19321), .ZN(n7451) );
  OR2_X1 U7971 ( .A1(n8076), .A2(n23481), .ZN(n21974) );
  INV_X1 U7972 ( .A(n23479), .ZN(n8076) );
  INV_X1 U7973 ( .A(n23306), .ZN(n6914) );
  AND2_X1 U7974 ( .A1(n20491), .A2(n20490), .ZN(n4240) );
  INV_X1 U7975 ( .A(n23160), .ZN(n21957) );
  AND4_X2 U7976 ( .A1(n5655), .A2(n5654), .A3(n21220), .A4(n21221), .ZN(n23171) );
  OR2_X1 U7977 ( .A1(n2456), .A2(n5284), .ZN(n5654) );
  AND2_X1 U7979 ( .A1(n21895), .A2(n21913), .ZN(n7522) );
  INV_X1 U7981 ( .A(n22165), .ZN(n19576) );
  INV_X1 U7982 ( .A(n22170), .ZN(n5311) );
  INV_X1 U7984 ( .A(n21074), .ZN(n21073) );
  INV_X1 U7985 ( .A(n23335), .ZN(n21742) );
  INV_X1 U7986 ( .A(n20868), .ZN(n21733) );
  OAI21_X1 U7987 ( .B1(n20085), .B2(n18324), .A(n16788), .ZN(n6316) );
  OAI21_X1 U7988 ( .B1(n19980), .B2(n20255), .A(n19979), .ZN(n8363) );
  AND3_X1 U7989 ( .A1(n2812), .A2(n2814), .A3(n2811), .ZN(n7628) );
  AND2_X1 U7990 ( .A1(n24324), .A2(n50990), .ZN(n3306) );
  XNOR2_X1 U7992 ( .A(n23107), .B(n24905), .ZN(n24691) );
  AND3_X1 U7994 ( .A1(n18367), .A2(n18366), .A3(n18365), .ZN(n3448) );
  INV_X1 U7995 ( .A(n23921), .ZN(n22805) );
  INV_X1 U7996 ( .A(n23925), .ZN(n23134) );
  INV_X1 U7998 ( .A(n21948), .ZN(n23154) );
  AND3_X1 U7999 ( .A1(n16494), .A2(n5854), .A3(n5853), .ZN(n7987) );
  OR2_X1 U8000 ( .A1(n2555), .A2(n21778), .ZN(n21129) );
  NOR2_X1 U8001 ( .A1(n3331), .A2(n4131), .ZN(n3330) );
  INV_X1 U8002 ( .A(n29472), .ZN(n27762) );
  XNOR2_X1 U8003 ( .A(n27467), .B(n26600), .ZN(n27263) );
  OR2_X1 U8004 ( .A1(n29555), .A2(n29546), .ZN(n26763) );
  INV_X1 U8005 ( .A(n27661), .ZN(n27071) );
  XNOR2_X1 U8006 ( .A(n25816), .B(n23187), .ZN(n26287) );
  XNOR2_X1 U8007 ( .A(n25144), .B(n24970), .ZN(n25220) );
  INV_X1 U8008 ( .A(n29764), .ZN(n29065) );
  XNOR2_X1 U8009 ( .A(n22339), .B(n4211), .ZN(n26804) );
  INV_X1 U8010 ( .A(n24392), .ZN(n4211) );
  XNOR2_X1 U8011 ( .A(n23524), .B(n8733), .ZN(n30788) );
  XNOR2_X1 U8012 ( .A(n25005), .B(n23745), .ZN(n5518) );
  INV_X1 U8013 ( .A(n28711), .ZN(n29282) );
  INV_X1 U8014 ( .A(n29899), .ZN(n27570) );
  XNOR2_X1 U8015 ( .A(n8281), .B(n2296), .ZN(n8280) );
  XNOR2_X1 U8016 ( .A(n25218), .B(n24826), .ZN(n8282) );
  AND2_X1 U8018 ( .A1(n5791), .A2(n5792), .ZN(n5790) );
  INV_X1 U8020 ( .A(n28849), .ZN(n30343) );
  XNOR2_X1 U8021 ( .A(n27239), .B(n2312), .ZN(n28796) );
  INV_X1 U8022 ( .A(n52147), .ZN(n6488) );
  INV_X1 U8024 ( .A(n30232), .ZN(n30227) );
  INV_X1 U8025 ( .A(n29183), .ZN(n29188) );
  INV_X1 U8026 ( .A(n29554), .ZN(n27702) );
  AND2_X1 U8027 ( .A1(n24563), .A2(n29467), .ZN(n27755) );
  XNOR2_X1 U8028 ( .A(n25012), .B(n22570), .ZN(n7944) );
  INV_X1 U8029 ( .A(n28529), .ZN(n27104) );
  AND2_X1 U8030 ( .A1(n5355), .A2(n28874), .ZN(n28872) );
  INV_X1 U8031 ( .A(n29029), .ZN(n5355) );
  AND2_X1 U8032 ( .A1(n27105), .A2(n29029), .ZN(n29039) );
  INV_X1 U8033 ( .A(n28874), .ZN(n27105) );
  OR2_X1 U8034 ( .A1(n26619), .A2(n28874), .ZN(n28881) );
  INV_X1 U8035 ( .A(n26937), .ZN(n3765) );
  INV_X1 U8036 ( .A(n29029), .ZN(n28883) );
  INV_X1 U8038 ( .A(n26393), .ZN(n7075) );
  XNOR2_X1 U8039 ( .A(n3470), .B(n28056), .ZN(n20887) );
  NOR2_X1 U8040 ( .A1(n31699), .A2(n31700), .ZN(n32120) );
  OR2_X1 U8041 ( .A1(n24878), .A2(n51748), .ZN(n27113) );
  INV_X1 U8042 ( .A(n29543), .ZN(n29567) );
  OR2_X1 U8043 ( .A1(n33034), .A2(n719), .ZN(n6984) );
  AND2_X1 U8044 ( .A1(n32867), .A2(n32876), .ZN(n4422) );
  OAI21_X1 U8045 ( .B1(n30433), .B2(n29867), .A(n5329), .ZN(n28334) );
  NAND2_X1 U8046 ( .A1(n29859), .A2(n1981), .ZN(n28335) );
  INV_X1 U8047 ( .A(n626), .ZN(n5417) );
  INV_X1 U8048 ( .A(n25626), .ZN(n29263) );
  OR2_X1 U8049 ( .A1(n27681), .A2(n27690), .ZN(n27678) );
  INV_X1 U8050 ( .A(n30601), .ZN(n30911) );
  INV_X1 U8052 ( .A(n30766), .ZN(n5769) );
  OR2_X1 U8053 ( .A1(n28507), .A2(n28458), .ZN(n28511) );
  AND2_X1 U8055 ( .A1(n30734), .A2(n1121), .ZN(n30364) );
  AND2_X1 U8056 ( .A1(n29882), .A2(n52181), .ZN(n3421) );
  AND3_X1 U8057 ( .A1(n25198), .A2(n30159), .A3(n30183), .ZN(n30303) );
  INV_X1 U8058 ( .A(n24878), .ZN(n30282) );
  AND2_X1 U8059 ( .A1(n28014), .A2(n28013), .ZN(n8185) );
  OR2_X1 U8060 ( .A1(n32822), .A2(n32816), .ZN(n32425) );
  OR2_X1 U8061 ( .A1(n33002), .A2(n31383), .ZN(n33013) );
  INV_X1 U8062 ( .A(n31443), .ZN(n32663) );
  INV_X1 U8063 ( .A(n29141), .ZN(n30307) );
  INV_X1 U8064 ( .A(n31700), .ZN(n31708) );
  NAND4_X1 U8065 ( .A1(n31712), .A2(n4381), .A3(n4379), .A4(n4539), .ZN(n26348) );
  AND2_X1 U8066 ( .A1(n26345), .A2(n26344), .ZN(n4539) );
  AOI21_X1 U8067 ( .B1(n26343), .B2(n29522), .A(n4380), .ZN(n4379) );
  INV_X1 U8068 ( .A(n30433), .ZN(n6770) );
  OR2_X1 U8069 ( .A1(n30342), .A2(n28849), .ZN(n30358) );
  NOR2_X1 U8070 ( .A1(n7383), .A2(n31850), .ZN(n31742) );
  NOR2_X1 U8071 ( .A1(n30881), .A2(n31986), .ZN(n31188) );
  OAI21_X1 U8072 ( .B1(n25514), .B2(n25515), .A(n29186), .ZN(n25517) );
  OR2_X1 U8073 ( .A1(n31550), .A2(n32666), .ZN(n31551) );
  AOI22_X1 U8074 ( .A1(n5865), .A2(n31542), .B1(n5864), .B2(n31543), .ZN(n5863) );
  INV_X1 U8075 ( .A(n34881), .ZN(n5998) );
  AND3_X1 U8076 ( .A1(n25969), .A2(n27899), .A3(n25971), .ZN(n6878) );
  INV_X1 U8078 ( .A(n35334), .ZN(n7291) );
  INV_X1 U8079 ( .A(n34856), .ZN(n5239) );
  XNOR2_X1 U8080 ( .A(n35686), .B(n37331), .ZN(n35693) );
  XNOR2_X1 U8081 ( .A(n33096), .B(n8619), .ZN(n38035) );
  INV_X1 U8082 ( .A(n33095), .ZN(n8619) );
  XNOR2_X1 U8084 ( .A(n35477), .B(n33686), .ZN(n35136) );
  INV_X1 U8085 ( .A(n34207), .ZN(n36375) );
  XNOR2_X1 U8086 ( .A(n35612), .B(n32751), .ZN(n6706) );
  NAND2_X1 U8087 ( .A1(n38212), .A2(n36305), .ZN(n35169) );
  XNOR2_X1 U8088 ( .A(n37249), .B(n35617), .ZN(n35666) );
  INV_X1 U8089 ( .A(n699), .ZN(n7851) );
  XNOR2_X1 U8090 ( .A(n33344), .B(n36796), .ZN(n35807) );
  OR2_X1 U8091 ( .A1(n37521), .A2(n35951), .ZN(n37532) );
  XNOR2_X1 U8092 ( .A(n36993), .B(n34623), .ZN(n8351) );
  INV_X1 U8094 ( .A(n7048), .ZN(n36885) );
  INV_X1 U8095 ( .A(n37764), .ZN(n37507) );
  INV_X1 U8096 ( .A(n38057), .ZN(n31621) );
  INV_X1 U8097 ( .A(n35405), .ZN(n37190) );
  INV_X1 U8099 ( .A(n38152), .ZN(n37571) );
  INV_X1 U8100 ( .A(n38587), .ZN(n38592) );
  INV_X1 U8101 ( .A(n38340), .ZN(n38329) );
  OR2_X1 U8103 ( .A1(n37667), .A2(n35405), .ZN(n38335) );
  INV_X1 U8104 ( .A(n37901), .ZN(n37900) );
  INV_X1 U8105 ( .A(n39027), .ZN(n39036) );
  XNOR2_X1 U8106 ( .A(n4602), .B(n36872), .ZN(n38937) );
  XNOR2_X1 U8107 ( .A(n7048), .B(n36886), .ZN(n38940) );
  INV_X1 U8108 ( .A(n38014), .ZN(n38189) );
  AND2_X1 U8109 ( .A1(n36598), .A2(n36600), .ZN(n8366) );
  OR2_X1 U8110 ( .A1(n36051), .A2(n696), .ZN(n36593) );
  NAND2_X1 U8111 ( .A1(n38565), .A2(n36105), .ZN(n38562) );
  AND2_X1 U8113 ( .A1(n1692), .A2(n36581), .ZN(n4279) );
  INV_X1 U8114 ( .A(n37759), .ZN(n37756) );
  INV_X1 U8115 ( .A(n37749), .ZN(n36239) );
  INV_X1 U8116 ( .A(n37765), .ZN(n37499) );
  XNOR2_X1 U8117 ( .A(n34162), .B(n34161), .ZN(n36473) );
  AND2_X1 U8118 ( .A1(n38188), .A2(n38177), .ZN(n38004) );
  INV_X1 U8119 ( .A(n37981), .ZN(n5712) );
  INV_X1 U8120 ( .A(n34948), .ZN(n2660) );
  NOR2_X1 U8121 ( .A1(n34208), .A2(n36372), .ZN(n38036) );
  INV_X1 U8122 ( .A(n35951), .ZN(n38501) );
  AND2_X1 U8123 ( .A1(n38188), .A2(n38001), .ZN(n3332) );
  INV_X1 U8124 ( .A(n37976), .ZN(n36351) );
  INV_X1 U8125 ( .A(n35017), .ZN(n5235) );
  INV_X1 U8126 ( .A(n38053), .ZN(n36342) );
  AND2_X1 U8128 ( .A1(n38566), .A2(n38560), .ZN(n38205) );
  OR2_X1 U8129 ( .A1(n38067), .A2(n51522), .ZN(n2959) );
  INV_X1 U8130 ( .A(n5236), .ZN(n38058) );
  INV_X1 U8131 ( .A(n38054), .ZN(n38148) );
  AND3_X1 U8132 ( .A1(n36632), .A2(n50984), .A3(n36312), .ZN(n34197) );
  AND2_X1 U8133 ( .A1(n36629), .A2(n34193), .ZN(n36638) );
  INV_X1 U8134 ( .A(n34960), .ZN(n38087) );
  INV_X1 U8135 ( .A(n36044), .ZN(n36456) );
  INV_X1 U8136 ( .A(n38214), .ZN(n38553) );
  INV_X1 U8137 ( .A(n51738), .ZN(n5846) );
  NOR2_X1 U8138 ( .A1(n41902), .A2(n41332), .ZN(n40729) );
  INV_X1 U8139 ( .A(n34656), .ZN(n8089) );
  AND2_X1 U8140 ( .A1(n35879), .A2(n36052), .ZN(n36585) );
  XNOR2_X1 U8141 ( .A(n37309), .B(n37308), .ZN(n37313) );
  INV_X1 U8142 ( .A(n39263), .ZN(n39016) );
  OR2_X1 U8143 ( .A1(n33458), .A2(n3048), .ZN(n35946) );
  AND2_X1 U8145 ( .A1(n4297), .A2(n38052), .ZN(n7513) );
  OR2_X1 U8146 ( .A1(n38290), .A2(n37624), .ZN(n37630) );
  AND4_X1 U8147 ( .A1(n34525), .A2(n38272), .A3(n37624), .A4(n37620), .ZN(
        n4418) );
  INV_X1 U8148 ( .A(n38284), .ZN(n36436) );
  AND2_X1 U8149 ( .A1(n40295), .A2(n42441), .ZN(n40051) );
  OR2_X1 U8150 ( .A1(n34807), .A2(n37720), .ZN(n3041) );
  AND2_X1 U8151 ( .A1(n39481), .A2(n39486), .ZN(n36212) );
  INV_X1 U8152 ( .A(n37990), .ZN(n36080) );
  AND2_X1 U8153 ( .A1(n37956), .A2(n36540), .ZN(n8012) );
  OR2_X1 U8154 ( .A1(n39767), .A2(n41446), .ZN(n40647) );
  INV_X1 U8155 ( .A(n36593), .ZN(n36591) );
  INV_X1 U8157 ( .A(n39968), .ZN(n7120) );
  NOR3_X1 U8158 ( .A1(n38313), .A2(n7772), .A3(n39299), .ZN(n38730) );
  AND2_X1 U8159 ( .A1(n32683), .A2(n32682), .ZN(n6552) );
  AND2_X1 U8160 ( .A1(n7268), .A2(n7267), .ZN(n40649) );
  AND2_X1 U8161 ( .A1(n39768), .A2(n41446), .ZN(n7267) );
  AND2_X1 U8162 ( .A1(n37961), .A2(n3625), .ZN(n3624) );
  OAI21_X1 U8163 ( .B1(n38487), .B2(n38486), .A(n38485), .ZN(n7749) );
  AND2_X1 U8164 ( .A1(n7932), .A2(n7931), .ZN(n7930) );
  AND2_X1 U8165 ( .A1(n35175), .A2(n31355), .ZN(n2719) );
  OR2_X1 U8168 ( .A1(n41670), .A2(n3489), .ZN(n41244) );
  AOI21_X1 U8169 ( .B1(n34903), .B2(n34904), .A(n6090), .ZN(n6089) );
  OAI211_X1 U8170 ( .C1(n39402), .C2(n37890), .A(n37884), .B(n39393), .ZN(
        n6087) );
  OR2_X1 U8171 ( .A1(n3738), .A2(n37894), .ZN(n37888) );
  XNOR2_X1 U8172 ( .A(n34077), .B(n34421), .ZN(n6292) );
  OR2_X1 U8173 ( .A1(n39576), .A2(n41004), .ZN(n43325) );
  OR2_X1 U8174 ( .A1(n39146), .A2(n38866), .ZN(n39705) );
  AND2_X1 U8175 ( .A1(n40565), .A2(n40156), .ZN(n6199) );
  XNOR2_X1 U8176 ( .A(n44974), .B(n5286), .ZN(n5285) );
  INV_X1 U8177 ( .A(n44973), .ZN(n5286) );
  XNOR2_X1 U8178 ( .A(n41458), .B(n44394), .ZN(n41759) );
  INV_X1 U8179 ( .A(n48273), .ZN(n6674) );
  XNOR2_X1 U8180 ( .A(n38400), .B(n2278), .ZN(n44665) );
  XNOR2_X1 U8181 ( .A(n44360), .B(n44361), .ZN(n44678) );
  XNOR2_X1 U8182 ( .A(n5883), .B(n5882), .ZN(n45560) );
  INV_X1 U8183 ( .A(n44168), .ZN(n5882) );
  XNOR2_X1 U8184 ( .A(n44167), .B(n7152), .ZN(n5883) );
  XNOR2_X1 U8185 ( .A(n44392), .B(n44166), .ZN(n7152) );
  INV_X1 U8187 ( .A(n43996), .ZN(n7036) );
  XNOR2_X1 U8188 ( .A(n43104), .B(n45068), .ZN(n43887) );
  XNOR2_X1 U8189 ( .A(n42955), .B(n44546), .ZN(n45439) );
  XNOR2_X1 U8190 ( .A(n4958), .B(n4957), .ZN(n4956) );
  INV_X1 U8191 ( .A(n46059), .ZN(n4957) );
  XNOR2_X1 U8192 ( .A(n41187), .B(n44541), .ZN(n4958) );
  XNOR2_X1 U8193 ( .A(n44505), .B(n2284), .ZN(n47096) );
  INV_X1 U8194 ( .A(n46781), .ZN(n6569) );
  OR2_X1 U8195 ( .A1(n52050), .A2(n52161), .ZN(n3959) );
  OR2_X1 U8196 ( .A1(n5322), .A2(n5323), .ZN(n5321) );
  INV_X1 U8197 ( .A(n48214), .ZN(n5323) );
  OR2_X1 U8198 ( .A1(n45547), .A2(n52161), .ZN(n45554) );
  AND2_X1 U8199 ( .A1(n48117), .A2(n46542), .ZN(n45611) );
  INV_X1 U8200 ( .A(n45614), .ZN(n8569) );
  INV_X1 U8201 ( .A(n46444), .ZN(n48459) );
  OR2_X1 U8203 ( .A1(n49168), .A2(n45649), .ZN(n45656) );
  OR2_X1 U8204 ( .A1(n46272), .A2(n46273), .ZN(n2825) );
  AND3_X1 U8205 ( .A1(n46249), .A2(n49170), .A3(n49177), .ZN(n45216) );
  INV_X1 U8206 ( .A(n49112), .ZN(n5662) );
  XNOR2_X1 U8207 ( .A(n45299), .B(n43526), .ZN(n7720) );
  OR2_X1 U8208 ( .A1(n47321), .A2(n50375), .ZN(n8534) );
  OR2_X1 U8209 ( .A1(n50385), .A2(n8532), .ZN(n8531) );
  INV_X1 U8210 ( .A(n6172), .ZN(n50010) );
  XNOR2_X1 U8211 ( .A(n3653), .B(n43506), .ZN(n3652) );
  AND2_X1 U8212 ( .A1(n45165), .A2(n44471), .ZN(n45157) );
  OR2_X1 U8213 ( .A1(n46840), .A2(n47126), .ZN(n4527) );
  AND2_X1 U8214 ( .A1(n3894), .A2(n3893), .ZN(n3889) );
  NAND3_X1 U8215 ( .A1(n3573), .A2(n28), .A3(n49642), .ZN(n49810) );
  NAND4_X1 U8217 ( .A1(n50303), .A2(n50296), .A3(n49942), .A4(n3572), .ZN(
        n3573) );
  AND2_X1 U8218 ( .A1(n46716), .A2(n46717), .ZN(n5410) );
  OR2_X1 U8219 ( .A1(n48112), .A2(n48100), .ZN(n48103) );
  AND2_X1 U8222 ( .A1(n48944), .A2(n48935), .ZN(n48954) );
  NOR2_X1 U8223 ( .A1(n49809), .A2(n49752), .ZN(n49705) );
  AND2_X1 U8224 ( .A1(n49648), .A2(n4250), .ZN(n50029) );
  AND2_X1 U8225 ( .A1(n49649), .A2(n49650), .ZN(n4250) );
  AND2_X1 U8226 ( .A1(n6172), .A2(n50325), .ZN(n49994) );
  AND2_X1 U8227 ( .A1(n52126), .A2(n50716), .ZN(n4039) );
  INV_X1 U8228 ( .A(n12057), .ZN(n7019) );
  INV_X1 U8230 ( .A(n12253), .ZN(n11339) );
  AOI21_X1 U8231 ( .B1(n3023), .B2(n3025), .A(n2954), .ZN(n11241) );
  INV_X1 U8234 ( .A(n12694), .ZN(n11125) );
  AND2_X1 U8235 ( .A1(n10741), .A2(n12260), .ZN(n7285) );
  INV_X1 U8236 ( .A(n10747), .ZN(n7286) );
  INV_X1 U8237 ( .A(n11648), .ZN(n5915) );
  NOR2_X1 U8238 ( .A1(n9585), .A2(n12169), .ZN(n12176) );
  INV_X1 U8239 ( .A(n12626), .ZN(n5220) );
  AND2_X1 U8240 ( .A1(n11186), .A2(n7341), .ZN(n12570) );
  AND2_X1 U8241 ( .A1(n12557), .A2(n2828), .ZN(n11572) );
  INV_X1 U8242 ( .A(n9234), .ZN(n10413) );
  XNOR2_X1 U8244 ( .A(Key[3]), .B(n9217), .ZN(n10360) );
  AND2_X1 U8245 ( .A1(n10921), .A2(n10920), .ZN(n3384) );
  INV_X1 U8246 ( .A(n12263), .ZN(n6267) );
  OAI21_X1 U8247 ( .B1(n12258), .B2(n11339), .A(n9646), .ZN(n10740) );
  NOR2_X1 U8248 ( .A1(n10739), .A2(n10738), .ZN(n10753) );
  AND2_X1 U8250 ( .A1(n11269), .A2(n10590), .ZN(n11672) );
  NOR2_X1 U8251 ( .A1(n11684), .A2(n11674), .ZN(n4186) );
  OR2_X1 U8252 ( .A1(n15358), .A2(n11853), .ZN(n13918) );
  OR2_X1 U8253 ( .A1(n13441), .A2(n13450), .ZN(n4210) );
  INV_X1 U8254 ( .A(n9927), .ZN(n11215) );
  INV_X1 U8255 ( .A(n11338), .ZN(n6067) );
  OR2_X1 U8256 ( .A1(n4797), .A2(n12292), .ZN(n7822) );
  NOR2_X1 U8257 ( .A1(n2347), .A2(n5358), .ZN(n5930) );
  AND2_X1 U8258 ( .A1(n5359), .A2(n12344), .ZN(n5358) );
  NOR2_X1 U8259 ( .A1(n12338), .A2(n10669), .ZN(n5359) );
  OR2_X1 U8260 ( .A1(n9378), .A2(n12054), .ZN(n10666) );
  OAI21_X1 U8261 ( .B1(n10665), .B2(n12051), .A(n10661), .ZN(n3807) );
  OR2_X1 U8262 ( .A1(n13316), .A2(n5176), .ZN(n13313) );
  INV_X1 U8263 ( .A(n15342), .ZN(n15332) );
  AND2_X1 U8264 ( .A1(n8840), .A2(n10926), .ZN(n5047) );
  AND2_X1 U8265 ( .A1(n10788), .A2(n10789), .ZN(n6385) );
  AND2_X1 U8266 ( .A1(n641), .A2(n12914), .ZN(n13087) );
  NOR2_X1 U8267 ( .A1(n15167), .A2(n51370), .ZN(n6320) );
  AND2_X1 U8268 ( .A1(n10161), .A2(n10000), .ZN(n3428) );
  OAI21_X1 U8269 ( .B1(n6294), .B2(n15306), .A(n15305), .ZN(n15311) );
  INV_X1 U8270 ( .A(n12453), .ZN(n7354) );
  NOR2_X1 U8271 ( .A1(n7354), .A2(n11082), .ZN(n12461) );
  INV_X1 U8272 ( .A(n8967), .ZN(n8965) );
  INV_X1 U8273 ( .A(n51760), .ZN(n12555) );
  AOI21_X1 U8274 ( .B1(n9130), .B2(n9131), .A(n8384), .ZN(n8383) );
  AND2_X1 U8275 ( .A1(n12557), .A2(n11525), .ZN(n8384) );
  INV_X1 U8276 ( .A(n12627), .ZN(n10462) );
  AND2_X1 U8277 ( .A1(n12245), .A2(n12244), .ZN(n4532) );
  AND2_X1 U8278 ( .A1(n12256), .A2(n12257), .ZN(n12271) );
  AND2_X1 U8279 ( .A1(n4351), .A2(n12330), .ZN(n12349) );
  OR2_X1 U8280 ( .A1(n11464), .A2(n11461), .ZN(n7968) );
  OAI21_X1 U8281 ( .B1(n454), .B2(n11635), .A(n11634), .ZN(n7964) );
  OAI21_X1 U8282 ( .B1(n11001), .B2(n9751), .A(n10246), .ZN(n7589) );
  AND2_X1 U8283 ( .A1(n9752), .A2(n10192), .ZN(n7588) );
  AND2_X1 U8284 ( .A1(n10286), .A2(n10673), .ZN(n10289) );
  AND2_X1 U8285 ( .A1(n8050), .A2(n12134), .ZN(n12146) );
  AND2_X1 U8286 ( .A1(n9605), .A2(n11410), .ZN(n12144) );
  NOR2_X1 U8287 ( .A1(n11374), .A2(n9632), .ZN(n10373) );
  INV_X1 U8288 ( .A(n15434), .ZN(n15448) );
  OR2_X1 U8289 ( .A1(n13367), .A2(n16039), .ZN(n13385) );
  INV_X1 U8290 ( .A(n14999), .ZN(n13709) );
  OAI211_X1 U8291 ( .C1(n9704), .C2(n12277), .A(n7080), .B(n10230), .ZN(n9399)
         );
  AND2_X1 U8292 ( .A1(n9376), .A2(n12053), .ZN(n4464) );
  OAI22_X1 U8294 ( .A1(n2701), .A2(n9748), .B1(n9032), .B2(n9031), .ZN(n2700)
         );
  INV_X1 U8295 ( .A(n11008), .ZN(n11000) );
  INV_X1 U8296 ( .A(n15378), .ZN(n14805) );
  INV_X1 U8297 ( .A(n3752), .ZN(n14821) );
  OR2_X1 U8298 ( .A1(n15279), .A2(n14962), .ZN(n14945) );
  OAI21_X1 U8301 ( .B1(n12315), .B2(n10302), .A(n12300), .ZN(n9765) );
  NOR2_X1 U8302 ( .A1(n10707), .A2(n4369), .ZN(n10713) );
  INV_X1 U8303 ( .A(n11315), .ZN(n7755) );
  AND2_X1 U8304 ( .A1(n2149), .A2(n14666), .ZN(n14673) );
  INV_X1 U8305 ( .A(n2151), .ZN(n14956) );
  OR2_X1 U8306 ( .A1(n14976), .A2(n14984), .ZN(n15100) );
  INV_X1 U8307 ( .A(n13917), .ZN(n13916) );
  AND2_X1 U8308 ( .A1(n4557), .A2(n14928), .ZN(n14931) );
  OR2_X1 U8309 ( .A1(n14930), .A2(n14929), .ZN(n4557) );
  INV_X1 U8310 ( .A(n15304), .ZN(n14924) );
  AND4_X1 U8311 ( .A1(n14920), .A2(n15766), .A3(n15067), .A4(n15307), .ZN(
        n4446) );
  OAI21_X1 U8312 ( .B1(n15767), .B2(n14922), .A(n14921), .ZN(n4445) );
  NOR2_X1 U8313 ( .A1(n8286), .A2(n5731), .ZN(n8288) );
  NOR2_X1 U8314 ( .A1(n14999), .A2(n5340), .ZN(n14992) );
  INV_X1 U8315 ( .A(n15131), .ZN(n5340) );
  INV_X1 U8316 ( .A(n9183), .ZN(n7538) );
  NOR2_X1 U8317 ( .A1(n15386), .A2(n15365), .ZN(n13917) );
  OR2_X1 U8319 ( .A1(n11157), .A2(n13103), .ZN(n12824) );
  NOR2_X1 U8320 ( .A1(n3317), .A2(n3316), .ZN(n3315) );
  OAI21_X1 U8322 ( .B1(n14036), .B2(n782), .A(n5733), .ZN(n5732) );
  NOR2_X1 U8323 ( .A1(n8568), .A2(n8567), .ZN(n8566) );
  AND2_X1 U8324 ( .A1(n9321), .A2(n9320), .ZN(n3078) );
  AND2_X1 U8325 ( .A1(n5002), .A2(n9314), .ZN(n3077) );
  AND2_X1 U8326 ( .A1(n5314), .A2(n9319), .ZN(n8329) );
  AND2_X1 U8327 ( .A1(n14149), .A2(n14164), .ZN(n13762) );
  OR2_X1 U8328 ( .A1(n6835), .A2(n14160), .ZN(n13764) );
  AND3_X1 U8329 ( .A1(n10080), .A2(n10075), .A3(n10076), .ZN(n4122) );
  OAI21_X1 U8330 ( .B1(n15335), .B2(n15435), .A(n15334), .ZN(n15339) );
  AND2_X1 U8331 ( .A1(n15327), .A2(n15445), .ZN(n3015) );
  OR2_X1 U8332 ( .A1(n3461), .A2(n14998), .ZN(n15000) );
  INV_X1 U8333 ( .A(n15003), .ZN(n5348) );
  AND2_X1 U8336 ( .A1(n10274), .A2(n12353), .ZN(n7594) );
  NOR2_X1 U8337 ( .A1(n15435), .A2(n15437), .ZN(n15443) );
  AND2_X1 U8339 ( .A1(n9330), .A2(n8296), .ZN(n7516) );
  OR2_X1 U8340 ( .A1(n14999), .A2(n15131), .ZN(n14260) );
  INV_X1 U8341 ( .A(n6494), .ZN(n6492) );
  OR2_X1 U8342 ( .A1(n6668), .A2(n13189), .ZN(n13192) );
  INV_X1 U8343 ( .A(n13377), .ZN(n13384) );
  INV_X1 U8344 ( .A(n14220), .ZN(n13219) );
  OR2_X1 U8345 ( .A1(n3672), .A2(n14368), .ZN(n14359) );
  OR2_X1 U8346 ( .A1(n13346), .A2(n14542), .ZN(n14365) );
  OAI21_X1 U8347 ( .B1(n8458), .B2(n10578), .A(n10584), .ZN(n8457) );
  OR2_X1 U8348 ( .A1(n12307), .A2(n12308), .ZN(n8561) );
  AND2_X1 U8349 ( .A1(n12306), .A2(n12305), .ZN(n8415) );
  NOR2_X1 U8350 ( .A1(n2392), .A2(n3932), .ZN(n12368) );
  NOR2_X1 U8351 ( .A1(n13091), .A2(n13088), .ZN(n3943) );
  INV_X1 U8352 ( .A(n10030), .ZN(n4450) );
  AND3_X1 U8354 ( .A1(n10405), .A2(n10404), .A3(n10403), .ZN(n4344) );
  AND3_X1 U8355 ( .A1(n10408), .A2(n10409), .A3(n10410), .ZN(n4441) );
  INV_X1 U8356 ( .A(n10535), .ZN(n7412) );
  INV_X1 U8357 ( .A(n2249), .ZN(n7253) );
  NOR2_X1 U8358 ( .A1(n11738), .A2(n9719), .ZN(n14477) );
  OR2_X1 U8359 ( .A1(n11750), .A2(n483), .ZN(n4232) );
  OR2_X1 U8360 ( .A1(n9730), .A2(n10142), .ZN(n5962) );
  OR2_X1 U8361 ( .A1(n9731), .A2(n10919), .ZN(n5963) );
  XNOR2_X1 U8362 ( .A(n14662), .B(n4511), .ZN(n15294) );
  INV_X1 U8363 ( .A(n17960), .ZN(n4511) );
  OR2_X1 U8364 ( .A1(n19078), .A2(n19077), .ZN(n19067) );
  XNOR2_X1 U8366 ( .A(n17234), .B(n15472), .ZN(n4534) );
  AND3_X1 U8367 ( .A1(n2957), .A2(n9532), .A3(n11168), .ZN(n4326) );
  AND2_X1 U8368 ( .A1(n9625), .A2(n9623), .ZN(n3405) );
  AND2_X1 U8369 ( .A1(n9624), .A2(n9629), .ZN(n3406) );
  AOI21_X1 U8370 ( .B1(n13132), .B2(n13137), .A(n3676), .ZN(n12910) );
  INV_X1 U8371 ( .A(n19534), .ZN(n19056) );
  XNOR2_X1 U8372 ( .A(n17178), .B(n15746), .ZN(n16093) );
  AND3_X1 U8373 ( .A1(n12978), .A2(n12979), .A3(n14438), .ZN(n2953) );
  INV_X1 U8374 ( .A(n16765), .ZN(n18714) );
  XNOR2_X1 U8376 ( .A(n19239), .B(n18436), .ZN(n5699) );
  XNOR2_X1 U8377 ( .A(n18553), .B(n15948), .ZN(n5700) );
  AND3_X1 U8378 ( .A1(n19378), .A2(n19376), .A3(n19377), .ZN(n5862) );
  INV_X1 U8379 ( .A(n19795), .ZN(n3683) );
  OR2_X1 U8381 ( .A1(n19636), .A2(n15630), .ZN(n7947) );
  OR2_X1 U8382 ( .A1(n20474), .A2(n20472), .ZN(n19381) );
  AND2_X1 U8383 ( .A1(n18330), .A2(n18062), .ZN(n17437) );
  INV_X1 U8384 ( .A(n19988), .ZN(n2861) );
  AND2_X1 U8386 ( .A1(n18043), .A2(n19410), .ZN(n3476) );
  AND2_X1 U8387 ( .A1(n20508), .A2(n489), .ZN(n18087) );
  INV_X1 U8388 ( .A(n18085), .ZN(n20504) );
  OR2_X1 U8389 ( .A1(n18030), .A2(n18029), .ZN(n21698) );
  AND2_X1 U8390 ( .A1(n19410), .A2(n18041), .ZN(n17559) );
  OAI21_X1 U8391 ( .B1(n19327), .B2(n50), .A(n2423), .ZN(n19178) );
  AND2_X1 U8392 ( .A1(n19331), .A2(n19330), .ZN(n3969) );
  NOR2_X1 U8393 ( .A1(n17045), .A2(n17447), .ZN(n3060) );
  INV_X1 U8394 ( .A(n18377), .ZN(n5881) );
  INV_X1 U8395 ( .A(n21441), .ZN(n21435) );
  INV_X1 U8396 ( .A(n21425), .ZN(n21442) );
  INV_X1 U8397 ( .A(n20838), .ZN(n20329) );
  OAI21_X1 U8398 ( .B1(n19071), .B2(n18344), .A(n20132), .ZN(n5458) );
  INV_X1 U8399 ( .A(n18053), .ZN(n20436) );
  AND2_X1 U8400 ( .A1(n20473), .A2(n20474), .ZN(n8592) );
  AND2_X1 U8401 ( .A1(n20375), .A2(n21388), .ZN(n20412) );
  OR2_X1 U8402 ( .A1(n20798), .A2(n581), .ZN(n3412) );
  OR2_X1 U8403 ( .A1(n6865), .A2(n20375), .ZN(n6864) );
  AND2_X1 U8404 ( .A1(n20641), .A2(n3189), .ZN(n20628) );
  INV_X1 U8405 ( .A(n20201), .ZN(n20623) );
  XNOR2_X1 U8406 ( .A(n4022), .B(n18395), .ZN(n18398) );
  NOR2_X1 U8407 ( .A1(n3885), .A2(n18962), .ZN(n17076) );
  INV_X1 U8408 ( .A(n3885), .ZN(n17083) );
  NOR2_X1 U8409 ( .A1(n24411), .A2(n24412), .ZN(n23518) );
  OR2_X1 U8410 ( .A1(n19955), .A2(n20838), .ZN(n3492) );
  INV_X1 U8411 ( .A(n20348), .ZN(n20351) );
  OR3_X2 U8412 ( .A1(n8139), .A2(n6934), .A3(n6935), .ZN(n23827) );
  AOI21_X1 U8413 ( .B1(n16111), .B2(n21512), .A(n20188), .ZN(n6935) );
  NOR2_X1 U8415 ( .A1(n19893), .A2(n19891), .ZN(n8354) );
  INV_X1 U8416 ( .A(n22989), .ZN(n3691) );
  INV_X1 U8417 ( .A(n23521), .ZN(n23732) );
  INV_X1 U8418 ( .A(n21251), .ZN(n3335) );
  INV_X1 U8419 ( .A(n21432), .ZN(n5146) );
  AND2_X1 U8420 ( .A1(n22937), .A2(n23044), .ZN(n8229) );
  OR2_X1 U8421 ( .A1(n23135), .A2(n3907), .ZN(n3906) );
  NAND4_X1 U8422 ( .A1(n2307), .A2(n19780), .A3(n19791), .A4(n19790), .ZN(
        n19901) );
  NOR2_X1 U8423 ( .A1(n22769), .A2(n19901), .ZN(n23102) );
  NAND2_X1 U8424 ( .A1(n25057), .A2(n23092), .ZN(n3042) );
  AND2_X1 U8425 ( .A1(n23417), .A2(n22046), .ZN(n7650) );
  AND2_X1 U8426 ( .A1(n6952), .A2(n18287), .ZN(n6949) );
  INV_X1 U8428 ( .A(n23304), .ZN(n8303) );
  NOR2_X1 U8429 ( .A1(n23303), .A2(n441), .ZN(n23318) );
  INV_X1 U8430 ( .A(n23317), .ZN(n8402) );
  AND2_X1 U8432 ( .A1(n8576), .A2(n8572), .ZN(n18225) );
  AND2_X1 U8434 ( .A1(n18004), .A2(n18005), .ZN(n2561) );
  OR2_X1 U8435 ( .A1(n21767), .A2(n758), .ZN(n21115) );
  AND3_X1 U8436 ( .A1(n21913), .A2(n21915), .A3(n7510), .ZN(n7511) );
  OAI211_X1 U8437 ( .C1(n6179), .C2(n19310), .A(n19306), .B(n6173), .ZN(n6178)
         );
  OR2_X1 U8438 ( .A1(n23136), .A2(n22521), .ZN(n21510) );
  INV_X1 U8439 ( .A(n19831), .ZN(n5244) );
  AND2_X1 U8440 ( .A1(n21174), .A2(n3088), .ZN(n3087) );
  AND2_X1 U8441 ( .A1(n3589), .A2(n19832), .ZN(n3088) );
  OAI21_X1 U8442 ( .B1(n19701), .B2(n19702), .A(n19704), .ZN(n3090) );
  OR2_X1 U8444 ( .A1(n23068), .A2(n17420), .ZN(n22268) );
  INV_X1 U8445 ( .A(n21974), .ZN(n23488) );
  NOR2_X1 U8446 ( .A1(n23143), .A2(n23924), .ZN(n23912) );
  AND2_X1 U8447 ( .A1(n22864), .A2(n22856), .ZN(n19612) );
  INV_X1 U8448 ( .A(n21975), .ZN(n7535) );
  AND2_X1 U8449 ( .A1(n20278), .A2(n20279), .ZN(n6745) );
  INV_X1 U8450 ( .A(n24237), .ZN(n21811) );
  NAND2_X1 U8452 ( .A1(n20325), .A2(n20326), .ZN(n20322) );
  OR2_X1 U8453 ( .A1(n23895), .A2(n3906), .ZN(n23925) );
  OR2_X1 U8454 ( .A1(n19513), .A2(n7049), .ZN(n16681) );
  AND2_X1 U8455 ( .A1(n51124), .A2(n22481), .ZN(n4719) );
  INV_X1 U8456 ( .A(n23568), .ZN(n8205) );
  NAND2_X1 U8457 ( .A1(n7689), .A2(n22586), .ZN(n23447) );
  AND2_X1 U8459 ( .A1(n51123), .A2(n21948), .ZN(n2930) );
  AND2_X1 U8460 ( .A1(n21948), .A2(n23153), .ZN(n19592) );
  OR2_X1 U8461 ( .A1(n22055), .A2(n23182), .ZN(n22535) );
  AND3_X1 U8462 ( .A1(n17876), .A2(n17877), .A3(n19434), .ZN(n5465) );
  AND3_X1 U8463 ( .A1(n17862), .A2(n17861), .A3(n17863), .ZN(n4144) );
  XNOR2_X1 U8464 ( .A(n18470), .B(n18469), .ZN(n18471) );
  XNOR2_X1 U8465 ( .A(n18458), .B(n6671), .ZN(n6670) );
  INV_X1 U8466 ( .A(n22334), .ZN(n22325) );
  NOR2_X1 U8467 ( .A1(n22412), .A2(n22411), .ZN(n22413) );
  AND2_X1 U8468 ( .A1(n4882), .A2(n23379), .ZN(n20707) );
  XNOR2_X1 U8469 ( .A(n25445), .B(n2623), .ZN(n4614) );
  NOR2_X1 U8470 ( .A1(n19817), .A2(n2256), .ZN(n7266) );
  INV_X1 U8471 ( .A(n22738), .ZN(n23815) );
  AND2_X1 U8472 ( .A1(n1497), .A2(n21810), .ZN(n23784) );
  NOR2_X1 U8473 ( .A1(n21866), .A2(n21860), .ZN(n22956) );
  AND2_X1 U8475 ( .A1(n22979), .A2(n22983), .ZN(n7910) );
  AND2_X1 U8476 ( .A1(n22997), .A2(n22996), .ZN(n3331) );
  OR2_X1 U8477 ( .A1(n22992), .A2(n22993), .ZN(n4132) );
  INV_X1 U8478 ( .A(n22983), .ZN(n22998) );
  INV_X1 U8479 ( .A(n21861), .ZN(n5539) );
  NOR2_X1 U8480 ( .A1(n23427), .A2(n5332), .ZN(n23430) );
  INV_X1 U8481 ( .A(n23424), .ZN(n5332) );
  AND2_X1 U8482 ( .A1(n22101), .A2(n24034), .ZN(n23666) );
  AND2_X1 U8483 ( .A1(n24026), .A2(n24041), .ZN(n22097) );
  AOI21_X1 U8484 ( .B1(n22640), .B2(n23076), .A(n5178), .ZN(n22647) );
  AND3_X1 U8485 ( .A1(n52155), .A2(n23066), .A3(n23075), .ZN(n5178) );
  NAND4_X1 U8486 ( .A1(n6063), .A2(n23594), .A3(n20559), .A4(n20558), .ZN(
        n24213) );
  OR2_X1 U8488 ( .A1(n21122), .A2(n21767), .ZN(n21770) );
  OAI21_X1 U8489 ( .B1(n8214), .B2(n8215), .A(n23166), .ZN(n8213) );
  AND3_X1 U8490 ( .A1(n23186), .A2(n23180), .A3(n23181), .ZN(n4230) );
  NAND4_X1 U8492 ( .A1(n15634), .A2(n8556), .A3(n5748), .A4(n15635), .ZN(n4973) );
  NOR2_X1 U8493 ( .A1(n2376), .A2(n2234), .ZN(n7619) );
  INV_X1 U8494 ( .A(n21810), .ZN(n21823) );
  INV_X1 U8495 ( .A(n22687), .ZN(n22688) );
  INV_X1 U8496 ( .A(n22275), .ZN(n22274) );
  OR2_X1 U8497 ( .A1(n22236), .A2(n23536), .ZN(n22237) );
  INV_X1 U8498 ( .A(n22068), .ZN(n8431) );
  AND3_X1 U8499 ( .A1(n22067), .A2(n22668), .A3(n5447), .ZN(n8432) );
  OAI21_X1 U8500 ( .B1(n2279), .B2(n3055), .A(n23166), .ZN(n22066) );
  NOR2_X1 U8502 ( .A1(n3762), .A2(n23537), .ZN(n3761) );
  AND2_X1 U8503 ( .A1(n23693), .A2(n5415), .ZN(n3759) );
  AND3_X1 U8504 ( .A1(n3425), .A2(n7111), .A3(n19566), .ZN(n19570) );
  OAI22_X1 U8506 ( .A1(n7520), .A2(n5896), .B1(n21083), .B2(n7519), .ZN(n7521)
         );
  INV_X1 U8507 ( .A(n7528), .ZN(n7352) );
  NAND4_X1 U8509 ( .A1(n21645), .A2(n23127), .A3(n24111), .A4(n24117), .ZN(
        n21679) );
  AND2_X1 U8510 ( .A1(n17514), .A2(n23329), .ZN(n4254) );
  INV_X1 U8511 ( .A(n24736), .ZN(n3669) );
  AND2_X1 U8513 ( .A1(n5259), .A2(n50990), .ZN(n7214) );
  AND3_X1 U8514 ( .A1(n23163), .A2(n6623), .A3(n7043), .ZN(n6622) );
  OR2_X1 U8517 ( .A1(n30664), .A2(n30661), .ZN(n2798) );
  AND3_X1 U8518 ( .A1(n23633), .A2(n20855), .A3(n20854), .ZN(n4658) );
  XNOR2_X1 U8519 ( .A(n28095), .B(n28094), .ZN(n8406) );
  XNOR2_X1 U8520 ( .A(n7229), .B(n28114), .ZN(n5693) );
  OAI21_X1 U8521 ( .B1(n27577), .B2(n3783), .A(n27679), .ZN(n26812) );
  OR2_X1 U8522 ( .A1(n29719), .A2(n28982), .ZN(n28983) );
  OR2_X1 U8523 ( .A1(n51489), .A2(n30346), .ZN(n28783) );
  AND2_X1 U8524 ( .A1(n514), .A2(n29764), .ZN(n5390) );
  XNOR2_X1 U8525 ( .A(n25126), .B(n25316), .ZN(n30179) );
  INV_X1 U8526 ( .A(n25317), .ZN(n25316) );
  INV_X1 U8527 ( .A(n27654), .ZN(n27653) );
  OR2_X1 U8528 ( .A1(n27067), .A2(n2642), .ZN(n6867) );
  INV_X1 U8529 ( .A(n28067), .ZN(n7899) );
  INV_X1 U8530 ( .A(n28508), .ZN(n29800) );
  INV_X1 U8532 ( .A(n28903), .ZN(n27128) );
  NOR2_X1 U8533 ( .A1(n27668), .A2(n3765), .ZN(n26950) );
  INV_X1 U8534 ( .A(n27067), .ZN(n26933) );
  INV_X1 U8535 ( .A(n26815), .ZN(n26814) );
  AND2_X1 U8536 ( .A1(n26775), .A2(n6449), .ZN(n26810) );
  AND2_X1 U8537 ( .A1(n27856), .A2(n3124), .ZN(n25842) );
  NOR2_X1 U8538 ( .A1(n29187), .A2(n4965), .ZN(n29189) );
  INV_X1 U8539 ( .A(n31624), .ZN(n4907) );
  OR2_X1 U8540 ( .A1(n29918), .A2(n3302), .ZN(n29920) );
  OR2_X1 U8541 ( .A1(n51746), .A2(n29867), .ZN(n28739) );
  OR2_X1 U8542 ( .A1(n6916), .A2(n29698), .ZN(n29862) );
  AND2_X1 U8543 ( .A1(n6708), .A2(n29153), .ZN(n27147) );
  INV_X1 U8544 ( .A(n29156), .ZN(n6708) );
  AND2_X1 U8545 ( .A1(n7783), .A2(n26745), .ZN(n7782) );
  INV_X1 U8546 ( .A(n29327), .ZN(n29324) );
  INV_X1 U8547 ( .A(n27918), .ZN(n30267) );
  INV_X1 U8548 ( .A(n26346), .ZN(n4380) );
  AND2_X1 U8549 ( .A1(n26723), .A2(n26066), .ZN(n4435) );
  NAND4_X1 U8550 ( .A1(n26201), .A2(n26200), .A3(n26199), .A4(n26198), .ZN(
        n26202) );
  XNOR2_X1 U8553 ( .A(n25390), .B(n25092), .ZN(n6643) );
  OR2_X1 U8554 ( .A1(n29123), .A2(n51114), .ZN(n4775) );
  AND2_X1 U8556 ( .A1(n30227), .A2(n29248), .ZN(n28664) );
  INV_X1 U8557 ( .A(n30873), .ZN(n7667) );
  AND3_X1 U8558 ( .A1(n26086), .A2(n26082), .A3(n26081), .ZN(n2928) );
  INV_X1 U8559 ( .A(n3783), .ZN(n26818) );
  INV_X1 U8560 ( .A(n30263), .ZN(n25415) );
  INV_X1 U8562 ( .A(n29185), .ZN(n27924) );
  AND2_X1 U8564 ( .A1(n29255), .A2(n29252), .ZN(n7391) );
  INV_X1 U8565 ( .A(n32874), .ZN(n7232) );
  AND3_X1 U8566 ( .A1(n6800), .A2(n26655), .A3(n26656), .ZN(n26665) );
  AND2_X1 U8567 ( .A1(n8418), .A2(n8417), .ZN(n8425) );
  OAI21_X1 U8568 ( .B1(n28710), .B2(n28711), .A(n8419), .ZN(n8418) );
  INV_X1 U8569 ( .A(n27015), .ZN(n7972) );
  INV_X1 U8570 ( .A(n32211), .ZN(n32209) );
  OR2_X1 U8571 ( .A1(n32194), .A2(n32211), .ZN(n32201) );
  INV_X1 U8572 ( .A(n32487), .ZN(n8344) );
  AND2_X1 U8573 ( .A1(n29437), .A2(n747), .ZN(n29454) );
  AND2_X1 U8574 ( .A1(n31067), .A2(n30924), .ZN(n30082) );
  OR2_X1 U8575 ( .A1(n29848), .A2(n27164), .ZN(n7645) );
  OAI21_X1 U8576 ( .B1(n28760), .B2(n28759), .A(n30384), .ZN(n5978) );
  OR2_X1 U8577 ( .A1(n27107), .A2(n6764), .ZN(n26622) );
  XNOR2_X1 U8578 ( .A(n25143), .B(n27396), .ZN(n7663) );
  AND2_X1 U8579 ( .A1(n30296), .A2(n28143), .ZN(n7604) );
  OR2_X1 U8580 ( .A1(n29998), .A2(n29096), .ZN(n30003) );
  NOR2_X1 U8581 ( .A1(n32882), .A2(n33026), .ZN(n5497) );
  AND2_X1 U8582 ( .A1(n30342), .A2(n29761), .ZN(n3722) );
  AND2_X1 U8583 ( .A1(n29766), .A2(n30343), .ZN(n3723) );
  AOI21_X1 U8584 ( .B1(n28798), .B2(n30407), .A(n3301), .ZN(n7691) );
  INV_X1 U8585 ( .A(n32299), .ZN(n4434) );
  NOR2_X1 U8588 ( .A1(n32356), .A2(n3703), .ZN(n32441) );
  OAI21_X1 U8589 ( .B1(n27742), .B2(n5276), .A(n29467), .ZN(n27771) );
  AOI21_X1 U8590 ( .B1(n27767), .B2(n27766), .A(n4298), .ZN(n27769) );
  AOI21_X1 U8591 ( .B1(n27683), .B2(n27684), .A(n2409), .ZN(n6283) );
  OAI21_X1 U8592 ( .B1(n27703), .B2(n3799), .A(n27702), .ZN(n6014) );
  NOR2_X1 U8593 ( .A1(n6016), .A2(n27699), .ZN(n6015) );
  INV_X1 U8594 ( .A(n31422), .ZN(n31146) );
  INV_X1 U8595 ( .A(n32909), .ZN(n6270) );
  OAI21_X1 U8596 ( .B1(n2845), .B2(n2844), .A(n29557), .ZN(n26686) );
  AND2_X1 U8597 ( .A1(n31033), .A2(n31043), .ZN(n4715) );
  AND2_X1 U8598 ( .A1(n30743), .A2(n30742), .ZN(n3967) );
  OR2_X1 U8600 ( .A1(n29677), .A2(n30873), .ZN(n30881) );
  AND4_X1 U8601 ( .A1(n26740), .A2(n26736), .A3(n29417), .A4(n29431), .ZN(
        n7682) );
  NAND2_X1 U8602 ( .A1(n26734), .A2(n26735), .ZN(n7681) );
  AND2_X1 U8603 ( .A1(n28161), .A2(n6244), .ZN(n7333) );
  INV_X1 U8604 ( .A(n26501), .ZN(n30293) );
  INV_X1 U8605 ( .A(n32719), .ZN(n32316) );
  OR2_X1 U8606 ( .A1(n26329), .A2(n2912), .ZN(n6079) );
  AOI22_X1 U8607 ( .A1(n29547), .A2(n27048), .B1(n5696), .B2(n29541), .ZN(
        n27063) );
  INV_X1 U8609 ( .A(n30073), .ZN(n31115) );
  INV_X1 U8610 ( .A(n32125), .ZN(n3096) );
  OR2_X1 U8611 ( .A1(n27072), .A2(n27652), .ZN(n8331) );
  AND2_X1 U8613 ( .A1(n30282), .A2(n2881), .ZN(n27110) );
  AND3_X1 U8614 ( .A1(n29553), .A2(n29552), .A3(n2518), .ZN(n7788) );
  INV_X1 U8615 ( .A(n4715), .ZN(n3581) );
  OR2_X1 U8616 ( .A1(n31668), .A2(n2091), .ZN(n32694) );
  INV_X1 U8617 ( .A(n31986), .ZN(n32508) );
  AND2_X1 U8618 ( .A1(n32960), .A2(n32957), .ZN(n8125) );
  OR2_X1 U8619 ( .A1(n32759), .A2(n32771), .ZN(n3339) );
  AND2_X1 U8620 ( .A1(n29506), .A2(n26983), .ZN(n7292) );
  OAI21_X1 U8621 ( .B1(n29277), .B2(n51116), .A(n2353), .ZN(n3125) );
  INV_X1 U8622 ( .A(n27678), .ZN(n27582) );
  AND2_X1 U8623 ( .A1(n27674), .A2(n27676), .ZN(n5339) );
  INV_X1 U8624 ( .A(n29684), .ZN(n31097) );
  NOR2_X1 U8625 ( .A1(n30593), .A2(n30598), .ZN(n31089) );
  NOR2_X1 U8626 ( .A1(n30593), .A2(n30912), .ZN(n31099) );
  INV_X1 U8627 ( .A(n31624), .ZN(n31638) );
  INV_X1 U8628 ( .A(n8272), .ZN(n8359) );
  OR2_X1 U8630 ( .A1(n27563), .A2(n30766), .ZN(n3662) );
  AND3_X1 U8631 ( .A1(n3225), .A2(n31496), .A3(n722), .ZN(n31495) );
  INV_X1 U8632 ( .A(n29622), .ZN(n2984) );
  AND2_X1 U8633 ( .A1(n28150), .A2(n3868), .ZN(n3867) );
  AOI22_X1 U8634 ( .A1(n7602), .A2(n3870), .B1(n28153), .B2(n28546), .ZN(n3869) );
  INV_X1 U8636 ( .A(n29609), .ZN(n5682) );
  INV_X1 U8637 ( .A(n31454), .ZN(n3847) );
  OR2_X1 U8638 ( .A1(n30797), .A2(n30798), .ZN(n6791) );
  NOR2_X1 U8639 ( .A1(n32765), .A2(n32960), .ZN(n6042) );
  OR2_X1 U8640 ( .A1(n32175), .A2(n32965), .ZN(n3811) );
  NOR2_X1 U8641 ( .A1(n5182), .A2(n26699), .ZN(n26704) );
  INV_X1 U8642 ( .A(n30740), .ZN(n30361) );
  NOR2_X1 U8643 ( .A1(n7040), .A2(n32299), .ZN(n7041) );
  NOR2_X1 U8645 ( .A1(n32214), .A2(n32210), .ZN(n32204) );
  NOR2_X1 U8646 ( .A1(n29626), .A2(n32491), .ZN(n2820) );
  NOR2_X1 U8647 ( .A1(n4100), .A2(n6539), .ZN(n8745) );
  AND3_X1 U8648 ( .A1(n32618), .A2(n51471), .A3(n31558), .ZN(n6539) );
  AND3_X1 U8649 ( .A1(n29506), .A2(n29539), .A3(n8740), .ZN(n3259) );
  AND2_X1 U8650 ( .A1(n31512), .A2(n30925), .ZN(n30081) );
  AND2_X1 U8651 ( .A1(n6836), .A2(n26729), .ZN(n4046) );
  INV_X1 U8652 ( .A(n32608), .ZN(n31471) );
  OR2_X1 U8653 ( .A1(n30748), .A2(n29886), .ZN(n28778) );
  OAI21_X1 U8654 ( .B1(n26474), .B2(n28905), .A(n6547), .ZN(n26482) );
  AND3_X1 U8655 ( .A1(n30679), .A2(n30678), .A3(n7804), .ZN(n30680) );
  INV_X1 U8656 ( .A(n36685), .ZN(n36857) );
  AND2_X1 U8657 ( .A1(n26327), .A2(n26319), .ZN(n4679) );
  INV_X1 U8658 ( .A(n8536), .ZN(n32417) );
  AND3_X1 U8659 ( .A1(n5030), .A2(n29786), .A3(n5029), .ZN(n5028) );
  XNOR2_X1 U8660 ( .A(n34156), .B(n34896), .ZN(n34359) );
  OR2_X1 U8661 ( .A1(n32732), .A2(n32724), .ZN(n32718) );
  XNOR2_X1 U8662 ( .A(n34360), .B(n32644), .ZN(n35282) );
  OR2_X1 U8663 ( .A1(n30428), .A2(n30433), .ZN(n6772) );
  AOI21_X1 U8664 ( .B1(n30437), .B2(n30438), .A(n6404), .ZN(n30439) );
  OR2_X1 U8665 ( .A1(n31658), .A2(n32327), .ZN(n5217) );
  INV_X1 U8666 ( .A(n32326), .ZN(n32325) );
  INV_X1 U8668 ( .A(n515), .ZN(n33386) );
  INV_X1 U8669 ( .A(n31892), .ZN(n29992) );
  AND2_X1 U8670 ( .A1(n6302), .A2(n6301), .ZN(n6300) );
  XNOR2_X1 U8671 ( .A(n34466), .B(n33753), .ZN(n35510) );
  XNOR2_X1 U8672 ( .A(n34425), .B(n36818), .ZN(n37019) );
  XNOR2_X1 U8674 ( .A(n6833), .B(n6832), .ZN(n35409) );
  INV_X1 U8675 ( .A(n37420), .ZN(n6637) );
  INV_X1 U8676 ( .A(n38562), .ZN(n38198) );
  INV_X1 U8677 ( .A(n36428), .ZN(n8090) );
  INV_X1 U8678 ( .A(n68), .ZN(n5989) );
  INV_X1 U8680 ( .A(n35530), .ZN(n3596) );
  OR2_X1 U8681 ( .A1(n37484), .A2(n37439), .ZN(n36159) );
  OR2_X1 U8683 ( .A1(n37893), .A2(n37894), .ZN(n38994) );
  XNOR2_X1 U8684 ( .A(n35402), .B(n3426), .ZN(n38340) );
  XNOR2_X1 U8685 ( .A(n34887), .B(n37151), .ZN(n34905) );
  NAND2_X1 U8686 ( .A1(n36781), .A2(n2100), .ZN(n39266) );
  AND2_X1 U8687 ( .A1(n696), .A2(n36459), .ZN(n35875) );
  XNOR2_X1 U8688 ( .A(n34044), .B(n2315), .ZN(n35348) );
  INV_X1 U8689 ( .A(n37667), .ZN(n37670) );
  AND4_X1 U8690 ( .A1(n7914), .A2(n7913), .A3(n7915), .A4(n7912), .ZN(n37625)
         );
  AND2_X1 U8691 ( .A1(n2741), .A2(n37624), .ZN(n7913) );
  OR2_X1 U8692 ( .A1(n38283), .A2(n37623), .ZN(n7912) );
  AND2_X1 U8693 ( .A1(n36492), .A2(n36012), .ZN(n2722) );
  AND2_X1 U8694 ( .A1(n39002), .A2(n39399), .ZN(n7407) );
  OR2_X1 U8695 ( .A1(n36472), .A2(n36558), .ZN(n36478) );
  AND2_X1 U8696 ( .A1(n36494), .A2(n35315), .ZN(n4300) );
  INV_X1 U8697 ( .A(n37977), .ZN(n36531) );
  INV_X1 U8698 ( .A(n5987), .ZN(n35431) );
  INV_X1 U8699 ( .A(n36161), .ZN(n8315) );
  INV_X1 U8700 ( .A(n36159), .ZN(n38515) );
  AND2_X1 U8701 ( .A1(n38199), .A2(n5312), .ZN(n6024) );
  OAI21_X1 U8702 ( .B1(n38592), .B2(n38164), .A(n7546), .ZN(n35690) );
  NOR3_X1 U8703 ( .A1(n38584), .A2(n38593), .A3(n38599), .ZN(n7546) );
  INV_X1 U8704 ( .A(n39483), .ZN(n39473) );
  OR2_X1 U8705 ( .A1(n38014), .A2(n35028), .ZN(n7072) );
  INV_X1 U8706 ( .A(n38475), .ZN(n38481) );
  AND2_X1 U8707 ( .A1(n2855), .A2(n40446), .ZN(n6852) );
  INV_X1 U8708 ( .A(n37569), .ZN(n38153) );
  AND2_X1 U8710 ( .A1(n3768), .A2(n40727), .ZN(n3682) );
  OR2_X1 U8711 ( .A1(n41902), .A2(n41316), .ZN(n3770) );
  OR2_X1 U8713 ( .A1(n38492), .A2(n38496), .ZN(n4062) );
  OR2_X1 U8714 ( .A1(n37384), .A2(n37385), .ZN(n2739) );
  OR2_X1 U8715 ( .A1(n35960), .A2(n3590), .ZN(n35963) );
  AND2_X1 U8716 ( .A1(n39377), .A2(n51102), .ZN(n4523) );
  OR2_X1 U8717 ( .A1(n39285), .A2(n39284), .ZN(n7021) );
  INV_X1 U8718 ( .A(n39647), .ZN(n40336) );
  NOR2_X1 U8719 ( .A1(n41539), .A2(n41395), .ZN(n40932) );
  AND2_X1 U8721 ( .A1(n3577), .A2(n38998), .ZN(n37884) );
  INV_X1 U8722 ( .A(n34906), .ZN(n3577) );
  NOR2_X1 U8723 ( .A1(n36604), .A2(n36430), .ZN(n34930) );
  OR2_X1 U8724 ( .A1(n39273), .A2(n5262), .ZN(n39269) );
  INV_X1 U8725 ( .A(n36115), .ZN(n37415) );
  AND2_X1 U8726 ( .A1(n37541), .A2(n37400), .ZN(n5805) );
  INV_X1 U8727 ( .A(n38535), .ZN(n38521) );
  OR2_X1 U8728 ( .A1(n38053), .A2(n38054), .ZN(n7515) );
  OR2_X1 U8729 ( .A1(n38056), .A2(n38050), .ZN(n38051) );
  INV_X1 U8730 ( .A(n38335), .ZN(n38332) );
  AND3_X1 U8732 ( .A1(n39337), .A2(n34691), .A3(n37778), .ZN(n4753) );
  OAI21_X1 U8733 ( .B1(n36542), .B2(n8016), .A(n37957), .ZN(n8015) );
  INV_X1 U8734 ( .A(n39097), .ZN(n38428) );
  OR2_X1 U8735 ( .A1(n41319), .A2(n41902), .ZN(n40732) );
  AND2_X1 U8736 ( .A1(n36056), .A2(n36055), .ZN(n7506) );
  NOR2_X1 U8737 ( .A1(n40940), .A2(n40939), .ZN(n5216) );
  AND2_X1 U8738 ( .A1(n41096), .A2(n41642), .ZN(n40623) );
  OR2_X1 U8739 ( .A1(n39101), .A2(n40014), .ZN(n37848) );
  AND2_X1 U8740 ( .A1(n6749), .A2(n39312), .ZN(n4338) );
  AND2_X1 U8741 ( .A1(n40388), .A2(n41150), .ZN(n4111) );
  NAND4_X1 U8742 ( .A1(n3158), .A2(n3157), .A3(n5603), .A4(n3156), .ZN(n8256)
         );
  AND2_X1 U8743 ( .A1(n38315), .A2(n39295), .ZN(n5603) );
  AND2_X1 U8744 ( .A1(n38316), .A2(n38320), .ZN(n3158) );
  AND2_X1 U8746 ( .A1(n36355), .A2(n36356), .ZN(n3434) );
  INV_X1 U8747 ( .A(n41352), .ZN(n8123) );
  AND2_X1 U8748 ( .A1(n36007), .A2(n36006), .ZN(n4367) );
  AND2_X1 U8750 ( .A1(n40009), .A2(n39094), .ZN(n6885) );
  AND2_X1 U8751 ( .A1(n41356), .A2(n41352), .ZN(n40358) );
  NOR2_X1 U8752 ( .A1(n40835), .A2(n40838), .ZN(n39515) );
  AND2_X1 U8753 ( .A1(n6114), .A2(n40503), .ZN(n3390) );
  INV_X1 U8754 ( .A(n40730), .ZN(n4703) );
  AND3_X1 U8755 ( .A1(n7401), .A2(n36345), .A3(n7399), .ZN(n7397) );
  INV_X1 U8756 ( .A(n36161), .ZN(n38522) );
  INV_X1 U8757 ( .A(n40662), .ZN(n40669) );
  AND2_X1 U8758 ( .A1(n35714), .A2(n35713), .ZN(n35715) );
  OR2_X1 U8759 ( .A1(n43669), .A2(n3550), .ZN(n40633) );
  INV_X1 U8760 ( .A(n40566), .ZN(n39653) );
  AND2_X1 U8761 ( .A1(n40458), .A2(n2855), .ZN(n40461) );
  AND2_X2 U8762 ( .A1(n2557), .A2(n36435), .ZN(n39955) );
  OR2_X1 U8763 ( .A1(n41353), .A2(n38740), .ZN(n38745) );
  AND3_X1 U8764 ( .A1(n6442), .A2(n6441), .A3(n36378), .ZN(n6440) );
  AOI22_X1 U8765 ( .A1(n38028), .A2(n36374), .B1(n6437), .B2(n38037), .ZN(
        n6436) );
  AND2_X1 U8766 ( .A1(n7225), .A2(n36366), .ZN(n7224) );
  INV_X1 U8767 ( .A(n36368), .ZN(n7223) );
  OR2_X1 U8768 ( .A1(n36367), .A2(n6541), .ZN(n6540) );
  INV_X1 U8769 ( .A(n41902), .ZN(n41329) );
  OR2_X1 U8770 ( .A1(n40633), .A2(n38815), .ZN(n41793) );
  AND2_X1 U8771 ( .A1(n35945), .A2(n35938), .ZN(n4205) );
  INV_X1 U8774 ( .A(n40729), .ZN(n39818) );
  AND3_X1 U8775 ( .A1(n39256), .A2(n39255), .A3(n39257), .ZN(n6334) );
  AND2_X1 U8776 ( .A1(n42441), .A2(n596), .ZN(n36286) );
  INV_X1 U8777 ( .A(n36057), .ZN(n4128) );
  INV_X1 U8778 ( .A(n34656), .ZN(n36427) );
  OR2_X1 U8779 ( .A1(n39098), .A2(n39099), .ZN(n40000) );
  INV_X1 U8780 ( .A(n38728), .ZN(n39302) );
  AND2_X1 U8781 ( .A1(n39259), .A2(n39019), .ZN(n37941) );
  AND2_X1 U8782 ( .A1(n6995), .A2(n37530), .ZN(n2934) );
  AND3_X1 U8783 ( .A1(n37695), .A2(n37696), .A3(n4105), .ZN(n37705) );
  INV_X1 U8784 ( .A(n8494), .ZN(n7818) );
  OAI21_X1 U8785 ( .B1(n37578), .B2(n37577), .A(n37576), .ZN(n7308) );
  AND2_X1 U8786 ( .A1(n37583), .A2(n37582), .ZN(n7307) );
  AND2_X1 U8787 ( .A1(n37599), .A2(n37601), .ZN(n8339) );
  AOI21_X1 U8788 ( .B1(n6938), .B2(n6940), .A(n40617), .ZN(n6939) );
  AND2_X1 U8790 ( .A1(n39216), .A2(n39215), .ZN(n5556) );
  OR2_X1 U8791 ( .A1(n36527), .A2(n3281), .ZN(n36079) );
  AND3_X1 U8792 ( .A1(n40280), .A2(n5071), .A3(n40083), .ZN(n5070) );
  AND2_X1 U8793 ( .A1(n41084), .A2(n41079), .ZN(n38875) );
  OR2_X1 U8794 ( .A1(n40615), .A2(n7637), .ZN(n7636) );
  NOR2_X1 U8795 ( .A1(n41975), .A2(n41642), .ZN(n7637) );
  AND2_X1 U8796 ( .A1(n41645), .A2(n41101), .ZN(n8108) );
  NOR2_X1 U8798 ( .A1(n41230), .A2(n41673), .ZN(n3858) );
  INV_X1 U8799 ( .A(n39316), .ZN(n3861) );
  NOR2_X1 U8800 ( .A1(n41243), .A2(n331), .ZN(n41248) );
  INV_X1 U8801 ( .A(n39943), .ZN(n39937) );
  INV_X1 U8802 ( .A(n8256), .ZN(n40525) );
  AND2_X1 U8803 ( .A1(n40098), .A2(n39587), .ZN(n5460) );
  AND3_X1 U8804 ( .A1(n41231), .A2(n2743), .A3(n41234), .ZN(n41669) );
  INV_X1 U8805 ( .A(n39157), .ZN(n7701) );
  NAND3_X2 U8806 ( .A1(n4094), .A2(n36043), .A3(n36041), .ZN(n40120) );
  AND2_X1 U8807 ( .A1(n36042), .A2(n36040), .ZN(n4094) );
  XNOR2_X1 U8808 ( .A(n3526), .B(n51100), .ZN(n3582) );
  NOR2_X1 U8809 ( .A1(n7848), .A2(n4954), .ZN(n40154) );
  INV_X1 U8810 ( .A(n40633), .ZN(n40639) );
  INV_X1 U8813 ( .A(n41932), .ZN(n41940) );
  INV_X1 U8814 ( .A(n41245), .ZN(n2743) );
  OR2_X1 U8815 ( .A1(n39316), .A2(n41670), .ZN(n41684) );
  NOR2_X1 U8816 ( .A1(n39140), .A2(n41083), .ZN(n41087) );
  AND3_X1 U8817 ( .A1(n34660), .A2(n37960), .A3(n4969), .ZN(n6597) );
  NAND2_X1 U8818 ( .A1(n45538), .A2(n52070), .ZN(n45542) );
  INV_X1 U8820 ( .A(n46267), .ZN(n44765) );
  XNOR2_X1 U8821 ( .A(n42871), .B(n7578), .ZN(n42886) );
  INV_X1 U8822 ( .A(n7842), .ZN(n46282) );
  INV_X1 U8823 ( .A(n43147), .ZN(n2790) );
  XNOR2_X1 U8824 ( .A(n43049), .B(n2301), .ZN(n46034) );
  INV_X1 U8825 ( .A(n50261), .ZN(n5617) );
  XNOR2_X1 U8826 ( .A(n44975), .B(n5285), .ZN(n4750) );
  INV_X1 U8827 ( .A(n46691), .ZN(n46908) );
  OAI21_X1 U8828 ( .B1(n46676), .B2(n46844), .A(n46842), .ZN(n2992) );
  AND2_X1 U8829 ( .A1(n46918), .A2(n46606), .ZN(n46694) );
  OAI22_X1 U8830 ( .A1(n45764), .A2(n46629), .B1(n45763), .B2(n46630), .ZN(
        n8157) );
  AND2_X1 U8831 ( .A1(n45763), .A2(n44868), .ZN(n5246) );
  AND2_X1 U8832 ( .A1(n45793), .A2(n46572), .ZN(n46707) );
  NAND2_X1 U8833 ( .A1(n41723), .A2(n45188), .ZN(n46744) );
  BUF_X1 U8834 ( .A(n44280), .Z(n45820) );
  OR2_X1 U8835 ( .A1(n44670), .A2(n44669), .ZN(n3571) );
  AND2_X1 U8836 ( .A1(n48410), .A2(n48412), .ZN(n4003) );
  NOR2_X1 U8837 ( .A1(n45547), .A2(n44263), .ZN(n45002) );
  XNOR2_X1 U8838 ( .A(n5435), .B(n41819), .ZN(n5434) );
  INV_X1 U8839 ( .A(n48434), .ZN(n48430) );
  AND2_X1 U8840 ( .A1(n48473), .A2(n8096), .ZN(n48311) );
  AND2_X1 U8841 ( .A1(n5561), .A2(n48437), .ZN(n48443) );
  OR2_X1 U8842 ( .A1(n48248), .A2(n6649), .ZN(n48475) );
  INV_X1 U8843 ( .A(n48479), .ZN(n6649) );
  OR2_X1 U8844 ( .A1(n48485), .A2(n48475), .ZN(n48309) );
  AND2_X1 U8845 ( .A1(n46219), .A2(n46220), .ZN(n4278) );
  XNOR2_X1 U8847 ( .A(n3756), .B(n42939), .ZN(n3755) );
  INV_X1 U8848 ( .A(n49231), .ZN(n49684) );
  INV_X1 U8849 ( .A(n45967), .ZN(n49216) );
  INV_X1 U8850 ( .A(n42886), .ZN(n49247) );
  INV_X1 U8851 ( .A(n49627), .ZN(n7798) );
  OR2_X1 U8852 ( .A1(n49659), .A2(n2726), .ZN(n46027) );
  XNOR2_X1 U8853 ( .A(n7036), .B(n43887), .ZN(n7035) );
  AND2_X1 U8854 ( .A1(n50322), .A2(n47368), .ZN(n50320) );
  INV_X1 U8855 ( .A(n46034), .ZN(n50287) );
  AND2_X1 U8856 ( .A1(n50268), .A2(n50267), .ZN(n50272) );
  INV_X1 U8857 ( .A(n47044), .ZN(n7824) );
  AND2_X1 U8858 ( .A1(n47046), .A2(n50251), .ZN(n50269) );
  AND2_X1 U8859 ( .A1(n47288), .A2(n47030), .ZN(n50349) );
  OR2_X1 U8860 ( .A1(n46810), .A2(n46828), .ZN(n45176) );
  NOR2_X1 U8861 ( .A1(n6992), .A2(n6991), .ZN(n4789) );
  NOR2_X1 U8862 ( .A1(n50331), .A2(n50321), .ZN(n6991) );
  INV_X1 U8863 ( .A(n47161), .ZN(n2753) );
  AND2_X1 U8865 ( .A1(n47574), .A2(n51286), .ZN(n47505) );
  OR2_X1 U8866 ( .A1(n5986), .A2(n47111), .ZN(n46727) );
  OR2_X1 U8867 ( .A1(n46788), .A2(n46787), .ZN(n3473) );
  INV_X1 U8868 ( .A(n6566), .ZN(n46788) );
  OR2_X1 U8869 ( .A1(n51340), .A2(n47599), .ZN(n47591) );
  AND3_X1 U8870 ( .A1(n47745), .A2(n47778), .A3(n47786), .ZN(n45869) );
  OAI21_X1 U8871 ( .B1(n46739), .B2(n46740), .A(n46738), .ZN(n7025) );
  AND2_X1 U8872 ( .A1(n47945), .A2(n52056), .ZN(n47899) );
  OR2_X1 U8873 ( .A1(n48074), .A2(n3076), .ZN(n44442) );
  INV_X1 U8874 ( .A(n44685), .ZN(n48244) );
  INV_X1 U8875 ( .A(n48100), .ZN(n5502) );
  AND3_X1 U8876 ( .A1(n45571), .A2(n45568), .A3(n46317), .ZN(n4179) );
  AND2_X2 U8877 ( .A1(n45536), .A2(n45537), .ZN(n48159) );
  INV_X1 U8878 ( .A(n51318), .ZN(n6987) );
  INV_X1 U8879 ( .A(n48353), .ZN(n4946) );
  OR2_X1 U8880 ( .A1(n6986), .A2(n51318), .ZN(n48366) );
  NOR2_X1 U8881 ( .A1(n51087), .A2(n48368), .ZN(n48364) );
  INV_X1 U8882 ( .A(n48380), .ZN(n8103) );
  AND2_X1 U8883 ( .A1(n48386), .A2(n48382), .ZN(n8102) );
  OAI21_X1 U8884 ( .B1(n48455), .B2(n7275), .A(n51732), .ZN(n48454) );
  OR2_X1 U8885 ( .A1(n8570), .A2(n46444), .ZN(n48458) );
  AND3_X1 U8886 ( .A1(n48470), .A2(n48452), .A3(n48453), .ZN(n8380) );
  NAND4_X1 U8887 ( .A1(n7275), .A2(n48451), .A3(n48455), .A4(n51732), .ZN(
        n48452) );
  NAND4_X1 U8888 ( .A1(n46509), .A2(n46507), .A3(n46508), .A4(n46506), .ZN(
        n47403) );
  INV_X1 U8891 ( .A(n48821), .ZN(n6664) );
  AND2_X1 U8892 ( .A1(n45693), .A2(n45697), .ZN(n3283) );
  AND2_X1 U8893 ( .A1(n46353), .A2(n46344), .ZN(n3633) );
  NOR2_X1 U8894 ( .A1(n45694), .A2(n46277), .ZN(n3634) );
  AOI21_X1 U8895 ( .B1(n45630), .B2(n45629), .A(n6096), .ZN(n45639) );
  INV_X1 U8896 ( .A(n49021), .ZN(n7161) );
  XNOR2_X1 U8897 ( .A(n42317), .B(n43504), .ZN(n42318) );
  INV_X1 U8898 ( .A(n49112), .ZN(n49081) );
  AND2_X1 U8899 ( .A1(n49127), .A2(n49112), .ZN(n49089) );
  INV_X1 U8900 ( .A(n7017), .ZN(n49492) );
  NOR2_X1 U8901 ( .A1(n2297), .A2(n2724), .ZN(n43444) );
  AND2_X1 U8902 ( .A1(n49850), .A2(n49854), .ZN(n49819) );
  AND2_X1 U8903 ( .A1(n6116), .A2(n49667), .ZN(n49652) );
  AND2_X1 U8905 ( .A1(n51480), .A2(n50187), .ZN(n4842) );
  OR2_X1 U8906 ( .A1(n50433), .A2(n50485), .ZN(n50451) );
  OAI211_X1 U8907 ( .C1(n50372), .C2(n50361), .A(n50359), .B(n50360), .ZN(
        n6957) );
  NOR2_X1 U8908 ( .A1(n50371), .A2(n50372), .ZN(n5162) );
  OR2_X1 U8909 ( .A1(n50366), .A2(n6811), .ZN(n6959) );
  OR2_X1 U8910 ( .A1(n50367), .A2(n50364), .ZN(n6960) );
  AND2_X1 U8911 ( .A1(n47014), .A2(n8534), .ZN(n8533) );
  AOI21_X1 U8912 ( .B1(n46965), .B2(n50006), .A(n2280), .ZN(n7880) );
  AND2_X1 U8913 ( .A1(n50641), .A2(n51029), .ZN(n50599) );
  INV_X1 U8914 ( .A(n47152), .ZN(n43683) );
  INV_X1 U8915 ( .A(n50641), .ZN(n50630) );
  INV_X1 U8917 ( .A(n7747), .ZN(n7744) );
  AND2_X1 U8918 ( .A1(n46971), .A2(n3610), .ZN(n46977) );
  NOR2_X1 U8919 ( .A1(n50902), .A2(n50955), .ZN(n8294) );
  OR2_X1 U8920 ( .A1(n49826), .A2(n49850), .ZN(n3549) );
  AND2_X1 U8921 ( .A1(n44709), .A2(n7419), .ZN(n6523) );
  AOI21_X1 U8922 ( .B1(n2686), .B2(n2688), .A(n46394), .ZN(n2685) );
  INV_X1 U8923 ( .A(n50482), .ZN(n50436) );
  INV_X1 U8924 ( .A(Key[173]), .ZN(n7747) );
  AND2_X1 U8925 ( .A1(n11367), .A2(n12117), .ZN(n10701) );
  AND2_X1 U8926 ( .A1(n11032), .A2(n10584), .ZN(n10165) );
  INV_X1 U8927 ( .A(n11376), .ZN(n12117) );
  INV_X1 U8928 ( .A(n12532), .ZN(n7264) );
  INV_X1 U8929 ( .A(n9786), .ZN(n9022) );
  INV_X1 U8931 ( .A(n11630), .ZN(n7812) );
  INV_X1 U8932 ( .A(n11346), .ZN(n12241) );
  INV_X1 U8933 ( .A(n8994), .ZN(n12267) );
  INV_X1 U8934 ( .A(n12243), .ZN(n6928) );
  NOR2_X1 U8935 ( .A1(n6047), .A2(n51433), .ZN(n6571) );
  INV_X1 U8936 ( .A(n12300), .ZN(n9762) );
  AND2_X1 U8937 ( .A1(n10983), .A2(n9787), .ZN(n10989) );
  INV_X1 U8939 ( .A(n10142), .ZN(n4161) );
  INV_X1 U8940 ( .A(n10701), .ZN(n12123) );
  INV_X1 U8941 ( .A(n10279), .ZN(n10671) );
  INV_X1 U8942 ( .A(n9057), .ZN(n12312) );
  INV_X1 U8943 ( .A(n9656), .ZN(n9772) );
  AND2_X1 U8944 ( .A1(n10267), .A2(n10262), .ZN(n10983) );
  INV_X1 U8945 ( .A(n11374), .ZN(n12114) );
  OR2_X1 U8946 ( .A1(n7694), .A2(n12516), .ZN(n7693) );
  AOI21_X1 U8947 ( .B1(n12245), .B2(n6928), .A(n12263), .ZN(n10745) );
  NOR2_X1 U8948 ( .A1(n10778), .A2(n9117), .ZN(n10786) );
  INV_X1 U8949 ( .A(n9185), .ZN(n7541) );
  AND2_X1 U8950 ( .A1(n11126), .A2(n12698), .ZN(n8314) );
  AND2_X1 U8951 ( .A1(n8313), .A2(n8312), .ZN(n2718) );
  AND2_X1 U8952 ( .A1(n10104), .A2(n10509), .ZN(n10106) );
  OAI21_X1 U8953 ( .B1(n10137), .B2(n10138), .A(n10919), .ZN(n7905) );
  AND3_X1 U8954 ( .A1(n9707), .A2(n9706), .A3(n9705), .ZN(n9708) );
  INV_X1 U8955 ( .A(n9548), .ZN(n12597) );
  AND2_X1 U8956 ( .A1(n12610), .A2(n11914), .ZN(n12589) );
  INV_X1 U8957 ( .A(n12710), .ZN(n12712) );
  OR2_X1 U8958 ( .A1(n12699), .A2(n12440), .ZN(n3711) );
  OR2_X1 U8959 ( .A1(n11122), .A2(n3712), .ZN(n12438) );
  OR2_X1 U8961 ( .A1(n6004), .A2(n10968), .ZN(n10119) );
  NOR2_X1 U8962 ( .A1(n11099), .A2(n9109), .ZN(n12535) );
  INV_X1 U8963 ( .A(n15278), .ZN(n14958) );
  INV_X1 U8964 ( .A(n13782), .ZN(n12417) );
  OAI21_X1 U8965 ( .B1(n8099), .B2(n2211), .A(n8098), .ZN(n11067) );
  INV_X1 U8966 ( .A(n9339), .ZN(n11275) );
  INV_X1 U8967 ( .A(n14322), .ZN(n13045) );
  INV_X1 U8968 ( .A(n2690), .ZN(n17246) );
  INV_X1 U8970 ( .A(n14573), .ZN(n8170) );
  INV_X1 U8971 ( .A(n15162), .ZN(n7715) );
  INV_X1 U8972 ( .A(n9573), .ZN(n10424) );
  OR2_X1 U8973 ( .A1(n12727), .A2(n10437), .ZN(n12733) );
  AND2_X1 U8974 ( .A1(n3377), .A2(n12597), .ZN(n11922) );
  INV_X1 U8976 ( .A(n12638), .ZN(n12632) );
  OR2_X1 U8977 ( .A1(n12176), .A2(n4008), .ZN(n9594) );
  INV_X1 U8978 ( .A(n14454), .ZN(n14444) );
  INV_X1 U8980 ( .A(n9921), .ZN(n10619) );
  INV_X1 U8981 ( .A(n10070), .ZN(n10605) );
  AND2_X1 U8982 ( .A1(n11705), .A2(n9926), .ZN(n11714) );
  AND3_X1 U8983 ( .A1(n11692), .A2(n11691), .A3(n11690), .ZN(n11693) );
  OAI21_X1 U8984 ( .B1(n9305), .B2(n11659), .A(n11662), .ZN(n11661) );
  OR2_X1 U8985 ( .A1(n9205), .A2(n10464), .ZN(n7150) );
  INV_X1 U8986 ( .A(n16036), .ZN(n16049) );
  AND2_X1 U8987 ( .A1(n7694), .A2(n12516), .ZN(n5845) );
  NOR2_X1 U8988 ( .A1(n12512), .A2(n12515), .ZN(n6684) );
  NAND4_X1 U8989 ( .A1(n14491), .A2(n11552), .A3(n14813), .A4(n14812), .ZN(
        n3752) );
  INV_X1 U8990 ( .A(n11536), .ZN(n14491) );
  INV_X1 U8991 ( .A(n11874), .ZN(n7356) );
  INV_X1 U8992 ( .A(n11872), .ZN(n3763) );
  OR2_X1 U8993 ( .A1(n12151), .A2(n12160), .ZN(n3451) );
  AND2_X1 U8994 ( .A1(n11322), .A2(n12171), .ZN(n10414) );
  AND2_X1 U8995 ( .A1(n10412), .A2(n11333), .ZN(n5366) );
  INV_X1 U8996 ( .A(n12790), .ZN(n13432) );
  AND2_X1 U8997 ( .A1(n11396), .A2(n5212), .ZN(n6478) );
  OR2_X1 U8998 ( .A1(n8227), .A2(n14311), .ZN(n13818) );
  OR2_X1 U8999 ( .A1(n13295), .A2(n14030), .ZN(n13289) );
  AND2_X1 U9000 ( .A1(n14257), .A2(n15131), .ZN(n13697) );
  INV_X1 U9001 ( .A(n3081), .ZN(n12912) );
  INV_X1 U9002 ( .A(n10449), .ZN(n7529) );
  OR2_X1 U9003 ( .A1(n11986), .A2(n10445), .ZN(n9181) );
  NOR2_X1 U9004 ( .A1(n12777), .A2(n3279), .ZN(n7767) );
  AND2_X1 U9005 ( .A1(n12780), .A2(n13481), .ZN(n3279) );
  OR2_X1 U9006 ( .A1(n10268), .A2(n10262), .ZN(n4175) );
  OR2_X1 U9008 ( .A1(n14160), .A2(n13761), .ZN(n10766) );
  AND2_X1 U9009 ( .A1(n5176), .A2(n13316), .ZN(n3399) );
  OR2_X1 U9010 ( .A1(n12419), .A2(n13173), .ZN(n12018) );
  INV_X1 U9011 ( .A(n15132), .ZN(n8514) );
  AND2_X1 U9012 ( .A1(n15132), .A2(n13697), .ZN(n13700) );
  NOR2_X1 U9013 ( .A1(n16049), .A2(n51018), .ZN(n14520) );
  INV_X1 U9014 ( .A(n13947), .ZN(n6668) );
  AND4_X1 U9015 ( .A1(n12141), .A2(n11423), .A3(n11411), .A4(n10392), .ZN(
        n8427) );
  NAND4_X1 U9016 ( .A1(n11483), .A2(n11482), .A3(n11481), .A4(n11480), .ZN(
        n11558) );
  AND3_X1 U9017 ( .A1(n5254), .A2(n5249), .A3(n5248), .ZN(n5253) );
  NAND3_X1 U9019 ( .A1(n3825), .A2(n3824), .A3(n10188), .ZN(n10208) );
  AND3_X1 U9020 ( .A1(n10189), .A2(n10180), .A3(n10175), .ZN(n3825) );
  OR2_X1 U9021 ( .A1(n15425), .A2(n2640), .ZN(n12031) );
  AND3_X1 U9022 ( .A1(n11799), .A2(n5907), .A3(n13817), .ZN(n5906) );
  INV_X1 U9023 ( .A(n12544), .ZN(n11447) );
  AOI21_X1 U9024 ( .B1(n12698), .B2(n12697), .A(n2156), .ZN(n2581) );
  NAND2_X1 U9025 ( .A1(n2585), .A2(n11933), .ZN(n2583) );
  OR2_X1 U9026 ( .A1(n12499), .A2(n12498), .ZN(n5179) );
  OR2_X1 U9027 ( .A1(n13148), .A2(n14178), .ZN(n14184) );
  NOR2_X1 U9029 ( .A1(n10198), .A2(n2455), .ZN(n6842) );
  NAND4_X1 U9030 ( .A1(n12564), .A2(n12562), .A3(n12580), .A4(n12563), .ZN(
        n2838) );
  INV_X1 U9031 ( .A(n13313), .ZN(n14609) );
  INV_X1 U9032 ( .A(n10208), .ZN(n13142) );
  INV_X1 U9033 ( .A(n14454), .ZN(n3260) );
  AND2_X1 U9034 ( .A1(n8844), .A2(n8845), .ZN(n4498) );
  INV_X1 U9035 ( .A(n9835), .ZN(n6319) );
  INV_X1 U9036 ( .A(n15438), .ZN(n15325) );
  OAI21_X1 U9037 ( .B1(n12437), .B2(n11926), .A(n12705), .ZN(n8470) );
  OR2_X1 U9038 ( .A1(n14547), .A2(n14550), .ZN(n4594) );
  INV_X1 U9039 ( .A(n13346), .ZN(n14543) );
  AND2_X1 U9040 ( .A1(n14030), .A2(n469), .ZN(n4158) );
  AOI22_X1 U9041 ( .A1(n14104), .A2(n14105), .B1(n14446), .B2(n14450), .ZN(
        n14109) );
  AND2_X1 U9042 ( .A1(n11910), .A2(n11897), .ZN(n5803) );
  INV_X1 U9043 ( .A(n18543), .ZN(n17161) );
  OAI22_X1 U9044 ( .A1(n13104), .A2(n13103), .B1(n13102), .B2(n3902), .ZN(
        n13106) );
  INV_X1 U9045 ( .A(n11157), .ZN(n3902) );
  NAND4_X1 U9046 ( .A1(n641), .A2(n13086), .A3(n13091), .A4(n3080), .ZN(n3802)
         );
  INV_X1 U9047 ( .A(n11821), .ZN(n13101) );
  NAND3_X1 U9048 ( .A1(n51369), .A2(n15168), .A3(n14579), .ZN(n5766) );
  INV_X1 U9049 ( .A(n8716), .ZN(n5765) );
  AND2_X1 U9050 ( .A1(n13226), .A2(n639), .ZN(n6641) );
  AOI21_X1 U9051 ( .B1(n8823), .B2(n11037), .A(n3428), .ZN(n8830) );
  NOR2_X1 U9052 ( .A1(n12733), .A2(n11942), .ZN(n6739) );
  OR3_X2 U9053 ( .A1(n3184), .A2(n3182), .A3(n5341), .ZN(n14999) );
  AND2_X1 U9054 ( .A1(n12624), .A2(n12069), .ZN(n5341) );
  AND2_X1 U9055 ( .A1(n14271), .A2(n15131), .ZN(n14998) );
  OR2_X1 U9056 ( .A1(n11874), .A2(n7354), .ZN(n11890) );
  OR2_X1 U9059 ( .A1(n9574), .A2(n6910), .ZN(n6908) );
  NOR2_X1 U9060 ( .A1(n6907), .A2(n2269), .ZN(n6909) );
  INV_X1 U9061 ( .A(n13343), .ZN(n14721) );
  OR2_X1 U9062 ( .A1(n9907), .A2(n10616), .ZN(n6119) );
  AND2_X1 U9064 ( .A1(n9814), .A2(n9815), .ZN(n4427) );
  AND2_X1 U9066 ( .A1(n51018), .A2(n16039), .ZN(n16045) );
  AND2_X1 U9067 ( .A1(n7967), .A2(n11637), .ZN(n7966) );
  INV_X1 U9068 ( .A(n13377), .ZN(n5925) );
  NAND2_X1 U9069 ( .A1(n3511), .A2(n6738), .ZN(n15134) );
  INV_X1 U9070 ( .A(n6739), .ZN(n6738) );
  NOR2_X1 U9071 ( .A1(n14257), .A2(n6737), .ZN(n3511) );
  AOI22_X1 U9072 ( .A1(n2702), .A2(n11000), .B1(n2700), .B2(n10252), .ZN(n5412) );
  INV_X1 U9073 ( .A(n14139), .ZN(n4345) );
  OR2_X1 U9074 ( .A1(n12031), .A2(n14880), .ZN(n15414) );
  AND2_X1 U9075 ( .A1(n10771), .A2(n10772), .ZN(n4169) );
  AND2_X1 U9076 ( .A1(n12761), .A2(n12760), .ZN(n8106) );
  INV_X1 U9077 ( .A(n14983), .ZN(n7802) );
  INV_X1 U9078 ( .A(n11853), .ZN(n7735) );
  OR2_X1 U9079 ( .A1(n10646), .A2(n14345), .ZN(n4231) );
  NOR2_X1 U9080 ( .A1(n11292), .A2(n5461), .ZN(n11301) );
  XNOR2_X1 U9081 ( .A(n17936), .B(n18795), .ZN(n15932) );
  INV_X1 U9083 ( .A(n14233), .ZN(n12921) );
  OR2_X1 U9084 ( .A1(n13220), .A2(n11834), .ZN(n5552) );
  AND2_X1 U9085 ( .A1(n15378), .A2(n15382), .ZN(n11852) );
  AND3_X1 U9086 ( .A1(n8892), .A2(n8893), .A3(n8891), .ZN(n4917) );
  AND3_X1 U9087 ( .A1(n12233), .A2(n7929), .A3(n12239), .ZN(n4011) );
  INV_X1 U9088 ( .A(n11433), .ZN(n14096) );
  XNOR2_X1 U9089 ( .A(n18464), .B(n17297), .ZN(n15454) );
  AND2_X1 U9090 ( .A1(n3349), .A2(n11170), .ZN(n4520) );
  INV_X1 U9091 ( .A(n14713), .ZN(n14716) );
  INV_X1 U9092 ( .A(n13948), .ZN(n13933) );
  INV_X1 U9093 ( .A(n37288), .ZN(n6412) );
  INV_X1 U9094 ( .A(n7756), .ZN(n12957) );
  AND2_X1 U9095 ( .A1(n778), .A2(n17499), .ZN(n18315) );
  XNOR2_X1 U9096 ( .A(n4938), .B(n15685), .ZN(n19673) );
  XNOR2_X1 U9097 ( .A(n18193), .B(n13893), .ZN(n18450) );
  INV_X1 U9098 ( .A(n18041), .ZN(n6332) );
  BUF_X1 U9099 ( .A(n18457), .Z(n18591) );
  OR2_X1 U9100 ( .A1(n18085), .A2(n51705), .ZN(n15535) );
  AND3_X1 U9101 ( .A1(n10911), .A2(n10912), .A3(n10910), .ZN(n6279) );
  XNOR2_X1 U9102 ( .A(n17754), .B(n6099), .ZN(n13267) );
  INV_X1 U9103 ( .A(n16624), .ZN(n6098) );
  INV_X1 U9104 ( .A(n543), .ZN(n3587) );
  XNOR2_X1 U9105 ( .A(n17132), .B(n17131), .ZN(n17195) );
  AOI21_X1 U9106 ( .B1(n14019), .B2(n11047), .A(n4822), .ZN(n6278) );
  XNOR2_X1 U9107 ( .A(n2579), .B(n14847), .ZN(n19258) );
  XNOR2_X1 U9108 ( .A(n17127), .B(n8211), .ZN(n2579) );
  AND3_X1 U9109 ( .A1(n17871), .A2(n8378), .A3(n19425), .ZN(n6529) );
  NOR2_X1 U9110 ( .A1(n20266), .A2(n20270), .ZN(n3371) );
  OAI21_X1 U9111 ( .B1(n6834), .B2(n14147), .A(n13765), .ZN(n7983) );
  INV_X1 U9113 ( .A(n18234), .ZN(n20212) );
  NOR2_X1 U9114 ( .A1(n6224), .A2(n21186), .ZN(n21177) );
  INV_X1 U9115 ( .A(n21181), .ZN(n6224) );
  INV_X1 U9116 ( .A(n19785), .ZN(n21271) );
  OR2_X1 U9117 ( .A1(n51374), .A2(n19410), .ZN(n4340) );
  AND2_X1 U9118 ( .A1(n19404), .A2(n5671), .ZN(n17870) );
  INV_X1 U9119 ( .A(n18085), .ZN(n4516) );
  XNOR2_X1 U9120 ( .A(n14505), .B(n14498), .ZN(n7641) );
  INV_X1 U9121 ( .A(n20678), .ZN(n20675) );
  XNOR2_X1 U9122 ( .A(n17831), .B(n8699), .ZN(n16765) );
  INV_X1 U9123 ( .A(n4960), .ZN(n4385) );
  OAI21_X1 U9124 ( .B1(n6667), .B2(n14231), .A(n14234), .ZN(n6666) );
  AND2_X1 U9125 ( .A1(n14364), .A2(n3460), .ZN(n14375) );
  NOR2_X1 U9126 ( .A1(n14355), .A2(n14354), .ZN(n6074) );
  OR2_X1 U9127 ( .A1(n14357), .A2(n14356), .ZN(n2873) );
  AND2_X1 U9128 ( .A1(n20101), .A2(n20094), .ZN(n17596) );
  INV_X1 U9129 ( .A(n21354), .ZN(n21603) );
  AND2_X1 U9130 ( .A1(n17496), .A2(n633), .ZN(n17532) );
  AND2_X1 U9131 ( .A1(n21463), .A2(n20493), .ZN(n21470) );
  XNOR2_X1 U9132 ( .A(n14679), .B(n15618), .ZN(n20478) );
  INV_X1 U9133 ( .A(n16294), .ZN(n8083) );
  OR2_X1 U9134 ( .A1(n17066), .A2(n51403), .ZN(n7038) );
  AND2_X1 U9135 ( .A1(n51126), .A2(n19544), .ZN(n19049) );
  INV_X1 U9136 ( .A(n20122), .ZN(n20109) );
  INV_X1 U9137 ( .A(n20354), .ZN(n20360) );
  XNOR2_X1 U9138 ( .A(n7270), .B(n18665), .ZN(n8490) );
  OR2_X1 U9140 ( .A1(n21355), .A2(n8490), .ZN(n21361) );
  INV_X1 U9141 ( .A(n20067), .ZN(n4459) );
  INV_X1 U9143 ( .A(n20052), .ZN(n19487) );
  INV_X1 U9144 ( .A(n16211), .ZN(n19499) );
  NOR2_X1 U9145 ( .A1(n17999), .A2(n18000), .ZN(n20471) );
  OR2_X1 U9146 ( .A1(n19388), .A2(n19396), .ZN(n17575) );
  INV_X1 U9147 ( .A(n20078), .ZN(n20076) );
  OR2_X1 U9148 ( .A1(n19143), .A2(n20073), .ZN(n19138) );
  AND2_X1 U9149 ( .A1(n6332), .A2(n19425), .ZN(n19417) );
  INV_X1 U9150 ( .A(n6711), .ZN(n7585) );
  INV_X1 U9151 ( .A(n18043), .ZN(n19412) );
  NAND2_X1 U9152 ( .A1(n6605), .A2(n17873), .ZN(n18043) );
  INV_X1 U9153 ( .A(n51704), .ZN(n8688) );
  AND2_X1 U9154 ( .A1(n15557), .A2(n6282), .ZN(n6281) );
  INV_X1 U9155 ( .A(n18023), .ZN(n18013) );
  INV_X1 U9156 ( .A(n17576), .ZN(n17568) );
  INV_X1 U9157 ( .A(n19801), .ZN(n19711) );
  INV_X1 U9159 ( .A(n21177), .ZN(n19704) );
  NAND2_X1 U9160 ( .A1(n19828), .A2(n19826), .ZN(n3589) );
  NOR2_X1 U9161 ( .A1(n23171), .A2(n22674), .ZN(n23176) );
  OAI211_X1 U9162 ( .C1(n51039), .C2(n19853), .A(n19642), .B(n19640), .ZN(
        n5342) );
  INV_X1 U9163 ( .A(n21654), .ZN(n20277) );
  AND2_X1 U9164 ( .A1(n20132), .A2(n51403), .ZN(n7844) );
  BUF_X1 U9165 ( .A(n16214), .Z(n18303) );
  AND2_X1 U9166 ( .A1(n18303), .A2(n16218), .ZN(n20061) );
  INV_X1 U9167 ( .A(n21382), .ZN(n21385) );
  INV_X1 U9169 ( .A(n20805), .ZN(n7836) );
  INV_X1 U9170 ( .A(n19514), .ZN(n17039) );
  INV_X1 U9171 ( .A(n17194), .ZN(n19522) );
  AND2_X1 U9172 ( .A1(n22107), .A2(n24041), .ZN(n8526) );
  NAND2_X1 U9173 ( .A1(n6721), .A2(n20658), .ZN(n18847) );
  INV_X1 U9174 ( .A(n19047), .ZN(n19544) );
  INV_X1 U9175 ( .A(n17090), .ZN(n19543) );
  OR2_X1 U9176 ( .A1(n19534), .A2(n20114), .ZN(n19047) );
  AND2_X1 U9177 ( .A1(n21286), .A2(n21287), .ZN(n8446) );
  AND2_X1 U9178 ( .A1(n18075), .A2(n19344), .ZN(n4347) );
  NOR2_X1 U9179 ( .A1(n21495), .A2(n2221), .ZN(n20829) );
  AND2_X1 U9180 ( .A1(n22464), .A2(n22471), .ZN(n20523) );
  OR2_X1 U9182 ( .A1(n19032), .A2(n51039), .ZN(n18268) );
  INV_X1 U9183 ( .A(n22851), .ZN(n19603) );
  NOR2_X1 U9184 ( .A1(n23254), .A2(n23247), .ZN(n23243) );
  INV_X1 U9185 ( .A(n412), .ZN(n22116) );
  OR2_X1 U9186 ( .A1(n20242), .A2(n21615), .ZN(n19984) );
  INV_X1 U9187 ( .A(n21639), .ZN(n19978) );
  OR2_X1 U9188 ( .A1(n25064), .A2(n51654), .ZN(n22207) );
  OR2_X1 U9189 ( .A1(n51654), .A2(n52175), .ZN(n22763) );
  OAI21_X1 U9190 ( .B1(n18888), .B2(n18999), .A(n18995), .ZN(n18889) );
  INV_X1 U9191 ( .A(n21360), .ZN(n21358) );
  NOR2_X1 U9192 ( .A1(n21349), .A2(n21364), .ZN(n19294) );
  INV_X1 U9193 ( .A(n21361), .ZN(n21350) );
  INV_X1 U9195 ( .A(n22740), .ZN(n2810) );
  OR2_X1 U9196 ( .A1(n457), .A2(n5415), .ZN(n23701) );
  OR2_X1 U9197 ( .A1(n24291), .A2(n24292), .ZN(n23503) );
  OR2_X1 U9198 ( .A1(n21782), .A2(n758), .ZN(n20534) );
  AND2_X1 U9199 ( .A1(n22144), .A2(n22157), .ZN(n21935) );
  AND2_X1 U9200 ( .A1(n17583), .A2(n17582), .ZN(n3637) );
  INV_X1 U9201 ( .A(n23102), .ZN(n4407) );
  OR2_X1 U9203 ( .A1(n20752), .A2(n20745), .ZN(n19936) );
  INV_X1 U9204 ( .A(n20197), .ZN(n21537) );
  OAI211_X1 U9205 ( .C1(n2861), .C2(n21413), .A(n21566), .B(n2860), .ZN(n19997) );
  INV_X1 U9206 ( .A(n22494), .ZN(n22835) );
  AND2_X1 U9207 ( .A1(n20020), .A2(n2647), .ZN(n2646) );
  OAI21_X1 U9209 ( .B1(n20018), .B2(n20011), .A(n2652), .ZN(n2651) );
  AND2_X1 U9210 ( .A1(n52048), .A2(n21700), .ZN(n19917) );
  OR2_X1 U9211 ( .A1(n21104), .A2(n4140), .ZN(n21707) );
  AND2_X1 U9212 ( .A1(n17558), .A2(n17559), .ZN(n4219) );
  INV_X1 U9213 ( .A(n23360), .ZN(n17074) );
  OAI211_X1 U9214 ( .C1(n20040), .C2(n20043), .A(n17044), .B(n20042), .ZN(
        n17052) );
  INV_X1 U9215 ( .A(n22735), .ZN(n3398) );
  AND3_X1 U9217 ( .A1(n21500), .A2(n21497), .A3(n21498), .ZN(n6206) );
  INV_X1 U9218 ( .A(n22524), .ZN(n23911) );
  INV_X1 U9219 ( .A(n23480), .ZN(n21977) );
  OAI21_X1 U9220 ( .B1(n21981), .B2(n5352), .A(n5351), .ZN(n21990) );
  OR2_X1 U9221 ( .A1(n23479), .A2(n23481), .ZN(n5351) );
  INV_X1 U9222 ( .A(n21877), .ZN(n5006) );
  AND2_X1 U9223 ( .A1(n21893), .A2(n21878), .ZN(n5000) );
  INV_X1 U9225 ( .A(n22784), .ZN(n22789) );
  INV_X1 U9226 ( .A(n22542), .ZN(n4549) );
  INV_X1 U9227 ( .A(n22548), .ZN(n5270) );
  AND3_X1 U9228 ( .A1(n23153), .A2(n23473), .A3(n23157), .ZN(n23470) );
  AND2_X1 U9229 ( .A1(n20417), .A2(n21382), .ZN(n3971) );
  INV_X1 U9230 ( .A(n21155), .ZN(n23570) );
  AND2_X1 U9231 ( .A1(n19304), .A2(n19302), .ZN(n3913) );
  AND2_X1 U9232 ( .A1(n23675), .A2(n8526), .ZN(n24023) );
  INV_X1 U9233 ( .A(n18846), .ZN(n16885) );
  AND2_X1 U9234 ( .A1(n22085), .A2(n23045), .ZN(n3505) );
  INV_X1 U9236 ( .A(n24333), .ZN(n23536) );
  INV_X1 U9237 ( .A(n23535), .ZN(n3822) );
  AND2_X1 U9238 ( .A1(n21723), .A2(n3636), .ZN(n22404) );
  OR2_X1 U9239 ( .A1(n23220), .A2(n18369), .ZN(n3636) );
  AND2_X1 U9240 ( .A1(n22605), .A2(n24187), .ZN(n4060) );
  OR2_X1 U9241 ( .A1(n24242), .A2(n24247), .ZN(n20879) );
  AND2_X1 U9242 ( .A1(n23153), .A2(n23467), .ZN(n8287) );
  NOR2_X1 U9243 ( .A1(n20523), .A2(n3777), .ZN(n3776) );
  INV_X1 U9244 ( .A(n22308), .ZN(n3777) );
  NOR2_X1 U9245 ( .A1(n19734), .A2(n19813), .ZN(n8036) );
  INV_X1 U9246 ( .A(n22639), .ZN(n23613) );
  AOI21_X1 U9247 ( .B1(n7169), .B2(n2262), .A(n19754), .ZN(n22555) );
  NOR2_X1 U9248 ( .A1(n22989), .A2(n22977), .ZN(n7169) );
  OR2_X1 U9249 ( .A1(n22979), .A2(n22983), .ZN(n22562) );
  NOR2_X1 U9250 ( .A1(n24413), .A2(n24409), .ZN(n24106) );
  OR2_X1 U9251 ( .A1(n24283), .A2(n5898), .ZN(n5897) );
  NOR2_X1 U9252 ( .A1(n755), .A2(n52433), .ZN(n21083) );
  NOR2_X1 U9253 ( .A1(n20989), .A2(n21085), .ZN(n7520) );
  OAI21_X1 U9254 ( .B1(n23811), .B2(n22729), .A(n5371), .ZN(n3483) );
  INV_X1 U9256 ( .A(n23871), .ZN(n24185) );
  OR2_X1 U9257 ( .A1(n24074), .A2(n24119), .ZN(n21674) );
  OR2_X1 U9258 ( .A1(n24105), .A2(n23129), .ZN(n23127) );
  NOR2_X1 U9259 ( .A1(n4324), .A2(n21689), .ZN(n4323) );
  AND2_X1 U9260 ( .A1(n18904), .A2(n18905), .ZN(n5534) );
  INV_X1 U9261 ( .A(n22317), .ZN(n23421) );
  NOR2_X1 U9262 ( .A1(n5146), .A2(n5145), .ZN(n5144) );
  AND2_X1 U9263 ( .A1(n24000), .A2(n23987), .ZN(n5116) );
  INV_X1 U9264 ( .A(n22427), .ZN(n23998) );
  INV_X1 U9265 ( .A(n22100), .ZN(n24042) );
  INV_X1 U9266 ( .A(n21715), .ZN(n22190) );
  OAI21_X1 U9267 ( .B1(n18866), .B2(n8298), .A(n498), .ZN(n18881) );
  AND3_X1 U9268 ( .A1(n18880), .A2(n18878), .A3(n18879), .ZN(n4430) );
  OR2_X1 U9270 ( .A1(n23310), .A2(n22249), .ZN(n6134) );
  OR2_X1 U9271 ( .A1(n23317), .A2(n23316), .ZN(n23320) );
  AND2_X1 U9272 ( .A1(n21767), .A2(n24452), .ZN(n22290) );
  AND2_X1 U9273 ( .A1(n23832), .A2(n1942), .ZN(n24160) );
  OR2_X1 U9274 ( .A1(n23599), .A2(n2610), .ZN(n24212) );
  INV_X1 U9275 ( .A(n23598), .ZN(n2610) );
  INV_X1 U9276 ( .A(n22837), .ZN(n6053) );
  NOR2_X1 U9277 ( .A1(n22189), .A2(n21700), .ZN(n5130) );
  INV_X1 U9278 ( .A(n21095), .ZN(n21094) );
  INV_X1 U9279 ( .A(n23992), .ZN(n3912) );
  INV_X1 U9280 ( .A(n22639), .ZN(n3170) );
  INV_X1 U9281 ( .A(n23595), .ZN(n22642) );
  AND2_X1 U9282 ( .A1(n23965), .A2(n23090), .ZN(n4061) );
  AOI22_X1 U9283 ( .A1(n4412), .A2(n4413), .B1(n21015), .B2(n23023), .ZN(n2847) );
  AND4_X1 U9284 ( .A1(n21977), .A2(n7535), .A3(n23489), .A4(n23479), .ZN(n8474) );
  AND2_X1 U9285 ( .A1(n23489), .A2(n21974), .ZN(n8475) );
  NOR2_X1 U9286 ( .A1(n23200), .A2(n24180), .ZN(n24179) );
  AND2_X1 U9287 ( .A1(n22602), .A2(n22603), .ZN(n4799) );
  OR2_X1 U9288 ( .A1(n19577), .A2(n22918), .ZN(n5543) );
  OR2_X1 U9289 ( .A1(n23466), .A2(n23473), .ZN(n23468) );
  OR2_X1 U9290 ( .A1(n22461), .A2(n2083), .ZN(n4718) );
  NOR2_X1 U9291 ( .A1(n23473), .A2(n6010), .ZN(n23156) );
  AND3_X1 U9292 ( .A1(n2996), .A2(n19593), .A3(n19594), .ZN(n19599) );
  OAI211_X1 U9293 ( .C1(n3646), .C2(n22121), .A(n7846), .B(n22118), .ZN(n22412) );
  AND2_X1 U9294 ( .A1(n18369), .A2(n413), .ZN(n3877) );
  AND2_X1 U9295 ( .A1(n22171), .A2(n22172), .ZN(n7940) );
  AND2_X1 U9296 ( .A1(n22337), .A2(n22335), .ZN(n4765) );
  OR2_X1 U9298 ( .A1(n20864), .A2(n22256), .ZN(n20866) );
  OR2_X1 U9299 ( .A1(n23641), .A2(n23950), .ZN(n23956) );
  AND2_X1 U9300 ( .A1(n23641), .A2(n22623), .ZN(n23622) );
  OR2_X1 U9301 ( .A1(n22909), .A2(n22914), .ZN(n5310) );
  NOR2_X1 U9302 ( .A1(n29156), .A2(n27145), .ZN(n5781) );
  XNOR2_X1 U9303 ( .A(n26176), .B(n25365), .ZN(n28361) );
  XNOR2_X1 U9304 ( .A(n28221), .B(n24949), .ZN(n28095) );
  AOI22_X1 U9305 ( .A1(n22896), .A2(n3022), .B1(n21039), .B2(n21038), .ZN(
        n21045) );
  INV_X1 U9306 ( .A(n7350), .ZN(n6601) );
  AND2_X1 U9307 ( .A1(n22949), .A2(n23063), .ZN(n22093) );
  XNOR2_X1 U9309 ( .A(n25798), .B(n51647), .ZN(n27491) );
  INV_X1 U9311 ( .A(n5384), .ZN(n22554) );
  AND2_X1 U9312 ( .A1(n29016), .A2(n28923), .ZN(n7146) );
  INV_X1 U9313 ( .A(n21030), .ZN(n21023) );
  AND2_X1 U9314 ( .A1(n28587), .A2(n3143), .ZN(n25298) );
  INV_X1 U9315 ( .A(n26775), .ZN(n24467) );
  INV_X1 U9316 ( .A(n23112), .ZN(n29851) );
  NOR2_X1 U9318 ( .A1(n8432), .A2(n8431), .ZN(n8430) );
  AND2_X1 U9319 ( .A1(n22897), .A2(n22365), .ZN(n7192) );
  NAND2_X1 U9320 ( .A1(n7973), .A2(n29462), .ZN(n29456) );
  INV_X1 U9321 ( .A(n26763), .ZN(n26760) );
  XNOR2_X1 U9322 ( .A(n26091), .B(n26089), .ZN(n8621) );
  INV_X1 U9323 ( .A(n26761), .ZN(n29556) );
  INV_X1 U9324 ( .A(n26197), .ZN(n29559) );
  NOR2_X1 U9325 ( .A1(n26761), .A2(n8454), .ZN(n8453) );
  OR2_X1 U9326 ( .A1(n29306), .A2(n29291), .ZN(n3407) );
  XNOR2_X1 U9327 ( .A(n24464), .B(n25154), .ZN(n5615) );
  INV_X1 U9328 ( .A(n2158), .ZN(n25075) );
  INV_X1 U9329 ( .A(n29153), .ZN(n6709) );
  OAI211_X1 U9331 ( .C1(n6925), .C2(n20288), .A(n6924), .B(n6923), .ZN(n8081)
         );
  OR2_X1 U9332 ( .A1(n20287), .A2(n43702), .ZN(n6925) );
  NAND2_X1 U9333 ( .A1(n24348), .A2(n29916), .ZN(n27556) );
  INV_X1 U9335 ( .A(n6265), .ZN(n3112) );
  INV_X1 U9336 ( .A(n26575), .ZN(n28056) );
  XNOR2_X1 U9337 ( .A(n23291), .B(n23292), .ZN(n24578) );
  NOR2_X1 U9338 ( .A1(n51706), .A2(n8422), .ZN(n8421) );
  AOI21_X1 U9339 ( .B1(n28710), .B2(n8242), .A(n29183), .ZN(n8419) );
  XNOR2_X1 U9341 ( .A(n24547), .B(n24546), .ZN(n27765) );
  INV_X1 U9343 ( .A(n24092), .ZN(n29940) );
  INV_X1 U9344 ( .A(n29039), .ZN(n27103) );
  NOR2_X1 U9345 ( .A1(n28015), .A2(n28923), .ZN(n4190) );
  OR2_X1 U9346 ( .A1(n29424), .A2(n51679), .ZN(n5141) );
  XNOR2_X1 U9347 ( .A(n25638), .B(n8335), .ZN(n6447) );
  AND2_X1 U9348 ( .A1(n29564), .A2(n27700), .ZN(n6016) );
  INV_X1 U9349 ( .A(n32609), .ZN(n7626) );
  INV_X1 U9350 ( .A(n29691), .ZN(n29690) );
  XNOR2_X1 U9351 ( .A(n7181), .B(n27495), .ZN(n7180) );
  XNOR2_X1 U9353 ( .A(n6719), .B(n25590), .ZN(n28437) );
  INV_X1 U9354 ( .A(n27450), .ZN(n6720) );
  INV_X1 U9355 ( .A(n51693), .ZN(n30458) );
  INV_X1 U9356 ( .A(n29000), .ZN(n29740) );
  OR2_X1 U9357 ( .A1(n27070), .A2(n26945), .ZN(n27068) );
  OR2_X1 U9358 ( .A1(n30724), .A2(n29853), .ZN(n27163) );
  XNOR2_X1 U9359 ( .A(n24840), .B(n2319), .ZN(n30283) );
  INV_X1 U9360 ( .A(n8723), .ZN(n5082) );
  INV_X1 U9361 ( .A(n27113), .ZN(n28551) );
  OR2_X1 U9362 ( .A1(n26288), .A2(n28623), .ZN(n29512) );
  XNOR2_X1 U9363 ( .A(n5679), .B(n5678), .ZN(n5677) );
  NOR2_X1 U9364 ( .A1(n7008), .A2(n2762), .ZN(n7007) );
  XNOR2_X1 U9365 ( .A(n3302), .B(n738), .ZN(n24352) );
  INV_X1 U9366 ( .A(n738), .ZN(n8377) );
  INV_X1 U9367 ( .A(n27562), .ZN(n5768) );
  INV_X1 U9368 ( .A(n24882), .ZN(n30289) );
  OR2_X1 U9369 ( .A1(n30172), .A2(n30168), .ZN(n30173) );
  INV_X1 U9370 ( .A(n547), .ZN(n30314) );
  AND2_X1 U9371 ( .A1(n30177), .A2(n547), .ZN(n3265) );
  INV_X1 U9372 ( .A(n29446), .ZN(n27038) );
  XNOR2_X1 U9373 ( .A(n27119), .B(n3143), .ZN(n27126) );
  INV_X1 U9374 ( .A(n27751), .ZN(n27750) );
  INV_X1 U9375 ( .A(n29550), .ZN(n8455) );
  INV_X1 U9376 ( .A(n31910), .ZN(n7723) );
  INV_X1 U9377 ( .A(n27660), .ZN(n27065) );
  INV_X1 U9378 ( .A(n30296), .ZN(n28548) );
  AND2_X1 U9380 ( .A1(n29350), .A2(n30206), .ZN(n7817) );
  INV_X1 U9381 ( .A(n29187), .ZN(n27930) );
  AND3_X1 U9382 ( .A1(n24776), .A2(n27671), .A3(n27662), .ZN(n27657) );
  INV_X1 U9383 ( .A(n29686), .ZN(n30597) );
  OR2_X1 U9384 ( .A1(n30662), .A2(n27609), .ZN(n4054) );
  NAND4_X1 U9385 ( .A1(n27616), .A2(n8358), .A3(n27626), .A4(n27617), .ZN(
        n8361) );
  AND2_X1 U9387 ( .A1(n28863), .A2(n2499), .ZN(n2706) );
  OAI21_X1 U9388 ( .B1(n30790), .B2(n30780), .A(n2774), .ZN(n30781) );
  AND3_X1 U9389 ( .A1(n30796), .A2(n3341), .A3(n3340), .ZN(n6792) );
  NOR2_X1 U9390 ( .A1(n28923), .A2(n29020), .ZN(n28019) );
  OAI222_X1 U9392 ( .A1(n28797), .A2(n30403), .B1(n30412), .B2(n28189), .C1(
        n28974), .C2(n28973), .ZN(n28190) );
  NOR2_X1 U9393 ( .A1(n30790), .A2(n51723), .ZN(n27409) );
  NOR2_X1 U9394 ( .A1(n32396), .A2(n32402), .ZN(n32404) );
  AND3_X1 U9395 ( .A1(n32816), .A2(n31904), .A3(n2759), .ZN(n2758) );
  AND2_X1 U9396 ( .A1(n32882), .A2(n32874), .ZN(n30969) );
  AND2_X1 U9397 ( .A1(n7082), .A2(n29245), .ZN(n5795) );
  AND2_X1 U9398 ( .A1(n29233), .A2(n29246), .ZN(n5794) );
  AND2_X1 U9399 ( .A1(n31447), .A2(n6188), .ZN(n5864) );
  OR2_X1 U9400 ( .A1(n32661), .A2(n32665), .ZN(n31550) );
  NAND4_X1 U9401 ( .A1(n25479), .A2(n51116), .A3(n377), .A4(n5522), .ZN(n27931) );
  OR2_X1 U9402 ( .A1(n2158), .A2(n6487), .ZN(n27969) );
  INV_X1 U9403 ( .A(n31096), .ZN(n30599) );
  AND2_X1 U9404 ( .A1(n7626), .A2(n32616), .ZN(n8277) );
  AND2_X1 U9405 ( .A1(n27857), .A2(n29498), .ZN(n4117) );
  AND2_X1 U9406 ( .A1(n29479), .A2(n27858), .ZN(n4362) );
  NOR2_X1 U9407 ( .A1(n32351), .A2(n32439), .ZN(n32355) );
  NOR2_X1 U9408 ( .A1(n28022), .A2(n30183), .ZN(n5743) );
  AND3_X1 U9409 ( .A1(n30254), .A2(n30252), .A3(n30253), .ZN(n2866) );
  INV_X1 U9410 ( .A(n30349), .ZN(n3716) );
  INV_X1 U9411 ( .A(n4267), .ZN(n30398) );
  OR2_X1 U9412 ( .A1(n31800), .A2(n31883), .ZN(n31797) );
  NOR2_X1 U9413 ( .A1(n31883), .A2(n3104), .ZN(n31874) );
  AND2_X1 U9414 ( .A1(n31668), .A2(n32691), .ZN(n31660) );
  INV_X1 U9415 ( .A(n30081), .ZN(n5326) );
  INV_X1 U9416 ( .A(n29643), .ZN(n31057) );
  AND2_X1 U9417 ( .A1(n23856), .A2(n23855), .ZN(n3536) );
  AND2_X1 U9420 ( .A1(n30855), .A2(n30857), .ZN(n2872) );
  AND3_X1 U9421 ( .A1(n32139), .A2(n32135), .A3(n32134), .ZN(n8222) );
  INV_X1 U9423 ( .A(n32503), .ZN(n7897) );
  NOR2_X1 U9424 ( .A1(n30877), .A2(n32511), .ZN(n8722) );
  NOR2_X1 U9425 ( .A1(n31535), .A2(n31534), .ZN(n34121) );
  INV_X1 U9426 ( .A(n8082), .ZN(n29171) );
  OR2_X1 U9427 ( .A1(n32821), .A2(n32822), .ZN(n4391) );
  NOR2_X1 U9428 ( .A1(n29287), .A2(n7375), .ZN(n7374) );
  AND2_X1 U9429 ( .A1(n29279), .A2(n51706), .ZN(n7375) );
  INV_X1 U9430 ( .A(n31608), .ZN(n32088) );
  INV_X1 U9431 ( .A(n32118), .ZN(n32131) );
  INV_X1 U9432 ( .A(n32404), .ZN(n5779) );
  OR2_X1 U9433 ( .A1(n33159), .A2(n32075), .ZN(n32069) );
  INV_X1 U9434 ( .A(n33013), .ZN(n33018) );
  OAI211_X1 U9435 ( .C1(n30997), .C2(n722), .A(n30996), .B(n31497), .ZN(n31001) );
  INV_X1 U9437 ( .A(n31489), .ZN(n31273) );
  INV_X1 U9438 ( .A(n32601), .ZN(n32596) );
  INV_X1 U9439 ( .A(n32586), .ZN(n32597) );
  OR2_X1 U9441 ( .A1(n7042), .A2(n8742), .ZN(n28208) );
  OR2_X1 U9442 ( .A1(n8390), .A2(n32761), .ZN(n32524) );
  INV_X1 U9443 ( .A(n31285), .ZN(n31284) );
  AND2_X1 U9444 ( .A1(n31280), .A2(n32394), .ZN(n4851) );
  INV_X1 U9445 ( .A(n32899), .ZN(n8228) );
  AND2_X1 U9446 ( .A1(n5976), .A2(n32908), .ZN(n32547) );
  OR2_X1 U9447 ( .A1(n29107), .A2(n5109), .ZN(n25409) );
  NOR2_X1 U9448 ( .A1(n31466), .A2(n32609), .ZN(n31561) );
  AND2_X1 U9449 ( .A1(n32066), .A2(n32402), .ZN(n6635) );
  OR2_X1 U9450 ( .A1(n714), .A2(n31947), .ZN(n32412) );
  INV_X1 U9451 ( .A(n34405), .ZN(n8248) );
  NOR2_X1 U9452 ( .A1(n3847), .A2(n5868), .ZN(n3846) );
  INV_X1 U9453 ( .A(n32918), .ZN(n32638) );
  AND2_X1 U9454 ( .A1(n8517), .A2(n31385), .ZN(n31010) );
  AND2_X1 U9455 ( .A1(n31676), .A2(n7598), .ZN(n30978) );
  OR2_X1 U9456 ( .A1(n27833), .A2(n6303), .ZN(n6302) );
  OR2_X1 U9457 ( .A1(n32457), .A2(n3237), .ZN(n32721) );
  INV_X1 U9458 ( .A(n6562), .ZN(n6561) );
  OR2_X1 U9459 ( .A1(n27889), .A2(n29329), .ZN(n6873) );
  INV_X1 U9460 ( .A(n31850), .ZN(n32303) );
  OAI21_X1 U9461 ( .B1(n31488), .B2(n31487), .A(n621), .ZN(n31494) );
  OAI21_X1 U9462 ( .B1(n30219), .B2(n30220), .A(n2747), .ZN(n30222) );
  OR2_X1 U9463 ( .A1(n30591), .A2(n30590), .ZN(n30909) );
  NOR2_X1 U9464 ( .A1(n30601), .A2(n29686), .ZN(n31086) );
  OR2_X1 U9466 ( .A1(n30852), .A2(n31030), .ZN(n6321) );
  NOR2_X1 U9467 ( .A1(n30983), .A2(n31680), .ZN(n30023) );
  OR2_X1 U9468 ( .A1(n2878), .A2(n30006), .ZN(n30008) );
  INV_X1 U9469 ( .A(n32175), .ZN(n32766) );
  NOR2_X1 U9470 ( .A1(n32600), .A2(n29618), .ZN(n6344) );
  NOR2_X1 U9471 ( .A1(n32957), .A2(n32760), .ZN(n32961) );
  INV_X1 U9473 ( .A(n32315), .ZN(n31644) );
  INV_X1 U9474 ( .A(n31332), .ZN(n4770) );
  AND2_X1 U9475 ( .A1(n30882), .A2(n31188), .ZN(n32000) );
  AOI21_X1 U9476 ( .B1(n31835), .B2(n32759), .A(n32533), .ZN(n3045) );
  OR2_X1 U9477 ( .A1(n31838), .A2(n3811), .ZN(n3046) );
  XNOR2_X1 U9478 ( .A(n2840), .B(n32997), .ZN(n36983) );
  INV_X1 U9479 ( .A(n35632), .ZN(n2840) );
  AND2_X1 U9480 ( .A1(n31831), .A2(n31832), .ZN(n6463) );
  AND2_X1 U9481 ( .A1(n31522), .A2(n31523), .ZN(n4266) );
  INV_X1 U9482 ( .A(n35749), .ZN(n5999) );
  INV_X1 U9483 ( .A(n5367), .ZN(n33815) );
  INV_X1 U9484 ( .A(n30901), .ZN(n32104) );
  AND3_X1 U9485 ( .A1(n29637), .A2(n5719), .A3(n29634), .ZN(n5718) );
  NAND2_X1 U9486 ( .A1(n29619), .A2(n30513), .ZN(n6243) );
  AND2_X1 U9487 ( .A1(n28726), .A2(n28725), .ZN(n4633) );
  INV_X1 U9488 ( .A(n31886), .ZN(n31799) );
  OR2_X1 U9489 ( .A1(n31028), .A2(n31798), .ZN(n6401) );
  INV_X1 U9490 ( .A(n31885), .ZN(n7838) );
  AND2_X1 U9491 ( .A1(n31789), .A2(n3122), .ZN(n3121) );
  OR2_X1 U9492 ( .A1(n52047), .A2(n3123), .ZN(n3122) );
  INV_X1 U9493 ( .A(n29687), .ZN(n31098) );
  INV_X1 U9494 ( .A(n31089), .ZN(n2944) );
  AND2_X1 U9495 ( .A1(n31638), .A2(n31637), .ZN(n7961) );
  INV_X1 U9496 ( .A(n37040), .ZN(n7271) );
  AND2_X1 U9497 ( .A1(n31497), .A2(n31489), .ZN(n5631) );
  NOR2_X1 U9498 ( .A1(n32601), .A2(n32976), .ZN(n6521) );
  OR2_X1 U9500 ( .A1(n27651), .A2(n2434), .ZN(n2822) );
  NAND3_X1 U9501 ( .A1(n29406), .A2(n29404), .A3(n29405), .ZN(n36847) );
  AND2_X1 U9502 ( .A1(n29596), .A2(n29595), .ZN(n4059) );
  OR2_X1 U9503 ( .A1(n29647), .A2(n30081), .ZN(n4108) );
  INV_X1 U9504 ( .A(n35282), .ZN(n34625) );
  XNOR2_X1 U9505 ( .A(n36758), .B(n35762), .ZN(n35477) );
  OR2_X1 U9506 ( .A1(n27874), .A2(n31424), .ZN(n6306) );
  AND2_X1 U9507 ( .A1(n32430), .A2(n2595), .ZN(n2594) );
  NOR2_X1 U9508 ( .A1(n6746), .A2(n2593), .ZN(n2592) );
  AND2_X1 U9510 ( .A1(n32320), .A2(n32321), .ZN(n5599) );
  INV_X1 U9511 ( .A(n32997), .ZN(n2842) );
  AND2_X1 U9512 ( .A1(n32448), .A2(n32449), .ZN(n3362) );
  INV_X1 U9513 ( .A(n37553), .ZN(n7011) );
  XNOR2_X1 U9514 ( .A(n33644), .B(n33643), .ZN(n5811) );
  AND2_X1 U9515 ( .A1(n32669), .A2(n32670), .ZN(n4573) );
  XNOR2_X1 U9516 ( .A(n37077), .B(n37284), .ZN(n7610) );
  INV_X1 U9517 ( .A(n38138), .ZN(n36341) );
  OR2_X1 U9518 ( .A1(n51429), .A2(n5037), .ZN(n38160) );
  AND2_X1 U9519 ( .A1(n5706), .A2(n28602), .ZN(n5705) );
  NAND4_X1 U9521 ( .A1(n31378), .A2(n3241), .A3(n31376), .A4(n6417), .ZN(n6418) );
  AND2_X1 U9522 ( .A1(n32514), .A2(n32516), .ZN(n5159) );
  XNOR2_X1 U9523 ( .A(n35606), .B(n34553), .ZN(n34726) );
  INV_X1 U9524 ( .A(n34958), .ZN(n7916) );
  INV_X1 U9525 ( .A(n33910), .ZN(n4260) );
  INV_X1 U9526 ( .A(n38323), .ZN(n37664) );
  AOI21_X1 U9527 ( .B1(n37730), .B2(n3738), .A(n3737), .ZN(n3736) );
  INV_X1 U9528 ( .A(n35736), .ZN(n3354) );
  OR2_X1 U9529 ( .A1(n37484), .A2(n617), .ZN(n38534) );
  INV_X1 U9530 ( .A(n37033), .ZN(n39380) );
  AND2_X1 U9531 ( .A1(n37688), .A2(n37219), .ZN(n3311) );
  OR2_X1 U9532 ( .A1(n51487), .A2(n37439), .ZN(n4137) );
  OAI21_X1 U9533 ( .B1(n35157), .B2(n35162), .A(n2661), .ZN(n33175) );
  OAI21_X1 U9534 ( .B1(n38290), .B2(n38271), .A(n38275), .ZN(n2787) );
  INV_X1 U9535 ( .A(n38345), .ZN(n6612) );
  INV_X1 U9536 ( .A(n39367), .ZN(n39189) );
  INV_X1 U9537 ( .A(n39369), .ZN(n38963) );
  AND2_X1 U9538 ( .A1(n36381), .A2(n35154), .ZN(n36384) );
  OAI211_X1 U9539 ( .C1(n38282), .C2(n35424), .A(n2487), .B(n6862), .ZN(n35426) );
  AND2_X1 U9540 ( .A1(n42018), .A2(n41587), .ZN(n7709) );
  INV_X1 U9543 ( .A(n36373), .ZN(n36371) );
  OR2_X1 U9544 ( .A1(n34937), .A2(n5152), .ZN(n34949) );
  OR2_X1 U9545 ( .A1(n36339), .A2(n611), .ZN(n7399) );
  NOR2_X1 U9546 ( .A1(n38056), .A2(n7403), .ZN(n7402) );
  INV_X1 U9547 ( .A(n35457), .ZN(n37372) );
  AND2_X1 U9548 ( .A1(n38562), .A2(n36106), .ZN(n35711) );
  OR2_X1 U9549 ( .A1(n38557), .A2(n51738), .ZN(n35170) );
  INV_X1 U9550 ( .A(n34958), .ZN(n36629) );
  INV_X1 U9551 ( .A(n584), .ZN(n40118) );
  AND2_X1 U9552 ( .A1(n41034), .A2(n41275), .ZN(n40423) );
  NOR2_X1 U9553 ( .A1(n36401), .A2(n51334), .ZN(n6264) );
  OAI21_X1 U9554 ( .B1(n37806), .B2(n37810), .A(n37809), .ZN(n37811) );
  AND3_X1 U9555 ( .A1(n37799), .A2(n38980), .A3(n38977), .ZN(n4997) );
  OR2_X1 U9556 ( .A1(n35942), .A2(n35939), .ZN(n37776) );
  INV_X1 U9557 ( .A(n36186), .ZN(n3070) );
  OR2_X1 U9558 ( .A1(n39206), .A2(n39429), .ZN(n38647) );
  NOR2_X1 U9559 ( .A1(n43327), .A2(n51146), .ZN(n40806) );
  INV_X1 U9560 ( .A(n43666), .ZN(n3550) );
  INV_X1 U9561 ( .A(n40689), .ZN(n38401) );
  NAND2_X1 U9563 ( .A1(n38339), .A2(n38341), .ZN(n2756) );
  INV_X1 U9565 ( .A(n38270), .ZN(n38276) );
  AND2_X1 U9566 ( .A1(n6778), .A2(n6777), .ZN(n6776) );
  AND2_X1 U9567 ( .A1(n3028), .A2(n35148), .ZN(n6782) );
  AND2_X1 U9568 ( .A1(n38566), .A2(n33062), .ZN(n6783) );
  AND2_X1 U9569 ( .A1(n36106), .A2(n481), .ZN(n6781) );
  AND3_X1 U9570 ( .A1(n38530), .A2(n3596), .A3(n38522), .ZN(n3595) );
  INV_X1 U9571 ( .A(n38534), .ZN(n38518) );
  NOR2_X1 U9572 ( .A1(n42205), .A2(n40250), .ZN(n40248) );
  XNOR2_X1 U9573 ( .A(n34251), .B(n34249), .ZN(n5909) );
  AND2_X1 U9574 ( .A1(n36604), .A2(n36428), .ZN(n36614) );
  NOR2_X1 U9575 ( .A1(n5990), .A2(n5989), .ZN(n5988) );
  NAND2_X1 U9576 ( .A1(n35310), .A2(n35305), .ZN(n5990) );
  OR2_X1 U9577 ( .A1(n39224), .A2(n3874), .ZN(n3873) );
  INV_X1 U9578 ( .A(n41004), .ZN(n5911) );
  OAI21_X1 U9579 ( .B1(n3707), .B2(n3706), .A(n38660), .ZN(n4887) );
  INV_X1 U9580 ( .A(n38994), .ZN(n38991) );
  OAI21_X1 U9581 ( .B1(n612), .B2(n37892), .A(n39401), .ZN(n3813) );
  INV_X1 U9582 ( .A(n38666), .ZN(n37210) );
  OR2_X1 U9583 ( .A1(n37665), .A2(n37667), .ZN(n4761) );
  AND2_X1 U9584 ( .A1(n51146), .A2(n43327), .ZN(n37605) );
  AND2_X1 U9585 ( .A1(n3985), .A2(n39390), .ZN(n7389) );
  NAND4_X1 U9586 ( .A1(n37769), .A2(n37771), .A3(n37772), .A4(n37770), .ZN(
        n37815) );
  OR2_X1 U9587 ( .A1(n37763), .A2(n37500), .ZN(n37770) );
  AND2_X1 U9588 ( .A1(n39429), .A2(n39423), .ZN(n39202) );
  OR2_X1 U9589 ( .A1(n38949), .A2(n38940), .ZN(n8186) );
  AND2_X1 U9590 ( .A1(n39009), .A2(n8478), .ZN(n8479) );
  INV_X1 U9591 ( .A(n38015), .ZN(n37996) );
  AND3_X1 U9592 ( .A1(n8644), .A2(n41268), .A3(n36786), .ZN(n4332) );
  AND2_X1 U9594 ( .A1(n38578), .A2(n38577), .ZN(n6820) );
  AND2_X1 U9595 ( .A1(n7977), .A2(n39834), .ZN(n40381) );
  INV_X1 U9596 ( .A(n37751), .ZN(n37510) );
  INV_X1 U9598 ( .A(n41113), .ZN(n41263) );
  INV_X1 U9599 ( .A(n40316), .ZN(n3043) );
  INV_X1 U9600 ( .A(n40806), .ZN(n39609) );
  AND2_X1 U9602 ( .A1(n38996), .A2(n38997), .ZN(n7406) );
  AND2_X1 U9603 ( .A1(n39938), .A2(n39955), .ZN(n7979) );
  OAI21_X1 U9604 ( .B1(n39236), .B2(n38302), .A(n39247), .ZN(n38305) );
  INV_X1 U9605 ( .A(n37802), .ZN(n39487) );
  NAND4_X2 U9606 ( .A1(n35322), .A2(n35323), .A3(n35321), .A4(n35324), .ZN(
        n39097) );
  NOR2_X1 U9607 ( .A1(n37892), .A2(n38998), .ZN(n39004) );
  INV_X1 U9608 ( .A(n38311), .ZN(n35853) );
  OR2_X1 U9609 ( .A1(n36542), .A2(n36540), .ZN(n36028) );
  AND2_X1 U9610 ( .A1(n3094), .A2(n40120), .ZN(n40124) );
  INV_X1 U9611 ( .A(n37639), .ZN(n5722) );
  OR2_X1 U9613 ( .A1(n38665), .A2(n38666), .ZN(n8134) );
  NOR2_X1 U9614 ( .A1(n4469), .A2(n38693), .ZN(n38694) );
  INV_X1 U9615 ( .A(n41200), .ZN(n40022) );
  AND2_X1 U9616 ( .A1(n5919), .A2(n41202), .ZN(n40668) );
  AOI22_X1 U9617 ( .A1(n38036), .A2(n2660), .B1(n35154), .B2(n38034), .ZN(
        n38047) );
  OAI21_X1 U9618 ( .B1(n40334), .B2(n40335), .A(n40336), .ZN(n40346) );
  OR2_X1 U9619 ( .A1(n36617), .A2(n36064), .ZN(n3838) );
  OR2_X1 U9620 ( .A1(n34925), .A2(n36062), .ZN(n3837) );
  AND3_X1 U9621 ( .A1(n34977), .A2(n34979), .A3(n38181), .ZN(n5873) );
  NOR2_X1 U9622 ( .A1(n37981), .A2(n594), .ZN(n5710) );
  NOR2_X1 U9623 ( .A1(n41195), .A2(n7955), .ZN(n41200) );
  INV_X1 U9624 ( .A(n41207), .ZN(n7955) );
  NOR2_X1 U9625 ( .A1(n51233), .A2(n40113), .ZN(n40122) );
  INV_X1 U9626 ( .A(n39551), .ZN(n40127) );
  OR2_X1 U9627 ( .A1(n40412), .A2(n5324), .ZN(n39734) );
  NOR2_X1 U9628 ( .A1(n685), .A2(n51052), .ZN(n5919) );
  INV_X1 U9629 ( .A(n40556), .ZN(n4302) );
  INV_X1 U9630 ( .A(n40565), .ZN(n40567) );
  AND2_X1 U9632 ( .A1(n35029), .A2(n7072), .ZN(n7071) );
  NOR2_X1 U9633 ( .A1(n41143), .A2(n40377), .ZN(n41146) );
  OR2_X1 U9635 ( .A1(n40782), .A2(n431), .ZN(n4777) );
  OR2_X1 U9636 ( .A1(n39800), .A2(n7015), .ZN(n40789) );
  AND2_X1 U9637 ( .A1(n39754), .A2(n39751), .ZN(n4251) );
  NAND4_X1 U9638 ( .A1(n41008), .A2(n43329), .A3(n39576), .A4(n38760), .ZN(
        n38761) );
  INV_X1 U9640 ( .A(n40801), .ZN(n7000) );
  OR2_X1 U9641 ( .A1(n42209), .A2(n2738), .ZN(n6980) );
  INV_X1 U9642 ( .A(n41617), .ZN(n41707) );
  AOI22_X1 U9643 ( .A1(n7660), .A2(n38549), .B1(n38551), .B2(n38550), .ZN(
        n8285) );
  AND2_X1 U9644 ( .A1(n38600), .A2(n38599), .ZN(n3230) );
  OAI22_X1 U9645 ( .A1(n34319), .A2(n40340), .B1(n52101), .B2(n40328), .ZN(
        n34324) );
  NOR2_X1 U9646 ( .A1(n36257), .A2(n34807), .ZN(n36254) );
  AND2_X1 U9647 ( .A1(n6961), .A2(n39103), .ZN(n40016) );
  AND2_X1 U9648 ( .A1(n39097), .A2(n6740), .ZN(n40011) );
  AND3_X1 U9649 ( .A1(n35946), .A2(n33465), .A3(n8719), .ZN(n6876) );
  NAND4_X2 U9650 ( .A1(n33565), .A2(n38510), .A3(n33563), .A4(n33564), .ZN(
        n41792) );
  AND2_X1 U9651 ( .A1(n6050), .A2(n33559), .ZN(n33565) );
  OR2_X1 U9652 ( .A1(n3647), .A2(n36241), .ZN(n36246) );
  NAND4_X2 U9653 ( .A1(n7513), .A2(n38069), .A3(n38070), .A4(n7514), .ZN(
        n40910) );
  AND2_X1 U9654 ( .A1(n7515), .A2(n38051), .ZN(n7514) );
  OR2_X1 U9655 ( .A1(n6940), .A2(n41104), .ZN(n41644) );
  NOR2_X1 U9656 ( .A1(n41096), .A2(n41642), .ZN(n41971) );
  INV_X1 U9657 ( .A(n39604), .ZN(n41052) );
  INV_X1 U9658 ( .A(n8317), .ZN(n39700) );
  AOI21_X1 U9660 ( .B1(n39394), .B2(n5050), .A(n5051), .ZN(n5049) );
  AND2_X1 U9661 ( .A1(n39393), .A2(n3737), .ZN(n5050) );
  NOR2_X1 U9662 ( .A1(n39396), .A2(n3737), .ZN(n5051) );
  INV_X1 U9664 ( .A(n41581), .ZN(n6236) );
  AND3_X1 U9666 ( .A1(n37723), .A2(n7373), .A3(n37724), .ZN(n7372) );
  NOR2_X1 U9667 ( .A1(n37815), .A2(n41770), .ZN(n42132) );
  OAI21_X1 U9668 ( .B1(n2433), .B2(n37720), .A(n3040), .ZN(n8494) );
  OR2_X1 U9669 ( .A1(n36257), .A2(n3041), .ZN(n3040) );
  INV_X1 U9670 ( .A(n40293), .ZN(n42050) );
  NOR2_X1 U9671 ( .A1(n41706), .A2(n41691), .ZN(n39873) );
  AND2_X1 U9672 ( .A1(n5475), .A2(n41690), .ZN(n41615) );
  INV_X1 U9673 ( .A(n41706), .ZN(n41703) );
  INV_X1 U9674 ( .A(n40647), .ZN(n40646) );
  NOR2_X1 U9678 ( .A1(n38414), .A2(n39927), .ZN(n5399) );
  AND2_X1 U9679 ( .A1(n35218), .A2(n35219), .ZN(n8376) );
  OR2_X1 U9680 ( .A1(n39889), .A2(n6469), .ZN(n5416) );
  NOR2_X1 U9681 ( .A1(n41692), .A2(n41690), .ZN(n40353) );
  OR2_X1 U9682 ( .A1(n40623), .A2(n41645), .ZN(n7638) );
  NAND4_X1 U9683 ( .A1(n40880), .A2(n40879), .A3(n40878), .A4(n40877), .ZN(
        n41308) );
  AND2_X1 U9684 ( .A1(n39873), .A2(n40353), .ZN(n41174) );
  AND2_X1 U9685 ( .A1(n4954), .A2(n40565), .ZN(n40559) );
  NAND4_X1 U9686 ( .A1(n4338), .A2(n4337), .A3(n38719), .A4(n3355), .ZN(n4626)
         );
  OAI21_X1 U9687 ( .B1(n39755), .B2(n39957), .A(n7979), .ZN(n6272) );
  INV_X1 U9690 ( .A(n41352), .ZN(n41360) );
  OAI211_X1 U9691 ( .C1(n39519), .C2(n39518), .A(n39517), .B(n39516), .ZN(
        n41968) );
  AND2_X1 U9692 ( .A1(n37960), .A2(n3624), .ZN(n37972) );
  NOR2_X1 U9693 ( .A1(n40910), .A2(n3655), .ZN(n40273) );
  NAND2_X1 U9694 ( .A1(n38511), .A2(n41319), .ZN(n3597) );
  OR2_X1 U9695 ( .A1(n41144), .A2(n41143), .ZN(n2638) );
  NOR2_X1 U9696 ( .A1(n51012), .A2(n41150), .ZN(n6550) );
  INV_X1 U9697 ( .A(n6345), .ZN(n42278) );
  INV_X1 U9698 ( .A(n42458), .ZN(n45357) );
  AND2_X1 U9700 ( .A1(n39859), .A2(n39860), .ZN(n8030) );
  INV_X1 U9701 ( .A(n43325), .ZN(n39611) );
  NOR2_X1 U9702 ( .A1(n6137), .A2(n51430), .ZN(n6136) );
  NAND2_X1 U9703 ( .A1(n41207), .A2(n40029), .ZN(n6137) );
  INV_X1 U9705 ( .A(n34668), .ZN(n7685) );
  NAND4_X1 U9706 ( .A1(n40466), .A2(n40465), .A3(n40463), .A4(n40464), .ZN(
        n42380) );
  AND2_X1 U9707 ( .A1(n36512), .A2(n36513), .ZN(n4574) );
  OR2_X1 U9708 ( .A1(n39752), .A2(n39943), .ZN(n39760) );
  AND2_X1 U9709 ( .A1(n4251), .A2(n2386), .ZN(n8070) );
  OAI21_X1 U9710 ( .B1(n41669), .B2(n8756), .A(n2771), .ZN(n2770) );
  OR2_X1 U9712 ( .A1(n41043), .A2(n5016), .ZN(n5012) );
  AND2_X1 U9713 ( .A1(n38886), .A2(n2789), .ZN(n38905) );
  INV_X1 U9714 ( .A(n37890), .ZN(n6088) );
  AOI22_X1 U9715 ( .A1(n6033), .A2(n34665), .B1(n34666), .B2(n6032), .ZN(n8110) );
  AND2_X1 U9716 ( .A1(n38810), .A2(n41792), .ZN(n41804) );
  INV_X1 U9718 ( .A(n7174), .ZN(n7173) );
  AND2_X1 U9719 ( .A1(n40207), .A2(n40208), .ZN(n5899) );
  INV_X1 U9720 ( .A(n8391), .ZN(n3862) );
  AOI21_X1 U9721 ( .B1(n41248), .B2(n41679), .A(n3860), .ZN(n3859) );
  OAI21_X1 U9722 ( .B1(n4894), .B2(n3858), .A(n8392), .ZN(n3857) );
  AND2_X1 U9723 ( .A1(n7029), .A2(n7031), .ZN(n5578) );
  INV_X1 U9725 ( .A(n45339), .ZN(n43344) );
  XNOR2_X1 U9726 ( .A(n42962), .B(n5353), .ZN(n41387) );
  INV_X1 U9727 ( .A(n43609), .ZN(n5353) );
  XNOR2_X1 U9728 ( .A(n41851), .B(n7102), .ZN(n42218) );
  AND2_X1 U9729 ( .A1(n48519), .A2(n46478), .ZN(n8685) );
  AND2_X1 U9730 ( .A1(n51451), .A2(n45562), .ZN(n8686) );
  INV_X1 U9731 ( .A(n49137), .ZN(n46287) );
  AND2_X1 U9732 ( .A1(n46280), .A2(n46292), .ZN(n3361) );
  INV_X1 U9733 ( .A(n46290), .ZN(n43427) );
  INV_X1 U9734 ( .A(n50378), .ZN(n49739) );
  AND2_X1 U9735 ( .A1(n50352), .A2(n47271), .ZN(n47275) );
  INV_X1 U9736 ( .A(n505), .ZN(n47278) );
  NOR2_X1 U9737 ( .A1(n2104), .A2(n46721), .ZN(n47094) );
  AND2_X1 U9738 ( .A1(n2159), .A2(n46565), .ZN(n7495) );
  OR2_X1 U9739 ( .A1(n46700), .A2(n46586), .ZN(n7680) );
  AND2_X1 U9740 ( .A1(n46583), .A2(n46584), .ZN(n7679) );
  NOR2_X1 U9741 ( .A1(n5170), .A2(n45780), .ZN(n45781) );
  AND2_X1 U9743 ( .A1(n44989), .A2(n46908), .ZN(n7700) );
  OR2_X1 U9744 ( .A1(n5562), .A2(n48437), .ZN(n44659) );
  INV_X1 U9745 ( .A(n48391), .ZN(n6986) );
  AND2_X1 U9746 ( .A1(n6194), .A2(n48165), .ZN(n48408) );
  OR2_X1 U9747 ( .A1(n46267), .A2(n45237), .ZN(n42602) );
  OR2_X1 U9748 ( .A1(n49205), .A2(n42702), .ZN(n4404) );
  OR2_X1 U9749 ( .A1(n8137), .A2(n49165), .ZN(n46248) );
  AND2_X1 U9750 ( .A1(n49170), .A2(n46255), .ZN(n8137) );
  AND2_X1 U9751 ( .A1(n46486), .A2(n4480), .ZN(n4698) );
  OR2_X1 U9752 ( .A1(n46505), .A2(n46380), .ZN(n4480) );
  AND2_X1 U9753 ( .A1(n49197), .A2(n45966), .ZN(n3842) );
  AND2_X1 U9755 ( .A1(n46282), .A2(n4460), .ZN(n45941) );
  OR2_X1 U9756 ( .A1(n49150), .A2(n49139), .ZN(n46286) );
  OAI21_X1 U9757 ( .B1(n45959), .B2(n50027), .A(n49671), .ZN(n45960) );
  AND3_X1 U9758 ( .A1(n43470), .A2(n42994), .A3(n42992), .ZN(n7796) );
  OR2_X1 U9759 ( .A1(n49663), .A2(n49667), .ZN(n50019) );
  INV_X1 U9760 ( .A(n47294), .ZN(n44608) );
  NAND2_X1 U9762 ( .A1(n50335), .A2(n505), .ZN(n50351) );
  INV_X1 U9763 ( .A(n44607), .ZN(n6669) );
  INV_X1 U9764 ( .A(n50339), .ZN(n47288) );
  INV_X1 U9765 ( .A(n47108), .ZN(n46570) );
  NOR2_X1 U9766 ( .A1(n2576), .A2(n47088), .ZN(n2575) );
  OR2_X1 U9767 ( .A1(n46568), .A2(n46878), .ZN(n46567) );
  INV_X1 U9768 ( .A(n47089), .ZN(n46878) );
  INV_X1 U9769 ( .A(n46830), .ZN(n47076) );
  AND2_X1 U9770 ( .A1(n46918), .A2(n46919), .ZN(n46922) );
  OR2_X1 U9772 ( .A1(n48701), .A2(n47410), .ZN(n48684) );
  INV_X1 U9774 ( .A(n47563), .ZN(n47574) );
  INV_X1 U9775 ( .A(n51289), .ZN(n47572) );
  AND2_X1 U9776 ( .A1(n45770), .A2(n45768), .ZN(n8158) );
  AND2_X1 U9777 ( .A1(n45796), .A2(n45797), .ZN(n4227) );
  NAND4_X1 U9778 ( .A1(n44863), .A2(n44862), .A3(n44861), .A4(n44860), .ZN(
        n45872) );
  AND3_X1 U9779 ( .A1(n45001), .A2(n45000), .A3(n44999), .ZN(n45005) );
  OAI21_X1 U9780 ( .B1(n45766), .B2(n44871), .A(n52153), .ZN(n6889) );
  INV_X1 U9781 ( .A(n47786), .ZN(n47762) );
  NOR2_X1 U9783 ( .A1(n47945), .A2(n47936), .ZN(n47981) );
  AOI21_X1 U9784 ( .B1(n44422), .B2(n44866), .A(n6756), .ZN(n6755) );
  INV_X1 U9785 ( .A(n45757), .ZN(n8646) );
  OR2_X1 U9786 ( .A1(n48077), .A2(n51092), .ZN(n48082) );
  AND2_X1 U9787 ( .A1(n8689), .A2(n48159), .ZN(n8065) );
  AND2_X1 U9788 ( .A1(n48103), .A2(n46535), .ZN(n8067) );
  NOR2_X1 U9789 ( .A1(n45611), .A2(n8689), .ZN(n48158) );
  NOR2_X1 U9790 ( .A1(n5502), .A2(n46542), .ZN(n48110) );
  NOR2_X1 U9791 ( .A1(n48156), .A2(n48159), .ZN(n48095) );
  INV_X1 U9792 ( .A(n48531), .ZN(n48547) );
  INV_X1 U9795 ( .A(n48540), .ZN(n46462) );
  OAI22_X1 U9796 ( .A1(n657), .A2(n46350), .B1(n46342), .B2(n46355), .ZN(
        n46366) );
  NOR2_X1 U9798 ( .A1(n46277), .A2(n46357), .ZN(n46350) );
  AND2_X1 U9799 ( .A1(n3247), .A2(n2266), .ZN(n6532) );
  INV_X1 U9800 ( .A(n48831), .ZN(n48796) );
  AND2_X1 U9801 ( .A1(n3247), .A2(n45213), .ZN(n3246) );
  OR2_X1 U9802 ( .A1(n46502), .A2(n46484), .ZN(n2687) );
  OR2_X1 U9803 ( .A1(n48912), .A2(n3782), .ZN(n5079) );
  NOR2_X1 U9804 ( .A1(n48908), .A2(n48912), .ZN(n48875) );
  INV_X1 U9805 ( .A(n48935), .ZN(n48958) );
  INV_X1 U9806 ( .A(n49020), .ZN(n49007) );
  NOR2_X1 U9807 ( .A1(n46265), .A2(n46264), .ZN(n2826) );
  INV_X1 U9808 ( .A(n49047), .ZN(n6391) );
  INV_X1 U9809 ( .A(n45216), .ZN(n45214) );
  AND2_X1 U9810 ( .A1(n44781), .A2(n44780), .ZN(n7213) );
  NOR2_X1 U9811 ( .A1(n44777), .A2(n7211), .ZN(n7210) );
  INV_X1 U9812 ( .A(n51729), .ZN(n49371) );
  INV_X1 U9813 ( .A(n2859), .ZN(n2858) );
  OR2_X1 U9814 ( .A1(n45993), .A2(n45997), .ZN(n7309) );
  OR2_X1 U9815 ( .A1(n6705), .A2(n6704), .ZN(n7310) );
  AOI21_X1 U9816 ( .B1(n45908), .B2(n52052), .A(n6160), .ZN(n6705) );
  AND2_X1 U9817 ( .A1(n52107), .A2(n49457), .ZN(n49393) );
  INV_X1 U9818 ( .A(n42905), .ZN(n5814) );
  AND2_X1 U9819 ( .A1(n43285), .A2(n3833), .ZN(n3832) );
  INV_X1 U9820 ( .A(n46032), .ZN(n5761) );
  AND2_X1 U9821 ( .A1(n50020), .A2(n5763), .ZN(n5762) );
  NOR2_X1 U9822 ( .A1(n51691), .A2(n7568), .ZN(n7567) );
  INV_X1 U9823 ( .A(n49638), .ZN(n7568) );
  INV_X1 U9824 ( .A(n50144), .ZN(n4203) );
  OR2_X1 U9825 ( .A1(n50145), .A2(n51645), .ZN(n50083) );
  INV_X1 U9826 ( .A(n50115), .ZN(n50101) );
  AND2_X1 U9827 ( .A1(n8508), .A2(n562), .ZN(n50098) );
  NOR2_X1 U9828 ( .A1(n50324), .A2(n1812), .ZN(n6416) );
  AND3_X1 U9830 ( .A1(n47347), .A2(n47346), .A3(n47348), .ZN(n2886) );
  INV_X1 U9831 ( .A(n50192), .ZN(n50226) );
  AOI21_X1 U9832 ( .B1(n52224), .B2(n47375), .A(n47374), .ZN(n47376) );
  NOR2_X1 U9833 ( .A1(n50482), .A2(n7114), .ZN(n50455) );
  OR2_X1 U9834 ( .A1(n49956), .A2(n50287), .ZN(n7141) );
  AND2_X1 U9835 ( .A1(n50638), .A2(n50598), .ZN(n50631) );
  INV_X1 U9836 ( .A(n50689), .ZN(n50692) );
  AND2_X1 U9837 ( .A1(n47068), .A2(n47063), .ZN(n6575) );
  AND3_X1 U9838 ( .A1(n47060), .A2(n47062), .A3(n47061), .ZN(n6574) );
  INV_X1 U9839 ( .A(n50772), .ZN(n50787) );
  OAI21_X1 U9840 ( .B1(n47146), .B2(n47145), .A(n47144), .ZN(n8668) );
  AND2_X1 U9841 ( .A1(n52093), .A2(n50886), .ZN(n50851) );
  AND2_X1 U9842 ( .A1(n50929), .A2(n50958), .ZN(n7323) );
  NOR2_X1 U9844 ( .A1(n46852), .A2(n3891), .ZN(n3890) );
  OR2_X1 U9845 ( .A1(n46845), .A2(n3892), .ZN(n3891) );
  NOR2_X1 U9846 ( .A1(n42396), .A2(n2267), .ZN(n6029) );
  INV_X1 U9847 ( .A(n42397), .ZN(n6028) );
  OR2_X1 U9848 ( .A1(n47570), .A2(n52045), .ZN(n47543) );
  AND3_X1 U9849 ( .A1(n46791), .A2(n46792), .A3(n6231), .ZN(n6230) );
  NOR2_X1 U9850 ( .A1(n47518), .A2(n47500), .ZN(n5992) );
  NOR2_X1 U9851 ( .A1(n47527), .A2(n47543), .ZN(n47521) );
  INV_X1 U9852 ( .A(n47539), .ZN(n47499) );
  NOR2_X1 U9853 ( .A1(n47557), .A2(n414), .ZN(n3019) );
  OR2_X1 U9854 ( .A1(n5573), .A2(n47591), .ZN(n47615) );
  AND3_X1 U9855 ( .A1(n47977), .A2(n47978), .A3(n6020), .ZN(n47999) );
  NAND4_X1 U9856 ( .A1(n646), .A2(n7766), .A3(n8061), .A4(n3911), .ZN(n3908)
         );
  AND2_X1 U9857 ( .A1(n48162), .A2(n48161), .ZN(n3909) );
  AND2_X2 U9858 ( .A1(n48186), .A2(n48187), .ZN(n8104) );
  INV_X1 U9859 ( .A(n48275), .ZN(n8259) );
  OR2_X1 U9860 ( .A1(n4946), .A2(n51728), .ZN(n48368) );
  OR2_X1 U9861 ( .A1(n48468), .A2(n48454), .ZN(n8379) );
  NOR2_X1 U9862 ( .A1(n4666), .A2(n655), .ZN(n7674) );
  AND2_X1 U9863 ( .A1(n7675), .A2(n4666), .ZN(n7673) );
  AND2_X1 U9864 ( .A1(n48880), .A2(n48886), .ZN(n5890) );
  AND2_X1 U9865 ( .A1(n49031), .A2(n49032), .ZN(n3792) );
  OAI21_X1 U9866 ( .B1(n49038), .B2(n49037), .A(n49039), .ZN(n3794) );
  AND4_X1 U9867 ( .A1(n5772), .A2(n49538), .A3(n49534), .A4(n49503), .ZN(n3897) );
  AND3_X1 U9868 ( .A1(n4983), .A2(n43488), .A3(n43489), .ZN(n4982) );
  OR2_X1 U9869 ( .A1(n49564), .A2(n6985), .ZN(n43416) );
  OR2_X1 U9870 ( .A1(n49682), .A2(n50029), .ZN(n6688) );
  INV_X1 U9871 ( .A(n49794), .ZN(n3944) );
  AND2_X1 U9872 ( .A1(n544), .A2(n50452), .ZN(n50466) );
  AND2_X1 U9873 ( .A1(n50440), .A2(n50439), .ZN(n2925) );
  NOR2_X1 U9875 ( .A1(n50563), .A2(n50508), .ZN(n5263) );
  AND2_X1 U9877 ( .A1(n50493), .A2(n50494), .ZN(n7473) );
  OAI21_X1 U9878 ( .B1(n6606), .B2(n50619), .A(n52061), .ZN(n50589) );
  NOR2_X1 U9879 ( .A1(n8018), .A2(n50599), .ZN(n6606) );
  OR2_X1 U9880 ( .A1(n50641), .A2(n44121), .ZN(n8616) );
  NOR2_X1 U9881 ( .A1(n50615), .A2(n52225), .ZN(n50619) );
  AND2_X1 U9882 ( .A1(n50625), .A2(n5838), .ZN(n5837) );
  NAND2_X1 U9883 ( .A1(n50613), .A2(n50614), .ZN(n5838) );
  NOR2_X1 U9884 ( .A1(n11467), .A2(n3024), .ZN(n3023) );
  OR2_X1 U9885 ( .A1(n7341), .A2(n11186), .ZN(n11568) );
  INV_X1 U9886 ( .A(n10037), .ZN(n6049) );
  AND2_X1 U9887 ( .A1(n10546), .A2(n10551), .ZN(n4077) );
  OAI21_X1 U9888 ( .B1(n11004), .B2(n876), .A(n7942), .ZN(n10255) );
  NOR2_X1 U9889 ( .A1(n10687), .A2(n6786), .ZN(n3611) );
  AND2_X1 U9890 ( .A1(n3079), .A2(n11662), .ZN(n9317) );
  BUF_X1 U9891 ( .A(n9178), .Z(n12660) );
  NOR2_X1 U9892 ( .A1(n12705), .A2(n11932), .ZN(n7781) );
  OR2_X1 U9893 ( .A1(n10279), .A2(n12328), .ZN(n10281) );
  OR2_X1 U9894 ( .A1(n11488), .A2(n11900), .ZN(n11063) );
  INV_X1 U9895 ( .A(n11908), .ZN(n11071) );
  XNOR2_X1 U9896 ( .A(Key[150]), .B(Ciphertext[119]), .ZN(n9459) );
  AND2_X1 U9897 ( .A1(n12573), .A2(n51760), .ZN(n2927) );
  AND2_X1 U9898 ( .A1(n2197), .A2(n10004), .ZN(n8407) );
  INV_X1 U9899 ( .A(n8885), .ZN(n5473) );
  INV_X1 U9900 ( .A(n11581), .ZN(n7340) );
  INV_X1 U9901 ( .A(n11569), .ZN(n11525) );
  OR2_X1 U9902 ( .A1(n12556), .A2(n11186), .ZN(n11510) );
  OR2_X1 U9903 ( .A1(n12256), .A2(n12255), .ZN(n4858) );
  OR2_X1 U9904 ( .A1(n11210), .A2(n643), .ZN(n11710) );
  NOR2_X1 U9905 ( .A1(n7993), .A2(n11621), .ZN(n7992) );
  OR2_X1 U9906 ( .A1(n9104), .A2(n9103), .ZN(n7993) );
  AND3_X1 U9907 ( .A1(n3250), .A2(n10816), .A3(n11590), .ZN(n3249) );
  INV_X1 U9909 ( .A(n9667), .ZN(n12337) );
  INV_X1 U9910 ( .A(n11032), .ZN(n10575) );
  INV_X1 U9911 ( .A(n11914), .ZN(n9538) );
  INV_X1 U9912 ( .A(n12496), .ZN(n8024) );
  OR2_X1 U9913 ( .A1(n8187), .A2(n13088), .ZN(n11161) );
  INV_X1 U9914 ( .A(n12914), .ZN(n8187) );
  AND2_X1 U9915 ( .A1(n9895), .A2(n11601), .ZN(n9280) );
  INV_X1 U9917 ( .A(n11269), .ZN(n11280) );
  INV_X1 U9919 ( .A(n5105), .ZN(n5107) );
  OR2_X1 U9920 ( .A1(n7019), .A2(n10662), .ZN(n11388) );
  NAND4_X1 U9921 ( .A1(n5687), .A2(n10356), .A3(n10362), .A4(n799), .ZN(n9389)
         );
  INV_X1 U9922 ( .A(n10664), .ZN(n3168) );
  AND2_X1 U9923 ( .A1(n10965), .A2(n10052), .ZN(n2865) );
  INV_X1 U9924 ( .A(n11600), .ZN(n11592) );
  AND2_X1 U9925 ( .A1(n8050), .A2(n12144), .ZN(n8049) );
  INV_X1 U9926 ( .A(n11276), .ZN(n4555) );
  INV_X1 U9927 ( .A(n9973), .ZN(n11274) );
  NOR2_X1 U9928 ( .A1(n11979), .A2(n797), .ZN(n10338) );
  INV_X1 U9929 ( .A(n10109), .ZN(n10026) );
  INV_X1 U9930 ( .A(n8818), .ZN(n10580) );
  NAND2_X1 U9931 ( .A1(n8639), .A2(n8818), .ZN(n11030) );
  INV_X1 U9933 ( .A(n12045), .ZN(n8349) );
  AOI22_X1 U9934 ( .A1(n10966), .A2(n10053), .B1(n10054), .B2(n10965), .ZN(
        n10059) );
  INV_X1 U9935 ( .A(n12532), .ZN(n6409) );
  INV_X1 U9936 ( .A(n12545), .ZN(n12537) );
  INV_X1 U9937 ( .A(n11402), .ZN(n10383) );
  INV_X1 U9938 ( .A(n14137), .ZN(n3564) );
  INV_X1 U9940 ( .A(n10124), .ZN(n3317) );
  INV_X1 U9941 ( .A(n10121), .ZN(n3316) );
  INV_X1 U9942 ( .A(n10956), .ZN(n10125) );
  NOR2_X1 U9943 ( .A1(n12481), .A2(n5252), .ZN(n5250) );
  AND2_X1 U9944 ( .A1(n10456), .A2(n12649), .ZN(n6423) );
  OR2_X1 U9945 ( .A1(n14410), .A2(n12961), .ZN(n14397) );
  INV_X1 U9946 ( .A(n11484), .ZN(n11065) );
  INV_X1 U9947 ( .A(n11941), .ZN(n11109) );
  AOI22_X1 U9948 ( .A1(n6445), .A2(n10976), .B1(n10986), .B2(n9023), .ZN(n6444) );
  AND2_X1 U9949 ( .A1(n9785), .A2(n10988), .ZN(n6445) );
  INV_X1 U9950 ( .A(n12341), .ZN(n12332) );
  AND2_X1 U9951 ( .A1(n9049), .A2(n3649), .ZN(n3648) );
  INV_X1 U9952 ( .A(n12478), .ZN(n12484) );
  INV_X1 U9953 ( .A(n10962), .ZN(n6004) );
  AND2_X1 U9954 ( .A1(n7340), .A2(n12555), .ZN(n12577) );
  INV_X1 U9955 ( .A(n12375), .ZN(n6712) );
  NAND2_X1 U9956 ( .A1(n2285), .A2(n12059), .ZN(n11395) );
  INV_X1 U9957 ( .A(n9515), .ZN(n11654) );
  OR2_X1 U9959 ( .A1(n7465), .A2(n14482), .ZN(n3289) );
  INV_X1 U9961 ( .A(n11268), .ZN(n10591) );
  INV_X1 U9962 ( .A(n14317), .ZN(n8227) );
  AND2_X1 U9964 ( .A1(n13854), .A2(n13841), .ZN(n7464) );
  OR2_X1 U9965 ( .A1(n12559), .A2(n5827), .ZN(n5826) );
  INV_X1 U9966 ( .A(n2828), .ZN(n11567) );
  NOR2_X1 U9967 ( .A1(n11191), .A2(n51760), .ZN(n11566) );
  AOI21_X1 U9969 ( .B1(n7236), .B2(n11920), .A(n4610), .ZN(n9545) );
  AND2_X1 U9970 ( .A1(n12589), .A2(n9543), .ZN(n4610) );
  OR2_X1 U9971 ( .A1(n12595), .A2(n9547), .ZN(n9548) );
  AND2_X1 U9972 ( .A1(n12384), .A2(n12373), .ZN(n12375) );
  OR2_X1 U9973 ( .A1(n12379), .A2(n12391), .ZN(n6479) );
  NAND2_X1 U9975 ( .A1(n9210), .A2(n12626), .ZN(n12617) );
  INV_X1 U9976 ( .A(n10633), .ZN(n6584) );
  OR2_X1 U9977 ( .A1(n10586), .A2(n11032), .ZN(n2911) );
  NOR2_X1 U9978 ( .A1(n10580), .A2(n11027), .ZN(n8458) );
  NOR2_X1 U9979 ( .A1(n15438), .A2(n15341), .ZN(n8140) );
  OR2_X1 U9980 ( .A1(n15421), .A2(n2640), .ZN(n13873) );
  NOR2_X1 U9981 ( .A1(n14342), .A2(n14339), .ZN(n14337) );
  OR2_X1 U9982 ( .A1(n11161), .A2(n13091), .ZN(n11820) );
  AND2_X1 U9983 ( .A1(n12755), .A2(n12756), .ZN(n14636) );
  AND3_X1 U9984 ( .A1(n10322), .A2(n10324), .A3(n10323), .ZN(n3459) );
  OR2_X1 U9985 ( .A1(n10563), .A2(n11639), .ZN(n4757) );
  AND2_X1 U9986 ( .A1(n11663), .A2(n11660), .ZN(n3883) );
  INV_X1 U9988 ( .A(n7865), .ZN(n12404) );
  AND2_X1 U9989 ( .A1(n13575), .A2(n13588), .ZN(n4209) );
  AND2_X1 U9990 ( .A1(n13560), .A2(n14472), .ZN(n3949) );
  INV_X1 U9991 ( .A(n14065), .ZN(n12868) );
  INV_X1 U9992 ( .A(n15286), .ZN(n14949) );
  OAI21_X1 U9993 ( .B1(n14660), .B2(n3563), .A(n12789), .ZN(n3562) );
  INV_X1 U9994 ( .A(n13990), .ZN(n3563) );
  INV_X1 U9995 ( .A(n4119), .ZN(n4118) );
  OAI21_X1 U9996 ( .B1(n10590), .B2(n11687), .A(n9341), .ZN(n4119) );
  OR2_X1 U9997 ( .A1(n14936), .A2(n15285), .ZN(n14063) );
  AND2_X1 U9998 ( .A1(n12834), .A2(n13633), .ZN(n7757) );
  INV_X1 U10000 ( .A(n15206), .ZN(n14763) );
  INV_X1 U10001 ( .A(n13299), .ZN(n12410) );
  INV_X1 U10002 ( .A(n13781), .ZN(n13776) );
  AND2_X1 U10004 ( .A1(n11660), .A2(n7185), .ZN(n3882) );
  INV_X1 U10005 ( .A(n12961), .ZN(n3512) );
  INV_X1 U10006 ( .A(n13939), .ZN(n4024) );
  AOI21_X1 U10007 ( .B1(n15135), .B2(n15134), .A(n13700), .ZN(n8386) );
  OAI21_X1 U10008 ( .B1(n14581), .B2(n15161), .A(n14580), .ZN(n5208) );
  AND2_X1 U10009 ( .A1(n14573), .A2(n14572), .ZN(n7714) );
  INV_X1 U10010 ( .A(n10766), .ZN(n13110) );
  OR2_X1 U10011 ( .A1(n12977), .A2(n14099), .ZN(n12848) );
  INV_X1 U10012 ( .A(n11048), .ZN(n12023) );
  NOR2_X1 U10013 ( .A1(n12252), .A2(n6067), .ZN(n8992) );
  AND3_X1 U10014 ( .A1(n8993), .A2(n8991), .A3(n12247), .ZN(n6213) );
  OR2_X1 U10016 ( .A1(n11014), .A2(n9743), .ZN(n3348) );
  AOI22_X1 U10017 ( .A1(n12671), .A2(n12672), .B1(n12674), .B2(n12673), .ZN(
        n12686) );
  INV_X1 U10019 ( .A(n12995), .ZN(n14597) );
  INV_X1 U10020 ( .A(n5175), .ZN(n5174) );
  OAI21_X1 U10021 ( .B1(n13169), .B2(n13179), .A(n13186), .ZN(n3628) );
  OR2_X1 U10022 ( .A1(n14710), .A2(n14200), .ZN(n14090) );
  INV_X1 U10024 ( .A(n13737), .ZN(n6726) );
  AND2_X1 U10025 ( .A1(n13575), .A2(n8397), .ZN(n12196) );
  OR2_X1 U10026 ( .A1(n13933), .A2(n13947), .ZN(n13202) );
  AND2_X1 U10027 ( .A1(n6668), .A2(n13930), .ZN(n13208) );
  NOR2_X1 U10028 ( .A1(n13207), .A2(n13948), .ZN(n13198) );
  NAND2_X1 U10029 ( .A1(n6299), .A2(n14178), .ZN(n6298) );
  AND2_X1 U10030 ( .A1(n3679), .A2(n13130), .ZN(n6296) );
  NOR2_X1 U10031 ( .A1(n14178), .A2(n12907), .ZN(n6295) );
  AND2_X1 U10032 ( .A1(n14178), .A2(n14186), .ZN(n10204) );
  INV_X1 U10034 ( .A(n14634), .ZN(n2763) );
  AND2_X1 U10035 ( .A1(n13412), .A2(n14344), .ZN(n13812) );
  OR2_X1 U10036 ( .A1(n14103), .A2(n14106), .ZN(n12976) );
  OR2_X1 U10037 ( .A1(n11433), .A2(n14453), .ZN(n12977) );
  OR2_X1 U10038 ( .A1(n784), .A2(n14285), .ZN(n12202) );
  AND2_X1 U10039 ( .A1(n15435), .A2(n8141), .ZN(n14860) );
  NOR2_X1 U10040 ( .A1(n14831), .A2(n15437), .ZN(n8141) );
  AND2_X1 U10041 ( .A1(n13124), .A2(n14164), .ZN(n5630) );
  OR2_X1 U10042 ( .A1(n15437), .A2(n15326), .ZN(n15439) );
  INV_X1 U10043 ( .A(n13529), .ZN(n13499) );
  NAND2_X1 U10044 ( .A1(n13533), .A2(n13532), .ZN(n4196) );
  OR2_X1 U10047 ( .A1(n14633), .A2(n13667), .ZN(n14632) );
  AND2_X1 U10048 ( .A1(n641), .A2(n13088), .ZN(n3350) );
  INV_X1 U10049 ( .A(n13040), .ZN(n12809) );
  OAI211_X1 U10050 ( .C1(n12378), .C2(n12090), .A(n4546), .B(n12089), .ZN(
        n12104) );
  OAI21_X1 U10051 ( .B1(n4601), .B2(n10373), .A(n10374), .ZN(n6054) );
  NOR2_X1 U10052 ( .A1(n3699), .A2(n3696), .ZN(n3695) );
  AND3_X1 U10053 ( .A1(n4707), .A2(n4708), .A3(n15416), .ZN(n13264) );
  OR2_X1 U10054 ( .A1(n13263), .A2(n13262), .ZN(n4708) );
  INV_X1 U10055 ( .A(n13036), .ZN(n14521) );
  AND2_X1 U10056 ( .A1(n7980), .A2(n7981), .ZN(n3987) );
  OR2_X1 U10057 ( .A1(n13075), .A2(n3834), .ZN(n7980) );
  INV_X1 U10058 ( .A(n13005), .ZN(n12007) );
  AOI21_X1 U10059 ( .B1(n13634), .B2(n13641), .A(n8350), .ZN(n12956) );
  AND2_X1 U10060 ( .A1(n9770), .A2(n9063), .ZN(n7561) );
  AND3_X1 U10061 ( .A1(n10979), .A2(n10980), .A3(n2454), .ZN(n4821) );
  INV_X1 U10062 ( .A(n14286), .ZN(n4424) );
  NOR2_X1 U10063 ( .A1(n14824), .A2(n14825), .ZN(n5258) );
  INV_X1 U10064 ( .A(n13526), .ZN(n13500) );
  INV_X1 U10065 ( .A(n11845), .ZN(n13515) );
  AND2_X1 U10067 ( .A1(n13091), .A2(n12914), .ZN(n4147) );
  AND2_X1 U10068 ( .A1(n14943), .A2(n14942), .ZN(n3084) );
  OR2_X1 U10070 ( .A1(n15259), .A2(n14784), .ZN(n15253) );
  INV_X1 U10071 ( .A(n13104), .ZN(n12917) );
  INV_X1 U10072 ( .A(n13587), .ZN(n14284) );
  INV_X1 U10073 ( .A(n14297), .ZN(n14295) );
  AND2_X1 U10074 ( .A1(n10907), .A2(n13774), .ZN(n13772) );
  OAI21_X1 U10075 ( .B1(n12994), .B2(n14003), .A(n14006), .ZN(n12999) );
  OAI21_X1 U10076 ( .B1(n12015), .B2(n12419), .A(n12014), .ZN(n12016) );
  XNOR2_X1 U10077 ( .A(n17133), .B(n3588), .ZN(n18150) );
  INV_X1 U10078 ( .A(n19196), .ZN(n3588) );
  OAI21_X1 U10079 ( .B1(n14172), .B2(n14171), .A(n5173), .ZN(n14173) );
  AND2_X1 U10080 ( .A1(n14663), .A2(n14664), .ZN(n5582) );
  OR2_X1 U10081 ( .A1(n13627), .A2(n7755), .ZN(n7754) );
  AND2_X1 U10082 ( .A1(n11314), .A2(n11319), .ZN(n5583) );
  OR4_X1 U10083 ( .A1(n13143), .A2(n14186), .A3(n13148), .A4(n14178), .ZN(
        n11176) );
  OAI21_X1 U10084 ( .B1(n11553), .B2(n11852), .A(n15385), .ZN(n11561) );
  AND2_X1 U10085 ( .A1(n15119), .A2(n352), .ZN(n2868) );
  AND3_X1 U10086 ( .A1(n13926), .A2(n13928), .A3(n13925), .ZN(n4819) );
  AOI21_X1 U10087 ( .B1(n13122), .B2(n14155), .A(n14156), .ZN(n2697) );
  OAI211_X1 U10088 ( .C1(n13574), .C2(n14298), .A(n5411), .B(n7135), .ZN(
        n11791) );
  INV_X1 U10089 ( .A(n13575), .ZN(n7135) );
  INV_X1 U10090 ( .A(n6794), .ZN(n11778) );
  AND2_X1 U10092 ( .A1(n13822), .A2(n13820), .ZN(n13605) );
  OR2_X1 U10094 ( .A1(n14914), .A2(n15063), .ZN(n3009) );
  INV_X1 U10095 ( .A(n12717), .ZN(n2589) );
  OAI21_X1 U10096 ( .B1(n2582), .B2(n2581), .A(n12700), .ZN(n2580) );
  INV_X1 U10097 ( .A(n13125), .ZN(n13759) );
  XNOR2_X1 U10098 ( .A(n3644), .B(n16701), .ZN(n15220) );
  INV_X1 U10099 ( .A(n9996), .ZN(n3644) );
  INV_X1 U10100 ( .A(n15294), .ZN(n19188) );
  AND3_X1 U10101 ( .A1(n14615), .A2(n14614), .A3(n14613), .ZN(n4652) );
  AND3_X1 U10102 ( .A1(n3016), .A2(n15328), .A3(n3015), .ZN(n15348) );
  NOR2_X1 U10103 ( .A1(n14997), .A2(n15126), .ZN(n5343) );
  INV_X1 U10104 ( .A(n21527), .ZN(n16859) );
  NOR2_X1 U10105 ( .A1(n16125), .A2(n21530), .ZN(n7420) );
  XNOR2_X1 U10106 ( .A(n4979), .B(n17257), .ZN(n17259) );
  INV_X1 U10108 ( .A(n14353), .ZN(n4310) );
  AND2_X1 U10109 ( .A1(n13008), .A2(n13425), .ZN(n4311) );
  AND2_X1 U10111 ( .A1(n14103), .A2(n14454), .ZN(n3263) );
  OAI211_X1 U10112 ( .C1(n14102), .C2(n14101), .A(n7887), .B(n7886), .ZN(n7885) );
  OAI211_X2 U10113 ( .C1(n12992), .C2(n10872), .A(n10880), .B(n8162), .ZN(
        n7191) );
  AND2_X1 U10114 ( .A1(n10879), .A2(n10878), .ZN(n8162) );
  OR2_X1 U10115 ( .A1(n13099), .A2(n8440), .ZN(n8439) );
  NOR2_X1 U10116 ( .A1(n13085), .A2(n3801), .ZN(n13109) );
  AND3_X1 U10117 ( .A1(n5765), .A2(n13456), .A3(n13460), .ZN(n5764) );
  XNOR2_X1 U10118 ( .A(n17145), .B(n15486), .ZN(n7643) );
  AOI22_X1 U10119 ( .A1(n13960), .A2(n13216), .B1(n9798), .B2(n13958), .ZN(
        n9802) );
  INV_X1 U10120 ( .A(n13701), .ZN(n5444) );
  NOR2_X1 U10121 ( .A1(n14268), .A2(n14269), .ZN(n2986) );
  INV_X1 U10123 ( .A(n14632), .ZN(n12754) );
  INV_X1 U10124 ( .A(n2827), .ZN(n7299) );
  OAI211_X1 U10126 ( .C1(n12880), .C2(n13206), .A(n11761), .B(n13192), .ZN(
        n4962) );
  INV_X1 U10127 ( .A(n13215), .ZN(n14226) );
  OR2_X1 U10128 ( .A1(n14234), .A2(n5540), .ZN(n14229) );
  NAND4_X1 U10129 ( .A1(n14222), .A2(n5825), .A3(n14233), .A4(n14223), .ZN(
        n14237) );
  AND2_X1 U10130 ( .A1(n12149), .A2(n12147), .ZN(n3674) );
  INV_X1 U10131 ( .A(n13881), .ZN(n15423) );
  NAND4_X1 U10132 ( .A1(n13341), .A2(n13342), .A3(n13340), .A4(n13339), .ZN(
        n14897) );
  AND2_X1 U10135 ( .A1(n14487), .A2(n14486), .ZN(n14496) );
  INV_X1 U10136 ( .A(n18888), .ZN(n3686) );
  NOR2_X1 U10137 ( .A1(n19793), .A2(n19792), .ZN(n7875) );
  INV_X1 U10138 ( .A(n20607), .ZN(n7160) );
  AND3_X1 U10139 ( .A1(n13156), .A2(n13155), .A3(n13154), .ZN(n13157) );
  NOR2_X1 U10140 ( .A1(n20474), .A2(n20478), .ZN(n18002) );
  XNOR2_X1 U10141 ( .A(n15220), .B(n3643), .ZN(n17648) );
  INV_X1 U10142 ( .A(n18643), .ZN(n3643) );
  INV_X1 U10143 ( .A(n16834), .ZN(n17440) );
  XNOR2_X1 U10144 ( .A(n15014), .B(n2314), .ZN(n18120) );
  AND2_X1 U10145 ( .A1(n4927), .A2(n10776), .ZN(n7194) );
  AND2_X1 U10146 ( .A1(n13375), .A2(n13374), .ZN(n13396) );
  XNOR2_X1 U10147 ( .A(n8237), .B(n16028), .ZN(n15604) );
  XNOR2_X1 U10148 ( .A(n15185), .B(n2311), .ZN(n8237) );
  OR2_X1 U10149 ( .A1(n19783), .A2(n19459), .ZN(n19127) );
  INV_X1 U10150 ( .A(n18352), .ZN(n7839) );
  AOI21_X1 U10151 ( .B1(n12921), .B2(n13244), .A(n4107), .ZN(n4106) );
  OR2_X1 U10153 ( .A1(n15237), .A2(n15236), .ZN(n14122) );
  AND2_X1 U10154 ( .A1(n14195), .A2(n14194), .ZN(n4929) );
  OAI21_X1 U10155 ( .B1(n6611), .B2(n6610), .A(n14185), .ZN(n4928) );
  NOR2_X1 U10156 ( .A1(n5715), .A2(n12033), .ZN(n12036) );
  INV_X1 U10157 ( .A(n21451), .ZN(n19362) );
  XNOR2_X1 U10158 ( .A(n6352), .B(n6351), .ZN(n16792) );
  INV_X1 U10159 ( .A(n16719), .ZN(n6352) );
  XNOR2_X1 U10160 ( .A(n16717), .B(n16718), .ZN(n6351) );
  OR2_X1 U10161 ( .A1(n20608), .A2(n21520), .ZN(n16867) );
  OR2_X1 U10162 ( .A1(n19521), .A2(n19520), .ZN(n4528) );
  INV_X1 U10163 ( .A(n20215), .ZN(n4681) );
  INV_X1 U10164 ( .A(n19774), .ZN(n5229) );
  NOR2_X1 U10165 ( .A1(n19459), .A2(n19461), .ZN(n3509) );
  INV_X1 U10166 ( .A(n18394), .ZN(n15642) );
  INV_X1 U10167 ( .A(n17999), .ZN(n20462) );
  INV_X1 U10168 ( .A(n16125), .ZN(n20614) );
  OR2_X1 U10169 ( .A1(n52213), .A2(n16125), .ZN(n20607) );
  AND3_X1 U10171 ( .A1(n14255), .A2(n14254), .A3(n14253), .ZN(n3382) );
  AND2_X1 U10172 ( .A1(n11061), .A2(n14787), .ZN(n4073) );
  INV_X1 U10173 ( .A(n16722), .ZN(n16321) );
  INV_X1 U10174 ( .A(n20628), .ZN(n21540) );
  OR2_X1 U10175 ( .A1(n16873), .A2(n20230), .ZN(n7951) );
  AND2_X1 U10176 ( .A1(n20672), .A2(n20231), .ZN(n8552) );
  AND2_X1 U10177 ( .A1(n17492), .A2(n2166), .ZN(n4467) );
  INV_X1 U10178 ( .A(n20474), .ZN(n20394) );
  NOR2_X1 U10180 ( .A1(n5953), .A2(n51711), .ZN(n21564) );
  OR2_X1 U10182 ( .A1(n18234), .A2(n18921), .ZN(n18239) );
  AND2_X1 U10183 ( .A1(n52213), .A2(n16125), .ZN(n18895) );
  NOR3_X1 U10184 ( .A1(n19800), .A2(n19793), .A3(n21300), .ZN(n7097) );
  AND2_X1 U10185 ( .A1(n21300), .A2(n18996), .ZN(n4521) );
  INV_X1 U10186 ( .A(n21231), .ZN(n8409) );
  OAI21_X1 U10187 ( .B1(n19110), .B2(n19109), .A(n19112), .ZN(n5626) );
  INV_X1 U10189 ( .A(n17057), .ZN(n20100) );
  OR2_X1 U10190 ( .A1(n20698), .A2(n21620), .ZN(n21622) );
  INV_X1 U10191 ( .A(n19681), .ZN(n20216) );
  INV_X1 U10192 ( .A(n21555), .ZN(n20601) );
  AND2_X1 U10193 ( .A1(n21584), .A2(n5192), .ZN(n21403) );
  INV_X1 U10194 ( .A(n21406), .ZN(n21583) );
  AOI21_X1 U10195 ( .B1(n21412), .B2(n18823), .A(n51710), .ZN(n21581) );
  XNOR2_X1 U10196 ( .A(n16753), .B(n2275), .ZN(n17059) );
  INV_X1 U10197 ( .A(n20097), .ZN(n6312) );
  NOR2_X1 U10198 ( .A1(n51128), .A2(n20207), .ZN(n7857) );
  AND2_X1 U10199 ( .A1(n4681), .A2(n19681), .ZN(n20218) );
  AND2_X1 U10200 ( .A1(n20225), .A2(n20214), .ZN(n4680) );
  INV_X1 U10201 ( .A(n18895), .ZN(n20609) );
  INV_X1 U10203 ( .A(n20478), .ZN(n3745) );
  XNOR2_X1 U10204 ( .A(n14051), .B(n2302), .ZN(n6989) );
  INV_X1 U10205 ( .A(n18070), .ZN(n18061) );
  OR2_X1 U10206 ( .A1(n7484), .A2(n20642), .ZN(n19933) );
  NAND2_X1 U10207 ( .A1(n3187), .A2(n7484), .ZN(n20737) );
  INV_X1 U10208 ( .A(n20638), .ZN(n3187) );
  NOR2_X1 U10209 ( .A1(n18997), .A2(n18999), .ZN(n8574) );
  AND2_X1 U10210 ( .A1(n18352), .A2(n19066), .ZN(n20136) );
  INV_X1 U10211 ( .A(n20044), .ZN(n20045) );
  INV_X1 U10212 ( .A(n20476), .ZN(n2560) );
  NOR2_X1 U10213 ( .A1(n3746), .A2(n17639), .ZN(n3747) );
  AND2_X1 U10214 ( .A1(n15093), .A2(n18288), .ZN(n17496) );
  INV_X1 U10215 ( .A(n23507), .ZN(n21902) );
  OR2_X1 U10216 ( .A1(n18011), .A2(n16846), .ZN(n8486) );
  AOI21_X1 U10217 ( .B1(n21538), .B2(n20749), .A(n6929), .ZN(n20750) );
  NOR2_X1 U10218 ( .A1(n3729), .A2(n25062), .ZN(n3728) );
  INV_X1 U10219 ( .A(n25055), .ZN(n3729) );
  INV_X1 U10220 ( .A(n19710), .ZN(n19708) );
  INV_X1 U10221 ( .A(n19636), .ZN(n5936) );
  AND2_X1 U10222 ( .A1(n51127), .A2(n5749), .ZN(n18246) );
  INV_X1 U10223 ( .A(n19892), .ZN(n5750) );
  XNOR2_X1 U10224 ( .A(n8501), .B(n15677), .ZN(n15867) );
  INV_X1 U10225 ( .A(n22624), .ZN(n23087) );
  NOR2_X1 U10226 ( .A1(n3371), .A2(n3370), .ZN(n3369) );
  OR2_X1 U10227 ( .A1(n760), .A2(n20230), .ZN(n8094) );
  NOR2_X1 U10228 ( .A1(n52174), .A2(n23101), .ZN(n7807) );
  INV_X1 U10229 ( .A(n20147), .ZN(n18362) );
  OR2_X1 U10230 ( .A1(n17412), .A2(n21234), .ZN(n19512) );
  INV_X1 U10231 ( .A(n18458), .ZN(n8623) );
  INV_X1 U10232 ( .A(n16792), .ZN(n20088) );
  NOR2_X1 U10233 ( .A1(n19047), .A2(n16490), .ZN(n17094) );
  AND2_X1 U10234 ( .A1(n7119), .A2(n21713), .ZN(n6260) );
  OR2_X1 U10235 ( .A1(n23244), .A2(n23257), .ZN(n22125) );
  AND2_X1 U10236 ( .A1(n23513), .A2(n52206), .ZN(n23507) );
  INV_X1 U10237 ( .A(n21283), .ZN(n6868) );
  INV_X1 U10238 ( .A(n22593), .ZN(n5041) );
  OAI21_X1 U10240 ( .B1(n5231), .B2(n21211), .A(n21195), .ZN(n5284) );
  INV_X1 U10241 ( .A(n23167), .ZN(n7811) );
  OAI211_X1 U10242 ( .C1(n17873), .C2(n5671), .A(n51374), .B(n19410), .ZN(
        n17874) );
  INV_X1 U10244 ( .A(n20434), .ZN(n19324) );
  AND2_X1 U10245 ( .A1(n20737), .A2(n20630), .ZN(n3188) );
  INV_X1 U10246 ( .A(n20630), .ZN(n20736) );
  INV_X1 U10247 ( .A(n18742), .ZN(n6671) );
  INV_X1 U10248 ( .A(n20029), .ZN(n6711) );
  NOR2_X1 U10249 ( .A1(n21543), .A2(n20197), .ZN(n20194) );
  OR2_X1 U10250 ( .A1(n17404), .A2(n21199), .ZN(n21204) );
  OR2_X1 U10251 ( .A1(n19472), .A2(n3885), .ZN(n17084) );
  AND2_X1 U10254 ( .A1(n23171), .A2(n23166), .ZN(n6462) );
  OR2_X1 U10255 ( .A1(n22983), .A2(n22977), .ZN(n22441) );
  AND2_X1 U10257 ( .A1(n18971), .A2(n18970), .ZN(n7189) );
  AND2_X1 U10258 ( .A1(n21133), .A2(n22466), .ZN(n6593) );
  OAI21_X1 U10259 ( .B1(n15630), .B2(n19893), .A(n19658), .ZN(n7258) );
  INV_X1 U10260 ( .A(n23341), .ZN(n21144) );
  INV_X1 U10261 ( .A(n22359), .ZN(n5542) );
  AND3_X1 U10262 ( .A1(n21526), .A2(n21527), .A3(n21528), .ZN(n6163) );
  OR2_X1 U10263 ( .A1(n21520), .A2(n21521), .ZN(n3345) );
  OR2_X1 U10264 ( .A1(n21245), .A2(n19477), .ZN(n2936) );
  OR2_X1 U10265 ( .A1(n19060), .A2(n20109), .ZN(n8266) );
  NOR2_X1 U10266 ( .A1(n3314), .A2(n6652), .ZN(n6650) );
  OR2_X1 U10267 ( .A1(n51200), .A2(n21756), .ZN(n23335) );
  OR2_X1 U10268 ( .A1(n22290), .A2(n21782), .ZN(n2884) );
  OR2_X1 U10269 ( .A1(n20795), .A2(n21389), .ZN(n4414) );
  INV_X1 U10270 ( .A(n18933), .ZN(n16881) );
  NOR2_X1 U10271 ( .A1(n7947), .A2(n19894), .ZN(n7946) );
  AND2_X1 U10272 ( .A1(n19894), .A2(n19892), .ZN(n8502) );
  AND2_X1 U10273 ( .A1(n7707), .A2(n24290), .ZN(n20984) );
  INV_X1 U10274 ( .A(n21318), .ZN(n22019) );
  INV_X1 U10275 ( .A(n23445), .ZN(n21319) );
  INV_X1 U10276 ( .A(n19131), .ZN(n19490) );
  INV_X1 U10277 ( .A(n19381), .ZN(n20480) );
  OR2_X1 U10278 ( .A1(n20471), .A2(n4098), .ZN(n14739) );
  AND2_X1 U10280 ( .A1(n17582), .A2(n8604), .ZN(n3638) );
  AND2_X1 U10281 ( .A1(n50992), .A2(n22140), .ZN(n21931) );
  AND2_X1 U10282 ( .A1(n22548), .A2(n5269), .ZN(n8215) );
  INV_X1 U10283 ( .A(n5610), .ZN(n23433) );
  INV_X1 U10284 ( .A(n20720), .ZN(n23363) );
  OR2_X1 U10285 ( .A1(n22687), .A2(n51033), .ZN(n23136) );
  INV_X1 U10286 ( .A(n23821), .ZN(n23826) );
  AND3_X1 U10287 ( .A1(n5559), .A2(n5557), .A3(n5560), .ZN(n6530) );
  OR2_X1 U10288 ( .A1(n5069), .A2(n23637), .ZN(n7617) );
  AND2_X1 U10289 ( .A1(n23086), .A2(n5068), .ZN(n5067) );
  AOI21_X1 U10290 ( .B1(n23087), .B2(n559), .A(n754), .ZN(n23089) );
  AND2_X1 U10291 ( .A1(n754), .A2(n23631), .ZN(n7820) );
  OAI21_X1 U10292 ( .B1(n18720), .B2(n18721), .A(n19290), .ZN(n8491) );
  OR2_X1 U10293 ( .A1(n20144), .A2(n7843), .ZN(n18349) );
  AND2_X1 U10294 ( .A1(n23209), .A2(n23230), .ZN(n18387) );
  OR2_X1 U10295 ( .A1(n23142), .A2(n23135), .ZN(n22687) );
  INV_X1 U10297 ( .A(n20084), .ZN(n23423) );
  NAND2_X1 U10298 ( .A1(n6261), .A2(n6260), .ZN(n6259) );
  AND2_X1 U10299 ( .A1(n21711), .A2(n21700), .ZN(n6261) );
  OR2_X1 U10302 ( .A1(n23986), .A2(n23981), .ZN(n5103) );
  OR2_X1 U10303 ( .A1(n6875), .A2(n23154), .ZN(n2894) );
  OR2_X1 U10304 ( .A1(n22110), .A2(n24026), .ZN(n7492) );
  OR2_X1 U10305 ( .A1(n23673), .A2(n24036), .ZN(n7491) );
  NOR2_X1 U10306 ( .A1(n23436), .A2(n22593), .ZN(n22018) );
  AND2_X1 U10307 ( .A1(n6930), .A2(n22586), .ZN(n19549) );
  OR2_X1 U10308 ( .A1(n22390), .A2(n50977), .ZN(n22733) );
  NOR2_X1 U10310 ( .A1(n21945), .A2(n21948), .ZN(n23465) );
  OR2_X1 U10311 ( .A1(n22145), .A2(n22151), .ZN(n19559) );
  AOI21_X1 U10313 ( .B1(n22986), .B2(n22562), .A(n22985), .ZN(n3690) );
  XNOR2_X1 U10314 ( .A(n28381), .B(n3031), .ZN(n28258) );
  AND2_X1 U10315 ( .A1(n24111), .A2(n5951), .ZN(n5950) );
  AND2_X1 U10316 ( .A1(n24413), .A2(n24411), .ZN(n5951) );
  AND2_X1 U10317 ( .A1(n23637), .A2(n23950), .ZN(n20847) );
  INV_X1 U10318 ( .A(n8353), .ZN(n22764) );
  OAI21_X1 U10319 ( .B1(n23835), .B2(n23833), .A(n630), .ZN(n4671) );
  NOR2_X1 U10320 ( .A1(n23821), .A2(n630), .ZN(n23268) );
  OAI22_X1 U10321 ( .A1(n22005), .A2(n22023), .B1(n23442), .B2(n23447), .ZN(
        n22006) );
  OR2_X1 U10322 ( .A1(n23832), .A2(n23825), .ZN(n2908) );
  INV_X1 U10323 ( .A(n23271), .ZN(n23831) );
  AND2_X1 U10324 ( .A1(n7076), .A2(n23823), .ZN(n23839) );
  NOR2_X1 U10325 ( .A1(n21067), .A2(n22832), .ZN(n22223) );
  OR2_X1 U10326 ( .A1(n22506), .A2(n20298), .ZN(n21067) );
  OAI211_X1 U10327 ( .C1(n23102), .C2(n23101), .A(n23100), .B(n6171), .ZN(
        n25061) );
  AND2_X1 U10328 ( .A1(n51654), .A2(n25064), .ZN(n6171) );
  INV_X1 U10330 ( .A(n24155), .ZN(n24145) );
  AND2_X1 U10331 ( .A1(n21780), .A2(n51081), .ZN(n20948) );
  OR2_X1 U10332 ( .A1(n20944), .A2(n22699), .ZN(n20946) );
  INV_X1 U10333 ( .A(n24106), .ZN(n23734) );
  OAI21_X1 U10334 ( .B1(n21715), .B2(n3872), .A(n19917), .ZN(n3871) );
  INV_X1 U10335 ( .A(n19916), .ZN(n3872) );
  NOR2_X1 U10336 ( .A1(n6655), .A2(n23261), .ZN(n8706) );
  NOR2_X1 U10337 ( .A1(n23259), .A2(n22654), .ZN(n6655) );
  OR2_X1 U10338 ( .A1(n22796), .A2(n4349), .ZN(n23915) );
  NOR2_X1 U10340 ( .A1(n21778), .A2(n22702), .ZN(n22704) );
  INV_X1 U10341 ( .A(n24284), .ZN(n4087) );
  INV_X1 U10342 ( .A(n21904), .ZN(n23504) );
  INV_X1 U10343 ( .A(n23345), .ZN(n3003) );
  INV_X1 U10344 ( .A(n23318), .ZN(n23319) );
  OAI21_X1 U10345 ( .B1(n22954), .B2(n22955), .A(n23317), .ZN(n23307) );
  OR2_X1 U10346 ( .A1(n21782), .A2(n24452), .ZN(n3017) );
  AND2_X1 U10347 ( .A1(n24001), .A2(n24000), .ZN(n22427) );
  INV_X1 U10348 ( .A(n23611), .ZN(n22644) );
  OR2_X1 U10349 ( .A1(n23698), .A2(n23697), .ZN(n3960) );
  OR2_X1 U10350 ( .A1(n21048), .A2(n23417), .ZN(n7648) );
  AND2_X1 U10351 ( .A1(n20081), .A2(n20080), .ZN(n3186) );
  OR2_X1 U10352 ( .A1(n24249), .A2(n21820), .ZN(n24251) );
  OAI21_X1 U10353 ( .B1(n23786), .B2(n23785), .A(n5296), .ZN(n24243) );
  INV_X1 U10354 ( .A(n23784), .ZN(n5296) );
  OR2_X1 U10355 ( .A1(n22703), .A2(n20948), .ZN(n22286) );
  INV_X1 U10356 ( .A(n22703), .ZN(n22698) );
  INV_X1 U10357 ( .A(n22260), .ZN(n7321) );
  NAND4_X1 U10360 ( .A1(n5007), .A2(n6631), .A3(n2832), .A4(n19402), .ZN(n2831) );
  INV_X1 U10361 ( .A(n19609), .ZN(n19611) );
  AND2_X1 U10363 ( .A1(n24029), .A2(n24026), .ZN(n23674) );
  AND3_X1 U10364 ( .A1(n5703), .A2(n23669), .A3(n23670), .ZN(n5702) );
  AND2_X1 U10365 ( .A1(n3192), .A2(n3191), .ZN(n3190) );
  INV_X1 U10366 ( .A(n21948), .ZN(n8416) );
  INV_X1 U10367 ( .A(n23156), .ZN(n7593) );
  INV_X1 U10368 ( .A(n22157), .ZN(n20952) );
  INV_X1 U10369 ( .A(n22034), .ZN(n23422) );
  AND2_X1 U10371 ( .A1(n6064), .A2(n20560), .ZN(n3929) );
  XNOR2_X1 U10372 ( .A(n51646), .B(n28038), .ZN(n25571) );
  XNOR2_X1 U10373 ( .A(n3110), .B(n3030), .ZN(n27201) );
  INV_X1 U10374 ( .A(n28048), .ZN(n3030) );
  INV_X1 U10375 ( .A(n24188), .ZN(n4328) );
  INV_X1 U10376 ( .A(n50977), .ZN(n22741) );
  AND3_X1 U10377 ( .A1(n4736), .A2(n19724), .A3(n4735), .ZN(n7347) );
  AOI22_X1 U10378 ( .A1(n3087), .A2(n3086), .B1(n21180), .B2(n19703), .ZN(
        n3085) );
  AND2_X1 U10379 ( .A1(n19742), .A2(n18909), .ZN(n5093) );
  INV_X1 U10380 ( .A(n6082), .ZN(n25673) );
  INV_X1 U10381 ( .A(n23912), .ZN(n23908) );
  NOR2_X1 U10382 ( .A1(n23141), .A2(n5143), .ZN(n8153) );
  INV_X1 U10383 ( .A(n2846), .ZN(n2795) );
  OR2_X1 U10384 ( .A1(n23023), .A2(n8370), .ZN(n8369) );
  XNOR2_X1 U10385 ( .A(n26304), .B(n25724), .ZN(n26552) );
  OR3_X2 U10386 ( .A1(n6513), .A2(n23355), .A3(n2273), .ZN(n28396) );
  XNOR2_X1 U10387 ( .A(n3031), .B(n25813), .ZN(n25691) );
  INV_X1 U10388 ( .A(n2667), .ZN(n26274) );
  INV_X1 U10390 ( .A(n23378), .ZN(n3815) );
  INV_X1 U10391 ( .A(n22586), .ZN(n23434) );
  INV_X1 U10392 ( .A(n22022), .ZN(n22021) );
  NOR2_X1 U10394 ( .A1(n22080), .A2(n23044), .ZN(n2913) );
  AOI22_X1 U10395 ( .A1(n22406), .A2(n22120), .B1(n20973), .B2(n23209), .ZN(
        n20978) );
  XNOR2_X1 U10396 ( .A(n7350), .B(n42918), .ZN(n24866) );
  AND3_X1 U10397 ( .A1(n22414), .A2(n22413), .A3(n6311), .ZN(n6309) );
  AOI21_X1 U10398 ( .B1(n20546), .B2(n22722), .A(n3776), .ZN(n20553) );
  INV_X1 U10399 ( .A(n25540), .ZN(n22747) );
  INV_X1 U10400 ( .A(n26523), .ZN(n7553) );
  OR2_X1 U10401 ( .A1(n22794), .A2(n22793), .ZN(n2621) );
  XNOR2_X1 U10402 ( .A(n25339), .B(n33429), .ZN(n4368) );
  XNOR2_X1 U10404 ( .A(n25540), .B(n26529), .ZN(n23941) );
  INV_X1 U10405 ( .A(n23941), .ZN(n27346) );
  XNOR2_X1 U10406 ( .A(n6159), .B(n6158), .ZN(n25317) );
  INV_X1 U10407 ( .A(n25125), .ZN(n6159) );
  INV_X1 U10408 ( .A(n25639), .ZN(n8281) );
  OR2_X1 U10409 ( .A1(n3120), .A2(n21867), .ZN(n3119) );
  OR2_X1 U10410 ( .A1(n22822), .A2(n320), .ZN(n22840) );
  XNOR2_X1 U10411 ( .A(n22973), .B(n2667), .ZN(n26575) );
  AND2_X1 U10412 ( .A1(n5134), .A2(n3748), .ZN(n5132) );
  MUX2_X1 U10413 ( .A(n21774), .B(n21773), .S(n21782), .Z(n21789) );
  AOI21_X1 U10414 ( .B1(n22267), .B2(n22642), .A(n2800), .ZN(n22271) );
  XNOR2_X1 U10415 ( .A(n24736), .B(n6601), .ZN(n24737) );
  XNOR2_X1 U10416 ( .A(n26531), .B(n26221), .ZN(n5613) );
  XNOR2_X1 U10417 ( .A(n28221), .B(n25493), .ZN(n26436) );
  INV_X1 U10418 ( .A(n28201), .ZN(n28927) );
  INV_X1 U10419 ( .A(n25915), .ZN(n25738) );
  XNOR2_X1 U10420 ( .A(n25804), .B(n25803), .ZN(n25840) );
  XNOR2_X1 U10421 ( .A(n7939), .B(n25173), .ZN(n25174) );
  INV_X1 U10422 ( .A(n25479), .ZN(n4965) );
  INV_X1 U10423 ( .A(n444), .ZN(n24911) );
  INV_X1 U10424 ( .A(n25259), .ZN(n7933) );
  INV_X1 U10425 ( .A(n27197), .ZN(n26573) );
  AOI22_X1 U10426 ( .A1(n23490), .A2(n8475), .B1(n21978), .B2(n8474), .ZN(
        n21994) );
  INV_X1 U10427 ( .A(n27303), .ZN(n26584) );
  INV_X1 U10429 ( .A(n24776), .ZN(n26743) );
  NOR2_X1 U10430 ( .A1(n27668), .A2(n2677), .ZN(n26742) );
  XNOR2_X1 U10431 ( .A(n28292), .B(n5726), .ZN(n26535) );
  OAI21_X1 U10432 ( .B1(n22718), .B2(n22308), .A(n2083), .ZN(n22310) );
  INV_X1 U10433 ( .A(n28194), .ZN(n28572) );
  XNOR2_X1 U10434 ( .A(n26272), .B(n26277), .ZN(n5678) );
  NOR2_X1 U10435 ( .A1(n30795), .A2(n51722), .ZN(n23660) );
  AND3_X1 U10436 ( .A1(n3760), .A2(n23545), .A3(n3758), .ZN(n6917) );
  INV_X1 U10437 ( .A(n22412), .ZN(n22410) );
  OAI21_X1 U10438 ( .B1(n21724), .B2(n3635), .A(n418), .ZN(n21729) );
  OR2_X1 U10439 ( .A1(n29485), .A2(n25841), .ZN(n29489) );
  INV_X1 U10440 ( .A(n30211), .ZN(n27876) );
  INV_X1 U10441 ( .A(n29428), .ZN(n26997) );
  XNOR2_X1 U10442 ( .A(n20886), .B(n20860), .ZN(n3470) );
  XNOR2_X1 U10443 ( .A(n27497), .B(n2288), .ZN(n28333) );
  INV_X1 U10445 ( .A(n28662), .ZN(n28657) );
  XNOR2_X1 U10446 ( .A(n7971), .B(n26565), .ZN(n25681) );
  INV_X1 U10447 ( .A(n28713), .ZN(n29271) );
  OR2_X1 U10448 ( .A1(n29184), .A2(n29185), .ZN(n29273) );
  INV_X1 U10449 ( .A(n29283), .ZN(n7370) );
  INV_X1 U10450 ( .A(n28291), .ZN(n5725) );
  XNOR2_X1 U10451 ( .A(n25503), .B(n25496), .ZN(n4366) );
  AND2_X1 U10452 ( .A1(n29259), .A2(n29252), .ZN(n28662) );
  INV_X1 U10453 ( .A(n28361), .ZN(n28357) );
  OR2_X1 U10454 ( .A1(n28948), .A2(n28965), .ZN(n7902) );
  INV_X1 U10455 ( .A(n29921), .ZN(n29915) );
  XNOR2_X1 U10456 ( .A(n24441), .B(n2320), .ZN(n26954) );
  XNOR2_X1 U10457 ( .A(n27502), .B(n6601), .ZN(n26401) );
  INV_X1 U10458 ( .A(n25935), .ZN(n8179) );
  INV_X1 U10459 ( .A(n23301), .ZN(n29900) );
  INV_X1 U10460 ( .A(n401), .ZN(n27525) );
  XNOR2_X1 U10461 ( .A(n25495), .B(n25493), .ZN(n8444) );
  OR2_X1 U10462 ( .A1(n28849), .A2(n29065), .ZN(n28779) );
  INV_X1 U10463 ( .A(n27993), .ZN(n28582) );
  INV_X1 U10464 ( .A(n28872), .ZN(n28877) );
  INV_X1 U10465 ( .A(n29006), .ZN(n28007) );
  XNOR2_X1 U10466 ( .A(n28311), .B(n5024), .ZN(n26397) );
  XNOR2_X1 U10467 ( .A(n23842), .B(n23841), .ZN(n25143) );
  INV_X1 U10468 ( .A(n26556), .ZN(n8322) );
  INV_X1 U10469 ( .A(n26175), .ZN(n5383) );
  XNOR2_X1 U10470 ( .A(n26436), .B(n28343), .ZN(n26596) );
  XNOR2_X1 U10471 ( .A(n26517), .B(n8627), .ZN(n26619) );
  NOR2_X1 U10472 ( .A1(n31547), .A2(n31546), .ZN(n4163) );
  INV_X1 U10473 ( .A(n29308), .ZN(n28684) );
  INV_X1 U10474 ( .A(n28695), .ZN(n28690) );
  INV_X1 U10475 ( .A(n26083), .ZN(n29294) );
  INV_X1 U10476 ( .A(n27847), .ZN(n3059) );
  XNOR2_X1 U10477 ( .A(n25638), .B(n28319), .ZN(n6807) );
  AND3_X1 U10479 ( .A1(n28989), .A2(n29018), .A3(n28933), .ZN(n4143) );
  INV_X1 U10480 ( .A(n28879), .ZN(n29038) );
  INV_X1 U10482 ( .A(n25841), .ZN(n3124) );
  OR2_X1 U10483 ( .A1(n29882), .A2(n29782), .ZN(n4320) );
  OR2_X1 U10484 ( .A1(n28623), .A2(n4075), .ZN(n29520) );
  INV_X1 U10485 ( .A(n28757), .ZN(n4493) );
  AND2_X1 U10487 ( .A1(n27956), .A2(n5168), .ZN(n8582) );
  INV_X1 U10488 ( .A(n41272), .ZN(n6927) );
  NOR2_X1 U10489 ( .A1(n30082), .A2(n3099), .ZN(n3394) );
  OAI21_X1 U10490 ( .B1(n27687), .B2(n2611), .A(n26956), .ZN(n26957) );
  AND2_X1 U10491 ( .A1(n30773), .A2(n29921), .ZN(n26930) );
  OAI211_X1 U10493 ( .C1(n27657), .C2(n2671), .A(n8290), .B(n27065), .ZN(n2670) );
  AND2_X1 U10494 ( .A1(n27070), .A2(n27671), .ZN(n2671) );
  INV_X1 U10497 ( .A(n6403), .ZN(n30425) );
  XNOR2_X1 U10498 ( .A(n28068), .B(n3234), .ZN(n30431) );
  XNOR2_X1 U10499 ( .A(n2255), .B(n27478), .ZN(n3234) );
  OR2_X1 U10500 ( .A1(n30412), .A2(n30403), .ZN(n30406) );
  INV_X1 U10501 ( .A(n30268), .ZN(n29110) );
  INV_X1 U10502 ( .A(n30226), .ZN(n29254) );
  XNOR2_X1 U10503 ( .A(n6943), .B(n26287), .ZN(n6945) );
  INV_X1 U10504 ( .A(n25934), .ZN(n6944) );
  AND2_X1 U10505 ( .A1(n32587), .A2(n29618), .ZN(n3952) );
  AND2_X1 U10506 ( .A1(n28659), .A2(n4724), .ZN(n29261) );
  NAND4_X1 U10508 ( .A1(n29311), .A2(n29310), .A3(n29308), .A4(n29309), .ZN(
        n3915) );
  OR2_X1 U10509 ( .A1(n32840), .A2(n31911), .ZN(n32836) );
  AND2_X1 U10511 ( .A1(n25418), .A2(n7123), .ZN(n8720) );
  AND2_X1 U10512 ( .A1(n32895), .A2(n32633), .ZN(n4173) );
  OR2_X1 U10513 ( .A1(n26843), .A2(n30769), .ZN(n29918) );
  AND2_X1 U10514 ( .A1(n26887), .A2(n27730), .ZN(n8055) );
  INV_X1 U10515 ( .A(n26458), .ZN(n29015) );
  NOR2_X1 U10516 ( .A1(n32089), .A2(n32107), .ZN(n32106) );
  INV_X1 U10517 ( .A(n30387), .ZN(n30394) );
  INV_X1 U10518 ( .A(n31497), .ZN(n3225) );
  INV_X1 U10519 ( .A(n31300), .ZN(n30644) );
  OAI21_X1 U10520 ( .B1(n26478), .B2(n28903), .A(n28905), .ZN(n6547) );
  OR2_X1 U10521 ( .A1(n27987), .A2(n51118), .ZN(n4751) );
  INV_X1 U10522 ( .A(n26619), .ZN(n29030) );
  INV_X1 U10523 ( .A(n30647), .ZN(n4607) );
  AND2_X1 U10525 ( .A1(n29438), .A2(n2213), .ZN(n7474) );
  INV_X1 U10526 ( .A(n6602), .ZN(n6303) );
  OR2_X1 U10527 ( .A1(n31538), .A2(n32665), .ZN(n31547) );
  AND2_X1 U10528 ( .A1(n32559), .A2(n32560), .ZN(n29355) );
  INV_X1 U10529 ( .A(n32204), .ZN(n31769) );
  AND2_X1 U10530 ( .A1(n30360), .A2(n29781), .ZN(n3433) );
  INV_X1 U10531 ( .A(n30125), .ZN(n28489) );
  AND2_X1 U10532 ( .A1(n30119), .A2(n3102), .ZN(n25986) );
  OAI21_X1 U10533 ( .B1(n31874), .B2(n31870), .A(n3103), .ZN(n3102) );
  AND2_X1 U10534 ( .A1(n31873), .A2(n31886), .ZN(n3103) );
  OR2_X1 U10535 ( .A1(n28953), .A2(n29789), .ZN(n4264) );
  NAND2_X1 U10536 ( .A1(n29327), .A2(n25975), .ZN(n29329) );
  NOR2_X1 U10537 ( .A1(n30602), .A2(n5278), .ZN(n30608) );
  INV_X1 U10538 ( .A(n30651), .ZN(n4936) );
  AND3_X1 U10539 ( .A1(n29891), .A2(n29888), .A3(n29889), .ZN(n4695) );
  OR4_X1 U10540 ( .A1(n32233), .A2(n32254), .A3(n32251), .A4(n32252), .ZN(
        n32234) );
  INV_X1 U10541 ( .A(n5442), .ZN(n5439) );
  AND2_X1 U10542 ( .A1(n32251), .A2(n32242), .ZN(n32239) );
  INV_X1 U10543 ( .A(n29372), .ZN(n32253) );
  OAI21_X1 U10544 ( .B1(n26947), .B2(n27659), .A(n27658), .ZN(n8691) );
  INV_X1 U10545 ( .A(n32239), .ZN(n31783) );
  OR2_X1 U10546 ( .A1(n32485), .A2(n32025), .ZN(n8345) );
  OAI21_X1 U10547 ( .B1(n5769), .B2(n5768), .A(n5767), .ZN(n32019) );
  INV_X1 U10548 ( .A(n31569), .ZN(n32617) );
  AND2_X1 U10549 ( .A1(n31055), .A2(n31512), .ZN(n4184) );
  OAI21_X1 U10551 ( .B1(n26884), .B2(n2983), .A(n2982), .ZN(n26886) );
  OR2_X1 U10552 ( .A1(n27627), .A2(n27623), .ZN(n2983) );
  NAND2_X1 U10554 ( .A1(n32986), .A2(n32595), .ZN(n2746) );
  INV_X1 U10555 ( .A(n32379), .ZN(n32380) );
  AND2_X1 U10556 ( .A1(n30915), .A2(n30911), .ZN(n30914) );
  AND2_X1 U10557 ( .A1(n26708), .A2(n30846), .ZN(n3687) );
  INV_X1 U10558 ( .A(n8517), .ZN(n31379) );
  AND2_X1 U10559 ( .A1(n4434), .A2(n435), .ZN(n31846) );
  AND2_X1 U10560 ( .A1(n51105), .A2(n30873), .ZN(n32502) );
  OR2_X1 U10561 ( .A1(n31608), .A2(n32558), .ZN(n30901) );
  OR2_X1 U10562 ( .A1(n29840), .A2(n30110), .ZN(n4848) );
  INV_X1 U10563 ( .A(n30940), .ZN(n30070) );
  AND2_X1 U10564 ( .A1(n33014), .A2(n31383), .ZN(n29635) );
  AND2_X1 U10565 ( .A1(n29620), .A2(n6242), .ZN(n6239) );
  INV_X1 U10566 ( .A(n30513), .ZN(n6242) );
  AND2_X1 U10567 ( .A1(n28723), .A2(n30853), .ZN(n3951) );
  AND2_X1 U10568 ( .A1(n33017), .A2(n8517), .ZN(n8516) );
  INV_X1 U10569 ( .A(n33019), .ZN(n7542) );
  AOI21_X1 U10570 ( .B1(n31794), .B2(n31793), .A(n31882), .ZN(n31795) );
  OAI21_X1 U10571 ( .B1(n32485), .B2(n32473), .A(n32472), .ZN(n32474) );
  INV_X1 U10572 ( .A(n32906), .ZN(n30822) );
  OR2_X1 U10574 ( .A1(n30576), .A2(n30846), .ZN(n30577) );
  NOR2_X1 U10575 ( .A1(n32215), .A2(n50981), .ZN(n31763) );
  AND2_X1 U10576 ( .A1(n31580), .A2(n31624), .ZN(n4905) );
  INV_X1 U10577 ( .A(n31298), .ZN(n29652) );
  AND2_X1 U10578 ( .A1(n30628), .A2(n30627), .ZN(n5817) );
  AOI21_X1 U10580 ( .B1(n30983), .B2(n26795), .A(n31680), .ZN(n29966) );
  INV_X1 U10581 ( .A(n30014), .ZN(n30013) );
  INV_X1 U10582 ( .A(n30975), .ZN(n31682) );
  INV_X1 U10583 ( .A(n31510), .ZN(n5698) );
  OR2_X1 U10585 ( .A1(n31161), .A2(n7626), .ZN(n4289) );
  AND2_X1 U10586 ( .A1(n32618), .A2(n31556), .ZN(n5481) );
  INV_X1 U10587 ( .A(n32660), .ZN(n30964) );
  NOR2_X1 U10588 ( .A1(n31385), .A2(n33002), .ZN(n3177) );
  NOR2_X1 U10589 ( .A1(n31385), .A2(n720), .ZN(n33004) );
  AND2_X1 U10591 ( .A1(n31418), .A2(n29655), .ZN(n29994) );
  INV_X1 U10592 ( .A(n29995), .ZN(n31151) );
  OAI21_X1 U10593 ( .B1(n27984), .B2(n27983), .A(n27982), .ZN(n7750) );
  NOR2_X1 U10594 ( .A1(n29685), .A2(n31089), .ZN(n6891) );
  AND3_X1 U10597 ( .A1(n32429), .A2(n32428), .A3(n32814), .ZN(n6746) );
  AND2_X1 U10598 ( .A1(n31218), .A2(n32210), .ZN(n29104) );
  INV_X1 U10599 ( .A(n32356), .ZN(n32453) );
  OAI21_X1 U10600 ( .B1(n32638), .B2(n32639), .A(n8088), .ZN(n32640) );
  INV_X1 U10601 ( .A(n32896), .ZN(n8088) );
  OR2_X1 U10603 ( .A1(n31558), .A2(n7064), .ZN(n5038) );
  OR2_X1 U10604 ( .A1(n31236), .A2(n32230), .ZN(n6118) );
  OAI211_X1 U10605 ( .C1(n8277), .C2(n31561), .A(n31558), .B(n31564), .ZN(
        n8276) );
  INV_X1 U10607 ( .A(n31561), .ZN(n30330) );
  OAI21_X1 U10608 ( .B1(n31026), .B2(n31874), .A(n31880), .ZN(n30124) );
  OR2_X1 U10609 ( .A1(n32848), .A2(n31910), .ZN(n30492) );
  AND2_X1 U10610 ( .A1(n32164), .A2(n3064), .ZN(n3063) );
  OR2_X1 U10611 ( .A1(n32798), .A2(n32797), .ZN(n4370) );
  NOR2_X1 U10612 ( .A1(n29212), .A2(n32395), .ZN(n3886) );
  INV_X1 U10613 ( .A(n31955), .ZN(n32042) );
  OR2_X1 U10614 ( .A1(n32770), .A2(n3303), .ZN(n32775) );
  AND3_X1 U10615 ( .A1(n32956), .A2(n32771), .A3(n3035), .ZN(n3810) );
  INV_X1 U10617 ( .A(n31793), .ZN(n31880) );
  OR2_X1 U10618 ( .A1(n31662), .A2(n32327), .ZN(n4334) );
  INV_X1 U10619 ( .A(n29648), .ZN(n31051) );
  NOR2_X1 U10620 ( .A1(n31055), .A2(n5326), .ZN(n31062) );
  INV_X1 U10621 ( .A(n31777), .ZN(n32226) );
  INV_X1 U10622 ( .A(n33711), .ZN(n33218) );
  INV_X1 U10623 ( .A(n30036), .ZN(n30033) );
  AND2_X1 U10624 ( .A1(n32133), .A2(n32140), .ZN(n8223) );
  AND3_X1 U10625 ( .A1(n26798), .A2(n26797), .A3(n30012), .ZN(n3420) );
  INV_X1 U10626 ( .A(n35656), .ZN(n37015) );
  OR2_X1 U10627 ( .A1(n8536), .A2(n51618), .ZN(n31400) );
  AND2_X1 U10628 ( .A1(n31904), .A2(n31401), .ZN(n7408) );
  AND2_X1 U10629 ( .A1(n8517), .A2(n51740), .ZN(n6420) );
  AND2_X1 U10631 ( .A1(n32190), .A2(n32188), .ZN(n4044) );
  INV_X1 U10632 ( .A(n32491), .ZN(n32483) );
  XNOR2_X1 U10633 ( .A(n33753), .B(n4737), .ZN(n3986) );
  AND2_X1 U10634 ( .A1(n6458), .A2(n6460), .ZN(n5123) );
  AND2_X1 U10635 ( .A1(n31952), .A2(n32069), .ZN(n4085) );
  INV_X1 U10637 ( .A(n31205), .ZN(n32492) );
  NOR2_X1 U10638 ( .A1(n30052), .A2(n2365), .ZN(n8292) );
  OR2_X1 U10639 ( .A1(n32661), .A2(n31538), .ZN(n31176) );
  NOR2_X1 U10640 ( .A1(n5868), .A2(n32665), .ZN(n31177) );
  NOR2_X1 U10641 ( .A1(n5867), .A2(n5868), .ZN(n31165) );
  AND2_X1 U10642 ( .A1(n32545), .A2(n32544), .ZN(n4234) );
  NOR2_X1 U10643 ( .A1(n31755), .A2(n31754), .ZN(n7829) );
  INV_X1 U10644 ( .A(n34116), .ZN(n36701) );
  AND2_X1 U10645 ( .A1(n32222), .A2(n32220), .ZN(n4318) );
  BUF_X1 U10646 ( .A(n33728), .Z(n35387) );
  XNOR2_X1 U10647 ( .A(n35282), .B(n51366), .ZN(n35490) );
  AND4_X1 U10648 ( .A1(n31008), .A2(n3920), .A3(n31004), .A4(n31009), .ZN(
        n3919) );
  INV_X1 U10649 ( .A(n31003), .ZN(n3923) );
  AND2_X1 U10650 ( .A1(n8538), .A2(n30479), .ZN(n8537) );
  XNOR2_X1 U10651 ( .A(n35240), .B(n34452), .ZN(n6858) );
  INV_X1 U10652 ( .A(n35403), .ZN(n3719) );
  INV_X1 U10653 ( .A(n33306), .ZN(n35289) );
  XNOR2_X1 U10654 ( .A(n4224), .B(n35586), .ZN(n35260) );
  INV_X1 U10655 ( .A(n32909), .ZN(n32894) );
  AND2_X1 U10656 ( .A1(n33006), .A2(n31383), .ZN(n30542) );
  OR2_X1 U10657 ( .A1(n33014), .A2(n31383), .ZN(n31012) );
  AND2_X1 U10658 ( .A1(n30986), .A2(n30987), .ZN(n2974) );
  OAI21_X1 U10659 ( .B1(n30977), .B2(n30978), .A(n30976), .ZN(n30989) );
  INV_X1 U10660 ( .A(n29650), .ZN(n31313) );
  INV_X1 U10661 ( .A(n30830), .ZN(n30835) );
  INV_X1 U10662 ( .A(n35586), .ZN(n33578) );
  INV_X1 U10663 ( .A(n6760), .ZN(n6559) );
  XNOR2_X1 U10664 ( .A(n35254), .B(n34811), .ZN(n36951) );
  INV_X1 U10665 ( .A(n37264), .ZN(n7360) );
  INV_X1 U10666 ( .A(n36248), .ZN(n7083) );
  AND2_X1 U10667 ( .A1(n6321), .A2(n31029), .ZN(n2843) );
  OR2_X1 U10668 ( .A1(n30012), .A2(n30983), .ZN(n30027) );
  INV_X1 U10669 ( .A(n37991), .ZN(n36534) );
  AND2_X1 U10670 ( .A1(n32137), .A2(n5100), .ZN(n6066) );
  INV_X1 U10671 ( .A(n31716), .ZN(n6065) );
  OR2_X1 U10672 ( .A1(n31644), .A2(n8548), .ZN(n8545) );
  XNOR2_X1 U10673 ( .A(n37269), .B(n37096), .ZN(n36962) );
  INV_X1 U10674 ( .A(n36328), .ZN(n7400) );
  NOR2_X1 U10675 ( .A1(n2321), .A2(n4770), .ZN(n4769) );
  INV_X1 U10676 ( .A(n35240), .ZN(n37114) );
  INV_X1 U10677 ( .A(n32000), .ZN(n2755) );
  XNOR2_X1 U10678 ( .A(n8595), .B(n34240), .ZN(n37256) );
  INV_X1 U10679 ( .A(n34533), .ZN(n8595) );
  XNOR2_X1 U10680 ( .A(n4421), .B(n34238), .ZN(n33489) );
  XNOR2_X1 U10681 ( .A(n35247), .B(n33326), .ZN(n4421) );
  XNOR2_X1 U10682 ( .A(n31575), .B(n31574), .ZN(n34810) );
  AND2_X1 U10683 ( .A1(n36122), .A2(n38599), .ZN(n3940) );
  INV_X1 U10685 ( .A(n37453), .ZN(n3211) );
  INV_X1 U10686 ( .A(n34535), .ZN(n33337) );
  XNOR2_X1 U10687 ( .A(n5648), .B(n5999), .ZN(n37134) );
  AND2_X1 U10689 ( .A1(n37731), .A2(n39003), .ZN(n4693) );
  INV_X1 U10690 ( .A(n36529), .ZN(n3654) );
  XNOR2_X1 U10691 ( .A(n34135), .B(n34130), .ZN(n7126) );
  NAND2_X1 U10692 ( .A1(n35943), .A2(n35940), .ZN(n6982) );
  INV_X1 U10693 ( .A(n38322), .ZN(n6615) );
  INV_X1 U10694 ( .A(n38290), .ZN(n37627) );
  AND2_X1 U10695 ( .A1(n36098), .A2(n35151), .ZN(n5312) );
  AND2_X1 U10696 ( .A1(n29658), .A2(n31420), .ZN(n4697) );
  INV_X1 U10697 ( .A(n39247), .ZN(n4258) );
  OAI211_X1 U10698 ( .C1(n31791), .C2(n3121), .A(n31023), .B(n31022), .ZN(
        n31024) );
  AND2_X1 U10699 ( .A1(n31101), .A2(n31100), .ZN(n2941) );
  AND3_X1 U10700 ( .A1(n31628), .A2(n31627), .A3(n31642), .ZN(n3998) );
  NOR2_X1 U10701 ( .A1(n6522), .A2(n6521), .ZN(n6520) );
  OAI21_X1 U10702 ( .B1(n32533), .B2(n32534), .A(n32963), .ZN(n32537) );
  INV_X1 U10703 ( .A(n34869), .ZN(n8460) );
  INV_X1 U10704 ( .A(n37637), .ZN(n37643) );
  INV_X1 U10705 ( .A(n37647), .ZN(n5588) );
  INV_X1 U10706 ( .A(n37648), .ZN(n5590) );
  AND2_X1 U10707 ( .A1(n6262), .A2(n37646), .ZN(n37645) );
  XNOR2_X1 U10708 ( .A(n34078), .B(n3113), .ZN(n33740) );
  INV_X1 U10709 ( .A(n5234), .ZN(n3113) );
  INV_X1 U10710 ( .A(n39429), .ZN(n36887) );
  INV_X1 U10711 ( .A(n33726), .ZN(n33718) );
  AND2_X1 U10714 ( .A1(n4948), .A2(n39450), .ZN(n36898) );
  INV_X1 U10715 ( .A(n39027), .ZN(n4948) );
  INV_X1 U10716 ( .A(n36898), .ZN(n36259) );
  INV_X1 U10717 ( .A(n39032), .ZN(n39441) );
  INV_X1 U10718 ( .A(n38953), .ZN(n38941) );
  INV_X1 U10719 ( .A(n35214), .ZN(n36054) );
  OR2_X1 U10720 ( .A1(n37664), .A2(n37665), .ZN(n4270) );
  OR2_X1 U10721 ( .A1(n51508), .A2(n6343), .ZN(n39247) );
  OR2_X1 U10722 ( .A1(n39173), .A2(n39172), .ZN(n39175) );
  INV_X1 U10723 ( .A(n8077), .ZN(n5571) );
  AND3_X1 U10724 ( .A1(n36410), .A2(n51334), .A3(n35732), .ZN(n37639) );
  NOR2_X1 U10725 ( .A1(n38270), .A2(n37624), .ZN(n6011) );
  AND2_X1 U10726 ( .A1(n38707), .A2(n39243), .ZN(n4238) );
  INV_X1 U10727 ( .A(n38241), .ZN(n3708) );
  INV_X1 U10728 ( .A(n39169), .ZN(n38245) );
  INV_X1 U10729 ( .A(n38283), .ZN(n36439) );
  XNOR2_X1 U10730 ( .A(n34856), .B(n34043), .ZN(n34044) );
  AND2_X1 U10731 ( .A1(n37964), .A2(n7851), .ZN(n7850) );
  INV_X1 U10732 ( .A(n40874), .ZN(n6525) );
  OR2_X1 U10733 ( .A1(n40863), .A2(n40862), .ZN(n40544) );
  INV_X1 U10734 ( .A(n6541), .ZN(n34969) );
  INV_X1 U10735 ( .A(n37585), .ZN(n37379) );
  INV_X1 U10736 ( .A(n38549), .ZN(n38227) );
  NOR2_X1 U10737 ( .A1(n36141), .A2(n38558), .ZN(n36300) );
  INV_X1 U10738 ( .A(n34193), .ZN(n34184) );
  INV_X1 U10739 ( .A(n36312), .ZN(n36628) );
  OR2_X1 U10740 ( .A1(n38593), .A2(n38585), .ZN(n37452) );
  AND2_X1 U10741 ( .A1(n36427), .A2(n36428), .ZN(n4576) );
  OR2_X1 U10742 ( .A1(n51360), .A2(n38630), .ZN(n3946) );
  OR2_X1 U10743 ( .A1(n2049), .A2(n34963), .ZN(n6904) );
  OR2_X1 U10744 ( .A1(n38549), .A2(n38214), .ZN(n5980) );
  OR2_X1 U10745 ( .A1(n38218), .A2(n36142), .ZN(n36309) );
  AND2_X1 U10746 ( .A1(n38810), .A2(n41796), .ZN(n38819) );
  INV_X1 U10747 ( .A(n6638), .ZN(n36398) );
  INV_X1 U10748 ( .A(n2714), .ZN(n5741) );
  INV_X1 U10749 ( .A(n38557), .ZN(n6735) );
  INV_X1 U10751 ( .A(n41332), .ZN(n41316) );
  AND3_X1 U10752 ( .A1(n39269), .A2(n39270), .A3(n39268), .ZN(n2570) );
  OR2_X1 U10753 ( .A1(n41693), .A2(n41692), .ZN(n41709) );
  INV_X1 U10754 ( .A(n34629), .ZN(n34632) );
  OR2_X1 U10755 ( .A1(n36586), .A2(n35209), .ZN(n35878) );
  XNOR2_X1 U10756 ( .A(n7364), .B(n7508), .ZN(n2691) );
  AND2_X1 U10757 ( .A1(n2855), .A2(n6851), .ZN(n39978) );
  AND2_X1 U10758 ( .A1(n37526), .A2(n38496), .ZN(n6996) );
  NAND2_X1 U10759 ( .A1(n37518), .A2(n38504), .ZN(n6109) );
  AND2_X1 U10760 ( .A1(n37532), .A2(n37531), .ZN(n6995) );
  OR2_X1 U10761 ( .A1(n37644), .A2(n37643), .ZN(n4352) );
  INV_X1 U10762 ( .A(n39227), .ZN(n38699) );
  INV_X1 U10763 ( .A(n39219), .ZN(n37697) );
  OR2_X1 U10764 ( .A1(n35972), .A2(n3044), .ZN(n37366) );
  AND2_X1 U10765 ( .A1(n40768), .A2(n40777), .ZN(n39800) );
  NOR2_X1 U10766 ( .A1(n38504), .A2(n37387), .ZN(n5729) );
  OR2_X1 U10767 ( .A1(n37385), .A2(n38496), .ZN(n5730) );
  NOR2_X1 U10768 ( .A1(n618), .A2(n38504), .ZN(n5808) );
  INV_X1 U10769 ( .A(n39204), .ZN(n39428) );
  AND2_X1 U10770 ( .A1(n36240), .A2(n37757), .ZN(n5942) );
  XNOR2_X1 U10771 ( .A(n35284), .B(n37005), .ZN(n38638) );
  AND2_X1 U10772 ( .A1(n36232), .A2(n35973), .ZN(n4235) );
  OR2_X1 U10773 ( .A1(n36320), .A2(n34187), .ZN(n4162) );
  OR2_X1 U10774 ( .A1(n40470), .A2(n41268), .ZN(n40482) );
  INV_X1 U10776 ( .A(n6980), .ZN(n40251) );
  INV_X1 U10777 ( .A(n41079), .ZN(n39144) );
  OR2_X1 U10778 ( .A1(n2787), .A2(n2784), .ZN(n2783) );
  INV_X1 U10780 ( .A(n40499), .ZN(n39131) );
  OR2_X1 U10781 ( .A1(n40453), .A2(n2848), .ZN(n39738) );
  OAI21_X1 U10782 ( .B1(n41698), .B2(n41693), .A(n7137), .ZN(n8192) );
  NOR2_X1 U10784 ( .A1(n40396), .A2(n6850), .ZN(n40400) );
  INV_X1 U10785 ( .A(n38909), .ZN(n40644) );
  INV_X1 U10786 ( .A(n41435), .ZN(n40655) );
  OAI21_X1 U10787 ( .B1(n40536), .B2(n40860), .A(n40535), .ZN(n5597) );
  OR2_X1 U10788 ( .A1(n40533), .A2(n40534), .ZN(n5596) );
  OR2_X1 U10789 ( .A1(n40526), .A2(n40869), .ZN(n40857) );
  AND2_X1 U10790 ( .A1(n40909), .A2(n40081), .ZN(n40275) );
  INV_X1 U10791 ( .A(n40909), .ZN(n3655) );
  INV_X1 U10792 ( .A(n40500), .ZN(n6392) );
  AND2_X1 U10793 ( .A1(n8256), .A2(n40862), .ZN(n39968) );
  INV_X1 U10794 ( .A(n40544), .ZN(n40540) );
  INV_X1 U10796 ( .A(n40903), .ZN(n5072) );
  INV_X1 U10797 ( .A(n40275), .ZN(n40097) );
  INV_X1 U10798 ( .A(n40785), .ZN(n40776) );
  AND2_X1 U10799 ( .A1(n40420), .A2(n41276), .ZN(n40421) );
  INV_X1 U10800 ( .A(n41039), .ZN(n8615) );
  INV_X1 U10801 ( .A(n40960), .ZN(n38885) );
  AOI22_X1 U10802 ( .A1(n35718), .A2(n40571), .B1(n35719), .B2(n40566), .ZN(
        n4068) );
  INV_X1 U10803 ( .A(n41902), .ZN(n8235) );
  AOI22_X1 U10804 ( .A1(n41325), .A2(n41326), .B1(n41327), .B2(n5316), .ZN(
        n41336) );
  AND2_X1 U10805 ( .A1(n40198), .A2(n40119), .ZN(n6185) );
  AND2_X1 U10806 ( .A1(n38773), .A2(n40125), .ZN(n2900) );
  NOR2_X1 U10807 ( .A1(n3831), .A2(n4943), .ZN(n2973) );
  INV_X1 U10808 ( .A(n41573), .ZN(n42002) );
  AND2_X1 U10809 ( .A1(n40738), .A2(n40739), .ZN(n40748) );
  INV_X1 U10810 ( .A(n41345), .ZN(n40357) );
  INV_X1 U10811 ( .A(n39768), .ZN(n7704) );
  OAI21_X1 U10812 ( .B1(n38931), .B2(n41931), .A(n41942), .ZN(n3029) );
  INV_X1 U10813 ( .A(n38809), .ZN(n6062) );
  AND2_X1 U10814 ( .A1(n38810), .A2(n38815), .ZN(n6061) );
  NOR2_X1 U10815 ( .A1(n43665), .A2(n3936), .ZN(n38820) );
  OR2_X1 U10816 ( .A1(n40632), .A2(n41792), .ZN(n3936) );
  INV_X1 U10817 ( .A(n41725), .ZN(n41726) );
  OR2_X1 U10818 ( .A1(n3771), .A2(n40366), .ZN(n3681) );
  INV_X1 U10820 ( .A(n39873), .ZN(n41609) );
  INV_X1 U10821 ( .A(n4683), .ZN(n4682) );
  OAI21_X1 U10822 ( .B1(n41695), .B2(n41702), .A(n41693), .ZN(n4683) );
  NOR2_X1 U10823 ( .A1(n41544), .A2(n40943), .ZN(n5215) );
  INV_X1 U10824 ( .A(n40981), .ZN(n40936) );
  INV_X1 U10825 ( .A(n41389), .ZN(n41388) );
  OR2_X1 U10827 ( .A1(n36457), .A2(n36585), .ZN(n34410) );
  AND2_X1 U10828 ( .A1(n41483), .A2(n42041), .ZN(n39067) );
  AND2_X1 U10829 ( .A1(n37660), .A2(n37662), .ZN(n7490) );
  OR2_X1 U10830 ( .A1(n36233), .A2(n37585), .ZN(n37380) );
  AND2_X1 U10831 ( .A1(n37402), .A2(n37401), .ZN(n5806) );
  OAI21_X1 U10832 ( .B1(n38533), .B2(n37435), .A(n37446), .ZN(n5964) );
  INV_X1 U10833 ( .A(n40986), .ZN(n41524) );
  OAI21_X1 U10834 ( .B1(n38925), .B2(n6580), .A(n2744), .ZN(n7174) );
  AND2_X1 U10835 ( .A1(n41065), .A2(n39129), .ZN(n41051) );
  INV_X1 U10836 ( .A(n41082), .ZN(n39140) );
  NOR2_X1 U10837 ( .A1(n42149), .A2(n41764), .ZN(n7424) );
  AND3_X1 U10838 ( .A1(n4399), .A2(n41766), .A3(n4398), .ZN(n6840) );
  OR2_X1 U10839 ( .A1(n34662), .A2(n8011), .ZN(n8010) );
  INV_X1 U10840 ( .A(n40342), .ZN(n40329) );
  OR2_X2 U10841 ( .A1(n34318), .A2(n34317), .ZN(n40338) );
  INV_X1 U10842 ( .A(n40016), .ZN(n3751) );
  OAI21_X1 U10843 ( .B1(n39127), .B2(n40511), .A(n39126), .ZN(n3440) );
  OR2_X1 U10845 ( .A1(n40120), .A2(n40204), .ZN(n3093) );
  AND2_X1 U10846 ( .A1(n40250), .A2(n2738), .ZN(n6580) );
  OR2_X1 U10847 ( .A1(n2738), .A2(n40250), .ZN(n2737) );
  NAND2_X1 U10848 ( .A1(n41051), .A2(n610), .ZN(n6212) );
  OR2_X1 U10849 ( .A1(n39759), .A2(n3231), .ZN(n41607) );
  INV_X1 U10850 ( .A(n8754), .ZN(n7986) );
  INV_X1 U10851 ( .A(n41539), .ZN(n40989) );
  AOI21_X1 U10852 ( .B1(n4561), .B2(n41736), .A(n41259), .ZN(n41632) );
  OR2_X1 U10853 ( .A1(n41706), .A2(n41692), .ZN(n41172) );
  AOI21_X1 U10854 ( .B1(n40015), .B2(n39097), .A(n39099), .ZN(n39666) );
  INV_X1 U10855 ( .A(n6884), .ZN(n2834) );
  AND3_X1 U10856 ( .A1(n41697), .A2(n41690), .A3(n2179), .ZN(n8194) );
  NAND2_X1 U10857 ( .A1(n39043), .A2(n40353), .ZN(n8195) );
  AND2_X1 U10858 ( .A1(n6370), .A2(n38840), .ZN(n6372) );
  AND2_X1 U10859 ( .A1(n6375), .A2(n38839), .ZN(n6374) );
  OR2_X1 U10860 ( .A1(n39943), .A2(n575), .ZN(n6375) );
  NOR2_X1 U10861 ( .A1(n51012), .A2(n40377), .ZN(n4116) );
  AND2_X1 U10862 ( .A1(n41802), .A2(n42105), .ZN(n8271) );
  INV_X1 U10863 ( .A(n41509), .ZN(n41504) );
  NOR2_X1 U10864 ( .A1(n51297), .A2(n39097), .ZN(n39095) );
  INV_X1 U10865 ( .A(n41268), .ZN(n41124) );
  AND2_X1 U10866 ( .A1(n41682), .A2(n41681), .ZN(n5576) );
  OR2_X1 U10867 ( .A1(n6886), .A2(n39100), .ZN(n6881) );
  NOR2_X1 U10868 ( .A1(n6427), .A2(n8673), .ZN(n8672) );
  OAI21_X1 U10869 ( .B1(n41579), .B2(n41578), .A(n41577), .ZN(n8671) );
  INV_X1 U10870 ( .A(n40751), .ZN(n39884) );
  XNOR2_X1 U10871 ( .A(n42560), .B(n7384), .ZN(n45250) );
  INV_X1 U10872 ( .A(n4647), .ZN(n7384) );
  INV_X1 U10873 ( .A(n43703), .ZN(n7101) );
  INV_X1 U10874 ( .A(n42135), .ZN(n41747) );
  NAND4_X1 U10875 ( .A1(n40244), .A2(n40246), .A3(n40243), .A4(n40245), .ZN(
        n5824) );
  INV_X1 U10876 ( .A(n35004), .ZN(n40502) );
  INV_X1 U10877 ( .A(n5884), .ZN(n41045) );
  INV_X1 U10878 ( .A(n41330), .ZN(n6325) );
  AND2_X1 U10879 ( .A1(n42018), .A2(n41589), .ZN(n41412) );
  OR2_X1 U10880 ( .A1(n41509), .A2(n41415), .ZN(n41420) );
  OAI21_X1 U10881 ( .B1(n5747), .B2(n40860), .A(n40535), .ZN(n39965) );
  AND2_X1 U10882 ( .A1(n41375), .A2(n40960), .ZN(n3796) );
  AND3_X1 U10883 ( .A1(n40093), .A2(n40092), .A3(n40091), .ZN(n40102) );
  INV_X1 U10884 ( .A(n40081), .ZN(n8597) );
  OR2_X1 U10885 ( .A1(n40130), .A2(n40131), .ZN(n4280) );
  NAND4_X1 U10886 ( .A1(n39734), .A2(n39732), .A3(n39733), .A4(n5436), .ZN(
        n39735) );
  OAI21_X1 U10887 ( .B1(n41804), .B2(n43669), .A(n40633), .ZN(n40634) );
  INV_X1 U10888 ( .A(n40968), .ZN(n41373) );
  INV_X1 U10889 ( .A(n40736), .ZN(n39882) );
  INV_X1 U10890 ( .A(n38745), .ZN(n39895) );
  INV_X1 U10891 ( .A(n40746), .ZN(n40744) );
  INV_X1 U10892 ( .A(n40653), .ZN(n41448) );
  AND2_X1 U10893 ( .A1(n4871), .A2(n2393), .ZN(n37176) );
  XNOR2_X1 U10894 ( .A(n45089), .B(n43110), .ZN(n43111) );
  XNOR2_X1 U10895 ( .A(n45091), .B(n44098), .ZN(n43360) );
  OR2_X1 U10896 ( .A1(n38620), .A2(n2653), .ZN(n33282) );
  AND2_X1 U10897 ( .A1(n6998), .A2(n39581), .ZN(n4096) );
  INV_X1 U10898 ( .A(n2597), .ZN(n40321) );
  NOR2_X1 U10899 ( .A1(n37824), .A2(n40250), .ZN(n42206) );
  INV_X1 U10900 ( .A(n4862), .ZN(n41930) );
  INV_X1 U10901 ( .A(n39902), .ZN(n39915) );
  NOR2_X1 U10902 ( .A1(n39907), .A2(n38445), .ZN(n39919) );
  INV_X1 U10903 ( .A(n43547), .ZN(n46049) );
  OAI21_X1 U10904 ( .B1(n4861), .B2(n41933), .A(n4236), .ZN(n40256) );
  AND2_X1 U10905 ( .A1(n41080), .A2(n8219), .ZN(n8218) );
  INV_X1 U10907 ( .A(n44217), .ZN(n43703) );
  OAI211_X1 U10908 ( .C1(n41977), .C2(n41971), .A(n41644), .B(n6939), .ZN(
        n5091) );
  AND2_X1 U10909 ( .A1(n5090), .A2(n41653), .ZN(n5092) );
  INV_X1 U10910 ( .A(n40534), .ZN(n40859) );
  INV_X1 U10911 ( .A(n42006), .ZN(n42015) );
  OR2_X1 U10913 ( .A1(n42006), .A2(n6236), .ZN(n6235) );
  AND3_X1 U10914 ( .A1(n33997), .A2(n36079), .A3(n33998), .ZN(n4355) );
  AND2_X1 U10915 ( .A1(n8608), .A2(n40340), .ZN(n37867) );
  AND2_X1 U10916 ( .A1(n39873), .A2(n2867), .ZN(n41611) );
  INV_X1 U10917 ( .A(n41615), .ZN(n5043) );
  AND3_X1 U10918 ( .A1(n38408), .A2(n38407), .A3(n5402), .ZN(n5401) );
  INV_X1 U10919 ( .A(n44176), .ZN(n45460) );
  AND2_X1 U10920 ( .A1(n34918), .A2(n8108), .ZN(n8107) );
  XNOR2_X1 U10921 ( .A(n43236), .B(n43954), .ZN(n42576) );
  OAI21_X1 U10922 ( .B1(n40314), .B2(n40566), .A(n4953), .ZN(n39656) );
  AND3_X1 U10923 ( .A1(n43334), .A2(n39618), .A3(n39619), .ZN(n6595) );
  AND2_X1 U10924 ( .A1(n4763), .A2(n40265), .ZN(n3471) );
  NOR2_X1 U10926 ( .A1(n52169), .A2(n51513), .ZN(n45844) );
  XNOR2_X1 U10927 ( .A(n42038), .B(n42037), .ZN(n42180) );
  INV_X1 U10928 ( .A(n45790), .ZN(n3108) );
  OR2_X1 U10929 ( .A1(n42181), .A2(n3627), .ZN(n44822) );
  XNOR2_X1 U10930 ( .A(n42278), .B(n2552), .ZN(n5435) );
  AND2_X1 U10931 ( .A1(n48259), .A2(n39812), .ZN(n48432) );
  XNOR2_X1 U10933 ( .A(n44338), .B(n7622), .ZN(n42486) );
  INV_X1 U10934 ( .A(n46471), .ZN(n46478) );
  AND2_X1 U10935 ( .A1(n40035), .A2(n41212), .ZN(n6145) );
  OR2_X1 U10936 ( .A1(n49137), .A2(n51515), .ZN(n7656) );
  XNOR2_X1 U10937 ( .A(n42636), .B(n6326), .ZN(n43377) );
  INV_X1 U10938 ( .A(n44147), .ZN(n6326) );
  AND2_X1 U10939 ( .A1(n37471), .A2(n39654), .ZN(n6198) );
  INV_X1 U10940 ( .A(n3149), .ZN(n3148) );
  OAI21_X1 U10941 ( .B1(n51684), .B2(n40632), .A(n43669), .ZN(n3149) );
  XNOR2_X1 U10942 ( .A(n42942), .B(n42941), .ZN(n3757) );
  INV_X1 U10943 ( .A(n43432), .ZN(n49199) );
  AND2_X1 U10944 ( .A1(n49979), .A2(n49989), .ZN(n3278) );
  OAI211_X1 U10945 ( .C1(n39760), .C2(n8070), .A(n39958), .B(n39957), .ZN(
        n5476) );
  OAI21_X1 U10946 ( .B1(n40039), .B2(n40038), .A(n41670), .ZN(n7609) );
  AND2_X1 U10947 ( .A1(n40041), .A2(n2768), .ZN(n2767) );
  NAND3_X1 U10949 ( .A1(n49731), .A2(n423), .A3(n51058), .ZN(n5089) );
  NOR2_X1 U10950 ( .A1(n49987), .A2(n49980), .ZN(n7640) );
  XNOR2_X1 U10951 ( .A(n42519), .B(n42518), .ZN(n46077) );
  AND2_X1 U10952 ( .A1(n5013), .A2(n5012), .ZN(n5010) );
  INV_X1 U10953 ( .A(n5017), .ZN(n5015) );
  OAI21_X1 U10954 ( .B1(n41231), .B2(n41681), .A(n331), .ZN(n39317) );
  XNOR2_X1 U10955 ( .A(n43547), .B(n2551), .ZN(n6425) );
  XNOR2_X1 U10956 ( .A(n7849), .B(n45327), .ZN(n43320) );
  NAND4_X1 U10957 ( .A1(n41974), .A2(n41100), .A3(n41983), .A4(n41099), .ZN(
        n6542) );
  AND2_X1 U10958 ( .A1(n41106), .A2(n41107), .ZN(n6543) );
  AND2_X1 U10959 ( .A1(n40018), .A2(n40017), .ZN(n8372) );
  OR2_X1 U10961 ( .A1(n43345), .A2(n43346), .ZN(n4813) );
  AND3_X1 U10962 ( .A1(n42437), .A2(n42439), .A3(n42440), .ZN(n42447) );
  INV_X1 U10963 ( .A(n44040), .ZN(n7871) );
  AND2_X1 U10964 ( .A1(n658), .A2(n50279), .ZN(n47065) );
  AND3_X1 U10965 ( .A1(n47076), .A2(n7046), .A3(n51404), .ZN(n5592) );
  NOR2_X1 U10966 ( .A1(n49278), .A2(n49266), .ZN(n6025) );
  INV_X1 U10967 ( .A(n46782), .ZN(n6567) );
  INV_X1 U10968 ( .A(n47596), .ZN(n8448) );
  NOR2_X1 U10969 ( .A1(n51344), .A2(n5356), .ZN(n5357) );
  INV_X1 U10970 ( .A(n44873), .ZN(n44654) );
  INV_X1 U10971 ( .A(n46458), .ZN(n44681) );
  OR2_X1 U10972 ( .A1(n44678), .A2(n48481), .ZN(n44685) );
  AND2_X1 U10973 ( .A1(n48546), .A2(n46464), .ZN(n3328) );
  NOR2_X1 U10975 ( .A1(n45574), .A2(n48412), .ZN(n7290) );
  NOR2_X1 U10976 ( .A1(n2341), .A2(n8686), .ZN(n8210) );
  INV_X1 U10979 ( .A(n48539), .ZN(n48237) );
  OR2_X1 U10980 ( .A1(n506), .A2(n48416), .ZN(n48403) );
  INV_X1 U10981 ( .A(n48416), .ZN(n8057) );
  INV_X1 U10983 ( .A(n42796), .ZN(n2716) );
  AND2_X1 U10984 ( .A1(n46380), .A2(n45661), .ZN(n46386) );
  INV_X1 U10987 ( .A(n49714), .ZN(n7797) );
  XNOR2_X1 U10989 ( .A(n44951), .B(n43596), .ZN(n46079) );
  OR2_X1 U10990 ( .A1(n50367), .A2(n3610), .ZN(n46970) );
  INV_X1 U10991 ( .A(n50262), .ZN(n8085) );
  AND2_X1 U10992 ( .A1(n50276), .A2(n50254), .ZN(n2805) );
  INV_X1 U10993 ( .A(n47341), .ZN(n44001) );
  INV_X1 U10994 ( .A(n50252), .ZN(n8451) );
  NAND2_X1 U10995 ( .A1(n6811), .A2(n43797), .ZN(n3610) );
  OR2_X1 U10996 ( .A1(n47139), .A2(n50372), .ZN(n46796) );
  AND2_X1 U10997 ( .A1(n46903), .A2(n46908), .ZN(n46689) );
  OR2_X1 U10998 ( .A1(n47468), .A2(n47586), .ZN(n47265) );
  OR2_X1 U10999 ( .A1(n47617), .A2(n47586), .ZN(n47462) );
  OAI211_X1 U11000 ( .C1(n3106), .C2(n3107), .A(n46713), .B(n44842), .ZN(
        n44844) );
  INV_X1 U11001 ( .A(n46710), .ZN(n3107) );
  AND2_X1 U11002 ( .A1(n44843), .A2(n51396), .ZN(n6888) );
  AND2_X1 U11003 ( .A1(n508), .A2(n47850), .ZN(n6679) );
  OR2_X1 U11004 ( .A1(n48074), .A2(n51092), .ZN(n48038) );
  AND2_X1 U11005 ( .A1(n46633), .A2(n44868), .ZN(n5245) );
  OR2_X1 U11006 ( .A1(n46542), .A2(n48100), .ZN(n48127) );
  NOR2_X1 U11007 ( .A1(n4946), .A2(n52172), .ZN(n48303) );
  INV_X1 U11008 ( .A(n48931), .ZN(n48970) );
  OR2_X1 U11010 ( .A1(n42310), .A2(n49177), .ZN(n7067) );
  AND2_X1 U11011 ( .A1(n49114), .A2(n49119), .ZN(n5661) );
  NOR2_X1 U11012 ( .A1(n49347), .A2(n51729), .ZN(n49363) );
  OR2_X1 U11013 ( .A1(n49347), .A2(n49302), .ZN(n49380) );
  NOR2_X1 U11014 ( .A1(n52107), .A2(n2858), .ZN(n49407) );
  OR2_X1 U11015 ( .A1(n49443), .A2(n51316), .ZN(n49451) );
  AND2_X1 U11016 ( .A1(n47195), .A2(n51091), .ZN(n47192) );
  INV_X1 U11017 ( .A(n49443), .ZN(n49450) );
  AND2_X1 U11018 ( .A1(n49511), .A2(n43490), .ZN(n4572) );
  INV_X1 U11019 ( .A(n43490), .ZN(n3322) );
  AND2_X1 U11020 ( .A1(n49652), .A2(n5763), .ZN(n49655) );
  NAND2_X1 U11021 ( .A1(n49671), .A2(n2725), .ZN(n49658) );
  INV_X1 U11022 ( .A(n49877), .ZN(n46179) );
  INV_X1 U11023 ( .A(n49916), .ZN(n47420) );
  INV_X1 U11025 ( .A(n7503), .ZN(n7502) );
  OR2_X1 U11026 ( .A1(n3864), .A2(n51727), .ZN(n50068) );
  INV_X1 U11027 ( .A(n50145), .ZN(n3864) );
  NAND2_X1 U11028 ( .A1(n8603), .A2(n50145), .ZN(n50142) );
  OR2_X1 U11030 ( .A1(n50192), .A2(n52099), .ZN(n50224) );
  INV_X1 U11032 ( .A(n50637), .ZN(n50578) );
  AND2_X1 U11033 ( .A1(n43579), .A2(n50332), .ZN(n6990) );
  NOR2_X1 U11034 ( .A1(n50779), .A2(n50798), .ZN(n50786) );
  XNOR2_X1 U11035 ( .A(n51730), .B(n51296), .ZN(n7441) );
  AND2_X1 U11036 ( .A1(n51312), .A2(n50837), .ZN(n50848) );
  NAND4_X1 U11037 ( .A1(n51287), .A2(n47572), .A3(n51302), .A4(n47538), .ZN(
        n47490) );
  INV_X1 U11038 ( .A(n47541), .ZN(n5282) );
  AND2_X1 U11039 ( .A1(n2628), .A2(n47265), .ZN(n2627) );
  OR2_X1 U11040 ( .A1(n47266), .A2(n46668), .ZN(n2628) );
  AND2_X1 U11041 ( .A1(n47601), .A2(n2630), .ZN(n2629) );
  AND3_X1 U11042 ( .A1(n47620), .A2(n51401), .A3(n47617), .ZN(n2631) );
  OR2_X1 U11043 ( .A1(n6831), .A2(n47613), .ZN(n5575) );
  AND2_X1 U11044 ( .A1(n47652), .A2(n47655), .ZN(n4223) );
  OR2_X1 U11045 ( .A1(n45858), .A2(n47687), .ZN(n45864) );
  NAND2_X1 U11047 ( .A1(n47676), .A2(n47695), .ZN(n5967) );
  OR2_X1 U11048 ( .A1(n47792), .A2(n47793), .ZN(n47794) );
  OR2_X1 U11049 ( .A1(n47839), .A2(n47873), .ZN(n4397) );
  AND3_X1 U11050 ( .A1(n44711), .A2(n44712), .A3(n5857), .ZN(n44721) );
  OAI21_X1 U11051 ( .B1(n48041), .B2(n48074), .A(n3076), .ZN(n48044) );
  OR2_X1 U11052 ( .A1(n48082), .A2(n48041), .ZN(n48086) );
  OR2_X1 U11053 ( .A1(n8059), .A2(n8062), .ZN(n8058) );
  AND2_X1 U11054 ( .A1(n48095), .A2(n48157), .ZN(n8062) );
  AND2_X1 U11055 ( .A1(n8066), .A2(n4155), .ZN(n8063) );
  OR2_X1 U11056 ( .A1(n48129), .A2(n7766), .ZN(n48139) );
  NAND4_X1 U11057 ( .A1(n3855), .A2(n48142), .A3(n48143), .A4(n3854), .ZN(
        n3856) );
  NOR2_X1 U11058 ( .A1(n48110), .A2(n8690), .ZN(n46540) );
  NOR2_X1 U11059 ( .A1(n48344), .A2(n6987), .ZN(n48319) );
  NOR2_X1 U11060 ( .A1(n8104), .A2(n51728), .ZN(n48351) );
  OAI21_X1 U11061 ( .B1(n48354), .B2(n6987), .A(n48396), .ZN(n48355) );
  AOI22_X1 U11062 ( .A1(n48363), .A2(n48364), .B1(n48361), .B2(n48362), .ZN(
        n48373) );
  AND2_X1 U11063 ( .A1(n48372), .A2(n48370), .ZN(n4632) );
  OAI21_X1 U11064 ( .B1(n48296), .B2(n8103), .A(n8102), .ZN(n8101) );
  INV_X1 U11065 ( .A(n48652), .ZN(n6788) );
  OR2_X1 U11066 ( .A1(n4321), .A2(n48583), .ZN(n48620) );
  INV_X1 U11067 ( .A(n48581), .ZN(n48624) );
  NOR2_X1 U11068 ( .A1(n48695), .A2(n7060), .ZN(n7059) );
  INV_X1 U11069 ( .A(n48696), .ZN(n7060) );
  INV_X1 U11070 ( .A(n994), .ZN(n48782) );
  OAI21_X1 U11071 ( .B1(n48759), .B2(n48734), .A(n52067), .ZN(n3145) );
  OR2_X1 U11072 ( .A1(n48730), .A2(n52067), .ZN(n3144) );
  AND2_X1 U11073 ( .A1(n48801), .A2(n48828), .ZN(n4873) );
  AND3_X1 U11074 ( .A1(n45517), .A2(n45516), .A3(n45741), .ZN(n45518) );
  AND2_X1 U11076 ( .A1(n48905), .A2(n5081), .ZN(n2637) );
  AND2_X1 U11077 ( .A1(n48899), .A2(n5079), .ZN(n48889) );
  AND2_X1 U11078 ( .A1(n48974), .A2(n3208), .ZN(n3210) );
  AND2_X1 U11079 ( .A1(n48957), .A2(n51510), .ZN(n3208) );
  AND2_X1 U11080 ( .A1(n46279), .A2(n49020), .ZN(n2969) );
  OR2_X1 U11081 ( .A1(n8133), .A2(n49019), .ZN(n8131) );
  AND3_X1 U11082 ( .A1(n48996), .A2(n48993), .A3(n49032), .ZN(n4436) );
  AND3_X1 U11083 ( .A1(n7599), .A2(n49101), .A3(n49114), .ZN(n49088) );
  AND2_X1 U11084 ( .A1(n49089), .A2(n49119), .ZN(n49091) );
  OR2_X1 U11085 ( .A1(n49390), .A2(n2859), .ZN(n49391) );
  OAI21_X1 U11086 ( .B1(n51091), .B2(n49432), .A(n2859), .ZN(n47201) );
  AND2_X1 U11087 ( .A1(n49441), .A2(n49440), .ZN(n3221) );
  NOR3_X1 U11088 ( .A1(n51316), .A2(n49442), .A3(n49432), .ZN(n49459) );
  OR2_X1 U11090 ( .A1(n49574), .A2(n49608), .ZN(n4544) );
  OAI21_X1 U11091 ( .B1(n49600), .B2(n49601), .A(n6814), .ZN(n6813) );
  OR2_X1 U11092 ( .A1(n49604), .A2(n49603), .ZN(n6812) );
  INV_X1 U11093 ( .A(n49770), .ZN(n6249) );
  AND2_X1 U11094 ( .A1(n562), .A2(n50143), .ZN(n2794) );
  NOR2_X1 U11095 ( .A1(n4202), .A2(n50064), .ZN(n50063) );
  AND2_X1 U11097 ( .A1(n50193), .A2(n50195), .ZN(n5797) );
  AND3_X1 U11098 ( .A1(n5224), .A2(n50398), .A3(n50410), .ZN(n5222) );
  OR2_X1 U11099 ( .A1(n50457), .A2(n50412), .ZN(n5224) );
  AND2_X1 U11100 ( .A1(n50480), .A2(n50481), .ZN(n8244) );
  OR2_X1 U11101 ( .A1(n50473), .A2(n50457), .ZN(n8243) );
  INV_X1 U11102 ( .A(n50533), .ZN(n50554) );
  INV_X1 U11103 ( .A(n50550), .ZN(n50520) );
  INV_X1 U11104 ( .A(n50521), .ZN(n6665) );
  OAI21_X1 U11105 ( .B1(n46967), .B2(n49994), .A(n7883), .ZN(n7882) );
  AND2_X1 U11106 ( .A1(n5849), .A2(n5850), .ZN(n5847) );
  AND3_X1 U11107 ( .A1(n44111), .A2(n7452), .A3(n46778), .ZN(n5742) );
  INV_X1 U11108 ( .A(n50679), .ZN(n2564) );
  NOR2_X1 U11109 ( .A1(n50678), .A2(n1467), .ZN(n6619) );
  AND2_X1 U11110 ( .A1(n50705), .A2(n50702), .ZN(n4079) );
  NOR2_X1 U11111 ( .A1(n50798), .A2(n2095), .ZN(n4562) );
  AND2_X1 U11112 ( .A1(n50751), .A2(n50787), .ZN(n4830) );
  OR2_X1 U11113 ( .A1(n52097), .A2(n50890), .ZN(n6818) );
  AOI22_X1 U11114 ( .A1(n50820), .A2(n50880), .B1(n50870), .B2(n52093), .ZN(
        n50824) );
  INV_X1 U11115 ( .A(n50831), .ZN(n50887) );
  OR2_X1 U11116 ( .A1(n50864), .A2(n50847), .ZN(n50897) );
  OR2_X1 U11117 ( .A1(n2731), .A2(n2732), .ZN(n2730) );
  INV_X1 U11118 ( .A(n50901), .ZN(n50916) );
  NOR2_X1 U11119 ( .A1(n50911), .A2(n2864), .ZN(n2863) );
  OAI21_X1 U11120 ( .B1(n7324), .B2(n7323), .A(n50934), .ZN(n47395) );
  AOI21_X1 U11121 ( .B1(n3547), .B2(n49804), .A(n3548), .ZN(n3543) );
  INV_X1 U11122 ( .A(n4515), .ZN(n6229) );
  NOR2_X1 U11123 ( .A1(n5992), .A2(n47521), .ZN(n4055) );
  OAI211_X1 U11124 ( .C1(n47805), .C2(n47804), .A(n47810), .B(n47811), .ZN(
        n47813) );
  AND2_X1 U11125 ( .A1(n3957), .A2(n47997), .ZN(n3956) );
  AND2_X1 U11126 ( .A1(n6354), .A2(n48052), .ZN(n48063) );
  NAND4_X1 U11127 ( .A1(n48163), .A2(n3909), .A3(n3990), .A4(n3908), .ZN(n3910) );
  OAI21_X1 U11128 ( .B1(n48327), .B2(n8104), .A(n51728), .ZN(n48337) );
  AND2_X1 U11129 ( .A1(n48608), .A2(n48609), .ZN(n6805) );
  AOI22_X1 U11130 ( .A1(n7676), .A2(n7674), .B1(n7670), .B2(n34420), .ZN(n7669) );
  AND2_X1 U11131 ( .A1(n8167), .A2(n8165), .ZN(n8163) );
  OAI21_X1 U11132 ( .B1(n48873), .B2(n48872), .A(n48881), .ZN(n5886) );
  INV_X1 U11133 ( .A(n4423), .ZN(n3793) );
  AND2_X1 U11134 ( .A1(n50447), .A2(n50460), .ZN(n4690) );
  OAI211_X1 U11135 ( .C1(n50456), .C2(n50476), .A(n7113), .B(n7112), .ZN(
        n50462) );
  NAND2_X1 U11136 ( .A1(n7748), .A2(n7747), .ZN(n7737) );
  AND2_X1 U11137 ( .A1(n50960), .A2(n50962), .ZN(n4504) );
  INV_X1 U11138 ( .A(n51052), .ZN(n40032) );
  INV_X1 U11139 ( .A(n21873), .ZN(n23303) );
  INV_X1 U11140 ( .A(n29191), .ZN(n5656) );
  INV_X1 U11141 ( .A(n36141), .ZN(n3817) );
  INV_X1 U11143 ( .A(n39299), .ZN(n5593) );
  INV_X1 U11144 ( .A(n11629), .ZN(n3024) );
  INV_X1 U11146 ( .A(n12612), .ZN(n3377) );
  XNOR2_X1 U11147 ( .A(n18185), .B(n18184), .ZN(n21304) );
  INV_X1 U11149 ( .A(n39395), .ZN(n3737) );
  AND4_X1 U11151 ( .A1(n23634), .A2(n23641), .A3(n23958), .A4(n23955), .ZN(
        n2234) );
  INV_X1 U11152 ( .A(n32439), .ZN(n3703) );
  INV_X1 U11153 ( .A(n12278), .ZN(n10724) );
  NAND4_X2 U11155 ( .A1(n5339), .A2(n27675), .A3(n5206), .A4(n5205), .ZN(
        n31096) );
  INV_X1 U11156 ( .A(n31096), .ZN(n5278) );
  INV_X1 U11157 ( .A(n23924), .ZN(n8149) );
  INV_X1 U11158 ( .A(n32478), .ZN(n3664) );
  INV_X1 U11159 ( .A(n13874), .ZN(n8437) );
  INV_X1 U11160 ( .A(n28333), .ZN(n5330) );
  INV_X1 U11161 ( .A(n46196), .ZN(n5783) );
  AND3_X1 U11162 ( .A1(n11260), .A2(n2504), .A3(n10834), .ZN(n2236) );
  INV_X1 U11163 ( .A(n11224), .ZN(n4150) );
  INV_X1 U11166 ( .A(n28143), .ZN(n7602) );
  AND2_X1 U11167 ( .A1(n29998), .A2(n30983), .ZN(n2237) );
  AND2_X1 U11168 ( .A1(n11993), .A2(n15341), .ZN(n2238) );
  AND4_X1 U11169 ( .A1(n19820), .A2(n21197), .A3(n19819), .A4(n21208), .ZN(
        n2239) );
  AND3_X1 U11170 ( .A1(n27800), .A2(n6058), .A3(n51747), .ZN(n2240) );
  OR2_X1 U11171 ( .A1(n15134), .A2(n15138), .ZN(n2241) );
  AND2_X1 U11172 ( .A1(n42994), .A2(n7797), .ZN(n2242) );
  OR2_X1 U11173 ( .A1(n37751), .A2(n3650), .ZN(n2243) );
  AND2_X1 U11174 ( .A1(n3270), .A2(n3269), .ZN(n2244) );
  AND2_X1 U11175 ( .A1(n36305), .A2(n38549), .ZN(n2245) );
  OR2_X1 U11176 ( .A1(n18906), .A2(n19640), .ZN(n2246) );
  AND2_X1 U11177 ( .A1(n29270), .A2(n29185), .ZN(n2247) );
  AND2_X1 U11178 ( .A1(n40652), .A2(n41446), .ZN(n2248) );
  INV_X1 U11179 ( .A(n11354), .ZN(n9369) );
  INV_X1 U11180 ( .A(n42181), .ZN(n42176) );
  INV_X1 U11182 ( .A(n34649), .ZN(n36430) );
  XOR2_X1 U11183 ( .A(n4627), .B(n4487), .Z(n2250) );
  AND2_X1 U11184 ( .A1(n4130), .A2(n4127), .ZN(n2251) );
  AND2_X1 U11185 ( .A1(n47076), .A2(n7046), .ZN(n2252) );
  AND2_X1 U11186 ( .A1(n640), .A2(n14453), .ZN(n2253) );
  INV_X1 U11187 ( .A(n24452), .ZN(n22702) );
  INV_X1 U11188 ( .A(n26905), .ZN(n7362) );
  INV_X1 U11189 ( .A(n30180), .ZN(n30182) );
  XOR2_X1 U11191 ( .A(n15627), .B(n16079), .Z(n2254) );
  INV_X1 U11192 ( .A(n15630), .ZN(n7259) );
  INV_X1 U11193 ( .A(n19336), .ZN(n20515) );
  INV_X1 U11194 ( .A(n21530), .ZN(n21513) );
  INV_X1 U11195 ( .A(n20422), .ZN(n6452) );
  INV_X1 U11196 ( .A(n11410), .ZN(n11423) );
  INV_X1 U11197 ( .A(n29686), .ZN(n6013) );
  INV_X1 U11198 ( .A(n21389), .ZN(n5923) );
  INV_X1 U11199 ( .A(n41150), .ZN(n7977) );
  INV_X1 U11200 ( .A(n31683), .ZN(n7598) );
  INV_X1 U11201 ( .A(n7616), .ZN(n50008) );
  INV_X1 U11202 ( .A(n37721), .ZN(n36901) );
  INV_X1 U11203 ( .A(n31538), .ZN(n5867) );
  INV_X1 U11204 ( .A(n2176), .ZN(n37805) );
  INV_X1 U11205 ( .A(n48140), .ZN(n8689) );
  INV_X1 U11206 ( .A(n32402), .ZN(n5665) );
  INV_X1 U11208 ( .A(n39273), .ZN(n36781) );
  INV_X1 U11210 ( .A(n38701), .ZN(n37911) );
  INV_X1 U11211 ( .A(n23142), .ZN(n3907) );
  INV_X1 U11212 ( .A(n41650), .ZN(n6938) );
  INV_X1 U11213 ( .A(n31496), .ZN(n3224) );
  INV_X1 U11215 ( .A(n12595), .ZN(n12602) );
  INV_X1 U11216 ( .A(n46880), .ZN(n7449) );
  INV_X1 U11218 ( .A(n27670), .ZN(n8290) );
  INV_X1 U11219 ( .A(n37519), .ZN(n7004) );
  AND2_X1 U11220 ( .A1(n20376), .A2(n5923), .ZN(n2257) );
  XNOR2_X1 U11221 ( .A(n28099), .B(n8405), .ZN(n28860) );
  INV_X1 U11222 ( .A(n28860), .ZN(n28867) );
  INV_X1 U11226 ( .A(n32900), .ZN(n8681) );
  INV_X1 U11227 ( .A(n5656), .ZN(n8422) );
  OR2_X1 U11228 ( .A1(n23487), .A2(n23486), .ZN(n2258) );
  AND4_X1 U11229 ( .A1(n3878), .A2(n3879), .A3(n3881), .A4(n3880), .ZN(n2259)
         );
  INV_X1 U11230 ( .A(n39184), .ZN(n7729) );
  XNOR2_X1 U11231 ( .A(n5717), .B(n37093), .ZN(n39184) );
  INV_X1 U11232 ( .A(n46721), .ZN(n7919) );
  INV_X1 U11233 ( .A(n23531), .ZN(n3816) );
  AND2_X1 U11234 ( .A1(n47066), .A2(n47067), .ZN(n2260) );
  AND4_X1 U11235 ( .A1(n12050), .A2(n9227), .A3(n2915), .A4(n2914), .ZN(n2261)
         );
  BUF_X1 U11236 ( .A(n30593), .Z(n30607) );
  INV_X1 U11238 ( .A(n40316), .ZN(n4000) );
  OR2_X1 U11239 ( .A1(n22982), .A2(n22983), .ZN(n2262) );
  XOR2_X1 U11240 ( .A(n52180), .B(n18821), .Z(n2263) );
  INV_X1 U11242 ( .A(n50708), .ZN(n7459) );
  OR2_X1 U11243 ( .A1(n23955), .A2(n5069), .ZN(n5068) );
  INV_X1 U11244 ( .A(n30592), .ZN(n30598) );
  XNOR2_X1 U11245 ( .A(n24466), .B(n28121), .ZN(n28297) );
  INV_X1 U11246 ( .A(n29488), .ZN(n26671) );
  AND2_X1 U11247 ( .A1(n23030), .A2(n19317), .ZN(n2264) );
  INV_X1 U11248 ( .A(n21652), .ZN(n6721) );
  XOR2_X1 U11249 ( .A(n18605), .B(n18604), .Z(n2265) );
  AND4_X1 U11250 ( .A1(n45656), .A2(n49181), .A3(n45217), .A4(n3229), .ZN(
        n2266) );
  AND3_X1 U11251 ( .A1(n42365), .A2(n46204), .A3(n666), .ZN(n2267) );
  AND2_X1 U11252 ( .A1(n3852), .A2(n48198), .ZN(n2268) );
  AND3_X1 U11253 ( .A1(n10439), .A2(n11941), .A3(n11957), .ZN(n2269) );
  INV_X1 U11254 ( .A(n14294), .ZN(n8397) );
  AND3_X1 U11255 ( .A1(n6259), .A2(n6258), .A3(n2554), .ZN(n2270) );
  AND3_X1 U11256 ( .A1(n19067), .A2(n7038), .A3(n7037), .ZN(n2271) );
  AND3_X1 U11257 ( .A1(n38178), .A2(n38179), .A3(n7903), .ZN(n2272) );
  AND2_X1 U11258 ( .A1(n22272), .A2(n7789), .ZN(n2273) );
  INV_X1 U11259 ( .A(n41082), .ZN(n2888) );
  XOR2_X1 U11261 ( .A(n18660), .B(n18397), .Z(n2275) );
  XNOR2_X1 U11262 ( .A(n16236), .B(n16235), .ZN(n18962) );
  INV_X1 U11263 ( .A(n18962), .ZN(n21252) );
  AND3_X1 U11264 ( .A1(n8780), .A2(n9028), .A3(n8779), .ZN(n2276) );
  INV_X1 U11265 ( .A(n39754), .ZN(n39942) );
  XOR2_X1 U11266 ( .A(n36832), .B(n36833), .Z(n2277) );
  INV_X1 U11267 ( .A(n48156), .ZN(n8061) );
  NAND2_X1 U11268 ( .A1(n25479), .A2(n29182), .ZN(n29272) );
  XOR2_X1 U11269 ( .A(n42222), .B(n40642), .Z(n2278) );
  OR2_X1 U11270 ( .A1(n22674), .A2(n51021), .ZN(n2279) );
  AND2_X1 U11271 ( .A1(n50321), .A2(n49994), .ZN(n2280) );
  INV_X1 U11272 ( .A(n10686), .ZN(n6786) );
  XNOR2_X1 U11273 ( .A(n25512), .B(n25511), .ZN(n28708) );
  AND3_X1 U11274 ( .A1(n3010), .A2(n31258), .A3(n32425), .ZN(n2281) );
  AND2_X1 U11275 ( .A1(n14063), .A2(n14062), .ZN(n2282) );
  INV_X1 U11276 ( .A(n39944), .ZN(n38838) );
  INV_X1 U11278 ( .A(n37406), .ZN(n5784) );
  XNOR2_X1 U11279 ( .A(n9242), .B(Key[31]), .ZN(n10398) );
  NOR2_X1 U11280 ( .A1(n31911), .A2(n31075), .ZN(n32844) );
  XOR2_X1 U11281 ( .A(n44504), .B(n44503), .Z(n2284) );
  AND2_X1 U11282 ( .A1(n11393), .A2(n9221), .ZN(n2285) );
  INV_X1 U11283 ( .A(n30854), .ZN(n31631) );
  AND2_X1 U11284 ( .A1(n47090), .A2(n2574), .ZN(n2286) );
  INV_X1 U11285 ( .A(n20660), .ZN(n3344) );
  AND3_X1 U11286 ( .A1(n8828), .A2(n8831), .A3(n8829), .ZN(n2287) );
  XNOR2_X1 U11287 ( .A(n43722), .B(n8669), .ZN(n43797) );
  INV_X1 U11288 ( .A(n667), .ZN(n3607) );
  XOR2_X1 U11289 ( .A(n27496), .B(n27495), .Z(n2288) );
  INV_X1 U11290 ( .A(n38937), .ZN(n5151) );
  AND2_X1 U11291 ( .A1(n3484), .A2(n31014), .ZN(n2289) );
  XOR2_X1 U11292 ( .A(n18659), .B(n2181), .Z(n2290) );
  INV_X1 U11293 ( .A(n20649), .ZN(n3370) );
  INV_X1 U11294 ( .A(n39576), .ZN(n41013) );
  XNOR2_X1 U11295 ( .A(n29983), .B(n29982), .ZN(n38543) );
  XOR2_X1 U11296 ( .A(n25084), .B(n23852), .Z(n2291) );
  INV_X1 U11297 ( .A(n36550), .ZN(n8016) );
  AND3_X1 U11298 ( .A1(n19918), .A2(n19919), .A3(n3871), .ZN(n2292) );
  INV_X1 U11299 ( .A(n12617), .ZN(n12069) );
  INV_X1 U11300 ( .A(n2222), .ZN(n19427) );
  XOR2_X1 U11301 ( .A(n25485), .B(n25604), .Z(n2293) );
  INV_X1 U11302 ( .A(n37740), .ZN(n3738) );
  XNOR2_X1 U11303 ( .A(n43709), .B(n45047), .ZN(n6811) );
  OR2_X1 U11304 ( .A1(n29514), .A2(n29508), .ZN(n2295) );
  XOR2_X1 U11305 ( .A(n51502), .B(n24817), .Z(n2296) );
  XNOR2_X1 U11306 ( .A(n25263), .B(n5663), .ZN(n27132) );
  AND2_X1 U11307 ( .A1(n46028), .A2(n49656), .ZN(n2297) );
  INV_X1 U11308 ( .A(n21303), .ZN(n18217) );
  INV_X1 U11309 ( .A(n591), .ZN(n7759) );
  XOR2_X1 U11310 ( .A(n16330), .B(n16746), .Z(n2298) );
  XNOR2_X1 U11311 ( .A(n8821), .B(Key[42]), .ZN(n10162) );
  OR2_X1 U11312 ( .A1(n19705), .A2(n18976), .ZN(n2299) );
  INV_X1 U11315 ( .A(n48944), .ZN(n47476) );
  INV_X1 U11316 ( .A(n31558), .ZN(n32620) );
  XNOR2_X1 U11319 ( .A(n23853), .B(n2291), .ZN(n23861) );
  INV_X1 U11320 ( .A(n23861), .ZN(n3819) );
  XOR2_X1 U11321 ( .A(n45368), .B(n43118), .Z(n2301) );
  XOR2_X1 U11323 ( .A(n14112), .B(n15682), .Z(n2302) );
  XOR2_X1 U11324 ( .A(n44984), .B(n44983), .Z(n2303) );
  XOR2_X1 U11325 ( .A(n33776), .B(n33775), .Z(n2304) );
  NAND2_X1 U11326 ( .A1(n20474), .A2(n20472), .ZN(n20468) );
  INV_X1 U11327 ( .A(n20468), .ZN(n4098) );
  XOR2_X1 U11328 ( .A(n26377), .B(n25124), .Z(n2305) );
  XNOR2_X1 U11329 ( .A(n24914), .B(n24913), .ZN(n27957) );
  AND2_X1 U11331 ( .A1(n19781), .A2(n19789), .ZN(n2307) );
  INV_X1 U11332 ( .A(n39270), .ZN(n36779) );
  XNOR2_X1 U11333 ( .A(n40765), .B(n40766), .ZN(n44652) );
  INV_X1 U11334 ( .A(n44652), .ZN(n5325) );
  INV_X1 U11336 ( .A(n37130), .ZN(n34069) );
  INV_X1 U11337 ( .A(n34069), .ZN(n3924) );
  OR3_X1 U11338 ( .A1(n48548), .A2(n45372), .A3(n52059), .ZN(n2308) );
  INV_X1 U11339 ( .A(n15631), .ZN(n19893) );
  XOR2_X1 U11340 ( .A(n36808), .B(n33707), .Z(n2309) );
  AND2_X1 U11341 ( .A1(n2999), .A2(n2998), .ZN(n2310) );
  INV_X1 U11342 ( .A(n10096), .ZN(n10530) );
  INV_X1 U11343 ( .A(n41587), .ZN(n3831) );
  XOR2_X1 U11344 ( .A(n33627), .B(n15603), .Z(n2311) );
  XOR2_X1 U11345 ( .A(n27482), .B(n27223), .Z(n2312) );
  XNOR2_X1 U11346 ( .A(n45398), .B(n45397), .ZN(n46336) );
  AND3_X1 U11347 ( .A1(n10293), .A2(n10945), .A3(n12314), .ZN(n2313) );
  INV_X1 U11348 ( .A(n19703), .ZN(n8311) );
  XOR2_X1 U11349 ( .A(n28729), .B(n4275), .Z(n2314) );
  INV_X1 U11350 ( .A(n46435), .ZN(n8585) );
  NAND3_X2 U11351 ( .A1(n5470), .A2(n28326), .A3(n28327), .ZN(n32960) );
  XOR2_X1 U11352 ( .A(n35347), .B(n35346), .Z(n2315) );
  INV_X1 U11353 ( .A(n19636), .ZN(n3033) );
  XOR2_X1 U11354 ( .A(n26127), .B(n26126), .Z(n2316) );
  XOR2_X1 U11355 ( .A(n16506), .B(n16505), .Z(n2317) );
  XOR2_X1 U11356 ( .A(n17850), .B(n17849), .Z(n2318) );
  XOR2_X1 U11357 ( .A(n24839), .B(n24838), .Z(n2319) );
  XOR2_X1 U11358 ( .A(n24440), .B(n24439), .Z(n2320) );
  AND3_X1 U11359 ( .A1(n30054), .A2(n30053), .A3(n31336), .ZN(n2321) );
  INV_X1 U11361 ( .A(n41539), .ZN(n3494) );
  INV_X1 U11362 ( .A(n8909), .ZN(n11500) );
  XOR2_X1 U11363 ( .A(n36858), .B(n34814), .Z(n2322) );
  XOR2_X1 U11364 ( .A(n17925), .B(n15945), .Z(n2323) );
  XNOR2_X1 U11365 ( .A(n2590), .B(n37268), .ZN(n37283) );
  INV_X1 U11366 ( .A(n37283), .ZN(n6343) );
  INV_X1 U11367 ( .A(n31122), .ZN(n31111) );
  INV_X1 U11368 ( .A(n41328), .ZN(n5859) );
  INV_X1 U11369 ( .A(n15386), .ZN(n15382) );
  INV_X1 U11370 ( .A(n11467), .ZN(n11621) );
  AND3_X1 U11371 ( .A1(n51325), .A2(n40120), .A3(n40119), .ZN(n2324) );
  NOR2_X1 U11372 ( .A1(n23112), .A2(n27158), .ZN(n30719) );
  AND3_X1 U11373 ( .A1(n36019), .A2(n36567), .A3(n36560), .ZN(n2325) );
  XOR2_X1 U11374 ( .A(n34632), .B(n37646), .Z(n2326) );
  XOR2_X1 U11375 ( .A(n51057), .B(n444), .Z(n2327) );
  INV_X1 U11376 ( .A(n9406), .ZN(n12125) );
  NAND2_X1 U11377 ( .A1(n30248), .A2(n30244), .ZN(n27145) );
  INV_X1 U11378 ( .A(n27145), .ZN(n5821) );
  XOR2_X1 U11379 ( .A(n18123), .B(n17733), .Z(n2329) );
  INV_X1 U11380 ( .A(n30345), .ZN(n30348) );
  XNOR2_X1 U11381 ( .A(n8562), .B(n24531), .ZN(n29459) );
  INV_X1 U11382 ( .A(n29459), .ZN(n7973) );
  OR3_X1 U11383 ( .A1(n613), .A2(n37619), .A3(n2123), .ZN(n2330) );
  AND2_X1 U11384 ( .A1(n36632), .A2(n695), .ZN(n2331) );
  AND3_X1 U11385 ( .A1(n50890), .A2(n601), .A3(n51312), .ZN(n2332) );
  INV_X1 U11386 ( .A(n31764), .ZN(n31219) );
  INV_X1 U11387 ( .A(n42209), .ZN(n7306) );
  INV_X1 U11388 ( .A(n21714), .ZN(n21713) );
  AND2_X1 U11389 ( .A1(n601), .A2(n50829), .ZN(n2333) );
  INV_X1 U11390 ( .A(n14139), .ZN(n14783) );
  INV_X1 U11391 ( .A(n47477), .ZN(n3209) );
  AND2_X1 U11392 ( .A1(n31746), .A2(n32303), .ZN(n2334) );
  INV_X1 U11393 ( .A(n12600), .ZN(n3692) );
  AND3_X1 U11394 ( .A1(n2220), .A2(n21495), .A3(n20441), .ZN(n2335) );
  AND3_X1 U11395 ( .A1(n44876), .A2(n44875), .A3(n44874), .ZN(n2336) );
  AND2_X1 U11396 ( .A1(n28508), .A2(n28862), .ZN(n2337) );
  INV_X1 U11397 ( .A(n30256), .ZN(n6486) );
  NOR2_X1 U11398 ( .A1(n10240), .A2(n10199), .ZN(n10244) );
  AND2_X1 U11399 ( .A1(n20840), .A2(n20322), .ZN(n4433) );
  XNOR2_X1 U11400 ( .A(n24813), .B(n24812), .ZN(n2338) );
  XOR2_X1 U11401 ( .A(n18619), .B(n18198), .Z(n2339) );
  OR2_X1 U11402 ( .A1(n39464), .A2(n7815), .ZN(n2340) );
  AND2_X1 U11403 ( .A1(n46475), .A2(n52203), .ZN(n2341) );
  INV_X1 U11404 ( .A(n50913), .ZN(n5365) );
  AND2_X1 U11405 ( .A1(n39236), .A2(n51063), .ZN(n2342) );
  XOR2_X1 U11406 ( .A(n51472), .B(n35790), .Z(n2343) );
  NOR2_X1 U11407 ( .A1(n51400), .A2(n46668), .ZN(n8449) );
  AND3_X1 U11408 ( .A1(n43328), .A2(n40801), .A3(n38763), .ZN(n2344) );
  INV_X1 U11409 ( .A(n45164), .ZN(n2751) );
  INV_X1 U11411 ( .A(n37962), .ZN(n3626) );
  OR2_X1 U11412 ( .A1(n48264), .A2(n6674), .ZN(n2346) );
  AND2_X1 U11413 ( .A1(n12344), .A2(n12340), .ZN(n2347) );
  AND4_X1 U11414 ( .A1(n12338), .A2(n12339), .A3(n12337), .A4(n12336), .ZN(
        n2348) );
  AND3_X1 U11415 ( .A1(n723), .A2(n3703), .A3(n32438), .ZN(n2349) );
  AND2_X1 U11416 ( .A1(n46029), .A2(n50020), .ZN(n2350) );
  OAI21_X1 U11417 ( .B1(n6249), .B2(n6248), .A(n49854), .ZN(n49842) );
  AND2_X1 U11418 ( .A1(n21630), .A2(n21639), .ZN(n2351) );
  AND2_X1 U11419 ( .A1(n22859), .A2(n22857), .ZN(n2352) );
  INV_X1 U11420 ( .A(n11635), .ZN(n11477) );
  AND2_X1 U11422 ( .A1(n27784), .A2(n28715), .ZN(n2353) );
  AND2_X1 U11423 ( .A1(n30034), .A2(n31333), .ZN(n2354) );
  XOR2_X1 U11424 ( .A(n18464), .B(n16559), .Z(n2355) );
  AND3_X1 U11425 ( .A1(n41153), .A2(n41152), .A3(n1931), .ZN(n2356) );
  OR2_X1 U11426 ( .A1(n37773), .A2(n37781), .ZN(n2357) );
  XNOR2_X1 U11427 ( .A(n33829), .B(n33828), .ZN(n33870) );
  INV_X1 U11428 ( .A(n33870), .ZN(n7159) );
  AND3_X1 U11429 ( .A1(n14652), .A2(n12785), .A3(n12794), .ZN(n2358) );
  OR2_X1 U11430 ( .A1(n32464), .A2(n2853), .ZN(n2359) );
  AND2_X1 U11431 ( .A1(n40014), .A2(n6961), .ZN(n2360) );
  AND2_X1 U11432 ( .A1(n14542), .A2(n14545), .ZN(n2361) );
  AND2_X1 U11433 ( .A1(n34806), .A2(n39450), .ZN(n2362) );
  AND3_X1 U11434 ( .A1(n5919), .A2(n41202), .A3(n41212), .ZN(n2363) );
  AND2_X1 U11435 ( .A1(n37561), .A2(n7011), .ZN(n2364) );
  AND2_X1 U11436 ( .A1(n31347), .A2(n31346), .ZN(n2365) );
  INV_X1 U11437 ( .A(n6515), .ZN(n20032) );
  OR2_X1 U11439 ( .A1(n31892), .A2(n31425), .ZN(n2366) );
  AND2_X1 U11440 ( .A1(n30690), .A2(n29940), .ZN(n2367) );
  OR2_X1 U11441 ( .A1(n20826), .A2(n2220), .ZN(n2368) );
  AND2_X1 U11442 ( .A1(n36461), .A2(n36045), .ZN(n2369) );
  INV_X1 U11443 ( .A(n12068), .ZN(n3347) );
  AND3_X1 U11444 ( .A1(n10570), .A2(n10565), .A3(n10572), .ZN(n2370) );
  XOR2_X1 U11445 ( .A(n43561), .B(n43830), .Z(n2371) );
  INV_X1 U11446 ( .A(n21945), .ZN(n6010) );
  AND3_X1 U11447 ( .A1(n37393), .A2(n37517), .A3(n5730), .ZN(n2372) );
  OR2_X1 U11448 ( .A1(n29893), .A2(n30785), .ZN(n2373) );
  INV_X1 U11449 ( .A(n49579), .ZN(n6985) );
  AND2_X1 U11450 ( .A1(n21434), .A2(n21431), .ZN(n2374) );
  XOR2_X1 U11451 ( .A(n17965), .B(n34495), .Z(n2375) );
  INV_X1 U11452 ( .A(n38317), .ZN(n6748) );
  AND2_X1 U11453 ( .A1(n23635), .A2(n23090), .ZN(n2376) );
  XOR2_X1 U11454 ( .A(n38005), .B(n35028), .Z(n2377) );
  AND2_X1 U11455 ( .A1(n12134), .A2(n11411), .ZN(n2378) );
  OR2_X1 U11456 ( .A1(n3597), .A2(n41328), .ZN(n2379) );
  AND2_X1 U11458 ( .A1(n8463), .A2(n15442), .ZN(n2380) );
  NAND2_X1 U11459 ( .A1(n21276), .A2(n19452), .ZN(n19455) );
  INV_X1 U11460 ( .A(n51755), .ZN(n5167) );
  INV_X1 U11461 ( .A(n21414), .ZN(n5192) );
  AND2_X1 U11462 ( .A1(n22201), .A2(n3505), .ZN(n2381) );
  AND2_X1 U11463 ( .A1(n51375), .A2(n42154), .ZN(n2382) );
  AND2_X1 U11464 ( .A1(n12699), .A2(n12710), .ZN(n2383) );
  INV_X1 U11465 ( .A(n15134), .ZN(n5347) );
  XOR2_X1 U11466 ( .A(n32752), .B(n16941), .Z(n2384) );
  OR2_X1 U11467 ( .A1(n32487), .A2(n32486), .ZN(n2385) );
  OR2_X1 U11468 ( .A1(n7449), .A2(n46869), .ZN(n47110) );
  AND2_X1 U11469 ( .A1(n575), .A2(n39955), .ZN(n2386) );
  XOR2_X1 U11470 ( .A(n33267), .B(n33056), .Z(n2387) );
  INV_X1 U11471 ( .A(n23171), .ZN(n3055) );
  INV_X1 U11472 ( .A(n50888), .ZN(n6817) );
  XNOR2_X1 U11473 ( .A(n6291), .B(n7722), .ZN(n6449) );
  AND2_X1 U11474 ( .A1(n32608), .A2(n31569), .ZN(n2388) );
  INV_X1 U11475 ( .A(n31112), .ZN(n7093) );
  INV_X1 U11477 ( .A(n28659), .ZN(n30218) );
  OR2_X1 U11478 ( .A1(n48267), .A2(n44665), .ZN(n2390) );
  AND2_X1 U11479 ( .A1(n20067), .A2(n18303), .ZN(n2391) );
  NOR2_X1 U11480 ( .A1(n12352), .A2(n8724), .ZN(n2392) );
  OR2_X1 U11481 ( .A1(n40468), .A2(n41115), .ZN(n2393) );
  AND2_X1 U11482 ( .A1(n12543), .A2(n442), .ZN(n2394) );
  OR2_X1 U11483 ( .A1(n51140), .A2(n11914), .ZN(n2395) );
  AND2_X1 U11484 ( .A1(n49092), .A2(n49068), .ZN(n2396) );
  OR2_X1 U11485 ( .A1(n48150), .A2(n4501), .ZN(n2397) );
  OR2_X1 U11486 ( .A1(n21452), .A2(n20488), .ZN(n2398) );
  INV_X1 U11487 ( .A(n39103), .ZN(n6740) );
  INV_X1 U11489 ( .A(n50847), .ZN(n5295) );
  OR2_X1 U11490 ( .A1(n26813), .A2(n27580), .ZN(n2400) );
  INV_X1 U11492 ( .A(n24105), .ZN(n4726) );
  OR2_X1 U11493 ( .A1(n30022), .A2(n51240), .ZN(n2402) );
  OR2_X1 U11494 ( .A1(n21470), .A2(n21450), .ZN(n2403) );
  INV_X1 U11495 ( .A(n51747), .ZN(n6059) );
  AND2_X1 U11497 ( .A1(n49291), .A2(n49289), .ZN(n2404) );
  AND2_X1 U11498 ( .A1(n42206), .A2(n37827), .ZN(n2405) );
  AND2_X1 U11499 ( .A1(n12266), .A2(n10748), .ZN(n2406) );
  XOR2_X1 U11500 ( .A(n16504), .B(n16503), .Z(n2407) );
  AND2_X1 U11501 ( .A1(n41211), .A2(n41202), .ZN(n2408) );
  AND2_X1 U11502 ( .A1(n27686), .A2(n27685), .ZN(n2409) );
  XOR2_X1 U11503 ( .A(n35841), .B(n36681), .Z(n2410) );
  OR2_X1 U11504 ( .A1(n9515), .A2(n9305), .ZN(n2411) );
  XOR2_X1 U11505 ( .A(n25946), .B(n24399), .Z(n2412) );
  AND2_X1 U11506 ( .A1(n41013), .A2(n51358), .ZN(n2413) );
  OR2_X1 U11507 ( .A1(n19399), .A2(n19396), .ZN(n2414) );
  AND2_X1 U11508 ( .A1(n47505), .A2(n51346), .ZN(n2415) );
  INV_X1 U11509 ( .A(n47309), .ZN(n47012) );
  AND2_X1 U11510 ( .A1(n46435), .A2(n51732), .ZN(n2416) );
  AND2_X1 U11511 ( .A1(n30065), .A2(n30066), .ZN(n2417) );
  AND3_X1 U11512 ( .A1(n32759), .A2(n32760), .A3(n32761), .ZN(n2418) );
  AND2_X1 U11513 ( .A1(n19659), .A2(n19658), .ZN(n2419) );
  AND2_X1 U11514 ( .A1(n29424), .A2(n26998), .ZN(n2420) );
  AND3_X1 U11515 ( .A1(n38629), .A2(n3947), .A3(n3946), .ZN(n2421) );
  AND2_X1 U11516 ( .A1(n46799), .A2(n46798), .ZN(n2422) );
  AND2_X1 U11517 ( .A1(n19176), .A2(n19175), .ZN(n2423) );
  AND2_X1 U11518 ( .A1(n26905), .A2(n26998), .ZN(n2424) );
  INV_X1 U11519 ( .A(n29905), .ZN(n29908) );
  OR2_X1 U11520 ( .A1(n12834), .A2(n11315), .ZN(n13620) );
  OR2_X1 U11521 ( .A1(n40147), .A2(n4950), .ZN(n2425) );
  AND2_X1 U11522 ( .A1(n20119), .A2(n19056), .ZN(n2426) );
  AND2_X1 U11523 ( .A1(n50369), .A2(n50370), .ZN(n2427) );
  AND2_X1 U11524 ( .A1(n3455), .A2(n3453), .ZN(n2428) );
  XOR2_X1 U11525 ( .A(n17160), .B(n17159), .Z(n2429) );
  OR2_X1 U11526 ( .A1(n26732), .A2(n2115), .ZN(n2430) );
  XOR2_X1 U11527 ( .A(n36973), .B(n36972), .Z(n2431) );
  NAND2_X1 U11528 ( .A1(n32787), .A2(n32788), .ZN(n2432) );
  AND2_X1 U11529 ( .A1(n39451), .A2(n36255), .ZN(n2433) );
  AND2_X1 U11530 ( .A1(n32481), .A2(n3664), .ZN(n2434) );
  OR2_X1 U11531 ( .A1(n4975), .A2(n12060), .ZN(n2435) );
  NOR2_X1 U11532 ( .A1(n38722), .A2(n38728), .ZN(n2436) );
  AND2_X1 U11533 ( .A1(n11342), .A2(n11335), .ZN(n2437) );
  OR2_X1 U11534 ( .A1(n30698), .A2(n30699), .ZN(n2438) );
  AND2_X1 U11535 ( .A1(n52137), .A2(n48968), .ZN(n2439) );
  AND2_X1 U11536 ( .A1(n49807), .A2(n49863), .ZN(n2440) );
  OR2_X1 U11537 ( .A1(n34639), .A2(n37640), .ZN(n2441) );
  AND2_X1 U11538 ( .A1(n29484), .A2(n25844), .ZN(n2442) );
  OR2_X1 U11539 ( .A1(n36576), .A2(n458), .ZN(n2443) );
  AND2_X1 U11540 ( .A1(n21519), .A2(n3345), .ZN(n2444) );
  OR2_X1 U11541 ( .A1(n44583), .A2(n50277), .ZN(n2445) );
  AND2_X1 U11542 ( .A1(n50492), .A2(n5483), .ZN(n2446) );
  INV_X1 U11545 ( .A(n24409), .ZN(n24411) );
  OR3_X2 U11546 ( .A1(n2824), .A2(n2826), .A3(n46278), .ZN(n49021) );
  OR2_X1 U11547 ( .A1(n48403), .A2(n48404), .ZN(n2447) );
  AND2_X1 U11548 ( .A1(n27671), .A2(n2642), .ZN(n2448) );
  AND2_X1 U11549 ( .A1(n32551), .A2(n32549), .ZN(n2449) );
  AND3_X1 U11550 ( .A1(n31422), .A2(n31893), .A3(n29992), .ZN(n2450) );
  OR3_X1 U11551 ( .A1(n47792), .A2(n45877), .A3(n45876), .ZN(n2451) );
  NAND2_X1 U11552 ( .A1(n10598), .A2(n10597), .ZN(n2452) );
  AND2_X1 U11553 ( .A1(n21190), .A2(n21191), .ZN(n2453) );
  OR2_X1 U11554 ( .A1(n10981), .A2(n10982), .ZN(n2454) );
  AND2_X1 U11555 ( .A1(n10194), .A2(n10195), .ZN(n2455) );
  AND2_X1 U11556 ( .A1(n21197), .A2(n21208), .ZN(n2456) );
  AND3_X1 U11557 ( .A1(n20984), .A2(n23511), .A3(n21085), .ZN(n2457) );
  AND2_X1 U11558 ( .A1(n28660), .A2(n6220), .ZN(n2458) );
  OR2_X1 U11559 ( .A1(n46189), .A2(n45661), .ZN(n2459) );
  INV_X1 U11560 ( .A(n29447), .ZN(n27040) );
  NAND2_X1 U11561 ( .A1(n49126), .A2(n49117), .ZN(n2460) );
  AND2_X1 U11562 ( .A1(n47126), .A2(n3892), .ZN(n2461) );
  XOR2_X1 U11563 ( .A(n31340), .B(n31338), .Z(n2462) );
  OR2_X1 U11564 ( .A1(n37387), .A2(n38494), .ZN(n2463) );
  INV_X1 U11565 ( .A(n30531), .ZN(n3242) );
  INV_X1 U11566 ( .A(n31452), .ZN(n5868) );
  AND2_X1 U11567 ( .A1(n47151), .A2(n46890), .ZN(n2464) );
  AND2_X1 U11568 ( .A1(n39467), .A2(n39438), .ZN(n2465) );
  INV_X1 U11569 ( .A(n41690), .ZN(n2867) );
  AND3_X1 U11570 ( .A1(n24687), .A2(n30670), .A3(n26909), .ZN(n2466) );
  AND2_X1 U11571 ( .A1(n46715), .A2(n51317), .ZN(n2467) );
  NAND2_X1 U11572 ( .A1(n10060), .A2(n5328), .ZN(n2468) );
  INV_X1 U11573 ( .A(n30245), .ZN(n5169) );
  OR2_X1 U11574 ( .A1(n46838), .A2(n2992), .ZN(n2469) );
  INV_X1 U11575 ( .A(n41938), .ZN(n41927) );
  INV_X1 U11576 ( .A(n8988), .ZN(n10741) );
  AND2_X1 U11577 ( .A1(n3254), .A2(n2114), .ZN(n2470) );
  INV_X1 U11578 ( .A(n41238), .ZN(n6335) );
  AND2_X1 U11579 ( .A1(n5630), .A2(n13764), .ZN(n2471) );
  OR2_X1 U11580 ( .A1(n36430), .A2(n51015), .ZN(n2472) );
  INV_X1 U11582 ( .A(n35953), .ZN(n37386) );
  NOR2_X1 U11583 ( .A1(n32761), .A2(n32765), .ZN(n2473) );
  AND2_X1 U11584 ( .A1(n38659), .A2(n37928), .ZN(n2474) );
  AND2_X1 U11585 ( .A1(n19663), .A2(n51127), .ZN(n2475) );
  NAND2_X1 U11586 ( .A1(n22140), .A2(n22157), .ZN(n2476) );
  NAND3_X1 U11587 ( .A1(n3275), .A2(n7910), .A3(n3274), .ZN(n2477) );
  AND2_X1 U11588 ( .A1(n3640), .A2(n8604), .ZN(n2478) );
  INV_X1 U11589 ( .A(n32966), .ZN(n3303) );
  AND2_X1 U11590 ( .A1(n30694), .A2(n30693), .ZN(n2479) );
  OR2_X1 U11591 ( .A1(n36887), .A2(n39211), .ZN(n2480) );
  OR2_X1 U11592 ( .A1(n22677), .A2(n23184), .ZN(n2481) );
  AND3_X1 U11593 ( .A1(n13814), .A2(n13815), .A3(n13813), .ZN(n2482) );
  OR2_X1 U11594 ( .A1(n32457), .A2(n31648), .ZN(n2483) );
  NAND2_X1 U11595 ( .A1(n26499), .A2(n26498), .ZN(n2484) );
  AND2_X1 U11596 ( .A1(n33026), .A2(n33027), .ZN(n2485) );
  AND2_X1 U11597 ( .A1(n31042), .A2(n5468), .ZN(n2486) );
  INV_X1 U11598 ( .A(n10438), .ZN(n12727) );
  NAND2_X1 U11599 ( .A1(n34529), .A2(n38270), .ZN(n2487) );
  NAND2_X1 U11600 ( .A1(n3637), .A2(n3639), .ZN(n2488) );
  INV_X1 U11601 ( .A(n9547), .ZN(n10474) );
  OR2_X2 U11602 ( .A1(n7988), .A2(n19707), .ZN(n22386) );
  INV_X1 U11603 ( .A(n22386), .ZN(n3270) );
  INV_X1 U11604 ( .A(n38370), .ZN(n40396) );
  OR2_X1 U11605 ( .A1(n49993), .A2(n52143), .ZN(n2489) );
  AND2_X1 U11606 ( .A1(n40862), .A2(n40863), .ZN(n2490) );
  INV_X1 U11607 ( .A(n24292), .ZN(n23510) );
  INV_X1 U11609 ( .A(n13780), .ZN(n13186) );
  OR2_X1 U11610 ( .A1(n38635), .A2(n51360), .ZN(n2491) );
  AND2_X1 U11611 ( .A1(n35978), .A2(n36231), .ZN(n2492) );
  OR2_X1 U11612 ( .A1(n20083), .A2(n20082), .ZN(n2493) );
  INV_X1 U11613 ( .A(n30168), .ZN(n3368) );
  AND2_X1 U11614 ( .A1(n12051), .A2(n799), .ZN(n2494) );
  INV_X1 U11615 ( .A(n40113), .ZN(n7239) );
  NAND3_X1 U11616 ( .A1(n5081), .A2(n48905), .A3(n48900), .ZN(n2495) );
  OR2_X1 U11617 ( .A1(n13873), .A2(n7245), .ZN(n3700) );
  AND2_X1 U11618 ( .A1(n31744), .A2(n435), .ZN(n2496) );
  OR2_X1 U11619 ( .A1(n46908), .A2(n46905), .ZN(n2497) );
  AND2_X1 U11620 ( .A1(n21888), .A2(n22856), .ZN(n2498) );
  AND2_X1 U11621 ( .A1(n29794), .A2(n2707), .ZN(n2499) );
  OR2_X1 U11622 ( .A1(n19851), .A2(n19647), .ZN(n2500) );
  XNOR2_X1 U11623 ( .A(n7079), .B(n9450), .ZN(n2501) );
  AND2_X1 U11624 ( .A1(n30805), .A2(n30799), .ZN(n2502) );
  OR2_X1 U11625 ( .A1(n11036), .A2(n11035), .ZN(n2503) );
  OR2_X1 U11626 ( .A1(n12525), .A2(n5180), .ZN(n2504) );
  OR2_X1 U11627 ( .A1(n45957), .A2(n6116), .ZN(n2505) );
  OR2_X1 U11628 ( .A1(n11325), .A2(n11324), .ZN(n2506) );
  AND3_X1 U11629 ( .A1(n39213), .A2(n36887), .A3(n5160), .ZN(n2507) );
  AND2_X1 U11630 ( .A1(n11027), .A2(n11023), .ZN(n2508) );
  OR2_X1 U11631 ( .A1(n32024), .A2(n32025), .ZN(n2509) );
  OR2_X1 U11632 ( .A1(n21880), .A2(n21875), .ZN(n2510) );
  OR2_X1 U11633 ( .A1(n5056), .A2(n2707), .ZN(n2511) );
  OR2_X1 U11634 ( .A1(n2611), .A2(n8481), .ZN(n2512) );
  OR2_X1 U11635 ( .A1(n39262), .A2(n8429), .ZN(n2513) );
  OR2_X1 U11636 ( .A1(n2756), .A2(n35889), .ZN(n2514) );
  XNOR2_X1 U11637 ( .A(n15898), .B(n15897), .ZN(n2515) );
  AND2_X1 U11638 ( .A1(n22721), .A2(n20528), .ZN(n2516) );
  AND2_X1 U11639 ( .A1(n10608), .A2(n9476), .ZN(n2517) );
  OR2_X1 U11640 ( .A1(n41395), .A2(n5216), .ZN(n41534) );
  INV_X1 U11641 ( .A(n41534), .ZN(n3559) );
  OR2_X1 U11642 ( .A1(n29554), .A2(n6339), .ZN(n2518) );
  BUF_X1 U11643 ( .A(n46173), .Z(n49894) );
  AND2_X1 U11644 ( .A1(n24330), .A2(n23373), .ZN(n2519) );
  AND2_X1 U11645 ( .A1(n51112), .A2(n26731), .ZN(n2520) );
  OR2_X1 U11646 ( .A1(n46572), .A2(n46710), .ZN(n2521) );
  INV_X1 U11647 ( .A(n44822), .ZN(n45523) );
  AND2_X1 U11648 ( .A1(n14471), .A2(n13849), .ZN(n2522) );
  AND2_X1 U11649 ( .A1(n5683), .A2(n52048), .ZN(n2523) );
  OR2_X1 U11650 ( .A1(n29288), .A2(n26083), .ZN(n29305) );
  AND2_X1 U11651 ( .A1(n26828), .A2(n30791), .ZN(n2524) );
  AND2_X1 U11652 ( .A1(n18913), .A2(n5342), .ZN(n2525) );
  INV_X1 U11653 ( .A(n2738), .ZN(n40249) );
  AND4_X2 U11654 ( .A1(n35959), .A2(n35956), .A3(n35957), .A4(n35958), .ZN(
        n2738) );
  AND2_X1 U11655 ( .A1(n6355), .A2(n48084), .ZN(n2526) );
  OR2_X1 U11656 ( .A1(n23961), .A2(n23950), .ZN(n2527) );
  INV_X1 U11657 ( .A(n20487), .ZN(n6180) );
  AND2_X1 U11658 ( .A1(n27795), .A2(n26308), .ZN(n2528) );
  INV_X1 U11659 ( .A(n40972), .ZN(n3775) );
  AND2_X1 U11660 ( .A1(n43666), .A2(n41792), .ZN(n2529) );
  OR2_X1 U11661 ( .A1(n31679), .A2(n2094), .ZN(n2530) );
  AND2_X1 U11662 ( .A1(n28865), .A2(n3826), .ZN(n2531) );
  INV_X1 U11664 ( .A(n27629), .ZN(n3282) );
  INV_X1 U11665 ( .A(n41446), .ZN(n39160) );
  AND2_X1 U11666 ( .A1(n45995), .A2(n43464), .ZN(n49711) );
  INV_X1 U11667 ( .A(n49711), .ZN(n6704) );
  INV_X1 U11669 ( .A(n32965), .ZN(n3035) );
  AND2_X1 U11670 ( .A1(n8803), .A2(n10055), .ZN(n9859) );
  INV_X1 U11671 ( .A(n40049), .ZN(n3290) );
  AND2_X1 U11672 ( .A1(n31306), .A2(n31311), .ZN(n30642) );
  OR2_X1 U11674 ( .A1(n35002), .A2(n35001), .ZN(n2532) );
  INV_X1 U11675 ( .A(n22605), .ZN(n24186) );
  INV_X1 U11676 ( .A(n11619), .ZN(n11470) );
  AND2_X1 U11677 ( .A1(n13102), .A2(n12914), .ZN(n3080) );
  AND2_X1 U11678 ( .A1(n10240), .A2(n10199), .ZN(n8781) );
  OR2_X1 U11679 ( .A1(n27856), .A2(n3124), .ZN(n2533) );
  OR2_X1 U11680 ( .A1(n22772), .A2(n7806), .ZN(n2534) );
  INV_X1 U11681 ( .A(n21698), .ZN(n21105) );
  OR2_X1 U11682 ( .A1(n33562), .A2(n38495), .ZN(n37516) );
  OR2_X1 U11683 ( .A1(n9083), .A2(n9278), .ZN(n2535) );
  OR2_X1 U11684 ( .A1(n49718), .A2(n46001), .ZN(n42992) );
  NAND3_X1 U11685 ( .A1(n39225), .A2(n51507), .A3(n38701), .ZN(n2536) );
  OR2_X1 U11686 ( .A1(n29342), .A2(n29341), .ZN(n2537) );
  OR2_X1 U11687 ( .A1(n10040), .A2(n10041), .ZN(n2538) );
  INV_X1 U11688 ( .A(n3685), .ZN(n7874) );
  NAND2_X1 U11689 ( .A1(n1456), .A2(n5177), .ZN(n2539) );
  OR2_X1 U11690 ( .A1(n12601), .A2(n11137), .ZN(n2540) );
  AND2_X1 U11691 ( .A1(n49432), .A2(n47195), .ZN(n49434) );
  XOR2_X1 U11692 ( .A(n27333), .B(n42824), .Z(n2541) );
  XOR2_X1 U11693 ( .A(n40849), .B(n17994), .Z(n2542) );
  XOR2_X1 U11694 ( .A(n26133), .B(n42592), .Z(n2543) );
  XOR2_X1 U11695 ( .A(n24943), .B(n42314), .Z(n2544) );
  XOR2_X1 U11696 ( .A(n45071), .B(n23774), .Z(n2545) );
  XOR2_X1 U11697 ( .A(n40222), .B(n24011), .Z(n2546) );
  XOR2_X1 U11698 ( .A(n35292), .B(n26360), .Z(n2547) );
  XOR2_X1 U11699 ( .A(n35655), .B(n35654), .Z(n2548) );
  XOR2_X1 U11700 ( .A(n35799), .B(n35798), .Z(n2549) );
  XOR2_X1 U11701 ( .A(n37291), .B(n37290), .Z(n2550) );
  XOR2_X1 U11702 ( .A(n43923), .B(n43922), .Z(n2551) );
  XOR2_X1 U11703 ( .A(n41818), .B(n41817), .Z(n2552) );
  INV_X1 U11704 ( .A(Key[189]), .ZN(n3111) );
  INV_X1 U11705 ( .A(n1341), .ZN(n6311) );
  INV_X1 U11706 ( .A(n4885), .ZN(n6327) );
  INV_X1 U11707 ( .A(n2183), .ZN(n6926) );
  NAND2_X1 U11708 ( .A1(n2553), .A2(n10676), .ZN(n5928) );
  INV_X1 U11711 ( .A(n2554), .ZN(n22182) );
  INV_X1 U11712 ( .A(n10959), .ZN(n10122) );
  NAND2_X1 U11713 ( .A1(n3315), .A2(n10125), .ZN(n9795) );
  NAND2_X1 U11714 ( .A1(n21114), .A2(n21113), .ZN(n2555) );
  INV_X1 U11715 ( .A(n2556), .ZN(n10313) );
  AOI21_X1 U11717 ( .B1(n2556), .B2(n14966), .A(n13124), .ZN(n12237) );
  NAND3_X1 U11718 ( .A1(n2659), .A2(n13116), .A3(n2556), .ZN(n13119) );
  XNOR2_X1 U11719 ( .A(n39955), .B(n38838), .ZN(n36470) );
  NAND2_X1 U11720 ( .A1(n34922), .A2(n34923), .ZN(n36435) );
  NOR2_X1 U11721 ( .A1(n36434), .A2(n36433), .ZN(n2557) );
  NOR2_X1 U11722 ( .A1(n18006), .A2(n2560), .ZN(n2559) );
  NAND2_X1 U11723 ( .A1(n20384), .A2(n20476), .ZN(n19385) );
  NAND2_X1 U11724 ( .A1(n20384), .A2(n2559), .ZN(n2558) );
  NAND2_X1 U11725 ( .A1(n2563), .A2(n18001), .ZN(n2562) );
  AND2_X1 U11726 ( .A1(n18000), .A2(n18003), .ZN(n2563) );
  NAND2_X1 U11728 ( .A1(n52083), .A2(n51012), .ZN(n39842) );
  NAND2_X1 U11730 ( .A1(n2564), .A2(n50708), .ZN(n50689) );
  NAND2_X1 U11731 ( .A1(n44590), .A2(n50251), .ZN(n2565) );
  NAND2_X1 U11732 ( .A1(n44592), .A2(n50277), .ZN(n2566) );
  NAND2_X1 U11733 ( .A1(n44584), .A2(n44585), .ZN(n2567) );
  NAND2_X1 U11734 ( .A1(n27140), .A2(n27995), .ZN(n28908) );
  NAND2_X1 U11735 ( .A1(n28897), .A2(n28588), .ZN(n2568) );
  OR2_X1 U11736 ( .A1(n27131), .A2(n27132), .ZN(n27139) );
  NOR2_X1 U11737 ( .A1(n40990), .A2(n2569), .ZN(n41556) );
  INV_X1 U11738 ( .A(n40932), .ZN(n2569) );
  NAND2_X1 U11739 ( .A1(n2570), .A2(n2571), .ZN(n39277) );
  NAND3_X1 U11740 ( .A1(n39013), .A2(n2571), .A3(n39274), .ZN(n38691) );
  NAND3_X1 U11741 ( .A1(n39286), .A2(n39015), .A3(n2571), .ZN(n39023) );
  NAND2_X1 U11743 ( .A1(n2572), .A2(n19884), .ZN(n15633) );
  NAND2_X1 U11744 ( .A1(n19886), .A2(n19636), .ZN(n2572) );
  OAI211_X1 U11745 ( .C1(n18930), .C2(n2573), .A(n18928), .B(n18929), .ZN(
        n18931) );
  INV_X1 U11746 ( .A(n19886), .ZN(n2573) );
  INV_X1 U11747 ( .A(n47111), .ZN(n2576) );
  NAND2_X1 U11748 ( .A1(n47109), .A2(n47111), .ZN(n2577) );
  INV_X1 U11749 ( .A(n2577), .ZN(n46569) );
  NAND2_X1 U11750 ( .A1(n47109), .A2(n2575), .ZN(n2574) );
  NAND3_X1 U11751 ( .A1(n2577), .A2(n7449), .A3(n47104), .ZN(n45141) );
  AOI22_X1 U11752 ( .A1(n46883), .A2(n2577), .B1(n46882), .B2(n46881), .ZN(
        n46884) );
  XNOR2_X1 U11753 ( .A(n15608), .B(n8233), .ZN(n2578) );
  AOI21_X1 U11754 ( .B1(n12708), .B2(n12712), .A(n2383), .ZN(n2582) );
  INV_X1 U11755 ( .A(n12700), .ZN(n2584) );
  NOR2_X1 U11756 ( .A1(n2588), .A2(n2587), .ZN(n2586) );
  OAI21_X1 U11757 ( .B1(n12708), .B2(n12709), .A(n12707), .ZN(n2587) );
  NOR2_X1 U11758 ( .A1(n1782), .A2(n12701), .ZN(n2588) );
  XNOR2_X1 U11759 ( .A(n37250), .B(n2591), .ZN(n2590) );
  INV_X1 U11760 ( .A(n37251), .ZN(n2591) );
  INV_X1 U11761 ( .A(n32425), .ZN(n2593) );
  NAND3_X2 U11762 ( .A1(n2592), .A2(n32431), .A3(n2594), .ZN(n35830) );
  NAND2_X1 U11763 ( .A1(n32427), .A2(n32426), .ZN(n2595) );
  XNOR2_X1 U11764 ( .A(n27276), .B(n27266), .ZN(n2596) );
  INV_X1 U11765 ( .A(n35966), .ZN(n38528) );
  AND3_X1 U11766 ( .A1(n2955), .A2(n28719), .A3(n28718), .ZN(n8423) );
  OR2_X1 U11767 ( .A1(n39210), .A2(n39426), .ZN(n5160) );
  OAI211_X1 U11768 ( .C1(n14312), .C2(n13824), .A(n14320), .B(n13819), .ZN(
        n14328) );
  OR2_X1 U11769 ( .A1(n44417), .A2(n46626), .ZN(n45769) );
  INV_X1 U11770 ( .A(n11066), .ZN(n8099) );
  XNOR2_X1 U11772 ( .A(n42797), .B(n2716), .ZN(n45659) );
  AND2_X1 U11773 ( .A1(n4954), .A2(n40572), .ZN(n2597) );
  INV_X1 U11774 ( .A(n51339), .ZN(n2788) );
  OR2_X1 U11775 ( .A1(n43455), .A2(n49987), .ZN(n2803) );
  INV_X1 U11776 ( .A(n23551), .ZN(n22276) );
  INV_X1 U11777 ( .A(n30171), .ZN(n2815) );
  OR2_X1 U11778 ( .A1(n32199), .A2(n3963), .ZN(n25407) );
  NOR2_X1 U11779 ( .A1(n13202), .A2(n13207), .ZN(n7591) );
  OAI21_X1 U11780 ( .B1(n38696), .B2(n39236), .A(n39245), .ZN(n38698) );
  AOI22_X1 U11781 ( .A1(n37701), .A2(n37341), .B1(n39245), .B2(n37340), .ZN(
        n37696) );
  NOR2_X1 U11782 ( .A1(n39245), .A2(n3873), .ZN(n37335) );
  AND2_X1 U11783 ( .A1(n51508), .A2(n39245), .ZN(n39223) );
  INV_X1 U11784 ( .A(n30705), .ZN(n27588) );
  NOR2_X1 U11785 ( .A1(n38666), .A2(n37924), .ZN(n3706) );
  NOR2_X1 U11786 ( .A1(n50732), .A2(n50727), .ZN(n4078) );
  INV_X1 U11787 ( .A(n27830), .ZN(n29448) );
  OR2_X1 U11788 ( .A1(n27830), .A2(n7826), .ZN(n27839) );
  INV_X1 U11789 ( .A(n25176), .ZN(n25892) );
  INV_X1 U11790 ( .A(n15400), .ZN(n6605) );
  XNOR2_X1 U11791 ( .A(n18216), .B(n15224), .ZN(n15400) );
  INV_X1 U11792 ( .A(n30925), .ZN(n31513) );
  AND2_X1 U11793 ( .A1(n11337), .A2(n11343), .ZN(n7280) );
  INV_X1 U11794 ( .A(n37097), .ZN(n2598) );
  NAND2_X1 U11795 ( .A1(n38301), .A2(n2342), .ZN(n38307) );
  XNOR2_X1 U11797 ( .A(n37303), .B(n34169), .ZN(n8482) );
  NOR2_X1 U11798 ( .A1(n353), .A2(n22375), .ZN(n22298) );
  NOR2_X1 U11800 ( .A1(n21293), .A2(n7655), .ZN(n7654) );
  INV_X1 U11801 ( .A(n21293), .ZN(n21302) );
  OR2_X1 U11802 ( .A1(n2118), .A2(n20215), .ZN(n7859) );
  OR2_X1 U11803 ( .A1(n37654), .A2(n38313), .ZN(n38319) );
  AND2_X1 U11804 ( .A1(n7532), .A2(n5417), .ZN(n7531) );
  AND3_X1 U11805 ( .A1(n14536), .A2(n14552), .A3(n14533), .ZN(n12982) );
  NOR2_X1 U11806 ( .A1(n32879), .A2(n32867), .ZN(n33030) );
  OAI22_X1 U11807 ( .A1(n48115), .A2(n48159), .B1(n48117), .B2(n48116), .ZN(
        n8201) );
  INV_X1 U11808 ( .A(n37019), .ZN(n37310) );
  OAI22_X1 U11809 ( .A1(n7052), .A2(n29270), .B1(n29272), .B2(n29187), .ZN(
        n28717) );
  INV_X1 U11810 ( .A(n29272), .ZN(n8242) );
  OR2_X2 U11811 ( .A1(n51138), .A2(n11354), .ZN(n12379) );
  AND3_X1 U11812 ( .A1(n28843), .A2(n28842), .A3(n4741), .ZN(n28845) );
  AND2_X1 U11813 ( .A1(n4198), .A2(n35850), .ZN(n35860) );
  AND2_X1 U11814 ( .A1(n12882), .A2(n13198), .ZN(n11861) );
  AND3_X2 U11816 ( .A1(n3378), .A2(n7189), .A3(n18972), .ZN(n22979) );
  INV_X1 U11817 ( .A(n23568), .ZN(n23562) );
  AOI21_X1 U11819 ( .B1(n49994), .B2(n50008), .A(n50329), .ZN(n7504) );
  OR2_X1 U11820 ( .A1(n38638), .A2(n38635), .ZN(n4816) );
  AND2_X1 U11822 ( .A1(n27669), .A2(n51117), .ZN(n27656) );
  OR2_X1 U11823 ( .A1(n27668), .A2(n51117), .ZN(n27654) );
  NOR2_X1 U11826 ( .A1(n12506), .A2(n51653), .ZN(n7694) );
  OR2_X1 U11827 ( .A1(n642), .A2(n51653), .ZN(n11255) );
  NOR2_X1 U11828 ( .A1(n40340), .A2(n40338), .ZN(n2665) );
  NOR2_X1 U11829 ( .A1(n39857), .A2(n40338), .ZN(n8608) );
  AOI21_X1 U11831 ( .B1(n36216), .B2(n37798), .A(n37806), .ZN(n36209) );
  INV_X1 U11832 ( .A(n36216), .ZN(n8198) );
  AND2_X1 U11833 ( .A1(n31385), .A2(n33005), .ZN(n33016) );
  OR2_X1 U11834 ( .A1(n3241), .A2(n33005), .ZN(n30531) );
  AND3_X1 U11835 ( .A1(n19985), .A2(n19986), .A3(n19984), .ZN(n8362) );
  XNOR2_X1 U11836 ( .A(n5613), .B(n51752), .ZN(n24735) );
  XNOR2_X1 U11838 ( .A(n51680), .B(n43623), .ZN(n45279) );
  AND2_X1 U11839 ( .A1(n9250), .A2(n9251), .ZN(n8653) );
  NOR2_X1 U11840 ( .A1(n3840), .A2(n3836), .ZN(n3835) );
  AND2_X1 U11841 ( .A1(n41557), .A2(n41559), .ZN(n5533) );
  AND2_X1 U11843 ( .A1(n46446), .A2(n42512), .ZN(n46434) );
  AND2_X1 U11845 ( .A1(n13354), .A2(n14553), .ZN(n14540) );
  AND2_X1 U11846 ( .A1(n24287), .A2(n24278), .ZN(n3950) );
  INV_X1 U11848 ( .A(n452), .ZN(n2676) );
  NOR2_X1 U11849 ( .A1(n17046), .A2(n17047), .ZN(n18375) );
  INV_X1 U11850 ( .A(n17046), .ZN(n17049) );
  AND3_X1 U11851 ( .A1(n41153), .A2(n41148), .A3(n41147), .ZN(n6551) );
  OAI211_X1 U11852 ( .C1(n35704), .C2(n6784), .A(n6782), .B(n6780), .ZN(n6779)
         );
  XNOR2_X2 U11853 ( .A(n4650), .B(n4295), .ZN(n43968) );
  XNOR2_X2 U11854 ( .A(n4654), .B(Key[82]), .ZN(n43105) );
  XNOR2_X2 U11855 ( .A(n4641), .B(n4932), .ZN(n23370) );
  XNOR2_X2 U11856 ( .A(n4931), .B(n4752), .ZN(n33653) );
  XNOR2_X2 U11857 ( .A(n4886), .B(n4208), .ZN(n43293) );
  INV_X1 U11858 ( .A(n43263), .ZN(n2600) );
  INV_X1 U11859 ( .A(n2600), .ZN(n2601) );
  XNOR2_X2 U11860 ( .A(n4827), .B(Key[28]), .ZN(n44483) );
  INV_X1 U11861 ( .A(n2250), .ZN(n2603) );
  XNOR2_X2 U11862 ( .A(n5016), .B(n4737), .ZN(n42322) );
  XNOR2_X2 U11863 ( .A(n4847), .B(n4880), .ZN(n25040) );
  XOR2_X1 U11864 ( .A(n48843), .B(Key[101]), .Z(n45050) );
  INV_X1 U11865 ( .A(n45050), .ZN(n2604) );
  XNOR2_X2 U11866 ( .A(n1341), .B(n6031), .ZN(n24992) );
  XNOR2_X2 U11867 ( .A(n4343), .B(n4868), .ZN(n45106) );
  XNOR2_X2 U11868 ( .A(n4655), .B(n4721), .ZN(n41367) );
  XNOR2_X1 U11869 ( .A(Key[174]), .B(Key[150]), .ZN(n2605) );
  XNOR2_X2 U11870 ( .A(n4618), .B(n3481), .ZN(n35815) );
  XNOR2_X2 U11871 ( .A(n4869), .B(n4429), .ZN(n45463) );
  XNOR2_X2 U11872 ( .A(Key[118]), .B(Key[94]), .ZN(n33474) );
  XNOR2_X2 U11873 ( .A(Key[9]), .B(n4896), .ZN(n35107) );
  XNOR2_X2 U11874 ( .A(n4667), .B(n4838), .ZN(n44493) );
  XNOR2_X2 U11875 ( .A(n42668), .B(n4650), .ZN(n24057) );
  XNOR2_X2 U11876 ( .A(n4649), .B(n4837), .ZN(n23943) );
  XNOR2_X2 U11877 ( .A(n4666), .B(n4885), .ZN(n45107) );
  INV_X1 U11878 ( .A(n42327), .ZN(n5382) );
  XNOR2_X2 U11879 ( .A(n4895), .B(n4824), .ZN(n42327) );
  XNOR2_X2 U11880 ( .A(n4668), .B(n4694), .ZN(n33374) );
  XNOR2_X2 U11881 ( .A(n2183), .B(n3014), .ZN(n43702) );
  XNOR2_X2 U11882 ( .A(n4706), .B(n4651), .ZN(n38626) );
  XNOR2_X2 U11883 ( .A(n4613), .B(n4687), .ZN(n42889) );
  XNOR2_X2 U11884 ( .A(n4665), .B(n4705), .ZN(n41567) );
  XNOR2_X2 U11885 ( .A(n4744), .B(n4884), .ZN(n34265) );
  XNOR2_X2 U11886 ( .A(n4597), .B(n4536), .ZN(n26541) );
  XNOR2_X2 U11887 ( .A(n33429), .B(n33049), .ZN(n45105) );
  XNOR2_X2 U11888 ( .A(n4554), .B(n4157), .ZN(n33049) );
  XNOR2_X2 U11889 ( .A(n4286), .B(n4879), .ZN(n32856) );
  XNOR2_X1 U11890 ( .A(n17960), .B(n31432), .ZN(n3013) );
  XNOR2_X2 U11891 ( .A(n4676), .B(n4518), .ZN(n31432) );
  XNOR2_X2 U11892 ( .A(Key[183]), .B(n2117), .ZN(n41155) );
  XNOR2_X1 U11894 ( .A(n4638), .B(n4565), .ZN(n2608) );
  NAND2_X1 U11895 ( .A1(n2609), .A2(n29995), .ZN(n29996) );
  NOR2_X1 U11896 ( .A1(n2609), .A2(n31892), .ZN(n31421) );
  OAI21_X1 U11897 ( .B1(n27868), .B2(n2609), .A(n31151), .ZN(n27869) );
  NAND2_X1 U11898 ( .A1(n24212), .A2(n23066), .ZN(n6064) );
  NAND2_X1 U11899 ( .A1(n30608), .A2(n31089), .ZN(n30595) );
  INV_X1 U11900 ( .A(n27686), .ZN(n2611) );
  NAND2_X1 U11901 ( .A1(n2612), .A2(n38228), .ZN(n2721) );
  OAI22_X1 U11902 ( .A1(n38227), .A2(n38226), .B1(n38552), .B2(n35175), .ZN(
        n2612) );
  NAND3_X1 U11903 ( .A1(n49607), .A2(n49606), .A3(n49605), .ZN(n2613) );
  NAND2_X1 U11904 ( .A1(n51088), .A2(n49569), .ZN(n49607) );
  NOR2_X1 U11905 ( .A1(n51394), .A2(n40972), .ZN(n2615) );
  NAND2_X1 U11906 ( .A1(n40971), .A2(n2614), .ZN(n40974) );
  NAND2_X1 U11907 ( .A1(n40959), .A2(n2615), .ZN(n2614) );
  OAI22_X1 U11908 ( .A1(n27677), .A2(n6290), .B1(n27678), .B2(n27685), .ZN(
        n8338) );
  NAND2_X1 U11909 ( .A1(n8481), .A2(n26954), .ZN(n26775) );
  INV_X1 U11910 ( .A(n27690), .ZN(n6290) );
  AND2_X1 U11911 ( .A1(n27681), .A2(n27690), .ZN(n26771) );
  NAND2_X1 U11912 ( .A1(n2616), .A2(n40269), .ZN(n40087) );
  INV_X1 U11913 ( .A(n40272), .ZN(n2616) );
  XNOR2_X1 U11914 ( .A(n6293), .B(n6292), .ZN(n2617) );
  OAI21_X1 U11916 ( .B1(n34993), .B2(n36029), .A(n37957), .ZN(n37968) );
  OAI21_X1 U11917 ( .B1(n2619), .B2(n26815), .A(n2618), .ZN(n26817) );
  OR2_X1 U11918 ( .A1(n3783), .A2(n27685), .ZN(n2618) );
  INV_X1 U11919 ( .A(n26813), .ZN(n2619) );
  NAND2_X1 U11920 ( .A1(n6290), .A2(n27681), .ZN(n3783) );
  INV_X1 U11921 ( .A(n6449), .ZN(n27681) );
  OR2_X1 U11922 ( .A1(n2620), .A2(n14205), .ZN(n4207) );
  NOR2_X1 U11923 ( .A1(n13334), .A2(n2620), .ZN(n14895) );
  NAND2_X1 U11924 ( .A1(n14718), .A2(n14719), .ZN(n2620) );
  INV_X1 U11925 ( .A(n25825), .ZN(n2623) );
  NAND2_X1 U11926 ( .A1(n22791), .A2(n22790), .ZN(n2622) );
  NAND2_X1 U11927 ( .A1(n3055), .A2(n51021), .ZN(n22784) );
  NAND2_X1 U11928 ( .A1(n46229), .A2(n49199), .ZN(n2626) );
  OAI21_X1 U11929 ( .B1(n49212), .B2(n46228), .A(n2624), .ZN(n45975) );
  NAND2_X1 U11930 ( .A1(n2625), .A2(n49209), .ZN(n2624) );
  NAND3_X1 U11931 ( .A1(n2626), .A2(n52106), .A3(n6502), .ZN(n2625) );
  OAI211_X1 U11932 ( .C1(n2627), .C2(n2632), .A(n2629), .B(n47615), .ZN(n2877)
         );
  NAND2_X1 U11933 ( .A1(n47589), .A2(n2631), .ZN(n2630) );
  NAND2_X1 U11934 ( .A1(n47608), .A2(n51340), .ZN(n47601) );
  NAND2_X1 U11935 ( .A1(n47595), .A2(n47588), .ZN(n2632) );
  NAND2_X1 U11936 ( .A1(n28557), .A2(n30280), .ZN(n28561) );
  AOI21_X1 U11937 ( .B1(n28546), .B2(n26502), .A(n2633), .ZN(n26503) );
  INV_X1 U11938 ( .A(n28557), .ZN(n2633) );
  INV_X1 U11939 ( .A(n28558), .ZN(n2634) );
  NAND3_X1 U11940 ( .A1(n2637), .A2(n48875), .A3(n48916), .ZN(n2635) );
  NAND2_X1 U11941 ( .A1(n48847), .A2(n48862), .ZN(n2636) );
  NOR2_X1 U11942 ( .A1(n48919), .A2(n48853), .ZN(n48916) );
  INV_X1 U11943 ( .A(n39831), .ZN(n2639) );
  OAI21_X2 U11944 ( .B1(n9265), .B2(n9266), .A(n4313), .ZN(n2640) );
  NAND2_X1 U11945 ( .A1(n2640), .A2(n13885), .ZN(n14873) );
  NAND2_X1 U11946 ( .A1(n2640), .A2(n3696), .ZN(n14876) );
  NAND2_X1 U11948 ( .A1(n2640), .A2(n14880), .ZN(n13262) );
  NAND2_X1 U11949 ( .A1(n13886), .A2(n2640), .ZN(n9268) );
  NAND3_X1 U11950 ( .A1(n15421), .A2(n14871), .A3(n2640), .ZN(n9270) );
  NAND2_X1 U11951 ( .A1(n1555), .A2(n2640), .ZN(n13875) );
  OAI21_X1 U11952 ( .B1(n7245), .B2(n2640), .A(n3705), .ZN(n9267) );
  NAND2_X1 U11953 ( .A1(n27668), .A2(n2641), .ZN(n27661) );
  INV_X1 U11954 ( .A(n26937), .ZN(n2641) );
  NAND2_X1 U11956 ( .A1(n20024), .A2(n18287), .ZN(n2644) );
  NAND2_X1 U11957 ( .A1(n20025), .A2(n2648), .ZN(n2647) );
  INV_X1 U11958 ( .A(n20010), .ZN(n2652) );
  NAND2_X1 U11959 ( .A1(n677), .A2(n41150), .ZN(n2653) );
  XNOR2_X2 U11960 ( .A(n8832), .B(Key[23]), .ZN(n10147) );
  NAND2_X1 U11961 ( .A1(n10216), .A2(n52189), .ZN(n10913) );
  AND2_X1 U11962 ( .A1(n10143), .A2(n9807), .ZN(n10216) );
  INV_X1 U11963 ( .A(n2654), .ZN(n13132) );
  NAND2_X1 U11964 ( .A1(n3678), .A2(n14186), .ZN(n2654) );
  NAND3_X1 U11965 ( .A1(n2654), .A2(n13145), .A3(n14178), .ZN(n12212) );
  OAI21_X1 U11966 ( .B1(n5502), .B2(n2655), .A(n48103), .ZN(n8064) );
  NAND2_X1 U11967 ( .A1(n48112), .A2(n48136), .ZN(n2655) );
  INV_X1 U11968 ( .A(n46387), .ZN(n2656) );
  OR2_X1 U11969 ( .A1(n46396), .A2(n2657), .ZN(n46400) );
  NAND2_X1 U11970 ( .A1(n46387), .A2(n991), .ZN(n2657) );
  NAND2_X1 U11971 ( .A1(n2658), .A2(n4246), .ZN(n34641) );
  NAND2_X1 U11972 ( .A1(n36565), .A2(n63), .ZN(n2658) );
  NAND2_X1 U11973 ( .A1(n34948), .A2(n38034), .ZN(n2661) );
  MUX2_X1 U11974 ( .A(n36386), .B(n36387), .S(n34948), .Z(n36388) );
  NAND2_X1 U11975 ( .A1(n2662), .A2(n46464), .ZN(n46470) );
  NAND3_X1 U11976 ( .A1(n48551), .A2(n45635), .A3(n48548), .ZN(n48549) );
  NAND2_X1 U11977 ( .A1(n48227), .A2(n2207), .ZN(n48548) );
  AND2_X1 U11978 ( .A1(n48546), .A2(n48531), .ZN(n45635) );
  NAND2_X1 U11979 ( .A1(n48540), .A2(n48239), .ZN(n2663) );
  NAND2_X1 U11981 ( .A1(n40334), .A2(n2665), .ZN(n39642) );
  OAI211_X1 U11982 ( .C1(n2665), .C2(n40337), .A(n39863), .B(n40334), .ZN(
        n39865) );
  NAND3_X1 U11983 ( .A1(n10213), .A2(n2666), .A3(n10930), .ZN(n4014) );
  NAND2_X1 U11984 ( .A1(n10215), .A2(n10219), .ZN(n10930) );
  NAND2_X1 U11985 ( .A1(n10216), .A2(n10921), .ZN(n2666) );
  XNOR2_X1 U11986 ( .A(n2667), .B(n25937), .ZN(n24514) );
  XNOR2_X1 U11987 ( .A(n26274), .B(n2543), .ZN(n26134) );
  INV_X1 U11988 ( .A(n587), .ZN(n2668) );
  NAND2_X1 U11989 ( .A1(n2669), .A2(n27071), .ZN(n2674) );
  OAI211_X1 U11990 ( .C1(n27659), .C2(n3765), .A(n2448), .B(n2673), .ZN(n2672)
         );
  NAND2_X1 U11991 ( .A1(n27068), .A2(n27067), .ZN(n2673) );
  NAND2_X1 U11992 ( .A1(n23421), .A2(n2675), .ZN(n23431) );
  NAND2_X1 U11993 ( .A1(n22034), .A2(n20084), .ZN(n2675) );
  NAND2_X1 U11994 ( .A1(n2676), .A2(n3506), .ZN(n20084) );
  NAND2_X1 U11997 ( .A1(n13332), .A2(n13333), .ZN(n14894) );
  NAND2_X1 U11999 ( .A1(n2677), .A2(n26944), .ZN(n26945) );
  NOR2_X1 U12000 ( .A1(n27070), .A2(n24774), .ZN(n3764) );
  NAND3_X1 U12001 ( .A1(n38363), .A2(n2679), .A3(n2678), .ZN(n4577) );
  OAI211_X1 U12002 ( .C1(n39707), .C2(n41084), .A(n39712), .B(n41085), .ZN(
        n2678) );
  OR2_X1 U12003 ( .A1(n8317), .A2(n39707), .ZN(n2679) );
  NAND2_X1 U12004 ( .A1(n17532), .A2(n20021), .ZN(n17537) );
  INV_X1 U12007 ( .A(n12324), .ZN(n2680) );
  NAND2_X1 U12008 ( .A1(n45658), .A2(n46494), .ZN(n2684) );
  NAND2_X1 U12009 ( .A1(n48912), .A2(n48908), .ZN(n48920) );
  NAND3_X1 U12010 ( .A1(n2687), .A2(n46190), .A3(n45660), .ZN(n2686) );
  INV_X1 U12011 ( .A(n36604), .ZN(n34928) );
  OAI21_X1 U12012 ( .B1(n36614), .B2(n34930), .A(n2689), .ZN(n34655) );
  INV_X1 U12013 ( .A(n36609), .ZN(n2689) );
  NAND2_X1 U12014 ( .A1(n698), .A2(n51716), .ZN(n36609) );
  XNOR2_X2 U12015 ( .A(n34278), .B(n34771), .ZN(n36604) );
  XNOR2_X1 U12017 ( .A(n2690), .B(n18427), .ZN(n18798) );
  XNOR2_X1 U12018 ( .A(n485), .B(n2690), .ZN(n16472) );
  NAND2_X1 U12019 ( .A1(n8160), .A2(n51153), .ZN(n21751) );
  NAND2_X1 U12020 ( .A1(n17468), .A2(n19404), .ZN(n2692) );
  INV_X1 U12021 ( .A(n12324), .ZN(n3649) );
  NAND3_X1 U12024 ( .A1(n2833), .A2(n2230), .A3(n2694), .ZN(n6697) );
  NAND2_X1 U12025 ( .A1(n49137), .A2(n2695), .ZN(n43401) );
  NAND3_X1 U12028 ( .A1(n11001), .A2(n11000), .A3(n10246), .ZN(n2696) );
  INV_X1 U12030 ( .A(n14972), .ZN(n14162) );
  OAI21_X1 U12031 ( .B1(n2697), .B2(n51175), .A(n2698), .ZN(n14972) );
  NAND2_X1 U12032 ( .A1(n14156), .A2(n14155), .ZN(n2698) );
  NAND2_X1 U12033 ( .A1(n2699), .A2(n2502), .ZN(n30800) );
  NAND2_X1 U12034 ( .A1(n11014), .A2(n51762), .ZN(n2701) );
  OAI211_X1 U12035 ( .C1(n9029), .C2(n8776), .A(n9753), .B(n2703), .ZN(n2702)
         );
  INV_X1 U12037 ( .A(n9743), .ZN(n2704) );
  INV_X1 U12038 ( .A(n2705), .ZN(n41541) );
  NAND3_X1 U12039 ( .A1(n41535), .A2(n3494), .A3(n40986), .ZN(n2705) );
  NAND2_X1 U12040 ( .A1(n2705), .A2(n5546), .ZN(n40935) );
  NAND2_X1 U12041 ( .A1(n28957), .A2(n2707), .ZN(n28507) );
  NAND2_X1 U12042 ( .A1(n28947), .A2(n2511), .ZN(n28858) );
  NAND3_X1 U12043 ( .A1(n29804), .A2(n29802), .A3(n2707), .ZN(n28463) );
  NAND2_X1 U12044 ( .A1(n28864), .A2(n2706), .ZN(n28868) );
  NAND2_X1 U12046 ( .A1(n50114), .A2(n50101), .ZN(n50062) );
  NAND2_X1 U12047 ( .A1(n49966), .A2(n49965), .ZN(n2709) );
  NAND3_X1 U12048 ( .A1(n49967), .A2(n49969), .A3(n49968), .ZN(n2710) );
  XNOR2_X1 U12050 ( .A(n6729), .B(n2548), .ZN(n35657) );
  NAND4_X2 U12051 ( .A1(n16883), .A2(n7948), .A3(n16879), .A4(n8506), .ZN(
        n24292) );
  NAND2_X1 U12052 ( .A1(n2712), .A2(n2711), .ZN(n3488) );
  NAND2_X1 U12053 ( .A1(n23513), .A2(n23510), .ZN(n2711) );
  AND2_X1 U12056 ( .A1(n18942), .A2(n5936), .ZN(n18933) );
  NAND3_X1 U12057 ( .A1(n37192), .A2(n2714), .A3(n4761), .ZN(n4760) );
  NAND3_X1 U12058 ( .A1(n38330), .A2(n2714), .A3(n38322), .ZN(n38325) );
  OAI21_X1 U12059 ( .B1(n2714), .B2(n38345), .A(n37195), .ZN(n3709) );
  NAND2_X1 U12060 ( .A1(n3256), .A2(n2714), .ZN(n38327) );
  NAND2_X1 U12061 ( .A1(n37673), .A2(n2714), .ZN(n37674) );
  NOR2_X1 U12062 ( .A1(n35897), .A2(n2714), .ZN(n5739) );
  NAND2_X1 U12063 ( .A1(n45220), .A2(n2715), .ZN(n45221) );
  NAND2_X1 U12064 ( .A1(n2688), .A2(n46503), .ZN(n2715) );
  AND2_X1 U12066 ( .A1(n11127), .A2(n5297), .ZN(n2717) );
  NAND2_X1 U12067 ( .A1(n4221), .A2(n5297), .ZN(n14766) );
  NAND3_X1 U12068 ( .A1(n8314), .A2(n2718), .A3(n11127), .ZN(n14765) );
  NAND2_X1 U12069 ( .A1(n38545), .A2(n3817), .ZN(n35173) );
  OR2_X1 U12071 ( .A1(n35173), .A2(n38228), .ZN(n2720) );
  NAND2_X1 U12072 ( .A1(n2723), .A2(n2722), .ZN(n36013) );
  NAND2_X1 U12073 ( .A1(n2723), .A2(n36491), .ZN(n7436) );
  INV_X1 U12074 ( .A(n36565), .ZN(n2723) );
  NAND3_X1 U12075 ( .A1(n6116), .A2(n52211), .A3(n2726), .ZN(n2724) );
  OR2_X1 U12076 ( .A1(n2726), .A2(n51733), .ZN(n46030) );
  NOR2_X1 U12077 ( .A1(n2726), .A2(n46028), .ZN(n49650) );
  NOR2_X1 U12078 ( .A1(n2726), .A2(n49672), .ZN(n50020) );
  NOR2_X1 U12079 ( .A1(n49663), .A2(n2726), .ZN(n49673) );
  AND2_X1 U12080 ( .A1(n49656), .A2(n49657), .ZN(n2725) );
  OAI211_X1 U12081 ( .C1(n2730), .C2(n2736), .A(n2728), .B(n2727), .ZN(
        Plaintext[185]) );
  NAND2_X1 U12082 ( .A1(n2736), .A2(n46932), .ZN(n2727) );
  OAI21_X1 U12083 ( .B1(n2732), .B2(n2729), .A(n46932), .ZN(n2728) );
  INV_X1 U12084 ( .A(n46931), .ZN(n2729) );
  NAND2_X1 U12085 ( .A1(n46931), .A2(n4890), .ZN(n2731) );
  NAND3_X1 U12086 ( .A1(n2735), .A2(n2734), .A3(n2733), .ZN(n2732) );
  NAND2_X1 U12087 ( .A1(n50872), .A2(n2332), .ZN(n2733) );
  OAI21_X1 U12088 ( .B1(n50872), .B2(n50882), .A(n50853), .ZN(n2734) );
  NAND3_X1 U12089 ( .A1(n46927), .A2(n52093), .A3(n5295), .ZN(n2735) );
  OAI211_X1 U12090 ( .C1(n50873), .C2(n52093), .A(n50823), .B(n46930), .ZN(
        n2736) );
  AND2_X1 U12091 ( .A1(n7306), .A2(n2738), .ZN(n41931) );
  NAND2_X1 U12092 ( .A1(n42201), .A2(n2738), .ZN(n37824) );
  AND2_X1 U12093 ( .A1(n42209), .A2(n2738), .ZN(n38928) );
  NAND3_X1 U12094 ( .A1(n41939), .A2(n2738), .A3(n41938), .ZN(n41941) );
  NAND2_X1 U12095 ( .A1(n41926), .A2(n2737), .ZN(n39540) );
  AOI21_X1 U12096 ( .B1(n680), .B2(n40250), .A(n2738), .ZN(n35994) );
  NAND2_X1 U12097 ( .A1(n2740), .A2(n4062), .ZN(n35954) );
  NAND2_X1 U12098 ( .A1(n2740), .A2(n2739), .ZN(n35955) );
  NAND2_X1 U12099 ( .A1(n38503), .A2(n2463), .ZN(n2740) );
  NAND2_X1 U12100 ( .A1(n8316), .A2(n41087), .ZN(n3095) );
  NOR2_X1 U12102 ( .A1(n38290), .A2(n2741), .ZN(n4417) );
  INV_X1 U12105 ( .A(n48413), .ZN(n2742) );
  NAND2_X1 U12106 ( .A1(n2743), .A2(n41670), .ZN(n41235) );
  XNOR2_X1 U12107 ( .A(n41683), .B(n2743), .ZN(n7030) );
  NAND3_X1 U12108 ( .A1(n41677), .A2(n41684), .A3(n2743), .ZN(n39318) );
  OAI21_X1 U12109 ( .B1(n41242), .B2(n2743), .A(n41241), .ZN(n8391) );
  NAND3_X1 U12110 ( .A1(n21523), .A2(n16858), .A3(n18899), .ZN(n16861) );
  NAND2_X1 U12111 ( .A1(n20612), .A2(n21528), .ZN(n21523) );
  NOR2_X2 U12112 ( .A1(n51048), .A2(n20188), .ZN(n21528) );
  XNOR2_X2 U12113 ( .A(n16110), .B(n16109), .ZN(n20188) );
  NAND3_X1 U12115 ( .A1(n41939), .A2(n6580), .A3(n41932), .ZN(n2744) );
  INV_X1 U12117 ( .A(n2745), .ZN(n30505) );
  OAI21_X1 U12118 ( .B1(n30502), .B2(n32590), .A(n2746), .ZN(n2745) );
  NAND2_X1 U12119 ( .A1(n29622), .A2(n32988), .ZN(n30502) );
  NAND2_X1 U12120 ( .A1(n29264), .A2(n51114), .ZN(n2747) );
  NAND2_X1 U12121 ( .A1(n2748), .A2(n27007), .ZN(n24567) );
  OAI22_X1 U12122 ( .A1(n2748), .A2(n29455), .B1(n29460), .B2(n29456), .ZN(
        n29458) );
  INV_X1 U12123 ( .A(n27755), .ZN(n2748) );
  OAI211_X1 U12124 ( .C1(n23502), .C2(n24292), .A(n2750), .B(n24287), .ZN(
        n2876) );
  NAND2_X1 U12125 ( .A1(n21081), .A2(n23510), .ZN(n2750) );
  NAND2_X1 U12126 ( .A1(n7519), .A2(n7247), .ZN(n23502) );
  NAND2_X1 U12127 ( .A1(n617), .A2(n37484), .ZN(n35966) );
  NAND2_X1 U12128 ( .A1(n2751), .A2(n47159), .ZN(n47160) );
  NAND2_X1 U12129 ( .A1(n47159), .A2(n2753), .ZN(n2752) );
  NAND2_X1 U12130 ( .A1(n2464), .A2(n2754), .ZN(n5849) );
  NAND4_X2 U12131 ( .A1(n30883), .A2(n30885), .A3(n2755), .A4(n30884), .ZN(
        n35345) );
  INV_X1 U12132 ( .A(n35889), .ZN(n2757) );
  NAND3_X1 U12133 ( .A1(n2757), .A2(n38330), .A3(n38323), .ZN(n8459) );
  AND2_X1 U12135 ( .A1(n32830), .A2(n31401), .ZN(n2759) );
  NAND2_X1 U12136 ( .A1(n2758), .A2(n51618), .ZN(n30474) );
  NAND3_X1 U12137 ( .A1(n30392), .A2(n30690), .A3(n2761), .ZN(n28754) );
  INV_X1 U12138 ( .A(n29938), .ZN(n2761) );
  NAND3_X1 U12139 ( .A1(n41202), .A2(n5919), .A3(n51430), .ZN(n41205) );
  NAND2_X1 U12140 ( .A1(n38572), .A2(n38205), .ZN(n38206) );
  NAND2_X1 U12142 ( .A1(n26833), .A2(n27408), .ZN(n2762) );
  XNOR2_X2 U12145 ( .A(n14470), .B(n14469), .ZN(n20474) );
  NAND2_X1 U12146 ( .A1(n13032), .A2(n2765), .ZN(n5221) );
  INV_X1 U12148 ( .A(n40210), .ZN(n41677) );
  INV_X1 U12149 ( .A(n41242), .ZN(n2772) );
  NAND2_X1 U12150 ( .A1(n41234), .A2(n52198), .ZN(n41242) );
  NAND4_X2 U12151 ( .A1(n2770), .A2(n2769), .A3(n7609), .A4(n2767), .ZN(n44963) );
  NAND2_X1 U12152 ( .A1(n40716), .A2(n41685), .ZN(n2768) );
  NAND2_X1 U12153 ( .A1(n2772), .A2(n41683), .ZN(n2769) );
  NAND2_X1 U12154 ( .A1(n41677), .A2(n41244), .ZN(n2771) );
  NAND2_X1 U12157 ( .A1(n20256), .A2(n21617), .ZN(n21619) );
  INV_X1 U12158 ( .A(n21632), .ZN(n2773) );
  NOR2_X1 U12159 ( .A1(n30780), .A2(n30792), .ZN(n29902) );
  NAND3_X1 U12160 ( .A1(n161), .A2(n29909), .A3(n2774), .ZN(n27574) );
  NAND2_X1 U12161 ( .A1(n27411), .A2(n2774), .ZN(n23663) );
  NAND2_X1 U12162 ( .A1(n27568), .A2(n2774), .ZN(n27569) );
  NAND3_X1 U12163 ( .A1(n38546), .A2(n2776), .A3(n2775), .ZN(n6968) );
  NAND2_X1 U12164 ( .A1(n38542), .A2(n38541), .ZN(n2775) );
  AOI22_X1 U12165 ( .A1(n2245), .A2(n38544), .B1(n38545), .B2(n38553), .ZN(
        n2776) );
  NAND2_X1 U12166 ( .A1(n26829), .A2(n30789), .ZN(n2778) );
  NAND3_X1 U12167 ( .A1(n2373), .A2(n29896), .A3(n2778), .ZN(n26830) );
  NOR2_X1 U12168 ( .A1(n51394), .A2(n41380), .ZN(n41383) );
  OAI21_X1 U12169 ( .B1(n37631), .B2(n2783), .A(n2779), .ZN(n3447) );
  OAI211_X1 U12170 ( .C1(n38283), .C2(n37630), .A(n2781), .B(n2780), .ZN(n2779) );
  NAND2_X1 U12171 ( .A1(n37628), .A2(n38284), .ZN(n2780) );
  NOR2_X1 U12173 ( .A1(n38288), .A2(n38291), .ZN(n2784) );
  NAND2_X1 U12174 ( .A1(n37629), .A2(n38272), .ZN(n2785) );
  NAND2_X1 U12175 ( .A1(n38288), .A2(n38272), .ZN(n2786) );
  NOR2_X1 U12176 ( .A1(n37623), .A2(n37624), .ZN(n37628) );
  NAND2_X1 U12177 ( .A1(n710), .A2(n32242), .ZN(n32233) );
  INV_X1 U12178 ( .A(n31781), .ZN(n32246) );
  NAND2_X1 U12179 ( .A1(n41383), .A2(n40970), .ZN(n2789) );
  NAND2_X1 U12180 ( .A1(n49973), .A2(n2790), .ZN(n43452) );
  NAND2_X1 U12181 ( .A1(n49989), .A2(n2790), .ZN(n49623) );
  NAND3_X1 U12182 ( .A1(n32347), .A2(n32438), .A3(n723), .ZN(n2792) );
  NAND2_X1 U12183 ( .A1(n2792), .A2(n32436), .ZN(n32043) );
  NAND2_X1 U12184 ( .A1(n2792), .A2(n2791), .ZN(n31322) );
  OR2_X1 U12185 ( .A1(n32444), .A2(n31320), .ZN(n2791) );
  OAI211_X1 U12186 ( .C1(n50102), .C2(n51442), .A(n50047), .B(n2793), .ZN(
        n50048) );
  NAND2_X1 U12187 ( .A1(n50083), .A2(n2794), .ZN(n2793) );
  INV_X1 U12188 ( .A(n51644), .ZN(n50114) );
  NAND2_X1 U12189 ( .A1(n2846), .A2(n2510), .ZN(n5591) );
  NAND3_X1 U12190 ( .A1(n8369), .A2(n23022), .A3(n2795), .ZN(n23024) );
  NAND3_X1 U12191 ( .A1(n10608), .A2(n10072), .A3(n10069), .ZN(n2796) );
  AND3_X1 U12192 ( .A1(n41013), .A2(n51358), .A3(n40807), .ZN(n43328) );
  NAND2_X1 U12194 ( .A1(n31788), .A2(n29372), .ZN(n2797) );
  NAND3_X1 U12195 ( .A1(n2799), .A2(n27601), .A3(n2798), .ZN(n23862) );
  NAND3_X1 U12196 ( .A1(n2799), .A2(n27601), .A3(n26911), .ZN(n30678) );
  NAND2_X1 U12197 ( .A1(n2801), .A2(n23068), .ZN(n23592) );
  NAND2_X1 U12198 ( .A1(n2801), .A2(n24211), .ZN(n17419) );
  AND2_X1 U12199 ( .A1(n52155), .A2(n2801), .ZN(n2800) );
  NOR2_X1 U12200 ( .A1(n3170), .A2(n17420), .ZN(n2801) );
  NOR2_X1 U12201 ( .A1(n727), .A2(n30449), .ZN(n28839) );
  NAND3_X1 U12202 ( .A1(n30444), .A2(n2328), .A3(n727), .ZN(n28445) );
  NOR2_X1 U12203 ( .A1(n50277), .A2(n51410), .ZN(n2804) );
  NAND2_X1 U12205 ( .A1(n50540), .A2(n50521), .ZN(n50517) );
  AND2_X1 U12206 ( .A1(n2807), .A2(n50540), .ZN(n50537) );
  NAND2_X1 U12207 ( .A1(n50563), .A2(n50536), .ZN(n2807) );
  NAND2_X1 U12210 ( .A1(n19020), .A2(n19777), .ZN(n2809) );
  NOR2_X1 U12211 ( .A1(n7657), .A2(n45936), .ZN(n4460) );
  NAND2_X1 U12212 ( .A1(n44730), .A2(n49139), .ZN(n45936) );
  OR2_X1 U12213 ( .A1(n46290), .A2(n51016), .ZN(n49139) );
  NAND3_X1 U12214 ( .A1(n2810), .A2(n22376), .A3(n23814), .ZN(n2811) );
  OAI21_X1 U12215 ( .B1(n2813), .B2(n2244), .A(n22736), .ZN(n2812) );
  INV_X1 U12216 ( .A(n21062), .ZN(n22731) );
  OAI21_X1 U12217 ( .B1(n22375), .B2(n22373), .A(n21062), .ZN(n2813) );
  NAND2_X1 U12218 ( .A1(n353), .A2(n22390), .ZN(n21062) );
  NAND3_X1 U12219 ( .A1(n22385), .A2(n753), .A3(n5371), .ZN(n2814) );
  AND2_X1 U12220 ( .A1(n8310), .A2(n353), .ZN(n22385) );
  NAND2_X1 U12221 ( .A1(n29622), .A2(n32986), .ZN(n32586) );
  NOR2_X1 U12222 ( .A1(n29618), .A2(n29616), .ZN(n32986) );
  NAND2_X1 U12223 ( .A1(n2815), .A2(n30163), .ZN(n28023) );
  NAND2_X1 U12224 ( .A1(n8091), .A2(n2816), .ZN(n27596) );
  NAND2_X1 U12225 ( .A1(n28800), .A2(n2817), .ZN(n2816) );
  NAND2_X1 U12226 ( .A1(n30725), .A2(n30716), .ZN(n2817) );
  AND2_X1 U12227 ( .A1(n30711), .A2(n2205), .ZN(n30725) );
  NAND2_X2 U12228 ( .A1(n52218), .A2(n30706), .ZN(n30723) );
  NAND2_X1 U12230 ( .A1(n19675), .A2(n18234), .ZN(n19676) );
  NAND2_X1 U12234 ( .A1(n27671), .A2(n24776), .ZN(n2819) );
  OAI22_X1 U12235 ( .A1(n27661), .A2(n748), .B1(n2819), .B2(n27670), .ZN(
        n24761) );
  NOR2_X1 U12236 ( .A1(n2821), .A2(n2820), .ZN(n2823) );
  NAND2_X1 U12237 ( .A1(n31003), .A2(n32025), .ZN(n2821) );
  OAI21_X2 U12238 ( .B1(n2823), .B2(n2822), .A(n27650), .ZN(n36940) );
  NAND3_X1 U12239 ( .A1(n46271), .A2(n2825), .A3(n46270), .ZN(n2824) );
  NAND2_X1 U12240 ( .A1(n49019), .A2(n51397), .ZN(n48984) );
  OAI21_X1 U12241 ( .B1(n13667), .B2(n13653), .A(n12755), .ZN(n2827) );
  NAND2_X1 U12242 ( .A1(n11514), .A2(n12573), .ZN(n2828) );
  NAND3_X1 U12243 ( .A1(n7341), .A2(n12574), .A3(n2828), .ZN(n11573) );
  NAND3_X1 U12244 ( .A1(n11575), .A2(n7341), .A3(n2828), .ZN(n11576) );
  NAND2_X1 U12245 ( .A1(n41797), .A2(n38812), .ZN(n42104) );
  NAND2_X1 U12246 ( .A1(n4734), .A2(n33787), .ZN(n38812) );
  XNOR2_X1 U12247 ( .A(n17240), .B(n2501), .ZN(n8512) );
  NAND2_X1 U12248 ( .A1(n22849), .A2(n23020), .ZN(n21877) );
  NAND2_X1 U12249 ( .A1(n6701), .A2(n49460), .ZN(n2833) );
  INV_X2 U12250 ( .A(n22329), .ZN(n22857) );
  NAND3_X1 U12251 ( .A1(n23023), .A2(n22334), .A3(n4413), .ZN(n22335) );
  NAND2_X1 U12252 ( .A1(n22849), .A2(n22329), .ZN(n23023) );
  NAND3_X1 U12253 ( .A1(n2834), .A2(n40002), .A3(n39668), .ZN(n39669) );
  NAND2_X1 U12254 ( .A1(n2836), .A2(n718), .ZN(n6155) );
  INV_X1 U12255 ( .A(n32048), .ZN(n2836) );
  NAND2_X1 U12256 ( .A1(n32048), .A2(n32438), .ZN(n2837) );
  NAND2_X1 U12257 ( .A1(n723), .A2(n32439), .ZN(n32048) );
  NAND2_X1 U12258 ( .A1(n4550), .A2(n12579), .ZN(n2839) );
  XNOR2_X1 U12259 ( .A(n32997), .B(n2841), .ZN(n5238) );
  XNOR2_X1 U12260 ( .A(n32997), .B(n33862), .ZN(n33863) );
  XNOR2_X1 U12261 ( .A(n32997), .B(n2550), .ZN(n37293) );
  XNOR2_X1 U12262 ( .A(n36792), .B(n2842), .ZN(n33352) );
  XNOR2_X1 U12263 ( .A(n34842), .B(n2842), .ZN(n33963) );
  XNOR2_X1 U12264 ( .A(n35800), .B(n2842), .ZN(n34436) );
  NOR2_X1 U12265 ( .A1(n27058), .A2(n27053), .ZN(n2844) );
  INV_X1 U12266 ( .A(n27053), .ZN(n27701) );
  OAI21_X1 U12267 ( .B1(n2847), .B2(n2846), .A(n23025), .ZN(n21017) );
  NOR2_X1 U12268 ( .A1(n2091), .A2(n32705), .ZN(n32707) );
  NOR2_X1 U12269 ( .A1(n32324), .A2(n2091), .ZN(n30141) );
  NAND2_X1 U12270 ( .A1(n1988), .A2(n2091), .ZN(n31666) );
  NAND2_X1 U12271 ( .A1(n29814), .A2(n2091), .ZN(n32331) );
  NOR2_X1 U12272 ( .A1(n32692), .A2(n2091), .ZN(n29816) );
  AOI21_X1 U12273 ( .B1(n32692), .B2(n32693), .A(n2091), .ZN(n32696) );
  OAI21_X1 U12274 ( .B1(n31661), .B2(n2091), .A(n4334), .ZN(n31673) );
  NAND2_X1 U12275 ( .A1(n40450), .A2(n39738), .ZN(n39741) );
  INV_X1 U12276 ( .A(n40447), .ZN(n2848) );
  NAND4_X2 U12277 ( .A1(n37206), .A2(n37208), .A3(n37207), .A4(n37205), .ZN(
        n40447) );
  INV_X1 U12278 ( .A(n49967), .ZN(n47276) );
  NAND2_X1 U12279 ( .A1(n2849), .A2(n2850), .ZN(n49967) );
  NAND2_X1 U12280 ( .A1(n50351), .A2(n50344), .ZN(n2849) );
  AND2_X1 U12281 ( .A1(n47270), .A2(n555), .ZN(n2850) );
  NAND2_X1 U12282 ( .A1(n2851), .A2(n30452), .ZN(n28518) );
  INV_X1 U12283 ( .A(n28517), .ZN(n2851) );
  NAND4_X1 U12284 ( .A1(n36047), .A2(n36052), .A3(n36590), .A4(n35879), .ZN(
        n36044) );
  NAND2_X1 U12285 ( .A1(n36591), .A2(n36456), .ZN(n7505) );
  NAND2_X1 U12286 ( .A1(n2852), .A2(n32727), .ZN(n32728) );
  INV_X1 U12287 ( .A(n32464), .ZN(n2852) );
  AND2_X2 U12288 ( .A1(n12403), .A2(n7865), .ZN(n14033) );
  NAND2_X1 U12289 ( .A1(n2855), .A2(n40453), .ZN(n40397) );
  NAND2_X1 U12291 ( .A1(n2854), .A2(n40450), .ZN(n3530) );
  INV_X1 U12292 ( .A(n40453), .ZN(n2854) );
  AND2_X1 U12293 ( .A1(n49462), .A2(n2859), .ZN(n49423) );
  INV_X1 U12294 ( .A(n49449), .ZN(n2857) );
  NAND3_X1 U12295 ( .A1(n49434), .A2(n49422), .A3(n2856), .ZN(n49426) );
  NAND2_X1 U12296 ( .A1(n2857), .A2(n49442), .ZN(n2856) );
  NAND2_X1 U12297 ( .A1(n49443), .A2(n2859), .ZN(n49420) );
  OR2_X2 U12298 ( .A1(n45975), .A2(n45974), .ZN(n2859) );
  NAND2_X1 U12299 ( .A1(n19988), .A2(n51755), .ZN(n2860) );
  NAND2_X1 U12300 ( .A1(n21556), .A2(n21555), .ZN(n21413) );
  INV_X1 U12301 ( .A(n50912), .ZN(n2862) );
  INV_X1 U12302 ( .A(n50920), .ZN(n2864) );
  NAND2_X1 U12303 ( .A1(n35704), .A2(n38566), .ZN(n33064) );
  NAND2_X1 U12305 ( .A1(n2867), .A2(n41692), .ZN(n41704) );
  OAI211_X1 U12306 ( .C1(n15106), .C2(n14252), .A(n13690), .B(n14977), .ZN(
        n8975) );
  NAND2_X1 U12307 ( .A1(n2868), .A2(n14251), .ZN(n13690) );
  NOR2_X1 U12308 ( .A1(n3458), .A2(n3457), .ZN(n2869) );
  NAND2_X1 U12310 ( .A1(n46605), .A2(n46604), .ZN(n2870) );
  NOR2_X1 U12313 ( .A1(n12809), .A2(n13034), .ZN(n2871) );
  NOR2_X1 U12314 ( .A1(n21769), .A2(n51081), .ZN(n21779) );
  NAND2_X1 U12315 ( .A1(n30550), .A2(n2872), .ZN(n30557) );
  NAND2_X1 U12316 ( .A1(n39098), .A2(n2360), .ZN(n37843) );
  NAND2_X1 U12318 ( .A1(n4907), .A2(n30856), .ZN(n31578) );
  NAND2_X1 U12319 ( .A1(n49165), .A2(n49164), .ZN(n2874) );
  NAND2_X1 U12320 ( .A1(n49166), .A2(n49167), .ZN(n2875) );
  NAND2_X1 U12321 ( .A1(n2876), .A2(n3937), .ZN(n21088) );
  NOR2_X1 U12322 ( .A1(n47267), .A2(n2877), .ZN(n47269) );
  NAND2_X1 U12323 ( .A1(n31680), .A2(n2094), .ZN(n30006) );
  NAND2_X1 U12324 ( .A1(n30007), .A2(n30983), .ZN(n2878) );
  NOR2_X1 U12325 ( .A1(n2539), .A2(n21233), .ZN(n2879) );
  INV_X1 U12327 ( .A(n39817), .ZN(n41333) );
  NAND2_X1 U12328 ( .A1(n41328), .A2(n52214), .ZN(n39817) );
  NAND2_X1 U12329 ( .A1(n2881), .A2(n2195), .ZN(n26501) );
  INV_X1 U12330 ( .A(n26494), .ZN(n2881) );
  OAI21_X1 U12334 ( .B1(n2883), .B2(n38516), .A(n38515), .ZN(n38526) );
  INV_X1 U12335 ( .A(n37446), .ZN(n2883) );
  NAND2_X1 U12336 ( .A1(n51735), .A2(n38535), .ZN(n37446) );
  AND2_X1 U12337 ( .A1(n11900), .A2(n800), .ZN(n11484) );
  NAND3_X1 U12338 ( .A1(n12727), .A2(n12729), .A3(n12728), .ZN(n12731) );
  OR2_X1 U12340 ( .A1(n11682), .A2(n2885), .ZN(n11691) );
  OAI21_X1 U12341 ( .B1(n11685), .B2(n11684), .A(n11683), .ZN(n2885) );
  NAND2_X1 U12343 ( .A1(n2888), .A2(n41079), .ZN(n38876) );
  AND2_X1 U12344 ( .A1(n34644), .A2(n34642), .ZN(n2887) );
  NAND2_X1 U12345 ( .A1(n38055), .A2(n38057), .ZN(n36336) );
  INV_X1 U12347 ( .A(n27783), .ZN(n29192) );
  INV_X1 U12348 ( .A(n29269), .ZN(n6660) );
  OAI21_X1 U12349 ( .B1(n31726), .B2(n6577), .A(n32282), .ZN(n32285) );
  AND2_X1 U12350 ( .A1(n21712), .A2(n22184), .ZN(n22189) );
  INV_X1 U12352 ( .A(n19778), .ZN(n19462) );
  NAND2_X1 U12353 ( .A1(n19118), .A2(n21276), .ZN(n19778) );
  NAND2_X1 U12354 ( .A1(n2890), .A2(n34664), .ZN(n6596) );
  NAND2_X1 U12355 ( .A1(n3578), .A2(n3580), .ZN(n2890) );
  NAND2_X1 U12357 ( .A1(n28332), .A2(n29859), .ZN(n28336) );
  NOR2_X1 U12359 ( .A1(n37624), .A2(n2123), .ZN(n35417) );
  INV_X1 U12360 ( .A(n44518), .ZN(n7900) );
  INV_X1 U12361 ( .A(n6965), .ZN(n6962) );
  NAND3_X1 U12362 ( .A1(n22469), .A2(n20527), .A3(n4718), .ZN(n22309) );
  NAND2_X1 U12363 ( .A1(n4719), .A2(n22721), .ZN(n22469) );
  NAND3_X1 U12364 ( .A1(n22874), .A2(n25056), .A3(n23101), .ZN(n21688) );
  NAND3_X1 U12366 ( .A1(n33459), .A2(n36195), .A3(n33460), .ZN(n33463) );
  OR2_X1 U12367 ( .A1(n14533), .A2(n14370), .ZN(n3672) );
  NAND2_X1 U12370 ( .A1(n4210), .A2(n13440), .ZN(n13442) );
  NAND2_X1 U12371 ( .A1(n31991), .A2(n2891), .ZN(n7666) );
  NAND2_X1 U12372 ( .A1(n31986), .A2(n29677), .ZN(n2891) );
  NAND2_X1 U12373 ( .A1(n7386), .A2(n9713), .ZN(n2892) );
  INV_X1 U12377 ( .A(n20041), .ZN(n2893) );
  NAND2_X1 U12378 ( .A1(n16814), .A2(n18377), .ZN(n20041) );
  NAND2_X1 U12379 ( .A1(n23470), .A2(n2894), .ZN(n21963) );
  INV_X1 U12381 ( .A(n38631), .ZN(n2896) );
  NAND2_X1 U12382 ( .A1(n3311), .A2(n38252), .ZN(n38627) );
  NAND3_X1 U12384 ( .A1(n13300), .A2(n13299), .A3(n14033), .ZN(n4634) );
  AND2_X1 U12385 ( .A1(n18381), .A2(n16814), .ZN(n16815) );
  NAND3_X1 U12386 ( .A1(n17609), .A2(n22156), .A3(n21026), .ZN(n5018) );
  NAND3_X1 U12387 ( .A1(n2897), .A2(n37957), .A3(n3554), .ZN(n36043) );
  NAND3_X1 U12388 ( .A1(n3555), .A2(n36028), .A3(n6218), .ZN(n2897) );
  NAND2_X1 U12390 ( .A1(n42799), .A2(n42800), .ZN(n2898) );
  AOI21_X1 U12392 ( .B1(n2901), .B2(n40200), .A(n2900), .ZN(n38388) );
  NAND2_X1 U12393 ( .A1(n40111), .A2(n40201), .ZN(n2901) );
  XNOR2_X1 U12394 ( .A(n2902), .B(n6229), .ZN(Plaintext[0]) );
  NAND3_X1 U12395 ( .A1(n6233), .A2(n6230), .A3(n6232), .ZN(n2902) );
  AND3_X1 U12397 ( .A1(n43578), .A2(n46010), .A3(n50328), .ZN(n4552) );
  NAND2_X1 U12398 ( .A1(n7823), .A2(n12276), .ZN(n9007) );
  AND2_X1 U12399 ( .A1(n32925), .A2(n32926), .ZN(n4702) );
  INV_X1 U12400 ( .A(n22935), .ZN(n22086) );
  NAND2_X1 U12401 ( .A1(n23044), .A2(n424), .ZN(n22935) );
  XNOR2_X1 U12403 ( .A(n15932), .B(n19244), .ZN(n17240) );
  AND3_X1 U12404 ( .A1(n39906), .A2(n37356), .A3(n6645), .ZN(n39788) );
  AND2_X1 U12406 ( .A1(n19706), .A2(n2299), .ZN(n8309) );
  OR2_X1 U12407 ( .A1(n39182), .A2(n38663), .ZN(n38678) );
  AND2_X1 U12409 ( .A1(n6340), .A2(n6337), .ZN(n6336) );
  AND2_X1 U12410 ( .A1(n13854), .A2(n14472), .ZN(n6793) );
  XNOR2_X1 U12412 ( .A(n33303), .B(n6729), .ZN(n35285) );
  XNOR2_X1 U12413 ( .A(n6846), .B(n43983), .ZN(n46380) );
  INV_X1 U12415 ( .A(n9057), .ZN(n2905) );
  AOI22_X1 U12416 ( .A1(n46502), .A2(n46499), .B1(n46500), .B2(n46501), .ZN(
        n46507) );
  INV_X1 U12417 ( .A(n13818), .ZN(n13598) );
  INV_X1 U12418 ( .A(n47477), .ZN(n48974) );
  NOR2_X1 U12419 ( .A1(n5776), .A2(n10289), .ZN(n9742) );
  INV_X1 U12420 ( .A(n42020), .ZN(n6654) );
  INV_X1 U12421 ( .A(n37195), .ZN(n38338) );
  INV_X1 U12422 ( .A(n30577), .ZN(n5181) );
  INV_X1 U12423 ( .A(n47554), .ZN(n5787) );
  XNOR2_X1 U12424 ( .A(n43937), .B(n43936), .ZN(n44505) );
  NAND2_X1 U12425 ( .A1(n2906), .A2(n31347), .ZN(n31332) );
  INV_X1 U12426 ( .A(n31334), .ZN(n2906) );
  XNOR2_X1 U12427 ( .A(n28046), .B(n7180), .ZN(n28622) );
  NAND3_X1 U12428 ( .A1(n11132), .A2(n51139), .A3(n10474), .ZN(n10478) );
  OR2_X2 U12430 ( .A1(n15141), .A2(n3439), .ZN(n16711) );
  AND2_X2 U12431 ( .A1(n36148), .A2(n31355), .ZN(n38557) );
  NAND2_X1 U12432 ( .A1(n16892), .A2(n16886), .ZN(n6629) );
  NAND2_X1 U12433 ( .A1(n5347), .A2(n14270), .ZN(n15128) );
  NAND2_X1 U12434 ( .A1(n26351), .A2(n26352), .ZN(n4685) );
  NAND2_X1 U12435 ( .A1(n23824), .A2(n2908), .ZN(n23830) );
  NOR2_X2 U12436 ( .A1(n23821), .A2(n23827), .ZN(n23824) );
  OAI21_X1 U12437 ( .B1(n41764), .B2(n42145), .A(n2909), .ZN(n40887) );
  NAND2_X1 U12438 ( .A1(n42145), .A2(n2382), .ZN(n2909) );
  NAND2_X1 U12440 ( .A1(n10585), .A2(n2911), .ZN(n2910) );
  NAND2_X1 U12441 ( .A1(n29498), .A2(n26666), .ZN(n2912) );
  NAND2_X1 U12442 ( .A1(n23254), .A2(n23247), .ZN(n22654) );
  INV_X1 U12443 ( .A(n11955), .ZN(n12724) );
  NAND3_X1 U12444 ( .A1(n4891), .A2(n20803), .A3(n20804), .ZN(n20808) );
  NOR2_X1 U12445 ( .A1(n2381), .A2(n2913), .ZN(n3495) );
  NAND2_X1 U12447 ( .A1(n9220), .A2(n6328), .ZN(n2914) );
  NAND2_X1 U12448 ( .A1(n9219), .A2(n10665), .ZN(n2915) );
  NAND2_X1 U12451 ( .A1(n39450), .A2(n39027), .ZN(n39448) );
  XNOR2_X2 U12452 ( .A(n34725), .B(n8504), .ZN(n39450) );
  NAND2_X2 U12453 ( .A1(n3313), .A2(n3733), .ZN(n8403) );
  NAND2_X1 U12456 ( .A1(n2918), .A2(n46908), .ZN(n45855) );
  NAND4_X1 U12458 ( .A1(n2920), .A2(n8193), .A3(n39042), .A4(n2919), .ZN(n8197) );
  NAND2_X1 U12459 ( .A1(n41703), .A2(n41170), .ZN(n2919) );
  INV_X1 U12460 ( .A(n8192), .ZN(n2920) );
  XNOR2_X1 U12462 ( .A(n2922), .B(n39725), .ZN(n39810) );
  XNOR2_X1 U12463 ( .A(n39661), .B(n39660), .ZN(n2922) );
  NAND3_X1 U12465 ( .A1(n38740), .A2(n40736), .A3(n40737), .ZN(n4496) );
  NAND2_X1 U12466 ( .A1(n10645), .A2(n10646), .ZN(n10651) );
  AND2_X2 U12467 ( .A1(n50366), .A2(n50364), .ZN(n46984) );
  NAND3_X1 U12470 ( .A1(n32774), .A2(n32775), .A3(n32764), .ZN(n2923) );
  NAND2_X1 U12471 ( .A1(n18731), .A2(n15998), .ZN(n21626) );
  NAND2_X1 U12473 ( .A1(n33015), .A2(n33016), .ZN(n2924) );
  INV_X1 U12474 ( .A(n21304), .ZN(n3685) );
  AND3_X2 U12475 ( .A1(n7363), .A2(n9428), .A3(n9427), .ZN(n12834) );
  NAND3_X1 U12476 ( .A1(n7476), .A2(n50438), .A3(n2925), .ZN(n50449) );
  OAI211_X1 U12477 ( .C1(n7891), .C2(n12087), .A(n12385), .B(n12389), .ZN(
        n2926) );
  NAND2_X1 U12478 ( .A1(n11188), .A2(n7341), .ZN(n5622) );
  NAND2_X1 U12479 ( .A1(n7340), .A2(n2927), .ZN(n11188) );
  OR2_X1 U12480 ( .A1(n38204), .A2(n38201), .ZN(n8578) );
  INV_X1 U12481 ( .A(n14724), .ZN(n13749) );
  NAND3_X1 U12482 ( .A1(n14717), .A2(n14724), .A3(n14712), .ZN(n14080) );
  AND2_X1 U12483 ( .A1(n14716), .A2(n14711), .ZN(n14724) );
  INV_X1 U12484 ( .A(n12835), .ZN(n14671) );
  OAI21_X1 U12485 ( .B1(n3228), .B2(n19849), .A(n19848), .ZN(n2929) );
  NAND2_X1 U12486 ( .A1(n21166), .A2(n2930), .ZN(n2996) );
  OR2_X1 U12487 ( .A1(n20357), .A2(n19170), .ZN(n18050) );
  INV_X1 U12488 ( .A(n18056), .ZN(n3351) );
  NAND3_X1 U12489 ( .A1(n4135), .A2(n30638), .A3(n5817), .ZN(n5816) );
  OAI21_X1 U12491 ( .B1(n3509), .B2(n5229), .A(n19786), .ZN(n2931) );
  INV_X1 U12492 ( .A(n11884), .ZN(n12458) );
  NAND2_X1 U12493 ( .A1(n24277), .A2(n20982), .ZN(n7527) );
  NAND3_X1 U12494 ( .A1(n30652), .A2(n31298), .A3(n31303), .ZN(n24784) );
  OAI22_X1 U12495 ( .A1(n39197), .A2(n39196), .B1(n39374), .B2(n39390), .ZN(
        n8393) );
  XNOR2_X2 U12496 ( .A(n52119), .B(n34754), .ZN(n36714) );
  XNOR2_X1 U12497 ( .A(n7900), .B(n44519), .ZN(n46565) );
  AOI22_X1 U12498 ( .A1(n16880), .A2(n7946), .B1(n8502), .B2(n7949), .ZN(n7948) );
  AND3_X1 U12499 ( .A1(n6594), .A2(n20492), .A3(n4240), .ZN(n20500) );
  INV_X1 U12500 ( .A(n19891), .ZN(n19658) );
  NOR2_X1 U12501 ( .A1(n20965), .A2(n20966), .ZN(n18369) );
  AND2_X1 U12502 ( .A1(n10005), .A2(n10000), .ZN(n9997) );
  INV_X1 U12503 ( .A(n47094), .ZN(n47106) );
  AND2_X1 U12504 ( .A1(n6176), .A2(n21475), .ZN(n6175) );
  INV_X1 U12506 ( .A(n23981), .ZN(n6967) );
  XNOR2_X1 U12507 ( .A(n25566), .B(n26364), .ZN(n7428) );
  INV_X1 U12508 ( .A(n29462), .ZN(n27758) );
  INV_X1 U12509 ( .A(n24292), .ZN(n7707) );
  INV_X1 U12510 ( .A(n41275), .ZN(n7218) );
  INV_X1 U12511 ( .A(n39377), .ZN(n37032) );
  OAI21_X1 U12512 ( .B1(n8077), .B2(n38727), .A(n5569), .ZN(n38725) );
  AOI22_X1 U12513 ( .A1(n1906), .A2(n30698), .B1(n30695), .B2(n30395), .ZN(
        n30397) );
  NAND4_X1 U12515 ( .A1(n24884), .A2(n30299), .A3(n24883), .A4(n2932), .ZN(
        n24888) );
  NAND2_X1 U12516 ( .A1(n2111), .A2(n27110), .ZN(n2932) );
  XNOR2_X2 U12518 ( .A(n15505), .B(n15506), .ZN(n18085) );
  NAND3_X1 U12519 ( .A1(n46346), .A2(n46343), .A3(n46356), .ZN(n4089) );
  NOR2_X1 U12520 ( .A1(n13488), .A2(n13486), .ZN(n12775) );
  NAND2_X1 U12521 ( .A1(n15044), .A2(n15048), .ZN(n13488) );
  NAND2_X1 U12522 ( .A1(n2933), .A2(n3036), .ZN(n28471) );
  NAND2_X1 U12524 ( .A1(n6993), .A2(n2934), .ZN(n38764) );
  OR2_X1 U12525 ( .A1(n37425), .A2(n38468), .ZN(n35144) );
  NAND2_X1 U12527 ( .A1(n31273), .A2(n621), .ZN(n31481) );
  INV_X1 U12528 ( .A(n22099), .ZN(n24024) );
  NOR2_X1 U12529 ( .A1(n22575), .A2(n354), .ZN(n4188) );
  XNOR2_X1 U12530 ( .A(n2935), .B(n47498), .ZN(Plaintext[1]) );
  NAND4_X1 U12531 ( .A1(n47497), .A2(n47496), .A3(n47494), .A4(n47495), .ZN(
        n2935) );
  NAND4_X2 U12532 ( .A1(n9728), .A2(n9727), .A3(n9726), .A4(n9725), .ZN(n17646) );
  AND2_X1 U12534 ( .A1(n5113), .A2(n6384), .ZN(n6383) );
  NAND3_X1 U12535 ( .A1(n19677), .A2(n20214), .A3(n19676), .ZN(n19697) );
  NAND3_X1 U12536 ( .A1(n19102), .A2(n2937), .A3(n2936), .ZN(n19104) );
  NAND2_X1 U12537 ( .A1(n21254), .A2(n21256), .ZN(n2937) );
  NAND3_X1 U12538 ( .A1(n50232), .A2(n50222), .A3(n50233), .ZN(n50157) );
  NAND3_X1 U12539 ( .A1(n14701), .A2(n14719), .A3(n14700), .ZN(n14707) );
  NAND3_X1 U12540 ( .A1(n9539), .A2(n3692), .A3(n11132), .ZN(n11130) );
  XNOR2_X2 U12541 ( .A(n6141), .B(n2938), .ZN(n27764) );
  XNOR2_X1 U12542 ( .A(n24560), .B(n24559), .ZN(n2938) );
  XNOR2_X2 U12543 ( .A(n2939), .B(n15028), .ZN(n6952) );
  XNOR2_X1 U12544 ( .A(n15709), .B(n15027), .ZN(n2939) );
  NAND2_X1 U12545 ( .A1(n52226), .A2(n50638), .ZN(n50622) );
  NAND4_X2 U12546 ( .A1(n2940), .A2(n38510), .A3(n38508), .A4(n38509), .ZN(
        n41319) );
  NAND2_X1 U12548 ( .A1(n8333), .A2(n2943), .ZN(n2942) );
  NAND2_X1 U12549 ( .A1(n2944), .A2(n6892), .ZN(n2943) );
  NAND3_X1 U12550 ( .A1(n14359), .A2(n14369), .A3(n3673), .ZN(n12434) );
  NAND2_X1 U12551 ( .A1(n14720), .A2(n14713), .ZN(n14199) );
  AND4_X2 U12552 ( .A1(n12347), .A2(n12349), .A3(n12348), .A4(n12346), .ZN(
        n14713) );
  NAND2_X1 U12553 ( .A1(n2946), .A2(n2945), .ZN(n5190) );
  NAND2_X1 U12554 ( .A1(n14948), .A2(n14949), .ZN(n2945) );
  NAND2_X1 U12555 ( .A1(n14947), .A2(n51724), .ZN(n2946) );
  NAND3_X1 U12556 ( .A1(n22916), .A2(n22363), .A3(n22908), .ZN(n21041) );
  NAND2_X1 U12557 ( .A1(n27795), .A2(n28618), .ZN(n29505) );
  XNOR2_X1 U12559 ( .A(n44338), .B(n43390), .ZN(n43394) );
  NAND3_X1 U12561 ( .A1(n44269), .A2(n48204), .A3(n45539), .ZN(n2949) );
  XNOR2_X1 U12562 ( .A(n25463), .B(n25049), .ZN(n2950) );
  INV_X1 U12563 ( .A(n35179), .ZN(n35178) );
  NOR2_X1 U12564 ( .A1(n14269), .A2(n15132), .ZN(n3461) );
  AND3_X2 U12565 ( .A1(n33466), .A2(n33455), .A3(n6876), .ZN(n38810) );
  OR2_X1 U12566 ( .A1(n12373), .A2(n12384), .ZN(n9679) );
  INV_X1 U12567 ( .A(n20046), .ZN(n16826) );
  OR2_X1 U12568 ( .A1(n22704), .A2(n2980), .ZN(n4860) );
  NAND2_X1 U12569 ( .A1(n29802), .A2(n2337), .ZN(n28510) );
  NAND2_X1 U12571 ( .A1(n6799), .A2(n14520), .ZN(n6798) );
  NAND2_X1 U12572 ( .A1(n15173), .A2(n15177), .ZN(n14124) );
  AND3_X1 U12573 ( .A1(n5621), .A2(n10864), .A3(n11512), .ZN(n5619) );
  INV_X1 U12574 ( .A(n25213), .ZN(n8368) );
  INV_X1 U12575 ( .A(n11579), .ZN(n11189) );
  AOI21_X1 U12576 ( .B1(n11278), .B2(n11277), .A(n4186), .ZN(n11285) );
  AND3_X1 U12577 ( .A1(n23915), .A2(n23916), .A3(n23917), .ZN(n4696) );
  INV_X1 U12578 ( .A(n14394), .ZN(n12872) );
  MUX2_X1 U12579 ( .A(n19602), .B(n22864), .S(n22857), .Z(n19608) );
  XNOR2_X1 U12581 ( .A(n2951), .B(n50400), .ZN(Plaintext[150]) );
  NAND3_X1 U12582 ( .A1(n5223), .A2(n5225), .A3(n5222), .ZN(n2951) );
  NAND3_X1 U12584 ( .A1(n31764), .A2(n50981), .A3(n32197), .ZN(n7250) );
  NAND2_X1 U12586 ( .A1(n629), .A2(n23341), .ZN(n21737) );
  NAND2_X1 U12587 ( .A1(n16798), .A2(n6363), .ZN(n5813) );
  INV_X1 U12589 ( .A(n11227), .ZN(n2954) );
  NAND3_X2 U12590 ( .A1(n5124), .A2(n5125), .A3(n40356), .ZN(n44979) );
  NAND3_X1 U12591 ( .A1(n31403), .A2(n31404), .A3(n31402), .ZN(n31405) );
  NAND3_X1 U12592 ( .A1(n28720), .A2(n28721), .A3(n8713), .ZN(n28722) );
  OAI21_X1 U12593 ( .B1(n7051), .B2(n29281), .A(n8421), .ZN(n2955) );
  NAND2_X1 U12594 ( .A1(n24113), .A2(n24106), .ZN(n24107) );
  NAND2_X1 U12595 ( .A1(n31931), .A2(n30053), .ZN(n30036) );
  NAND2_X1 U12596 ( .A1(n19488), .A2(n20052), .ZN(n3197) );
  NOR2_X1 U12597 ( .A1(n30424), .A2(n487), .ZN(n6771) );
  AOI21_X1 U12598 ( .B1(n22243), .B2(n23964), .A(n4061), .ZN(n22248) );
  INV_X1 U12600 ( .A(n39450), .ZN(n3479) );
  INV_X1 U12601 ( .A(n12893), .ZN(n4949) );
  NAND3_X1 U12602 ( .A1(n13669), .A2(n3254), .A3(n13667), .ZN(n13645) );
  NAND2_X2 U12603 ( .A1(n4586), .A2(n9093), .ZN(n13667) );
  NAND3_X1 U12604 ( .A1(n29034), .A2(n28875), .A3(n27104), .ZN(n27102) );
  INV_X1 U12605 ( .A(n12678), .ZN(n11879) );
  NAND2_X1 U12606 ( .A1(n11082), .A2(n11884), .ZN(n12678) );
  NAND2_X1 U12607 ( .A1(n28545), .A2(n28148), .ZN(n28559) );
  NAND2_X1 U12608 ( .A1(n3292), .A2(n13082), .ZN(n2957) );
  NAND2_X1 U12609 ( .A1(n2958), .A2(n38132), .ZN(n32148) );
  OAI21_X1 U12610 ( .B1(n36329), .B2(n38136), .A(n2959), .ZN(n2958) );
  OAI21_X1 U12612 ( .B1(n29938), .B2(n51113), .A(n2960), .ZN(n28750) );
  NAND2_X1 U12613 ( .A1(n30688), .A2(n51113), .ZN(n2960) );
  NAND3_X1 U12614 ( .A1(n2962), .A2(n9128), .A3(n2961), .ZN(n8382) );
  NAND2_X1 U12615 ( .A1(n5826), .A2(n9127), .ZN(n2961) );
  OR2_X1 U12616 ( .A1(n14529), .A2(n13377), .ZN(n13390) );
  NAND4_X2 U12617 ( .A1(n6225), .A2(n19531), .A3(n19532), .A4(n19533), .ZN(
        n23445) );
  INV_X1 U12618 ( .A(n31283), .ZN(n7907) );
  XOR2_X1 U12619 ( .A(n27263), .B(n26608), .Z(n8120) );
  XNOR2_X1 U12620 ( .A(n18150), .B(n3587), .ZN(n17142) );
  NAND2_X1 U12621 ( .A1(n7077), .A2(n23832), .ZN(n2963) );
  NAND2_X1 U12623 ( .A1(n2965), .A2(n20032), .ZN(n16830) );
  OAI211_X1 U12624 ( .C1(n16826), .C2(n16823), .A(n20039), .B(n16825), .ZN(
        n2965) );
  AOI21_X1 U12625 ( .B1(n3659), .B2(n30852), .A(n3658), .ZN(n3657) );
  NAND2_X1 U12626 ( .A1(n2966), .A2(n31021), .ZN(n3151) );
  NAND2_X1 U12627 ( .A1(n3152), .A2(n2967), .ZN(n2966) );
  XNOR2_X2 U12628 ( .A(n6921), .B(n33360), .ZN(n3675) );
  NAND2_X2 U12629 ( .A1(n30131), .A2(n30132), .ZN(n6921) );
  NAND3_X1 U12630 ( .A1(n30572), .A2(n3688), .A3(n3687), .ZN(n26710) );
  OR2_X1 U12631 ( .A1(n28978), .A2(n28979), .ZN(n28980) );
  NAND2_X1 U12633 ( .A1(n6661), .A2(n2968), .ZN(n12247) );
  OAI211_X1 U12634 ( .C1(n48991), .C2(n48990), .A(n49036), .B(n48989), .ZN(
        n48992) );
  NAND2_X1 U12635 ( .A1(n49034), .A2(n2969), .ZN(n48989) );
  NAND2_X1 U12638 ( .A1(n6037), .A2(n6036), .ZN(n2970) );
  NAND4_X2 U12639 ( .A1(n12192), .A2(n12191), .A3(n14529), .A4(n12190), .ZN(
        n18689) );
  NAND3_X1 U12640 ( .A1(n2971), .A2(n41351), .A3(n41350), .ZN(n8122) );
  NAND2_X1 U12641 ( .A1(n41347), .A2(n8123), .ZN(n2971) );
  INV_X1 U12643 ( .A(n6571), .ZN(n12074) );
  INV_X1 U12645 ( .A(n25708), .ZN(n25605) );
  XNOR2_X1 U12646 ( .A(n25708), .B(n51719), .ZN(n24790) );
  NAND3_X1 U12648 ( .A1(n41573), .A2(n42015), .A3(n2973), .ZN(n41508) );
  NAND3_X1 U12649 ( .A1(n2975), .A2(n17409), .A3(n17408), .ZN(n7792) );
  OAI21_X1 U12650 ( .B1(n17407), .B2(n18112), .A(n19734), .ZN(n2975) );
  NAND3_X1 U12651 ( .A1(n10845), .A2(n10844), .A3(n10843), .ZN(n10857) );
  NAND3_X1 U12652 ( .A1(n11469), .A2(n11629), .A3(n11634), .ZN(n11472) );
  INV_X1 U12653 ( .A(n9103), .ZN(n2976) );
  OAI211_X1 U12654 ( .C1(n14548), .C2(n14368), .A(n2978), .B(n2977), .ZN(
        n12984) );
  NAND2_X1 U12655 ( .A1(n14363), .A2(n14544), .ZN(n2977) );
  NAND2_X1 U12656 ( .A1(n14536), .A2(n3038), .ZN(n2978) );
  NAND2_X1 U12658 ( .A1(n45205), .A2(n48461), .ZN(n2979) );
  INV_X1 U12659 ( .A(n22705), .ZN(n2980) );
  INV_X1 U12661 ( .A(n30283), .ZN(n28148) );
  XNOR2_X1 U12662 ( .A(n15575), .B(n13720), .ZN(n16834) );
  INV_X1 U12663 ( .A(n18071), .ZN(n18072) );
  NAND3_X1 U12664 ( .A1(n45235), .A2(n46274), .A3(n45236), .ZN(n45249) );
  NAND4_X2 U12666 ( .A1(n15058), .A2(n15057), .A3(n2981), .A4(n15056), .ZN(
        n16754) );
  NAND2_X1 U12670 ( .A1(n27627), .A2(n27623), .ZN(n2982) );
  INV_X1 U12671 ( .A(n24803), .ZN(n8498) );
  XOR2_X1 U12672 ( .A(n51668), .B(n13535), .Z(n5136) );
  NAND2_X1 U12674 ( .A1(n2984), .A2(n32974), .ZN(n32601) );
  AND2_X1 U12677 ( .A1(n2987), .A2(n21555), .ZN(n4363) );
  NAND2_X1 U12678 ( .A1(n3752), .A2(n15364), .ZN(n14806) );
  INV_X1 U12679 ( .A(n10262), .ZN(n4176) );
  NAND3_X1 U12680 ( .A1(n4834), .A2(n45906), .A3(n49714), .ZN(n3300) );
  XNOR2_X1 U12681 ( .A(n2988), .B(n37001), .ZN(n37002) );
  XNOR2_X1 U12682 ( .A(n37000), .B(n36999), .ZN(n2988) );
  NAND2_X1 U12683 ( .A1(n10013), .A2(n11663), .ZN(n11657) );
  INV_X1 U12684 ( .A(n32395), .ZN(n31290) );
  AND2_X1 U12687 ( .A1(n33160), .A2(n33162), .ZN(n3984) );
  NAND3_X1 U12688 ( .A1(n51683), .A2(n13526), .A3(n11841), .ZN(n8002) );
  NAND4_X1 U12690 ( .A1(n2989), .A2(n28524), .A3(n30449), .A4(n29737), .ZN(
        n28525) );
  OAI21_X1 U12691 ( .B1(n28521), .B2(n30458), .A(n28523), .ZN(n2989) );
  NAND3_X1 U12692 ( .A1(n20479), .A2(n20478), .A3(n20480), .ZN(n20481) );
  NOR2_X1 U12694 ( .A1(n13255), .A2(n13260), .ZN(n2990) );
  NAND2_X1 U12695 ( .A1(n2991), .A2(n30422), .ZN(n3374) );
  NAND2_X1 U12696 ( .A1(n30420), .A2(n30421), .ZN(n2991) );
  NAND3_X1 U12697 ( .A1(n31909), .A2(n31261), .A3(n32421), .ZN(n31262) );
  OAI211_X1 U12698 ( .C1(n31260), .C2(n8536), .A(n31259), .B(n31258), .ZN(
        n31909) );
  NAND2_X1 U12699 ( .A1(n46654), .A2(n47118), .ZN(n46838) );
  INV_X1 U12701 ( .A(n30497), .ZN(n2993) );
  OAI21_X1 U12702 ( .B1(n28941), .B2(n28940), .A(n28939), .ZN(n2994) );
  OAI22_X1 U12703 ( .A1(n29065), .A2(n5389), .B1(n30354), .B2(n29061), .ZN(
        n28851) );
  NAND2_X1 U12704 ( .A1(n28936), .A2(n28937), .ZN(n4142) );
  NAND2_X1 U12705 ( .A1(n28687), .A2(n28686), .ZN(n2995) );
  NAND2_X1 U12706 ( .A1(n30940), .A2(n7957), .ZN(n30942) );
  NAND2_X1 U12707 ( .A1(n7659), .A2(n31110), .ZN(n30940) );
  NAND2_X1 U12708 ( .A1(n8941), .A2(n12538), .ZN(n10778) );
  AND3_X1 U12709 ( .A1(n9374), .A2(n9373), .A3(n9375), .ZN(n2997) );
  NAND2_X1 U12710 ( .A1(n36266), .A2(n33676), .ZN(n36281) );
  NAND2_X1 U12711 ( .A1(n49423), .A2(n49424), .ZN(n49425) );
  INV_X1 U12712 ( .A(n41691), .ZN(n5475) );
  NAND2_X1 U12713 ( .A1(n31082), .A2(n31918), .ZN(n2998) );
  NAND2_X1 U12714 ( .A1(n32839), .A2(n32844), .ZN(n2999) );
  INV_X1 U12715 ( .A(n49420), .ZN(n49418) );
  INV_X1 U12716 ( .A(n15562), .ZN(n6285) );
  XNOR2_X1 U12717 ( .A(n5999), .B(n34780), .ZN(n34875) );
  OAI22_X1 U12718 ( .A1(n41616), .A2(n5043), .B1(n41706), .B2(n41617), .ZN(
        n41618) );
  NOR2_X2 U12719 ( .A1(n24008), .A2(n24007), .ZN(n25682) );
  NAND4_X1 U12720 ( .A1(n41325), .A2(n38604), .A3(n40729), .A4(n52214), .ZN(
        n38605) );
  AND2_X1 U12723 ( .A1(n4277), .A2(n20998), .ZN(n7353) );
  NAND2_X1 U12724 ( .A1(n3000), .A2(n19927), .ZN(n3475) );
  NAND2_X1 U12725 ( .A1(n20758), .A2(n19285), .ZN(n3000) );
  INV_X1 U12726 ( .A(n36305), .ZN(n6734) );
  NAND2_X1 U12727 ( .A1(n3100), .A2(n23507), .ZN(n24285) );
  OAI22_X1 U12729 ( .A1(n10986), .A2(n9782), .B1(n10987), .B2(n10990), .ZN(
        n3001) );
  INV_X1 U12730 ( .A(n35409), .ZN(n3251) );
  INV_X1 U12731 ( .A(n50019), .ZN(n46029) );
  AND3_X1 U12734 ( .A1(n13872), .A2(n12029), .A3(n12035), .ZN(n3359) );
  INV_X1 U12735 ( .A(n43580), .ZN(n50315) );
  XNOR2_X1 U12736 ( .A(n36961), .B(n36960), .ZN(n3061) );
  INV_X1 U12737 ( .A(n34604), .ZN(n6581) );
  NAND4_X1 U12739 ( .A1(n27912), .A2(n29340), .A3(n27909), .A4(n27906), .ZN(
        n30623) );
  AND3_X1 U12740 ( .A1(n11130), .A2(n11129), .A3(n2540), .ZN(n11142) );
  INV_X1 U12741 ( .A(n12145), .ZN(n11411) );
  INV_X1 U12742 ( .A(n23825), .ZN(n3520) );
  XNOR2_X1 U12743 ( .A(n37262), .B(n36940), .ZN(n34128) );
  INV_X1 U12744 ( .A(n2174), .ZN(n5737) );
  INV_X1 U12745 ( .A(n13277), .ZN(n15188) );
  INV_X1 U12746 ( .A(n21355), .ZN(n19284) );
  INV_X1 U12748 ( .A(n14434), .ZN(n14102) );
  NOR2_X1 U12749 ( .A1(n23955), .A2(n5069), .ZN(n23623) );
  NAND4_X1 U12750 ( .A1(n11427), .A2(n11426), .A3(n11425), .A4(n6477), .ZN(
        n11433) );
  INV_X1 U12751 ( .A(n22157), .ZN(n3423) );
  NOR2_X1 U12752 ( .A1(n50329), .A2(n50316), .ZN(n6992) );
  INV_X1 U12753 ( .A(n40125), .ZN(n3094) );
  NOR2_X1 U12754 ( .A1(n14762), .A2(n15206), .ZN(n14764) );
  NOR2_X1 U12755 ( .A1(n30698), .A2(n30694), .ZN(n4267) );
  XNOR2_X1 U12756 ( .A(n35360), .B(n35359), .ZN(n6833) );
  AOI22_X1 U12757 ( .A1(n36001), .A2(n36002), .B1(n36003), .B2(n37635), .ZN(
        n36007) );
  NAND2_X1 U12758 ( .A1(n7938), .A2(n20984), .ZN(n3938) );
  NAND2_X1 U12760 ( .A1(n20981), .A2(n20984), .ZN(n21913) );
  NAND3_X1 U12761 ( .A1(n3003), .A2(n23341), .A3(n23342), .ZN(n3002) );
  XNOR2_X1 U12762 ( .A(n3004), .B(n16703), .ZN(n16705) );
  XNOR2_X1 U12763 ( .A(n16702), .B(n16701), .ZN(n3004) );
  NAND2_X1 U12765 ( .A1(n9052), .A2(n9051), .ZN(n3005) );
  XNOR2_X2 U12766 ( .A(n42979), .B(n44160), .ZN(n44394) );
  XNOR2_X1 U12767 ( .A(n34111), .B(n3006), .ZN(n3365) );
  XNOR2_X1 U12768 ( .A(n34119), .B(n34120), .ZN(n3006) );
  NAND2_X1 U12769 ( .A1(n7369), .A2(n29282), .ZN(n29284) );
  NAND4_X1 U12770 ( .A1(n37502), .A2(n36244), .A3(n37500), .A4(n3527), .ZN(
        n3528) );
  NAND2_X1 U12771 ( .A1(n3007), .A2(n29528), .ZN(n27804) );
  NAND4_X1 U12772 ( .A1(n23707), .A2(n23703), .A3(n5415), .A4(n23536), .ZN(
        n22239) );
  NAND2_X1 U12773 ( .A1(n3008), .A2(n39212), .ZN(n39216) );
  OAI22_X1 U12774 ( .A1(n37907), .A2(n39208), .B1(n39206), .B2(n39207), .ZN(
        n3008) );
  NAND2_X1 U12775 ( .A1(n3715), .A2(n18021), .ZN(n19402) );
  NAND2_X1 U12776 ( .A1(n7997), .A2(n28546), .ZN(n28554) );
  NAND2_X1 U12777 ( .A1(n15306), .A2(n3009), .ZN(n13791) );
  NAND2_X1 U12778 ( .A1(n25199), .A2(n30178), .ZN(n29141) );
  OR3_X1 U12779 ( .A1(n10003), .A2(n11023), .A3(n10005), .ZN(n9998) );
  INV_X1 U12780 ( .A(n32426), .ZN(n3011) );
  AND4_X1 U12781 ( .A1(n12425), .A2(n12426), .A3(n12428), .A4(n12427), .ZN(
        n3012) );
  NAND2_X1 U12782 ( .A1(n15330), .A2(n15329), .ZN(n3016) );
  NAND2_X1 U12783 ( .A1(n13352), .A2(n14370), .ZN(n14551) );
  XNOR2_X1 U12784 ( .A(n3018), .B(n44966), .ZN(n44968) );
  XNOR2_X1 U12785 ( .A(n44961), .B(n44960), .ZN(n3018) );
  OAI21_X1 U12786 ( .B1(n2415), .B2(n3019), .A(n51302), .ZN(n47506) );
  NOR2_X1 U12788 ( .A1(n8058), .A2(n7764), .ZN(n3020) );
  AOI22_X1 U12789 ( .A1(n3021), .A2(n41577), .B1(n41412), .B2(n42021), .ZN(
        n41423) );
  INV_X1 U12790 ( .A(n41414), .ZN(n3021) );
  NAND2_X1 U12791 ( .A1(n42011), .A2(n42006), .ZN(n41414) );
  XOR2_X1 U12792 ( .A(n34357), .B(n36713), .Z(n7732) );
  NAND4_X2 U12794 ( .A1(n12875), .A2(n12874), .A3(n12873), .A4(n12962), .ZN(
        n17665) );
  NAND2_X1 U12795 ( .A1(n4149), .A2(n11632), .ZN(n3025) );
  NAND2_X2 U12796 ( .A1(n27866), .A2(n27867), .ZN(n31892) );
  NAND4_X1 U12797 ( .A1(n20834), .A2(n20832), .A3(n20831), .A4(n20833), .ZN(
        n3026) );
  AOI21_X1 U12798 ( .B1(n6553), .B2(n36895), .A(n39035), .ZN(n3027) );
  NAND2_X1 U12799 ( .A1(n26933), .A2(n27652), .ZN(n7784) );
  NAND2_X1 U12800 ( .A1(n35150), .A2(n6783), .ZN(n3028) );
  NAND3_X2 U12801 ( .A1(n34432), .A2(n7730), .A3(n7595), .ZN(n41084) );
  INV_X1 U12802 ( .A(n41035), .ZN(n39115) );
  NAND2_X1 U12804 ( .A1(n23165), .A2(n3032), .ZN(n8214) );
  NAND2_X1 U12805 ( .A1(n23176), .A2(n51021), .ZN(n3032) );
  MUX2_X1 U12806 ( .A(n19893), .B(n19892), .S(n3033), .Z(n19895) );
  AND2_X1 U12807 ( .A1(n19894), .A2(n3033), .ZN(n19666) );
  NAND2_X1 U12808 ( .A1(n19658), .A2(n5936), .ZN(n18944) );
  AOI21_X1 U12809 ( .B1(n19657), .B2(n51127), .A(n3033), .ZN(n19661) );
  AOI22_X1 U12810 ( .A1(n18938), .A2(n19894), .B1(n51127), .B2(n3033), .ZN(
        n16882) );
  INV_X2 U12811 ( .A(n32761), .ZN(n32962) );
  NAND2_X2 U12812 ( .A1(n28193), .A2(n8714), .ZN(n32761) );
  NAND3_X1 U12814 ( .A1(n32765), .A2(n32761), .A3(n32766), .ZN(n3036) );
  NAND2_X1 U12815 ( .A1(n14551), .A2(n14542), .ZN(n6069) );
  INV_X1 U12816 ( .A(n11376), .ZN(n3039) );
  NAND2_X1 U12817 ( .A1(n3039), .A2(n51391), .ZN(n11374) );
  NAND3_X1 U12818 ( .A1(n12112), .A2(n12113), .A3(n12114), .ZN(n12115) );
  NAND2_X1 U12819 ( .A1(n39448), .A2(n51737), .ZN(n36257) );
  NAND2_X1 U12820 ( .A1(n39035), .A2(n39036), .ZN(n39451) );
  INV_X1 U12822 ( .A(n3042), .ZN(n22211) );
  NAND3_X1 U12823 ( .A1(n3042), .A2(n8353), .A3(n22207), .ZN(n4468) );
  NAND2_X1 U12824 ( .A1(n37596), .A2(n37378), .ZN(n3044) );
  NAND2_X1 U12825 ( .A1(n37592), .A2(n3044), .ZN(n3129) );
  INV_X1 U12826 ( .A(n32182), .ZN(n32533) );
  NAND2_X1 U12827 ( .A1(n32962), .A2(n32957), .ZN(n32182) );
  NAND3_X1 U12828 ( .A1(n37775), .A2(n37778), .A3(n37774), .ZN(n3048) );
  NAND2_X1 U12829 ( .A1(n3050), .A2(n37782), .ZN(n3049) );
  NAND4_X1 U12830 ( .A1(n6982), .A2(n6981), .A3(n2357), .A4(n35941), .ZN(n3050) );
  INV_X1 U12831 ( .A(n5844), .ZN(n42179) );
  NAND2_X1 U12832 ( .A1(n42175), .A2(n45521), .ZN(n5844) );
  NAND2_X1 U12833 ( .A1(n3052), .A2(n44283), .ZN(n3051) );
  NAND2_X1 U12834 ( .A1(n3053), .A2(n44282), .ZN(n3052) );
  NAND2_X1 U12835 ( .A1(n45820), .A2(n45521), .ZN(n3053) );
  NAND2_X1 U12836 ( .A1(n44817), .A2(n42179), .ZN(n3054) );
  NAND2_X1 U12837 ( .A1(n3055), .A2(n23166), .ZN(n22673) );
  XNOR2_X1 U12838 ( .A(n3056), .B(n48018), .ZN(Plaintext[36]) );
  NAND3_X1 U12839 ( .A1(n48017), .A2(n3058), .A3(n3057), .ZN(n3056) );
  NAND2_X1 U12840 ( .A1(n48072), .A2(n2526), .ZN(n3057) );
  AND2_X1 U12841 ( .A1(n48016), .A2(n48015), .ZN(n3058) );
  NAND2_X1 U12842 ( .A1(n48003), .A2(n48038), .ZN(n48072) );
  NAND2_X1 U12844 ( .A1(n28688), .A2(n51518), .ZN(n26084) );
  INV_X1 U12845 ( .A(n3060), .ZN(n17454) );
  NAND2_X1 U12848 ( .A1(n32798), .A2(n32787), .ZN(n3064) );
  NAND3_X1 U12849 ( .A1(n32150), .A2(n32153), .A3(n3064), .ZN(n32155) );
  OAI22_X1 U12850 ( .A1(n32782), .A2(n3064), .B1(n2432), .B2(n32791), .ZN(
        n32783) );
  NAND3_X1 U12851 ( .A1(n32165), .A2(n32166), .A3(n3063), .ZN(n32167) );
  XNOR2_X1 U12852 ( .A(n3065), .B(n33605), .ZN(n35337) );
  INV_X1 U12853 ( .A(n33382), .ZN(n3065) );
  XNOR2_X1 U12854 ( .A(n35072), .B(n3066), .ZN(n35073) );
  INV_X1 U12855 ( .A(n33605), .ZN(n3066) );
  NOR2_X1 U12856 ( .A1(n3067), .A2(n29715), .ZN(n28182) );
  OAI21_X1 U12857 ( .B1(n30418), .B2(n30419), .A(n3067), .ZN(n30420) );
  OR2_X1 U12858 ( .A1(n5405), .A2(n37991), .ZN(n3068) );
  NAND3_X1 U12861 ( .A1(n37782), .A2(n52054), .A3(n39335), .ZN(n3072) );
  INV_X1 U12863 ( .A(n17546), .ZN(n3073) );
  INV_X1 U12865 ( .A(n48077), .ZN(n3076) );
  INV_X1 U12866 ( .A(n48083), .ZN(n3075) );
  NAND2_X1 U12868 ( .A1(n13525), .A2(n51683), .ZN(n11845) );
  INV_X1 U12869 ( .A(n10563), .ZN(n3079) );
  NAND3_X1 U12871 ( .A1(n10899), .A2(n10898), .A3(n13170), .ZN(n13774) );
  NAND2_X1 U12872 ( .A1(n11157), .A2(n3081), .ZN(n13095) );
  NAND3_X1 U12873 ( .A1(n37750), .A2(n36251), .A3(n37759), .ZN(n35925) );
  NAND2_X1 U12874 ( .A1(n3082), .A2(n36408), .ZN(n35997) );
  AOI21_X1 U12875 ( .B1(n5722), .B2(n3082), .A(n37648), .ZN(n35203) );
  NAND2_X1 U12876 ( .A1(n37644), .A2(n36397), .ZN(n3082) );
  OAI21_X1 U12877 ( .B1(n19705), .B2(n19834), .A(n19704), .ZN(n3086) );
  NAND3_X1 U12879 ( .A1(n3090), .A2(n21171), .A3(n21188), .ZN(n3089) );
  NAND3_X1 U12880 ( .A1(n40195), .A2(n3092), .A3(n3091), .ZN(n39559) );
  NAND2_X1 U12881 ( .A1(n40124), .A2(n40110), .ZN(n3091) );
  MUX2_X1 U12883 ( .A(n32128), .B(n26315), .S(n32125), .Z(n26328) );
  NAND2_X1 U12885 ( .A1(n29974), .A2(n3097), .ZN(n29981) );
  NAND2_X1 U12886 ( .A1(n32125), .A2(n721), .ZN(n3097) );
  MUX2_X1 U12887 ( .A(n32122), .B(n32123), .S(n32125), .Z(n32141) );
  NOR2_X1 U12890 ( .A1(n52433), .A2(n3100), .ZN(n24282) );
  OAI21_X1 U12891 ( .B1(n23509), .B2(n23511), .A(n3100), .ZN(n23515) );
  NOR2_X1 U12892 ( .A1(n21896), .A2(n3100), .ZN(n21897) );
  OR2_X1 U12893 ( .A1(n25858), .A2(n5912), .ZN(n3101) );
  NAND3_X1 U12894 ( .A1(n31879), .A2(n31876), .A3(n3101), .ZN(n30119) );
  INV_X1 U12896 ( .A(n31876), .ZN(n3104) );
  AND2_X1 U12897 ( .A1(n26677), .A2(n26679), .ZN(n3105) );
  NAND3_X1 U12899 ( .A1(n2294), .A2(n26677), .A3(n27859), .ZN(n29484) );
  NAND2_X1 U12900 ( .A1(n46714), .A2(n46595), .ZN(n3106) );
  INV_X1 U12901 ( .A(n45790), .ZN(n46710) );
  XNOR2_X1 U12902 ( .A(n52100), .B(n3111), .ZN(n28383) );
  XNOR2_X1 U12903 ( .A(n3112), .B(n52100), .ZN(n28055) );
  XNOR2_X1 U12904 ( .A(n52100), .B(n2547), .ZN(n26361) );
  XNOR2_X1 U12905 ( .A(n52100), .B(n2546), .ZN(n24012) );
  NAND2_X1 U12906 ( .A1(n3114), .A2(n32537), .ZN(n34504) );
  INV_X1 U12907 ( .A(n22251), .ZN(n23322) );
  NAND2_X1 U12908 ( .A1(n3115), .A2(n23320), .ZN(n3118) );
  NAND3_X2 U12912 ( .A1(n3118), .A2(n6133), .A3(n3119), .ZN(n25889) );
  NAND2_X1 U12913 ( .A1(n22255), .A2(n23310), .ZN(n3120) );
  INV_X1 U12914 ( .A(n52047), .ZN(n31019) );
  NAND2_X1 U12915 ( .A1(n31876), .A2(n31870), .ZN(n3123) );
  INV_X1 U12916 ( .A(n37377), .ZN(n3126) );
  NAND2_X1 U12918 ( .A1(n3127), .A2(n3126), .ZN(n3130) );
  NAND2_X1 U12919 ( .A1(n37376), .A2(n37597), .ZN(n3127) );
  NAND2_X1 U12920 ( .A1(n3129), .A2(n37377), .ZN(n3128) );
  AOI21_X1 U12921 ( .B1(n37365), .B2(n37366), .A(n1006), .ZN(n37370) );
  NAND2_X1 U12922 ( .A1(n31297), .A2(n3131), .ZN(n3133) );
  INV_X1 U12923 ( .A(n30652), .ZN(n3131) );
  NAND4_X2 U12924 ( .A1(n3134), .A2(n3133), .A3(n29654), .A4(n3132), .ZN(
        n37318) );
  OAI21_X1 U12925 ( .B1(n29653), .B2(n29396), .A(n30643), .ZN(n3132) );
  NAND3_X1 U12926 ( .A1(n29651), .A2(n31313), .A3(n3135), .ZN(n3134) );
  NAND2_X1 U12927 ( .A1(n30640), .A2(n31298), .ZN(n3135) );
  NAND3_X1 U12928 ( .A1(n3138), .A2(n3137), .A3(n32119), .ZN(n3136) );
  NAND2_X1 U12929 ( .A1(n29975), .A2(n30814), .ZN(n3137) );
  NAND2_X1 U12930 ( .A1(n30816), .A2(n29975), .ZN(n3138) );
  XNOR2_X2 U12931 ( .A(n16488), .B(n16487), .ZN(n20114) );
  INV_X1 U12932 ( .A(n26640), .ZN(n26639) );
  NAND2_X1 U12933 ( .A1(n26065), .A2(n27835), .ZN(n26640) );
  NAND2_X1 U12934 ( .A1(n3140), .A2(n14338), .ZN(n14350) );
  NAND2_X1 U12935 ( .A1(n14336), .A2(n3141), .ZN(n3140) );
  NAND2_X1 U12936 ( .A1(n6073), .A2(n14337), .ZN(n3141) );
  NAND2_X1 U12937 ( .A1(n13425), .A2(n14341), .ZN(n14336) );
  INV_X2 U12938 ( .A(n10639), .ZN(n13425) );
  XNOR2_X1 U12939 ( .A(n18592), .B(n3142), .ZN(n15995) );
  XNOR2_X1 U12940 ( .A(n16388), .B(n3142), .ZN(n16389) );
  XNOR2_X1 U12941 ( .A(n3142), .B(n18605), .ZN(n15028) );
  XNOR2_X1 U12942 ( .A(n16483), .B(n3142), .ZN(n16484) );
  XNOR2_X1 U12943 ( .A(n16766), .B(n3142), .ZN(n18458) );
  XNOR2_X1 U12944 ( .A(n14377), .B(n3142), .ZN(n15617) );
  XNOR2_X2 U12945 ( .A(n44918), .B(n44917), .ZN(n45848) );
  NAND2_X1 U12947 ( .A1(n27132), .A2(n3143), .ZN(n28894) );
  NAND2_X1 U12948 ( .A1(n27119), .A2(n3143), .ZN(n27993) );
  AND2_X1 U12949 ( .A1(n27119), .A2(n28897), .ZN(n26478) );
  NAND3_X1 U12951 ( .A1(n48760), .A2(n3145), .A3(n3144), .ZN(n46429) );
  NAND2_X2 U12952 ( .A1(n6554), .A2(n24420), .ZN(n25554) );
  NAND2_X1 U12953 ( .A1(n4725), .A2(n24111), .ZN(n24115) );
  NAND2_X1 U12954 ( .A1(n40635), .A2(n3146), .ZN(n4308) );
  NAND3_X1 U12955 ( .A1(n43670), .A2(n3148), .A3(n3147), .ZN(n3146) );
  NAND2_X1 U12956 ( .A1(n43667), .A2(n43665), .ZN(n3147) );
  NAND3_X1 U12957 ( .A1(n41799), .A2(n51684), .A3(n42109), .ZN(n43670) );
  INV_X1 U12958 ( .A(n31881), .ZN(n3152) );
  NAND2_X1 U12959 ( .A1(n31798), .A2(n31028), .ZN(n31881) );
  NAND2_X1 U12960 ( .A1(n3151), .A2(n3150), .ZN(n30132) );
  NAND2_X1 U12961 ( .A1(n30119), .A2(n30118), .ZN(n3150) );
  NAND2_X1 U12963 ( .A1(n29238), .A2(n29242), .ZN(n3154) );
  INV_X1 U12964 ( .A(n46597), .ZN(n3155) );
  NAND3_X1 U12965 ( .A1(n44838), .A2(n46583), .A3(n46701), .ZN(n44839) );
  NAND2_X1 U12966 ( .A1(n38312), .A2(n38728), .ZN(n3156) );
  INV_X1 U12967 ( .A(n26458), .ZN(n3160) );
  NAND2_X1 U12968 ( .A1(n29015), .A2(n3159), .ZN(n3161) );
  NAND2_X1 U12969 ( .A1(n28923), .A2(n29006), .ZN(n26459) );
  NAND2_X1 U12970 ( .A1(n28916), .A2(n28926), .ZN(n29006) );
  NAND2_X1 U12971 ( .A1(n3162), .A2(n21473), .ZN(n7994) );
  NAND2_X1 U12972 ( .A1(n19353), .A2(n2398), .ZN(n3162) );
  NAND2_X1 U12973 ( .A1(n19351), .A2(n19357), .ZN(n19353) );
  NAND2_X1 U12975 ( .A1(n23048), .A2(n23052), .ZN(n22944) );
  NAND2_X1 U12976 ( .A1(n5876), .A2(n33649), .ZN(n37403) );
  INV_X1 U12977 ( .A(n37396), .ZN(n3164) );
  INV_X1 U12978 ( .A(n37403), .ZN(n37539) );
  NAND2_X1 U12979 ( .A1(n3164), .A2(n525), .ZN(n3165) );
  NAND2_X1 U12980 ( .A1(n20648), .A2(n20647), .ZN(n3167) );
  OAI22_X1 U12981 ( .A1(n8349), .A2(n12051), .B1(n12059), .B2(n3168), .ZN(
        n12044) );
  NAND2_X1 U12982 ( .A1(n5307), .A2(n10664), .ZN(n6019) );
  OAI211_X1 U12983 ( .C1(n12046), .C2(n3168), .A(n9386), .B(n9385), .ZN(n9387)
         );
  NOR2_X1 U12986 ( .A1(n3174), .A2(n3171), .ZN(n3175) );
  NAND2_X1 U12987 ( .A1(n3173), .A2(n3172), .ZN(n3171) );
  NAND2_X1 U12988 ( .A1(n24185), .A2(n23766), .ZN(n3172) );
  NAND2_X1 U12989 ( .A1(n23767), .A2(n24190), .ZN(n3173) );
  NAND2_X1 U12990 ( .A1(n23204), .A2(n23205), .ZN(n3174) );
  NAND4_X1 U12991 ( .A1(n6940), .A2(n40617), .A3(n41985), .A4(n41645), .ZN(
        n5933) );
  OR2_X2 U12992 ( .A1(n34809), .A2(n34808), .ZN(n41645) );
  NOR2_X1 U12993 ( .A1(n12516), .A2(n8024), .ZN(n8023) );
  OAI21_X1 U12994 ( .B1(n20375), .B2(n21389), .A(n20408), .ZN(n20798) );
  OR2_X1 U12995 ( .A1(n20795), .A2(n20376), .ZN(n20408) );
  OAI21_X1 U12996 ( .B1(n19045), .B2(n19544), .A(n20123), .ZN(n17101) );
  NAND2_X1 U12997 ( .A1(n30528), .A2(n51740), .ZN(n3179) );
  NAND2_X1 U12998 ( .A1(n3486), .A2(n3176), .ZN(n3485) );
  NAND2_X1 U12999 ( .A1(n30528), .A2(n3177), .ZN(n3176) );
  OAI21_X1 U13001 ( .B1(n31380), .B2(n33017), .A(n3179), .ZN(n6758) );
  NAND2_X1 U13002 ( .A1(n3180), .A2(n2519), .ZN(n23384) );
  NAND2_X1 U13005 ( .A1(n10469), .A2(n3183), .ZN(n3182) );
  NAND2_X1 U13006 ( .A1(n10464), .A2(n51432), .ZN(n3183) );
  NAND2_X1 U13007 ( .A1(n10470), .A2(n3185), .ZN(n3184) );
  NAND2_X1 U13008 ( .A1(n8718), .A2(n10463), .ZN(n3185) );
  INV_X1 U13009 ( .A(n20201), .ZN(n3189) );
  INV_X1 U13010 ( .A(n20638), .ZN(n21543) );
  NAND2_X1 U13011 ( .A1(n21533), .A2(n3188), .ZN(n20631) );
  NAND2_X1 U13012 ( .A1(n46699), .A2(n46700), .ZN(n46706) );
  OR2_X1 U13013 ( .A1(n46707), .A2(n46580), .ZN(n46700) );
  AND3_X2 U13016 ( .A1(n3193), .A2(n3190), .A3(n6021), .ZN(n23160) );
  NAND2_X1 U13017 ( .A1(n16213), .A2(n20076), .ZN(n3192) );
  NOR2_X1 U13018 ( .A1(n3196), .A2(n3194), .ZN(n3193) );
  OAI22_X1 U13019 ( .A1(n19498), .A2(n3195), .B1(n19138), .B2(n20075), .ZN(
        n3194) );
  NAND2_X1 U13020 ( .A1(n19491), .A2(n19494), .ZN(n20065) );
  NOR2_X1 U13021 ( .A1(n51478), .A2(n52137), .ZN(n48976) );
  NAND2_X1 U13024 ( .A1(n48937), .A2(n2439), .ZN(n47483) );
  NAND4_X1 U13025 ( .A1(n47476), .A2(n48971), .A3(n48972), .A4(n52137), .ZN(
        n48979) );
  NOR2_X1 U13026 ( .A1(n24351), .A2(n738), .ZN(n3200) );
  NAND2_X1 U13027 ( .A1(n51697), .A2(n29924), .ZN(n26843) );
  NAND2_X1 U13028 ( .A1(n51696), .A2(n3200), .ZN(n24349) );
  NAND3_X1 U13029 ( .A1(n27556), .A2(n3201), .A3(n24349), .ZN(n30767) );
  NAND2_X1 U13030 ( .A1(n30767), .A2(n30766), .ZN(n30778) );
  NAND3_X1 U13031 ( .A1(n30801), .A2(n3204), .A3(n3203), .ZN(n3202) );
  NAND2_X1 U13032 ( .A1(n31168), .A2(n381), .ZN(n3203) );
  NAND3_X1 U13033 ( .A1(n30802), .A2(n32669), .A3(n32662), .ZN(n3204) );
  NAND3_X1 U13034 ( .A1(n47484), .A2(n46954), .A3(n48960), .ZN(n3205) );
  AND2_X1 U13035 ( .A1(n3205), .A2(n47485), .ZN(n3206) );
  NAND2_X1 U13038 ( .A1(n3209), .A2(n48957), .ZN(n48931) );
  NAND2_X1 U13039 ( .A1(n46945), .A2(n3210), .ZN(n46946) );
  NAND3_X1 U13041 ( .A1(n37571), .A2(n3211), .A3(n37576), .ZN(n35697) );
  NAND2_X1 U13042 ( .A1(n38593), .A2(n35693), .ZN(n37453) );
  AND3_X1 U13043 ( .A1(n49454), .A2(n49437), .A3(n49439), .ZN(n3219) );
  NAND3_X1 U13044 ( .A1(n3216), .A2(n3215), .A3(n3212), .ZN(Plaintext[111]) );
  NAND4_X1 U13045 ( .A1(n3214), .A2(n3213), .A3(n49453), .A4(n3219), .ZN(n3212) );
  NOR2_X1 U13046 ( .A1(n3220), .A2(n49455), .ZN(n3213) );
  INV_X1 U13047 ( .A(n3221), .ZN(n3214) );
  NAND2_X1 U13048 ( .A1(n3221), .A2(n49455), .ZN(n3215) );
  INV_X1 U13053 ( .A(n5083), .ZN(n3222) );
  INV_X1 U13054 ( .A(n5083), .ZN(n19846) );
  NAND2_X1 U13055 ( .A1(n22736), .A2(n753), .ZN(n5094) );
  OR2_X2 U13056 ( .A1(n19743), .A2(n5093), .ZN(n22736) );
  NAND2_X1 U13057 ( .A1(n22146), .A2(n22142), .ZN(n3223) );
  INV_X1 U13058 ( .A(n3223), .ZN(n19568) );
  NAND3_X1 U13059 ( .A1(n3223), .A2(n21024), .A3(n50992), .ZN(n17611) );
  NAND2_X1 U13060 ( .A1(n3225), .A2(n30102), .ZN(n3790) );
  NAND2_X1 U13061 ( .A1(n722), .A2(n3226), .ZN(n30107) );
  INV_X1 U13062 ( .A(n5913), .ZN(n3226) );
  NOR2_X1 U13063 ( .A1(n722), .A2(n621), .ZN(n31492) );
  AOI22_X1 U13064 ( .A1(n30991), .A2(n30992), .B1(n31483), .B2(n621), .ZN(
        n31002) );
  MUX2_X1 U13065 ( .A(n31267), .B(n31268), .S(n30102), .Z(n31279) );
  NAND2_X1 U13066 ( .A1(n19871), .A2(n19639), .ZN(n3227) );
  INV_X1 U13068 ( .A(n19853), .ZN(n19847) );
  INV_X1 U13069 ( .A(n19871), .ZN(n19863) );
  NAND2_X1 U13070 ( .A1(n45216), .A2(n45215), .ZN(n3229) );
  OAI21_X1 U13071 ( .B1(n45640), .B2(n46239), .A(n3229), .ZN(n45641) );
  NOR2_X1 U13072 ( .A1(n38832), .A2(n52094), .ZN(n3231) );
  OR2_X1 U13073 ( .A1(n39759), .A2(n39942), .ZN(n39114) );
  NAND2_X1 U13074 ( .A1(n37856), .A2(n52073), .ZN(n39759) );
  XNOR2_X1 U13075 ( .A(n28083), .B(n27443), .ZN(n3232) );
  INV_X1 U13076 ( .A(n30431), .ZN(n3233) );
  NAND3_X2 U13077 ( .A1(n3235), .A2(n51780), .A3(n23648), .ZN(n3236) );
  OR2_X1 U13078 ( .A1(n23650), .A2(n23649), .ZN(n3235) );
  XNOR2_X2 U13079 ( .A(n3236), .B(n23651), .ZN(n27439) );
  XNOR2_X1 U13080 ( .A(n3236), .B(n47679), .ZN(n26234) );
  XNOR2_X1 U13081 ( .A(n3236), .B(n28214), .ZN(n28341) );
  XNOR2_X1 U13082 ( .A(n3236), .B(n25760), .ZN(n25761) );
  NAND2_X1 U13083 ( .A1(n32729), .A2(n32732), .ZN(n3237) );
  NOR2_X1 U13085 ( .A1(n32457), .A2(n32717), .ZN(n3238) );
  NAND2_X1 U13086 ( .A1(n32457), .A2(n31648), .ZN(n3239) );
  NAND2_X1 U13087 ( .A1(n3240), .A2(n31578), .ZN(n30864) );
  INV_X1 U13089 ( .A(n20698), .ZN(n19981) );
  XNOR2_X2 U13090 ( .A(n15963), .B(n15962), .ZN(n20698) );
  INV_X1 U13091 ( .A(n21618), .ZN(n20253) );
  NAND2_X1 U13092 ( .A1(n21630), .A2(n19981), .ZN(n21618) );
  INV_X1 U13093 ( .A(n51050), .ZN(n20615) );
  INV_X1 U13094 ( .A(n20188), .ZN(n18898) );
  NAND2_X1 U13095 ( .A1(n5409), .A2(n3244), .ZN(n5536) );
  AND2_X1 U13096 ( .A1(n18895), .A2(n3245), .ZN(n3244) );
  NAND2_X1 U13097 ( .A1(n51050), .A2(n21513), .ZN(n3245) );
  NAND2_X1 U13098 ( .A1(n18894), .A2(n18903), .ZN(n5409) );
  NAND3_X1 U13099 ( .A1(n6528), .A2(n49162), .A3(n6527), .ZN(n3247) );
  INV_X1 U13100 ( .A(n37976), .ZN(n3248) );
  NAND2_X1 U13102 ( .A1(n3249), .A2(n11591), .ZN(n11595) );
  INV_X1 U13103 ( .A(n16039), .ZN(n14527) );
  NAND2_X1 U13104 ( .A1(n16039), .A2(n13377), .ZN(n13036) );
  NAND3_X2 U13105 ( .A1(n7965), .A2(n7966), .A3(n11638), .ZN(n13377) );
  NAND2_X1 U13106 ( .A1(n37191), .A2(n3251), .ZN(n38339) );
  NAND2_X2 U13107 ( .A1(n36468), .A2(n3251), .ZN(n38330) );
  NAND2_X1 U13108 ( .A1(n41332), .A2(n40730), .ZN(n39821) );
  NAND4_X1 U13109 ( .A1(n41317), .A2(n41332), .A3(n41319), .A4(n40730), .ZN(
        n40725) );
  NAND2_X1 U13110 ( .A1(n3252), .A2(n41318), .ZN(n39631) );
  AOI22_X1 U13111 ( .A1(n13650), .A2(n12754), .B1(n3253), .B2(n12753), .ZN(
        n12761) );
  NAND2_X1 U13112 ( .A1(n12753), .A2(n14642), .ZN(n13651) );
  NOR2_X1 U13113 ( .A1(n3254), .A2(n13667), .ZN(n3253) );
  NAND2_X1 U13114 ( .A1(n35889), .A2(n35407), .ZN(n35893) );
  INV_X1 U13115 ( .A(n35890), .ZN(n3255) );
  NOR2_X1 U13116 ( .A1(n35889), .A2(n3257), .ZN(n3256) );
  INV_X1 U13117 ( .A(n36468), .ZN(n3257) );
  NAND3_X1 U13119 ( .A1(n3284), .A2(n19292), .A3(n19291), .ZN(n19300) );
  INV_X1 U13120 ( .A(n14761), .ZN(n15205) );
  NAND3_X2 U13122 ( .A1(n3259), .A2(n29540), .A3(n29538), .ZN(n30931) );
  AOI21_X1 U13123 ( .B1(n32905), .B2(n32906), .A(n32904), .ZN(n32927) );
  INV_X1 U13124 ( .A(n29512), .ZN(n29528) );
  NOR2_X1 U13125 ( .A1(n33029), .A2(n33040), .ZN(n3264) );
  NAND2_X1 U13126 ( .A1(n3260), .A2(n14103), .ZN(n14433) );
  OAI21_X1 U13128 ( .B1(n28018), .B2(n28017), .A(n28194), .ZN(n7336) );
  INV_X1 U13129 ( .A(n14438), .ZN(n4358) );
  NAND3_X1 U13130 ( .A1(n30049), .A2(n30047), .A3(n30048), .ZN(n30050) );
  NAND2_X1 U13131 ( .A1(n37649), .A2(n3261), .ZN(n37650) );
  NAND2_X1 U13133 ( .A1(n2370), .A2(n9516), .ZN(n3583) );
  NAND2_X1 U13134 ( .A1(n19567), .A2(n21018), .ZN(n3425) );
  NAND2_X1 U13136 ( .A1(n14445), .A2(n3263), .ZN(n3262) );
  NOR2_X1 U13137 ( .A1(n3264), .A2(n2485), .ZN(n3294) );
  NAND2_X1 U13139 ( .A1(n30186), .A2(n3265), .ZN(n30310) );
  NAND3_X1 U13140 ( .A1(n23198), .A2(n23197), .A3(n23199), .ZN(n3266) );
  NAND2_X1 U13141 ( .A1(n41111), .A2(n41123), .ZN(n40476) );
  AND4_X2 U13142 ( .A1(n36916), .A2(n36914), .A3(n36913), .A4(n36915), .ZN(
        n41111) );
  XNOR2_X2 U13144 ( .A(n34758), .B(n34757), .ZN(n39438) );
  NAND2_X1 U13145 ( .A1(n14871), .A2(n14880), .ZN(n13881) );
  INV_X1 U13146 ( .A(Ciphertext[11]), .ZN(n8656) );
  OAI21_X1 U13147 ( .B1(n9149), .B2(n3267), .A(n11204), .ZN(n7486) );
  NOR2_X1 U13148 ( .A1(n11211), .A2(n11198), .ZN(n3267) );
  NOR2_X1 U13151 ( .A1(n16891), .A2(n16890), .ZN(n3268) );
  NOR2_X1 U13152 ( .A1(n353), .A2(n22390), .ZN(n3269) );
  NAND2_X2 U13155 ( .A1(n4241), .A2(n6501), .ZN(n22983) );
  NOR2_X2 U13156 ( .A1(n11587), .A2(n11586), .ZN(n11723) );
  OAI21_X1 U13157 ( .B1(n30022), .B2(n29998), .A(n3272), .ZN(n26796) );
  NAND2_X1 U13158 ( .A1(n2237), .A2(n30004), .ZN(n3272) );
  NOR2_X1 U13160 ( .A1(n31342), .A2(n5682), .ZN(n3273) );
  NAND2_X1 U13161 ( .A1(n22434), .A2(n22985), .ZN(n3274) );
  NAND2_X1 U13162 ( .A1(n23002), .A2(n22982), .ZN(n3275) );
  NAND2_X1 U13163 ( .A1(n7007), .A2(n7006), .ZN(n24363) );
  NAND3_X1 U13165 ( .A1(n35454), .A2(n35455), .A3(n35456), .ZN(n35463) );
  AND2_X1 U13166 ( .A1(n40564), .A2(n40556), .ZN(n40314) );
  INV_X1 U13167 ( .A(n32486), .ZN(n32489) );
  XOR2_X1 U13168 ( .A(n36951), .B(n33185), .Z(n6902) );
  INV_X1 U13169 ( .A(n31778), .ZN(n32244) );
  NAND2_X1 U13170 ( .A1(n20817), .A2(n20813), .ZN(n19283) );
  NAND3_X1 U13171 ( .A1(n38213), .A2(n38557), .A3(n38543), .ZN(n31356) );
  NAND4_X1 U13172 ( .A1(n31445), .A2(n30800), .A3(n30806), .A4(n30807), .ZN(
        n7242) );
  OAI211_X1 U13173 ( .C1(n30997), .C2(n3785), .A(n31484), .B(n30990), .ZN(
        n3784) );
  NAND2_X1 U13174 ( .A1(n41934), .A2(n3277), .ZN(n7305) );
  NAND2_X1 U13175 ( .A1(n40249), .A2(n41938), .ZN(n3277) );
  NAND2_X1 U13176 ( .A1(n49597), .A2(n49596), .ZN(n6006) );
  NAND4_X1 U13177 ( .A1(n49590), .A2(n49589), .A3(n49588), .A4(n49587), .ZN(
        n49597) );
  NAND2_X1 U13178 ( .A1(n32877), .A2(n8544), .ZN(n33029) );
  NAND2_X1 U13179 ( .A1(n14783), .A2(n14784), .ZN(n14785) );
  NOR2_X1 U13180 ( .A1(n12246), .A2(n2406), .ZN(n8995) );
  INV_X1 U13181 ( .A(n30695), .ZN(n6256) );
  NAND2_X1 U13182 ( .A1(n11908), .A2(n11484), .ZN(n12491) );
  NAND3_X1 U13183 ( .A1(n7487), .A2(n6517), .A3(n32603), .ZN(n6518) );
  NAND4_X2 U13187 ( .A1(n17029), .A2(n17034), .A3(n17030), .A4(n17028), .ZN(
        n23568) );
  NAND3_X1 U13188 ( .A1(n37418), .A2(n37419), .A3(n38120), .ZN(n4571) );
  NAND3_X1 U13189 ( .A1(n6669), .A2(n50336), .A3(n50337), .ZN(n50340) );
  NAND2_X1 U13190 ( .A1(n37977), .A2(n37983), .ZN(n3281) );
  NAND2_X1 U13191 ( .A1(n36521), .A2(n37980), .ZN(n36527) );
  OAI21_X1 U13192 ( .B1(n38779), .B2(n38780), .A(n584), .ZN(n38790) );
  NAND3_X1 U13194 ( .A1(n26890), .A2(n27631), .A3(n3282), .ZN(n8274) );
  NOR2_X1 U13195 ( .A1(n21359), .A2(n19289), .ZN(n19286) );
  NAND2_X1 U13196 ( .A1(n21603), .A2(n21605), .ZN(n21359) );
  BUF_X2 U13197 ( .A(n47435), .Z(n48778) );
  NAND3_X1 U13198 ( .A1(n46343), .A2(n45687), .A3(n3283), .ZN(n45692) );
  NAND3_X1 U13199 ( .A1(n2495), .A2(n5890), .A3(n3285), .ZN(n5887) );
  INV_X1 U13200 ( .A(n48915), .ZN(n3285) );
  NAND2_X1 U13201 ( .A1(n12313), .A2(n12315), .ZN(n12309) );
  NAND2_X1 U13202 ( .A1(n20227), .A2(n20677), .ZN(n5463) );
  INV_X1 U13203 ( .A(n38555), .ZN(n35177) );
  NAND2_X1 U13204 ( .A1(n35175), .A2(n38550), .ZN(n38555) );
  OAI21_X1 U13207 ( .B1(n38092), .B2(n36629), .A(n6904), .ZN(n36318) );
  NAND2_X1 U13208 ( .A1(n3287), .A2(n23811), .ZN(n3286) );
  NAND2_X1 U13209 ( .A1(n22298), .A2(n5371), .ZN(n3287) );
  NAND2_X1 U13210 ( .A1(n20575), .A2(n22736), .ZN(n3288) );
  NAND2_X1 U13211 ( .A1(n13556), .A2(n3289), .ZN(n13557) );
  NAND2_X1 U13212 ( .A1(n29324), .A2(n29330), .ZN(n27821) );
  NAND2_X1 U13214 ( .A1(n40294), .A2(n42061), .ZN(n41491) );
  XNOR2_X1 U13215 ( .A(n3291), .B(n45986), .ZN(Plaintext[113]) );
  NAND3_X1 U13216 ( .A1(n45983), .A2(n3299), .A3(n45985), .ZN(n3291) );
  INV_X1 U13217 ( .A(n12821), .ZN(n3292) );
  NAND2_X1 U13218 ( .A1(n46881), .A2(n47106), .ZN(n46568) );
  NAND2_X1 U13219 ( .A1(n33035), .A2(n33036), .ZN(n33037) );
  NOR2_X1 U13220 ( .A1(n27841), .A2(n7825), .ZN(n27843) );
  AND2_X1 U13221 ( .A1(n31416), .A2(n31415), .ZN(n5635) );
  AND2_X1 U13222 ( .A1(n3731), .A2(n14931), .ZN(n3730) );
  NAND4_X2 U13223 ( .A1(n3293), .A2(n3294), .A3(n33028), .A4(n33043), .ZN(
        n33303) );
  NAND2_X1 U13224 ( .A1(n51063), .A2(n39224), .ZN(n39221) );
  NAND2_X1 U13225 ( .A1(n3978), .A2(n38054), .ZN(n3977) );
  AND3_X1 U13226 ( .A1(n20032), .A2(n18373), .A3(n51440), .ZN(n7580) );
  INV_X1 U13227 ( .A(n13449), .ZN(n3552) );
  NAND2_X1 U13228 ( .A1(n38298), .A2(n3874), .ZN(n39227) );
  NAND2_X1 U13229 ( .A1(n38887), .A2(n40967), .ZN(n41377) );
  AOI21_X1 U13230 ( .B1(n7499), .B2(n41247), .A(n41679), .ZN(n3860) );
  NAND4_X2 U13231 ( .A1(n39750), .A2(n39965), .A3(n39749), .A4(n39748), .ZN(
        n44561) );
  NAND2_X1 U13233 ( .A1(n18472), .A2(n21547), .ZN(n3295) );
  NAND3_X1 U13234 ( .A1(n2361), .A2(n14535), .A3(n3296), .ZN(n14539) );
  NAND2_X1 U13235 ( .A1(n14534), .A2(n14533), .ZN(n3296) );
  NAND2_X1 U13236 ( .A1(n20308), .A2(n417), .ZN(n3297) );
  NAND2_X1 U13237 ( .A1(n20307), .A2(n23230), .ZN(n3298) );
  NAND3_X2 U13238 ( .A1(n8255), .A2(n23770), .A3(n23771), .ZN(n26159) );
  INV_X1 U13239 ( .A(n28979), .ZN(n3301) );
  INV_X1 U13240 ( .A(n30768), .ZN(n3302) );
  NOR2_X1 U13241 ( .A1(n39422), .A2(n39206), .ZN(n39205) );
  NAND2_X1 U13242 ( .A1(n32962), .A2(n32767), .ZN(n32770) );
  NAND2_X1 U13243 ( .A1(n51374), .A2(n18040), .ZN(n18034) );
  NAND3_X1 U13244 ( .A1(n47589), .A2(n47618), .A3(n47617), .ZN(n47590) );
  NAND3_X1 U13245 ( .A1(n7679), .A2(n46585), .A3(n46582), .ZN(n3304) );
  NAND3_X1 U13246 ( .A1(n4777), .A2(n40779), .A3(n40780), .ZN(n40790) );
  NAND3_X1 U13247 ( .A1(n3305), .A2(n11951), .A3(n11950), .ZN(n11952) );
  NAND3_X1 U13248 ( .A1(n11949), .A2(n11948), .A3(n8882), .ZN(n3305) );
  NAND2_X1 U13249 ( .A1(n23703), .A2(n3306), .ZN(n24328) );
  NOR2_X1 U13250 ( .A1(n7361), .A2(n15437), .ZN(n8663) );
  NAND2_X1 U13253 ( .A1(n3309), .A2(n23464), .ZN(n23476) );
  NAND2_X1 U13254 ( .A1(n3310), .A2(n23463), .ZN(n3309) );
  NAND2_X1 U13255 ( .A1(n16688), .A2(n51123), .ZN(n23463) );
  INV_X1 U13256 ( .A(n23465), .ZN(n3310) );
  NAND2_X1 U13257 ( .A1(n3994), .A2(n3991), .ZN(n3415) );
  NAND4_X2 U13258 ( .A1(n46039), .A2(n7569), .A3(n7566), .A4(n46038), .ZN(
        n49916) );
  AOI21_X1 U13259 ( .B1(n21781), .B2(n51695), .A(n4225), .ZN(n21784) );
  OAI21_X1 U13260 ( .B1(n31281), .B2(n32409), .A(n4850), .ZN(n31293) );
  INV_X1 U13261 ( .A(n3312), .ZN(n21240) );
  OAI211_X1 U13262 ( .C1(n21231), .C2(n21230), .A(n21228), .B(n21229), .ZN(
        n3312) );
  NAND3_X1 U13263 ( .A1(n37204), .A2(n39016), .A3(n37203), .ZN(n37206) );
  NAND2_X1 U13264 ( .A1(n6651), .A2(n19052), .ZN(n3314) );
  OAI21_X1 U13265 ( .B1(n40622), .B2(n34919), .A(n41975), .ZN(n8109) );
  NOR2_X1 U13266 ( .A1(n31219), .A2(n31763), .ZN(n31776) );
  OAI21_X1 U13267 ( .B1(n26074), .B2(n29295), .A(n28686), .ZN(n26088) );
  XNOR2_X2 U13268 ( .A(n33669), .B(n33670), .ZN(n36272) );
  INV_X1 U13269 ( .A(n7378), .ZN(n6941) );
  NOR2_X1 U13270 ( .A1(n29465), .A2(n29456), .ZN(n5276) );
  INV_X1 U13271 ( .A(n19510), .ZN(n16677) );
  NAND2_X1 U13272 ( .A1(n8735), .A2(n29537), .ZN(n29538) );
  AND2_X1 U13273 ( .A1(n9923), .A2(n4006), .ZN(n8177) );
  INV_X1 U13274 ( .A(n28623), .ZN(n29526) );
  INV_X1 U13275 ( .A(n17418), .ZN(n23080) );
  XNOR2_X1 U13277 ( .A(n3318), .B(n28080), .ZN(n28081) );
  XNOR2_X1 U13278 ( .A(n28079), .B(n28240), .ZN(n3318) );
  NAND2_X1 U13279 ( .A1(n3812), .A2(n32776), .ZN(n3319) );
  NAND2_X1 U13280 ( .A1(n23693), .A2(n23536), .ZN(n3821) );
  NAND4_X2 U13281 ( .A1(n20619), .A2(n20622), .A3(n20620), .A4(n20621), .ZN(
        n23535) );
  NAND4_X1 U13282 ( .A1(n47678), .A2(n3320), .A3(n47677), .A4(n5967), .ZN(
        n5965) );
  NAND2_X1 U13283 ( .A1(n49492), .A2(n2193), .ZN(n3321) );
  NAND2_X1 U13284 ( .A1(n3322), .A2(n49514), .ZN(n7017) );
  AOI21_X1 U13285 ( .B1(n22414), .B2(n22413), .A(n6311), .ZN(n6310) );
  NAND2_X1 U13286 ( .A1(n3323), .A2(n44837), .ZN(n6102) );
  NAND3_X1 U13287 ( .A1(n44836), .A2(n4394), .A3(n44835), .ZN(n3323) );
  INV_X1 U13288 ( .A(n40250), .ZN(n6617) );
  NAND2_X1 U13289 ( .A1(n3664), .A2(n32027), .ZN(n3663) );
  NAND3_X1 U13290 ( .A1(n44707), .A2(n51396), .A3(n44845), .ZN(n44709) );
  NAND3_X1 U13291 ( .A1(n11005), .A2(n10251), .A3(n10195), .ZN(n9028) );
  OAI22_X1 U13292 ( .A1(n45025), .A2(n49494), .B1(n49479), .B2(n3325), .ZN(
        n3900) );
  NAND3_X1 U13293 ( .A1(n45024), .A2(n49521), .A3(n49503), .ZN(n3325) );
  OAI21_X1 U13294 ( .B1(n40314), .B2(n52160), .A(n40570), .ZN(n40317) );
  NOR2_X1 U13295 ( .A1(n12119), .A2(n3326), .ZN(n12128) );
  NAND3_X1 U13296 ( .A1(n12115), .A2(n4166), .A3(n12116), .ZN(n3326) );
  OR2_X1 U13297 ( .A1(n28496), .A2(n28953), .ZN(n28954) );
  NAND2_X1 U13298 ( .A1(n29794), .A2(n3827), .ZN(n28496) );
  OR2_X1 U13299 ( .A1(n46591), .A2(n51317), .ZN(n44706) );
  NAND3_X1 U13300 ( .A1(n48231), .A2(n48230), .A3(n3327), .ZN(n48232) );
  OR2_X1 U13301 ( .A1(n48550), .A2(n48239), .ZN(n3327) );
  NAND2_X1 U13302 ( .A1(n48238), .A2(n3328), .ZN(n48230) );
  NAND2_X1 U13303 ( .A1(n23112), .A2(n27158), .ZN(n30724) );
  NAND2_X2 U13304 ( .A1(n3329), .A2(n6842), .ZN(n12907) );
  INV_X1 U13305 ( .A(n21377), .ZN(n20410) );
  NOR2_X1 U13307 ( .A1(n23395), .A2(n8524), .ZN(n22108) );
  NAND2_X1 U13308 ( .A1(n35027), .A2(n3332), .ZN(n38181) );
  NAND2_X1 U13309 ( .A1(n5041), .A2(n20903), .ZN(n21318) );
  INV_X1 U13311 ( .A(n3334), .ZN(n19486) );
  AOI21_X1 U13312 ( .B1(n16306), .B2(n3335), .A(n21248), .ZN(n3334) );
  NAND2_X1 U13313 ( .A1(n17079), .A2(n16305), .ZN(n16306) );
  NAND2_X1 U13314 ( .A1(n3337), .A2(n20930), .ZN(n20937) );
  OAI21_X1 U13315 ( .B1(n20929), .B2(n21836), .A(n20928), .ZN(n3337) );
  NAND2_X1 U13316 ( .A1(n31482), .A2(n31483), .ZN(n31485) );
  NAND2_X1 U13321 ( .A1(n19122), .A2(n19023), .ZN(n3968) );
  NAND2_X1 U13322 ( .A1(n30792), .A2(n23658), .ZN(n3341) );
  NAND2_X1 U13323 ( .A1(n15425), .A2(n13874), .ZN(n13888) );
  INV_X1 U13324 ( .A(n19955), .ZN(n3342) );
  AOI22_X1 U13326 ( .A1(n29059), .A2(n30355), .B1(n29057), .B2(n29058), .ZN(
        n8189) );
  INV_X1 U13327 ( .A(n12435), .ZN(n12708) );
  OAI211_X1 U13328 ( .C1(n20650), .C2(n21654), .A(n21653), .B(n3343), .ZN(
        n15837) );
  NAND4_X2 U13330 ( .A1(n21347), .A2(n21348), .A3(n21346), .A4(n21345), .ZN(
        n25308) );
  NAND2_X1 U13331 ( .A1(n18903), .A2(n21521), .ZN(n21519) );
  AND2_X1 U13332 ( .A1(n14793), .A2(n14794), .ZN(n8342) );
  NAND2_X1 U13333 ( .A1(n10664), .A2(n11389), .ZN(n3805) );
  NOR2_X1 U13334 ( .A1(n8354), .A2(n19889), .ZN(n4470) );
  INV_X1 U13335 ( .A(n12073), .ZN(n4041) );
  AND3_X1 U13336 ( .A1(n19910), .A2(n19908), .A3(n19909), .ZN(n3346) );
  OR2_X1 U13337 ( .A1(n13346), .A2(n14534), .ZN(n13358) );
  XNOR2_X1 U13338 ( .A(n43774), .B(n46092), .ZN(n3653) );
  NAND2_X1 U13339 ( .A1(n11169), .A2(n3350), .ZN(n3349) );
  NAND3_X1 U13340 ( .A1(n36131), .A2(n36130), .A3(n36129), .ZN(n36140) );
  NAND3_X1 U13341 ( .A1(n32728), .A2(n32729), .A3(n32730), .ZN(n32734) );
  NAND2_X1 U13342 ( .A1(n35869), .A2(n2123), .ZN(n3352) );
  NAND2_X1 U13343 ( .A1(n5120), .A2(n11423), .ZN(n12133) );
  NAND2_X1 U13345 ( .A1(n3709), .A2(n38327), .ZN(n4253) );
  OAI211_X1 U13346 ( .C1(n47075), .C2(n46824), .A(n47071), .B(n46823), .ZN(
        n44452) );
  NAND2_X1 U13347 ( .A1(n47076), .A2(n45176), .ZN(n47071) );
  NOR2_X1 U13348 ( .A1(n438), .A2(n51141), .ZN(n11400) );
  AOI22_X1 U13350 ( .A1(n4071), .A2(n9531), .B1(n13076), .B2(n13105), .ZN(
        n9532) );
  NAND2_X1 U13353 ( .A1(n3354), .A2(n37637), .ZN(n36400) );
  OAI211_X1 U13354 ( .C1(n22503), .C2(n22228), .A(n22227), .B(n22226), .ZN(
        n22230) );
  NOR2_X1 U13355 ( .A1(n20213), .A2(n7857), .ZN(n7856) );
  NAND2_X1 U13356 ( .A1(n51734), .A2(n38805), .ZN(n41788) );
  NAND4_X4 U13357 ( .A1(n20108), .A2(n20106), .A3(n6722), .A4(n20107), .ZN(
        n23411) );
  NAND2_X1 U13358 ( .A1(n38717), .A2(n38718), .ZN(n3355) );
  OAI21_X1 U13360 ( .B1(n21989), .B2(n21990), .A(n21988), .ZN(n21992) );
  NAND2_X1 U13361 ( .A1(n23207), .A2(n412), .ZN(n23225) );
  NAND2_X1 U13362 ( .A1(n21349), .A2(n21350), .ZN(n21353) );
  AOI21_X1 U13364 ( .B1(n8348), .B2(n12047), .A(n3356), .ZN(n10366) );
  NAND2_X1 U13365 ( .A1(n32504), .A2(n32503), .ZN(n3358) );
  XNOR2_X1 U13367 ( .A(n8465), .B(n16576), .ZN(n5349) );
  INV_X1 U13369 ( .A(n50771), .ZN(n50779) );
  NOR2_X1 U13370 ( .A1(n7581), .A2(n7580), .ZN(n7579) );
  INV_X1 U13371 ( .A(n12601), .ZN(n11132) );
  INV_X1 U13372 ( .A(n7532), .ZN(n30251) );
  AOI21_X1 U13373 ( .B1(n18234), .B2(n19687), .A(n19671), .ZN(n3538) );
  XNOR2_X1 U13374 ( .A(n16782), .B(n8083), .ZN(n3472) );
  NAND2_X1 U13375 ( .A1(n45943), .A2(n3361), .ZN(n45947) );
  NAND2_X1 U13376 ( .A1(n29994), .A2(n29995), .ZN(n31150) );
  OR2_X1 U13378 ( .A1(n38005), .A2(n34971), .ZN(n35023) );
  INV_X1 U13379 ( .A(n41292), .ZN(n8291) );
  NAND4_X2 U13380 ( .A1(n9274), .A2(n9272), .A3(n9271), .A4(n9273), .ZN(n15677) );
  NAND3_X2 U13382 ( .A1(n7347), .A2(n7346), .A3(n19723), .ZN(n22375) );
  NAND2_X1 U13383 ( .A1(n27123), .A2(n28590), .ZN(n25300) );
  NAND2_X1 U13384 ( .A1(n47162), .A2(n8655), .ZN(n45156) );
  AND2_X1 U13385 ( .A1(n19296), .A2(n21362), .ZN(n3474) );
  NAND4_X2 U13386 ( .A1(n32451), .A2(n32456), .A3(n32450), .A4(n3362), .ZN(
        n36841) );
  NAND2_X1 U13387 ( .A1(n37158), .A2(n37924), .ZN(n38662) );
  NAND4_X2 U13388 ( .A1(n41397), .A2(n41398), .A3(n41396), .A4(n41399), .ZN(
        n45089) );
  NAND2_X1 U13389 ( .A1(n5480), .A2(n32616), .ZN(n3363) );
  OAI21_X1 U13390 ( .B1(n24417), .B2(n24418), .A(n24416), .ZN(n3364) );
  OR2_X1 U13391 ( .A1(n31463), .A2(n31558), .ZN(n6966) );
  NAND4_X2 U13392 ( .A1(n25302), .A2(n25303), .A3(n28890), .A4(n25304), .ZN(
        n32210) );
  INV_X1 U13393 ( .A(n23191), .ZN(n23746) );
  NAND4_X2 U13395 ( .A1(n38791), .A2(n38790), .A3(n38789), .A4(n51164), .ZN(
        n44534) );
  NAND2_X1 U13396 ( .A1(n41544), .A2(n40943), .ZN(n41389) );
  NAND4_X2 U13397 ( .A1(n23790), .A2(n6736), .A3(n23788), .A4(n23789), .ZN(
        n25483) );
  INV_X1 U13399 ( .A(n38959), .ZN(n7998) );
  NAND2_X1 U13401 ( .A1(n10047), .A2(n6005), .ZN(n7179) );
  NAND2_X1 U13402 ( .A1(n41791), .A2(n38810), .ZN(n42109) );
  NAND2_X2 U13403 ( .A1(n6685), .A2(n49228), .ZN(n49370) );
  NAND2_X1 U13404 ( .A1(n21459), .A2(n3366), .ZN(n6173) );
  XNOR2_X2 U13406 ( .A(n15788), .B(n15787), .ZN(n20270) );
  XNOR2_X1 U13407 ( .A(n46052), .B(n51337), .ZN(n3756) );
  XNOR2_X1 U13408 ( .A(n3757), .B(n3755), .ZN(n42945) );
  NAND2_X1 U13409 ( .A1(n30181), .A2(n1771), .ZN(n30172) );
  NAND2_X1 U13410 ( .A1(n20274), .A2(n3369), .ZN(n20268) );
  NAND3_X1 U13411 ( .A1(n31533), .A2(n32883), .A3(n32874), .ZN(n29077) );
  NAND2_X1 U13412 ( .A1(n40537), .A2(n40533), .ZN(n3372) );
  NAND2_X1 U13414 ( .A1(n21465), .A2(n21451), .ZN(n19356) );
  NAND3_X1 U13415 ( .A1(n31427), .A2(n5634), .A3(n5635), .ZN(n5633) );
  NOR2_X1 U13416 ( .A1(n21968), .A2(n21969), .ZN(n21973) );
  NOR2_X1 U13418 ( .A1(n3375), .A2(n3374), .ZN(n3373) );
  INV_X1 U13419 ( .A(n30423), .ZN(n3375) );
  NOR2_X1 U13420 ( .A1(n22956), .A2(n4514), .ZN(n21871) );
  NAND2_X1 U13421 ( .A1(n12613), .A2(n3377), .ZN(n3376) );
  NOR2_X1 U13422 ( .A1(n51429), .A2(n36133), .ZN(n38158) );
  NAND4_X1 U13423 ( .A1(n12503), .A2(n8024), .A3(n12514), .A4(n12502), .ZN(
        n12509) );
  NOR2_X1 U13424 ( .A1(n47152), .A2(n46888), .ZN(n46890) );
  INV_X1 U13425 ( .A(n21556), .ZN(n20783) );
  NAND2_X2 U13426 ( .A1(n7045), .A2(n777), .ZN(n21556) );
  NAND2_X1 U13427 ( .A1(n4656), .A2(n19087), .ZN(n3378) );
  XNOR2_X1 U13428 ( .A(n3380), .B(n16171), .ZN(n16175) );
  XNOR2_X1 U13429 ( .A(n16170), .B(n16169), .ZN(n3380) );
  AND3_X1 U13431 ( .A1(n19694), .A2(n19692), .A3(n19693), .ZN(n3381) );
  NAND2_X1 U13432 ( .A1(n14256), .A2(n3382), .ZN(n17691) );
  NAND2_X1 U13434 ( .A1(n3413), .A2(n30069), .ZN(n4730) );
  NAND2_X1 U13435 ( .A1(n3386), .A2(n651), .ZN(n3385) );
  NAND2_X1 U13437 ( .A1(n17082), .A2(n19094), .ZN(n17086) );
  OR2_X2 U13439 ( .A1(n31800), .A2(n31873), .ZN(n31882) );
  NAND2_X1 U13441 ( .A1(n5251), .A2(n2116), .ZN(n12475) );
  INV_X1 U13442 ( .A(n20561), .ZN(n7222) );
  XNOR2_X1 U13443 ( .A(n13811), .B(n8176), .ZN(n8175) );
  OR2_X1 U13444 ( .A1(n19296), .A2(n19289), .ZN(n21595) );
  INV_X1 U13445 ( .A(n36519), .ZN(n34985) );
  NAND3_X1 U13446 ( .A1(n24094), .A2(n24095), .A3(n28761), .ZN(n24096) );
  NAND3_X1 U13447 ( .A1(n30394), .A2(n28757), .A3(n5300), .ZN(n28761) );
  NAND2_X1 U13448 ( .A1(n29464), .A2(n29463), .ZN(n3388) );
  NAND4_X1 U13451 ( .A1(n40518), .A2(n40517), .A3(n3390), .A4(n40519), .ZN(
        n4395) );
  AOI21_X1 U13452 ( .B1(n7839), .B2(n51756), .A(n5458), .ZN(n5457) );
  NAND2_X1 U13453 ( .A1(n3391), .A2(n30015), .ZN(n29094) );
  NAND2_X1 U13454 ( .A1(n31689), .A2(n2530), .ZN(n3391) );
  INV_X1 U13455 ( .A(Ciphertext[141]), .ZN(n3392) );
  NOR2_X1 U13456 ( .A1(n31511), .A2(n3394), .ZN(n3393) );
  INV_X1 U13457 ( .A(n10615), .ZN(n9920) );
  NAND2_X1 U13458 ( .A1(n9908), .A2(n9915), .ZN(n10615) );
  XNOR2_X1 U13459 ( .A(n35667), .B(n36873), .ZN(n35671) );
  INV_X1 U13460 ( .A(n13841), .ZN(n7465) );
  INV_X1 U13461 ( .A(n12211), .ZN(n13136) );
  NAND2_X1 U13462 ( .A1(n6793), .A2(n13853), .ZN(n6794) );
  INV_X1 U13463 ( .A(n22733), .ZN(n6277) );
  NAND3_X1 U13464 ( .A1(n6402), .A2(n31027), .A3(n6401), .ZN(n6399) );
  NAND3_X1 U13465 ( .A1(n15188), .A2(n15243), .A3(n15234), .ZN(n13272) );
  NAND3_X1 U13467 ( .A1(n9944), .A2(n11655), .A3(n5917), .ZN(n9314) );
  AND3_X2 U13468 ( .A1(n10560), .A2(n7413), .A3(n10561), .ZN(n14342) );
  NAND2_X1 U13469 ( .A1(n31669), .A2(n32688), .ZN(n28602) );
  NAND2_X1 U13470 ( .A1(n32705), .A2(n32327), .ZN(n32332) );
  NAND3_X1 U13471 ( .A1(n37782), .A2(n37780), .A3(n33462), .ZN(n39337) );
  NAND2_X1 U13472 ( .A1(n3629), .A2(n12020), .ZN(n3395) );
  NAND3_X1 U13473 ( .A1(n36565), .A2(n36558), .A3(n36496), .ZN(n6397) );
  OR3_X1 U13474 ( .A1(n27994), .A2(n27993), .A3(n28577), .ZN(n28585) );
  INV_X1 U13476 ( .A(n19371), .ZN(n20390) );
  NAND2_X1 U13477 ( .A1(n20466), .A2(n20472), .ZN(n19371) );
  NAND2_X1 U13478 ( .A1(n22023), .A2(n23445), .ZN(n22022) );
  OR2_X1 U13479 ( .A1(n19652), .A2(n19651), .ZN(n19743) );
  NAND3_X1 U13480 ( .A1(n7772), .A2(n38727), .A3(n38731), .ZN(n39301) );
  NAND2_X1 U13481 ( .A1(n29785), .A2(n30736), .ZN(n29786) );
  NOR2_X1 U13482 ( .A1(n18088), .A2(n17627), .ZN(n20511) );
  NAND2_X1 U13483 ( .A1(n22734), .A2(n3397), .ZN(n22746) );
  NAND3_X1 U13484 ( .A1(n22729), .A2(n3398), .A3(n22730), .ZN(n3397) );
  NAND2_X1 U13485 ( .A1(n14611), .A2(n3399), .ZN(n14595) );
  OR2_X1 U13488 ( .A1(n30411), .A2(n28982), .ZN(n28178) );
  AND2_X1 U13491 ( .A1(n19026), .A2(n19025), .ZN(n7188) );
  OR2_X1 U13492 ( .A1(n32151), .A2(n31724), .ZN(n32152) );
  INV_X1 U13493 ( .A(n23464), .ZN(n21953) );
  INV_X1 U13494 ( .A(n9632), .ZN(n11368) );
  INV_X1 U13495 ( .A(n19016), .ZN(n19776) );
  XNOR2_X1 U13496 ( .A(n24578), .B(n8322), .ZN(n8323) );
  INV_X1 U13497 ( .A(n30434), .ZN(n28329) );
  INV_X1 U13498 ( .A(n39305), .ZN(n5553) );
  INV_X1 U13499 ( .A(n22360), .ZN(n22913) );
  INV_X1 U13500 ( .A(n41670), .ZN(n3490) );
  INV_X1 U13501 ( .A(n9632), .ZN(n6677) );
  NAND4_X1 U13502 ( .A1(n9369), .A2(n12097), .A3(n51138), .A4(n12380), .ZN(
        n9677) );
  NAND2_X1 U13503 ( .A1(n3403), .A2(n3402), .ZN(n20499) );
  NAND2_X1 U13504 ( .A1(n20498), .A2(n774), .ZN(n3402) );
  NAND2_X1 U13505 ( .A1(n3404), .A2(n6180), .ZN(n3403) );
  NAND2_X1 U13506 ( .A1(n22309), .A2(n2516), .ZN(n20529) );
  NAND2_X1 U13507 ( .A1(n51300), .A2(n51313), .ZN(n49638) );
  NAND2_X1 U13508 ( .A1(n19700), .A2(n17200), .ZN(n3409) );
  NAND2_X1 U13509 ( .A1(n17198), .A2(n17199), .ZN(n3410) );
  NAND2_X1 U13510 ( .A1(n5916), .A2(n2411), .ZN(n9313) );
  NAND3_X1 U13511 ( .A1(n20379), .A2(n20378), .A3(n3412), .ZN(n3411) );
  NOR2_X1 U13512 ( .A1(n7658), .A2(n30940), .ZN(n3413) );
  XNOR2_X1 U13513 ( .A(n3414), .B(n47459), .ZN(Plaintext[67]) );
  NAND4_X1 U13514 ( .A1(n47458), .A2(n47455), .A3(n47457), .A4(n47456), .ZN(
        n3414) );
  NAND3_X1 U13515 ( .A1(n3415), .A2(n49890), .A3(n46174), .ZN(n46183) );
  NAND2_X1 U13516 ( .A1(n35727), .A2(n35726), .ZN(n3416) );
  NAND2_X1 U13517 ( .A1(n10192), .A2(n10250), .ZN(n9743) );
  NAND3_X2 U13518 ( .A1(n3417), .A2(n37715), .A3(n37714), .ZN(n42907) );
  INV_X1 U13519 ( .A(n23706), .ZN(n24336) );
  NAND2_X1 U13520 ( .A1(n3419), .A2(n3418), .ZN(n13237) );
  NOR2_X1 U13522 ( .A1(n29887), .A2(n3421), .ZN(n30365) );
  NAND3_X1 U13523 ( .A1(n22120), .A2(n22121), .A3(n22116), .ZN(n18384) );
  NAND3_X1 U13524 ( .A1(n37510), .A2(n37501), .A3(n37762), .ZN(n37497) );
  XNOR2_X1 U13525 ( .A(n3422), .B(n48999), .ZN(Plaintext[91]) );
  NAND3_X1 U13526 ( .A1(n48997), .A2(n4436), .A3(n48998), .ZN(n3422) );
  XNOR2_X1 U13528 ( .A(n3424), .B(n32272), .ZN(n32274) );
  XNOR2_X1 U13529 ( .A(n32273), .B(n36723), .ZN(n3424) );
  NAND3_X1 U13530 ( .A1(n38101), .A2(n40097), .A3(n40910), .ZN(n38103) );
  XNOR2_X1 U13531 ( .A(n3718), .B(n35401), .ZN(n3426) );
  NAND2_X1 U13532 ( .A1(n30911), .A2(n29686), .ZN(n29684) );
  NAND2_X1 U13533 ( .A1(n39667), .A2(n40003), .ZN(n39100) );
  NAND2_X1 U13534 ( .A1(n47093), .A2(n47104), .ZN(n46877) );
  INV_X1 U13538 ( .A(n31549), .ZN(n32667) );
  NAND3_X1 U13539 ( .A1(n12917), .A2(n13103), .A3(n12916), .ZN(n12918) );
  INV_X1 U13540 ( .A(n12211), .ZN(n3679) );
  NAND3_X1 U13541 ( .A1(n37195), .A2(n38323), .A3(n38339), .ZN(n38326) );
  NAND3_X2 U13542 ( .A1(n13724), .A2(n8145), .A3(n13726), .ZN(n17902) );
  NAND2_X1 U13543 ( .A1(n12702), .A2(n11123), .ZN(n12699) );
  NAND2_X1 U13545 ( .A1(n785), .A2(n3427), .ZN(n12948) );
  INV_X1 U13546 ( .A(Ciphertext[136]), .ZN(n7140) );
  NAND2_X1 U13547 ( .A1(n3432), .A2(n3429), .ZN(n37361) );
  NAND2_X1 U13548 ( .A1(n3431), .A2(n3430), .ZN(n3429) );
  INV_X1 U13549 ( .A(n39565), .ZN(n3430) );
  NAND3_X1 U13550 ( .A1(n39566), .A2(n39908), .A3(n38445), .ZN(n3431) );
  NAND2_X1 U13551 ( .A1(n37359), .A2(n39565), .ZN(n3432) );
  NAND2_X1 U13552 ( .A1(n30370), .A2(n3433), .ZN(n5029) );
  XNOR2_X2 U13554 ( .A(n9198), .B(Key[129]), .ZN(n12635) );
  INV_X1 U13555 ( .A(n4007), .ZN(n15260) );
  NOR2_X1 U13556 ( .A1(n39307), .A2(n38317), .ZN(n35854) );
  AOI22_X1 U13557 ( .A1(n46890), .A2(n44471), .B1(n47150), .B2(n47153), .ZN(
        n44472) );
  NOR2_X1 U13558 ( .A1(n30043), .A2(n31339), .ZN(n30052) );
  INV_X1 U13559 ( .A(n29226), .ZN(n25420) );
  NAND2_X1 U13562 ( .A1(n4192), .A2(n5712), .ZN(n3435) );
  INV_X1 U13563 ( .A(n12018), .ZN(n13167) );
  NAND3_X1 U13565 ( .A1(n47743), .A2(n47771), .A3(n47789), .ZN(n47779) );
  OAI211_X1 U13566 ( .C1(n49514), .C2(n49511), .A(n49510), .B(n3437), .ZN(
        n49517) );
  INV_X1 U13567 ( .A(n49530), .ZN(n3437) );
  AND2_X1 U13569 ( .A1(n46244), .A2(n46252), .ZN(n49178) );
  NAND2_X1 U13570 ( .A1(n13608), .A2(n13609), .ZN(n13616) );
  NAND2_X1 U13571 ( .A1(n30850), .A2(n30582), .ZN(n30585) );
  AND2_X1 U13576 ( .A1(n14991), .A2(n14992), .ZN(n15137) );
  NAND3_X1 U13577 ( .A1(n8387), .A2(n8386), .A3(n15140), .ZN(n3439) );
  OR2_X1 U13578 ( .A1(n17619), .A2(n8558), .ZN(n8559) );
  NAND2_X1 U13579 ( .A1(n40967), .A2(n40972), .ZN(n40921) );
  AND2_X1 U13580 ( .A1(n37518), .A2(n33558), .ZN(n33559) );
  XNOR2_X1 U13581 ( .A(n33263), .B(n37134), .ZN(n31351) );
  NAND2_X1 U13582 ( .A1(n28614), .A2(n398), .ZN(n29515) );
  INV_X1 U13583 ( .A(n30673), .ZN(n26855) );
  AND2_X1 U13584 ( .A1(n38988), .A2(n38987), .ZN(n7207) );
  AND2_X1 U13585 ( .A1(n50199), .A2(n50227), .ZN(n4570) );
  INV_X1 U13586 ( .A(n51751), .ZN(n7999) );
  INV_X1 U13587 ( .A(n28882), .ZN(n28530) );
  INV_X1 U13588 ( .A(n33005), .ZN(n31380) );
  INV_X1 U13589 ( .A(n41692), .ZN(n41621) );
  INV_X1 U13590 ( .A(n18060), .ZN(n18326) );
  AOI22_X1 U13592 ( .A1(n7571), .A2(n14923), .B1(n15300), .B2(n14924), .ZN(
        n3731) );
  OAI21_X1 U13593 ( .B1(n9021), .B2(n9020), .A(n9783), .ZN(n6443) );
  NOR2_X1 U13594 ( .A1(n6157), .A2(n32609), .ZN(n32618) );
  INV_X1 U13595 ( .A(n13822), .ZN(n8226) );
  NOR2_X1 U13597 ( .A1(n22901), .A2(n5737), .ZN(n5736) );
  INV_X1 U13598 ( .A(n13819), .ZN(n7304) );
  XNOR2_X1 U13599 ( .A(n13976), .B(n17113), .ZN(n14381) );
  XNOR2_X1 U13600 ( .A(n26393), .B(n26395), .ZN(n4801) );
  XOR2_X1 U13601 ( .A(n42263), .B(n42473), .Z(n8138) );
  OAI211_X1 U13602 ( .C1(n6153), .C2(n10420), .A(n5366), .B(n2506), .ZN(n6152)
         );
  NAND2_X1 U13603 ( .A1(n36629), .A2(n38092), .ZN(n36635) );
  NAND3_X1 U13604 ( .A1(n45522), .A2(n45534), .A3(n45521), .ZN(n4428) );
  NOR2_X1 U13605 ( .A1(n2345), .A2(n3440), .ZN(n39137) );
  XNOR2_X1 U13606 ( .A(n3441), .B(n48108), .ZN(Plaintext[42]) );
  NAND4_X1 U13607 ( .A1(n8308), .A2(n48107), .A3(n48106), .A4(n48105), .ZN(
        n3441) );
  OR2_X1 U13610 ( .A1(n3506), .A2(n452), .ZN(n21053) );
  INV_X1 U13612 ( .A(n7823), .ZN(n9699) );
  NAND2_X1 U13613 ( .A1(n3443), .A2(n10234), .ZN(n9702) );
  NAND2_X1 U13614 ( .A1(n7823), .A2(n12280), .ZN(n3443) );
  INV_X1 U13615 ( .A(n12278), .ZN(n3444) );
  INV_X1 U13616 ( .A(n5335), .ZN(n3445) );
  NAND3_X1 U13617 ( .A1(n13856), .A2(n13841), .A3(n14883), .ZN(n9724) );
  NAND2_X1 U13619 ( .A1(n32302), .A2(n7041), .ZN(n3446) );
  INV_X1 U13620 ( .A(n3507), .ZN(n18222) );
  AOI21_X1 U13621 ( .B1(n7164), .B2(n9781), .A(n9782), .ZN(n7163) );
  NAND2_X2 U13623 ( .A1(n3448), .A2(n18368), .ZN(n23207) );
  NAND2_X1 U13624 ( .A1(n3599), .A2(n2368), .ZN(n3598) );
  OR2_X1 U13625 ( .A1(n46637), .A2(n52154), .ZN(n3449) );
  NAND2_X1 U13626 ( .A1(n46642), .A2(n45761), .ZN(n44421) );
  XNOR2_X1 U13628 ( .A(n15868), .B(n16896), .ZN(n15869) );
  NOR2_X1 U13629 ( .A1(n11022), .A2(n2508), .ZN(n11024) );
  INV_X1 U13630 ( .A(n32911), .ZN(n32907) );
  NAND3_X1 U13632 ( .A1(n45800), .A2(n46756), .A3(n46738), .ZN(n41813) );
  NAND3_X1 U13633 ( .A1(n2858), .A2(n47195), .A3(n49432), .ZN(n49452) );
  OR2_X2 U13634 ( .A1(n3452), .A2(n39522), .ZN(n43609) );
  OAI211_X1 U13635 ( .C1(n222), .C2(n39296), .A(n39294), .B(n39295), .ZN(
        n39306) );
  NAND2_X1 U13636 ( .A1(n37182), .A2(n39293), .ZN(n39295) );
  XNOR2_X2 U13638 ( .A(n16061), .B(n16381), .ZN(n21530) );
  NAND2_X1 U13639 ( .A1(n30367), .A2(n3454), .ZN(n3453) );
  INV_X1 U13640 ( .A(n30734), .ZN(n3454) );
  NAND2_X1 U13641 ( .A1(n30734), .A2(n30368), .ZN(n3455) );
  NAND2_X1 U13642 ( .A1(n6637), .A2(n38475), .ZN(n37416) );
  NAND3_X1 U13643 ( .A1(n3456), .A2(n44582), .A3(n2445), .ZN(n44584) );
  NAND2_X1 U13644 ( .A1(n50276), .A2(n50280), .ZN(n3456) );
  NAND2_X1 U13645 ( .A1(n16857), .A2(n18905), .ZN(n3457) );
  INV_X1 U13647 ( .A(n10471), .ZN(n10472) );
  NAND3_X1 U13648 ( .A1(n48613), .A2(n6803), .A3(n6804), .ZN(n6802) );
  NOR2_X1 U13649 ( .A1(n48593), .A2(n48640), .ZN(n48613) );
  NAND2_X1 U13651 ( .A1(n47154), .A2(n2178), .ZN(n4290) );
  INV_X1 U13652 ( .A(n35369), .ZN(n8504) );
  NAND2_X1 U13653 ( .A1(n14362), .A2(n14550), .ZN(n3460) );
  NAND2_X1 U13654 ( .A1(n43898), .A2(n43899), .ZN(n43903) );
  NAND2_X1 U13655 ( .A1(n51382), .A2(n48633), .ZN(n48639) );
  INV_X1 U13656 ( .A(n14640), .ZN(n11303) );
  NAND4_X2 U13657 ( .A1(n39806), .A2(n39805), .A3(n40589), .A4(n39804), .ZN(
        n43206) );
  NAND2_X1 U13659 ( .A1(n11582), .A2(n11579), .ZN(n9127) );
  INV_X1 U13660 ( .A(n44113), .ZN(n50609) );
  INV_X1 U13661 ( .A(n7015), .ZN(n40783) );
  INV_X1 U13662 ( .A(n20828), .ZN(n20830) );
  XNOR2_X1 U13663 ( .A(n33581), .B(n33580), .ZN(n7190) );
  NAND3_X1 U13664 ( .A1(n36330), .A2(n35012), .A3(n31621), .ZN(n35014) );
  AND2_X1 U13665 ( .A1(n15560), .A2(n15559), .ZN(n22708) );
  NAND2_X1 U13666 ( .A1(n41792), .A2(n41796), .ZN(n42105) );
  NAND2_X1 U13668 ( .A1(n36562), .A2(n36558), .ZN(n36014) );
  NAND2_X1 U13669 ( .A1(n23039), .A2(n23040), .ZN(n23041) );
  NAND2_X1 U13670 ( .A1(n5671), .A2(n51374), .ZN(n17869) );
  NAND2_X1 U13671 ( .A1(n34183), .A2(n7116), .ZN(n7118) );
  AND2_X1 U13672 ( .A1(n13766), .A2(n13767), .ZN(n4350) );
  NAND3_X1 U13673 ( .A1(n21295), .A2(n766), .A3(n19796), .ZN(n7098) );
  NAND3_X1 U13674 ( .A1(n18065), .A2(n18326), .A3(n18071), .ZN(n14386) );
  INV_X1 U13675 ( .A(Ciphertext[173]), .ZN(n7708) );
  INV_X1 U13676 ( .A(n30571), .ZN(n30579) );
  INV_X1 U13677 ( .A(n19795), .ZN(n19792) );
  AND2_X1 U13678 ( .A1(n21695), .A2(n22211), .ZN(n4324) );
  AND2_X1 U13679 ( .A1(n45909), .A2(n49717), .ZN(n45910) );
  INV_X1 U13681 ( .A(n10055), .ZN(n10967) );
  INV_X1 U13682 ( .A(n48156), .ZN(n46547) );
  XNOR2_X1 U13683 ( .A(n35760), .B(n37329), .ZN(n7048) );
  INV_X1 U13684 ( .A(n23982), .ZN(n24002) );
  INV_X1 U13686 ( .A(n27680), .ZN(n27577) );
  INV_X1 U13687 ( .A(n11084), .ZN(n11083) );
  NAND2_X1 U13688 ( .A1(n7354), .A2(n12675), .ZN(n11084) );
  INV_X1 U13689 ( .A(n39417), .ZN(n39414) );
  INV_X1 U13690 ( .A(n14149), .ZN(n6835) );
  XNOR2_X1 U13691 ( .A(n6851), .B(n6852), .ZN(n5664) );
  XNOR2_X1 U13692 ( .A(n8118), .B(n18186), .ZN(n4635) );
  XNOR2_X1 U13693 ( .A(n33946), .B(n5367), .ZN(n33555) );
  OAI21_X1 U13694 ( .B1(n27660), .B2(n27670), .A(n27654), .ZN(n5477) );
  MUX2_X1 U13695 ( .A(n17502), .B(n17501), .S(n18318), .Z(n17509) );
  NOR2_X1 U13696 ( .A1(n45848), .A2(n46614), .ZN(n3999) );
  NAND3_X1 U13697 ( .A1(n4859), .A2(n4858), .A3(n12254), .ZN(n12262) );
  INV_X1 U13698 ( .A(n49771), .ZN(n6248) );
  INV_X1 U13699 ( .A(n45898), .ZN(n49708) );
  INV_X1 U13700 ( .A(n49842), .ZN(n49784) );
  OAI22_X1 U13701 ( .A1(n12268), .A2(n12267), .B1(n12266), .B2(n6928), .ZN(
        n12270) );
  OAI21_X1 U13702 ( .B1(n37594), .B2(n36222), .A(n37366), .ZN(n36223) );
  XNOR2_X2 U13703 ( .A(n18523), .B(n16722), .ZN(n19210) );
  XNOR2_X1 U13704 ( .A(n3466), .B(n18445), .ZN(n18452) );
  XNOR2_X1 U13705 ( .A(n18446), .B(n18444), .ZN(n3466) );
  NAND2_X1 U13706 ( .A1(n49393), .A2(n49465), .ZN(n6472) );
  NAND2_X1 U13707 ( .A1(n36488), .A2(n36490), .ZN(n35311) );
  XNOR2_X1 U13708 ( .A(n4292), .B(n18769), .ZN(n3467) );
  NOR2_X1 U13709 ( .A1(n32018), .A2(n32471), .ZN(n32034) );
  OAI211_X1 U13711 ( .C1(n48588), .C2(n48641), .A(n3468), .B(n48583), .ZN(
        n48578) );
  NAND2_X1 U13712 ( .A1(n23562), .A2(n51676), .ZN(n20720) );
  NAND3_X1 U13714 ( .A1(n40959), .A2(n40963), .A3(n40970), .ZN(n3469) );
  XNOR2_X1 U13717 ( .A(n3472), .B(n15719), .ZN(n17284) );
  NAND2_X1 U13718 ( .A1(n30268), .A2(n52102), .ZN(n29239) );
  NAND2_X1 U13719 ( .A1(n5787), .A2(n3473), .ZN(n47557) );
  OAI21_X1 U13720 ( .B1(n3475), .B2(n3474), .A(n21604), .ZN(n4912) );
  NAND2_X2 U13721 ( .A1(n8737), .A2(n21111), .ZN(n24891) );
  NAND2_X1 U13722 ( .A1(n19411), .A2(n3476), .ZN(n18044) );
  NAND2_X1 U13724 ( .A1(n23436), .A2(n22593), .ZN(n23440) );
  XNOR2_X1 U13727 ( .A(n3478), .B(n35629), .ZN(n35631) );
  XNOR2_X1 U13728 ( .A(n35620), .B(n35621), .ZN(n3478) );
  XNOR2_X2 U13729 ( .A(n34740), .B(n8503), .ZN(n39027) );
  NAND4_X1 U13730 ( .A1(n8559), .A2(n8560), .A3(n17617), .A4(n19349), .ZN(
        n17618) );
  NAND2_X1 U13733 ( .A1(n3483), .A2(n3482), .ZN(n20580) );
  NAND2_X1 U13734 ( .A1(n20579), .A2(n22386), .ZN(n3482) );
  NOR2_X1 U13735 ( .A1(n26754), .A2(n27697), .ZN(n3799) );
  INV_X1 U13736 ( .A(n3604), .ZN(n19712) );
  OAI211_X1 U13737 ( .C1(n3241), .C2(n31010), .A(n3485), .B(n31380), .ZN(n3484) );
  NAND2_X1 U13738 ( .A1(n3487), .A2(n31385), .ZN(n3486) );
  INV_X1 U13739 ( .A(n8260), .ZN(n3487) );
  OR2_X2 U13740 ( .A1(n26504), .A2(n26505), .ZN(n31385) );
  NAND2_X1 U13741 ( .A1(n21906), .A2(n3488), .ZN(n21915) );
  INV_X1 U13742 ( .A(n41245), .ZN(n3489) );
  OAI211_X1 U13743 ( .C1(n20330), .C2(n3492), .A(n3491), .B(n21432), .ZN(
        n20331) );
  OR2_X1 U13744 ( .A1(n20840), .A2(n20838), .ZN(n21432) );
  INV_X1 U13745 ( .A(n19957), .ZN(n21426) );
  NAND2_X1 U13747 ( .A1(n3494), .A2(n40943), .ZN(n41530) );
  NAND2_X1 U13749 ( .A1(n3495), .A2(n22088), .ZN(n3496) );
  NAND2_X1 U13752 ( .A1(n3501), .A2(n15436), .ZN(n15344) );
  NAND3_X1 U13753 ( .A1(n15446), .A2(n15342), .A3(n15341), .ZN(n3501) );
  INV_X2 U13754 ( .A(n32473), .ZN(n32487) );
  NAND2_X1 U13756 ( .A1(n3503), .A2(n27569), .ZN(n27644) );
  OAI21_X1 U13757 ( .B1(n3504), .B2(n15299), .A(n15302), .ZN(n15313) );
  NOR2_X1 U13758 ( .A1(n15301), .A2(n15300), .ZN(n3504) );
  NAND2_X1 U13759 ( .A1(n15766), .A2(n12742), .ZN(n15299) );
  OR2_X2 U13760 ( .A1(n20332), .A2(n20331), .ZN(n23045) );
  NAND2_X1 U13761 ( .A1(n23414), .A2(n3506), .ZN(n23424) );
  OAI21_X1 U13762 ( .B1(n21293), .B2(n3686), .A(n3507), .ZN(n18986) );
  AOI21_X1 U13763 ( .B1(n7654), .B2(n21305), .A(n3507), .ZN(n21306) );
  NAND2_X1 U13764 ( .A1(n21308), .A2(n3507), .ZN(n7346) );
  INV_X1 U13766 ( .A(n3509), .ZN(n21282) );
  AOI21_X1 U13767 ( .B1(n19122), .B2(n5229), .A(n3509), .ZN(n19791) );
  NAND2_X1 U13768 ( .A1(n15134), .A2(n14269), .ZN(n3510) );
  NAND3_X1 U13769 ( .A1(n12872), .A2(n12870), .A3(n12871), .ZN(n12962) );
  INV_X1 U13770 ( .A(n23447), .ZN(n22012) );
  INV_X1 U13771 ( .A(n23436), .ZN(n3513) );
  INV_X1 U13772 ( .A(n23436), .ZN(n7689) );
  XNOR2_X2 U13773 ( .A(Key[90]), .B(Ciphertext[83]), .ZN(n11467) );
  NOR2_X1 U13774 ( .A1(n6578), .A2(n3514), .ZN(n7172) );
  AOI22_X1 U13775 ( .A1(n41932), .A2(n41933), .B1(n3514), .B2(n41934), .ZN(
        n41935) );
  AOI21_X1 U13776 ( .B1(n39540), .B2(n41934), .A(n3514), .ZN(n39546) );
  NAND3_X1 U13777 ( .A1(n12007), .A2(n13412), .A3(n3515), .ZN(n12012) );
  AOI21_X1 U13778 ( .B1(n29635), .B2(n31385), .A(n3242), .ZN(n29638) );
  OAI21_X1 U13779 ( .B1(n18898), .B2(n16125), .A(n20615), .ZN(n3518) );
  NAND2_X1 U13780 ( .A1(n3517), .A2(n3516), .ZN(n8139) );
  NAND2_X1 U13781 ( .A1(n21531), .A2(n20608), .ZN(n3516) );
  NAND2_X1 U13782 ( .A1(n16127), .A2(n3518), .ZN(n3517) );
  INV_X1 U13783 ( .A(Ciphertext[130]), .ZN(n8696) );
  AND2_X1 U13784 ( .A1(n13426), .A2(n13407), .ZN(n3519) );
  XNOR2_X2 U13785 ( .A(n18668), .B(n18756), .ZN(n16722) );
  OAI22_X1 U13786 ( .A1(n23276), .A2(n23833), .B1(n24157), .B2(n630), .ZN(
        n23278) );
  OR2_X2 U13787 ( .A1(n3521), .A2(n3522), .ZN(n48077) );
  AOI21_X1 U13788 ( .B1(n52178), .B2(n44430), .A(n3523), .ZN(n3522) );
  NAND2_X1 U13789 ( .A1(n44431), .A2(n48434), .ZN(n3523) );
  XNOR2_X1 U13790 ( .A(n51427), .B(n45401), .ZN(n36723) );
  XNOR2_X1 U13791 ( .A(n51427), .B(n37107), .ZN(n37109) );
  XNOR2_X1 U13792 ( .A(n51427), .B(n32859), .ZN(n33085) );
  XNOR2_X1 U13793 ( .A(n51427), .B(n35820), .ZN(n35821) );
  NAND3_X1 U13794 ( .A1(n3525), .A2(n30537), .A3(n33002), .ZN(n30538) );
  XNOR2_X1 U13795 ( .A(n3526), .B(n8515), .ZN(n43132) );
  XNOR2_X1 U13796 ( .A(n3526), .B(n44314), .ZN(n42928) );
  NAND2_X1 U13797 ( .A1(n37762), .A2(n37757), .ZN(n3527) );
  OAI21_X1 U13798 ( .B1(n3529), .B2(n37749), .A(n3528), .ZN(n5608) );
  NAND3_X1 U13799 ( .A1(n40458), .A2(n3531), .A3(n3530), .ZN(n37350) );
  XNOR2_X1 U13800 ( .A(n40397), .B(n40446), .ZN(n3531) );
  NAND2_X1 U13801 ( .A1(n26855), .A2(n3533), .ZN(n3532) );
  NOR2_X1 U13802 ( .A1(n24687), .A2(n30664), .ZN(n3533) );
  NAND4_X4 U13803 ( .A1(n3535), .A2(n5008), .A3(n3536), .A4(n3534), .ZN(n32251) );
  NAND2_X1 U13804 ( .A1(n2466), .A2(n26855), .ZN(n3534) );
  NAND2_X1 U13805 ( .A1(n22188), .A2(n22186), .ZN(n20561) );
  NAND2_X1 U13806 ( .A1(n3537), .A2(n19681), .ZN(n8079) );
  INV_X1 U13807 ( .A(n49705), .ZN(n49704) );
  NAND2_X1 U13808 ( .A1(n49948), .A2(n50288), .ZN(n3539) );
  NAND2_X1 U13809 ( .A1(n49615), .A2(n49614), .ZN(n3540) );
  NAND4_X1 U13810 ( .A1(n3544), .A2(n3543), .A3(n3542), .A4(n3541), .ZN(n49818) );
  NAND3_X1 U13811 ( .A1(n49816), .A2(n49815), .A3(n2440), .ZN(n3541) );
  NAND2_X1 U13812 ( .A1(n49804), .A2(n49829), .ZN(n3542) );
  INV_X1 U13814 ( .A(n49816), .ZN(n3545) );
  INV_X1 U13816 ( .A(n49803), .ZN(n3547) );
  NOR2_X1 U13817 ( .A1(n3549), .A2(n49841), .ZN(n3548) );
  NAND2_X1 U13818 ( .A1(n3944), .A2(n49841), .ZN(n49816) );
  NAND4_X2 U13819 ( .A1(n29947), .A2(n4444), .A3(n29946), .A4(n29945), .ZN(
        n32356) );
  NAND2_X1 U13820 ( .A1(n3552), .A2(n483), .ZN(n12793) );
  NAND2_X1 U13821 ( .A1(n12791), .A2(n3551), .ZN(n12897) );
  AND2_X1 U13822 ( .A1(n3552), .A2(n13429), .ZN(n3551) );
  OAI21_X1 U13823 ( .B1(n14652), .B2(n3552), .A(n13434), .ZN(n13435) );
  NAND3_X1 U13824 ( .A1(n51695), .A2(n3553), .A3(n20942), .ZN(n21774) );
  OAI211_X1 U13825 ( .C1(n36031), .C2(n37962), .A(n36030), .B(n37966), .ZN(
        n3554) );
  NAND2_X1 U13826 ( .A1(n5218), .A2(n37965), .ZN(n37966) );
  INV_X1 U13827 ( .A(n36539), .ZN(n5218) );
  NAND2_X1 U13829 ( .A1(n3559), .A2(n3557), .ZN(n41399) );
  NAND2_X1 U13830 ( .A1(n41393), .A2(n3558), .ZN(n3557) );
  NAND2_X1 U13831 ( .A1(n41535), .A2(n41540), .ZN(n3558) );
  INV_X1 U13832 ( .A(n23609), .ZN(n7774) );
  NAND2_X1 U13833 ( .A1(n9259), .A2(n12611), .ZN(n9537) );
  NAND2_X1 U13834 ( .A1(n9540), .A2(n9541), .ZN(n3560) );
  INV_X1 U13835 ( .A(n14660), .ZN(n12786) );
  NAND4_X2 U13836 ( .A1(n3561), .A2(n12802), .A3(n12800), .A4(n12801), .ZN(
        n16023) );
  NOR2_X1 U13837 ( .A1(n2358), .A2(n3562), .ZN(n3561) );
  NAND2_X1 U13839 ( .A1(n3567), .A2(n3566), .ZN(n3569) );
  NAND3_X1 U13840 ( .A1(n3567), .A2(n3566), .A3(n49867), .ZN(n49874) );
  NAND2_X1 U13841 ( .A1(n49845), .A2(n49844), .ZN(n3566) );
  NAND2_X1 U13842 ( .A1(n49846), .A2(n49793), .ZN(n3567) );
  NAND4_X1 U13844 ( .A1(n49859), .A2(n49857), .A3(n49858), .A4(n3569), .ZN(
        n49876) );
  NAND3_X1 U13845 ( .A1(n44668), .A2(n3571), .A3(n3570), .ZN(n44671) );
  NAND2_X1 U13847 ( .A1(n48430), .A2(n48438), .ZN(n45595) );
  OR2_X1 U13849 ( .A1(n51313), .A2(n49956), .ZN(n3572) );
  INV_X1 U13850 ( .A(n49956), .ZN(n50289) );
  OAI22_X1 U13852 ( .A1(n10715), .A2(n12290), .B1(n3576), .B2(n7823), .ZN(
        n10717) );
  INV_X1 U13853 ( .A(n3576), .ZN(n10725) );
  NAND2_X1 U13854 ( .A1(n9698), .A2(n12282), .ZN(n3576) );
  NAND2_X1 U13855 ( .A1(n37892), .A2(n37884), .ZN(n38997) );
  XNOR2_X2 U13856 ( .A(n8650), .B(n34848), .ZN(n38998) );
  INV_X1 U13857 ( .A(n34906), .ZN(n37739) );
  NAND2_X1 U13858 ( .A1(n3579), .A2(n6218), .ZN(n3578) );
  NAND2_X1 U13859 ( .A1(n5688), .A2(n34661), .ZN(n3579) );
  NAND2_X1 U13860 ( .A1(n34662), .A2(n36027), .ZN(n3580) );
  NAND2_X1 U13861 ( .A1(n8202), .A2(n8012), .ZN(n34662) );
  NAND3_X1 U13862 ( .A1(n31827), .A2(n31826), .A3(n3581), .ZN(n31832) );
  NAND3_X1 U13863 ( .A1(n30579), .A2(n31821), .A3(n3581), .ZN(n26713) );
  XNOR2_X1 U13864 ( .A(n3582), .B(n41858), .ZN(n41860) );
  XNOR2_X1 U13865 ( .A(n34330), .B(n3582), .ZN(n42353) );
  XNOR2_X1 U13866 ( .A(n44315), .B(n3582), .ZN(n44316) );
  NAND4_X1 U13869 ( .A1(n36308), .A2(n5979), .A3(n36309), .A4(n3586), .ZN(
        n36310) );
  OAI22_X1 U13870 ( .A1(n17203), .A2(n18973), .B1(n19704), .B2(n3589), .ZN(
        n17204) );
  NAND2_X1 U13871 ( .A1(n3589), .A2(n51434), .ZN(n18973) );
  NAND2_X1 U13872 ( .A1(n38521), .A2(n38532), .ZN(n3590) );
  OAI21_X1 U13873 ( .B1(n35961), .B2(n3591), .A(n51735), .ZN(n35965) );
  INV_X1 U13874 ( .A(n35960), .ZN(n3591) );
  NAND2_X1 U13875 ( .A1(n3634), .A2(n3593), .ZN(n3592) );
  INV_X1 U13876 ( .A(n45695), .ZN(n3593) );
  NAND2_X1 U13877 ( .A1(n30231), .A2(n4724), .ZN(n3594) );
  NAND2_X1 U13878 ( .A1(n51735), .A2(n3596), .ZN(n4977) );
  NAND3_X1 U13879 ( .A1(n38532), .A2(n3596), .A3(n38512), .ZN(n37433) );
  NAND2_X1 U13880 ( .A1(n38521), .A2(n3595), .ZN(n38524) );
  NAND2_X1 U13881 ( .A1(n37439), .A2(n37484), .ZN(n35530) );
  NAND2_X1 U13882 ( .A1(n3597), .A2(n41328), .ZN(n39814) );
  NAND3_X1 U13883 ( .A1(n3769), .A2(n5859), .A3(n3597), .ZN(n3768) );
  NAND3_X1 U13884 ( .A1(n51364), .A2(n39628), .A3(n3597), .ZN(n39630) );
  NAND2_X1 U13885 ( .A1(n20829), .A2(n20441), .ZN(n3599) );
  INV_X1 U13886 ( .A(n20829), .ZN(n20824) );
  OAI211_X1 U13887 ( .C1(n9080), .C2(n3601), .A(n9079), .B(n9078), .ZN(n9081)
         );
  INV_X1 U13888 ( .A(n9281), .ZN(n3601) );
  NAND2_X1 U13889 ( .A1(n22968), .A2(n51858), .ZN(n22969) );
  NAND2_X1 U13890 ( .A1(n23317), .A2(n21873), .ZN(n21010) );
  NAND2_X1 U13891 ( .A1(n19794), .A2(n3604), .ZN(n7876) );
  NAND2_X1 U13892 ( .A1(n19712), .A2(n766), .ZN(n3605) );
  OAI21_X1 U13893 ( .B1(n43798), .B2(n7426), .A(n3610), .ZN(n47146) );
  NAND2_X1 U13894 ( .A1(n50359), .A2(n3606), .ZN(n46806) );
  AOI21_X1 U13895 ( .B1(n50368), .B2(n3607), .A(n50361), .ZN(n3606) );
  NAND4_X1 U13896 ( .A1(n46975), .A2(n50367), .A3(n44595), .A4(n3610), .ZN(
        n44596) );
  NAND2_X1 U13897 ( .A1(n47143), .A2(n3608), .ZN(n43799) );
  INV_X1 U13898 ( .A(n3609), .ZN(n3608) );
  OAI21_X1 U13899 ( .B1(n50367), .B2(n3607), .A(n3610), .ZN(n3609) );
  NAND2_X1 U13902 ( .A1(n31828), .A2(n3612), .ZN(n3656) );
  NAND2_X1 U13903 ( .A1(n3614), .A2(n3621), .ZN(n3613) );
  NAND2_X1 U13904 ( .A1(n11328), .A2(n3615), .ZN(n3614) );
  INV_X1 U13906 ( .A(n11327), .ZN(n3619) );
  INV_X1 U13907 ( .A(n11324), .ZN(n3621) );
  NAND2_X1 U13908 ( .A1(n3622), .A2(n5452), .ZN(n5111) );
  NAND3_X1 U13910 ( .A1(n3623), .A2(n32638), .A3(n32541), .ZN(n32551) );
  NAND2_X1 U13911 ( .A1(n3626), .A2(n36542), .ZN(n3625) );
  NAND3_X1 U13912 ( .A1(n36548), .A2(n36553), .A3(n37964), .ZN(n37960) );
  INV_X1 U13914 ( .A(n44825), .ZN(n3627) );
  NAND3_X1 U13915 ( .A1(n45524), .A2(n45534), .A3(n45523), .ZN(n45833) );
  OR2_X1 U13916 ( .A1(n3628), .A2(n10904), .ZN(n10090) );
  INV_X1 U13917 ( .A(n10904), .ZN(n3629) );
  INV_X1 U13919 ( .A(n48919), .ZN(n3631) );
  NAND2_X1 U13921 ( .A1(n45696), .A2(n3633), .ZN(n3632) );
  INV_X1 U13922 ( .A(n22404), .ZN(n3635) );
  AND2_X1 U13923 ( .A1(n17583), .A2(n17571), .ZN(n3641) );
  NAND2_X1 U13924 ( .A1(n3642), .A2(n17581), .ZN(n3639) );
  NAND4_X2 U13925 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n22144) );
  INV_X1 U13926 ( .A(n17571), .ZN(n17612) );
  AOI22_X1 U13928 ( .A1(n12216), .A2(n13139), .B1(n3645), .B2(n12900), .ZN(
        n12219) );
  OAI211_X1 U13929 ( .C1(n18385), .C2(n413), .A(n18384), .B(n3646), .ZN(n18386) );
  NAND2_X1 U13930 ( .A1(n23219), .A2(n51355), .ZN(n3646) );
  NAND2_X1 U13931 ( .A1(n5942), .A2(n3647), .ZN(n5941) );
  NAND2_X1 U13932 ( .A1(n36239), .A2(n37750), .ZN(n3647) );
  NAND2_X1 U13933 ( .A1(n3649), .A2(n12325), .ZN(n9044) );
  NAND2_X1 U13934 ( .A1(n10669), .A2(n3648), .ZN(n9048) );
  AOI21_X1 U13935 ( .B1(n12337), .B2(n10669), .A(n3649), .ZN(n10670) );
  OAI21_X1 U13936 ( .B1(n10667), .B2(n3649), .A(n51462), .ZN(n10677) );
  NAND2_X1 U13937 ( .A1(n37745), .A2(n3650), .ZN(n37746) );
  NAND2_X1 U13938 ( .A1(n37750), .A2(n3650), .ZN(n37752) );
  OAI21_X1 U13939 ( .B1(n37502), .B2(n3650), .A(n37501), .ZN(n37503) );
  MUX2_X1 U13941 ( .A(n45869), .B(n47730), .S(n47771), .Z(n45009) );
  NAND2_X1 U13942 ( .A1(n44819), .A2(n44820), .ZN(n3651) );
  XNOR2_X2 U13943 ( .A(n3652), .B(n45344), .ZN(n50325) );
  NAND2_X1 U13944 ( .A1(n3654), .A2(n37977), .ZN(n36528) );
  NAND2_X1 U13946 ( .A1(n40910), .A2(n3655), .ZN(n38795) );
  NAND2_X1 U13947 ( .A1(n40903), .A2(n3655), .ZN(n40899) );
  NAND2_X1 U13948 ( .A1(n40901), .A2(n3655), .ZN(n38801) );
  NOR2_X1 U13949 ( .A1(n30581), .A2(n31816), .ZN(n3658) );
  NOR2_X1 U13950 ( .A1(n29382), .A2(n3660), .ZN(n3659) );
  NAND2_X1 U13952 ( .A1(n3663), .A2(n3661), .ZN(n32030) );
  NAND2_X1 U13953 ( .A1(n32483), .A2(n32478), .ZN(n3661) );
  NAND3_X1 U13954 ( .A1(n17611), .A2(n17610), .A3(n5018), .ZN(n3666) );
  INV_X1 U13955 ( .A(n24319), .ZN(n25440) );
  NAND3_X1 U13957 ( .A1(n17988), .A2(n17990), .A3(n17989), .ZN(n3668) );
  XNOR2_X1 U13958 ( .A(n3670), .B(n27345), .ZN(n27360) );
  XNOR2_X2 U13959 ( .A(n23744), .B(n3670), .ZN(n27609) );
  XNOR2_X1 U13960 ( .A(n24872), .B(n28398), .ZN(n3670) );
  NAND4_X1 U13961 ( .A1(n12504), .A2(n12514), .A3(n8024), .A4(n12512), .ZN(
        n3948) );
  NAND3_X1 U13962 ( .A1(n13354), .A2(n14542), .A3(n13346), .ZN(n14369) );
  NAND2_X1 U13963 ( .A1(n14370), .A2(n14552), .ZN(n13346) );
  AND2_X1 U13964 ( .A1(n14550), .A2(n14552), .ZN(n3673) );
  XNOR2_X1 U13966 ( .A(n636), .B(n576), .ZN(n15410) );
  XNOR2_X1 U13967 ( .A(n636), .B(n15707), .ZN(n16190) );
  XNOR2_X1 U13968 ( .A(n35065), .B(n3675), .ZN(n35066) );
  XNOR2_X1 U13969 ( .A(n33618), .B(n3675), .ZN(n33517) );
  XNOR2_X1 U13970 ( .A(n33371), .B(n3675), .ZN(n33381) );
  XNOR2_X1 U13971 ( .A(n3675), .B(n33364), .ZN(n33367) );
  XNOR2_X1 U13972 ( .A(n34275), .B(n3675), .ZN(n6205) );
  XNOR2_X1 U13973 ( .A(n3675), .B(n34596), .ZN(n34597) );
  INV_X1 U13974 ( .A(n14187), .ZN(n14193) );
  OR2_X1 U13975 ( .A1(n13152), .A2(n12211), .ZN(n14187) );
  NOR2_X1 U13976 ( .A1(n13152), .A2(n3677), .ZN(n3676) );
  NAND2_X1 U13977 ( .A1(n13136), .A2(n14186), .ZN(n3677) );
  INV_X1 U13978 ( .A(n12211), .ZN(n3678) );
  NAND2_X1 U13979 ( .A1(n3684), .A2(n21303), .ZN(n7655) );
  NAND2_X1 U13980 ( .A1(n18888), .A2(n3685), .ZN(n3684) );
  NAND3_X1 U13981 ( .A1(n18995), .A2(n19716), .A3(n3686), .ZN(n19002) );
  NAND2_X1 U13982 ( .A1(n31039), .A2(n31821), .ZN(n3688) );
  OAI21_X1 U13983 ( .B1(n6461), .B2(n3688), .A(n26688), .ZN(n26707) );
  NAND2_X1 U13984 ( .A1(n3689), .A2(n10372), .ZN(n9635) );
  NAND2_X1 U13985 ( .A1(n11372), .A2(n6676), .ZN(n3689) );
  INV_X2 U13986 ( .A(n22979), .ZN(n22995) );
  NAND3_X1 U13987 ( .A1(n11915), .A2(n3692), .A3(n3377), .ZN(n9544) );
  NOR2_X1 U13988 ( .A1(n11915), .A2(n9547), .ZN(n10480) );
  OAI21_X1 U13989 ( .B1(n1307), .B2(n12602), .A(n3693), .ZN(n9263) );
  NAND2_X1 U13990 ( .A1(n12603), .A2(n3693), .ZN(n12607) );
  INV_X1 U13991 ( .A(n11915), .ZN(n3693) );
  AOI22_X1 U13993 ( .A1(n14875), .A2(n3695), .B1(n13252), .B2(n14871), .ZN(
        n3694) );
  INV_X1 U13994 ( .A(n8437), .ZN(n3696) );
  NAND3_X1 U13995 ( .A1(n7245), .A2(n15421), .A3(n15425), .ZN(n3699) );
  NOR2_X1 U13996 ( .A1(n3701), .A2(n32441), .ZN(n32443) );
  NAND2_X1 U13997 ( .A1(n3702), .A2(n32438), .ZN(n3701) );
  NAND2_X1 U13998 ( .A1(n15425), .A2(n14871), .ZN(n3704) );
  AND2_X1 U13999 ( .A1(n13261), .A2(n14870), .ZN(n3705) );
  MUX2_X1 U14000 ( .A(n13887), .B(n13888), .S(n14875), .Z(n13889) );
  INV_X1 U14001 ( .A(n38664), .ZN(n38670) );
  INV_X1 U14002 ( .A(n35890), .ZN(n35407) );
  XNOR2_X1 U14003 ( .A(n3710), .B(n43702), .ZN(n14079) );
  XNOR2_X1 U14004 ( .A(n3710), .B(n2183), .ZN(n16471) );
  XNOR2_X1 U14005 ( .A(n3710), .B(n18207), .ZN(n18209) );
  NAND2_X1 U14006 ( .A1(n802), .A2(n12705), .ZN(n3712) );
  NAND2_X1 U14007 ( .A1(n3713), .A2(n17576), .ZN(n13542) );
  NAND2_X1 U14008 ( .A1(n19392), .A2(n3714), .ZN(n3713) );
  INV_X1 U14009 ( .A(n17569), .ZN(n3714) );
  INV_X1 U14010 ( .A(n19392), .ZN(n3715) );
  NAND2_X1 U14011 ( .A1(n17575), .A2(n17484), .ZN(n19392) );
  NAND2_X1 U14012 ( .A1(n2077), .A2(n29882), .ZN(n30748) );
  NAND3_X1 U14013 ( .A1(n28300), .A2(n3716), .A3(n7721), .ZN(n28299) );
  INV_X1 U14014 ( .A(n23175), .ZN(n3717) );
  NAND2_X1 U14015 ( .A1(n3717), .A2(n51021), .ZN(n22055) );
  XNOR2_X1 U14016 ( .A(n35404), .B(n3719), .ZN(n3718) );
  NAND2_X1 U14017 ( .A1(n32725), .A2(n32716), .ZN(n31645) );
  AOI21_X1 U14019 ( .B1(n29762), .B2(n3722), .A(n514), .ZN(n3724) );
  NAND3_X1 U14020 ( .A1(n29772), .A2(n29771), .A3(n29773), .ZN(n3725) );
  NAND2_X1 U14021 ( .A1(n3727), .A2(n514), .ZN(n3726) );
  NAND2_X1 U14022 ( .A1(n29756), .A2(n29757), .ZN(n3727) );
  AND3_X1 U14024 ( .A1(n37920), .A2(n37919), .A3(n3734), .ZN(n8554) );
  NAND3_X1 U14025 ( .A1(n37702), .A2(n37701), .A3(n39240), .ZN(n3734) );
  NAND2_X1 U14026 ( .A1(n37730), .A2(n3735), .ZN(n4152) );
  NAND3_X1 U14027 ( .A1(n37735), .A2(n39401), .A3(n612), .ZN(n37738) );
  NAND2_X1 U14028 ( .A1(n37732), .A2(n3736), .ZN(n37733) );
  NAND2_X1 U14030 ( .A1(n47424), .A2(n49877), .ZN(n3739) );
  OR2_X2 U14031 ( .A1(n7565), .A2(n7564), .ZN(n49932) );
  NAND2_X1 U14032 ( .A1(n25735), .A2(n25736), .ZN(n3741) );
  AND2_X1 U14033 ( .A1(n28857), .A2(n3742), .ZN(n3743) );
  NAND2_X1 U14034 ( .A1(n28851), .A2(n29070), .ZN(n3742) );
  NAND2_X1 U14035 ( .A1(n30343), .A2(n28850), .ZN(n3744) );
  NAND2_X1 U14037 ( .A1(n20478), .A2(n20474), .ZN(n3746) );
  AOI21_X1 U14038 ( .B1(n17998), .B2(n20460), .A(n3747), .ZN(n18005) );
  XNOR2_X2 U14039 ( .A(n15617), .B(n14737), .ZN(n17639) );
  NAND3_X1 U14040 ( .A1(n22189), .A2(n7119), .A3(n21700), .ZN(n3748) );
  OAI21_X1 U14041 ( .B1(n35417), .B2(n36436), .A(n3749), .ZN(n36445) );
  NAND2_X1 U14042 ( .A1(n36436), .A2(n38277), .ZN(n3749) );
  NAND2_X1 U14043 ( .A1(n38425), .A2(n3750), .ZN(n38427) );
  NAND2_X1 U14044 ( .A1(n39667), .A2(n3751), .ZN(n3750) );
  NAND2_X1 U14045 ( .A1(n15372), .A2(n3752), .ZN(n14487) );
  INV_X1 U14046 ( .A(n32760), .ZN(n3754) );
  NAND2_X1 U14047 ( .A1(n28331), .A2(n28330), .ZN(n3753) );
  NAND2_X1 U14049 ( .A1(n49722), .A2(n49711), .ZN(n49718) );
  NAND4_X1 U14050 ( .A1(n23537), .A2(n3759), .A3(n20706), .A4(n23694), .ZN(
        n3758) );
  NAND2_X1 U14051 ( .A1(n24336), .A2(n457), .ZN(n23694) );
  OAI21_X1 U14052 ( .B1(n3761), .B2(n5649), .A(n23703), .ZN(n3760) );
  INV_X1 U14053 ( .A(n23379), .ZN(n3762) );
  NAND2_X1 U14054 ( .A1(n12670), .A2(n3763), .ZN(n12688) );
  NAND2_X1 U14055 ( .A1(n11491), .A2(n3763), .ZN(n11507) );
  NAND2_X1 U14056 ( .A1(n26950), .A2(n3764), .ZN(n26869) );
  NAND2_X1 U14057 ( .A1(n3767), .A2(n31488), .ZN(n31271) );
  NAND2_X1 U14058 ( .A1(n40728), .A2(n40729), .ZN(n3771) );
  NAND2_X1 U14060 ( .A1(n40732), .A2(n5859), .ZN(n40366) );
  XNOR2_X1 U14061 ( .A(n5221), .B(n3772), .ZN(n16172) );
  XNOR2_X1 U14062 ( .A(n3772), .B(n17321), .ZN(n14859) );
  XNOR2_X1 U14063 ( .A(n3772), .B(n16610), .ZN(n16611) );
  XNOR2_X1 U14064 ( .A(n511), .B(n3772), .ZN(n15805) );
  INV_X1 U14065 ( .A(n21473), .ZN(n3774) );
  INV_X1 U14066 ( .A(n21473), .ZN(n21450) );
  OAI21_X1 U14067 ( .B1(n20487), .B2(n21458), .A(n21452), .ZN(n20489) );
  NAND2_X1 U14068 ( .A1(n3774), .A2(n20314), .ZN(n21458) );
  INV_X1 U14069 ( .A(n20447), .ZN(n20453) );
  NAND2_X1 U14070 ( .A1(n21492), .A2(n21480), .ZN(n20447) );
  NAND3_X1 U14072 ( .A1(n38159), .A2(n38160), .A3(n38585), .ZN(n38161) );
  NAND2_X1 U14074 ( .A1(n41374), .A2(n40960), .ZN(n41378) );
  NAND2_X1 U14075 ( .A1(n40957), .A2(n41375), .ZN(n41386) );
  NAND4_X2 U14076 ( .A1(n38171), .A2(n7954), .A3(n38169), .A4(n38170), .ZN(
        n40960) );
  NAND2_X1 U14078 ( .A1(n23702), .A2(n50990), .ZN(n3780) );
  NOR2_X1 U14079 ( .A1(n24336), .A2(n23531), .ZN(n3778) );
  NAND2_X1 U14080 ( .A1(n3780), .A2(n24332), .ZN(n24335) );
  AOI21_X1 U14081 ( .B1(n3781), .B2(n48905), .A(n48908), .ZN(n5080) );
  NAND3_X1 U14082 ( .A1(n3782), .A2(n48912), .A3(n48853), .ZN(n3781) );
  INV_X1 U14083 ( .A(n48853), .ZN(n5078) );
  XNOR2_X2 U14084 ( .A(n9451), .B(Key[19]), .ZN(n10037) );
  NAND2_X1 U14085 ( .A1(n3787), .A2(n3784), .ZN(n8483) );
  OAI21_X1 U14086 ( .B1(n31497), .B2(n31496), .A(n3786), .ZN(n3785) );
  NAND2_X1 U14087 ( .A1(n30998), .A2(n31496), .ZN(n3786) );
  NAND2_X1 U14088 ( .A1(n3788), .A2(n26881), .ZN(n3787) );
  XNOR2_X1 U14089 ( .A(n3791), .B(n3793), .ZN(Plaintext[93]) );
  NAND4_X1 U14090 ( .A1(n339), .A2(n3792), .A3(n3794), .A4(n3795), .ZN(n3791)
         );
  NAND2_X1 U14091 ( .A1(n49027), .A2(n49026), .ZN(n3795) );
  NAND2_X1 U14092 ( .A1(n41380), .A2(n40960), .ZN(n40239) );
  NAND2_X1 U14093 ( .A1(n41380), .A2(n3796), .ZN(n40968) );
  NAND2_X1 U14095 ( .A1(n41379), .A2(n40968), .ZN(n42086) );
  OAI21_X1 U14096 ( .B1(n47825), .B2(n51470), .A(n47880), .ZN(n3797) );
  INV_X1 U14097 ( .A(n372), .ZN(n3798) );
  NOR2_X1 U14098 ( .A1(n29330), .A2(n29327), .ZN(n27818) );
  INV_X1 U14099 ( .A(n27822), .ZN(n27819) );
  NAND2_X1 U14100 ( .A1(n27890), .A2(n27818), .ZN(n27822) );
  NAND2_X1 U14101 ( .A1(n35103), .A2(n38464), .ZN(n38467) );
  OAI211_X1 U14102 ( .C1(n35103), .C2(n38477), .A(n38468), .B(n38471), .ZN(
        n35141) );
  NAND2_X1 U14103 ( .A1(n3799), .A2(n26755), .ZN(n26759) );
  NAND2_X1 U14104 ( .A1(n3800), .A2(n27679), .ZN(n7785) );
  NAND2_X1 U14105 ( .A1(n26961), .A2(n2512), .ZN(n3800) );
  NAND3_X1 U14106 ( .A1(n13084), .A2(n13083), .A3(n3802), .ZN(n3801) );
  NAND3_X2 U14107 ( .A1(n3803), .A2(n10666), .A3(n3808), .ZN(n14601) );
  NAND3_X1 U14108 ( .A1(n11388), .A2(n10664), .A3(n10665), .ZN(n3804) );
  INV_X1 U14109 ( .A(n12051), .ZN(n11389) );
  NAND3_X1 U14110 ( .A1(n10660), .A2(n8712), .A3(n11387), .ZN(n3806) );
  NAND2_X1 U14111 ( .A1(n3809), .A2(n799), .ZN(n3808) );
  NAND2_X1 U14112 ( .A1(n11395), .A2(n10663), .ZN(n3809) );
  AOI21_X1 U14113 ( .B1(n3811), .B2(n2418), .A(n3810), .ZN(n3812) );
  NAND2_X1 U14114 ( .A1(n3813), .A2(n39406), .ZN(n37897) );
  NOR2_X1 U14115 ( .A1(n39002), .A2(n39395), .ZN(n39406) );
  NAND2_X1 U14116 ( .A1(n37740), .A2(n39400), .ZN(n39002) );
  NAND2_X1 U14117 ( .A1(n34908), .A2(n51474), .ZN(n37740) );
  NAND3_X1 U14118 ( .A1(n20606), .A2(n21560), .A3(n3814), .ZN(n7221) );
  OAI21_X1 U14119 ( .B1(n20783), .B2(n5167), .A(n21581), .ZN(n3814) );
  NAND3_X1 U14120 ( .A1(n23379), .A2(n3815), .A3(n23536), .ZN(n4442) );
  NAND2_X1 U14121 ( .A1(n3816), .A2(n50990), .ZN(n23378) );
  OR2_X1 U14122 ( .A1(n3818), .A2(n38545), .ZN(n38210) );
  INV_X1 U14123 ( .A(n38212), .ZN(n3818) );
  INV_X1 U14124 ( .A(n30669), .ZN(n26912) );
  NAND2_X1 U14125 ( .A1(n3819), .A2(n30665), .ZN(n30669) );
  AOI22_X1 U14126 ( .A1(n26913), .A2(n26912), .B1(n26910), .B2(n26911), .ZN(
        n26924) );
  AND2_X1 U14129 ( .A1(n10181), .A2(n10176), .ZN(n3824) );
  INV_X1 U14130 ( .A(n28948), .ZN(n3826) );
  OAI21_X1 U14131 ( .B1(n29797), .B2(n3827), .A(n29800), .ZN(n29798) );
  NAND2_X1 U14132 ( .A1(n3829), .A2(n3828), .ZN(n20629) );
  NAND2_X1 U14133 ( .A1(n20628), .A2(n20627), .ZN(n3828) );
  NAND2_X1 U14134 ( .A1(n20736), .A2(n20642), .ZN(n3829) );
  XNOR2_X1 U14135 ( .A(n3830), .B(n28217), .ZN(n28219) );
  XNOR2_X1 U14136 ( .A(n23937), .B(n3830), .ZN(n23781) );
  XNOR2_X1 U14137 ( .A(n25005), .B(n23745), .ZN(n3830) );
  OAI211_X1 U14139 ( .C1(n3831), .C2(n41581), .A(n42018), .B(n42006), .ZN(
        n41590) );
  NAND2_X1 U14140 ( .A1(n43284), .A2(n43283), .ZN(n3833) );
  OAI21_X1 U14141 ( .B1(n50028), .B2(n50027), .A(n3833), .ZN(n50030) );
  NAND3_X1 U14142 ( .A1(n49665), .A2(n49664), .A3(n3833), .ZN(n49679) );
  NAND3_X2 U14143 ( .A1(n43286), .A2(n43287), .A3(n3832), .ZN(n49608) );
  NOR3_X1 U14144 ( .A1(n38174), .A2(n38014), .A3(n38190), .ZN(n38191) );
  NAND2_X1 U14145 ( .A1(n6335), .A2(n3490), .ZN(n41228) );
  NAND2_X1 U14146 ( .A1(n13091), .A2(n13088), .ZN(n3834) );
  NOR2_X1 U14147 ( .A1(n13090), .A2(n3834), .ZN(n4182) );
  OAI22_X1 U14148 ( .A1(n8225), .A2(n12823), .B1(n12912), .B2(n3834), .ZN(
        n9529) );
  OAI22_X1 U14149 ( .A1(n13079), .A2(n13078), .B1(n13080), .B2(n3834), .ZN(
        n13085) );
  NAND3_X1 U14150 ( .A1(n3839), .A2(n3838), .A3(n3837), .ZN(n3836) );
  NAND3_X1 U14152 ( .A1(n34936), .A2(n34934), .A3(n3841), .ZN(n3840) );
  NAND2_X1 U14153 ( .A1(n34926), .A2(n36057), .ZN(n3841) );
  NAND3_X1 U14155 ( .A1(n49207), .A2(n49197), .A3(n49198), .ZN(n3845) );
  AND2_X2 U14156 ( .A1(n49201), .A2(n49197), .ZN(n46229) );
  NAND2_X1 U14157 ( .A1(n3842), .A2(n49201), .ZN(n3844) );
  NAND2_X1 U14158 ( .A1(n3843), .A2(n49216), .ZN(n4677) );
  NAND2_X1 U14159 ( .A1(n3845), .A2(n3844), .ZN(n3843) );
  NOR2_X1 U14160 ( .A1(n10539), .A2(n3850), .ZN(n3849) );
  INV_X1 U14161 ( .A(n51761), .ZN(n3850) );
  OAI21_X1 U14162 ( .B1(n45564), .B2(n45565), .A(n3851), .ZN(n45572) );
  NAND3_X1 U14163 ( .A1(n45563), .A2(n8684), .A3(n8685), .ZN(n3851) );
  NAND4_X1 U14164 ( .A1(n45563), .A2(n8684), .A3(n8685), .A4(n3853), .ZN(n3852) );
  INV_X1 U14165 ( .A(n48518), .ZN(n3853) );
  NAND2_X2 U14166 ( .A1(n2268), .A2(n48199), .ZN(n48381) );
  NAND2_X1 U14167 ( .A1(n7766), .A2(n8061), .ZN(n3854) );
  NAND2_X1 U14168 ( .A1(n48129), .A2(n8061), .ZN(n3855) );
  OAI21_X1 U14169 ( .B1(n48147), .B2(n3856), .A(n48146), .ZN(n48148) );
  AND3_X2 U14170 ( .A1(n3862), .A2(n3859), .A3(n3857), .ZN(n44923) );
  NAND2_X1 U14171 ( .A1(n50145), .A2(n51727), .ZN(n50064) );
  NAND2_X1 U14172 ( .A1(n3864), .A2(n51442), .ZN(n50079) );
  NAND2_X1 U14173 ( .A1(n50088), .A2(n3864), .ZN(n50069) );
  NOR2_X1 U14174 ( .A1(n3866), .A2(n17479), .ZN(n16843) );
  NAND2_X1 U14175 ( .A1(n3865), .A2(n19396), .ZN(n18022) );
  AOI21_X1 U14176 ( .B1(n18015), .B2(n18009), .A(n3866), .ZN(n17566) );
  OAI21_X1 U14177 ( .B1(n17567), .B2(n3866), .A(n18015), .ZN(n18008) );
  INV_X1 U14178 ( .A(n19396), .ZN(n3866) );
  NAND2_X1 U14180 ( .A1(n28563), .A2(n28548), .ZN(n3868) );
  INV_X1 U14181 ( .A(n51062), .ZN(n3874) );
  INV_X1 U14183 ( .A(n30692), .ZN(n28758) );
  INV_X1 U14184 ( .A(n23177), .ZN(n3876) );
  NAND2_X1 U14185 ( .A1(n3880), .A2(n3881), .ZN(n22411) );
  NAND3_X1 U14186 ( .A1(n21726), .A2(n51355), .A3(n8732), .ZN(n3880) );
  NAND3_X1 U14187 ( .A1(n21726), .A2(n22120), .A3(n3877), .ZN(n3881) );
  NAND2_X1 U14188 ( .A1(n22405), .A2(n21728), .ZN(n3878) );
  NAND2_X1 U14189 ( .A1(n21727), .A2(n22406), .ZN(n3879) );
  INV_X1 U14190 ( .A(n20501), .ZN(n8687) );
  NAND2_X1 U14192 ( .A1(n3883), .A2(n9942), .ZN(n9948) );
  AND2_X1 U14193 ( .A1(n7784), .A2(n26744), .ZN(n3884) );
  XNOR2_X2 U14194 ( .A(n16249), .B(n16544), .ZN(n3885) );
  NAND2_X1 U14195 ( .A1(n51222), .A2(n3885), .ZN(n19474) );
  NAND2_X1 U14196 ( .A1(n21252), .A2(n3885), .ZN(n19087) );
  NAND3_X1 U14197 ( .A1(n21249), .A2(n19482), .A3(n3885), .ZN(n19483) );
  INV_X1 U14198 ( .A(n3886), .ZN(n31282) );
  NOR2_X1 U14199 ( .A1(n29213), .A2(n3886), .ZN(n29218) );
  NAND2_X1 U14200 ( .A1(n45194), .A2(n50950), .ZN(n47236) );
  NAND4_X1 U14202 ( .A1(n3888), .A2(n46857), .A3(n45140), .A4(n3889), .ZN(
        n3887) );
  NAND2_X1 U14203 ( .A1(n3895), .A2(n45139), .ZN(n3888) );
  NAND2_X1 U14204 ( .A1(n46838), .A2(n4527), .ZN(n3895) );
  NAND2_X1 U14205 ( .A1(n46654), .A2(n46842), .ZN(n3893) );
  NOR2_X1 U14206 ( .A1(n46852), .A2(n46845), .ZN(n45775) );
  INV_X1 U14207 ( .A(n46844), .ZN(n3892) );
  NAND2_X1 U14208 ( .A1(n45137), .A2(n46840), .ZN(n3894) );
  NAND2_X1 U14209 ( .A1(n39462), .A2(n39035), .ZN(n39033) );
  NOR2_X1 U14210 ( .A1(n3897), .A2(n45026), .ZN(n3896) );
  NOR2_X1 U14211 ( .A1(n3901), .A2(n3900), .ZN(n3899) );
  NOR2_X1 U14213 ( .A1(n5167), .A2(n51711), .ZN(n3903) );
  AND2_X1 U14215 ( .A1(n21405), .A2(n21404), .ZN(n21410) );
  NAND2_X1 U14216 ( .A1(n21406), .A2(n3903), .ZN(n21404) );
  NOR2_X1 U14217 ( .A1(n777), .A2(n21584), .ZN(n21406) );
  OAI21_X1 U14218 ( .B1(n3906), .B2(n3904), .A(n23923), .ZN(n23927) );
  NAND2_X1 U14220 ( .A1(n23913), .A2(n23142), .ZN(n22799) );
  NOR2_X1 U14221 ( .A1(n48116), .A2(n48156), .ZN(n48152) );
  XNOR2_X1 U14222 ( .A(n3910), .B(n48164), .ZN(Plaintext[46]) );
  INV_X1 U14223 ( .A(n48117), .ZN(n3911) );
  AND2_X1 U14224 ( .A1(n24000), .A2(n3912), .ZN(n24003) );
  NAND2_X1 U14225 ( .A1(n23984), .A2(n23992), .ZN(n4485) );
  NOR2_X1 U14226 ( .A1(n23996), .A2(n3912), .ZN(n19447) );
  AOI22_X1 U14227 ( .A1(n1230), .A2(n23033), .B1(n5118), .B2(n3912), .ZN(n5117) );
  NAND3_X1 U14228 ( .A1(n23990), .A2(n23986), .A3(n3912), .ZN(n19448) );
  AND3_X2 U14229 ( .A1(n7009), .A2(n19303), .A3(n3913), .ZN(n23992) );
  NAND4_X1 U14230 ( .A1(n29312), .A2(n3917), .A3(n3916), .A4(n3915), .ZN(n3914) );
  OAI211_X1 U14231 ( .C1(n29295), .C2(n29294), .A(n29293), .B(n29292), .ZN(
        n3916) );
  OAI21_X1 U14232 ( .B1(n29304), .B2(n3918), .A(n26654), .ZN(n3917) );
  INV_X1 U14233 ( .A(n29306), .ZN(n3918) );
  INV_X1 U14234 ( .A(n32016), .ZN(n3921) );
  NAND2_X1 U14235 ( .A1(n3922), .A2(n3919), .ZN(n35088) );
  NAND2_X1 U14236 ( .A1(n3921), .A2(n32486), .ZN(n3920) );
  NAND3_X1 U14237 ( .A1(n31204), .A2(n3923), .A3(n32484), .ZN(n3922) );
  NAND2_X1 U14238 ( .A1(n8343), .A2(n8344), .ZN(n31003) );
  XNOR2_X1 U14239 ( .A(n34070), .B(n34364), .ZN(n3925) );
  XNOR2_X2 U14240 ( .A(n3925), .B(n3924), .ZN(n36027) );
  XNOR2_X1 U14241 ( .A(n34340), .B(n36800), .ZN(n3926) );
  INV_X1 U14242 ( .A(n36458), .ZN(n3927) );
  XNOR2_X1 U14243 ( .A(n33326), .B(n2154), .ZN(n32372) );
  NAND3_X1 U14244 ( .A1(n28840), .A2(n29747), .A3(n28830), .ZN(n28831) );
  NAND3_X1 U14246 ( .A1(n45511), .A2(n48831), .A3(n52091), .ZN(n45512) );
  XNOR2_X1 U14247 ( .A(n28347), .B(n3928), .ZN(n27313) );
  XNOR2_X1 U14248 ( .A(n27307), .B(n27308), .ZN(n3928) );
  NAND3_X1 U14249 ( .A1(n4215), .A2(n45518), .A3(n4214), .ZN(n4524) );
  NAND2_X1 U14252 ( .A1(n3931), .A2(n4069), .ZN(n4057) );
  NAND2_X1 U14253 ( .A1(n7022), .A2(n7021), .ZN(n3931) );
  NAND2_X1 U14254 ( .A1(n4080), .A2(n12353), .ZN(n3932) );
  NAND2_X1 U14256 ( .A1(n44823), .A2(n45817), .ZN(n3933) );
  NAND4_X1 U14257 ( .A1(n3935), .A2(n35572), .A3(n37532), .A4(n38494), .ZN(
        n35574) );
  NAND2_X1 U14258 ( .A1(n37520), .A2(n38506), .ZN(n3935) );
  AND2_X1 U14259 ( .A1(n41294), .A2(n41295), .ZN(n8583) );
  AND2_X1 U14260 ( .A1(n9801), .A2(n13225), .ZN(n5009) );
  AOI22_X1 U14261 ( .A1(n12904), .A2(n14191), .B1(n12905), .B2(n12906), .ZN(
        n12909) );
  INV_X1 U14263 ( .A(n35360), .ZN(n8503) );
  AND2_X1 U14264 ( .A1(n21574), .A2(n21409), .ZN(n7220) );
  INV_X1 U14265 ( .A(n33461), .ZN(n39340) );
  INV_X1 U14266 ( .A(n9291), .ZN(n10077) );
  INV_X1 U14268 ( .A(n12338), .ZN(n10277) );
  INV_X1 U14269 ( .A(n7577), .ZN(n49232) );
  INV_X1 U14270 ( .A(n13530), .ZN(n12938) );
  OAI21_X1 U14271 ( .B1(n9874), .B2(n7727), .A(n7726), .ZN(n8568) );
  XNOR2_X1 U14272 ( .A(n45081), .B(n46095), .ZN(n45771) );
  NAND2_X1 U14274 ( .A1(n23105), .A2(n22768), .ZN(n22771) );
  NAND2_X1 U14276 ( .A1(n38189), .A2(n38173), .ZN(n38175) );
  INV_X1 U14279 ( .A(n28297), .ZN(n7722) );
  INV_X1 U14280 ( .A(n12315), .ZN(n10945) );
  INV_X1 U14281 ( .A(n22868), .ZN(n19616) );
  INV_X1 U14282 ( .A(n11112), .ZN(n11113) );
  AND2_X1 U14285 ( .A1(n15925), .A2(n18867), .ZN(n4596) );
  NAND2_X1 U14287 ( .A1(n38592), .A2(n3940), .ZN(n36123) );
  NAND2_X1 U14289 ( .A1(n3942), .A2(n13104), .ZN(n12919) );
  AOI21_X1 U14290 ( .B1(n13090), .B2(n13075), .A(n3943), .ZN(n3942) );
  INV_X1 U14291 ( .A(n49841), .ZN(n49828) );
  NAND2_X2 U14292 ( .A1(n49705), .A2(n49706), .ZN(n49841) );
  NAND2_X1 U14293 ( .A1(n3945), .A2(n33884), .ZN(n33885) );
  NAND2_X1 U14294 ( .A1(n41788), .A2(n5604), .ZN(n3945) );
  NAND3_X1 U14296 ( .A1(n38637), .A2(n38628), .A3(n38635), .ZN(n3947) );
  XNOR2_X2 U14297 ( .A(n8913), .B(Key[67]), .ZN(n10831) );
  NAND2_X1 U14298 ( .A1(n31679), .A2(n29998), .ZN(n30975) );
  NAND2_X1 U14299 ( .A1(n45628), .A2(n46464), .ZN(n48539) );
  INV_X1 U14300 ( .A(n20421), .ZN(n19173) );
  NAND2_X1 U14301 ( .A1(n20427), .A2(n20359), .ZN(n20421) );
  OAI21_X1 U14302 ( .B1(n11255), .B2(n11258), .A(n3948), .ZN(n11257) );
  AND2_X2 U14303 ( .A1(n28650), .A2(n29260), .ZN(n29264) );
  NAND2_X1 U14304 ( .A1(n29802), .A2(n28508), .ZN(n28963) );
  AOI22_X1 U14305 ( .A1(n14477), .A2(n13856), .B1(n13559), .B2(n3949), .ZN(
        n9727) );
  NAND2_X1 U14306 ( .A1(n22901), .A2(n22359), .ZN(n22169) );
  NAND2_X1 U14307 ( .A1(n20656), .A2(n20270), .ZN(n20649) );
  NAND2_X1 U14308 ( .A1(n24277), .A2(n3950), .ZN(n7706) );
  NAND3_X1 U14309 ( .A1(n28904), .A2(n28583), .A3(n28895), .ZN(n27996) );
  NAND2_X1 U14310 ( .A1(n32596), .A2(n3952), .ZN(n28170) );
  NOR2_X1 U14311 ( .A1(n3954), .A2(n3953), .ZN(n50422) );
  NAND3_X1 U14312 ( .A1(n50410), .A2(n50441), .A3(n50409), .ZN(n3953) );
  INV_X1 U14313 ( .A(n50411), .ZN(n3954) );
  INV_X1 U14315 ( .A(n36267), .ZN(n36266) );
  XNOR2_X1 U14316 ( .A(n16937), .B(n15616), .ZN(n8488) );
  NOR2_X1 U14318 ( .A1(n358), .A2(n5923), .ZN(n5922) );
  OAI21_X1 U14319 ( .B1(n15986), .B2(n21631), .A(n18729), .ZN(n6728) );
  OAI211_X1 U14320 ( .C1(n26856), .C2(n26864), .A(n24683), .B(n26860), .ZN(
        n23857) );
  NAND4_X1 U14321 ( .A1(n47999), .A2(n3956), .A3(n47998), .A4(n3955), .ZN(
        n48001) );
  NAND2_X1 U14322 ( .A1(n47994), .A2(n52056), .ZN(n3955) );
  NAND2_X1 U14323 ( .A1(n47992), .A2(n47991), .ZN(n3957) );
  XNOR2_X2 U14324 ( .A(n16571), .B(n17947), .ZN(n18701) );
  NAND2_X1 U14325 ( .A1(n48210), .A2(n3959), .ZN(n44691) );
  OAI22_X1 U14326 ( .A1(n27668), .A2(n27669), .B1(n27671), .B2(n27670), .ZN(
        n27673) );
  XNOR2_X2 U14327 ( .A(n24719), .B(n24720), .ZN(n27652) );
  NAND3_X1 U14328 ( .A1(n49624), .A2(n43178), .A3(n49988), .ZN(n43179) );
  NAND3_X1 U14329 ( .A1(n23696), .A2(n24328), .A3(n3960), .ZN(n23699) );
  XNOR2_X1 U14333 ( .A(n3962), .B(n43420), .ZN(Plaintext[120]) );
  INV_X1 U14334 ( .A(n27768), .ZN(n4298) );
  OAI21_X1 U14335 ( .B1(n11852), .B2(n11851), .A(n15375), .ZN(n7156) );
  NAND2_X1 U14336 ( .A1(n32207), .A2(n32194), .ZN(n3963) );
  NOR2_X1 U14337 ( .A1(n18848), .A2(n18849), .ZN(n18855) );
  OAI21_X1 U14338 ( .B1(n23434), .B2(n23435), .A(n5610), .ZN(n23437) );
  NAND2_X1 U14339 ( .A1(n23442), .A2(n22593), .ZN(n23435) );
  NAND2_X1 U14340 ( .A1(n3965), .A2(n30435), .ZN(n30428) );
  NAND2_X1 U14341 ( .A1(n30424), .A2(n30434), .ZN(n3965) );
  XNOR2_X1 U14342 ( .A(n28262), .B(n8723), .ZN(n3966) );
  INV_X1 U14343 ( .A(n20119), .ZN(n19538) );
  INV_X1 U14344 ( .A(n50982), .ZN(n7317) );
  MUX2_X1 U14345 ( .A(n32898), .B(n32897), .S(n32896), .Z(n32905) );
  NAND2_X1 U14347 ( .A1(n19467), .A2(n3968), .ZN(n21281) );
  NAND2_X1 U14348 ( .A1(n19783), .A2(n8441), .ZN(n19467) );
  OR2_X1 U14349 ( .A1(n47404), .A2(n46530), .ZN(n7058) );
  NAND3_X1 U14350 ( .A1(n46437), .A2(n46436), .A3(n2416), .ZN(n46438) );
  NAND2_X1 U14351 ( .A1(n19328), .A2(n20428), .ZN(n3970) );
  OR2_X1 U14352 ( .A1(n11089), .A2(n11443), .ZN(n8948) );
  INV_X1 U14353 ( .A(n28764), .ZN(n30382) );
  INV_X1 U14354 ( .A(n32540), .ZN(n5976) );
  INV_X1 U14355 ( .A(n26677), .ZN(n29494) );
  XNOR2_X1 U14356 ( .A(n37133), .B(n7318), .ZN(n36754) );
  INV_X1 U14357 ( .A(n36869), .ZN(n7298) );
  INV_X1 U14358 ( .A(n15161), .ZN(n5113) );
  INV_X1 U14359 ( .A(n49717), .ZN(n42957) );
  XNOR2_X1 U14360 ( .A(n26032), .B(n24494), .ZN(n7945) );
  NAND3_X1 U14361 ( .A1(n29800), .A2(n28962), .A3(n5057), .ZN(n28498) );
  NOR2_X1 U14362 ( .A1(n31346), .A2(n30037), .ZN(n30054) );
  NAND2_X1 U14363 ( .A1(n21448), .A2(n5500), .ZN(n3972) );
  NAND2_X1 U14364 ( .A1(n8479), .A2(n39010), .ZN(n3973) );
  OAI21_X1 U14365 ( .B1(n31822), .B2(n31826), .A(n3974), .ZN(n30573) );
  NAND3_X1 U14366 ( .A1(n31829), .A2(n30849), .A3(n31033), .ZN(n3974) );
  NAND3_X2 U14367 ( .A1(n7618), .A2(n23091), .A3(n7619), .ZN(n27373) );
  INV_X1 U14368 ( .A(n11710), .ZN(n11712) );
  XNOR2_X2 U14369 ( .A(n24792), .B(n5384), .ZN(n25883) );
  NAND4_X1 U14370 ( .A1(n46284), .A2(n3975), .A3(n46285), .A4(n46286), .ZN(
        n46296) );
  NAND2_X1 U14371 ( .A1(n46282), .A2(n46283), .ZN(n3975) );
  NAND2_X1 U14372 ( .A1(n3977), .A2(n3976), .ZN(n38150) );
  NAND2_X1 U14373 ( .A1(n38148), .A2(n38149), .ZN(n3976) );
  NAND2_X1 U14374 ( .A1(n38144), .A2(n38143), .ZN(n3978) );
  NAND2_X1 U14376 ( .A1(n8071), .A2(n39763), .ZN(n3979) );
  NAND2_X1 U14377 ( .A1(n29846), .A2(n29847), .ZN(n32628) );
  XNOR2_X2 U14378 ( .A(Key[104]), .B(Ciphertext[85]), .ZN(n11608) );
  NAND2_X1 U14379 ( .A1(n50352), .A2(n47294), .ZN(n7177) );
  AOI21_X1 U14381 ( .B1(n41943), .B2(n41944), .A(n6545), .ZN(n6544) );
  NAND2_X1 U14382 ( .A1(n6013), .A2(n30592), .ZN(n30915) );
  NAND4_X1 U14383 ( .A1(n3981), .A2(n37446), .A3(n36155), .A4(n35968), .ZN(
        n35969) );
  NAND2_X1 U14384 ( .A1(n35967), .A2(n38532), .ZN(n3981) );
  NAND3_X1 U14385 ( .A1(n47213), .A2(n47212), .A3(n47606), .ZN(n47214) );
  NAND3_X1 U14386 ( .A1(n19848), .A2(n19870), .A3(n19874), .ZN(n4371) );
  NAND3_X2 U14387 ( .A1(n3982), .A2(n37463), .A3(n5422), .ZN(n43123) );
  OR2_X1 U14389 ( .A1(n21215), .A2(n19819), .ZN(n19737) );
  NAND2_X1 U14390 ( .A1(n7645), .A2(n8183), .ZN(n8182) );
  NAND2_X1 U14391 ( .A1(n28713), .A2(n29270), .ZN(n3983) );
  NOR2_X1 U14395 ( .A1(n30322), .A2(n8746), .ZN(n30336) );
  XNOR2_X1 U14396 ( .A(n34141), .B(n3986), .ZN(n32757) );
  NAND4_X2 U14397 ( .A1(n5003), .A2(n3987), .A3(n11827), .A4(n11828), .ZN(
        n18690) );
  NOR2_X1 U14398 ( .A1(n6377), .A2(n22729), .ZN(n6376) );
  AND2_X1 U14399 ( .A1(n34211), .A2(n34212), .ZN(n6714) );
  INV_X1 U14400 ( .A(n13282), .ZN(n15245) );
  INV_X1 U14401 ( .A(n26092), .ZN(n6922) );
  NAND2_X1 U14402 ( .A1(n23924), .A2(n23895), .ZN(n23921) );
  OAI21_X1 U14403 ( .B1(n20195), .B2(n20194), .A(n6929), .ZN(n20196) );
  OAI22_X1 U14405 ( .A1(n15178), .A2(n5766), .B1(n13459), .B2(n6320), .ZN(
        n4443) );
  NAND3_X1 U14408 ( .A1(n48158), .A2(n48156), .A3(n48157), .ZN(n3990) );
  XNOR2_X1 U14409 ( .A(n51664), .B(n34839), .ZN(n8022) );
  OAI21_X2 U14410 ( .B1(n27974), .B2(n27973), .A(n27972), .ZN(n31746) );
  AOI21_X1 U14411 ( .B1(n3993), .B2(n3992), .A(n49933), .ZN(n3991) );
  INV_X1 U14412 ( .A(n49909), .ZN(n3992) );
  INV_X1 U14413 ( .A(n47425), .ZN(n3993) );
  OAI21_X1 U14414 ( .B1(n46179), .B2(n47423), .A(n49934), .ZN(n3994) );
  INV_X1 U14415 ( .A(n23307), .ZN(n22957) );
  NAND2_X1 U14416 ( .A1(n21227), .A2(n3995), .ZN(n17314) );
  NAND2_X1 U14417 ( .A1(n8246), .A2(n8910), .ZN(n3996) );
  INV_X1 U14419 ( .A(n41553), .ZN(n6505) );
  INV_X1 U14420 ( .A(n22535), .ZN(n22541) );
  NAND3_X2 U14421 ( .A1(n7959), .A2(n3998), .A3(n7960), .ZN(n35468) );
  NAND2_X1 U14422 ( .A1(n19529), .A2(n19826), .ZN(n5273) );
  NAND2_X1 U14423 ( .A1(n21531), .A2(n21530), .ZN(n6165) );
  NAND2_X1 U14424 ( .A1(n23871), .A2(n22605), .ZN(n6718) );
  INV_X1 U14425 ( .A(n34313), .ZN(n36067) );
  NAND2_X1 U14426 ( .A1(n46901), .A2(n3999), .ZN(n46900) );
  NOR2_X2 U14427 ( .A1(n45585), .A2(n45586), .ZN(n46542) );
  NAND2_X1 U14428 ( .A1(n20415), .A2(n5923), .ZN(n21375) );
  NAND3_X1 U14429 ( .A1(n21380), .A2(n21381), .A3(n4002), .ZN(n4001) );
  NAND2_X1 U14430 ( .A1(n48411), .A2(n4003), .ZN(n45581) );
  NAND2_X1 U14431 ( .A1(n4004), .A2(n2738), .ZN(n4236) );
  NAND2_X1 U14432 ( .A1(n40248), .A2(n40247), .ZN(n4004) );
  XNOR2_X1 U14433 ( .A(n28250), .B(n4293), .ZN(n25338) );
  NOR2_X1 U14434 ( .A1(n27619), .A2(n26803), .ZN(n27739) );
  NAND3_X1 U14435 ( .A1(n13844), .A2(n13856), .A3(n9690), .ZN(n9692) );
  XNOR2_X1 U14436 ( .A(n4005), .B(n33940), .ZN(n33941) );
  XNOR2_X1 U14437 ( .A(n37021), .B(n34078), .ZN(n4005) );
  NAND2_X1 U14438 ( .A1(n50863), .A2(n50886), .ZN(n50864) );
  OAI21_X1 U14439 ( .B1(n9919), .B2(n9920), .A(n10609), .ZN(n4006) );
  AOI21_X1 U14440 ( .B1(n4007), .B2(n14791), .A(n14790), .ZN(n14792) );
  NAND3_X1 U14441 ( .A1(n45976), .A2(n49445), .A3(n49442), .ZN(n47202) );
  NAND2_X1 U14442 ( .A1(n10418), .A2(n52132), .ZN(n4008) );
  NAND2_X1 U14443 ( .A1(n32244), .A2(n32254), .ZN(n29364) );
  NAND2_X1 U14444 ( .A1(n4332), .A2(n41112), .ZN(n40468) );
  NAND3_X2 U14445 ( .A1(n5194), .A2(n5193), .A3(n5198), .ZN(n21756) );
  NAND2_X1 U14446 ( .A1(n4010), .A2(n2520), .ZN(n5140) );
  NAND2_X1 U14447 ( .A1(n27715), .A2(n29407), .ZN(n4010) );
  NAND2_X1 U14448 ( .A1(n30602), .A2(n30592), .ZN(n29687) );
  NOR2_X1 U14449 ( .A1(n4014), .A2(n4013), .ZN(n4012) );
  OAI22_X1 U14450 ( .A1(n7326), .A2(n10935), .B1(n10214), .B2(n10929), .ZN(
        n4013) );
  XNOR2_X1 U14451 ( .A(n34487), .B(n35404), .ZN(n6018) );
  AOI21_X1 U14452 ( .B1(n6344), .B2(n32601), .A(n712), .ZN(n7147) );
  NAND2_X1 U14453 ( .A1(n21435), .A2(n19156), .ZN(n19955) );
  OAI21_X1 U14454 ( .B1(n9738), .B2(n10678), .A(n10676), .ZN(n5994) );
  INV_X1 U14457 ( .A(Ciphertext[166]), .ZN(n4015) );
  MUX2_X1 U14458 ( .A(n9860), .B(n10956), .S(n10965), .Z(n13227) );
  NAND3_X1 U14459 ( .A1(n9742), .A2(n9741), .A3(n4273), .ZN(n5831) );
  NAND2_X1 U14460 ( .A1(n30071), .A2(n31121), .ZN(n26969) );
  OAI21_X1 U14461 ( .B1(n6829), .B2(n38370), .A(n4016), .ZN(n6828) );
  INV_X1 U14462 ( .A(n382), .ZN(n6188) );
  NAND2_X1 U14464 ( .A1(n21771), .A2(n21782), .ZN(n4017) );
  NAND2_X1 U14465 ( .A1(n4019), .A2(n4018), .ZN(n30728) );
  NAND2_X1 U14466 ( .A1(n30720), .A2(n30719), .ZN(n4018) );
  NAND2_X1 U14467 ( .A1(n4021), .A2(n4020), .ZN(n4019) );
  INV_X1 U14468 ( .A(n30719), .ZN(n4020) );
  NAND3_X1 U14469 ( .A1(n30717), .A2(n30724), .A3(n30716), .ZN(n4021) );
  INV_X1 U14470 ( .A(n6201), .ZN(n6200) );
  NAND2_X1 U14472 ( .A1(n30692), .A2(n29933), .ZN(n30694) );
  XNOR2_X2 U14473 ( .A(n7074), .B(n24087), .ZN(n30692) );
  NAND2_X1 U14474 ( .A1(n5593), .A2(n39291), .ZN(n39307) );
  XNOR2_X1 U14475 ( .A(n18396), .B(n18397), .ZN(n4022) );
  NAND3_X1 U14476 ( .A1(n13938), .A2(n13937), .A3(n4023), .ZN(n13956) );
  NAND2_X1 U14477 ( .A1(n4024), .A2(n13207), .ZN(n4023) );
  NAND4_X1 U14478 ( .A1(n12070), .A2(n12071), .A3(n51433), .A4(n12635), .ZN(
        n12072) );
  OR2_X1 U14479 ( .A1(n23834), .A2(n23821), .ZN(n4025) );
  NAND2_X1 U14481 ( .A1(n12660), .A2(n10457), .ZN(n10444) );
  NAND3_X1 U14482 ( .A1(n7494), .A2(n354), .A3(n22107), .ZN(n5701) );
  INV_X1 U14483 ( .A(n31387), .ZN(n6197) );
  OAI21_X1 U14484 ( .B1(n6253), .B2(n4267), .A(n30399), .ZN(n30400) );
  XNOR2_X2 U14485 ( .A(n16644), .B(n16643), .ZN(n19510) );
  XNOR2_X1 U14486 ( .A(n4027), .B(n17942), .ZN(n17946) );
  XNOR2_X1 U14487 ( .A(n17940), .B(n17941), .ZN(n4027) );
  XNOR2_X1 U14488 ( .A(n4028), .B(n16627), .ZN(n18770) );
  XNOR2_X1 U14489 ( .A(n16626), .B(n16625), .ZN(n4028) );
  INV_X1 U14490 ( .A(n46872), .ZN(n7332) );
  OAI22_X1 U14493 ( .A1(n21582), .A2(n21583), .B1(n21585), .B2(n21584), .ZN(
        n21586) );
  OAI21_X1 U14494 ( .B1(n7273), .B2(n5429), .A(n48461), .ZN(n7272) );
  INV_X1 U14496 ( .A(n40423), .ZN(n5436) );
  NAND2_X1 U14497 ( .A1(n23100), .A2(n22874), .ZN(n19882) );
  INV_X1 U14498 ( .A(n24026), .ZN(n24036) );
  AND2_X1 U14499 ( .A1(n31196), .A2(n31199), .ZN(n5746) );
  NOR2_X1 U14500 ( .A1(n19818), .A2(n2239), .ZN(n7265) );
  OR2_X1 U14501 ( .A1(n31195), .A2(n32501), .ZN(n4411) );
  NOR2_X1 U14502 ( .A1(n8126), .A2(n8127), .ZN(n14649) );
  AND2_X1 U14503 ( .A1(n19180), .A2(n7233), .ZN(n5646) );
  OR2_X1 U14504 ( .A1(n13438), .A2(n12894), .ZN(n13436) );
  INV_X1 U14505 ( .A(n25927), .ZN(n7103) );
  OR2_X1 U14506 ( .A1(n12903), .A2(n14190), .ZN(n12902) );
  INV_X1 U14507 ( .A(n19344), .ZN(n20503) );
  INV_X1 U14508 ( .A(n32242), .ZN(n31244) );
  AOI22_X1 U14509 ( .A1(n5833), .A2(n50992), .B1(n52381), .B2(n19563), .ZN(
        n19571) );
  INV_X1 U14510 ( .A(n49274), .ZN(n45670) );
  INV_X1 U14511 ( .A(n33470), .ZN(n37072) );
  XNOR2_X1 U14512 ( .A(n17837), .B(n17836), .ZN(n17856) );
  INV_X1 U14513 ( .A(n15077), .ZN(n7571) );
  XNOR2_X1 U14514 ( .A(n33306), .B(n52164), .ZN(n35747) );
  AOI21_X1 U14515 ( .B1(n6390), .B2(n48990), .A(n51310), .ZN(n6386) );
  XNOR2_X1 U14516 ( .A(n4030), .B(n47890), .ZN(Plaintext[29]) );
  NAND2_X1 U14518 ( .A1(n36093), .A2(n4032), .ZN(n36096) );
  INV_X1 U14519 ( .A(n4033), .ZN(n4032) );
  OAI21_X1 U14520 ( .B1(n40114), .B2(n40120), .A(n40203), .ZN(n4033) );
  NAND2_X1 U14521 ( .A1(n23755), .A2(n24180), .ZN(n24189) );
  INV_X1 U14522 ( .A(n41283), .ZN(n39730) );
  NAND2_X1 U14523 ( .A1(n41275), .A2(n41029), .ZN(n41283) );
  NAND3_X1 U14524 ( .A1(n36609), .A2(n36616), .A3(n34313), .ZN(n34311) );
  NAND2_X1 U14525 ( .A1(n34650), .A2(n51015), .ZN(n34313) );
  XNOR2_X1 U14526 ( .A(n35265), .B(n33190), .ZN(n33191) );
  XNOR2_X2 U14527 ( .A(n37062), .B(n36932), .ZN(n35265) );
  NAND2_X1 U14531 ( .A1(n4037), .A2(n4036), .ZN(n36039) );
  NAND2_X1 U14532 ( .A1(n36552), .A2(n37965), .ZN(n4036) );
  NAND2_X1 U14533 ( .A1(n37964), .A2(n36540), .ZN(n4037) );
  NOR2_X1 U14534 ( .A1(n4038), .A2(n5240), .ZN(n5241) );
  AND2_X1 U14535 ( .A1(n30208), .A2(n30207), .ZN(n4038) );
  NAND2_X1 U14537 ( .A1(n1467), .A2(n50679), .ZN(n50717) );
  OAI211_X1 U14538 ( .C1(n40964), .C2(n51394), .A(n40962), .B(n40961), .ZN(
        n4040) );
  NAND2_X1 U14539 ( .A1(n6047), .A2(n51432), .ZN(n12638) );
  NAND2_X1 U14541 ( .A1(n3075), .A2(n51092), .ZN(n48085) );
  AOI22_X1 U14543 ( .A1(n4043), .A2(n48465), .B1(n48467), .B2(n48466), .ZN(
        n48472) );
  NAND2_X1 U14544 ( .A1(n48464), .A2(n48463), .ZN(n4043) );
  NAND3_X1 U14545 ( .A1(n7452), .A2(n44454), .A3(n44455), .ZN(n44456) );
  NAND3_X1 U14546 ( .A1(n44110), .A2(n45176), .A3(n399), .ZN(n7452) );
  NAND2_X1 U14548 ( .A1(n39554), .A2(n40194), .ZN(n39555) );
  INV_X1 U14549 ( .A(n22898), .ZN(n22896) );
  NAND2_X1 U14550 ( .A1(n32634), .A2(n32900), .ZN(n32918) );
  NAND3_X1 U14551 ( .A1(n15100), .A2(n15112), .A3(n15101), .ZN(n4249) );
  OAI211_X1 U14552 ( .C1(n11625), .C2(n11629), .A(n4508), .B(n11466), .ZN(
        n10845) );
  NAND2_X1 U14553 ( .A1(n9773), .A2(n9762), .ZN(n12308) );
  NAND3_X2 U14554 ( .A1(n32191), .A2(n4044), .A3(n32189), .ZN(n35333) );
  INV_X1 U14555 ( .A(Ciphertext[160]), .ZN(n7563) );
  INV_X1 U14556 ( .A(n11875), .ZN(n11497) );
  NAND2_X1 U14557 ( .A1(n5361), .A2(n19674), .ZN(n16998) );
  NAND2_X1 U14558 ( .A1(n40450), .A2(n40403), .ZN(n39737) );
  NAND2_X1 U14559 ( .A1(n21899), .A2(n23507), .ZN(n23508) );
  NAND4_X1 U14560 ( .A1(n22404), .A2(n22401), .A3(n22402), .A4(n418), .ZN(
        n4047) );
  NAND2_X1 U14561 ( .A1(n22072), .A2(n22201), .ZN(n22088) );
  NAND4_X2 U14562 ( .A1(n20341), .A2(n20342), .A3(n20339), .A4(n20340), .ZN(
        n22748) );
  OR2_X1 U14563 ( .A1(n39233), .A2(n37283), .ZN(n4675) );
  NAND3_X1 U14564 ( .A1(n19668), .A2(n19669), .A3(n4049), .ZN(n19709) );
  NAND2_X1 U14565 ( .A1(n19637), .A2(n18942), .ZN(n4049) );
  NAND2_X2 U14566 ( .A1(n4050), .A2(n7628), .ZN(n26152) );
  INV_X1 U14567 ( .A(n4052), .ZN(n4051) );
  OAI21_X1 U14568 ( .B1(n22742), .B2(n22732), .A(n22390), .ZN(n4052) );
  NAND2_X1 U14569 ( .A1(n27610), .A2(n4053), .ZN(n27611) );
  NAND2_X1 U14570 ( .A1(n27608), .A2(n4054), .ZN(n4053) );
  INV_X1 U14571 ( .A(n11030), .ZN(n8410) );
  NAND4_X1 U14572 ( .A1(n47508), .A2(n5993), .A3(n4055), .A4(n47506), .ZN(
        n47510) );
  NOR2_X1 U14573 ( .A1(n37942), .A2(n39270), .ZN(n39011) );
  NAND2_X1 U14574 ( .A1(n21369), .A2(n20805), .ZN(n21393) );
  AND2_X1 U14575 ( .A1(n47786), .A2(n47777), .ZN(n47743) );
  OR2_X1 U14576 ( .A1(n23193), .A2(n23194), .ZN(n23198) );
  NAND2_X2 U14579 ( .A1(n4056), .A2(n8328), .ZN(n13514) );
  INV_X1 U14580 ( .A(n26552), .ZN(n27226) );
  INV_X1 U14582 ( .A(n8051), .ZN(n5920) );
  NAND4_X2 U14583 ( .A1(n20667), .A2(n20666), .A3(n20665), .A4(n20664), .ZN(
        n23531) );
  XNOR2_X1 U14586 ( .A(n7102), .B(n51448), .ZN(n43660) );
  INV_X1 U14587 ( .A(n11409), .ZN(n12139) );
  INV_X1 U14588 ( .A(n40822), .ZN(n40817) );
  INV_X1 U14589 ( .A(Ciphertext[133]), .ZN(n4771) );
  OR2_X1 U14590 ( .A1(n10956), .A2(n10955), .ZN(n9852) );
  XNOR2_X1 U14591 ( .A(n24308), .B(n8385), .ZN(n24354) );
  INV_X1 U14592 ( .A(n12705), .ZN(n12702) );
  INV_X1 U14593 ( .A(n37430), .ZN(n37491) );
  INV_X1 U14594 ( .A(n18847), .ZN(n21657) );
  INV_X1 U14595 ( .A(n14672), .ZN(n13629) );
  INV_X1 U14596 ( .A(n22145), .ZN(n8695) );
  INV_X1 U14597 ( .A(n31113), .ZN(n7957) );
  XNOR2_X1 U14598 ( .A(n28349), .B(n28348), .ZN(n28449) );
  XNOR2_X2 U14599 ( .A(n42639), .B(n44571), .ZN(n49197) );
  XNOR2_X2 U14600 ( .A(n45305), .B(n45445), .ZN(n43751) );
  NAND3_X2 U14601 ( .A1(n39624), .A2(n39623), .A3(n39625), .ZN(n45305) );
  NAND2_X1 U14602 ( .A1(n17509), .A2(n5195), .ZN(n4058) );
  OR3_X1 U14603 ( .A1(n26944), .A2(n51117), .A3(n27652), .ZN(n26948) );
  NAND2_X1 U14605 ( .A1(n24183), .A2(n4060), .ZN(n24177) );
  INV_X1 U14606 ( .A(Ciphertext[125]), .ZN(n7415) );
  OAI22_X1 U14607 ( .A1(n22504), .A2(n22498), .B1(n22834), .B2(n22497), .ZN(
        n22499) );
  NAND2_X1 U14608 ( .A1(n1145), .A2(n22830), .ZN(n22504) );
  NAND2_X1 U14609 ( .A1(n29530), .A2(n29531), .ZN(n29537) );
  INV_X1 U14612 ( .A(n21605), .ZN(n4063) );
  INV_X1 U14613 ( .A(n32510), .ZN(n5158) );
  NAND2_X1 U14614 ( .A1(n6847), .A2(n37696), .ZN(n4064) );
  NAND2_X1 U14615 ( .A1(n18072), .A2(n18330), .ZN(n14385) );
  XOR2_X1 U14616 ( .A(n13770), .B(n16330), .Z(n8176) );
  XNOR2_X1 U14617 ( .A(n17671), .B(n16024), .ZN(n15800) );
  NAND3_X1 U14618 ( .A1(n21548), .A2(n21540), .A3(n21541), .ZN(n21546) );
  NAND2_X1 U14619 ( .A1(n15263), .A2(n14783), .ZN(n11055) );
  NAND2_X1 U14620 ( .A1(n20376), .A2(n20795), .ZN(n20791) );
  NAND3_X1 U14621 ( .A1(n20891), .A2(n23426), .A3(n23412), .ZN(n20892) );
  INV_X1 U14622 ( .A(n27860), .ZN(n25841) );
  NAND2_X1 U14624 ( .A1(n5120), .A2(n11408), .ZN(n11399) );
  NAND2_X1 U14625 ( .A1(n36410), .A2(n51334), .ZN(n37632) );
  AND3_X1 U14627 ( .A1(n22633), .A2(n22631), .A3(n22632), .ZN(n4066) );
  AND2_X2 U14628 ( .A1(n4067), .A2(n17088), .ZN(n17418) );
  NAND2_X1 U14630 ( .A1(n23950), .A2(n22623), .ZN(n22624) );
  NAND2_X1 U14632 ( .A1(n21269), .A2(n51013), .ZN(n19466) );
  INV_X1 U14634 ( .A(n11825), .ZN(n4071) );
  NAND2_X1 U14635 ( .A1(n13089), .A2(n12914), .ZN(n11825) );
  NAND3_X1 U14636 ( .A1(n5718), .A2(n29639), .A3(n29638), .ZN(n32644) );
  NOR2_X1 U14637 ( .A1(n49597), .A2(n4072), .ZN(n49591) );
  NAND3_X2 U14638 ( .A1(n4074), .A2(n11060), .A3(n4073), .ZN(n18466) );
  INV_X1 U14639 ( .A(n29520), .ZN(n29519) );
  MUX2_X1 U14640 ( .A(n36610), .B(n36057), .S(n36065), .Z(n34923) );
  INV_X1 U14642 ( .A(n17351), .ZN(n8033) );
  INV_X1 U14643 ( .A(n22716), .ZN(n20548) );
  XOR2_X1 U14644 ( .A(n16925), .B(n16924), .Z(n8034) );
  INV_X1 U14645 ( .A(n38998), .ZN(n6825) );
  NAND2_X1 U14646 ( .A1(n10179), .A2(n4077), .ZN(n9457) );
  NAND2_X1 U14647 ( .A1(n42145), .A2(n42136), .ZN(n41760) );
  XNOR2_X2 U14648 ( .A(n18167), .B(n18166), .ZN(n19801) );
  OAI21_X1 U14649 ( .B1(n4079), .B2(n4078), .A(n50703), .ZN(n4303) );
  NAND4_X4 U14651 ( .A1(n9470), .A2(n9467), .A3(n9469), .A4(n9468), .ZN(n13091) );
  INV_X1 U14652 ( .A(n20157), .ZN(n4081) );
  INV_X1 U14654 ( .A(n14452), .ZN(n5652) );
  AOI22_X1 U14655 ( .A1(n11394), .A2(n12053), .B1(n6464), .B2(n10665), .ZN(
        n11396) );
  NAND3_X1 U14656 ( .A1(n30235), .A2(n29255), .A3(n29252), .ZN(n25637) );
  NAND2_X1 U14657 ( .A1(n28641), .A2(n383), .ZN(n29331) );
  INV_X1 U14658 ( .A(n39451), .ZN(n39442) );
  NOR2_X1 U14661 ( .A1(n38182), .A2(n38183), .ZN(n4083) );
  NAND2_X1 U14662 ( .A1(n723), .A2(n32356), .ZN(n32047) );
  NAND3_X1 U14663 ( .A1(n5780), .A2(n5779), .A3(n31949), .ZN(n4084) );
  XNOR2_X1 U14664 ( .A(n23894), .B(n23930), .ZN(n8443) );
  NOR2_X1 U14665 ( .A1(n21976), .A2(n23483), .ZN(n23490) );
  XNOR2_X1 U14666 ( .A(n39591), .B(n39590), .ZN(n39811) );
  AND3_X1 U14668 ( .A1(n30238), .A2(n30237), .A3(n30236), .ZN(n7065) );
  OR2_X1 U14669 ( .A1(n24244), .A2(n20875), .ZN(n21815) );
  AND2_X1 U14670 ( .A1(n10925), .A2(n9807), .ZN(n10922) );
  OR2_X1 U14671 ( .A1(n29715), .A2(n28983), .ZN(n28183) );
  XNOR2_X1 U14672 ( .A(n4086), .B(n17175), .ZN(n15888) );
  XNOR2_X1 U14673 ( .A(n15876), .B(n4762), .ZN(n4086) );
  XNOR2_X1 U14674 ( .A(n6732), .B(n23893), .ZN(n24092) );
  INV_X1 U14675 ( .A(n28025), .ZN(n26467) );
  NAND3_X1 U14676 ( .A1(n9907), .A2(n9922), .A3(n9908), .ZN(n9910) );
  NOR2_X1 U14677 ( .A1(n36606), .A2(n8090), .ZN(n34653) );
  NAND2_X1 U14678 ( .A1(n9289), .A2(n9291), .ZN(n10610) );
  NAND4_X1 U14680 ( .A1(n5557), .A2(n5559), .A3(n5560), .A4(n19435), .ZN(
        n21016) );
  AND2_X1 U14681 ( .A1(n52193), .A2(n41286), .ZN(n40412) );
  NAND2_X1 U14683 ( .A1(n695), .A2(n34189), .ZN(n34193) );
  INV_X1 U14684 ( .A(n24283), .ZN(n21085) );
  AND2_X1 U14685 ( .A1(n37533), .A2(n34679), .ZN(n7377) );
  NAND3_X1 U14686 ( .A1(n4087), .A2(n23514), .A3(n23515), .ZN(n23516) );
  NOR2_X1 U14688 ( .A1(n8550), .A2(n8549), .ZN(n7923) );
  INV_X1 U14689 ( .A(n29261), .ZN(n29251) );
  INV_X1 U14690 ( .A(n41642), .ZN(n41985) );
  INV_X1 U14691 ( .A(n24289), .ZN(n23509) );
  INV_X1 U14692 ( .A(n22263), .ZN(n23334) );
  NOR2_X1 U14693 ( .A1(n19610), .A2(n22859), .ZN(n22868) );
  INV_X1 U14694 ( .A(n31384), .ZN(n8260) );
  XNOR2_X1 U14695 ( .A(n25605), .B(n25483), .ZN(n25291) );
  XNOR2_X1 U14696 ( .A(n42486), .B(n7623), .ZN(n40631) );
  NAND3_X2 U14697 ( .A1(n4088), .A2(n10654), .A3(n10653), .ZN(n18791) );
  NAND2_X1 U14698 ( .A1(n4089), .A2(n45242), .ZN(n45243) );
  AOI21_X2 U14701 ( .B1(n8973), .B2(n8972), .A(n8971), .ZN(n14982) );
  NAND2_X1 U14702 ( .A1(n4090), .A2(n12383), .ZN(n4307) );
  NAND3_X1 U14703 ( .A1(n12101), .A2(n6479), .A3(n9370), .ZN(n4090) );
  NAND3_X1 U14704 ( .A1(n35925), .A2(n37507), .A3(n4092), .ZN(n4091) );
  NAND4_X1 U14705 ( .A1(n4093), .A2(n48584), .A3(n48609), .A4(n48620), .ZN(
        n48586) );
  OAI22_X1 U14706 ( .A1(n48578), .A2(n48579), .B1(n48577), .B2(n48576), .ZN(
        n4093) );
  NOR2_X1 U14707 ( .A1(n7488), .A2(n40823), .ZN(n39693) );
  NOR2_X1 U14708 ( .A1(n11502), .A2(n7356), .ZN(n11503) );
  NAND2_X1 U14710 ( .A1(n39576), .A2(n43323), .ZN(n39616) );
  NAND3_X2 U14711 ( .A1(n7307), .A2(n7308), .A3(n37584), .ZN(n43323) );
  NAND3_X1 U14712 ( .A1(n4095), .A2(n36208), .A3(n36207), .ZN(n36211) );
  NAND2_X2 U14713 ( .A1(n50286), .A2(n8763), .ZN(n50482) );
  NAND2_X1 U14715 ( .A1(n6997), .A2(n4096), .ZN(n41875) );
  NAND2_X1 U14716 ( .A1(n39580), .A2(n39579), .ZN(n7002) );
  NAND3_X1 U14718 ( .A1(n39577), .A2(n40800), .A3(n41004), .ZN(n39578) );
  INV_X1 U14719 ( .A(n28031), .ZN(n28033) );
  NAND2_X1 U14720 ( .A1(n3368), .A2(n547), .ZN(n28031) );
  OAI21_X1 U14721 ( .B1(n19592), .B2(n4099), .A(n23467), .ZN(n21163) );
  OAI21_X1 U14722 ( .B1(n21957), .B2(n21948), .A(n21945), .ZN(n4099) );
  NAND3_X1 U14723 ( .A1(n29052), .A2(n29051), .A3(n31530), .ZN(n29074) );
  NAND3_X1 U14725 ( .A1(n34653), .A2(n36066), .A3(n36062), .ZN(n36623) );
  NAND2_X1 U14726 ( .A1(n30198), .A2(n30199), .ZN(n30201) );
  NAND3_X1 U14727 ( .A1(n6394), .A2(n31559), .A3(n31560), .ZN(n4100) );
  OAI22_X1 U14728 ( .A1(n11897), .A2(n12483), .B1(n12481), .B2(n12478), .ZN(
        n11069) );
  NAND2_X1 U14729 ( .A1(n8667), .A2(n11908), .ZN(n11897) );
  XNOR2_X1 U14732 ( .A(n15605), .B(n16896), .ZN(n8233) );
  OAI21_X1 U14733 ( .B1(n38476), .B2(n38475), .A(n38474), .ZN(n4103) );
  INV_X1 U14734 ( .A(n19891), .ZN(n6043) );
  NAND3_X1 U14737 ( .A1(n23155), .A2(n23464), .A3(n2076), .ZN(n23163) );
  NAND2_X1 U14738 ( .A1(n37917), .A2(n38697), .ZN(n4105) );
  NAND2_X1 U14739 ( .A1(n7157), .A2(n5552), .ZN(n4107) );
  NAND3_X2 U14741 ( .A1(n4109), .A2(n4108), .A3(n29646), .ZN(n35762) );
  INV_X1 U14742 ( .A(n4110), .ZN(n4109) );
  OAI21_X1 U14743 ( .B1(n29649), .B2(n29648), .A(n29645), .ZN(n4110) );
  XNOR2_X1 U14746 ( .A(n18700), .B(n7381), .ZN(n7380) );
  NAND3_X1 U14747 ( .A1(n18317), .A2(n16788), .A3(n18316), .ZN(n18320) );
  OAI21_X1 U14748 ( .B1(n29035), .B2(n28874), .A(n28879), .ZN(n28878) );
  NOR2_X2 U14749 ( .A1(n8364), .A2(n28882), .ZN(n28879) );
  INV_X1 U14750 ( .A(n39843), .ZN(n38613) );
  NAND3_X1 U14752 ( .A1(n45643), .A2(n45644), .A3(n49161), .ZN(n45645) );
  XNOR2_X2 U14753 ( .A(n24504), .B(n24503), .ZN(n29467) );
  AND3_X2 U14754 ( .A1(n4112), .A2(n16692), .A3(n16693), .ZN(n28126) );
  NAND2_X1 U14755 ( .A1(n16695), .A2(n16694), .ZN(n4112) );
  INV_X1 U14756 ( .A(n24116), .ZN(n23731) );
  XNOR2_X1 U14757 ( .A(n26551), .B(n8657), .ZN(n26553) );
  INV_X1 U14758 ( .A(n14485), .ZN(n14807) );
  NAND2_X1 U14759 ( .A1(n15380), .A2(n15358), .ZN(n14485) );
  XNOR2_X1 U14760 ( .A(n4114), .B(n45020), .ZN(Plaintext[19]) );
  NAND4_X1 U14761 ( .A1(n45019), .A2(n45018), .A3(n45016), .A4(n45017), .ZN(
        n4114) );
  XNOR2_X1 U14762 ( .A(n17249), .B(n2225), .ZN(n17250) );
  XNOR2_X2 U14763 ( .A(n33385), .B(n33384), .ZN(n35939) );
  NAND4_X1 U14764 ( .A1(n39831), .A2(n4115), .A3(n38623), .A4(n38622), .ZN(
        n38624) );
  NAND3_X1 U14765 ( .A1(n10047), .A2(n10962), .A3(n10965), .ZN(n9848) );
  NAND2_X1 U14766 ( .A1(n11279), .A2(n4118), .ZN(n9523) );
  NOR2_X1 U14767 ( .A1(n27539), .A2(n27542), .ZN(n4758) );
  NAND3_X1 U14768 ( .A1(n37910), .A2(n38701), .A3(n37702), .ZN(n37695) );
  NAND3_X2 U14769 ( .A1(n4122), .A2(n10079), .A3(n10081), .ZN(n13779) );
  INV_X1 U14770 ( .A(Ciphertext[17]), .ZN(n8680) );
  INV_X1 U14772 ( .A(n21433), .ZN(n5145) );
  NAND3_X1 U14776 ( .A1(n27145), .A2(n4123), .A3(n27146), .ZN(n24988) );
  NAND3_X1 U14777 ( .A1(n29147), .A2(n626), .A3(n51473), .ZN(n4123) );
  XNOR2_X1 U14778 ( .A(n4124), .B(n48859), .ZN(Plaintext[78]) );
  NOR2_X1 U14779 ( .A1(n4363), .A2(n5407), .ZN(n5406) );
  INV_X1 U14780 ( .A(n12757), .ZN(n11304) );
  NAND2_X1 U14782 ( .A1(n19520), .A2(n598), .ZN(n17036) );
  NAND2_X1 U14783 ( .A1(n18389), .A2(n23217), .ZN(n6576) );
  NAND2_X1 U14784 ( .A1(n14082), .A2(n4125), .ZN(n13333) );
  NAND2_X1 U14785 ( .A1(n14197), .A2(n14200), .ZN(n4125) );
  XNOR2_X1 U14787 ( .A(n18754), .B(n18743), .ZN(n4126) );
  NAND2_X1 U14788 ( .A1(n4129), .A2(n4128), .ZN(n4127) );
  NAND2_X1 U14789 ( .A1(n34924), .A2(n34646), .ZN(n4129) );
  NAND2_X1 U14790 ( .A1(n34647), .A2(n36057), .ZN(n4130) );
  INV_X1 U14791 ( .A(n21564), .ZN(n20782) );
  NAND2_X1 U14792 ( .A1(n23003), .A2(n4132), .ZN(n4131) );
  XNOR2_X2 U14793 ( .A(n4133), .B(n4729), .ZN(n38475) );
  NAND2_X1 U14796 ( .A1(n29094), .A2(n29093), .ZN(n4134) );
  INV_X1 U14797 ( .A(n28023), .ZN(n28021) );
  OAI211_X1 U14798 ( .C1(n7545), .C2(n23351), .A(n6514), .B(n17075), .ZN(n6513) );
  INV_X1 U14799 ( .A(n21154), .ZN(n4849) );
  XNOR2_X1 U14800 ( .A(n34262), .B(n34250), .ZN(n5910) );
  AND3_X1 U14802 ( .A1(n8544), .A2(n33030), .A3(n33041), .ZN(n8113) );
  INV_X1 U14803 ( .A(n47586), .ZN(n8450) );
  INV_X1 U14804 ( .A(n9464), .ZN(n10184) );
  OAI22_X1 U14806 ( .A1(n760), .A2(n20679), .B1(n20678), .B2(n20677), .ZN(
        n20680) );
  NAND2_X1 U14807 ( .A1(n22145), .A2(n22157), .ZN(n19562) );
  NAND2_X1 U14809 ( .A1(n46586), .A2(n2521), .ZN(n44703) );
  NAND4_X4 U14810 ( .A1(n6796), .A2(n6795), .A3(n37197), .A4(n36469), .ZN(
        n39754) );
  NAND3_X1 U14811 ( .A1(n47361), .A2(n49990), .A3(n49989), .ZN(n47351) );
  NAND2_X1 U14814 ( .A1(n21319), .A2(n22586), .ZN(n23441) );
  OR2_X1 U14815 ( .A1(n11346), .A2(n9417), .ZN(n10737) );
  NAND2_X1 U14816 ( .A1(n37200), .A2(n37201), .ZN(n37207) );
  NOR2_X1 U14817 ( .A1(n39015), .A2(n39265), .ZN(n37200) );
  INV_X1 U14818 ( .A(n12893), .ZN(n4383) );
  NAND2_X1 U14819 ( .A1(n37430), .A2(n4137), .ZN(n37431) );
  OR2_X1 U14820 ( .A1(n2192), .A2(n49511), .ZN(n49529) );
  NAND2_X1 U14821 ( .A1(n19826), .A2(n19834), .ZN(n19524) );
  AOI21_X1 U14822 ( .B1(n19841), .B2(n19703), .A(n21185), .ZN(n19526) );
  NAND3_X1 U14823 ( .A1(n7649), .A2(n7648), .A3(n21047), .ZN(n21049) );
  OAI21_X1 U14824 ( .B1(n17853), .B2(n4138), .A(n17852), .ZN(n17854) );
  NAND2_X1 U14825 ( .A1(n19326), .A2(n20360), .ZN(n4138) );
  NAND3_X1 U14826 ( .A1(n46651), .A2(n5360), .A3(n2461), .ZN(n46677) );
  NAND2_X1 U14827 ( .A1(n4742), .A2(n38636), .ZN(n4139) );
  NAND2_X1 U14828 ( .A1(n14345), .A2(n13412), .ZN(n12227) );
  INV_X1 U14829 ( .A(n21707), .ZN(n21708) );
  NAND2_X1 U14830 ( .A1(n22186), .A2(n21712), .ZN(n4140) );
  NOR2_X1 U14831 ( .A1(n4143), .A2(n4142), .ZN(n4141) );
  INV_X1 U14832 ( .A(n30338), .ZN(n29062) );
  NAND2_X1 U14833 ( .A1(n29061), .A2(n28298), .ZN(n30338) );
  NAND2_X2 U14834 ( .A1(n4144), .A2(n17864), .ZN(n22918) );
  NAND2_X1 U14835 ( .A1(n28588), .A2(n51118), .ZN(n28903) );
  NAND3_X1 U14836 ( .A1(n10601), .A2(n10072), .A3(n10604), .ZN(n9909) );
  OAI21_X1 U14837 ( .B1(n22133), .B2(n21847), .A(n23255), .ZN(n21848) );
  NAND3_X2 U14838 ( .A1(n4640), .A2(n19484), .A3(n19485), .ZN(n22593) );
  OR2_X1 U14839 ( .A1(n26668), .A2(n27860), .ZN(n27854) );
  NAND2_X1 U14840 ( .A1(n22919), .A2(n22367), .ZN(n22898) );
  OAI211_X1 U14841 ( .C1(n51796), .C2(n32409), .A(n51640), .B(n33157), .ZN(
        n4145) );
  NAND2_X1 U14842 ( .A1(n4456), .A2(n4147), .ZN(n4146) );
  NAND2_X1 U14844 ( .A1(n31244), .A2(n31781), .ZN(n31229) );
  NAND2_X1 U14845 ( .A1(n33058), .A2(n38562), .ZN(n33059) );
  NAND3_X1 U14846 ( .A1(n19078), .A2(n19076), .A3(n19061), .ZN(n18348) );
  NAND2_X1 U14847 ( .A1(n11470), .A2(n4150), .ZN(n4149) );
  NAND3_X1 U14848 ( .A1(n4151), .A2(n15165), .A3(n51452), .ZN(n14125) );
  NAND2_X1 U14849 ( .A1(n14124), .A2(n7715), .ZN(n4151) );
  NAND4_X1 U14850 ( .A1(n4153), .A2(n47900), .A3(n47945), .A4(n567), .ZN(
        n47901) );
  OAI21_X1 U14851 ( .B1(n47988), .B2(n47937), .A(n51805), .ZN(n4153) );
  XNOR2_X1 U14853 ( .A(n7329), .B(n2329), .ZN(n4154) );
  NAND3_X1 U14854 ( .A1(n8064), .A2(n48128), .A3(n8065), .ZN(n4155) );
  NAND2_X1 U14855 ( .A1(n6091), .A2(n4156), .ZN(n27587) );
  NAND3_X1 U14856 ( .A1(n10863), .A2(n11565), .A3(n51760), .ZN(n10864) );
  NAND2_X1 U14857 ( .A1(n13089), .A2(n13102), .ZN(n11821) );
  XNOR2_X2 U14858 ( .A(n44323), .B(n44322), .ZN(n48479) );
  NOR2_X1 U14859 ( .A1(n24123), .A2(n4726), .ZN(n4725) );
  INV_X1 U14860 ( .A(n39575), .ZN(n41003) );
  AOI22_X1 U14861 ( .A1(n46547), .A2(n48159), .B1(n52344), .B2(n48100), .ZN(
        n48153) );
  NAND2_X1 U14863 ( .A1(n19380), .A2(n4098), .ZN(n20465) );
  NAND2_X1 U14864 ( .A1(n14031), .A2(n4158), .ZN(n14040) );
  NAND2_X1 U14866 ( .A1(n7864), .A2(n4159), .ZN(n7865) );
  NAND3_X1 U14867 ( .A1(n10917), .A2(n10918), .A3(n4160), .ZN(n4159) );
  NAND3_X1 U14868 ( .A1(n8030), .A2(n8031), .A3(n39861), .ZN(n39868) );
  NAND2_X1 U14869 ( .A1(n38078), .A2(n4162), .ZN(n34188) );
  NAND2_X1 U14870 ( .A1(n5541), .A2(n20240), .ZN(n20242) );
  NOR2_X1 U14872 ( .A1(n4163), .A2(n31452), .ZN(n7394) );
  NAND3_X1 U14873 ( .A1(n4164), .A2(n38134), .A3(n38133), .ZN(n38141) );
  NAND2_X1 U14874 ( .A1(n38131), .A2(n38055), .ZN(n4164) );
  NAND3_X1 U14875 ( .A1(n18732), .A2(n18733), .A3(n20692), .ZN(n18735) );
  XNOR2_X2 U14877 ( .A(n8900), .B(Key[44]), .ZN(n11501) );
  NAND2_X1 U14878 ( .A1(n44845), .A2(n2467), .ZN(n46716) );
  NAND2_X1 U14879 ( .A1(n30021), .A2(n2402), .ZN(n30024) );
  NAND2_X1 U14881 ( .A1(n10374), .A2(n4167), .ZN(n4166) );
  INV_X1 U14882 ( .A(n12117), .ZN(n4167) );
  NAND3_X1 U14883 ( .A1(n30067), .A2(n30068), .A3(n2417), .ZN(n30077) );
  NAND2_X1 U14884 ( .A1(n20649), .A2(n20650), .ZN(n21647) );
  NAND2_X1 U14885 ( .A1(n29457), .A2(n27015), .ZN(n26787) );
  NAND3_X2 U14886 ( .A1(n7194), .A2(n10777), .A3(n4168), .ZN(n17829) );
  NAND3_X1 U14887 ( .A1(n10773), .A2(n10774), .A3(n4169), .ZN(n4168) );
  NAND3_X1 U14888 ( .A1(n2500), .A2(n4371), .A3(n19646), .ZN(n19652) );
  XNOR2_X1 U14889 ( .A(n23501), .B(n23500), .ZN(n23524) );
  NAND2_X1 U14890 ( .A1(n49207), .A2(n45967), .ZN(n6502) );
  NAND2_X1 U14891 ( .A1(n4171), .A2(n5270), .ZN(n22552) );
  NAND2_X1 U14892 ( .A1(n22793), .A2(n4549), .ZN(n4171) );
  NAND4_X2 U14893 ( .A1(n44758), .A2(n44759), .A3(n44757), .A4(n44756), .ZN(
        n49126) );
  OR2_X1 U14895 ( .A1(n39166), .A2(n8048), .ZN(n8047) );
  NAND3_X1 U14896 ( .A1(n41641), .A2(n6938), .A3(n41977), .ZN(n41974) );
  NAND2_X1 U14897 ( .A1(n11279), .A2(n11673), .ZN(n7445) );
  NAND2_X1 U14898 ( .A1(n32837), .A2(n4172), .ZN(n32849) );
  NAND2_X1 U14899 ( .A1(n31078), .A2(n32836), .ZN(n4172) );
  NAND2_X1 U14900 ( .A1(n32909), .A2(n4173), .ZN(n28812) );
  NOR2_X1 U14902 ( .A1(n9782), .A2(n4175), .ZN(n10259) );
  OR2_X1 U14903 ( .A1(n36325), .A2(n36338), .ZN(n38144) );
  INV_X1 U14904 ( .A(n19122), .ZN(n19775) );
  NOR2_X1 U14905 ( .A1(n6511), .A2(n13782), .ZN(n6510) );
  XNOR2_X1 U14906 ( .A(n4178), .B(n43644), .ZN(n43646) );
  XNOR2_X1 U14907 ( .A(n43638), .B(n43639), .ZN(n4178) );
  XNOR2_X1 U14908 ( .A(n45159), .B(n43683), .ZN(n44470) );
  NAND2_X1 U14909 ( .A1(n7640), .A2(n49973), .ZN(n49976) );
  NAND3_X2 U14910 ( .A1(n45572), .A2(n4179), .A3(n45573), .ZN(n48112) );
  NAND2_X1 U14911 ( .A1(n39871), .A2(n41695), .ZN(n5960) );
  NAND3_X1 U14912 ( .A1(n9521), .A2(n9522), .A3(n9523), .ZN(n4181) );
  NOR2_X1 U14913 ( .A1(n4183), .A2(n4182), .ZN(n12920) );
  INV_X1 U14914 ( .A(n13095), .ZN(n4183) );
  INV_X1 U14915 ( .A(n27818), .ZN(n29316) );
  XNOR2_X1 U14916 ( .A(n36844), .B(n36843), .ZN(n36846) );
  NAND3_X1 U14918 ( .A1(n39310), .A2(n39311), .A3(n39309), .ZN(n39313) );
  NAND2_X1 U14919 ( .A1(n11400), .A2(n12134), .ZN(n9430) );
  AND2_X1 U14921 ( .A1(n29334), .A2(n29335), .ZN(n6287) );
  INV_X1 U14923 ( .A(n33097), .ZN(n8135) );
  NAND2_X1 U14924 ( .A1(n23092), .A2(n25056), .ZN(n8353) );
  NAND2_X1 U14925 ( .A1(n47137), .A2(n46799), .ZN(n46800) );
  NAND2_X1 U14926 ( .A1(n50853), .A2(n2333), .ZN(n50823) );
  AND3_X1 U14927 ( .A1(n41989), .A2(n41987), .A3(n41988), .ZN(n4187) );
  NAND2_X1 U14929 ( .A1(n32324), .A2(n52182), .ZN(n32326) );
  INV_X1 U14930 ( .A(n12902), .ZN(n12899) );
  OAI211_X1 U14931 ( .C1(n24025), .C2(n24036), .A(n4188), .B(n23393), .ZN(
        n5801) );
  INV_X1 U14932 ( .A(n36680), .ZN(n35268) );
  NOR2_X1 U14933 ( .A1(n4190), .A2(n4189), .ZN(n28018) );
  NAND2_X1 U14934 ( .A1(n28016), .A2(n29018), .ZN(n4189) );
  XNOR2_X2 U14935 ( .A(n17326), .B(n4191), .ZN(n21181) );
  XNOR2_X1 U14936 ( .A(n17157), .B(n17156), .ZN(n4191) );
  NAND2_X1 U14937 ( .A1(n41433), .A2(n40651), .ZN(n40653) );
  NAND2_X1 U14939 ( .A1(n36349), .A2(n36348), .ZN(n4192) );
  NAND2_X1 U14940 ( .A1(n51175), .A2(n14160), .ZN(n12231) );
  NAND2_X1 U14941 ( .A1(n19406), .A2(n2222), .ZN(n4194) );
  NAND3_X1 U14942 ( .A1(n30314), .A2(n30177), .A3(n4197), .ZN(n25200) );
  OR2_X1 U14943 ( .A1(n30181), .A2(n30163), .ZN(n4197) );
  XNOR2_X2 U14946 ( .A(n8771), .B(Key[65]), .ZN(n11011) );
  NAND2_X1 U14947 ( .A1(n11593), .A2(n11604), .ZN(n10806) );
  NAND3_X1 U14949 ( .A1(n5110), .A2(n32214), .A3(n51103), .ZN(n29107) );
  NOR2_X1 U14950 ( .A1(n4201), .A2(n4200), .ZN(n9345) );
  OAI21_X1 U14951 ( .B1(n9344), .B2(n9522), .A(n9342), .ZN(n4200) );
  INV_X1 U14952 ( .A(n9343), .ZN(n4201) );
  NAND2_X1 U14953 ( .A1(n50098), .A2(n4203), .ZN(n4202) );
  NAND4_X1 U14954 ( .A1(n50422), .A2(n50421), .A3(n50423), .A4(n50420), .ZN(
        n4390) );
  NAND2_X1 U14955 ( .A1(n42049), .A2(n42441), .ZN(n42053) );
  NAND2_X1 U14956 ( .A1(n12766), .A2(n13529), .ZN(n7711) );
  NAND2_X1 U14957 ( .A1(n39545), .A2(n39546), .ZN(n4206) );
  NAND3_X1 U14958 ( .A1(n14204), .A2(n14203), .A3(n4207), .ZN(n14206) );
  OAI21_X1 U14959 ( .B1(n11208), .B2(n9352), .A(n9499), .ZN(n8328) );
  XNOR2_X1 U14960 ( .A(n43947), .B(n43948), .ZN(n6918) );
  XOR2_X1 U14961 ( .A(n16575), .B(n5350), .Z(n8465) );
  INV_X1 U14962 ( .A(n47064), .ZN(n8084) );
  INV_X1 U14963 ( .A(n22585), .ZN(n22584) );
  OAI21_X1 U14964 ( .B1(n21777), .B2(n21117), .A(n21115), .ZN(n5446) );
  NAND4_X1 U14965 ( .A1(n26727), .A2(n27839), .A3(n26646), .A4(n29450), .ZN(
        n26647) );
  INV_X1 U14968 ( .A(n6461), .ZN(n31817) );
  XNOR2_X2 U14969 ( .A(n8557), .B(n15742), .ZN(n21664) );
  NAND2_X1 U14970 ( .A1(n17603), .A2(n17504), .ZN(n18322) );
  XNOR2_X2 U14972 ( .A(Key[180]), .B(n8878), .ZN(n12728) );
  NAND2_X1 U14973 ( .A1(n11964), .A2(n12720), .ZN(n9573) );
  INV_X1 U14974 ( .A(n19504), .ZN(n5177) );
  AND2_X1 U14975 ( .A1(n40774), .A2(n426), .ZN(n40596) );
  AND4_X1 U14976 ( .A1(n46526), .A2(n46525), .A3(n7062), .A4(n7063), .ZN(n7061) );
  NAND2_X1 U14977 ( .A1(n12314), .A2(n10296), .ZN(n12299) );
  NAND3_X1 U14978 ( .A1(n9026), .A2(n10245), .A3(n10195), .ZN(n9027) );
  NAND2_X1 U14979 ( .A1(n10245), .A2(n8781), .ZN(n9026) );
  AND3_X1 U14980 ( .A1(n50256), .A2(n50258), .A3(n50257), .ZN(n50274) );
  XNOR2_X1 U14981 ( .A(n44208), .B(n44911), .ZN(n45263) );
  INV_X1 U14982 ( .A(n7107), .ZN(n7106) );
  OR2_X1 U14983 ( .A1(n32389), .A2(n32843), .ZN(n32848) );
  INV_X1 U14984 ( .A(n22874), .ZN(n23105) );
  INV_X1 U14985 ( .A(n6921), .ZN(n33617) );
  INV_X1 U14986 ( .A(n45515), .ZN(n4214) );
  INV_X1 U14987 ( .A(n45514), .ZN(n4215) );
  NAND2_X1 U14989 ( .A1(n30390), .A2(n30394), .ZN(n4217) );
  INV_X1 U14990 ( .A(n41029), .ZN(n40420) );
  XNOR2_X1 U14991 ( .A(n18407), .B(n14427), .ZN(n16953) );
  INV_X1 U14992 ( .A(n18669), .ZN(n19203) );
  INV_X1 U14993 ( .A(n50343), .ZN(n50335) );
  NAND3_X1 U14994 ( .A1(n7258), .A2(n19892), .A3(n19887), .ZN(n7261) );
  INV_X1 U14995 ( .A(n29794), .ZN(n29802) );
  INV_X1 U14997 ( .A(n14137), .ZN(n13069) );
  OAI21_X1 U14998 ( .B1(n5400), .B2(n5399), .A(n51022), .ZN(n5398) );
  NOR2_X1 U14999 ( .A1(n13129), .A2(n7853), .ZN(n7852) );
  INV_X1 U15000 ( .A(n38135), .ZN(n5464) );
  AOI21_X1 U15001 ( .B1(n13122), .B2(n14159), .A(n14966), .ZN(n13116) );
  NOR2_X1 U15002 ( .A1(n38073), .A2(n2331), .ZN(n36634) );
  XNOR2_X1 U15003 ( .A(n45421), .B(n46059), .ZN(n45428) );
  XNOR2_X1 U15004 ( .A(n4218), .B(n18803), .ZN(n18808) );
  XNOR2_X1 U15005 ( .A(n18800), .B(n18799), .ZN(n4218) );
  NAND2_X1 U15007 ( .A1(n19427), .A2(n4219), .ZN(n15461) );
  NAND3_X1 U15008 ( .A1(n23984), .A2(n22427), .A3(n23981), .ZN(n24006) );
  NAND2_X1 U15009 ( .A1(n12538), .A2(n6409), .ZN(n10787) );
  INV_X1 U15010 ( .A(n21767), .ZN(n6167) );
  NAND2_X1 U15012 ( .A1(n38050), .A2(n36167), .ZN(n36329) );
  NAND2_X1 U15014 ( .A1(n38611), .A2(n40380), .ZN(n41142) );
  INV_X1 U15015 ( .A(n11954), .ZN(n6912) );
  NAND2_X1 U15016 ( .A1(n12435), .A2(n12440), .ZN(n11937) );
  NAND2_X1 U15017 ( .A1(n5299), .A2(n12709), .ZN(n4221) );
  OAI21_X1 U15018 ( .B1(n29063), .B2(n29768), .A(n4222), .ZN(n29059) );
  NAND2_X1 U15019 ( .A1(n29063), .A2(n28300), .ZN(n4222) );
  XNOR2_X1 U15020 ( .A(n34491), .B(n35503), .ZN(n4224) );
  NAND3_X2 U15021 ( .A1(n45798), .A2(n4226), .A3(n4227), .ZN(n47686) );
  NAND2_X1 U15022 ( .A1(n45789), .A2(n45790), .ZN(n4226) );
  INV_X1 U15023 ( .A(n7985), .ZN(n41394) );
  NAND2_X1 U15024 ( .A1(n19348), .A2(n20515), .ZN(n6282) );
  OR2_X1 U15025 ( .A1(n41539), .A2(n40943), .ZN(n41390) );
  NAND2_X1 U15027 ( .A1(n4228), .A2(n32478), .ZN(n31210) );
  NAND2_X1 U15028 ( .A1(n709), .A2(n29625), .ZN(n29627) );
  NAND2_X1 U15029 ( .A1(n24411), .A2(n24412), .ZN(n24074) );
  AND4_X2 U15031 ( .A1(n46377), .A2(n46379), .A3(n46378), .A4(n48556), .ZN(
        n48769) );
  NAND2_X1 U15032 ( .A1(n9586), .A2(n6147), .ZN(n4229) );
  INV_X1 U15033 ( .A(n21674), .ZN(n24072) );
  INV_X1 U15034 ( .A(n10733), .ZN(n14172) );
  NAND2_X1 U15035 ( .A1(n9636), .A2(n6677), .ZN(n6676) );
  OAI211_X1 U15036 ( .C1(n48394), .C2(n48360), .A(n48299), .B(n48347), .ZN(
        n48300) );
  NAND3_X1 U15037 ( .A1(n6986), .A2(n52172), .A3(n48381), .ZN(n48394) );
  XNOR2_X2 U15038 ( .A(n8801), .B(Key[84]), .ZN(n10968) );
  NAND3_X1 U15039 ( .A1(n8040), .A2(n27517), .A3(n29698), .ZN(n27518) );
  NAND2_X1 U15040 ( .A1(n11660), .A2(n9515), .ZN(n10565) );
  NAND2_X1 U15041 ( .A1(n11639), .A2(n9306), .ZN(n9515) );
  OAI21_X1 U15042 ( .B1(n11751), .B2(n786), .A(n4232), .ZN(n4960) );
  NAND2_X1 U15043 ( .A1(n11209), .A2(n51650), .ZN(n9927) );
  INV_X1 U15044 ( .A(Ciphertext[66]), .ZN(n8913) );
  NAND4_X4 U15045 ( .A1(n39025), .A2(n39022), .A3(n39024), .A4(n39023), .ZN(
        n41706) );
  XNOR2_X1 U15046 ( .A(n4233), .B(n18767), .ZN(n18772) );
  XNOR2_X1 U15047 ( .A(n18768), .B(n18766), .ZN(n4233) );
  NAND2_X1 U15048 ( .A1(n39285), .A2(n39271), .ZN(n8461) );
  AOI21_X1 U15049 ( .B1(n8194), .B2(n41707), .A(n41174), .ZN(n8196) );
  NAND3_X1 U15050 ( .A1(n27621), .A2(n27728), .A3(n26890), .ZN(n27723) );
  NAND2_X1 U15052 ( .A1(n26468), .A2(n30312), .ZN(n26466) );
  NAND2_X1 U15054 ( .A1(n32507), .A2(n30873), .ZN(n30877) );
  XNOR2_X2 U15055 ( .A(Key[164]), .B(Ciphertext[121]), .ZN(n10101) );
  NAND2_X1 U15056 ( .A1(n42205), .A2(n42209), .ZN(n4862) );
  INV_X1 U15057 ( .A(n11393), .ZN(n6465) );
  NAND2_X1 U15058 ( .A1(n38708), .A2(n4238), .ZN(n38710) );
  NAND2_X1 U15059 ( .A1(n39246), .A2(n39236), .ZN(n38708) );
  XNOR2_X1 U15060 ( .A(n20887), .B(n25338), .ZN(n4239) );
  NAND2_X1 U15061 ( .A1(n45550), .A2(n45549), .ZN(n5437) );
  NAND2_X1 U15062 ( .A1(n29270), .A2(n29272), .ZN(n27782) );
  NOR2_X1 U15063 ( .A1(n19865), .A2(n19650), .ZN(n4242) );
  NAND3_X1 U15064 ( .A1(n45851), .A2(n45850), .A3(n2497), .ZN(n45852) );
  INV_X1 U15065 ( .A(n14159), .ZN(n13124) );
  NAND2_X1 U15066 ( .A1(n48535), .A2(n48527), .ZN(n6097) );
  NAND4_X2 U15068 ( .A1(n15209), .A2(n15211), .A3(n15210), .A4(n15208), .ZN(
        n18427) );
  INV_X1 U15069 ( .A(n10262), .ZN(n12356) );
  NAND4_X2 U15070 ( .A1(n22193), .A2(n22194), .A3(n22192), .A4(n22195), .ZN(
        n25481) );
  NAND2_X1 U15071 ( .A1(n31326), .A2(n32352), .ZN(n4245) );
  INV_X1 U15072 ( .A(n44841), .ZN(n6101) );
  AND2_X1 U15074 ( .A1(n47581), .A2(n47567), .ZN(n4581) );
  INV_X1 U15075 ( .A(n46686), .ZN(n46904) );
  NAND2_X1 U15076 ( .A1(n26676), .A2(n26671), .ZN(n8744) );
  INV_X1 U15078 ( .A(n6048), .ZN(n30756) );
  AND3_X1 U15080 ( .A1(n45373), .A2(n45371), .A3(n48554), .ZN(n7376) );
  XNOR2_X1 U15081 ( .A(n37066), .B(n36847), .ZN(n35509) );
  AND2_X1 U15082 ( .A1(n29928), .A2(n30777), .ZN(n8507) );
  NOR2_X1 U15083 ( .A1(n680), .A2(n40250), .ZN(n41933) );
  INV_X1 U15084 ( .A(n38876), .ZN(n41088) );
  INV_X1 U15085 ( .A(n46609), .ZN(n46921) );
  INV_X1 U15086 ( .A(n15414), .ZN(n5715) );
  INV_X1 U15087 ( .A(n20611), .ZN(n21514) );
  XNOR2_X1 U15088 ( .A(n5611), .B(n17381), .ZN(n16653) );
  OAI21_X1 U15089 ( .B1(n39937), .B2(n2386), .A(n4251), .ZN(n38836) );
  NAND2_X1 U15091 ( .A1(n12954), .A2(n12953), .ZN(n4252) );
  NAND2_X1 U15092 ( .A1(n4253), .A2(n38330), .ZN(n6796) );
  INV_X1 U15093 ( .A(n39112), .ZN(n38827) );
  NAND2_X1 U15094 ( .A1(n39754), .A2(n39752), .ZN(n39112) );
  XNOR2_X2 U15095 ( .A(n13056), .B(n13055), .ZN(n17484) );
  NAND4_X2 U15096 ( .A1(n6898), .A2(n17515), .A3(n4254), .A4(n6896), .ZN(
        n24344) );
  NAND2_X1 U15098 ( .A1(n12750), .A2(n14643), .ZN(n13659) );
  OAI21_X1 U15099 ( .B1(n33018), .B2(n33019), .A(n8516), .ZN(n33020) );
  XNOR2_X1 U15100 ( .A(n24871), .B(n7613), .ZN(n7612) );
  OAI21_X1 U15101 ( .B1(n51686), .B2(n15263), .A(n4611), .ZN(n14782) );
  NAND2_X1 U15102 ( .A1(n4256), .A2(n4255), .ZN(n22346) );
  NAND2_X1 U15103 ( .A1(n27618), .A2(n27732), .ZN(n4255) );
  NAND2_X1 U15104 ( .A1(n26891), .A2(n737), .ZN(n4256) );
  NAND2_X1 U15105 ( .A1(n23446), .A2(n23445), .ZN(n19554) );
  NAND2_X1 U15110 ( .A1(n47477), .A2(n48957), .ZN(n48930) );
  XNOR2_X1 U15111 ( .A(n35775), .B(n4260), .ZN(n5531) );
  NAND4_X1 U15113 ( .A1(n32067), .A2(n32068), .A3(n32074), .A4(n7430), .ZN(
        n4261) );
  INV_X1 U15114 ( .A(n18969), .ZN(n19098) );
  INV_X1 U15115 ( .A(n9405), .ZN(n10375) );
  INV_X1 U15116 ( .A(n32608), .ZN(n7625) );
  OAI21_X1 U15117 ( .B1(n14170), .B2(n14595), .A(n4262), .ZN(n10765) );
  XNOR2_X1 U15118 ( .A(n15877), .B(n356), .ZN(n4762) );
  XNOR2_X1 U15119 ( .A(n17250), .B(n17251), .ZN(n4263) );
  NAND2_X1 U15120 ( .A1(n29790), .A2(n3826), .ZN(n4265) );
  NAND2_X1 U15121 ( .A1(n28950), .A2(n28862), .ZN(n28953) );
  NAND2_X1 U15122 ( .A1(n39072), .A2(n39073), .ZN(n39089) );
  NAND3_X1 U15124 ( .A1(n31394), .A2(n32823), .A3(n31404), .ZN(n31252) );
  NAND2_X1 U15125 ( .A1(n37941), .A2(n38689), .ZN(n36774) );
  NAND2_X1 U15126 ( .A1(n4711), .A2(n4266), .ZN(n31524) );
  NAND2_X2 U15127 ( .A1(n5137), .A2(n4268), .ZN(n18407) );
  AND3_X1 U15128 ( .A1(n13073), .A2(n4269), .A3(n13074), .ZN(n4268) );
  AOI21_X1 U15129 ( .B1(n13068), .B2(n14795), .A(n13067), .ZN(n4269) );
  NAND2_X1 U15130 ( .A1(n37663), .A2(n4270), .ZN(n37666) );
  OR2_X1 U15131 ( .A1(n35162), .A2(n38037), .ZN(n38033) );
  INV_X1 U15132 ( .A(n49932), .ZN(n49892) );
  AND2_X2 U15133 ( .A1(n37809), .A2(n2176), .ZN(n39481) );
  NAND4_X2 U15134 ( .A1(n38048), .A2(n38046), .A3(n38047), .A4(n38045), .ZN(
        n40269) );
  XNOR2_X1 U15135 ( .A(n42699), .B(n42698), .ZN(n43432) );
  XNOR2_X1 U15136 ( .A(n4271), .B(n27396), .ZN(n27397) );
  XNOR2_X1 U15137 ( .A(n27394), .B(n27395), .ZN(n4271) );
  NAND2_X1 U15138 ( .A1(n28764), .A2(n30376), .ZN(n29774) );
  INV_X1 U15140 ( .A(n17521), .ZN(n17534) );
  NAND2_X1 U15141 ( .A1(n20013), .A2(n17522), .ZN(n17521) );
  INV_X1 U15142 ( .A(n38723), .ZN(n37182) );
  AND2_X1 U15143 ( .A1(n38723), .A2(n37183), .ZN(n39311) );
  NAND2_X1 U15144 ( .A1(n39289), .A2(n39290), .ZN(n38723) );
  XNOR2_X1 U15146 ( .A(n4272), .B(n28119), .ZN(n24632) );
  XNOR2_X1 U15147 ( .A(n24630), .B(n25385), .ZN(n4272) );
  NAND2_X1 U15148 ( .A1(n6107), .A2(n30846), .ZN(n6461) );
  NAND2_X1 U15149 ( .A1(n5947), .A2(n5946), .ZN(n4273) );
  INV_X1 U15150 ( .A(n46636), .ZN(n4274) );
  XNOR2_X1 U15152 ( .A(n37001), .B(n36873), .ZN(n36875) );
  INV_X1 U15153 ( .A(n9918), .ZN(n8528) );
  INV_X1 U15154 ( .A(n27715), .ZN(n27714) );
  XNOR2_X1 U15155 ( .A(n4276), .B(n34304), .ZN(n34308) );
  XNOR2_X1 U15156 ( .A(n34622), .B(n8037), .ZN(n4276) );
  NAND2_X1 U15159 ( .A1(n51761), .A2(n10556), .ZN(n10547) );
  NAND2_X1 U15160 ( .A1(n11670), .A2(n11673), .ZN(n11278) );
  AND3_X1 U15163 ( .A1(n31226), .A2(n7252), .A3(n7250), .ZN(n7251) );
  INV_X1 U15164 ( .A(n13087), .ZN(n13081) );
  NAND2_X1 U15165 ( .A1(n36125), .A2(n38155), .ZN(n36130) );
  INV_X1 U15166 ( .A(n22390), .ZN(n5370) );
  NAND2_X1 U15167 ( .A1(n14700), .A2(n13335), .ZN(n13342) );
  XNOR2_X1 U15168 ( .A(n4281), .B(n44551), .ZN(n44552) );
  XNOR2_X1 U15169 ( .A(n44927), .B(n44550), .ZN(n4281) );
  NAND3_X1 U15170 ( .A1(n693), .A2(n36132), .A3(n38589), .ZN(n7954) );
  OR2_X1 U15171 ( .A1(n47105), .A2(n47089), .ZN(n6586) );
  NAND2_X1 U15172 ( .A1(n6049), .A2(n803), .ZN(n10045) );
  AND2_X1 U15173 ( .A1(n12268), .A2(n12257), .ZN(n12252) );
  NAND2_X1 U15174 ( .A1(n9985), .A2(n9986), .ZN(n9987) );
  NAND2_X1 U15175 ( .A1(n51669), .A2(n14709), .ZN(n14197) );
  AND3_X1 U15176 ( .A1(n11839), .A2(n11833), .A3(n11838), .ZN(n5551) );
  NAND2_X1 U15177 ( .A1(n14123), .A2(n15161), .ZN(n14577) );
  NAND2_X1 U15178 ( .A1(n49639), .A2(n50294), .ZN(n46035) );
  NAND2_X1 U15179 ( .A1(n49946), .A2(n51313), .ZN(n49639) );
  INV_X1 U15180 ( .A(n20211), .ZN(n19678) );
  OR2_X1 U15181 ( .A1(n7117), .A2(n52101), .ZN(n39643) );
  INV_X1 U15182 ( .A(n26436), .ZN(n27258) );
  OR2_X1 U15183 ( .A1(n41685), .A2(n41670), .ZN(n7034) );
  OR2_X1 U15188 ( .A1(n41202), .A2(n51430), .ZN(n4284) );
  NAND2_X1 U15189 ( .A1(n12068), .A2(n12066), .ZN(n12627) );
  INV_X1 U15190 ( .A(n49993), .ZN(n50009) );
  INV_X1 U15192 ( .A(n46869), .ZN(n44578) );
  INV_X1 U15193 ( .A(n51250), .ZN(n23150) );
  NOR2_X1 U15194 ( .A1(n33786), .A2(n33785), .ZN(n4734) );
  NAND2_X1 U15195 ( .A1(n354), .A2(n24030), .ZN(n22100) );
  INV_X1 U15196 ( .A(n32633), .ZN(n32908) );
  NOR2_X2 U15197 ( .A1(n13718), .A2(n13717), .ZN(n18756) );
  OAI21_X1 U15199 ( .B1(n22274), .B2(n23352), .A(n22276), .ZN(n23355) );
  INV_X1 U15200 ( .A(n22379), .ZN(n23813) );
  INV_X1 U15201 ( .A(n10047), .ZN(n9858) );
  INV_X1 U15202 ( .A(n18823), .ZN(n7045) );
  INV_X1 U15203 ( .A(n30459), .ZN(n28523) );
  INV_X1 U15204 ( .A(n41195), .ZN(n39502) );
  INV_X1 U15205 ( .A(Ciphertext[68]), .ZN(n8638) );
  INV_X1 U15206 ( .A(n10601), .ZN(n10606) );
  INV_X1 U15207 ( .A(n21945), .ZN(n6875) );
  INV_X1 U15208 ( .A(n28923), .ZN(n7226) );
  OR2_X1 U15209 ( .A1(n28915), .A2(n7226), .ZN(n29012) );
  OAI21_X1 U15210 ( .B1(n29931), .B2(n30688), .A(n30699), .ZN(n24093) );
  INV_X1 U15211 ( .A(n51677), .ZN(n8224) );
  NAND4_X2 U15212 ( .A1(n8928), .A2(n8927), .A3(n8929), .A4(n8926), .ZN(n14983) );
  AND3_X1 U15213 ( .A1(n46548), .A2(n46550), .A3(n46549), .ZN(n4288) );
  INV_X1 U15214 ( .A(n28547), .ZN(n28550) );
  NAND2_X1 U15215 ( .A1(n30285), .A2(n30280), .ZN(n28547) );
  INV_X1 U15216 ( .A(n381), .ZN(n31455) );
  NAND2_X1 U15217 ( .A1(n31160), .A2(n4289), .ZN(n31162) );
  OR2_X1 U15218 ( .A1(n39259), .A2(n551), .ZN(n38686) );
  INV_X1 U15219 ( .A(n21567), .ZN(n21557) );
  NAND3_X1 U15220 ( .A1(n2527), .A2(n5069), .A3(n23638), .ZN(n22628) );
  NAND4_X2 U15221 ( .A1(n19571), .A2(n19570), .A3(n19569), .A4(n19572), .ZN(
        n28103) );
  XOR2_X1 U15222 ( .A(n34770), .B(n32040), .Z(n8609) );
  XNOR2_X1 U15223 ( .A(n4291), .B(n45277), .ZN(n41366) );
  XNOR2_X1 U15224 ( .A(n41310), .B(n41309), .ZN(n4291) );
  NAND3_X1 U15225 ( .A1(n13446), .A2(n13447), .A3(n13445), .ZN(n13453) );
  XNOR2_X1 U15226 ( .A(n18768), .B(n17886), .ZN(n4292) );
  INV_X1 U15227 ( .A(n45657), .ZN(n5690) );
  INV_X1 U15228 ( .A(n32014), .ZN(n32481) );
  XNOR2_X1 U15230 ( .A(n17179), .B(n51014), .ZN(n17188) );
  XNOR2_X1 U15231 ( .A(n25681), .B(n20572), .ZN(n4293) );
  NOR2_X1 U15233 ( .A1(n7002), .A2(n4294), .ZN(n6997) );
  NOR2_X1 U15234 ( .A1(n39613), .A2(n6999), .ZN(n4294) );
  INV_X1 U15235 ( .A(n8968), .ZN(n8469) );
  NAND2_X1 U15236 ( .A1(n35015), .A2(n611), .ZN(n38052) );
  NAND2_X1 U15237 ( .A1(n38068), .A2(n38138), .ZN(n4297) );
  INV_X1 U15238 ( .A(n32412), .ZN(n32411) );
  INV_X1 U15239 ( .A(n48267), .ZN(n5561) );
  NOR2_X1 U15240 ( .A1(n48887), .A2(n48888), .ZN(n5709) );
  NAND3_X1 U15241 ( .A1(n37485), .A2(n37432), .A3(n37490), .ZN(n37434) );
  NAND2_X1 U15242 ( .A1(n23674), .A2(n23667), .ZN(n22098) );
  NOR2_X1 U15244 ( .A1(n13646), .A2(n13667), .ZN(n8127) );
  INV_X1 U15245 ( .A(n31099), .ZN(n30916) );
  INV_X1 U15246 ( .A(n19132), .ZN(n19488) );
  INV_X1 U15247 ( .A(n711), .ZN(n4299) );
  NAND2_X1 U15248 ( .A1(n435), .A2(n386), .ZN(n31366) );
  NAND3_X1 U15250 ( .A1(n15260), .A2(n51685), .A3(n15263), .ZN(n15261) );
  NAND2_X1 U15251 ( .A1(n20063), .A2(n16217), .ZN(n19131) );
  NAND2_X1 U15252 ( .A1(n36558), .A2(n4300), .ZN(n36480) );
  XNOR2_X1 U15253 ( .A(n4301), .B(n48815), .ZN(Plaintext[76]) );
  INV_X1 U15254 ( .A(n22018), .ZN(n22590) );
  AND2_X1 U15255 ( .A1(n19486), .A2(n19483), .ZN(n4640) );
  NAND4_X1 U15256 ( .A1(n4303), .A2(n50711), .A3(n50713), .A4(n50712), .ZN(
        n50715) );
  NAND2_X1 U15257 ( .A1(n47307), .A2(n49639), .ZN(n50309) );
  NAND3_X1 U15258 ( .A1(n9114), .A2(n11449), .A3(n9113), .ZN(n9115) );
  XNOR2_X1 U15259 ( .A(n4304), .B(n26171), .ZN(n26020) );
  XNOR2_X1 U15260 ( .A(n6308), .B(n26018), .ZN(n4304) );
  INV_X1 U15261 ( .A(n4305), .ZN(n8105) );
  OAI211_X1 U15262 ( .C1(n12759), .C2(n13658), .A(n12758), .B(n13654), .ZN(
        n4305) );
  NAND2_X1 U15263 ( .A1(n46574), .A2(n46705), .ZN(n44840) );
  NAND2_X1 U15264 ( .A1(n11461), .A2(n11467), .ZN(n11625) );
  NAND2_X1 U15266 ( .A1(n19639), .A2(n585), .ZN(n19032) );
  NOR2_X1 U15267 ( .A1(n30737), .A2(n4306), .ZN(n30380) );
  NAND2_X1 U15268 ( .A1(n1121), .A2(n29883), .ZN(n4306) );
  NAND2_X1 U15269 ( .A1(n4310), .A2(n14341), .ZN(n4309) );
  NAND3_X1 U15270 ( .A1(n39016), .A2(n39285), .A3(n39269), .ZN(n39017) );
  NAND2_X1 U15271 ( .A1(n13526), .A2(n51066), .ZN(n13530) );
  NAND4_X1 U15273 ( .A1(n11130), .A2(n9263), .A3(n11919), .A4(n9264), .ZN(
        n4313) );
  INV_X1 U15274 ( .A(n21768), .ZN(n21765) );
  INV_X1 U15275 ( .A(n21114), .ZN(n4314) );
  NAND2_X1 U15276 ( .A1(n22291), .A2(n21122), .ZN(n4315) );
  INV_X1 U15277 ( .A(n5734), .ZN(n5733) );
  INV_X1 U15278 ( .A(n9679), .ZN(n8643) );
  INV_X1 U15279 ( .A(n22533), .ZN(n5118) );
  INV_X1 U15280 ( .A(n20483), .ZN(n17636) );
  NAND3_X1 U15282 ( .A1(n11714), .A2(n11707), .A3(n11203), .ZN(n9502) );
  NAND2_X1 U15284 ( .A1(n32200), .A2(n32199), .ZN(n4319) );
  INV_X1 U15286 ( .A(n11344), .ZN(n11348) );
  NAND2_X1 U15287 ( .A1(n12258), .A2(n12257), .ZN(n11344) );
  NAND2_X1 U15288 ( .A1(n4407), .A2(n22879), .ZN(n22882) );
  NOR2_X1 U15289 ( .A1(n40663), .A2(n40664), .ZN(n5064) );
  NAND2_X1 U15290 ( .A1(n27400), .A2(n4320), .ZN(n28771) );
  NAND2_X1 U15291 ( .A1(n52042), .A2(n48567), .ZN(n48583) );
  NAND2_X1 U15292 ( .A1(n48640), .A2(n48604), .ZN(n4321) );
  OAI21_X1 U15293 ( .B1(n32714), .B2(n32715), .A(n32716), .ZN(n32736) );
  NAND4_X2 U15294 ( .A1(n4323), .A2(n4322), .A3(n21696), .A4(n21697), .ZN(
        n27291) );
  NAND2_X1 U15295 ( .A1(n21691), .A2(n21690), .ZN(n4322) );
  AOI21_X1 U15296 ( .B1(n36097), .B2(n38573), .A(n6024), .ZN(n36111) );
  XOR2_X1 U15297 ( .A(n33354), .B(n33864), .Z(n6143) );
  INV_X1 U15298 ( .A(n14952), .ZN(n14060) );
  XNOR2_X1 U15299 ( .A(n19232), .B(n19231), .ZN(n19969) );
  NAND2_X1 U15300 ( .A1(n22831), .A2(n22491), .ZN(n21074) );
  OAI21_X1 U15301 ( .B1(n11539), .B2(n51653), .A(n12516), .ZN(n12517) );
  NAND2_X1 U15302 ( .A1(n5370), .A2(n22375), .ZN(n22740) );
  INV_X1 U15304 ( .A(n13669), .ZN(n8121) );
  NAND2_X1 U15305 ( .A1(n7264), .A2(n12545), .ZN(n9117) );
  NAND3_X1 U15306 ( .A1(n32246), .A2(n32244), .A3(n32239), .ZN(n29373) );
  NAND3_X1 U15307 ( .A1(n28663), .A2(n28664), .A3(n30228), .ZN(n25853) );
  NAND3_X2 U15308 ( .A1(n4327), .A2(n34991), .A3(n2389), .ZN(n41063) );
  NAND2_X1 U15309 ( .A1(n34986), .A2(n36535), .ZN(n4327) );
  INV_X1 U15310 ( .A(n23196), .ZN(n22609) );
  OAI21_X1 U15312 ( .B1(n39427), .B2(n39205), .A(n38941), .ZN(n37905) );
  INV_X1 U15313 ( .A(Ciphertext[124]), .ZN(n8626) );
  AND3_X1 U15314 ( .A1(n28518), .A2(n28832), .A3(n28519), .ZN(n6716) );
  INV_X1 U15315 ( .A(n37881), .ZN(n38962) );
  INV_X1 U15316 ( .A(n14945), .ZN(n14935) );
  XNOR2_X1 U15318 ( .A(n42938), .B(n6327), .ZN(n42636) );
  NAND4_X2 U15319 ( .A1(n38824), .A2(n4738), .A3(n38823), .A4(n38822), .ZN(
        n44189) );
  XNOR2_X1 U15320 ( .A(n4330), .B(n23779), .ZN(n23780) );
  XNOR2_X1 U15321 ( .A(n23778), .B(n23777), .ZN(n4330) );
  NAND2_X1 U15322 ( .A1(n21085), .A2(n24290), .ZN(n24280) );
  INV_X1 U15323 ( .A(n49149), .ZN(n49141) );
  NAND2_X1 U15324 ( .A1(n43421), .A2(n49146), .ZN(n49149) );
  XNOR2_X1 U15325 ( .A(n4331), .B(n49293), .ZN(Plaintext[102]) );
  NAND3_X1 U15326 ( .A1(n49292), .A2(n49290), .A3(n2404), .ZN(n4331) );
  INV_X1 U15327 ( .A(n40468), .ZN(n40469) );
  OAI21_X1 U15328 ( .B1(n4335), .B2(n49145), .A(n7657), .ZN(n49156) );
  NAND2_X1 U15329 ( .A1(n49144), .A2(n49143), .ZN(n4335) );
  XNOR2_X1 U15332 ( .A(n4336), .B(n34769), .ZN(n34772) );
  XNOR2_X1 U15333 ( .A(n34768), .B(n34770), .ZN(n4336) );
  XNOR2_X1 U15334 ( .A(n19194), .B(n2515), .ZN(n5667) );
  OAI21_X1 U15335 ( .B1(n49282), .B2(n49367), .A(n49380), .ZN(n49283) );
  NAND3_X1 U15336 ( .A1(n12495), .A2(n10832), .A3(n642), .ZN(n8927) );
  INV_X1 U15337 ( .A(n38726), .ZN(n4337) );
  NAND3_X1 U15338 ( .A1(n10782), .A2(n11446), .A3(n9118), .ZN(n8937) );
  NAND3_X1 U15339 ( .A1(n17875), .A2(n17874), .A3(n4339), .ZN(n17876) );
  NAND2_X1 U15340 ( .A1(n19412), .A2(n4340), .ZN(n4339) );
  INV_X1 U15342 ( .A(n19577), .ZN(n22904) );
  NAND2_X1 U15343 ( .A1(n37488), .A2(n36161), .ZN(n38529) );
  NAND2_X1 U15344 ( .A1(n1206), .A2(n13885), .ZN(n15417) );
  NAND2_X1 U15345 ( .A1(n33034), .A2(n32874), .ZN(n32870) );
  NAND2_X1 U15347 ( .A1(n40372), .A2(n41332), .ZN(n4341) );
  NAND2_X1 U15348 ( .A1(n39823), .A2(n39822), .ZN(n4342) );
  NAND3_X2 U15351 ( .A1(n6909), .A2(n6908), .A3(n9583), .ZN(n13061) );
  NAND3_X1 U15352 ( .A1(n8592), .A2(n20475), .A3(n20476), .ZN(n8591) );
  OAI21_X1 U15353 ( .B1(n9206), .B2(n7150), .A(n10463), .ZN(n6036) );
  XNOR2_X1 U15354 ( .A(n32656), .B(n35768), .ZN(n33686) );
  NAND4_X2 U15355 ( .A1(n30336), .A2(n30334), .A3(n30333), .A4(n30335), .ZN(
        n34760) );
  NAND2_X1 U15356 ( .A1(n41674), .A2(n41227), .ZN(n41247) );
  NAND2_X1 U15358 ( .A1(n17621), .A2(n4347), .ZN(n4346) );
  XNOR2_X2 U15359 ( .A(n44525), .B(n42576), .ZN(n44320) );
  OAI22_X1 U15361 ( .A1(n45593), .A2(n45594), .B1(n45592), .B2(n48436), .ZN(
        n4348) );
  NAND2_X1 U15362 ( .A1(n646), .A2(n48135), .ZN(n46538) );
  NAND2_X1 U15363 ( .A1(n6860), .A2(n39100), .ZN(n35434) );
  NAND3_X2 U15364 ( .A1(n7983), .A2(n4350), .A3(n7982), .ZN(n17901) );
  XNOR2_X1 U15365 ( .A(n18148), .B(n18149), .ZN(n18151) );
  XNOR2_X2 U15366 ( .A(n18519), .B(n18755), .ZN(n18148) );
  NAND2_X1 U15367 ( .A1(n29123), .A2(n29260), .ZN(n29249) );
  XNOR2_X2 U15369 ( .A(n9042), .B(Key[102]), .ZN(n12340) );
  INV_X1 U15371 ( .A(Ciphertext[151]), .ZN(n7751) );
  OAI21_X1 U15372 ( .B1(n5260), .B2(n23705), .A(n23704), .ZN(n5259) );
  XNOR2_X1 U15373 ( .A(n43240), .B(n2228), .ZN(n43241) );
  OR2_X2 U15374 ( .A1(n32117), .A2(n32116), .ZN(n34869) );
  INV_X1 U15375 ( .A(n21680), .ZN(n25729) );
  NAND2_X1 U15376 ( .A1(n30171), .A2(n30163), .ZN(n30312) );
  XNOR2_X2 U15377 ( .A(n7664), .B(n7663), .ZN(n30163) );
  NAND3_X1 U15378 ( .A1(n4354), .A2(n29882), .A3(n1121), .ZN(n5843) );
  NAND2_X1 U15379 ( .A1(n30377), .A2(n30378), .ZN(n4354) );
  NAND2_X1 U15380 ( .A1(n23099), .A2(n22890), .ZN(n19883) );
  INV_X1 U15382 ( .A(n32429), .ZN(n31397) );
  NAND2_X1 U15383 ( .A1(n34912), .A2(n37500), .ZN(n36240) );
  NAND2_X1 U15385 ( .A1(n4357), .A2(n26468), .ZN(n26470) );
  OAI22_X1 U15386 ( .A1(n26467), .A2(n6084), .B1(n29140), .B2(n30306), .ZN(
        n4357) );
  NAND2_X1 U15387 ( .A1(n12549), .A2(n12547), .ZN(n11449) );
  INV_X1 U15388 ( .A(n30767), .ZN(n24350) );
  AOI22_X1 U15389 ( .A1(n4358), .A2(n14442), .B1(n9), .B2(n11811), .ZN(n11438)
         );
  NAND2_X1 U15391 ( .A1(n27855), .A2(n2956), .ZN(n4359) );
  NAND2_X1 U15392 ( .A1(n4362), .A2(n4361), .ZN(n4360) );
  NAND2_X1 U15393 ( .A1(n29485), .A2(n28667), .ZN(n4361) );
  OAI211_X1 U15394 ( .C1(n42049), .C2(n39062), .A(n4364), .B(n42043), .ZN(
        n39063) );
  NAND3_X1 U15395 ( .A1(n42049), .A2(n40049), .A3(n40295), .ZN(n4364) );
  NAND4_X2 U15396 ( .A1(n12859), .A2(n12860), .A3(n12858), .A4(n12857), .ZN(
        n16228) );
  NAND3_X2 U15397 ( .A1(n40161), .A2(n5770), .A3(n40160), .ZN(n43106) );
  XNOR2_X2 U15398 ( .A(n9364), .B(Key[8]), .ZN(n11353) );
  NAND2_X2 U15399 ( .A1(n9674), .A2(n4410), .ZN(n14472) );
  NAND4_X2 U15400 ( .A1(n22215), .A2(n22216), .A3(n22217), .A4(n22214), .ZN(
        n25778) );
  NOR2_X1 U15401 ( .A1(n45936), .A2(n43424), .ZN(n5938) );
  XNOR2_X1 U15402 ( .A(n16287), .B(n16190), .ZN(n7136) );
  NOR2_X1 U15403 ( .A1(n754), .A2(n23090), .ZN(n20852) );
  INV_X1 U15404 ( .A(n9015), .ZN(n7020) );
  INV_X1 U15405 ( .A(n9015), .ZN(n5335) );
  NAND4_X2 U15406 ( .A1(n22566), .A2(n4365), .A3(n22567), .A4(n22565), .ZN(
        n26264) );
  NAND2_X1 U15407 ( .A1(n22564), .A2(n22981), .ZN(n4365) );
  INV_X1 U15408 ( .A(n10586), .ZN(n5645) );
  NAND2_X1 U15409 ( .A1(n12258), .A2(n12255), .ZN(n4859) );
  NAND3_X1 U15410 ( .A1(n22073), .A2(n22932), .A3(n22074), .ZN(n22077) );
  INV_X1 U15411 ( .A(n48103), .ZN(n7766) );
  XNOR2_X1 U15412 ( .A(n28223), .B(n4366), .ZN(n25505) );
  INV_X1 U15413 ( .A(n28708), .ZN(n7909) );
  XNOR2_X1 U15415 ( .A(n17264), .B(n6583), .ZN(n16910) );
  XNOR2_X1 U15418 ( .A(n27196), .B(n4368), .ZN(n28047) );
  INV_X1 U15419 ( .A(n10708), .ZN(n4369) );
  NAND3_X1 U15420 ( .A1(n32796), .A2(n32795), .A3(n4370), .ZN(n32799) );
  NAND4_X4 U15421 ( .A1(n34202), .A2(n5526), .A3(n5525), .A4(n34201), .ZN(
        n40327) );
  NOR2_X1 U15424 ( .A1(n39411), .A2(n39207), .ZN(n39427) );
  INV_X1 U15425 ( .A(n27839), .ZN(n7825) );
  NAND4_X1 U15426 ( .A1(n7227), .A2(n12608), .A3(n4374), .A4(n4373), .ZN(n7228) );
  NAND2_X1 U15427 ( .A1(n12591), .A2(n12592), .ZN(n4373) );
  NAND2_X1 U15428 ( .A1(n12594), .A2(n12593), .ZN(n4374) );
  INV_X1 U15429 ( .A(n29989), .ZN(n31419) );
  NAND2_X1 U15431 ( .A1(n4375), .A2(n27719), .ZN(n24576) );
  OAI22_X1 U15432 ( .A1(n24569), .A2(n27720), .B1(n27627), .B2(n26803), .ZN(
        n4375) );
  NAND2_X1 U15434 ( .A1(n4377), .A2(n4376), .ZN(n37373) );
  NAND2_X1 U15435 ( .A1(n37371), .A2(n37587), .ZN(n4376) );
  NAND2_X1 U15436 ( .A1(n37372), .A2(n36232), .ZN(n4377) );
  XNOR2_X1 U15437 ( .A(n34810), .B(n2322), .ZN(n34828) );
  NOR3_X1 U15438 ( .A1(n49058), .A2(n2396), .A3(n4378), .ZN(n49061) );
  NAND4_X4 U15440 ( .A1(n8522), .A2(n5025), .A3(n19626), .A4(n8519), .ZN(
        n28311) );
  NAND2_X1 U15441 ( .A1(n2240), .A2(n27797), .ZN(n4381) );
  NAND2_X1 U15442 ( .A1(n12478), .A2(n12486), .ZN(n12479) );
  OAI21_X1 U15443 ( .B1(n40673), .B2(n40674), .A(n40672), .ZN(n40681) );
  NAND4_X1 U15445 ( .A1(n33011), .A2(n33012), .A3(n33010), .A4(n33009), .ZN(
        n33023) );
  INV_X1 U15447 ( .A(n27860), .ZN(n6346) );
  OAI21_X1 U15448 ( .B1(n4382), .B2(n2351), .A(n20695), .ZN(n20705) );
  NAND2_X1 U15449 ( .A1(n20693), .A2(n20694), .ZN(n4382) );
  NAND2_X1 U15450 ( .A1(n4383), .A2(n12787), .ZN(n13445) );
  NAND3_X2 U15451 ( .A1(n4384), .A2(n4385), .A3(n11758), .ZN(n17821) );
  INV_X1 U15452 ( .A(n4959), .ZN(n4384) );
  NAND3_X1 U15453 ( .A1(n4386), .A2(n30931), .A3(n29641), .ZN(n29580) );
  INV_X1 U15454 ( .A(n21613), .ZN(n8367) );
  NAND2_X1 U15455 ( .A1(n36552), .A2(n36541), .ZN(n8202) );
  XNOR2_X2 U15456 ( .A(n43935), .B(n43934), .ZN(n47058) );
  XNOR2_X1 U15458 ( .A(n4387), .B(n33426), .ZN(n6763) );
  XNOR2_X1 U15459 ( .A(n36868), .B(n37251), .ZN(n4387) );
  NAND2_X1 U15460 ( .A1(n4388), .A2(n30763), .ZN(n26845) );
  OAI22_X1 U15461 ( .A1(n27557), .A2(n30756), .B1(n30757), .B2(n30770), .ZN(
        n4388) );
  INV_X1 U15462 ( .A(n23701), .ZN(n23538) );
  NAND2_X1 U15464 ( .A1(n29054), .A2(n51490), .ZN(n30339) );
  NAND2_X1 U15465 ( .A1(n9313), .A2(n9316), .ZN(n5002) );
  OAI21_X1 U15467 ( .B1(n2419), .B2(n4389), .A(n19661), .ZN(n19669) );
  NAND2_X1 U15468 ( .A1(n19660), .A2(n19893), .ZN(n4389) );
  XNOR2_X1 U15469 ( .A(n4390), .B(n50424), .ZN(Plaintext[151]) );
  NAND2_X1 U15470 ( .A1(n32820), .A2(n4391), .ZN(n32824) );
  XNOR2_X1 U15471 ( .A(n4392), .B(n50770), .ZN(Plaintext[176]) );
  NAND2_X1 U15472 ( .A1(n50769), .A2(n50768), .ZN(n4392) );
  NAND4_X2 U15473 ( .A1(n22292), .A2(n22295), .A3(n22293), .A4(n22294), .ZN(
        n24757) );
  NOR2_X1 U15474 ( .A1(n44806), .A2(n4393), .ZN(n44807) );
  NAND3_X1 U15475 ( .A1(n44804), .A2(n49124), .A3(n44805), .ZN(n4393) );
  OR2_X1 U15476 ( .A1(n46596), .A2(n3107), .ZN(n4394) );
  XOR2_X1 U15477 ( .A(n15665), .B(n15664), .Z(n7863) );
  NAND2_X1 U15478 ( .A1(n6167), .A2(n21782), .ZN(n22703) );
  OR2_X2 U15479 ( .A1(n4395), .A2(n40509), .ZN(n42284) );
  NOR2_X1 U15480 ( .A1(n10784), .A2(n4439), .ZN(n6382) );
  OAI21_X1 U15481 ( .B1(n50786), .B2(n50762), .A(n50761), .ZN(n50763) );
  NAND3_X1 U15482 ( .A1(n4396), .A2(n11614), .A3(n2535), .ZN(n9284) );
  OAI21_X1 U15483 ( .B1(n11249), .B2(n11608), .A(n9277), .ZN(n4396) );
  NAND2_X1 U15484 ( .A1(n29173), .A2(n29156), .ZN(n27953) );
  NAND2_X1 U15485 ( .A1(n23518), .A2(n24414), .ZN(n24070) );
  NAND2_X1 U15486 ( .A1(n42158), .A2(n52092), .ZN(n4398) );
  NAND2_X1 U15487 ( .A1(n37819), .A2(n37818), .ZN(n4399) );
  NAND4_X2 U15488 ( .A1(n21826), .A2(n21827), .A3(n21825), .A4(n21824), .ZN(
        n25353) );
  INV_X1 U15489 ( .A(n52198), .ZN(n4400) );
  OAI211_X1 U15491 ( .C1(n12093), .C2(n12379), .A(n9687), .B(n12380), .ZN(
        n9688) );
  NAND4_X1 U15492 ( .A1(n20324), .A2(n4401), .A3(n20323), .A4(n21444), .ZN(
        n20332) );
  NAND2_X1 U15493 ( .A1(n21430), .A2(n4433), .ZN(n4401) );
  NAND2_X1 U15494 ( .A1(n8264), .A2(n37606), .ZN(n37607) );
  NAND4_X2 U15495 ( .A1(n27080), .A2(n27079), .A3(n27077), .A4(n27078), .ZN(
        n35503) );
  NAND4_X1 U15496 ( .A1(n46220), .A2(n4404), .A3(n4403), .A4(n4402), .ZN(
        n42709) );
  NAND2_X1 U15497 ( .A1(n42700), .A2(n46229), .ZN(n4402) );
  NAND2_X1 U15498 ( .A1(n49203), .A2(n46226), .ZN(n4403) );
  NOR2_X2 U15499 ( .A1(n14605), .A2(n13316), .ZN(n14603) );
  NOR2_X1 U15500 ( .A1(n30207), .A2(n29204), .ZN(n4405) );
  XNOR2_X1 U15501 ( .A(n4406), .B(n16325), .ZN(n16329) );
  XNOR2_X1 U15502 ( .A(n16727), .B(n16324), .ZN(n4406) );
  INV_X1 U15503 ( .A(n30048), .ZN(n7066) );
  OAI21_X1 U15504 ( .B1(n41201), .B2(n41202), .A(n41200), .ZN(n41204) );
  NAND2_X1 U15505 ( .A1(n10050), .A2(n9863), .ZN(n9864) );
  NAND3_X1 U15506 ( .A1(n9856), .A2(n10120), .A3(n6005), .ZN(n9863) );
  NAND4_X1 U15507 ( .A1(n4408), .A2(n40561), .A3(n40560), .A4(n40562), .ZN(
        n40579) );
  OAI21_X1 U15508 ( .B1(n40552), .B2(n40551), .A(n40550), .ZN(n4408) );
  NAND2_X1 U15509 ( .A1(n38587), .A2(n38599), .ZN(n38590) );
  XNOR2_X1 U15512 ( .A(n16953), .B(n16952), .ZN(n16954) );
  NAND2_X1 U15515 ( .A1(n40564), .A2(n40566), .ZN(n40310) );
  OR3_X1 U15516 ( .A1(n13947), .A2(n2173), .A3(n13948), .ZN(n4595) );
  NOR2_X1 U15517 ( .A1(n19612), .A2(n2352), .ZN(n4412) );
  NAND3_X1 U15518 ( .A1(n20794), .A2(n21388), .A3(n4414), .ZN(n20796) );
  NAND4_X2 U15519 ( .A1(n21031), .A2(n21032), .A3(n21034), .A4(n21033), .ZN(
        n26540) );
  OR2_X2 U15520 ( .A1(n41478), .A2(n41477), .ZN(n47841) );
  XOR2_X1 U15521 ( .A(n27377), .B(n27481), .Z(n5663) );
  NOR2_X1 U15523 ( .A1(n4418), .A2(n4417), .ZN(n4416) );
  NAND4_X1 U15525 ( .A1(n21371), .A2(n21373), .A3(n21372), .A4(n21389), .ZN(
        n21381) );
  NAND2_X1 U15526 ( .A1(n6207), .A2(n23902), .ZN(n23141) );
  NAND3_X1 U15527 ( .A1(n10136), .A2(n10135), .A3(n10913), .ZN(n10141) );
  NAND2_X1 U15528 ( .A1(n21253), .A2(n17079), .ZN(n19093) );
  NAND3_X1 U15530 ( .A1(n6039), .A2(n13902), .A3(n6038), .ZN(n4420) );
  NAND2_X1 U15531 ( .A1(n5498), .A2(n4422), .ZN(n31528) );
  XNOR2_X2 U15532 ( .A(n9174), .B(Key[185]), .ZN(n11978) );
  INV_X1 U15533 ( .A(n28487), .ZN(n5912) );
  NAND2_X1 U15534 ( .A1(n30463), .A2(n30464), .ZN(n30465) );
  NAND2_X1 U15535 ( .A1(n4424), .A2(n13587), .ZN(n13591) );
  XNOR2_X1 U15536 ( .A(n27225), .B(n8657), .ZN(n27227) );
  XNOR2_X2 U15537 ( .A(n4425), .B(n28281), .ZN(n30346) );
  XNOR2_X1 U15538 ( .A(n28282), .B(n28280), .ZN(n4425) );
  NOR2_X1 U15539 ( .A1(n5813), .A2(n20014), .ZN(n15091) );
  NOR2_X1 U15540 ( .A1(n8794), .A2(n7055), .ZN(n7053) );
  NAND2_X1 U15541 ( .A1(n6217), .A2(n8016), .ZN(n6216) );
  NAND2_X1 U15542 ( .A1(n47089), .A2(n47095), .ZN(n5275) );
  NAND4_X1 U15543 ( .A1(n45526), .A2(n4428), .A3(n45833), .A4(n45525), .ZN(
        n45529) );
  NAND3_X1 U15544 ( .A1(n6215), .A2(n34999), .A3(n34998), .ZN(n35000) );
  XNOR2_X2 U15545 ( .A(n9286), .B(Key[183]), .ZN(n10072) );
  INV_X1 U15546 ( .A(n39291), .ZN(n7772) );
  NAND2_X2 U15547 ( .A1(n4430), .A2(n18881), .ZN(n23317) );
  INV_X1 U15548 ( .A(n35973), .ZN(n37371) );
  INV_X1 U15549 ( .A(n21227), .ZN(n19113) );
  BUF_X1 U15550 ( .A(n35004), .Z(n39129) );
  INV_X1 U15551 ( .A(n10915), .ZN(n8840) );
  INV_X1 U15552 ( .A(n20230), .ZN(n15928) );
  INV_X1 U15553 ( .A(n34720), .ZN(n33187) );
  XNOR2_X1 U15554 ( .A(n15867), .B(n15866), .ZN(n15868) );
  AOI22_X1 U15555 ( .A1(n7475), .A2(n26721), .B1(n29444), .B2(n27026), .ZN(
        n6839) );
  AND3_X1 U15556 ( .A1(n27842), .A2(n6839), .A3(n6838), .ZN(n6837) );
  NAND2_X1 U15557 ( .A1(n22933), .A2(n4432), .ZN(n22939) );
  NAND3_X1 U15558 ( .A1(n22930), .A2(n22943), .A3(n23049), .ZN(n4432) );
  NAND2_X1 U15559 ( .A1(n6681), .A2(n4435), .ZN(n26067) );
  INV_X1 U15560 ( .A(n15279), .ZN(n14938) );
  NAND2_X1 U15562 ( .A1(n19475), .A2(n18969), .ZN(n16308) );
  NAND4_X2 U15563 ( .A1(n32141), .A2(n8222), .A3(n8223), .A4(n32132), .ZN(
        n35331) );
  INV_X1 U15567 ( .A(n5430), .ZN(n4567) );
  NAND2_X1 U15568 ( .A1(n13475), .A2(n15044), .ZN(n13794) );
  NAND2_X1 U15569 ( .A1(n4438), .A2(n32883), .ZN(n29052) );
  NAND2_X1 U15572 ( .A1(n12640), .A2(n6571), .ZN(n12625) );
  NAND3_X1 U15573 ( .A1(n21407), .A2(n21567), .A3(n21568), .ZN(n21409) );
  INV_X1 U15574 ( .A(n11575), .ZN(n11528) );
  NAND4_X2 U15575 ( .A1(n6281), .A2(n15558), .A3(n6280), .A4(n15556), .ZN(
        n24452) );
  NAND2_X1 U15576 ( .A1(n6385), .A2(n4440), .ZN(n4439) );
  NAND2_X1 U15577 ( .A1(n10786), .A2(n10785), .ZN(n4440) );
  NAND3_X1 U15581 ( .A1(n4442), .A2(n24328), .A3(n23380), .ZN(n23381) );
  AOI21_X1 U15583 ( .B1(n4906), .B2(n51545), .A(n4905), .ZN(n31582) );
  NAND4_X1 U15584 ( .A1(n29943), .A2(n29944), .A3(n30387), .A4(n30698), .ZN(
        n4444) );
  INV_X1 U15585 ( .A(n10514), .ZN(n10111) );
  NAND2_X1 U15586 ( .A1(n9482), .A2(n10096), .ZN(n10514) );
  NAND2_X2 U15587 ( .A1(n5406), .A2(n20786), .ZN(n23950) );
  NOR2_X1 U15588 ( .A1(n4446), .A2(n4445), .ZN(n14932) );
  NOR2_X1 U15590 ( .A1(n4449), .A2(n4448), .ZN(n4447) );
  NOR2_X1 U15591 ( .A1(n20851), .A2(n20850), .ZN(n4448) );
  INV_X1 U15593 ( .A(n21563), .ZN(n20781) );
  NAND2_X1 U15594 ( .A1(n20600), .A2(n51755), .ZN(n21563) );
  XNOR2_X1 U15595 ( .A(n51097), .B(n42635), .ZN(n8269) );
  INV_X1 U15596 ( .A(n28898), .ZN(n27997) );
  NAND2_X1 U15597 ( .A1(n37557), .A2(n37560), .ZN(n36267) );
  NAND2_X1 U15598 ( .A1(n27720), .A2(n27721), .ZN(n27722) );
  NAND4_X2 U15599 ( .A1(n4773), .A2(n7893), .A3(n7892), .A4(n11356), .ZN(
        n14454) );
  NAND2_X1 U15600 ( .A1(n21968), .A2(n20994), .ZN(n4452) );
  NAND2_X1 U15601 ( .A1(n21971), .A2(n20993), .ZN(n4453) );
  XNOR2_X2 U15602 ( .A(n44950), .B(n44949), .ZN(n46693) );
  XNOR2_X1 U15604 ( .A(n4455), .B(n27182), .ZN(n27184) );
  XNOR2_X1 U15605 ( .A(n27181), .B(n27180), .ZN(n4455) );
  NAND2_X1 U15606 ( .A1(n6634), .A2(n13100), .ZN(n4456) );
  NAND2_X1 U15608 ( .A1(n20068), .A2(n20067), .ZN(n4457) );
  NAND2_X1 U15609 ( .A1(n20069), .A2(n4459), .ZN(n4458) );
  NAND2_X1 U15610 ( .A1(n4461), .A2(n14149), .ZN(n14145) );
  INV_X1 U15611 ( .A(n5994), .ZN(n5832) );
  NOR2_X1 U15612 ( .A1(n29868), .A2(n30429), .ZN(n29864) );
  AOI22_X1 U15613 ( .A1(n718), .A2(n2349), .B1(n32436), .B2(n32437), .ZN(
        n32451) );
  NAND2_X1 U15614 ( .A1(n4462), .A2(n23191), .ZN(n4877) );
  NAND2_X1 U15615 ( .A1(n24190), .A2(n23866), .ZN(n23191) );
  XOR2_X1 U15616 ( .A(n24870), .B(n24869), .Z(n7613) );
  XNOR2_X1 U15618 ( .A(n14569), .B(n14113), .ZN(n5956) );
  NAND4_X4 U15619 ( .A1(n9392), .A2(n9390), .A3(n9391), .A4(n4463), .ZN(n14664) );
  INV_X1 U15621 ( .A(n21584), .ZN(n21412) );
  NAND2_X1 U15622 ( .A1(n17529), .A2(n4467), .ZN(n17493) );
  XNOR2_X1 U15623 ( .A(n6581), .B(n37304), .ZN(n7828) );
  NAND2_X1 U15624 ( .A1(n40203), .A2(n40119), .ZN(n39551) );
  XNOR2_X1 U15625 ( .A(n34177), .B(n34176), .ZN(n7827) );
  NAND2_X1 U15626 ( .A1(n32962), .A2(n8125), .ZN(n5227) );
  NAND2_X1 U15627 ( .A1(n23606), .A2(n17418), .ZN(n23614) );
  NAND2_X1 U15628 ( .A1(n3550), .A2(n43669), .ZN(n38805) );
  NAND2_X1 U15629 ( .A1(n8885), .A2(n8886), .ZN(n11108) );
  NAND2_X1 U15630 ( .A1(n4468), .A2(n22880), .ZN(n22217) );
  NAND3_X1 U15631 ( .A1(n38690), .A2(n38691), .A3(n38692), .ZN(n4469) );
  INV_X1 U15632 ( .A(n8948), .ZN(n11454) );
  NAND2_X1 U15633 ( .A1(n4470), .A2(n19890), .ZN(n7256) );
  XNOR2_X1 U15634 ( .A(n4472), .B(n44488), .ZN(n44490) );
  XNOR2_X1 U15635 ( .A(n45076), .B(n44482), .ZN(n4472) );
  NOR2_X1 U15636 ( .A1(n46430), .A2(n4473), .ZN(n46431) );
  NAND4_X1 U15637 ( .A1(n46427), .A2(n48720), .A3(n46429), .A4(n46428), .ZN(
        n4473) );
  AOI22_X1 U15638 ( .A1(n48850), .A2(n48920), .B1(n48851), .B2(n48852), .ZN(
        n48857) );
  NAND2_X1 U15639 ( .A1(n33175), .A2(n36375), .ZN(n4474) );
  NAND3_X1 U15640 ( .A1(n5380), .A2(n13512), .A3(n13511), .ZN(n13517) );
  NAND2_X1 U15641 ( .A1(n740), .A2(n51109), .ZN(n29203) );
  INV_X1 U15642 ( .A(n50482), .ZN(n4692) );
  NAND2_X1 U15643 ( .A1(n30752), .A2(n30751), .ZN(n4475) );
  NAND2_X1 U15644 ( .A1(n30753), .A2(n24348), .ZN(n4476) );
  NAND4_X2 U15645 ( .A1(n11285), .A2(n11286), .A3(n11284), .A4(n11283), .ZN(
        n14393) );
  XNOR2_X1 U15646 ( .A(n4477), .B(n25356), .ZN(n25364) );
  XNOR2_X1 U15647 ( .A(n25362), .B(n25355), .ZN(n4477) );
  NAND3_X1 U15648 ( .A1(n32800), .A2(n32799), .A3(n4478), .ZN(n5632) );
  AOI22_X1 U15649 ( .A1(n32792), .A2(n32791), .B1(n32789), .B2(n32790), .ZN(
        n4478) );
  NAND2_X1 U15650 ( .A1(n23997), .A2(n24002), .ZN(n4479) );
  XNOR2_X1 U15651 ( .A(n4481), .B(n33381), .ZN(n33385) );
  XNOR2_X1 U15652 ( .A(n35337), .B(n33380), .ZN(n4481) );
  INV_X1 U15653 ( .A(n32669), .ZN(n31180) );
  NAND2_X1 U15654 ( .A1(n31169), .A2(n31454), .ZN(n32669) );
  NAND2_X1 U15655 ( .A1(n21253), .A2(n19472), .ZN(n19089) );
  OAI21_X1 U15656 ( .B1(n12546), .B2(n12545), .A(n12544), .ZN(n12550) );
  XNOR2_X1 U15657 ( .A(n4483), .B(n44516), .ZN(n41659) );
  XNOR2_X1 U15658 ( .A(n41602), .B(n43006), .ZN(n4483) );
  NAND2_X1 U15659 ( .A1(n7936), .A2(n10199), .ZN(n7942) );
  NAND2_X1 U15660 ( .A1(n14633), .A2(n13667), .ZN(n13658) );
  NAND3_X1 U15662 ( .A1(n22425), .A2(n22424), .A3(n4485), .ZN(n4484) );
  NAND2_X1 U15663 ( .A1(n39252), .A2(n39253), .ZN(n39254) );
  NAND2_X1 U15664 ( .A1(n12516), .A2(n51709), .ZN(n11549) );
  NAND4_X2 U15665 ( .A1(n4488), .A2(n13365), .A3(n13363), .A4(n13364), .ZN(
        n16628) );
  NAND2_X1 U15666 ( .A1(n13350), .A2(n13354), .ZN(n4488) );
  NAND2_X1 U15667 ( .A1(n32841), .A2(n31911), .ZN(n32851) );
  XNOR2_X1 U15668 ( .A(n8282), .B(n28113), .ZN(n4491) );
  INV_X1 U15669 ( .A(Ciphertext[14]), .ZN(n8396) );
  INV_X1 U15670 ( .A(n28145), .ZN(n30285) );
  NAND2_X1 U15671 ( .A1(n46873), .A2(n47110), .ZN(n6587) );
  XNOR2_X2 U15672 ( .A(Key[80]), .B(Ciphertext[109]), .ZN(n10065) );
  NAND2_X1 U15673 ( .A1(n13449), .A2(n12790), .ZN(n13441) );
  XNOR2_X1 U15675 ( .A(n35474), .B(n4828), .ZN(n4492) );
  NOR2_X1 U15676 ( .A1(n5750), .A2(n19636), .ZN(n5749) );
  NAND2_X1 U15677 ( .A1(n4493), .A2(n28758), .ZN(n29943) );
  XNOR2_X1 U15680 ( .A(n17650), .B(n17649), .ZN(n4495) );
  NAND4_X1 U15683 ( .A1(n6475), .A2(n6474), .A3(n38749), .A4(n4496), .ZN(n5488) );
  NAND3_X2 U15684 ( .A1(n4497), .A2(n4498), .A3(n8846), .ZN(n14287) );
  NAND2_X1 U15685 ( .A1(n8837), .A2(n10217), .ZN(n4497) );
  NAND3_X1 U15686 ( .A1(n4499), .A2(n30734), .A3(n30733), .ZN(n30735) );
  INV_X1 U15687 ( .A(n30732), .ZN(n4499) );
  NAND2_X1 U15688 ( .A1(n30382), .A2(n30376), .ZN(n30732) );
  NAND2_X1 U15689 ( .A1(n8049), .A2(n2378), .ZN(n11416) );
  XNOR2_X2 U15691 ( .A(n31674), .B(n33728), .ZN(n37023) );
  XNOR2_X1 U15692 ( .A(n4500), .B(n16726), .ZN(n16728) );
  XNOR2_X1 U15693 ( .A(n16721), .B(n16722), .ZN(n4500) );
  AND3_X1 U15694 ( .A1(n12940), .A2(n12939), .A3(n12942), .ZN(n4717) );
  INV_X1 U15695 ( .A(n13708), .ZN(n10500) );
  NOR2_X1 U15696 ( .A1(n5038), .A2(n51106), .ZN(n5040) );
  XNOR2_X1 U15697 ( .A(n4503), .B(n50964), .ZN(Plaintext[191]) );
  INV_X1 U15699 ( .A(n18240), .ZN(n4505) );
  XNOR2_X1 U15701 ( .A(n16438), .B(n15721), .ZN(n4506) );
  NAND2_X1 U15702 ( .A1(n30931), .A2(n31067), .ZN(n31509) );
  INV_X1 U15703 ( .A(n15542), .ZN(n18483) );
  INV_X1 U15705 ( .A(n35402), .ZN(n4993) );
  INV_X1 U15706 ( .A(n49138), .ZN(n49151) );
  NOR2_X1 U15707 ( .A1(n13709), .A2(n15131), .ZN(n14993) );
  OAI211_X1 U15708 ( .C1(n36283), .C2(n39064), .A(n40287), .B(n7158), .ZN(
        n36284) );
  NAND3_X1 U15709 ( .A1(n21358), .A2(n20768), .A3(n21599), .ZN(n19926) );
  XNOR2_X1 U15712 ( .A(n4507), .B(n43322), .ZN(n43351) );
  XNOR2_X1 U15713 ( .A(n43321), .B(n45070), .ZN(n4507) );
  NAND2_X1 U15714 ( .A1(n38522), .A2(n51487), .ZN(n38513) );
  INV_X1 U15715 ( .A(n23675), .ZN(n6103) );
  INV_X1 U15716 ( .A(n8490), .ZN(n5150) );
  NAND2_X1 U15717 ( .A1(n25789), .A2(n26668), .ZN(n26679) );
  NAND2_X1 U15718 ( .A1(n7812), .A2(n11234), .ZN(n4508) );
  XNOR2_X1 U15719 ( .A(n35549), .B(n35548), .ZN(n5516) );
  XNOR2_X1 U15720 ( .A(n4509), .B(n44056), .ZN(n8293) );
  XNOR2_X1 U15721 ( .A(n44068), .B(n44067), .ZN(n4509) );
  NAND2_X1 U15722 ( .A1(n5486), .A2(n38618), .ZN(n5485) );
  BUF_X1 U15723 ( .A(n25352), .Z(n25504) );
  XNOR2_X2 U15724 ( .A(n24858), .B(n5082), .ZN(n30296) );
  XNOR2_X1 U15725 ( .A(n15294), .B(n15293), .ZN(n15297) );
  INV_X1 U15726 ( .A(n39427), .ZN(n39432) );
  INV_X1 U15727 ( .A(n37618), .ZN(n4512) );
  NOR2_X2 U15728 ( .A1(n7780), .A2(n12690), .ZN(n12440) );
  NAND2_X1 U15729 ( .A1(n31162), .A2(n32620), .ZN(n4513) );
  NAND2_X1 U15732 ( .A1(n4516), .A2(n19344), .ZN(n20514) );
  XNOR2_X2 U15733 ( .A(n7125), .B(n15548), .ZN(n19344) );
  NAND2_X1 U15734 ( .A1(n8963), .A2(n11928), .ZN(n8967) );
  NOR2_X1 U15735 ( .A1(n52121), .A2(n7957), .ZN(n29950) );
  AOI21_X1 U15736 ( .B1(n40941), .B2(n41534), .A(n5215), .ZN(n5214) );
  NAND2_X1 U15737 ( .A1(n19122), .A2(n19455), .ZN(n19783) );
  NAND2_X1 U15739 ( .A1(n6346), .A2(n6080), .ZN(n29479) );
  XNOR2_X1 U15740 ( .A(n43802), .B(n43063), .ZN(n43064) );
  OAI211_X1 U15741 ( .C1(n22548), .C2(n5290), .A(n22067), .B(n5289), .ZN(
        n21313) );
  NAND2_X1 U15742 ( .A1(n18990), .A2(n4521), .ZN(n18994) );
  XNOR2_X1 U15743 ( .A(n43394), .B(n43393), .ZN(n4522) );
  NAND2_X1 U15744 ( .A1(n39361), .A2(n4523), .ZN(n39191) );
  NAND2_X1 U15745 ( .A1(n9162), .A2(n14633), .ZN(n13662) );
  XNOR2_X1 U15746 ( .A(n4524), .B(n45519), .ZN(Plaintext[75]) );
  XNOR2_X2 U15747 ( .A(n7813), .B(n18417), .ZN(n7484) );
  XNOR2_X1 U15750 ( .A(n35477), .B(n4525), .ZN(n35487) );
  XNOR2_X1 U15751 ( .A(n35478), .B(n35485), .ZN(n4525) );
  INV_X1 U15752 ( .A(n23956), .ZN(n22241) );
  INV_X1 U15753 ( .A(n48791), .ZN(n48833) );
  NAND2_X1 U15754 ( .A1(n29642), .A2(n3099), .ZN(n29643) );
  XNOR2_X1 U15755 ( .A(n40467), .B(n43915), .ZN(n7622) );
  XNOR2_X2 U15756 ( .A(n18599), .B(n17822), .ZN(n17378) );
  NOR2_X1 U15757 ( .A1(n20075), .A2(n4459), .ZN(n19493) );
  XNOR2_X1 U15758 ( .A(n24911), .B(n7182), .ZN(n7181) );
  XNOR2_X1 U15760 ( .A(n42625), .B(n42624), .ZN(n4530) );
  NAND2_X1 U15763 ( .A1(n27755), .A2(n27764), .ZN(n27757) );
  NAND2_X1 U15765 ( .A1(n12241), .A2(n12257), .ZN(n4533) );
  XNOR2_X1 U15766 ( .A(n16720), .B(n4534), .ZN(n15474) );
  NAND2_X1 U15768 ( .A1(n18224), .A2(n21291), .ZN(n8576) );
  NOR2_X1 U15769 ( .A1(n23664), .A2(n8524), .ZN(n23665) );
  NAND4_X2 U15770 ( .A1(n27770), .A2(n27769), .A3(n27771), .A4(n5261), .ZN(
        n30593) );
  NAND2_X1 U15771 ( .A1(n4538), .A2(n38447), .ZN(n37363) );
  NAND4_X2 U15773 ( .A1(n46966), .A2(n7880), .A3(n7882), .A4(n7881), .ZN(
        n50542) );
  INV_X1 U15774 ( .A(n47371), .ZN(n50007) );
  XNOR2_X1 U15775 ( .A(n25936), .B(n25952), .ZN(n7834) );
  NAND3_X1 U15777 ( .A1(n47098), .A2(n47094), .A3(n669), .ZN(n47101) );
  OAI22_X1 U15778 ( .A1(n47108), .A2(n7919), .B1(n44578), .B2(n47109), .ZN(
        n47114) );
  NAND2_X1 U15779 ( .A1(n13297), .A2(n13729), .ZN(n11048) );
  XNOR2_X1 U15780 ( .A(n11035), .B(n10008), .ZN(n4540) );
  AND2_X1 U15781 ( .A1(n4673), .A2(n29073), .ZN(n4925) );
  NAND2_X1 U15782 ( .A1(n4541), .A2(n47000), .ZN(n46896) );
  OAI22_X1 U15783 ( .A1(n46892), .A2(n47159), .B1(n46891), .B2(n47154), .ZN(
        n4541) );
  AND2_X1 U15784 ( .A1(n10139), .A2(n10922), .ZN(n4593) );
  XNOR2_X1 U15785 ( .A(n42383), .B(n42382), .ZN(n44055) );
  INV_X1 U15786 ( .A(n30344), .ZN(n30354) );
  NAND2_X1 U15787 ( .A1(n12549), .A2(n12532), .ZN(n11096) );
  NOR2_X1 U15788 ( .A1(n30249), .A2(n6730), .ZN(n29148) );
  INV_X1 U15789 ( .A(n38998), .ZN(n5520) );
  XNOR2_X1 U15790 ( .A(n6170), .B(n6169), .ZN(n35890) );
  INV_X1 U15791 ( .A(n7905), .ZN(n7904) );
  INV_X1 U15792 ( .A(n11052), .ZN(n4822) );
  INV_X1 U15793 ( .A(n22832), .ZN(n8586) );
  XNOR2_X1 U15794 ( .A(n43642), .B(n42768), .ZN(n5532) );
  NAND3_X1 U15795 ( .A1(n49576), .A2(n49575), .A3(n4543), .ZN(n49578) );
  NAND2_X1 U15796 ( .A1(n49573), .A2(n4544), .ZN(n4543) );
  NAND3_X1 U15797 ( .A1(n42992), .A2(n2242), .A3(n42993), .ZN(n4545) );
  NOR2_X1 U15798 ( .A1(n39515), .A2(n40828), .ZN(n39074) );
  NAND2_X1 U15799 ( .A1(n640), .A2(n14454), .ZN(n14099) );
  NAND2_X1 U15800 ( .A1(n12166), .A2(n9589), .ZN(n11324) );
  INV_X1 U15801 ( .A(n14547), .ZN(n13361) );
  NAND2_X1 U15802 ( .A1(n14370), .A2(n14533), .ZN(n14547) );
  NAND2_X1 U15803 ( .A1(n14664), .A2(n11315), .ZN(n12950) );
  XNOR2_X2 U15804 ( .A(n9362), .B(Key[111]), .ZN(n12373) );
  NOR2_X1 U15805 ( .A1(n5354), .A2(n39523), .ZN(n4547) );
  XNOR2_X1 U15806 ( .A(n43162), .B(n43161), .ZN(n43181) );
  OAI211_X1 U15808 ( .C1(n37656), .C2(n37655), .A(n6748), .B(n39301), .ZN(
        n7489) );
  NAND2_X1 U15809 ( .A1(n8824), .A2(n10162), .ZN(n11023) );
  NAND2_X1 U15811 ( .A1(n30241), .A2(n7548), .ZN(n30242) );
  NAND2_X1 U15812 ( .A1(n30251), .A2(n5169), .ZN(n30241) );
  NAND2_X1 U15813 ( .A1(n9495), .A2(n11704), .ZN(n11203) );
  OAI21_X1 U15815 ( .B1(n29072), .B2(n29071), .A(n29070), .ZN(n8188) );
  NAND2_X1 U15816 ( .A1(n23184), .A2(n23167), .ZN(n22793) );
  INV_X1 U15818 ( .A(n29158), .ZN(n29167) );
  NAND2_X1 U15819 ( .A1(n29147), .A2(n626), .ZN(n29158) );
  NAND2_X1 U15820 ( .A1(n12571), .A2(n12570), .ZN(n4550) );
  NAND2_X1 U15821 ( .A1(n4551), .A2(n29171), .ZN(n29178) );
  NAND3_X1 U15822 ( .A1(n29168), .A2(n29170), .A3(n29169), .ZN(n4551) );
  OR2_X1 U15823 ( .A1(n26348), .A2(n29085), .ZN(n32134) );
  NAND4_X2 U15824 ( .A1(n11156), .A2(n11155), .A3(n11154), .A4(n11153), .ZN(
        n17965) );
  AND2_X1 U15825 ( .A1(n4553), .A2(n41583), .ZN(n41585) );
  NAND3_X1 U15826 ( .A1(n42011), .A2(n41582), .A3(n7709), .ZN(n4553) );
  XNOR2_X1 U15827 ( .A(n29385), .B(n35265), .ZN(n35517) );
  INV_X1 U15828 ( .A(Ciphertext[161]), .ZN(n8563) );
  INV_X1 U15830 ( .A(n12317), .ZN(n4617) );
  XNOR2_X1 U15831 ( .A(n27477), .B(n42266), .ZN(n4688) );
  XNOR2_X1 U15832 ( .A(n4556), .B(n33695), .ZN(n33780) );
  XNOR2_X1 U15833 ( .A(n34161), .B(n33694), .ZN(n4556) );
  OR2_X2 U15834 ( .A1(n13330), .A2(n13329), .ZN(n18755) );
  NAND2_X1 U15835 ( .A1(n12654), .A2(n12653), .ZN(n4559) );
  NAND2_X1 U15836 ( .A1(n12656), .A2(n12655), .ZN(n4560) );
  NAND2_X1 U15838 ( .A1(n6565), .A2(n6570), .ZN(n6564) );
  NAND2_X1 U15839 ( .A1(n11780), .A2(n13841), .ZN(n9691) );
  NAND3_X1 U15840 ( .A1(n13677), .A2(n13024), .A3(n13025), .ZN(n14244) );
  INV_X1 U15842 ( .A(n41734), .ZN(n4561) );
  NOR3_X1 U15843 ( .A1(n50767), .A2(n4563), .A3(n4562), .ZN(n50768) );
  INV_X1 U15844 ( .A(n50766), .ZN(n4563) );
  XNOR2_X2 U15845 ( .A(n42778), .B(n41494), .ZN(n43929) );
  AOI21_X1 U15846 ( .B1(n22417), .B2(n23032), .A(n5102), .ZN(n22433) );
  INV_X1 U15847 ( .A(n6329), .ZN(n12047) );
  NAND2_X1 U15848 ( .A1(n15047), .A2(n13483), .ZN(n15033) );
  XNOR2_X1 U15850 ( .A(n7872), .B(n7871), .ZN(n7870) );
  NAND3_X2 U15851 ( .A1(n4567), .A2(n4566), .A3(n38236), .ZN(n44209) );
  XNOR2_X1 U15852 ( .A(n16650), .B(n356), .ZN(n16651) );
  NAND3_X1 U15853 ( .A1(n5292), .A2(n5291), .A3(n21847), .ZN(n5293) );
  OR2_X2 U15854 ( .A1(n24199), .A2(n24198), .ZN(n25937) );
  NAND2_X1 U15855 ( .A1(n4569), .A2(n36427), .ZN(n6598) );
  NAND3_X1 U15856 ( .A1(n36060), .A2(n34654), .A3(n34655), .ZN(n4569) );
  INV_X1 U15857 ( .A(n30575), .ZN(n31830) );
  NAND2_X1 U15858 ( .A1(n31816), .A2(n31033), .ZN(n30575) );
  NAND4_X2 U15860 ( .A1(n23064), .A2(n23065), .A3(n23063), .A4(n23062), .ZN(
        n28038) );
  AOI21_X1 U15862 ( .B1(n36432), .B2(n4575), .A(n36431), .ZN(n36433) );
  NAND3_X1 U15863 ( .A1(n2472), .A2(n36617), .A3(n4576), .ZN(n4575) );
  NAND4_X2 U15864 ( .A1(n19152), .A2(n19154), .A3(n19155), .A4(n19153), .ZN(
        n28287) );
  INV_X1 U15865 ( .A(Ciphertext[116]), .ZN(n6123) );
  NOR2_X1 U15866 ( .A1(n26787), .A2(n26691), .ZN(n27742) );
  NAND3_X1 U15867 ( .A1(n11464), .A2(n11470), .A3(n11234), .ZN(n9325) );
  XNOR2_X1 U15869 ( .A(n4580), .B(n6131), .ZN(n35269) );
  XNOR2_X1 U15870 ( .A(n35266), .B(n35267), .ZN(n4580) );
  OAI22_X1 U15872 ( .A1(n35899), .A2(n38262), .B1(n6457), .B2(n38257), .ZN(
        n4582) );
  INV_X1 U15873 ( .A(n9981), .ZN(n11670) );
  OR2_X1 U15874 ( .A1(n29187), .A2(n25479), .ZN(n8424) );
  INV_X1 U15875 ( .A(n20451), .ZN(n20336) );
  INV_X1 U15876 ( .A(n8015), .ZN(n8014) );
  NAND3_X1 U15877 ( .A1(n22965), .A2(n22963), .A3(n22964), .ZN(n22970) );
  XNOR2_X1 U15878 ( .A(n4583), .B(n27341), .ZN(n23980) );
  XNOR2_X1 U15879 ( .A(n25475), .B(n25466), .ZN(n4583) );
  NAND2_X1 U15880 ( .A1(n4584), .A2(n14598), .ZN(n6350) );
  NAND2_X1 U15882 ( .A1(n719), .A2(n32883), .ZN(n32865) );
  INV_X1 U15883 ( .A(n6945), .ZN(n6658) );
  INV_X1 U15884 ( .A(n22441), .ZN(n22445) );
  NAND3_X1 U15886 ( .A1(n20605), .A2(n5167), .A3(n19988), .ZN(n19990) );
  NAND3_X1 U15887 ( .A1(n46703), .A2(n46699), .A3(n46701), .ZN(n44835) );
  XNOR2_X1 U15888 ( .A(n33148), .B(n2387), .ZN(n33057) );
  XNOR2_X1 U15889 ( .A(n33645), .B(n33048), .ZN(n33148) );
  XNOR2_X1 U15890 ( .A(n15294), .B(n4590), .ZN(n14677) );
  XNOR2_X1 U15891 ( .A(n16770), .B(n15295), .ZN(n4590) );
  NAND2_X1 U15892 ( .A1(n29883), .A2(n29784), .ZN(n30360) );
  XNOR2_X1 U15893 ( .A(n33452), .B(n33451), .ZN(n4591) );
  AND3_X1 U15894 ( .A1(n9571), .A2(n9566), .A3(n12625), .ZN(n8497) );
  XNOR2_X1 U15895 ( .A(n17819), .B(n16148), .ZN(n4592) );
  AOI21_X1 U15896 ( .B1(n10141), .B2(n10140), .A(n4593), .ZN(n10156) );
  NAND2_X1 U15897 ( .A1(n12384), .A2(n11354), .ZN(n12088) );
  NAND2_X1 U15898 ( .A1(n14546), .A2(n4594), .ZN(n14549) );
  NAND2_X1 U15899 ( .A1(n4595), .A2(n13932), .ZN(n9883) );
  NAND2_X1 U15900 ( .A1(n786), .A2(n12893), .ZN(n12791) );
  XNOR2_X2 U15902 ( .A(n28132), .B(n28133), .ZN(n28862) );
  AND3_X1 U15903 ( .A1(n20773), .A2(n20772), .A3(n20771), .ZN(n7288) );
  NAND2_X1 U15904 ( .A1(n23143), .A2(n23135), .ZN(n22796) );
  OAI21_X1 U15905 ( .B1(n27038), .B2(n26071), .A(n26639), .ZN(n5544) );
  NAND2_X1 U15907 ( .A1(n20354), .A2(n20427), .ZN(n20348) );
  OR2_X2 U15909 ( .A1(n6435), .A2(n9066), .ZN(n8670) );
  AND2_X1 U15910 ( .A1(n11808), .A2(n7767), .ZN(n7769) );
  NAND2_X1 U15911 ( .A1(n16841), .A2(n2414), .ZN(n13539) );
  NAND2_X1 U15912 ( .A1(n19387), .A2(n18012), .ZN(n16841) );
  NAND2_X1 U15913 ( .A1(n50447), .A2(n7114), .ZN(n50415) );
  NAND2_X1 U15914 ( .A1(n11372), .A2(n10709), .ZN(n4601) );
  OR2_X2 U15915 ( .A1(n26779), .A2(n29467), .ZN(n29460) );
  OAI21_X1 U15916 ( .B1(n13817), .B2(n8227), .A(n14310), .ZN(n5338) );
  INV_X1 U15917 ( .A(n36617), .ZN(n36421) );
  XNOR2_X2 U15919 ( .A(n9000), .B(Key[13]), .ZN(n12278) );
  INV_X1 U15920 ( .A(n10234), .ZN(n4797) );
  XNOR2_X1 U15921 ( .A(n7358), .B(n36867), .ZN(n4602) );
  NAND2_X1 U15922 ( .A1(n5151), .A2(n39429), .ZN(n39207) );
  NAND2_X1 U15923 ( .A1(n28470), .A2(n4603), .ZN(n28477) );
  NAND2_X1 U15924 ( .A1(n28469), .A2(n8390), .ZN(n4603) );
  NAND2_X1 U15925 ( .A1(n32962), .A2(n32771), .ZN(n28469) );
  INV_X1 U15926 ( .A(Ciphertext[10]), .ZN(n8487) );
  INV_X1 U15927 ( .A(n21615), .ZN(n20697) );
  INV_X1 U15928 ( .A(n10569), .ZN(n10015) );
  INV_X1 U15929 ( .A(n9763), .ZN(n4604) );
  INV_X2 U15930 ( .A(n49114), .ZN(n49127) );
  XNOR2_X1 U15932 ( .A(n4606), .B(n21080), .ZN(n21681) );
  XNOR2_X1 U15933 ( .A(n21139), .B(n23718), .ZN(n4606) );
  OAI211_X1 U15935 ( .C1(n2616), .C2(n40910), .A(n40274), .B(n40275), .ZN(
        n40277) );
  NAND2_X1 U15936 ( .A1(n9546), .A2(n357), .ZN(n4608) );
  NAND2_X1 U15937 ( .A1(n15264), .A2(n14784), .ZN(n4611) );
  AND2_X1 U15938 ( .A1(n24367), .A2(n6117), .ZN(n4972) );
  INV_X1 U15939 ( .A(n14488), .ZN(n14495) );
  INV_X1 U15940 ( .A(n17065), .ZN(n19078) );
  NAND2_X1 U15941 ( .A1(n46796), .A2(n46797), .ZN(n4625) );
  INV_X1 U15942 ( .A(n30393), .ZN(n5300) );
  INV_X1 U15943 ( .A(n34240), .ZN(n34402) );
  XNOR2_X1 U15944 ( .A(n34402), .B(n2410), .ZN(n33890) );
  NOR2_X1 U15945 ( .A1(n6111), .A2(n8648), .ZN(n6110) );
  XNOR2_X2 U15947 ( .A(n24647), .B(n24648), .ZN(n27711) );
  XNOR2_X1 U15948 ( .A(n4614), .B(n24456), .ZN(n24463) );
  NAND2_X1 U15949 ( .A1(n9061), .A2(n4615), .ZN(n7562) );
  NAND3_X1 U15950 ( .A1(n10950), .A2(n12308), .A3(n4616), .ZN(n4615) );
  NOR2_X1 U15951 ( .A1(n2313), .A2(n4617), .ZN(n4616) );
  INV_X1 U15952 ( .A(n4620), .ZN(n4619) );
  OAI211_X1 U15953 ( .C1(n21955), .C2(n21956), .A(n21954), .B(n21967), .ZN(
        n4620) );
  OAI21_X1 U15954 ( .B1(n5269), .B2(n23178), .A(n4621), .ZN(n22792) );
  INV_X1 U15955 ( .A(n5289), .ZN(n4621) );
  NAND2_X1 U15956 ( .A1(n23171), .A2(n4622), .ZN(n5289) );
  NOR2_X1 U15957 ( .A1(n22674), .A2(n51021), .ZN(n4622) );
  XNOR2_X1 U15958 ( .A(n24465), .B(n5615), .ZN(n5614) );
  XNOR2_X1 U15959 ( .A(n5614), .B(n24735), .ZN(n6291) );
  XNOR2_X1 U15961 ( .A(n17363), .B(n2226), .ZN(n17367) );
  NAND2_X1 U15963 ( .A1(n10740), .A2(n9418), .ZN(n7363) );
  NAND3_X1 U15964 ( .A1(n41212), .A2(n41207), .A3(n41211), .ZN(n41203) );
  INV_X1 U15965 ( .A(n47519), .ZN(n5991) );
  NAND3_X2 U15966 ( .A1(n36290), .A2(n5675), .A3(n36289), .ZN(n43954) );
  NAND2_X1 U15967 ( .A1(n10354), .A2(n799), .ZN(n5105) );
  INV_X1 U15968 ( .A(n39336), .ZN(n39334) );
  NOR2_X1 U15969 ( .A1(n8689), .A2(n48156), .ZN(n48124) );
  NAND2_X1 U15970 ( .A1(n7548), .A2(n26488), .ZN(n26489) );
  NAND2_X1 U15971 ( .A1(n38640), .A2(n38262), .ZN(n38256) );
  NAND2_X1 U15973 ( .A1(n40617), .A2(n41975), .ZN(n41981) );
  OR2_X2 U15977 ( .A1(n11730), .A2(n11732), .ZN(n13856) );
  INV_X1 U15978 ( .A(n5695), .ZN(n5694) );
  XNOR2_X1 U15981 ( .A(n4630), .B(n4694), .ZN(Plaintext[167]) );
  NAND2_X1 U15982 ( .A1(n8499), .A2(n44129), .ZN(n4630) );
  NAND2_X1 U15983 ( .A1(n7025), .A2(n46732), .ZN(n7024) );
  NAND2_X1 U15984 ( .A1(n32489), .A2(n32491), .ZN(n32017) );
  NAND2_X1 U15985 ( .A1(n4631), .A2(n48885), .ZN(n14901) );
  NAND2_X1 U15986 ( .A1(n8412), .A2(n14892), .ZN(n4631) );
  NAND2_X1 U15987 ( .A1(n20123), .A2(n19050), .ZN(n16494) );
  NAND3_X1 U15988 ( .A1(n48373), .A2(n48371), .A3(n4632), .ZN(n48375) );
  NAND3_X2 U15989 ( .A1(n28728), .A2(n4633), .A3(n28727), .ZN(n35512) );
  NAND3_X1 U15990 ( .A1(n37929), .A2(n37930), .A3(n2474), .ZN(n37931) );
  OR2_X1 U15991 ( .A1(n29018), .A2(n51115), .ZN(n28008) );
  NAND3_X2 U15992 ( .A1(n28682), .A2(n28680), .A3(n28681), .ZN(n30854) );
  XOR2_X1 U15994 ( .A(n25153), .B(n24276), .Z(n8385) );
  INV_X1 U15995 ( .A(Ciphertext[162]), .ZN(n7775) );
  INV_X1 U15996 ( .A(n31584), .ZN(n31634) );
  NAND3_X1 U15997 ( .A1(n10914), .A2(n10142), .A3(n10913), .ZN(n7864) );
  NAND2_X1 U15998 ( .A1(n19832), .A2(n21188), .ZN(n17194) );
  AND2_X1 U15999 ( .A1(n11236), .A2(n11235), .ZN(n11239) );
  INV_X1 U16001 ( .A(n4642), .ZN(n35937) );
  OAI211_X1 U16002 ( .C1(n35932), .C2(n35931), .A(n35929), .B(n35930), .ZN(
        n4642) );
  NAND2_X1 U16003 ( .A1(n12619), .A2(n10465), .ZN(n12637) );
  NAND2_X1 U16004 ( .A1(n19603), .A2(n19403), .ZN(n19436) );
  INV_X1 U16006 ( .A(n9213), .ZN(n7151) );
  XNOR2_X1 U16007 ( .A(n4643), .B(n25543), .ZN(n25547) );
  XNOR2_X1 U16008 ( .A(n25544), .B(n25542), .ZN(n4643) );
  XNOR2_X1 U16009 ( .A(n4644), .B(n36939), .ZN(n33575) );
  XNOR2_X1 U16010 ( .A(n33572), .B(n7550), .ZN(n4644) );
  NAND2_X1 U16011 ( .A1(n10192), .A2(n11015), .ZN(n9032) );
  OAI21_X1 U16013 ( .B1(n5933), .B2(n6938), .A(n7636), .ZN(n4646) );
  NAND2_X1 U16015 ( .A1(n7733), .A2(n15357), .ZN(n14486) );
  XNOR2_X1 U16016 ( .A(n18581), .B(n16590), .ZN(n4648) );
  INV_X1 U16018 ( .A(n51344), .ZN(n46755) );
  INV_X1 U16019 ( .A(n12359), .ZN(n10987) );
  INV_X1 U16022 ( .A(n22742), .ZN(n22297) );
  INV_X1 U16024 ( .A(n19800), .ZN(n21305) );
  XNOR2_X1 U16025 ( .A(n18139), .B(n15609), .ZN(n16937) );
  INV_X1 U16026 ( .A(n36606), .ZN(n36064) );
  INV_X1 U16027 ( .A(n42109), .ZN(n43667) );
  INV_X1 U16029 ( .A(n11488), .ZN(n11487) );
  NAND2_X1 U16031 ( .A1(n45877), .A2(n47795), .ZN(n47782) );
  AND4_X2 U16032 ( .A1(n45005), .A2(n45006), .A3(n48212), .A4(n45004), .ZN(
        n47795) );
  XNOR2_X1 U16033 ( .A(n18543), .B(n2429), .ZN(n17326) );
  XNOR2_X1 U16034 ( .A(n44085), .B(n41759), .ZN(n5362) );
  NAND2_X1 U16035 ( .A1(n21424), .A2(n21427), .ZN(n20840) );
  NAND3_X1 U16036 ( .A1(n12243), .A2(n12260), .A3(n12258), .ZN(n11338) );
  NAND3_X1 U16037 ( .A1(n36474), .A2(n36490), .A3(n36488), .ZN(n34640) );
  INV_X1 U16038 ( .A(n29032), .ZN(n26626) );
  NAND2_X1 U16039 ( .A1(n28160), .A2(n29032), .ZN(n28536) );
  INV_X1 U16042 ( .A(n11340), .ZN(n7284) );
  XOR2_X1 U16043 ( .A(n44903), .B(n43660), .Z(n7578) );
  INV_X1 U16044 ( .A(n14599), .ZN(n8039) );
  NAND3_X1 U16045 ( .A1(n44845), .A2(n51317), .A3(n46699), .ZN(n44836) );
  NAND2_X1 U16046 ( .A1(n18967), .A2(n19089), .ZN(n4656) );
  NAND2_X1 U16047 ( .A1(n21731), .A2(n22260), .ZN(n20863) );
  INV_X1 U16050 ( .A(n10046), .ZN(n10044) );
  NAND4_X4 U16051 ( .A1(n2232), .A2(n8078), .A3(n18241), .A4(n18242), .ZN(
        n22832) );
  INV_X1 U16054 ( .A(n47179), .ZN(n50774) );
  NAND2_X1 U16055 ( .A1(n50808), .A2(n51730), .ZN(n47179) );
  INV_X1 U16056 ( .A(n21578), .ZN(n5953) );
  XOR2_X1 U16057 ( .A(n16732), .B(n15467), .Z(n5672) );
  AOI22_X1 U16058 ( .A1(n32922), .A2(n5976), .B1(n4660), .B2(n32916), .ZN(
        n28826) );
  OAI21_X1 U16059 ( .B1(n31603), .B2(n32634), .A(n28812), .ZN(n4660) );
  NAND2_X1 U16060 ( .A1(n22765), .A2(n25064), .ZN(n5723) );
  OAI21_X1 U16061 ( .B1(n21025), .B2(n21931), .A(n21024), .ZN(n21029) );
  NAND2_X1 U16062 ( .A1(n19565), .A2(n22145), .ZN(n21024) );
  NAND3_X1 U16063 ( .A1(n4661), .A2(n327), .A3(n30105), .ZN(n30114) );
  OAI21_X1 U16064 ( .B1(n30103), .B2(n31502), .A(n31497), .ZN(n4661) );
  INV_X1 U16065 ( .A(n41274), .ZN(n7217) );
  INV_X1 U16067 ( .A(n4663), .ZN(n4662) );
  OAI211_X1 U16068 ( .C1(n7876), .C2(n3685), .A(n19805), .B(n7873), .ZN(n4663)
         );
  NOR2_X1 U16069 ( .A1(n14160), .A2(n14159), .ZN(n13763) );
  NAND3_X1 U16070 ( .A1(n30288), .A2(n30286), .A3(n30287), .ZN(n4664) );
  NAND2_X1 U16071 ( .A1(n10008), .A2(n580), .ZN(n10002) );
  NAND3_X1 U16072 ( .A1(n27627), .A2(n26890), .A3(n27618), .ZN(n26800) );
  NAND2_X2 U16073 ( .A1(n17544), .A2(n772), .ZN(n18342) );
  INV_X1 U16074 ( .A(n14368), .ZN(n4794) );
  NOR2_X1 U16075 ( .A1(n21285), .A2(n8446), .ZN(n8445) );
  XOR2_X1 U16076 ( .A(n15148), .B(n15147), .Z(n8118) );
  NAND3_X1 U16077 ( .A1(n21145), .A2(n22263), .A3(n21744), .ZN(n23329) );
  NAND4_X2 U16079 ( .A1(n23347), .A2(n23349), .A3(n23346), .A4(n23348), .ZN(
        n28430) );
  INV_X1 U16081 ( .A(n11033), .ZN(n8641) );
  OAI211_X1 U16082 ( .C1(n3876), .C2(n23182), .A(n22058), .B(n23171), .ZN(
        n7937) );
  OAI22_X1 U16083 ( .A1(n29716), .A2(n29715), .B1(n29714), .B2(n51108), .ZN(
        n29717) );
  NAND3_X1 U16084 ( .A1(n780), .A2(n15103), .A3(n15104), .ZN(n4669) );
  NAND2_X1 U16085 ( .A1(n12504), .A2(n51709), .ZN(n8154) );
  NAND2_X1 U16086 ( .A1(n24413), .A2(n23129), .ZN(n24123) );
  NAND2_X1 U16087 ( .A1(n10566), .A2(n11650), .ZN(n9511) );
  NAND2_X1 U16088 ( .A1(n26630), .A2(n26631), .ZN(n26632) );
  OAI21_X1 U16089 ( .B1(n23786), .B2(n4670), .A(n24246), .ZN(n21812) );
  NAND2_X1 U16090 ( .A1(n21823), .A2(n24245), .ZN(n4670) );
  NAND2_X1 U16091 ( .A1(n6654), .A2(n42018), .ZN(n42008) );
  NAND2_X1 U16092 ( .A1(n4672), .A2(n4671), .ZN(n21805) );
  NAND2_X1 U16093 ( .A1(n21791), .A2(n23827), .ZN(n4672) );
  NAND2_X2 U16095 ( .A1(n2336), .A2(n6889), .ZN(n47745) );
  OAI21_X1 U16096 ( .B1(n29767), .B2(n29064), .A(n30343), .ZN(n4673) );
  INV_X1 U16097 ( .A(n25106), .ZN(n29234) );
  NAND3_X1 U16098 ( .A1(n47782), .A2(n47730), .A3(n45877), .ZN(n45878) );
  INV_X1 U16099 ( .A(n47341), .ZN(n5237) );
  INV_X1 U16100 ( .A(n6356), .ZN(n6357) );
  INV_X1 U16101 ( .A(n20508), .ZN(n8001) );
  NAND4_X2 U16102 ( .A1(n11194), .A2(n11196), .A3(n11197), .A4(n11195), .ZN(
        n14070) );
  INV_X1 U16103 ( .A(n17747), .ZN(n5716) );
  NAND4_X1 U16106 ( .A1(n4677), .A2(n45973), .A3(n45971), .A4(n45972), .ZN(
        n45974) );
  NAND2_X1 U16107 ( .A1(n10221), .A2(n8839), .ZN(n10223) );
  NAND2_X1 U16108 ( .A1(n13846), .A2(n13847), .ZN(n13861) );
  XNOR2_X1 U16109 ( .A(n4678), .B(n17351), .ZN(n17114) );
  XNOR2_X1 U16110 ( .A(n17111), .B(n17112), .ZN(n4678) );
  NAND4_X2 U16111 ( .A1(n4679), .A2(n26326), .A3(n8209), .A4(n27901), .ZN(
        n31712) );
  OAI21_X1 U16112 ( .B1(n9772), .B2(n10296), .A(n9770), .ZN(n9653) );
  NAND2_X1 U16113 ( .A1(n10939), .A2(n9758), .ZN(n9770) );
  NAND4_X2 U16114 ( .A1(n4680), .A2(n7859), .A3(n20226), .A4(n7854), .ZN(
        n24237) );
  NAND4_X2 U16116 ( .A1(n20885), .A2(n20884), .A3(n20883), .A4(n20882), .ZN(
        n25946) );
  NOR2_X2 U16117 ( .A1(n44456), .A2(n44457), .ZN(n44468) );
  NOR2_X1 U16118 ( .A1(n5457), .A2(n5456), .ZN(n5455) );
  OAI211_X1 U16119 ( .C1(n38620), .C2(n38619), .A(n38616), .B(n38615), .ZN(
        n5487) );
  NAND3_X1 U16120 ( .A1(n13169), .A2(n13167), .A3(n13168), .ZN(n13183) );
  NAND3_X1 U16121 ( .A1(n10531), .A2(n10513), .A3(n10508), .ZN(n10032) );
  NAND2_X1 U16122 ( .A1(n41703), .A2(n4682), .ZN(n39872) );
  INV_X1 U16123 ( .A(n13184), .ZN(n4686) );
  XNOR2_X2 U16124 ( .A(n43272), .B(n44394), .ZN(n45344) );
  AOI22_X1 U16125 ( .A1(n38837), .A2(n6374), .B1(n52073), .B2(n38827), .ZN(
        n6373) );
  NAND2_X1 U16126 ( .A1(n7368), .A2(n29186), .ZN(n27929) );
  NAND3_X1 U16127 ( .A1(n42015), .A2(n42021), .A3(n41589), .ZN(n41584) );
  XNOR2_X1 U16128 ( .A(n25608), .B(n4688), .ZN(n24926) );
  NAND2_X1 U16133 ( .A1(n39394), .A2(n4693), .ZN(n37732) );
  INV_X1 U16134 ( .A(n29203), .ZN(n27888) );
  NAND2_X1 U16135 ( .A1(n9636), .A2(n11379), .ZN(n11365) );
  NAND2_X2 U16137 ( .A1(n4695), .A2(n29890), .ZN(n32438) );
  INV_X1 U16138 ( .A(n17619), .ZN(n18088) );
  NOR2_X1 U16139 ( .A1(n40528), .A2(n40539), .ZN(n5594) );
  NAND3_X1 U16140 ( .A1(n11025), .A2(n10578), .A3(n10000), .ZN(n10577) );
  NAND3_X1 U16141 ( .A1(n27938), .A2(n29263), .A3(n51114), .ZN(n30230) );
  NOR2_X1 U16142 ( .A1(n4699), .A2(n4698), .ZN(n8473) );
  NOR2_X1 U16143 ( .A1(n46407), .A2(n46193), .ZN(n4699) );
  NAND2_X1 U16145 ( .A1(n16842), .A2(n19389), .ZN(n4701) );
  NAND3_X2 U16146 ( .A1(n32927), .A2(n4702), .A3(n32924), .ZN(n33702) );
  INV_X1 U16147 ( .A(n12202), .ZN(n13017) );
  XNOR2_X1 U16149 ( .A(n42720), .B(n44397), .ZN(n4704) );
  OAI21_X1 U16150 ( .B1(n38684), .B2(n37944), .A(n37943), .ZN(n5265) );
  NAND4_X1 U16151 ( .A1(n7589), .A2(n9753), .A3(n9754), .A4(n7587), .ZN(n13229) );
  OR2_X2 U16152 ( .A1(n30952), .A2(n31109), .ZN(n35536) );
  NAND2_X1 U16153 ( .A1(n37539), .A2(n37551), .ZN(n37533) );
  NAND2_X1 U16154 ( .A1(n4709), .A2(n755), .ZN(n17011) );
  NOR2_X2 U16156 ( .A1(n32854), .A2(n32853), .ZN(n35761) );
  OAI21_X1 U16157 ( .B1(n31520), .B2(n31521), .A(n31519), .ZN(n4711) );
  INV_X1 U16158 ( .A(n32848), .ZN(n32839) );
  INV_X1 U16160 ( .A(n21632), .ZN(n21617) );
  NAND2_X1 U16161 ( .A1(n38762), .A2(n38761), .ZN(n5893) );
  XNOR2_X1 U16162 ( .A(n4713), .B(n16645), .ZN(n8408) );
  XNOR2_X1 U16163 ( .A(n16651), .B(n16652), .ZN(n4713) );
  NAND2_X1 U16164 ( .A1(n21082), .A2(n755), .ZN(n24296) );
  NOR2_X1 U16165 ( .A1(n23504), .A2(n24290), .ZN(n21082) );
  NAND2_X1 U16166 ( .A1(n29251), .A2(n28662), .ZN(n30223) );
  NAND2_X1 U16169 ( .A1(n9859), .A2(n10962), .ZN(n10051) );
  NAND3_X1 U16171 ( .A1(n31032), .A2(n31031), .A3(n31830), .ZN(n31049) );
  NAND3_X1 U16172 ( .A1(n4715), .A2(n31816), .A3(n31821), .ZN(n31029) );
  XNOR2_X1 U16173 ( .A(n4716), .B(n28215), .ZN(n28217) );
  XNOR2_X1 U16174 ( .A(n28216), .B(n28214), .ZN(n4716) );
  AOI21_X1 U16175 ( .B1(n7294), .B2(n18060), .A(n18327), .ZN(n7752) );
  OAI21_X1 U16178 ( .B1(n5244), .B2(n5243), .A(n19529), .ZN(n19706) );
  INV_X1 U16179 ( .A(Ciphertext[76]), .ZN(n5623) );
  OAI21_X1 U16180 ( .B1(n6819), .B2(n21470), .A(n52146), .ZN(n20498) );
  INV_X1 U16181 ( .A(n13646), .ZN(n14631) );
  INV_X1 U16182 ( .A(n29568), .ZN(n5267) );
  AOI21_X1 U16184 ( .B1(n23764), .B2(n23765), .A(n4722), .ZN(n23769) );
  NOR2_X1 U16185 ( .A1(n44869), .A2(n44870), .ZN(n45766) );
  NAND2_X1 U16186 ( .A1(n46633), .A2(n44864), .ZN(n44869) );
  INV_X1 U16187 ( .A(n40951), .ZN(n6741) );
  INV_X1 U16188 ( .A(n23937), .ZN(n5955) );
  INV_X1 U16189 ( .A(n32622), .ZN(n31562) );
  NAND2_X1 U16190 ( .A1(n22830), .A2(n22492), .ZN(n22822) );
  XNOR2_X1 U16191 ( .A(n2155), .B(n37252), .ZN(n31575) );
  INV_X1 U16192 ( .A(n30233), .ZN(n4724) );
  NOR2_X1 U16193 ( .A1(n22310), .A2(n22311), .ZN(n6822) );
  XNOR2_X1 U16194 ( .A(n15876), .B(n15454), .ZN(n17694) );
  OAI21_X1 U16195 ( .B1(n8574), .B2(n8573), .A(n19797), .ZN(n8572) );
  NAND4_X2 U16196 ( .A1(n20521), .A2(n20520), .A3(n20519), .A4(n20518), .ZN(
        n22470) );
  XNOR2_X1 U16198 ( .A(n8248), .B(n33504), .ZN(n8247) );
  XOR2_X1 U16199 ( .A(n46118), .B(n43721), .Z(n8669) );
  XNOR2_X1 U16200 ( .A(n5318), .B(n39822), .ZN(n41325) );
  OR2_X1 U16201 ( .A1(n11137), .A2(n52140), .ZN(n9259) );
  AND3_X1 U16202 ( .A1(n31695), .A2(n31698), .A3(n31696), .ZN(n8086) );
  NAND2_X2 U16203 ( .A1(n36238), .A2(n36237), .ZN(n42061) );
  NOR2_X1 U16204 ( .A1(n37416), .A2(n38468), .ZN(n38110) );
  INV_X1 U16205 ( .A(n33686), .ZN(n34622) );
  NAND4_X1 U16206 ( .A1(n41493), .A2(n41492), .A3(n41491), .A4(n41490), .ZN(
        n42778) );
  INV_X1 U16207 ( .A(n29410), .ZN(n27717) );
  AOI21_X1 U16208 ( .B1(n44618), .B2(n47294), .A(n44617), .ZN(n44619) );
  NAND2_X2 U16209 ( .A1(n4728), .A2(n2430), .ZN(n30983) );
  XNOR2_X1 U16210 ( .A(n35120), .B(n35118), .ZN(n4729) );
  OAI21_X1 U16211 ( .B1(n30070), .B2(n31104), .A(n4730), .ZN(n30075) );
  NAND2_X1 U16212 ( .A1(n4732), .A2(n4731), .ZN(n7866) );
  NAND2_X1 U16213 ( .A1(n45183), .A2(n45799), .ZN(n4731) );
  NAND2_X1 U16214 ( .A1(n46735), .A2(n46738), .ZN(n4732) );
  NAND2_X1 U16215 ( .A1(n9708), .A2(n9709), .ZN(n9720) );
  INV_X1 U16216 ( .A(n7957), .ZN(n7658) );
  NOR2_X1 U16217 ( .A1(n7481), .A2(n7480), .ZN(n7479) );
  OAI21_X1 U16218 ( .B1(n41680), .B2(n41684), .A(n41679), .ZN(n41682) );
  NAND2_X1 U16222 ( .A1(n19720), .A2(n19794), .ZN(n4735) );
  NAND2_X1 U16223 ( .A1(n19719), .A2(n19718), .ZN(n4736) );
  NAND4_X2 U16224 ( .A1(n13672), .A2(n13675), .A3(n13673), .A4(n13674), .ZN(
        n17234) );
  NAND2_X1 U16225 ( .A1(n20067), .A2(n20075), .ZN(n19132) );
  NAND2_X1 U16226 ( .A1(n31171), .A2(n31546), .ZN(n32661) );
  NAND2_X1 U16228 ( .A1(n31033), .A2(n30846), .ZN(n6105) );
  NAND3_X1 U16229 ( .A1(n32251), .A2(n31778), .A3(n1037), .ZN(n31236) );
  INV_X1 U16230 ( .A(n49984), .ZN(n7639) );
  OAI21_X1 U16231 ( .B1(n38737), .B2(n38736), .A(n6150), .ZN(n6149) );
  NAND2_X1 U16233 ( .A1(n40387), .A2(n40386), .ZN(n4740) );
  OAI21_X1 U16234 ( .B1(n11874), .B2(n50997), .A(n7355), .ZN(n11871) );
  NAND2_X1 U16235 ( .A1(n28839), .A2(n29746), .ZN(n4741) );
  NAND4_X2 U16236 ( .A1(n32393), .A2(n32392), .A3(n32391), .A4(n32390), .ZN(
        n35829) );
  NAND2_X1 U16238 ( .A1(n38633), .A2(n2491), .ZN(n4742) );
  NAND2_X1 U16239 ( .A1(n38262), .A2(n38259), .ZN(n38633) );
  INV_X1 U16240 ( .A(n8469), .ZN(n7780) );
  OAI21_X1 U16241 ( .B1(n48207), .B2(n48206), .A(n4743), .ZN(n48209) );
  OAI21_X1 U16242 ( .B1(n48204), .B2(n48205), .A(n48203), .ZN(n4743) );
  NAND2_X1 U16243 ( .A1(n47979), .A2(n47965), .ZN(n47927) );
  NAND2_X1 U16244 ( .A1(n40296), .A2(n40297), .ZN(n40298) );
  NAND2_X1 U16245 ( .A1(n4745), .A2(n37364), .ZN(n35453) );
  NAND2_X1 U16246 ( .A1(n35451), .A2(n35452), .ZN(n4745) );
  XOR2_X1 U16247 ( .A(n33761), .B(n34737), .Z(n6680) );
  NAND3_X2 U16248 ( .A1(n7353), .A2(n4922), .A3(n7352), .ZN(n28257) );
  XNOR2_X2 U16251 ( .A(n2196), .B(n46068), .ZN(n43522) );
  NAND2_X1 U16254 ( .A1(n37469), .A2(n6199), .ZN(n39654) );
  INV_X1 U16255 ( .A(n5813), .ZN(n20023) );
  NOR2_X1 U16256 ( .A1(n42053), .A2(n8758), .ZN(n5943) );
  INV_X1 U16257 ( .A(n10231), .ZN(n10230) );
  NAND2_X1 U16258 ( .A1(n12291), .A2(n12280), .ZN(n10231) );
  NAND2_X1 U16259 ( .A1(n13117), .A2(n13125), .ZN(n10776) );
  NAND2_X1 U16260 ( .A1(n14160), .A2(n14164), .ZN(n13125) );
  NAND2_X1 U16261 ( .A1(n22736), .A2(n22741), .ZN(n22738) );
  INV_X1 U16262 ( .A(n15617), .ZN(n6563) );
  NAND2_X1 U16263 ( .A1(n652), .A2(n49923), .ZN(n46175) );
  OAI21_X1 U16265 ( .B1(n28000), .B2(n28903), .A(n4751), .ZN(n26477) );
  OAI21_X1 U16267 ( .B1(n6704), .B2(n45993), .A(n45992), .ZN(n7564) );
  NAND2_X1 U16268 ( .A1(n4756), .A2(n49650), .ZN(n7167) );
  OAI21_X1 U16269 ( .B1(n4870), .B2(n50021), .A(n49659), .ZN(n4756) );
  NAND3_X1 U16270 ( .A1(n9944), .A2(n9507), .A3(n4757), .ZN(n9946) );
  NAND2_X1 U16272 ( .A1(n42152), .A2(n42144), .ZN(n4764) );
  NAND2_X1 U16273 ( .A1(n2846), .A2(n22333), .ZN(n4766) );
  INV_X1 U16274 ( .A(n24283), .ZN(n7247) );
  XNOR2_X2 U16275 ( .A(n5108), .B(n43596), .ZN(n45325) );
  XNOR2_X1 U16276 ( .A(n45320), .B(n43658), .ZN(n4767) );
  INV_X1 U16277 ( .A(n7827), .ZN(n6169) );
  NOR2_X1 U16278 ( .A1(n19409), .A2(n5558), .ZN(n5557) );
  NAND3_X2 U16281 ( .A1(n30056), .A2(n30055), .A3(n4769), .ZN(n37108) );
  NAND3_X1 U16282 ( .A1(n4772), .A2(n34634), .A3(n34633), .ZN(n34635) );
  NAND3_X1 U16283 ( .A1(n36396), .A2(n36410), .A3(n37640), .ZN(n4772) );
  XNOR2_X2 U16284 ( .A(n41523), .B(n41522), .ZN(n46730) );
  NAND2_X1 U16285 ( .A1(n11355), .A2(n12383), .ZN(n4773) );
  NAND2_X1 U16286 ( .A1(n4774), .A2(n28700), .ZN(n6800) );
  OAI22_X1 U16287 ( .A1(n5469), .A2(n29309), .B1(n26649), .B2(n29291), .ZN(
        n4774) );
  NAND3_X1 U16288 ( .A1(n46612), .A2(n46613), .A3(n51513), .ZN(n46617) );
  NAND2_X1 U16289 ( .A1(n4776), .A2(n40213), .ZN(n40211) );
  NOR2_X1 U16290 ( .A1(n331), .A2(n41231), .ZN(n4776) );
  XNOR2_X1 U16292 ( .A(n16909), .B(n16898), .ZN(n8513) );
  OAI211_X1 U16293 ( .C1(n5650), .C2(n14107), .A(n14434), .B(n14106), .ZN(
        n14108) );
  OAI21_X1 U16295 ( .B1(n47694), .B2(n47683), .A(n47667), .ZN(n4904) );
  OAI21_X1 U16296 ( .B1(n12110), .B2(n12109), .A(n4778), .ZN(n12119) );
  XNOR2_X1 U16297 ( .A(n4779), .B(n36856), .ZN(n37250) );
  XNOR2_X1 U16298 ( .A(n36865), .B(n35832), .ZN(n4779) );
  NAND2_X1 U16299 ( .A1(n11105), .A2(n10422), .ZN(n11961) );
  INV_X1 U16300 ( .A(n23535), .ZN(n23702) );
  AND2_X1 U16301 ( .A1(n8017), .A2(n50593), .ZN(n4941) );
  INV_X1 U16302 ( .A(n23477), .ZN(n20994) );
  INV_X1 U16304 ( .A(n47163), .ZN(n4780) );
  NAND2_X1 U16305 ( .A1(n46890), .A2(n45161), .ZN(n47163) );
  AND2_X1 U16306 ( .A1(n19035), .A2(n19034), .ZN(n6501) );
  AOI22_X1 U16307 ( .A1(n6069), .A2(n4794), .B1(n12983), .B2(n14553), .ZN(
        n6068) );
  INV_X1 U16308 ( .A(n50640), .ZN(n50611) );
  XNOR2_X1 U16309 ( .A(n42696), .B(n43352), .ZN(n43937) );
  INV_X1 U16310 ( .A(n6384), .ZN(n15162) );
  INV_X1 U16311 ( .A(n15338), .ZN(n15442) );
  INV_X1 U16312 ( .A(n8323), .ZN(n25991) );
  INV_X1 U16313 ( .A(n12464), .ZN(n8908) );
  AOI21_X1 U16315 ( .B1(n51699), .B2(n14826), .A(n15443), .ZN(n6039) );
  INV_X1 U16316 ( .A(n41354), .ZN(n6468) );
  NOR2_X1 U16317 ( .A1(n6432), .A2(n6431), .ZN(n6430) );
  INV_X1 U16318 ( .A(n21633), .ZN(n20692) );
  NOR2_X1 U16319 ( .A1(n2428), .A2(n5842), .ZN(n5841) );
  XNOR2_X1 U16320 ( .A(n18488), .B(n15744), .ZN(n15618) );
  XNOR2_X1 U16322 ( .A(n34079), .B(n34251), .ZN(n6293) );
  XNOR2_X1 U16323 ( .A(n33356), .B(n6143), .ZN(n6142) );
  XNOR2_X1 U16326 ( .A(n4783), .B(n44326), .ZN(n44341) );
  XNOR2_X1 U16327 ( .A(n44324), .B(n44325), .ZN(n4783) );
  NAND2_X1 U16328 ( .A1(n20013), .A2(n6952), .ZN(n17533) );
  NAND2_X1 U16329 ( .A1(n18294), .A2(n18288), .ZN(n20013) );
  INV_X1 U16332 ( .A(n40420), .ZN(n5324) );
  NAND4_X2 U16333 ( .A1(n4787), .A2(n46460), .A3(n336), .A4(n46461), .ZN(
        n48674) );
  NAND2_X1 U16334 ( .A1(n11460), .A2(n11634), .ZN(n9322) );
  NAND2_X1 U16335 ( .A1(n24412), .A2(n24409), .ZN(n21671) );
  AND4_X2 U16336 ( .A1(n21667), .A2(n21668), .A3(n21665), .A4(n21666), .ZN(
        n24409) );
  INV_X1 U16337 ( .A(n8069), .ZN(n8068) );
  OAI21_X1 U16339 ( .B1(n10571), .B2(n10570), .A(n7184), .ZN(n10573) );
  NAND2_X1 U16340 ( .A1(n6112), .A2(n29652), .ZN(n29402) );
  NAND2_X1 U16341 ( .A1(n47085), .A2(n46832), .ZN(n44467) );
  INV_X1 U16343 ( .A(n14059), .ZN(n14680) );
  NAND2_X1 U16344 ( .A1(n661), .A2(n46810), .ZN(n44458) );
  INV_X1 U16345 ( .A(n13458), .ZN(n15174) );
  XNOR2_X2 U16346 ( .A(n8930), .B(Key[156]), .ZN(n12545) );
  XNOR2_X1 U16347 ( .A(n16456), .B(n16455), .ZN(n16459) );
  XNOR2_X1 U16348 ( .A(n24086), .B(n25639), .ZN(n7074) );
  OAI21_X1 U16349 ( .B1(n684), .B2(n39751), .A(n39754), .ZN(n36508) );
  NAND2_X1 U16350 ( .A1(n39111), .A2(n38831), .ZN(n38837) );
  NAND2_X1 U16351 ( .A1(n45611), .A2(n48124), .ZN(n48162) );
  NAND3_X1 U16352 ( .A1(n5720), .A2(n5721), .A3(n33017), .ZN(n5719) );
  OAI22_X1 U16353 ( .A1(n12093), .A2(n12389), .B1(n12095), .B2(n12094), .ZN(
        n4790) );
  NAND2_X1 U16354 ( .A1(n19521), .A2(n6226), .ZN(n4791) );
  NAND3_X1 U16355 ( .A1(n4792), .A2(n13178), .A3(n13782), .ZN(n13181) );
  INV_X1 U16356 ( .A(n13177), .ZN(n4792) );
  NAND2_X1 U16357 ( .A1(n13161), .A2(n13170), .ZN(n13177) );
  XNOR2_X1 U16358 ( .A(n27240), .B(n26171), .ZN(n5386) );
  NAND2_X1 U16359 ( .A1(n9508), .A2(n11649), .ZN(n5658) );
  XNOR2_X1 U16360 ( .A(n51523), .B(n27309), .ZN(n24763) );
  XNOR2_X1 U16361 ( .A(n4795), .B(n49387), .ZN(Plaintext[107]) );
  AND3_X1 U16362 ( .A1(n49385), .A2(n49383), .A3(n49384), .ZN(n4796) );
  XNOR2_X1 U16363 ( .A(n4798), .B(n28056), .ZN(n28064) );
  XNOR2_X1 U16364 ( .A(n28062), .B(n28055), .ZN(n4798) );
  NAND2_X1 U16365 ( .A1(n4063), .A2(n21354), .ZN(n18724) );
  OR3_X1 U16366 ( .A1(n52094), .A2(n575), .A3(n39754), .ZN(n36505) );
  NAND2_X1 U16367 ( .A1(n23868), .A2(n4799), .ZN(n22613) );
  NAND3_X1 U16369 ( .A1(n5066), .A2(n5067), .A3(n7617), .ZN(n5065) );
  XNOR2_X1 U16371 ( .A(n28438), .B(n4801), .ZN(n28317) );
  NAND3_X1 U16372 ( .A1(n4804), .A2(n10318), .A3(n10317), .ZN(n10327) );
  NAND2_X1 U16373 ( .A1(n12079), .A2(n12635), .ZN(n4804) );
  INV_X1 U16374 ( .A(n13475), .ZN(n15054) );
  INV_X1 U16375 ( .A(n9210), .ZN(n6047) );
  NAND3_X1 U16376 ( .A1(n10604), .A2(n9915), .A3(n9914), .ZN(n9916) );
  NAND2_X1 U16377 ( .A1(n9380), .A2(n10665), .ZN(n9378) );
  NAND2_X1 U16378 ( .A1(n7019), .A2(n10662), .ZN(n9380) );
  NAND2_X1 U16380 ( .A1(n10607), .A2(n10065), .ZN(n10064) );
  AOI21_X1 U16381 ( .B1(n9878), .B2(n8528), .A(n8527), .ZN(n9924) );
  NAND3_X1 U16382 ( .A1(n2119), .A2(n48200), .A3(n45545), .ZN(n4808) );
  NAND2_X1 U16383 ( .A1(n52050), .A2(n52161), .ZN(n4809) );
  INV_X1 U16384 ( .A(n31996), .ZN(n31993) );
  NAND2_X1 U16385 ( .A1(n32509), .A2(n32503), .ZN(n31996) );
  INV_X1 U16386 ( .A(n17484), .ZN(n7956) );
  OAI21_X1 U16387 ( .B1(n11310), .B2(n12952), .A(n13627), .ZN(n7756) );
  NAND2_X1 U16388 ( .A1(n51736), .A2(n38704), .ZN(n38303) );
  NAND2_X1 U16389 ( .A1(n36123), .A2(n37448), .ZN(n36124) );
  NAND3_X2 U16390 ( .A1(n4810), .A2(n8982), .A3(n8980), .ZN(n18795) );
  NAND3_X1 U16391 ( .A1(n4811), .A2(n13703), .A3(n14257), .ZN(n13704) );
  INV_X1 U16392 ( .A(n14993), .ZN(n4811) );
  NAND2_X1 U16393 ( .A1(n4812), .A2(n43347), .ZN(n43348) );
  NAND3_X1 U16394 ( .A1(n43344), .A2(n43343), .A3(n4813), .ZN(n4812) );
  OAI21_X1 U16395 ( .B1(n22395), .B2(n22297), .A(n6376), .ZN(n19745) );
  NAND2_X1 U16396 ( .A1(n4815), .A2(n35305), .ZN(n35900) );
  NAND2_X1 U16397 ( .A1(n37680), .A2(n4816), .ZN(n4815) );
  NAND2_X1 U16398 ( .A1(n28852), .A2(n30340), .ZN(n28787) );
  NAND2_X1 U16399 ( .A1(n47122), .A2(n47128), .ZN(n47121) );
  NAND3_X1 U16401 ( .A1(n32091), .A2(n32092), .A3(n32090), .ZN(n32100) );
  AND2_X1 U16402 ( .A1(n21477), .A2(n21475), .ZN(n8395) );
  INV_X1 U16403 ( .A(n13778), .ZN(n7498) );
  NAND3_X2 U16404 ( .A1(n4925), .A2(n8189), .A3(n8188), .ZN(n33026) );
  INV_X1 U16405 ( .A(n22016), .ZN(n22008) );
  NAND2_X1 U16406 ( .A1(n22011), .A2(n21329), .ZN(n22016) );
  NAND3_X1 U16408 ( .A1(n47087), .A2(n7449), .A3(n7918), .ZN(n8523) );
  INV_X1 U16409 ( .A(n25680), .ZN(n28250) );
  NAND3_X1 U16410 ( .A1(n38686), .A2(n39271), .A3(n2513), .ZN(n38687) );
  NAND2_X2 U16411 ( .A1(n7390), .A2(n10238), .ZN(n14160) );
  OR2_X1 U16412 ( .A1(n27024), .A2(n29447), .ZN(n27028) );
  XNOR2_X1 U16413 ( .A(n16606), .B(n8729), .ZN(n16678) );
  INV_X1 U16414 ( .A(n39259), .ZN(n39282) );
  XNOR2_X1 U16415 ( .A(n17138), .B(n18522), .ZN(n15396) );
  BUF_X1 U16416 ( .A(Key[91]), .Z(n4818) );
  NOR2_X1 U16417 ( .A1(n12692), .A2(n12709), .ZN(n5298) );
  NAND3_X2 U16419 ( .A1(n36395), .A2(n36394), .A3(n36393), .ZN(n43950) );
  XNOR2_X2 U16420 ( .A(n15688), .B(n17786), .ZN(n18617) );
  NOR2_X1 U16421 ( .A1(n2457), .A2(n7526), .ZN(n7525) );
  NAND2_X1 U16422 ( .A1(n28548), .A2(n30283), .ZN(n27111) );
  XNOR2_X1 U16425 ( .A(n43349), .B(n8046), .ZN(n41893) );
  XNOR2_X1 U16426 ( .A(n25463), .B(n25462), .ZN(n6659) );
  INV_X1 U16427 ( .A(n40476), .ZN(n40470) );
  NAND3_X1 U16429 ( .A1(n19990), .A2(n21404), .A3(n21560), .ZN(n4825) );
  NAND2_X1 U16430 ( .A1(n41317), .A2(n41902), .ZN(n40726) );
  NAND2_X1 U16431 ( .A1(n6510), .A2(n13178), .ZN(n13786) );
  AND2_X2 U16432 ( .A1(n24570), .A2(n26804), .ZN(n26890) );
  INV_X1 U16433 ( .A(n13171), .ZN(n6511) );
  NAND3_X1 U16434 ( .A1(n30124), .A2(n30122), .A3(n30123), .ZN(n30130) );
  XNOR2_X1 U16435 ( .A(n35472), .B(n35473), .ZN(n4828) );
  INV_X1 U16436 ( .A(n17005), .ZN(n21900) );
  NAND2_X2 U16437 ( .A1(n52191), .A2(n38483), .ZN(n38468) );
  XNOR2_X1 U16438 ( .A(n4829), .B(n47924), .ZN(Plaintext[31]) );
  NAND4_X1 U16439 ( .A1(n47922), .A2(n47923), .A3(n47920), .A4(n47921), .ZN(
        n4829) );
  AND2_X1 U16440 ( .A1(n10558), .A2(n10559), .ZN(n7413) );
  OAI211_X1 U16441 ( .C1(n50804), .C2(n47187), .A(n50811), .B(n4830), .ZN(
        n47188) );
  NAND2_X1 U16442 ( .A1(n22481), .A2(n22479), .ZN(n22716) );
  NAND2_X1 U16443 ( .A1(n21527), .A2(n20611), .ZN(n18893) );
  NOR2_X2 U16444 ( .A1(n6903), .A2(n16125), .ZN(n20611) );
  INV_X1 U16445 ( .A(n43184), .ZN(n7216) );
  NAND2_X2 U16446 ( .A1(n5033), .A2(n35724), .ZN(n5032) );
  XNOR2_X1 U16447 ( .A(n45122), .B(n6012), .ZN(n45132) );
  XNOR2_X1 U16448 ( .A(n4833), .B(n36935), .ZN(n33415) );
  XNOR2_X1 U16449 ( .A(n35517), .B(n33411), .ZN(n4833) );
  NAND2_X1 U16450 ( .A1(n19806), .A2(n19801), .ZN(n18996) );
  NAND2_X1 U16451 ( .A1(n11921), .A2(n12612), .ZN(n12601) );
  NAND2_X1 U16453 ( .A1(n45904), .A2(n45905), .ZN(n4834) );
  NAND4_X2 U16455 ( .A1(n29969), .A2(n29971), .A3(n29972), .A4(n29970), .ZN(
        n5616) );
  NAND3_X2 U16457 ( .A1(n6877), .A2(n6878), .A3(n25979), .ZN(n31886) );
  NAND2_X1 U16458 ( .A1(n23314), .A2(n23306), .ZN(n22251) );
  INV_X1 U16459 ( .A(n12371), .ZN(n12369) );
  XNOR2_X1 U16460 ( .A(n25102), .B(n25103), .ZN(n6644) );
  OAI22_X1 U16461 ( .A1(n49016), .A2(n8131), .B1(n46310), .B2(n49019), .ZN(
        n8130) );
  XNOR2_X1 U16463 ( .A(n4839), .B(n50203), .ZN(Plaintext[147]) );
  NAND3_X1 U16464 ( .A1(n50202), .A2(n50200), .A3(n50201), .ZN(n4839) );
  OAI21_X1 U16467 ( .B1(n4842), .B2(n4841), .A(n50233), .ZN(n5798) );
  NAND2_X1 U16468 ( .A1(n5799), .A2(n50208), .ZN(n4841) );
  NAND3_X1 U16469 ( .A1(n37622), .A2(n2330), .A3(n4843), .ZN(n37626) );
  NAND2_X1 U16470 ( .A1(n37621), .A2(n37620), .ZN(n4843) );
  NAND2_X1 U16471 ( .A1(n29412), .A2(n4844), .ZN(n29414) );
  OR2_X1 U16472 ( .A1(n26731), .A2(n29413), .ZN(n4844) );
  XNOR2_X2 U16474 ( .A(n34460), .B(n34461), .ZN(n38270) );
  XNOR2_X2 U16476 ( .A(n43026), .B(n43025), .ZN(n50294) );
  NOR2_X1 U16477 ( .A1(n51635), .A2(n51691), .ZN(n7203) );
  NAND3_X1 U16478 ( .A1(n40817), .A2(n40815), .A3(n52151), .ZN(n6507) );
  XNOR2_X1 U16479 ( .A(n4846), .B(n34160), .ZN(n34162) );
  XNOR2_X1 U16480 ( .A(n34151), .B(n34152), .ZN(n4846) );
  INV_X1 U16481 ( .A(n39646), .ZN(n38842) );
  NAND2_X1 U16482 ( .A1(n40342), .A2(n39855), .ZN(n39646) );
  NOR2_X1 U16483 ( .A1(n11410), .A2(n438), .ZN(n10390) );
  XOR2_X1 U16484 ( .A(n28294), .B(n28293), .Z(n5313) );
  NAND4_X1 U16485 ( .A1(n49195), .A2(n46004), .A3(n46003), .A4(n6810), .ZN(
        n7565) );
  NOR2_X1 U16486 ( .A1(n34181), .A2(n36557), .ZN(n7434) );
  XNOR2_X1 U16487 ( .A(n40581), .B(n40524), .ZN(n7623) );
  NAND3_X1 U16488 ( .A1(n4849), .A2(n23570), .A3(n23350), .ZN(n6514) );
  NAND2_X1 U16490 ( .A1(n4851), .A2(n32409), .ZN(n4850) );
  OAI21_X1 U16491 ( .B1(n37888), .B2(n6088), .A(n6087), .ZN(n6086) );
  INV_X1 U16492 ( .A(n14596), .ZN(n8038) );
  XNOR2_X1 U16493 ( .A(n4852), .B(n34872), .ZN(n34874) );
  XNOR2_X1 U16494 ( .A(n34864), .B(n34863), .ZN(n4852) );
  NAND2_X1 U16495 ( .A1(n5669), .A2(n32301), .ZN(n30636) );
  NAND3_X2 U16496 ( .A1(n41558), .A2(n41560), .A3(n5533), .ZN(n44547) );
  INV_X1 U16498 ( .A(n41390), .ZN(n41542) );
  OAI211_X1 U16500 ( .C1(n15165), .C2(n15158), .A(n4853), .B(n15157), .ZN(
        n15160) );
  INV_X1 U16501 ( .A(n15159), .ZN(n4853) );
  INV_X1 U16502 ( .A(n14453), .ZN(n14442) );
  NAND3_X1 U16503 ( .A1(n40507), .A2(n40508), .A3(n4854), .ZN(n40509) );
  NAND3_X1 U16504 ( .A1(n40505), .A2(n40506), .A3(n41063), .ZN(n4854) );
  AND2_X1 U16505 ( .A1(n11349), .A2(n11336), .ZN(n7281) );
  AND2_X1 U16506 ( .A1(n29543), .A2(n27053), .ZN(n27703) );
  XNOR2_X1 U16507 ( .A(n43562), .B(n2371), .ZN(n43580) );
  INV_X1 U16508 ( .A(n34945), .ZN(n5153) );
  INV_X1 U16509 ( .A(n29545), .ZN(n27056) );
  AOI21_X1 U16510 ( .B1(n49924), .B2(n49925), .A(n5959), .ZN(n5958) );
  INV_X1 U16511 ( .A(n41395), .ZN(n40938) );
  BUF_X1 U16512 ( .A(Key[55]), .Z(n4855) );
  OAI21_X1 U16513 ( .B1(n7504), .B2(n50316), .A(n50328), .ZN(n7503) );
  NAND2_X1 U16514 ( .A1(n5278), .A2(n29686), .ZN(n31088) );
  NAND4_X2 U16515 ( .A1(n18116), .A2(n18115), .A3(n18114), .A4(n18113), .ZN(
        n22506) );
  XNOR2_X1 U16516 ( .A(n35283), .B(n36766), .ZN(n34305) );
  XNOR2_X1 U16517 ( .A(n26215), .B(n4856), .ZN(n26217) );
  XNOR2_X1 U16518 ( .A(n26213), .B(n26214), .ZN(n4856) );
  XNOR2_X1 U16519 ( .A(n4857), .B(n28401), .ZN(n28403) );
  XNOR2_X1 U16520 ( .A(n28399), .B(n28400), .ZN(n4857) );
  NAND2_X1 U16521 ( .A1(n22344), .A2(n27638), .ZN(n27728) );
  NAND4_X1 U16522 ( .A1(n4860), .A2(n22707), .A3(n22706), .A4(n22708), .ZN(
        n22727) );
  NAND4_X2 U16523 ( .A1(n40603), .A2(n7106), .A3(n40601), .A4(n40602), .ZN(
        n45284) );
  NAND2_X1 U16524 ( .A1(n40249), .A2(n4862), .ZN(n4861) );
  INV_X1 U16525 ( .A(n41291), .ZN(n5086) );
  NAND3_X2 U16527 ( .A1(n4863), .A2(n12392), .A3(n6710), .ZN(n14720) );
  NAND2_X1 U16528 ( .A1(n12374), .A2(n12373), .ZN(n4863) );
  INV_X1 U16529 ( .A(n13338), .ZN(n13337) );
  NAND2_X1 U16530 ( .A1(n15091), .A2(n2166), .ZN(n4867) );
  NAND3_X1 U16531 ( .A1(n35965), .A2(n35963), .A3(n35964), .ZN(n35970) );
  NOR2_X1 U16532 ( .A1(n31870), .A2(n28487), .ZN(n30125) );
  XNOR2_X1 U16533 ( .A(n18489), .B(n15901), .ZN(n19194) );
  INV_X1 U16535 ( .A(n30712), .ZN(n28801) );
  INV_X1 U16536 ( .A(n49647), .ZN(n4870) );
  NAND2_X1 U16537 ( .A1(n45957), .A2(n6116), .ZN(n49647) );
  XNOR2_X1 U16539 ( .A(n4872), .B(n48803), .ZN(Plaintext[74]) );
  NAND3_X1 U16540 ( .A1(n48802), .A2(n48800), .A3(n4873), .ZN(n4872) );
  NAND2_X1 U16541 ( .A1(n45749), .A2(n48808), .ZN(n48791) );
  AOI21_X1 U16542 ( .B1(n39012), .B2(n36780), .A(n36779), .ZN(n8462) );
  NAND2_X1 U16543 ( .A1(n35139), .A2(n38116), .ZN(n4875) );
  NAND2_X1 U16544 ( .A1(n39730), .A2(n41278), .ZN(n41028) );
  NOR2_X1 U16545 ( .A1(n40373), .A2(n41317), .ZN(n4876) );
  NAND2_X1 U16546 ( .A1(n28810), .A2(n30705), .ZN(n30717) );
  NAND3_X1 U16547 ( .A1(n50009), .A2(n50322), .A3(n47369), .ZN(n43578) );
  NAND2_X1 U16548 ( .A1(n50564), .A2(n50533), .ZN(n50497) );
  NAND4_X4 U16551 ( .A1(n28763), .A2(n28762), .A3(n5978), .A4(n5977), .ZN(
        n32909) );
  NAND3_X1 U16552 ( .A1(n48607), .A2(n48649), .A3(n51382), .ZN(n48603) );
  NAND2_X2 U16553 ( .A1(n5017), .A2(n41043), .ZN(n43102) );
  INV_X1 U16554 ( .A(n20416), .ZN(n7835) );
  XNOR2_X2 U16555 ( .A(n41820), .B(n44190), .ZN(n43197) );
  OAI211_X1 U16556 ( .C1(n786), .C2(n13436), .A(n4878), .B(n13435), .ZN(n13437) );
  NAND4_X1 U16557 ( .A1(n13431), .A2(n13994), .A3(n13432), .A4(n13433), .ZN(
        n4878) );
  OAI21_X1 U16558 ( .B1(n46969), .B2(n46984), .A(n50360), .ZN(n46973) );
  NAND2_X1 U16559 ( .A1(n48611), .A2(n48646), .ZN(n6806) );
  INV_X1 U16560 ( .A(n38815), .ZN(n38816) );
  NAND2_X1 U16561 ( .A1(n41792), .A2(n41800), .ZN(n38815) );
  XOR2_X1 U16562 ( .A(n28318), .B(n26516), .Z(n8627) );
  OAI211_X1 U16563 ( .C1(n6062), .C2(n41801), .A(n6061), .B(n5604), .ZN(n6060)
         );
  XOR2_X1 U16564 ( .A(n24530), .B(n28409), .Z(n8562) );
  NAND2_X1 U16565 ( .A1(n39710), .A2(n39711), .ZN(n39716) );
  NAND2_X1 U16566 ( .A1(n7011), .A2(n37545), .ZN(n37405) );
  NAND2_X1 U16567 ( .A1(n31116), .A2(n30073), .ZN(n29587) );
  NAND2_X1 U16568 ( .A1(n1497), .A2(n24237), .ZN(n20875) );
  NOR2_X2 U16571 ( .A1(n8367), .A2(n21620), .ZN(n21639) );
  NAND2_X1 U16573 ( .A1(n13765), .A2(n14159), .ZN(n7928) );
  OAI21_X1 U16574 ( .B1(n10287), .B2(n5776), .A(n12334), .ZN(n5927) );
  INV_X1 U16575 ( .A(n34087), .ZN(n8011) );
  INV_X1 U16577 ( .A(n15061), .ZN(n6294) );
  INV_X1 U16578 ( .A(n13659), .ZN(n14637) );
  NOR2_X1 U16579 ( .A1(n6559), .A2(n6558), .ZN(n6557) );
  NAND2_X1 U16580 ( .A1(n11999), .A2(n14394), .ZN(n11296) );
  INV_X1 U16581 ( .A(n45834), .ZN(n42175) );
  NAND2_X1 U16582 ( .A1(n45828), .A2(n42180), .ZN(n45834) );
  NAND4_X1 U16583 ( .A1(n48437), .A2(n48434), .A3(n48259), .A4(n48264), .ZN(
        n45587) );
  NAND4_X1 U16585 ( .A1(n11241), .A2(n11240), .A3(n11239), .A4(n11238), .ZN(
        n11293) );
  NOR2_X1 U16586 ( .A1(n11530), .A2(n11581), .ZN(n11508) );
  XNOR2_X2 U16588 ( .A(n37152), .B(n37151), .ZN(n38664) );
  NAND2_X1 U16589 ( .A1(n50297), .A2(n49637), .ZN(n49613) );
  XNOR2_X1 U16591 ( .A(n41306), .B(n41305), .ZN(n4888) );
  AOI21_X1 U16592 ( .B1(n4889), .B2(n975), .A(n22156), .ZN(n20954) );
  NAND2_X1 U16593 ( .A1(n20958), .A2(n22140), .ZN(n4889) );
  NAND3_X1 U16594 ( .A1(n14060), .A2(n15273), .A3(n14950), .ZN(n14061) );
  NAND4_X2 U16596 ( .A1(n20963), .A2(n20962), .A3(n20964), .A4(n21023), .ZN(
        n27419) );
  OAI211_X1 U16598 ( .C1(n37511), .C2(n37760), .A(n36250), .B(n36249), .ZN(
        n5940) );
  NOR2_X1 U16599 ( .A1(n20802), .A2(n20801), .ZN(n4891) );
  NAND2_X1 U16602 ( .A1(n754), .A2(n23955), .ZN(n20848) );
  NAND2_X1 U16603 ( .A1(n4893), .A2(n14576), .ZN(n7713) );
  NAND2_X1 U16604 ( .A1(n7714), .A2(n15178), .ZN(n4893) );
  NAND2_X1 U16605 ( .A1(n41233), .A2(n41232), .ZN(n4894) );
  INV_X1 U16606 ( .A(n41227), .ZN(n41229) );
  AND2_X1 U16608 ( .A1(n20565), .A2(n20564), .ZN(n20570) );
  AND2_X1 U16609 ( .A1(n38231), .A2(n38896), .ZN(n5431) );
  BUF_X1 U16610 ( .A(Key[33]), .Z(n4896) );
  OAI21_X1 U16612 ( .B1(n5138), .B2(n13063), .A(n13062), .ZN(n5137) );
  INV_X1 U16613 ( .A(n21605), .ZN(n21364) );
  INV_X1 U16614 ( .A(n14738), .ZN(n20383) );
  NOR2_X1 U16615 ( .A1(n18728), .A2(n8493), .ZN(n8492) );
  INV_X1 U16617 ( .A(n13057), .ZN(n14795) );
  INV_X1 U16618 ( .A(n9859), .ZN(n6005) );
  INV_X1 U16619 ( .A(n5312), .ZN(n38569) );
  INV_X1 U16620 ( .A(n40730), .ZN(n5318) );
  INV_X1 U16621 ( .A(n16834), .ZN(n5519) );
  INV_X1 U16622 ( .A(n28738), .ZN(n5199) );
  XNOR2_X1 U16623 ( .A(n33095), .B(n2309), .ZN(n7337) );
  OAI211_X1 U16624 ( .C1(n37731), .C2(n5520), .A(n37739), .B(n3735), .ZN(
        n37726) );
  OAI211_X1 U16625 ( .C1(n30629), .C2(n31747), .A(n5820), .B(n5819), .ZN(n5818) );
  XNOR2_X1 U16626 ( .A(n4898), .B(n18152), .ZN(n18167) );
  XNOR2_X1 U16627 ( .A(n18151), .B(n18150), .ZN(n4898) );
  XNOR2_X1 U16630 ( .A(n4900), .B(n43297), .ZN(n43299) );
  XNOR2_X1 U16631 ( .A(n43979), .B(n43296), .ZN(n4900) );
  XNOR2_X1 U16632 ( .A(n4901), .B(n8444), .ZN(n8442) );
  XNOR2_X1 U16633 ( .A(n23935), .B(n23936), .ZN(n4901) );
  XNOR2_X1 U16634 ( .A(n45376), .B(n4902), .ZN(n38400) );
  XNOR2_X1 U16635 ( .A(n37831), .B(n37832), .ZN(n4902) );
  AOI21_X1 U16637 ( .B1(n10272), .B2(n10991), .A(n9785), .ZN(n9021) );
  NAND2_X1 U16638 ( .A1(n4176), .A2(n10267), .ZN(n10991) );
  NAND2_X1 U16639 ( .A1(n4176), .A2(n9782), .ZN(n12352) );
  NAND2_X1 U16640 ( .A1(n6262), .A2(n36000), .ZN(n37644) );
  OR2_X2 U16641 ( .A1(n5684), .A2(n5938), .ZN(n49511) );
  NAND2_X1 U16642 ( .A1(n4903), .A2(n49343), .ZN(n49360) );
  OAI211_X1 U16643 ( .C1(n47664), .C2(n47668), .A(n4904), .B(n45887), .ZN(
        n45894) );
  INV_X1 U16645 ( .A(n31578), .ZN(n4906) );
  NAND3_X2 U16646 ( .A1(n37515), .A2(n37514), .A3(n5637), .ZN(n43327) );
  NAND2_X1 U16647 ( .A1(n18376), .A2(n20028), .ZN(n17046) );
  NAND2_X1 U16648 ( .A1(n51669), .A2(n14712), .ZN(n13343) );
  XNOR2_X1 U16649 ( .A(n26139), .B(n26138), .ZN(n26158) );
  NAND3_X1 U16650 ( .A1(n23472), .A2(n21957), .A3(n21945), .ZN(n23469) );
  NAND4_X1 U16651 ( .A1(n15325), .A2(n51700), .A3(n15324), .A4(n15437), .ZN(
        n15328) );
  XNOR2_X1 U16652 ( .A(n4910), .B(n26382), .ZN(n26383) );
  XNOR2_X1 U16653 ( .A(n26381), .B(n26380), .ZN(n4910) );
  NAND2_X1 U16655 ( .A1(n41621), .A2(n41693), .ZN(n41699) );
  NAND2_X1 U16656 ( .A1(n4912), .A2(n18727), .ZN(n18728) );
  INV_X1 U16657 ( .A(n22118), .ZN(n20972) );
  XNOR2_X1 U16658 ( .A(n4913), .B(n42452), .ZN(Plaintext[32]) );
  NAND2_X1 U16659 ( .A1(n46642), .A2(n44652), .ZN(n46631) );
  NAND2_X1 U16660 ( .A1(n14244), .A2(n14243), .ZN(n14256) );
  NAND3_X1 U16661 ( .A1(n4914), .A2(n39047), .A3(n41711), .ZN(n39048) );
  NAND2_X1 U16662 ( .A1(n39046), .A2(n41706), .ZN(n4914) );
  NAND2_X1 U16663 ( .A1(n11064), .A2(n11902), .ZN(n4915) );
  XNOR2_X2 U16664 ( .A(n32860), .B(n35333), .ZN(n37097) );
  NAND3_X2 U16666 ( .A1(n4917), .A2(n8895), .A3(n8894), .ZN(n14252) );
  OAI211_X1 U16667 ( .C1(n34321), .C2(n34322), .A(n34320), .B(n8607), .ZN(
        n34323) );
  NAND2_X1 U16668 ( .A1(n12470), .A2(n12488), .ZN(n11488) );
  NAND2_X1 U16670 ( .A1(n32401), .A2(n32066), .ZN(n32075) );
  NAND2_X1 U16671 ( .A1(n6378), .A2(n15377), .ZN(n15389) );
  INV_X1 U16672 ( .A(n10051), .ZN(n9862) );
  NAND2_X1 U16673 ( .A1(n4920), .A2(n6996), .ZN(n6108) );
  NAND2_X1 U16674 ( .A1(n37525), .A2(n37516), .ZN(n4920) );
  INV_X1 U16675 ( .A(n15358), .ZN(n7906) );
  XNOR2_X1 U16676 ( .A(n17336), .B(n17335), .ZN(n4921) );
  NAND2_X1 U16677 ( .A1(n5656), .A2(n29278), .ZN(n29183) );
  XNOR2_X2 U16678 ( .A(n25445), .B(n24976), .ZN(n25829) );
  XNOR2_X1 U16679 ( .A(n25441), .B(n4924), .ZN(n25453) );
  XNOR2_X1 U16680 ( .A(n25440), .B(n25443), .ZN(n4924) );
  NAND2_X1 U16681 ( .A1(n44001), .A2(n50259), .ZN(n47064) );
  NAND3_X2 U16682 ( .A1(n7265), .A2(n19825), .A3(n7266), .ZN(n25056) );
  NAND2_X1 U16683 ( .A1(n11322), .A2(n11329), .ZN(n11328) );
  NAND2_X1 U16684 ( .A1(n31533), .A2(n33030), .ZN(n33028) );
  NAND3_X1 U16685 ( .A1(n8584), .A2(n14966), .A3(n13124), .ZN(n4927) );
  NAND4_X4 U16686 ( .A1(n31390), .A2(n6422), .A3(n6419), .A4(n6418), .ZN(
        n37067) );
  NAND3_X2 U16687 ( .A1(n4929), .A2(n4928), .A3(n14196), .ZN(n17731) );
  INV_X1 U16688 ( .A(n31417), .ZN(n5634) );
  OAI21_X1 U16690 ( .B1(n20421), .B2(n20422), .A(n19330), .ZN(n4933) );
  NAND2_X1 U16692 ( .A1(n40617), .A2(n41647), .ZN(n41641) );
  NAND2_X1 U16693 ( .A1(n24191), .A2(n24188), .ZN(n23200) );
  NAND3_X1 U16694 ( .A1(n8306), .A2(n48093), .A3(n48094), .ZN(n8305) );
  NAND2_X1 U16695 ( .A1(n23036), .A2(n23035), .ZN(n4935) );
  NAND2_X1 U16696 ( .A1(n9120), .A2(n11095), .ZN(n9121) );
  NAND2_X1 U16697 ( .A1(n38687), .A2(n38688), .ZN(n38693) );
  XNOR2_X1 U16699 ( .A(n17253), .B(n15684), .ZN(n4938) );
  NOR2_X1 U16700 ( .A1(n41374), .A2(n41380), .ZN(n40242) );
  NAND3_X1 U16702 ( .A1(n4941), .A2(n50647), .A3(n50646), .ZN(n50649) );
  NAND4_X1 U16703 ( .A1(n4942), .A2(n12605), .A3(n12604), .A4(n1307), .ZN(
        n12606) );
  NAND3_X1 U16704 ( .A1(n12596), .A2(n11913), .A3(n4942), .ZN(n11918) );
  NAND2_X1 U16705 ( .A1(n12600), .A2(n3377), .ZN(n4942) );
  NAND2_X1 U16706 ( .A1(n683), .A2(n42006), .ZN(n42013) );
  NOR2_X1 U16707 ( .A1(n41587), .A2(n6654), .ZN(n41589) );
  INV_X1 U16708 ( .A(n42020), .ZN(n4943) );
  NAND3_X1 U16709 ( .A1(n42011), .A2(n6236), .A3(n3831), .ZN(n42012) );
  AOI21_X1 U16710 ( .B1(n41509), .B2(n3831), .A(n42014), .ZN(n40700) );
  NAND2_X1 U16711 ( .A1(n39493), .A2(n4944), .ZN(n39494) );
  NAND2_X1 U16712 ( .A1(n10069), .A2(n10607), .ZN(n10616) );
  NAND3_X1 U16713 ( .A1(n10069), .A2(n10607), .A3(n52185), .ZN(n10620) );
  OAI21_X1 U16715 ( .B1(n9921), .B2(n10618), .A(n10620), .ZN(n4945) );
  NAND4_X2 U16716 ( .A1(n29711), .A2(n29709), .A3(n29710), .A4(n29712), .ZN(
        n32724) );
  NAND2_X1 U16717 ( .A1(n39616), .A2(n51357), .ZN(n39577) );
  NAND2_X1 U16718 ( .A1(n21304), .A2(n19801), .ZN(n18999) );
  INV_X1 U16720 ( .A(n12799), .ZN(n12785) );
  NAND2_X1 U16721 ( .A1(n4949), .A2(n13449), .ZN(n12799) );
  NAND3_X2 U16722 ( .A1(n8177), .A2(n9925), .A3(n9924), .ZN(n13449) );
  NAND2_X1 U16723 ( .A1(n40549), .A2(n4950), .ZN(n4955) );
  INV_X1 U16726 ( .A(n40572), .ZN(n4951) );
  NAND2_X1 U16727 ( .A1(n4954), .A2(n40558), .ZN(n40555) );
  NAND3_X1 U16728 ( .A1(n4951), .A2(n4000), .A3(n4954), .ZN(n37464) );
  NAND2_X1 U16729 ( .A1(n40157), .A2(n4954), .ZN(n40311) );
  OAI211_X1 U16730 ( .C1(n40563), .C2(n4954), .A(n4952), .B(n40153), .ZN(
        n40155) );
  NAND3_X1 U16731 ( .A1(n40567), .A2(n40556), .A3(n4954), .ZN(n4952) );
  AND2_X1 U16732 ( .A1(n4954), .A2(n40549), .ZN(n4953) );
  NAND3_X1 U16733 ( .A1(n40319), .A2(n4955), .A3(n52160), .ZN(n39658) );
  NAND3_X1 U16736 ( .A1(n40496), .A2(n41057), .A3(n39129), .ZN(n35008) );
  NAND2_X1 U16739 ( .A1(n28715), .A2(n4965), .ZN(n27925) );
  NOR2_X1 U16740 ( .A1(n4966), .A2(n509), .ZN(n18989) );
  NAND2_X1 U16741 ( .A1(n3685), .A2(n18997), .ZN(n4966) );
  INV_X1 U16743 ( .A(n51716), .ZN(n4967) );
  NOR2_X1 U16744 ( .A1(n46869), .A2(n2159), .ZN(n47098) );
  NAND2_X1 U16746 ( .A1(n31039), .A2(n50986), .ZN(n30571) );
  OAI211_X1 U16747 ( .C1(n37963), .C2(n36548), .A(n3626), .B(n4968), .ZN(n4969) );
  NAND2_X1 U16748 ( .A1(n36542), .A2(n34090), .ZN(n4968) );
  INV_X1 U16749 ( .A(n36542), .ZN(n37963) );
  NAND2_X1 U16750 ( .A1(n23111), .A2(n30725), .ZN(n4970) );
  NAND3_X1 U16751 ( .A1(n28808), .A2(n30722), .A3(n30717), .ZN(n4971) );
  XNOR2_X2 U16752 ( .A(n35254), .B(n35833), .ZN(n34240) );
  NOR2_X1 U16754 ( .A1(n51127), .A2(n19892), .ZN(n19889) );
  XNOR2_X2 U16755 ( .A(n15586), .B(n4974), .ZN(n19892) );
  AND2_X1 U16756 ( .A1(n52147), .A2(n29110), .ZN(n25411) );
  INV_X1 U16757 ( .A(n12057), .ZN(n5687) );
  INV_X1 U16758 ( .A(n10662), .ZN(n10356) );
  NAND2_X1 U16759 ( .A1(n52211), .A2(n49656), .ZN(n45957) );
  NAND2_X1 U16760 ( .A1(n4978), .A2(n4976), .ZN(n38537) );
  NAND2_X1 U16761 ( .A1(n4977), .A2(n38512), .ZN(n4976) );
  NAND2_X1 U16762 ( .A1(n38531), .A2(n38530), .ZN(n4978) );
  XNOR2_X1 U16763 ( .A(n4979), .B(n16710), .ZN(n16713) );
  XNOR2_X1 U16764 ( .A(n4979), .B(n14591), .ZN(n14593) );
  XNOR2_X1 U16765 ( .A(n4979), .B(n18443), .ZN(n17108) );
  XNOR2_X1 U16766 ( .A(n4980), .B(n43495), .ZN(Plaintext[117]) );
  NAND3_X1 U16767 ( .A1(n43494), .A2(n4982), .A3(n4981), .ZN(n4980) );
  NAND2_X1 U16768 ( .A1(n338), .A2(n7209), .ZN(n4981) );
  NAND2_X1 U16769 ( .A1(n4984), .A2(n45021), .ZN(n4983) );
  XNOR2_X2 U16770 ( .A(n9072), .B(Key[29]), .ZN(n11611) );
  XNOR2_X2 U16771 ( .A(Key[153]), .B(Ciphertext[188]), .ZN(n11375) );
  NAND2_X1 U16772 ( .A1(n21339), .A2(n23489), .ZN(n4986) );
  NAND2_X1 U16773 ( .A1(n21339), .A2(n4985), .ZN(n8518) );
  NOR2_X1 U16774 ( .A1(n21977), .A2(n23485), .ZN(n4985) );
  INV_X1 U16775 ( .A(n23020), .ZN(n4987) );
  NAND2_X1 U16776 ( .A1(n4987), .A2(n21885), .ZN(n22862) );
  NAND2_X1 U16777 ( .A1(n19338), .A2(n8687), .ZN(n4989) );
  XNOR2_X1 U16778 ( .A(n4990), .B(n52138), .ZN(n37237) );
  XNOR2_X1 U16779 ( .A(n4990), .B(n34384), .ZN(n34386) );
  XNOR2_X1 U16780 ( .A(n4990), .B(n34020), .ZN(n34021) );
  XNOR2_X1 U16781 ( .A(n4990), .B(n33484), .ZN(n33485) );
  XNOR2_X2 U16782 ( .A(n36931), .B(n32801), .ZN(n4990) );
  NAND2_X1 U16783 ( .A1(n37189), .A2(n35407), .ZN(n4991) );
  XNOR2_X1 U16784 ( .A(n33813), .B(n33814), .ZN(n4995) );
  OAI22_X1 U16785 ( .A1(n4996), .A2(n46903), .B1(n44986), .B2(n46913), .ZN(
        n5023) );
  OAI21_X1 U16786 ( .B1(n603), .B2(n4996), .A(n46610), .ZN(n46611) );
  NAND2_X1 U16787 ( .A1(n45847), .A2(n4996), .ZN(n45849) );
  NAND2_X1 U16789 ( .A1(n5006), .A2(n2498), .ZN(n4999) );
  NAND4_X1 U16790 ( .A1(n5001), .A2(n29792), .A3(n28136), .A4(n28135), .ZN(
        n5932) );
  NAND2_X1 U16791 ( .A1(n5004), .A2(n13086), .ZN(n5003) );
  NAND2_X1 U16792 ( .A1(n12818), .A2(n13091), .ZN(n5004) );
  NOR2_X1 U16793 ( .A1(n30506), .A2(n32983), .ZN(n5935) );
  NAND2_X1 U16794 ( .A1(n712), .A2(n32590), .ZN(n32983) );
  NAND3_X1 U16795 ( .A1(n21892), .A2(n21890), .A3(n21891), .ZN(n5005) );
  OAI21_X1 U16796 ( .B1(n19397), .B2(n19396), .A(n19395), .ZN(n5007) );
  AOI21_X1 U16797 ( .B1(n17578), .B2(n17577), .A(n17576), .ZN(n19397) );
  NAND2_X1 U16798 ( .A1(n23857), .A2(n26912), .ZN(n5008) );
  NAND4_X2 U16799 ( .A1(n5009), .A2(n6640), .A3(n9800), .A4(n9802), .ZN(n5996)
         );
  XNOR2_X1 U16800 ( .A(n9803), .B(n557), .ZN(n10094) );
  XNOR2_X1 U16801 ( .A(n7339), .B(n44391), .ZN(n5011) );
  NAND2_X1 U16802 ( .A1(n5014), .A2(n5010), .ZN(n7339) );
  XNOR2_X1 U16803 ( .A(n46081), .B(n5011), .ZN(n41954) );
  NAND3_X1 U16804 ( .A1(n41043), .A2(n5017), .A3(n5016), .ZN(n5013) );
  NAND2_X1 U16805 ( .A1(n5015), .A2(n48064), .ZN(n5014) );
  OAI21_X1 U16806 ( .B1(n23140), .B2(n23139), .A(n23138), .ZN(n5019) );
  NAND2_X1 U16810 ( .A1(n46920), .A2(n46609), .ZN(n46604) );
  OAI21_X1 U16811 ( .B1(n46915), .B2(n44988), .A(n46919), .ZN(n5022) );
  XNOR2_X1 U16812 ( .A(n25747), .B(n26509), .ZN(n5024) );
  NAND3_X1 U16813 ( .A1(n5026), .A2(n30374), .A3(n30740), .ZN(n5030) );
  INV_X1 U16814 ( .A(n29884), .ZN(n5026) );
  NAND2_X1 U16815 ( .A1(n29779), .A2(n30733), .ZN(n5027) );
  NAND2_X2 U16816 ( .A1(n5031), .A2(n35698), .ZN(n40556) );
  XNOR2_X1 U16817 ( .A(n46113), .B(n5032), .ZN(n42730) );
  XNOR2_X1 U16818 ( .A(n44314), .B(n5032), .ZN(n42233) );
  XNOR2_X1 U16819 ( .A(n44240), .B(n5032), .ZN(n44241) );
  XNOR2_X1 U16820 ( .A(n46111), .B(n5032), .ZN(n42650) );
  XNOR2_X1 U16821 ( .A(n42358), .B(n5032), .ZN(n42359) );
  XNOR2_X1 U16822 ( .A(n42411), .B(n5032), .ZN(n42412) );
  NAND2_X1 U16824 ( .A1(n19447), .A2(n23987), .ZN(n23030) );
  NAND2_X1 U16825 ( .A1(n23032), .A2(n23983), .ZN(n5035) );
  INV_X1 U16827 ( .A(n35666), .ZN(n38165) );
  INV_X1 U16828 ( .A(n36122), .ZN(n5037) );
  NAND2_X1 U16829 ( .A1(n32615), .A2(n5040), .ZN(n32623) );
  NAND2_X1 U16830 ( .A1(n547), .A2(n29140), .ZN(n30160) );
  NAND2_X1 U16831 ( .A1(n39035), .A2(n51737), .ZN(n39439) );
  INV_X1 U16832 ( .A(n39452), .ZN(n39026) );
  INV_X1 U16833 ( .A(n39439), .ZN(n39437) );
  NAND2_X1 U16834 ( .A1(n39454), .A2(n5042), .ZN(n39041) );
  NAND2_X1 U16835 ( .A1(n39452), .A2(n39439), .ZN(n5042) );
  XNOR2_X1 U16837 ( .A(n5045), .B(n33857), .ZN(n33858) );
  XNOR2_X1 U16838 ( .A(n5045), .B(n5598), .ZN(n37294) );
  XNOR2_X1 U16839 ( .A(n5045), .B(n35537), .ZN(n36986) );
  NAND3_X2 U16840 ( .A1(n17022), .A2(n17023), .A3(n5046), .ZN(n23547) );
  INV_X1 U16841 ( .A(n17017), .ZN(n5046) );
  OAI211_X1 U16843 ( .C1(n28502), .C2(n28501), .A(n28500), .B(n5052), .ZN(
        n28516) );
  OAI211_X1 U16844 ( .C1(n29802), .C2(n28505), .A(n5053), .B(n28866), .ZN(
        n5052) );
  NAND2_X1 U16845 ( .A1(n5054), .A2(n29803), .ZN(n5053) );
  INV_X1 U16846 ( .A(n29796), .ZN(n5057) );
  NAND2_X1 U16848 ( .A1(n5061), .A2(n5060), .ZN(n5059) );
  NAND2_X1 U16849 ( .A1(n40662), .A2(n40661), .ZN(n5063) );
  NAND2_X1 U16850 ( .A1(n40662), .A2(n40032), .ZN(n5061) );
  NAND3_X1 U16852 ( .A1(n5065), .A2(n23089), .A3(n23088), .ZN(n7618) );
  INV_X1 U16853 ( .A(n23957), .ZN(n5069) );
  NAND2_X1 U16854 ( .A1(n5073), .A2(n40893), .ZN(n40280) );
  INV_X1 U16855 ( .A(n40893), .ZN(n40896) );
  NAND2_X1 U16856 ( .A1(n40893), .A2(n40274), .ZN(n5071) );
  INV_X1 U16858 ( .A(n40096), .ZN(n5076) );
  NAND2_X1 U16859 ( .A1(n48912), .A2(n48853), .ZN(n48886) );
  NAND4_X1 U16860 ( .A1(n7607), .A2(n48918), .A3(n5080), .A4(n5079), .ZN(n7606) );
  NAND4_X4 U16861 ( .A1(n5690), .A2(n5692), .A3(n5689), .A4(n5691), .ZN(n48919) );
  NAND2_X1 U16862 ( .A1(n5083), .A2(n16986), .ZN(n19640) );
  NAND2_X1 U16863 ( .A1(n45185), .A2(n46749), .ZN(n5084) );
  NAND2_X1 U16866 ( .A1(n41029), .A2(n41292), .ZN(n41291) );
  NAND2_X1 U16869 ( .A1(n50033), .A2(n5088), .ZN(n46160) );
  NOR2_X1 U16870 ( .A1(n50390), .A2(n5089), .ZN(n5088) );
  NAND4_X2 U16871 ( .A1(n5092), .A2(n41654), .A3(n41652), .A4(n5091), .ZN(
        n44510) );
  INV_X1 U16872 ( .A(n50976), .ZN(n5095) );
  OR2_X2 U16873 ( .A1(n19696), .A2(n19697), .ZN(n22390) );
  NAND4_X2 U16874 ( .A1(n11719), .A2(n11716), .A3(n11717), .A4(n11718), .ZN(
        n16036) );
  NAND2_X1 U16876 ( .A1(n2257), .A2(n20412), .ZN(n20373) );
  NAND2_X1 U16877 ( .A1(n11186), .A2(n7340), .ZN(n10859) );
  NAND2_X1 U16878 ( .A1(n13373), .A2(n5098), .ZN(n13374) );
  INV_X1 U16879 ( .A(n13371), .ZN(n5098) );
  OAI21_X1 U16882 ( .B1(n31709), .B2(n31712), .A(n5101), .ZN(n5100) );
  AOI21_X1 U16883 ( .B1(n31708), .B2(n31711), .A(n30814), .ZN(n5101) );
  NAND2_X1 U16884 ( .A1(n27852), .A2(n27858), .ZN(n26334) );
  OAI21_X1 U16886 ( .B1(n29487), .B2(n27852), .A(n29486), .ZN(n29491) );
  XNOR2_X1 U16887 ( .A(n33057), .B(n36754), .ZN(n33067) );
  INV_X1 U16888 ( .A(n33067), .ZN(n33062) );
  AND2_X1 U16889 ( .A1(n24000), .A2(n23992), .ZN(n22420) );
  NAND2_X1 U16890 ( .A1(n11389), .A2(n5107), .ZN(n5212) );
  NAND3_X1 U16891 ( .A1(n5106), .A2(n9221), .A3(n5104), .ZN(n9390) );
  NAND3_X1 U16892 ( .A1(n5105), .A2(n9388), .A3(n9389), .ZN(n5104) );
  NAND3_X1 U16893 ( .A1(n12051), .A2(n9389), .A3(n9388), .ZN(n5106) );
  XNOR2_X1 U16894 ( .A(n42715), .B(n51393), .ZN(n40979) );
  XNOR2_X1 U16895 ( .A(n51393), .B(n41924), .ZN(n41946) );
  XNOR2_X1 U16896 ( .A(n51393), .B(n44164), .ZN(n42501) );
  XNOR2_X1 U16897 ( .A(n51392), .B(n45327), .ZN(n42717) );
  XNOR2_X1 U16898 ( .A(n44074), .B(n51392), .ZN(n42554) );
  XNOR2_X1 U16899 ( .A(n44076), .B(n51392), .ZN(n44478) );
  INV_X1 U16900 ( .A(n32201), .ZN(n5110) );
  NAND2_X1 U16901 ( .A1(n5111), .A2(n32633), .ZN(n32917) );
  NAND3_X1 U16903 ( .A1(n32543), .A2(n32634), .A3(n5976), .ZN(n32544) );
  NOR2_X1 U16904 ( .A1(n14579), .A2(n15161), .ZN(n14572) );
  OAI21_X1 U16905 ( .B1(n51369), .B2(n5113), .A(n15177), .ZN(n13463) );
  NAND4_X1 U16906 ( .A1(n13458), .A2(n14579), .A3(n15163), .A4(n5113), .ZN(
        n13459) );
  NAND2_X1 U16907 ( .A1(n13457), .A2(n5112), .ZN(n10879) );
  OR2_X1 U16908 ( .A1(n14575), .A2(n5113), .ZN(n5112) );
  AND4_X4 U16909 ( .A1(n10824), .A2(n10823), .A3(n10822), .A4(n10821), .ZN(
        n15161) );
  NAND2_X1 U16910 ( .A1(n5116), .A2(n1230), .ZN(n5114) );
  NAND2_X1 U16911 ( .A1(n22429), .A2(n22430), .ZN(n22532) );
  NAND2_X1 U16912 ( .A1(n23032), .A2(n23036), .ZN(n5119) );
  AND2_X2 U16913 ( .A1(n12139), .A2(n438), .ZN(n5120) );
  NAND2_X1 U16914 ( .A1(n793), .A2(n5120), .ZN(n11418) );
  NAND2_X1 U16915 ( .A1(n8049), .A2(n5120), .ZN(n9606) );
  OAI21_X1 U16916 ( .B1(n793), .B2(n5120), .A(n11406), .ZN(n11415) );
  NAND2_X1 U16917 ( .A1(n12137), .A2(n5120), .ZN(n11406) );
  NAND3_X1 U16918 ( .A1(n5154), .A2(n32513), .A3(n5157), .ZN(n5121) );
  AND2_X1 U16919 ( .A1(n6459), .A2(n29395), .ZN(n5122) );
  NAND2_X1 U16920 ( .A1(n40355), .A2(n40354), .ZN(n5124) );
  NAND2_X1 U16923 ( .A1(n5131), .A2(n5129), .ZN(n5133) );
  AOI21_X1 U16924 ( .B1(n21100), .B2(n5130), .A(n21714), .ZN(n5129) );
  NAND3_X1 U16925 ( .A1(n21703), .A2(n21100), .A3(n20568), .ZN(n5131) );
  INV_X1 U16927 ( .A(n22189), .ZN(n20568) );
  NAND2_X1 U16928 ( .A1(n20567), .A2(n21094), .ZN(n5134) );
  NAND3_X1 U16930 ( .A1(n5139), .A2(n13058), .A3(n51685), .ZN(n5138) );
  NAND3_X1 U16933 ( .A1(n5147), .A2(n32620), .A3(n7626), .ZN(n32621) );
  INV_X1 U16934 ( .A(n31463), .ZN(n5147) );
  OR2_X1 U16935 ( .A1(n31463), .A2(n32620), .ZN(n31559) );
  OR2_X1 U16936 ( .A1(n50631), .A2(n50624), .ZN(n8017) );
  NAND2_X1 U16938 ( .A1(n5149), .A2(n47762), .ZN(n5148) );
  NOR2_X1 U16939 ( .A1(n47711), .A2(n47797), .ZN(n5149) );
  OAI22_X1 U16940 ( .A1(n8489), .A2(n21362), .B1(n21355), .B2(n21351), .ZN(
        n21352) );
  NAND2_X1 U16941 ( .A1(n5153), .A2(n33173), .ZN(n35162) );
  NAND3_X1 U16942 ( .A1(n36376), .A2(n36372), .A3(n5153), .ZN(n34950) );
  NAND2_X1 U16943 ( .A1(n36372), .A2(n35155), .ZN(n5152) );
  NAND2_X1 U16944 ( .A1(n35159), .A2(n5153), .ZN(n34937) );
  NAND3_X1 U16945 ( .A1(n5155), .A2(n32509), .A3(n32506), .ZN(n5154) );
  NAND2_X1 U16946 ( .A1(n32512), .A2(n51105), .ZN(n5155) );
  NAND2_X1 U16947 ( .A1(n32004), .A2(n32507), .ZN(n32506) );
  OAI21_X1 U16948 ( .B1(n32512), .B2(n5158), .A(n32511), .ZN(n5157) );
  NAND2_X1 U16949 ( .A1(n2480), .A2(n38649), .ZN(n36888) );
  NAND2_X1 U16950 ( .A1(n36887), .A2(n38940), .ZN(n38649) );
  NAND2_X2 U16951 ( .A1(n7493), .A2(n22113), .ZN(n28221) );
  INV_X1 U16952 ( .A(n51459), .ZN(n16911) );
  XNOR2_X1 U16953 ( .A(n15946), .B(n5161), .ZN(n15948) );
  XNOR2_X1 U16954 ( .A(n2323), .B(n51459), .ZN(n5161) );
  NAND3_X1 U16955 ( .A1(n5164), .A2(n6959), .A3(n50365), .ZN(n5163) );
  NAND2_X1 U16956 ( .A1(n6960), .A2(n50363), .ZN(n5164) );
  INV_X1 U16957 ( .A(n21810), .ZN(n5166) );
  NOR2_X1 U16958 ( .A1(n5166), .A2(n23785), .ZN(n5165) );
  NAND2_X1 U16959 ( .A1(n21403), .A2(n631), .ZN(n21558) );
  INV_X1 U16960 ( .A(n40087), .ZN(n40089) );
  NAND2_X1 U16961 ( .A1(n5169), .A2(n27145), .ZN(n5168) );
  NAND2_X1 U16962 ( .A1(n41268), .A2(n41265), .ZN(n41725) );
  OAI21_X2 U16963 ( .B1(n39422), .B2(n36894), .A(n36893), .ZN(n41268) );
  AND2_X1 U16964 ( .A1(n5171), .A2(n47127), .ZN(n5170) );
  NAND3_X1 U16965 ( .A1(n46862), .A2(n46861), .A3(n5171), .ZN(n46864) );
  OAI211_X1 U16966 ( .C1(n46682), .C2(n46681), .A(n46680), .B(n5171), .ZN(
        n46683) );
  NAND2_X1 U16967 ( .A1(n46854), .A2(n46840), .ZN(n5171) );
  NOR2_X1 U16969 ( .A1(n13323), .A2(n5176), .ZN(n14167) );
  OAI21_X1 U16970 ( .B1(n14600), .B2(n14011), .A(n5176), .ZN(n13324) );
  NAND3_X1 U16971 ( .A1(n13321), .A2(n14603), .A3(n5172), .ZN(n13328) );
  OR2_X1 U16972 ( .A1(n14170), .A2(n5176), .ZN(n5172) );
  AND2_X1 U16973 ( .A1(n5176), .A2(n14170), .ZN(n5173) );
  NAND2_X1 U16974 ( .A1(n14007), .A2(n5174), .ZN(n14014) );
  OAI21_X1 U16975 ( .B1(n14610), .B2(n5176), .A(n14605), .ZN(n5175) );
  NAND2_X1 U16976 ( .A1(n16673), .A2(n16678), .ZN(n21227) );
  NAND2_X1 U16977 ( .A1(n17313), .A2(n19113), .ZN(n19519) );
  OAI21_X1 U16979 ( .B1(n12515), .B2(n51709), .A(n5180), .ZN(n11545) );
  AOI21_X1 U16981 ( .B1(n12511), .B2(n5180), .A(n12525), .ZN(n11263) );
  OAI21_X1 U16982 ( .B1(n12513), .B2(n5180), .A(n12512), .ZN(n12519) );
  INV_X1 U16984 ( .A(n28616), .ZN(n5183) );
  OAI211_X1 U16986 ( .C1(n14963), .C2(n14962), .A(n14960), .B(n14961), .ZN(
        n5188) );
  XNOR2_X1 U16987 ( .A(n16265), .B(n18414), .ZN(n16272) );
  OAI211_X2 U16988 ( .C1(n17891), .C2(n19199), .A(n5187), .B(n5186), .ZN(
        n18414) );
  NAND2_X1 U16989 ( .A1(n17891), .A2(n5190), .ZN(n5187) );
  INV_X1 U16992 ( .A(n21413), .ZN(n21575) );
  NAND2_X1 U16993 ( .A1(n18823), .A2(n19989), .ZN(n21555) );
  NAND2_X1 U16994 ( .A1(n21758), .A2(n21756), .ZN(n23342) );
  NAND2_X1 U16995 ( .A1(n5196), .A2(n7129), .ZN(n5193) );
  NAND2_X1 U16996 ( .A1(n18323), .A2(n20090), .ZN(n5195) );
  NAND2_X1 U16997 ( .A1(n5197), .A2(n16788), .ZN(n5196) );
  NAND2_X1 U16998 ( .A1(n17500), .A2(n8624), .ZN(n5198) );
  INV_X1 U17000 ( .A(n16707), .ZN(n5200) );
  XNOR2_X1 U17001 ( .A(n5202), .B(n16706), .ZN(n5201) );
  XNOR2_X1 U17002 ( .A(n16705), .B(n17239), .ZN(n5202) );
  INV_X1 U17003 ( .A(n24030), .ZN(n5204) );
  NAND2_X1 U17004 ( .A1(n24028), .A2(n23675), .ZN(n22572) );
  NAND2_X1 U17005 ( .A1(n5207), .A2(n27655), .ZN(n5205) );
  OAI21_X1 U17006 ( .B1(n27657), .B2(n27656), .A(n27658), .ZN(n5206) );
  NOR2_X1 U17007 ( .A1(n5477), .A2(n27658), .ZN(n5207) );
  NAND2_X1 U17008 ( .A1(n5210), .A2(n14578), .ZN(n5209) );
  NOR2_X1 U17009 ( .A1(n15171), .A2(n7715), .ZN(n5210) );
  NAND2_X1 U17010 ( .A1(n10877), .A2(n14579), .ZN(n15171) );
  INV_X1 U17011 ( .A(n6403), .ZN(n5211) );
  INV_X1 U17012 ( .A(n30290), .ZN(n7997) );
  NAND2_X1 U17014 ( .A1(n40942), .A2(n5214), .ZN(n40944) );
  NAND4_X2 U17015 ( .A1(n31665), .A2(n5704), .A3(n5705), .A4(n28603), .ZN(
        n33753) );
  NAND2_X1 U17016 ( .A1(n5218), .A2(n36553), .ZN(n34995) );
  NAND2_X1 U17017 ( .A1(n37957), .A2(n5219), .ZN(n36544) );
  NAND2_X1 U17018 ( .A1(n36539), .A2(n37965), .ZN(n5219) );
  NAND2_X1 U17019 ( .A1(n34090), .A2(n34089), .ZN(n36539) );
  AND2_X1 U17020 ( .A1(n3347), .A2(n51432), .ZN(n9201) );
  NAND4_X1 U17021 ( .A1(n10468), .A2(n9564), .A3(n12637), .A4(n5220), .ZN(
        n9566) );
  XNOR2_X1 U17022 ( .A(n5221), .B(n51758), .ZN(n17320) );
  XNOR2_X1 U17023 ( .A(n17321), .B(n5221), .ZN(n15577) );
  OAI21_X1 U17024 ( .B1(n5226), .B2(n50396), .A(n50433), .ZN(n5223) );
  NAND2_X1 U17025 ( .A1(n50411), .A2(n50358), .ZN(n5226) );
  NAND2_X1 U17026 ( .A1(n50399), .A2(n50466), .ZN(n5225) );
  OAI211_X1 U17027 ( .C1(n32962), .C2(n32186), .A(n32965), .B(n5227), .ZN(
        n32178) );
  INV_X1 U17028 ( .A(n51107), .ZN(n29326) );
  NOR2_X1 U17029 ( .A1(n21196), .A2(n5231), .ZN(n17407) );
  NAND2_X1 U17030 ( .A1(n14999), .A2(n15131), .ZN(n10501) );
  XNOR2_X1 U17031 ( .A(n5232), .B(n25370), .ZN(n5233) );
  XNOR2_X1 U17032 ( .A(n25369), .B(n8208), .ZN(n5232) );
  XNOR2_X2 U17033 ( .A(n5233), .B(n25379), .ZN(n30209) );
  XNOR2_X1 U17034 ( .A(n5234), .B(n37137), .ZN(n37146) );
  XNOR2_X1 U17035 ( .A(n5234), .B(n37015), .ZN(n33791) );
  NAND2_X1 U17036 ( .A1(n36337), .A2(n5235), .ZN(n5236) );
  INV_X1 U17037 ( .A(n35017), .ZN(n38145) );
  NAND2_X1 U17038 ( .A1(n5236), .A2(n36167), .ZN(n36169) );
  INV_X1 U17039 ( .A(n50279), .ZN(n50253) );
  AND2_X1 U17040 ( .A1(n28669), .A2(n27852), .ZN(n27856) );
  XNOR2_X1 U17041 ( .A(n5239), .B(n33395), .ZN(n33726) );
  XNOR2_X1 U17042 ( .A(n5238), .B(n35095), .ZN(n33395) );
  NAND2_X1 U17043 ( .A1(n31039), .A2(n31826), .ZN(n31030) );
  NAND2_X1 U17044 ( .A1(n30206), .A2(n30216), .ZN(n5240) );
  NAND2_X1 U17045 ( .A1(n5242), .A2(n36638), .ZN(n36646) );
  NAND2_X1 U17046 ( .A1(n5242), .A2(n34199), .ZN(n34200) );
  NAND2_X1 U17047 ( .A1(n34198), .A2(n38093), .ZN(n5242) );
  NAND2_X1 U17049 ( .A1(n19700), .A2(n19699), .ZN(n5243) );
  AOI22_X1 U17050 ( .A1(n45759), .A2(n46622), .B1(n44423), .B2(n5246), .ZN(
        n45770) );
  NAND2_X1 U17051 ( .A1(n44423), .A2(n5245), .ZN(n6750) );
  NAND2_X1 U17052 ( .A1(n5247), .A2(n12484), .ZN(n5255) );
  OAI22_X1 U17053 ( .A1(n12471), .A2(n12475), .B1(n12483), .B2(n12486), .ZN(
        n5247) );
  AND2_X1 U17054 ( .A1(n2116), .A2(n11485), .ZN(n11895) );
  NAND2_X1 U17055 ( .A1(n11484), .A2(n11487), .ZN(n5248) );
  AOI22_X1 U17056 ( .A1(n11487), .A2(n11486), .B1(n2116), .B2(n5250), .ZN(
        n5249) );
  INV_X1 U17057 ( .A(n11485), .ZN(n5251) );
  INV_X1 U17058 ( .A(n11489), .ZN(n5252) );
  NAND2_X1 U17059 ( .A1(n510), .A2(n11908), .ZN(n5254) );
  NAND3_X1 U17060 ( .A1(n21533), .A2(n21543), .A3(n6929), .ZN(n21536) );
  NAND2_X1 U17061 ( .A1(n21548), .A2(n6929), .ZN(n19939) );
  XNOR2_X1 U17062 ( .A(n5256), .B(n34570), .ZN(n15515) );
  XNOR2_X1 U17063 ( .A(n16142), .B(n5256), .ZN(n18580) );
  XNOR2_X1 U17065 ( .A(n5256), .B(n16237), .ZN(n17652) );
  NAND2_X1 U17066 ( .A1(n27754), .A2(n29468), .ZN(n5261) );
  NAND2_X1 U17067 ( .A1(n26788), .A2(n29456), .ZN(n27751) );
  OR2_X1 U17068 ( .A1(n36778), .A2(n2100), .ZN(n36780) );
  OAI21_X1 U17069 ( .B1(n39282), .B2(n39273), .A(n2100), .ZN(n37204) );
  NAND2_X1 U17070 ( .A1(n38684), .A2(n2100), .ZN(n38695) );
  NOR2_X1 U17071 ( .A1(n50548), .A2(n50508), .ZN(n5264) );
  NAND2_X1 U17075 ( .A1(n40943), .A2(n40986), .ZN(n40990) );
  NAND3_X2 U17076 ( .A1(n5265), .A2(n37946), .A3(n37945), .ZN(n40986) );
  INV_X1 U17077 ( .A(n5266), .ZN(n22753) );
  NAND2_X1 U17078 ( .A1(n23048), .A2(n23045), .ZN(n5266) );
  NAND2_X1 U17079 ( .A1(n22754), .A2(n5266), .ZN(n22756) );
  NAND2_X1 U17080 ( .A1(n26197), .A2(n5267), .ZN(n29546) );
  NAND2_X1 U17081 ( .A1(n11539), .A2(n642), .ZN(n12522) );
  NAND2_X1 U17082 ( .A1(n14938), .A2(n14957), .ZN(n14952) );
  INV_X1 U17083 ( .A(n19702), .ZN(n5271) );
  OR2_X1 U17084 ( .A1(n51434), .A2(n19702), .ZN(n21174) );
  NAND2_X1 U17085 ( .A1(n5274), .A2(n5273), .ZN(n5272) );
  XNOR2_X1 U17086 ( .A(n14509), .B(n19250), .ZN(n14511) );
  NAND3_X1 U17087 ( .A1(n27777), .A2(n30597), .A3(n5277), .ZN(n27778) );
  NAND2_X1 U17088 ( .A1(n31089), .A2(n30599), .ZN(n5277) );
  OR2_X1 U17089 ( .A1(n5283), .A2(n5281), .ZN(n47548) );
  NAND2_X1 U17090 ( .A1(n47557), .A2(n51346), .ZN(n5283) );
  OR2_X1 U17091 ( .A1(n5279), .A2(n5283), .ZN(n47494) );
  NAND2_X1 U17092 ( .A1(n51303), .A2(n47579), .ZN(n5281) );
  NAND2_X1 U17093 ( .A1(n47518), .A2(n5280), .ZN(n5279) );
  AND2_X1 U17094 ( .A1(n51286), .A2(n52045), .ZN(n5280) );
  NAND2_X1 U17095 ( .A1(n5283), .A2(n5282), .ZN(n47534) );
  OAI21_X1 U17096 ( .B1(n5287), .B2(n50728), .A(n50650), .ZN(n50651) );
  NAND2_X1 U17097 ( .A1(n50665), .A2(n50721), .ZN(n5287) );
  AOI21_X1 U17098 ( .B1(n44600), .B2(n46797), .A(n43798), .ZN(n5288) );
  NAND2_X1 U17099 ( .A1(n22673), .A2(n22674), .ZN(n5290) );
  NAND2_X1 U17100 ( .A1(n628), .A2(n52133), .ZN(n5291) );
  NAND2_X1 U17101 ( .A1(n19151), .A2(n5293), .ZN(n19152) );
  INV_X1 U17102 ( .A(n23247), .ZN(n5294) );
  NAND2_X1 U17103 ( .A1(n11121), .A2(n5298), .ZN(n5297) );
  NAND2_X1 U17104 ( .A1(n11937), .A2(n12438), .ZN(n5299) );
  NAND4_X2 U17105 ( .A1(n27021), .A2(n27022), .A3(n27019), .A4(n27020), .ZN(
        n31340) );
  NAND4_X2 U17106 ( .A1(n27060), .A2(n27063), .A3(n27062), .A4(n27061), .ZN(
        n29602) );
  NAND2_X1 U17107 ( .A1(n30823), .A2(n5914), .ZN(n5301) );
  NAND3_X1 U17108 ( .A1(n5304), .A2(n6268), .A3(n5303), .ZN(n5302) );
  NAND2_X1 U17109 ( .A1(n32634), .A2(n32639), .ZN(n5303) );
  NAND3_X1 U17110 ( .A1(n5306), .A2(n30813), .A3(n5305), .ZN(n32944) );
  NAND3_X1 U17111 ( .A1(n30812), .A2(n31701), .A3(n32126), .ZN(n5306) );
  INV_X1 U17112 ( .A(n5687), .ZN(n5307) );
  NAND3_X1 U17113 ( .A1(n5307), .A2(n10356), .A3(n10354), .ZN(n9386) );
  OR2_X2 U17114 ( .A1(n5308), .A2(n5964), .ZN(n40774) );
  OAI211_X1 U17115 ( .C1(n46625), .C2(n46626), .A(n5309), .B(n46624), .ZN(
        n46647) );
  NAND4_X1 U17116 ( .A1(n6755), .A2(n6753), .A3(n44419), .A4(n5309), .ZN(n6752) );
  INV_X1 U17117 ( .A(n22169), .ZN(n22369) );
  NAND2_X1 U17118 ( .A1(n38560), .A2(n5312), .ZN(n38564) );
  NAND2_X1 U17119 ( .A1(n6774), .A2(n5312), .ZN(n5504) );
  NAND3_X1 U17120 ( .A1(n10018), .A2(n11663), .A3(n11649), .ZN(n5315) );
  NAND3_X1 U17121 ( .A1(n11644), .A2(n11663), .A3(n11655), .ZN(n11646) );
  NAND3_X1 U17123 ( .A1(n45965), .A2(n45963), .A3(n45964), .ZN(n47193) );
  NAND2_X1 U17124 ( .A1(n41324), .A2(n52215), .ZN(n5316) );
  NAND2_X1 U17125 ( .A1(n5317), .A2(n41902), .ZN(n41324) );
  NOR2_X1 U17126 ( .A1(n41319), .A2(n4703), .ZN(n5317) );
  INV_X1 U17127 ( .A(n41319), .ZN(n39822) );
  OR2_X1 U17128 ( .A1(n45542), .A2(n48205), .ZN(n5322) );
  NAND2_X1 U17129 ( .A1(n45544), .A2(n45543), .ZN(n5320) );
  NAND2_X1 U17130 ( .A1(n44873), .A2(n52154), .ZN(n45757) );
  NAND3_X1 U17131 ( .A1(n44873), .A2(n52153), .A3(n5325), .ZN(n47907) );
  NAND2_X1 U17132 ( .A1(n33150), .A2(n38043), .ZN(n5327) );
  NOR2_X1 U17133 ( .A1(n5330), .A2(n51746), .ZN(n5329) );
  NAND2_X1 U17134 ( .A1(n28329), .A2(n1981), .ZN(n27513) );
  INV_X1 U17136 ( .A(n23414), .ZN(n23426) );
  NAND2_X1 U17137 ( .A1(n590), .A2(n17523), .ZN(n16801) );
  INV_X1 U17138 ( .A(n6363), .ZN(n17523) );
  NOR2_X1 U17139 ( .A1(n6363), .A2(n18287), .ZN(n5333) );
  INV_X1 U17140 ( .A(n5334), .ZN(n30923) );
  OAI21_X1 U17141 ( .B1(n30910), .B2(n31099), .A(n30909), .ZN(n5334) );
  NAND2_X1 U17142 ( .A1(n5334), .A2(n31092), .ZN(n31102) );
  INV_X1 U17143 ( .A(n19396), .ZN(n5336) );
  NAND2_X1 U17144 ( .A1(n19398), .A2(n17575), .ZN(n19387) );
  NAND2_X1 U17145 ( .A1(n27660), .A2(n736), .ZN(n26874) );
  NAND2_X1 U17146 ( .A1(n19917), .A2(n21715), .ZN(n21101) );
  NAND2_X1 U17149 ( .A1(n5338), .A2(n13049), .ZN(n5337) );
  NAND2_X1 U17150 ( .A1(n6013), .A2(n31096), .ZN(n30591) );
  XNOR2_X1 U17152 ( .A(n15542), .B(n2384), .ZN(n16942) );
  NAND2_X1 U17155 ( .A1(n5348), .A2(n5347), .ZN(n5346) );
  NAND3_X1 U17156 ( .A1(n20135), .A2(n17065), .A3(n19061), .ZN(n18358) );
  XNOR2_X2 U17157 ( .A(n5349), .B(n16577), .ZN(n20132) );
  XNOR2_X2 U17158 ( .A(n8656), .B(Key[162]), .ZN(n11410) );
  XNOR2_X1 U17159 ( .A(n563), .B(n16568), .ZN(n5350) );
  INV_X1 U17161 ( .A(n23481), .ZN(n5352) );
  NAND2_X1 U17162 ( .A1(n23487), .A2(n21974), .ZN(n21971) );
  NAND2_X1 U17163 ( .A1(n21981), .A2(n23481), .ZN(n23487) );
  INV_X1 U17164 ( .A(n39966), .ZN(n5354) );
  NAND3_X1 U17165 ( .A1(n27104), .A2(n28872), .A3(n29032), .ZN(n29043) );
  NAND2_X1 U17166 ( .A1(n2092), .A2(n46730), .ZN(n5356) );
  NAND2_X1 U17167 ( .A1(n41811), .A2(n5357), .ZN(n46732) );
  NAND3_X1 U17168 ( .A1(n13759), .A2(n13760), .A3(n13761), .ZN(n7982) );
  INV_X1 U17169 ( .A(n35405), .ZN(n5482) );
  OAI21_X1 U17170 ( .B1(n35407), .B2(n35405), .A(n37667), .ZN(n37668) );
  NAND3_X1 U17171 ( .A1(n38339), .A2(n35405), .A3(n38329), .ZN(n37187) );
  NAND2_X1 U17172 ( .A1(n24034), .A2(n22097), .ZN(n22099) );
  NAND2_X1 U17173 ( .A1(n19970), .A2(n20829), .ZN(n19971) );
  OAI22_X1 U17174 ( .A1(n18239), .A2(n18236), .B1(n20211), .B2(n20209), .ZN(
        n5361) );
  NAND3_X1 U17175 ( .A1(n51344), .A2(n2092), .A3(n45188), .ZN(n46554) );
  NAND3_X1 U17177 ( .A1(n24289), .A2(n24290), .A3(n24291), .ZN(n5363) );
  OAI211_X1 U17178 ( .C1(n24296), .C2(n24295), .A(n24294), .B(n5363), .ZN(
        n24297) );
  NAND2_X1 U17179 ( .A1(n38503), .A2(n38505), .ZN(n38490) );
  OAI22_X1 U17180 ( .A1(n38493), .A2(n37516), .B1(n37517), .B2(n37392), .ZN(
        n38491) );
  NAND2_X1 U17181 ( .A1(n38494), .A2(n37385), .ZN(n37392) );
  NAND2_X1 U17183 ( .A1(n5364), .A2(n38494), .ZN(n38505) );
  INV_X1 U17184 ( .A(n38495), .ZN(n5364) );
  NAND3_X1 U17185 ( .A1(n50934), .A2(n50901), .A3(n50955), .ZN(n47398) );
  NAND3_X1 U17186 ( .A1(n12178), .A2(n10418), .A3(n12177), .ZN(n11333) );
  XNOR2_X1 U17187 ( .A(n33540), .B(n33542), .ZN(n5367) );
  NAND2_X1 U17188 ( .A1(n51256), .A2(n10368), .ZN(n5368) );
  OAI21_X1 U17189 ( .B1(n12118), .B2(n5368), .A(n9638), .ZN(n9695) );
  AOI21_X1 U17190 ( .B1(n10696), .B2(n5368), .A(n12118), .ZN(n10697) );
  NAND2_X1 U17191 ( .A1(n30715), .A2(n5639), .ZN(n5369) );
  NAND2_X1 U17192 ( .A1(n32478), .A2(n32473), .ZN(n32016) );
  AND2_X1 U17193 ( .A1(n23813), .A2(n3270), .ZN(n22739) );
  MUX2_X1 U17194 ( .A(n27696), .B(n29549), .S(n29543), .Z(n6017) );
  INV_X1 U17195 ( .A(n5373), .ZN(n20227) );
  NAND3_X1 U17196 ( .A1(n20686), .A2(n5373), .A3(n20672), .ZN(n18104) );
  NOR2_X1 U17197 ( .A1(n5373), .A2(n18101), .ZN(n15923) );
  OR2_X1 U17198 ( .A1(n8301), .A2(n5373), .ZN(n8300) );
  OAI21_X1 U17199 ( .B1(n760), .B2(n5373), .A(n20686), .ZN(n5695) );
  XNOR2_X1 U17200 ( .A(n43259), .B(n5374), .ZN(n43180) );
  XNOR2_X1 U17201 ( .A(n5375), .B(n5376), .ZN(n5374) );
  XNOR2_X1 U17202 ( .A(n43360), .B(n52085), .ZN(n5375) );
  XNOR2_X1 U17203 ( .A(n43115), .B(n43114), .ZN(n5376) );
  XNOR2_X1 U17204 ( .A(n37262), .B(n33818), .ZN(n8283) );
  NAND2_X1 U17205 ( .A1(n5378), .A2(n27778), .ZN(n5377) );
  NAND3_X1 U17206 ( .A1(n27776), .A2(n30605), .A3(n29683), .ZN(n5378) );
  XNOR2_X1 U17207 ( .A(n45284), .B(n5379), .ZN(n42272) );
  XNOR2_X1 U17208 ( .A(n5379), .B(n42386), .ZN(n42387) );
  XNOR2_X1 U17209 ( .A(n46069), .B(n5379), .ZN(n42626) );
  XNOR2_X2 U17210 ( .A(n9094), .B(Key[165]), .ZN(n11634) );
  INV_X1 U17211 ( .A(n11464), .ZN(n11633) );
  INV_X1 U17212 ( .A(n10889), .ZN(n5380) );
  NAND2_X1 U17213 ( .A1(n13501), .A2(n13514), .ZN(n10889) );
  NAND4_X1 U17214 ( .A1(n22552), .A2(n22550), .A3(n22551), .A4(n22553), .ZN(
        n5384) );
  XNOR2_X1 U17215 ( .A(n22554), .B(n5381), .ZN(n24140) );
  INV_X1 U17216 ( .A(n7939), .ZN(n5381) );
  XNOR2_X1 U17217 ( .A(n22554), .B(n5382), .ZN(n25613) );
  XNOR2_X1 U17218 ( .A(n5383), .B(n22554), .ZN(n24619) );
  NAND2_X1 U17219 ( .A1(n20044), .A2(n771), .ZN(n17447) );
  INV_X1 U17220 ( .A(n16395), .ZN(n5385) );
  XNOR2_X1 U17221 ( .A(n24764), .B(n24773), .ZN(n5387) );
  NAND3_X1 U17222 ( .A1(n21144), .A2(n21744), .A3(n23336), .ZN(n21734) );
  NAND4_X1 U17223 ( .A1(n48796), .A2(n48817), .A3(n48799), .A4(n48829), .ZN(
        n5391) );
  AND2_X1 U17224 ( .A1(n52434), .A2(n48808), .ZN(n48799) );
  OAI21_X1 U17225 ( .B1(n52090), .B2(n45745), .A(n5393), .ZN(n5392) );
  AOI21_X1 U17226 ( .B1(n45746), .B2(n52090), .A(n8340), .ZN(n5393) );
  NAND3_X1 U17227 ( .A1(n5395), .A2(n14128), .A3(n10865), .ZN(n10866) );
  NAND2_X1 U17228 ( .A1(n13457), .A2(n5394), .ZN(n13460) );
  NOR2_X1 U17229 ( .A1(n15168), .A2(n15163), .ZN(n5394) );
  NAND2_X1 U17230 ( .A1(n10876), .A2(n5395), .ZN(n10880) );
  INV_X1 U17231 ( .A(n15168), .ZN(n5395) );
  XNOR2_X1 U17232 ( .A(n2168), .B(n35809), .ZN(n34272) );
  XNOR2_X1 U17233 ( .A(n35618), .B(n2167), .ZN(n35621) );
  XNOR2_X1 U17234 ( .A(n2167), .B(n35237), .ZN(n34343) );
  XNOR2_X1 U17235 ( .A(n2598), .B(n2168), .ZN(n36959) );
  NAND2_X1 U17236 ( .A1(n397), .A2(n41276), .ZN(n41035) );
  NAND2_X1 U17237 ( .A1(n35172), .A2(n38228), .ZN(n5396) );
  NAND2_X1 U17238 ( .A1(n35173), .A2(n35174), .ZN(n5397) );
  NAND2_X1 U17239 ( .A1(n38413), .A2(n38412), .ZN(n5400) );
  NAND2_X1 U17240 ( .A1(n7778), .A2(n38405), .ZN(n5404) );
  NOR2_X1 U17241 ( .A1(n36516), .A2(n37976), .ZN(n5405) );
  XNOR2_X2 U17242 ( .A(n26253), .B(n26252), .ZN(n28623) );
  XNOR2_X2 U17243 ( .A(n18772), .B(n18771), .ZN(n21584) );
  NAND2_X1 U17244 ( .A1(n20784), .A2(n20785), .ZN(n5407) );
  INV_X1 U17246 ( .A(n8781), .ZN(n5408) );
  OAI211_X1 U17248 ( .C1(n20614), .C2(n5409), .A(n21523), .B(n20183), .ZN(
        n20184) );
  INV_X1 U17251 ( .A(n352), .ZN(n5414) );
  NAND2_X1 U17252 ( .A1(n51116), .A2(n25479), .ZN(n29190) );
  NAND2_X1 U17253 ( .A1(n7909), .A2(n377), .ZN(n29187) );
  OAI21_X1 U17254 ( .B1(n41347), .B2(n5416), .A(n39887), .ZN(n39888) );
  NAND2_X1 U17256 ( .A1(n23480), .A2(n23477), .ZN(n20996) );
  NAND2_X2 U17257 ( .A1(n16813), .A2(n16812), .ZN(n23479) );
  INV_X1 U17258 ( .A(n39266), .ZN(n38689) );
  NAND2_X1 U17260 ( .A1(n10063), .A2(n13787), .ZN(n10901) );
  NAND2_X1 U17261 ( .A1(n13174), .A2(n13161), .ZN(n13787) );
  AOI21_X1 U17262 ( .B1(n29276), .B2(n29277), .A(n51706), .ZN(n5418) );
  INV_X1 U17263 ( .A(n5418), .ZN(n5419) );
  NAND2_X1 U17264 ( .A1(n32105), .A2(n32107), .ZN(n30898) );
  NAND3_X1 U17265 ( .A1(n27935), .A2(n27934), .A3(n27933), .ZN(n5420) );
  NAND3_X1 U17266 ( .A1(n30625), .A2(n30624), .A3(n32303), .ZN(n31747) );
  INV_X1 U17267 ( .A(n38135), .ZN(n38055) );
  XNOR2_X1 U17270 ( .A(n5423), .B(n33938), .ZN(n31103) );
  XNOR2_X1 U17271 ( .A(n2133), .B(n36748), .ZN(n33790) );
  XNOR2_X1 U17272 ( .A(n2133), .B(n33433), .ZN(n33434) );
  XNOR2_X1 U17273 ( .A(n34608), .B(n5423), .ZN(n34609) );
  XNOR2_X1 U17274 ( .A(n2133), .B(n35471), .ZN(n35119) );
  XNOR2_X1 U17275 ( .A(n5423), .B(n35296), .ZN(n35756) );
  AOI21_X1 U17276 ( .B1(n25516), .B2(n28714), .A(n8242), .ZN(n29279) );
  NAND2_X1 U17277 ( .A1(n5424), .A2(n29192), .ZN(n28714) );
  NOR2_X1 U17278 ( .A1(n5425), .A2(n5522), .ZN(n5424) );
  INV_X1 U17279 ( .A(n51116), .ZN(n5425) );
  XNOR2_X1 U17280 ( .A(n5426), .B(n42451), .ZN(n42457) );
  XNOR2_X1 U17281 ( .A(n5427), .B(n42449), .ZN(n5426) );
  XNOR2_X1 U17282 ( .A(n5428), .B(n42448), .ZN(n5427) );
  XNOR2_X1 U17283 ( .A(n42662), .B(n44216), .ZN(n5428) );
  OAI211_X1 U17284 ( .C1(n38232), .C2(n40924), .A(n41386), .B(n5431), .ZN(
        n5430) );
  XNOR2_X1 U17285 ( .A(n42129), .B(n41821), .ZN(n5433) );
  INV_X1 U17286 ( .A(n30866), .ZN(n5438) );
  OAI21_X1 U17287 ( .B1(n5438), .B2(n31155), .A(n31160), .ZN(n5442) );
  NAND2_X1 U17288 ( .A1(n5441), .A2(n2388), .ZN(n5440) );
  NAND2_X1 U17289 ( .A1(n31462), .A2(n32618), .ZN(n5441) );
  NAND2_X1 U17290 ( .A1(n47334), .A2(n47335), .ZN(n47046) );
  INV_X1 U17291 ( .A(n38132), .ZN(n36340) );
  XNOR2_X2 U17292 ( .A(n31964), .B(n31965), .ZN(n38132) );
  INV_X1 U17293 ( .A(n35010), .ZN(n5443) );
  NAND2_X1 U17295 ( .A1(n10499), .A2(n14999), .ZN(n13701) );
  XNOR2_X1 U17296 ( .A(n50982), .B(n5445), .ZN(n32606) );
  XNOR2_X1 U17297 ( .A(n36818), .B(n5445), .ZN(n31657) );
  XNOR2_X1 U17298 ( .A(n34419), .B(n5445), .ZN(n34423) );
  XNOR2_X1 U17299 ( .A(n35296), .B(n5445), .ZN(n5810) );
  XNOR2_X1 U17300 ( .A(n34876), .B(n5445), .ZN(n34877) );
  NAND3_X1 U17302 ( .A1(n5446), .A2(n20943), .A3(n51081), .ZN(n20947) );
  AND2_X1 U17303 ( .A1(n23178), .A2(n23172), .ZN(n22067) );
  NAND2_X1 U17304 ( .A1(n23175), .A2(n23167), .ZN(n23172) );
  NAND2_X1 U17305 ( .A1(n3717), .A2(n23171), .ZN(n5447) );
  NAND3_X1 U17306 ( .A1(n31470), .A2(n31471), .A3(n32609), .ZN(n31156) );
  INV_X1 U17308 ( .A(n40686), .ZN(n40675) );
  NOR2_X1 U17309 ( .A1(n39931), .A2(n39929), .ZN(n40674) );
  NAND2_X1 U17310 ( .A1(n35215), .A2(n36051), .ZN(n35880) );
  AND2_X1 U17311 ( .A1(n39354), .A2(n39355), .ZN(n5450) );
  INV_X1 U17313 ( .A(n47356), .ZN(n5451) );
  NAND3_X1 U17314 ( .A1(n5451), .A2(n47354), .A3(n49982), .ZN(n49618) );
  NOR2_X1 U17315 ( .A1(n5453), .A2(n5640), .ZN(n5452) );
  INV_X1 U17316 ( .A(n28811), .ZN(n5453) );
  XNOR2_X1 U17317 ( .A(n37039), .B(n2154), .ZN(n37041) );
  XNOR2_X1 U17318 ( .A(n2155), .B(n34720), .ZN(n34721) );
  XNOR2_X1 U17319 ( .A(n34238), .B(n2155), .ZN(n33188) );
  XNOR2_X1 U17320 ( .A(n2155), .B(n36952), .ZN(n36953) );
  MUX2_X1 U17321 ( .A(n5459), .B(n22505), .S(n22504), .Z(n22511) );
  NAND2_X1 U17322 ( .A1(n5462), .A2(n11291), .ZN(n5461) );
  OAI21_X1 U17323 ( .B1(n14400), .B2(n11289), .A(n12861), .ZN(n5462) );
  AND2_X1 U17324 ( .A1(n14410), .A2(n14393), .ZN(n12861) );
  NAND2_X1 U17325 ( .A1(n8916), .A2(n10831), .ZN(n12506) );
  AND2_X1 U17326 ( .A1(n5737), .A2(n22359), .ZN(n22167) );
  XNOR2_X2 U17327 ( .A(n9172), .B(Key[96]), .ZN(n12659) );
  NAND2_X1 U17328 ( .A1(n35894), .A2(n37195), .ZN(n38328) );
  INV_X1 U17329 ( .A(n23440), .ZN(n22587) );
  OAI21_X1 U17330 ( .B1(n19554), .B2(n23435), .A(n21999), .ZN(n19555) );
  NAND2_X1 U17331 ( .A1(n5466), .A2(n30846), .ZN(n5468) );
  NAND2_X1 U17332 ( .A1(n5467), .A2(n30576), .ZN(n5466) );
  NAND2_X1 U17333 ( .A1(n31826), .A2(n31033), .ZN(n5467) );
  NAND2_X1 U17335 ( .A1(n26711), .A2(n50986), .ZN(n30581) );
  INV_X1 U17336 ( .A(n29288), .ZN(n26077) );
  NAND2_X1 U17337 ( .A1(n29294), .A2(n51518), .ZN(n5469) );
  NAND2_X1 U17338 ( .A1(n51517), .A2(n26083), .ZN(n26649) );
  NAND2_X1 U17339 ( .A1(n50269), .A2(n50262), .ZN(n47068) );
  NAND2_X1 U17340 ( .A1(n28324), .A2(n29763), .ZN(n5471) );
  NAND2_X1 U17341 ( .A1(n28323), .A2(n29063), .ZN(n5472) );
  NAND2_X1 U17343 ( .A1(n11941), .A2(n5473), .ZN(n11112) );
  XNOR2_X1 U17344 ( .A(n7132), .B(n2343), .ZN(n5474) );
  NAND2_X1 U17345 ( .A1(n8429), .A2(n39272), .ZN(n39263) );
  OAI21_X1 U17346 ( .B1(n31561), .B2(n31475), .A(n6966), .ZN(n5480) );
  NAND2_X1 U17347 ( .A1(n5481), .A2(n32616), .ZN(n5479) );
  NAND2_X1 U17348 ( .A1(n50565), .A2(n50539), .ZN(n5483) );
  INV_X1 U17349 ( .A(n8881), .ZN(n11107) );
  INV_X1 U17350 ( .A(n8882), .ZN(n5484) );
  NOR2_X1 U17351 ( .A1(n5487), .A2(n5485), .ZN(n5489) );
  NOR2_X1 U17352 ( .A1(n38750), .A2(n5488), .ZN(n5490) );
  AND2_X2 U17353 ( .A1(n5490), .A2(n38751), .ZN(n43909) );
  OAI21_X1 U17354 ( .B1(n5665), .B2(n32407), .A(n5495), .ZN(n5496) );
  NAND3_X1 U17355 ( .A1(n7430), .A2(n32407), .A3(n32066), .ZN(n5495) );
  INV_X1 U17356 ( .A(n19156), .ZN(n5499) );
  NAND2_X1 U17357 ( .A1(n5500), .A2(n21425), .ZN(n20837) );
  NAND2_X1 U17359 ( .A1(n48156), .A2(n5502), .ZN(n48102) );
  NAND2_X1 U17360 ( .A1(n48112), .A2(n5502), .ZN(n48160) );
  AND4_X2 U17361 ( .A1(n45608), .A2(n45607), .A3(n45605), .A4(n45606), .ZN(
        n48100) );
  NAND4_X1 U17362 ( .A1(n35152), .A2(n5504), .A3(n6776), .A4(n5503), .ZN(n6775) );
  NAND2_X1 U17363 ( .A1(n38198), .A2(n35146), .ZN(n5505) );
  NAND2_X1 U17364 ( .A1(n5506), .A2(n47355), .ZN(n43454) );
  INV_X1 U17365 ( .A(n11399), .ZN(n9601) );
  NAND2_X1 U17366 ( .A1(n11399), .A2(n5507), .ZN(n5509) );
  INV_X1 U17367 ( .A(n11400), .ZN(n5507) );
  NAND2_X1 U17368 ( .A1(n5509), .A2(n9607), .ZN(n5508) );
  NAND2_X1 U17369 ( .A1(n9434), .A2(n11423), .ZN(n5512) );
  XNOR2_X1 U17370 ( .A(n24489), .B(n21998), .ZN(n5517) );
  NAND2_X1 U17371 ( .A1(n18061), .A2(n18071), .ZN(n18341) );
  NOR2_X1 U17372 ( .A1(n39397), .A2(n2139), .ZN(n37895) );
  AOI21_X1 U17373 ( .B1(n5521), .B2(n45203), .A(n48463), .ZN(n45621) );
  OAI211_X1 U17374 ( .C1(n46415), .C2(n45207), .A(n48470), .B(n5521), .ZN(
        n42513) );
  NAND3_X1 U17375 ( .A1(n17433), .A2(n18332), .A3(n403), .ZN(n17434) );
  NAND2_X1 U17376 ( .A1(n5656), .A2(n5522), .ZN(n27780) );
  INV_X1 U17377 ( .A(n28708), .ZN(n5522) );
  NAND2_X1 U17378 ( .A1(n34194), .A2(n36319), .ZN(n5523) );
  NAND2_X1 U17379 ( .A1(n34195), .A2(n34196), .ZN(n5524) );
  NAND2_X1 U17380 ( .A1(n5527), .A2(n36317), .ZN(n5526) );
  NAND2_X1 U17381 ( .A1(n38072), .A2(n34185), .ZN(n5527) );
  AND3_X1 U17382 ( .A1(n17443), .A2(n17445), .A3(n17444), .ZN(n5529) );
  NAND2_X1 U17384 ( .A1(n36628), .A2(n5530), .ZN(n33274) );
  NOR2_X1 U17385 ( .A1(n36628), .A2(n5530), .ZN(n36631) );
  OR2_X1 U17386 ( .A1(n34960), .A2(n5530), .ZN(n36641) );
  OAI22_X1 U17387 ( .A1(n695), .A2(n36320), .B1(n1360), .B2(n5530), .ZN(n36321) );
  XNOR2_X1 U17388 ( .A(n51522), .B(n38132), .ZN(n38138) );
  XNOR2_X1 U17389 ( .A(n42776), .B(n5532), .ZN(n42777) );
  NAND2_X1 U17390 ( .A1(n18901), .A2(n21519), .ZN(n5537) );
  NAND2_X1 U17391 ( .A1(n18902), .A2(n21521), .ZN(n5538) );
  OR2_X1 U17392 ( .A1(n36547), .A2(n37962), .ZN(n6184) );
  NAND2_X1 U17393 ( .A1(n36541), .A2(n699), .ZN(n37962) );
  XNOR2_X2 U17394 ( .A(Key[135]), .B(Ciphertext[158]), .ZN(n10296) );
  NAND2_X1 U17395 ( .A1(n22960), .A2(n23314), .ZN(n21861) );
  INV_X1 U17396 ( .A(n13968), .ZN(n5540) );
  NAND2_X1 U17397 ( .A1(n5540), .A2(n639), .ZN(n14221) );
  INV_X1 U17398 ( .A(n5541), .ZN(n21637) );
  NAND2_X1 U17399 ( .A1(n5541), .A2(n21620), .ZN(n20250) );
  NAND2_X1 U17400 ( .A1(n20692), .A2(n5541), .ZN(n20693) );
  NAND2_X1 U17401 ( .A1(n5542), .A2(n2175), .ZN(n19577) );
  INV_X1 U17402 ( .A(n22918), .ZN(n22907) );
  OAI22_X1 U17403 ( .A1(n22164), .A2(n5543), .B1(n22350), .B2(n22914), .ZN(
        n19575) );
  NAND2_X1 U17404 ( .A1(n29976), .A2(n31700), .ZN(n6678) );
  NAND2_X1 U17405 ( .A1(n52120), .A2(n41539), .ZN(n5546) );
  NAND2_X1 U17407 ( .A1(n52198), .A2(n41245), .ZN(n41680) );
  INV_X1 U17408 ( .A(n39306), .ZN(n5555) );
  NAND2_X1 U17409 ( .A1(n48432), .A2(n48264), .ZN(n5562) );
  NAND2_X1 U17410 ( .A1(n5563), .A2(n52144), .ZN(n5564) );
  INV_X1 U17411 ( .A(n25410), .ZN(n5563) );
  INV_X1 U17412 ( .A(n25410), .ZN(n25418) );
  NAND2_X1 U17413 ( .A1(n38942), .A2(n39412), .ZN(n5565) );
  OAI211_X1 U17414 ( .C1(n41620), .C2(n41691), .A(n41697), .B(n41619), .ZN(
        n41624) );
  NAND2_X1 U17415 ( .A1(n26647), .A2(n26068), .ZN(n5566) );
  NAND2_X1 U17416 ( .A1(n27738), .A2(n27739), .ZN(n5567) );
  NAND2_X1 U17418 ( .A1(n38723), .A2(n616), .ZN(n5569) );
  NAND3_X1 U17419 ( .A1(n35851), .A2(n39288), .A3(n5571), .ZN(n35856) );
  INV_X1 U17420 ( .A(n47591), .ZN(n47206) );
  NAND2_X1 U17421 ( .A1(n5572), .A2(n47616), .ZN(n47624) );
  OAI211_X1 U17422 ( .C1(n5575), .C2(n47614), .A(n5574), .B(n47615), .ZN(n5572) );
  NAND2_X1 U17423 ( .A1(n51400), .A2(n47620), .ZN(n5573) );
  OR2_X1 U17424 ( .A1(n6831), .A2(n47619), .ZN(n5574) );
  NOR2_X1 U17425 ( .A1(n5577), .A2(n5576), .ZN(n5579) );
  NOR2_X1 U17426 ( .A1(n7030), .A2(n7033), .ZN(n5577) );
  NAND3_X2 U17427 ( .A1(n5579), .A2(n7032), .A3(n5578), .ZN(n43244) );
  NAND2_X1 U17428 ( .A1(n14561), .A2(n13669), .ZN(n5580) );
  NAND4_X2 U17429 ( .A1(n11321), .A2(n5583), .A3(n11320), .A4(n5581), .ZN(
        n17297) );
  NAND2_X1 U17430 ( .A1(n5582), .A2(n13629), .ZN(n5581) );
  INV_X1 U17431 ( .A(n39208), .ZN(n38951) );
  NAND3_X1 U17432 ( .A1(n5586), .A2(n46730), .A3(n5585), .ZN(n46564) );
  NAND2_X1 U17433 ( .A1(n46554), .A2(n46731), .ZN(n5585) );
  NAND2_X1 U17434 ( .A1(n46735), .A2(n46554), .ZN(n5586) );
  NAND2_X1 U17435 ( .A1(n32209), .A2(n32194), .ZN(n31218) );
  NAND2_X1 U17436 ( .A1(n2326), .A2(n5588), .ZN(n5587) );
  NAND2_X1 U17437 ( .A1(n37645), .A2(n5590), .ZN(n5589) );
  NAND3_X1 U17439 ( .A1(n46812), .A2(n5592), .A3(n46811), .ZN(n46815) );
  NAND2_X1 U17440 ( .A1(n2252), .A2(n47069), .ZN(n46770) );
  NAND3_X1 U17441 ( .A1(n2252), .A2(n51404), .A3(n46823), .ZN(n44105) );
  NAND3_X1 U17442 ( .A1(n5592), .A2(n51292), .A3(n51304), .ZN(n46813) );
  NAND2_X1 U17443 ( .A1(n45172), .A2(n2252), .ZN(n44463) );
  NAND2_X1 U17444 ( .A1(n44462), .A2(n5592), .ZN(n44464) );
  NAND2_X2 U17445 ( .A1(n45182), .A2(n45181), .ZN(n50913) );
  XNOR2_X2 U17446 ( .A(n5788), .B(n35807), .ZN(n39299) );
  NAND3_X2 U17448 ( .A1(n40548), .A2(n5595), .A3(n5594), .ZN(n43781) );
  XNOR2_X1 U17449 ( .A(n5598), .B(n4800), .ZN(n34434) );
  XNOR2_X1 U17450 ( .A(n33967), .B(n5598), .ZN(n34288) );
  NAND2_X1 U17451 ( .A1(n29759), .A2(n29760), .ZN(n29761) );
  NAND2_X1 U17452 ( .A1(n17440), .A2(n17553), .ZN(n18327) );
  OAI21_X1 U17453 ( .B1(n18064), .B2(n17436), .A(n5600), .ZN(n5602) );
  NAND2_X1 U17454 ( .A1(n17440), .A2(n5601), .ZN(n5600) );
  NOR2_X1 U17455 ( .A1(n17544), .A2(n18063), .ZN(n5601) );
  NAND2_X1 U17457 ( .A1(n38817), .A2(n41792), .ZN(n5604) );
  NAND2_X1 U17458 ( .A1(n20122), .A2(n20166), .ZN(n19542) );
  NOR2_X1 U17459 ( .A1(n5607), .A2(n5606), .ZN(n5605) );
  OAI21_X1 U17460 ( .B1(n37498), .B2(n37747), .A(n36242), .ZN(n5606) );
  AOI21_X1 U17461 ( .B1(n37763), .B2(n2243), .A(n36251), .ZN(n5607) );
  NAND2_X1 U17462 ( .A1(n37501), .A2(n37745), .ZN(n37498) );
  INV_X1 U17463 ( .A(n22586), .ZN(n5609) );
  NAND2_X1 U17464 ( .A1(n5609), .A2(n20903), .ZN(n5610) );
  XNOR2_X1 U17465 ( .A(n5611), .B(n17831), .ZN(n17382) );
  XNOR2_X1 U17466 ( .A(n5611), .B(n15738), .ZN(n15409) );
  XNOR2_X1 U17467 ( .A(n5611), .B(n18593), .ZN(n18594) );
  NAND3_X1 U17468 ( .A1(n20105), .A2(n17057), .A3(n778), .ZN(n16790) );
  XNOR2_X1 U17469 ( .A(n34608), .B(n5612), .ZN(n5648) );
  XNOR2_X1 U17470 ( .A(n33303), .B(n5612), .ZN(n34421) );
  XNOR2_X1 U17471 ( .A(n35752), .B(n5612), .ZN(n37307) );
  XNOR2_X1 U17472 ( .A(n5616), .B(n35273), .ZN(n35274) );
  XNOR2_X1 U17473 ( .A(n5616), .B(n37317), .ZN(n37321) );
  XNOR2_X1 U17474 ( .A(n35482), .B(n5616), .ZN(n33942) );
  NAND2_X1 U17475 ( .A1(n26985), .A2(n2424), .ZN(n29431) );
  INV_X1 U17476 ( .A(n37484), .ZN(n37490) );
  NAND3_X1 U17477 ( .A1(n658), .A2(n5617), .A3(n50280), .ZN(n50283) );
  NAND2_X1 U17478 ( .A1(n44001), .A2(n47044), .ZN(n50261) );
  NAND2_X1 U17481 ( .A1(n6384), .A2(n15163), .ZN(n14573) );
  NAND2_X1 U17482 ( .A1(n10862), .A2(n5622), .ZN(n5621) );
  INV_X1 U17484 ( .A(n22654), .ZN(n21852) );
  NAND2_X1 U17485 ( .A1(n8409), .A2(n21232), .ZN(n5624) );
  NAND4_X2 U17486 ( .A1(n19107), .A2(n5627), .A3(n19106), .A4(n19105), .ZN(
        n23247) );
  AOI22_X1 U17487 ( .A1(n19090), .A2(n19099), .B1(n19091), .B2(n19092), .ZN(
        n5627) );
  NAND3_X1 U17488 ( .A1(n5629), .A2(n14967), .A3(n10766), .ZN(n5628) );
  OAI21_X1 U17489 ( .B1(n14156), .B2(n14164), .A(n14150), .ZN(n5629) );
  NAND3_X1 U17490 ( .A1(n14455), .A2(n14441), .A3(n51383), .ZN(n11430) );
  NAND2_X1 U17491 ( .A1(n29841), .A2(n31497), .ZN(n30999) );
  NAND3_X1 U17492 ( .A1(n722), .A2(n29841), .A3(n5631), .ZN(n31276) );
  OR2_X2 U17493 ( .A1(n5632), .A2(n32783), .ZN(n36931) );
  OR2_X2 U17494 ( .A1(n5633), .A2(n7736), .ZN(n33911) );
  NAND2_X1 U17497 ( .A1(n37496), .A2(n37759), .ZN(n37751) );
  NAND3_X1 U17498 ( .A1(n29992), .A2(n29991), .A3(n31425), .ZN(n31426) );
  NAND2_X1 U17499 ( .A1(n41008), .A2(n39576), .ZN(n39575) );
  NAND2_X1 U17500 ( .A1(n5639), .A2(n30712), .ZN(n5638) );
  INV_X1 U17501 ( .A(n30707), .ZN(n5639) );
  INV_X1 U17502 ( .A(n30722), .ZN(n28807) );
  OAI22_X1 U17503 ( .A1(n28808), .A2(n5641), .B1(n30707), .B2(n30722), .ZN(
        n5640) );
  NAND2_X1 U17504 ( .A1(n28810), .A2(n52218), .ZN(n5641) );
  NAND3_X1 U17505 ( .A1(n5878), .A2(n23027), .A3(n23998), .ZN(n5642) );
  NAND2_X1 U17506 ( .A1(n5643), .A2(n11037), .ZN(n11038) );
  NAND2_X1 U17507 ( .A1(n5644), .A2(n2197), .ZN(n9825) );
  NOR2_X1 U17508 ( .A1(n22426), .A2(n23983), .ZN(n23029) );
  NAND4_X2 U17509 ( .A1(n19181), .A2(n5646), .A3(n19179), .A4(n7234), .ZN(
        n24000) );
  NAND2_X1 U17511 ( .A1(n49003), .A2(n49008), .ZN(n49031) );
  NOR2_X1 U17512 ( .A1(n23536), .A2(n23535), .ZN(n5649) );
  NAND2_X1 U17513 ( .A1(n2253), .A2(n11813), .ZN(n7887) );
  NAND2_X1 U17514 ( .A1(n5651), .A2(n14451), .ZN(n14460) );
  NAND2_X1 U17515 ( .A1(n5652), .A2(n11813), .ZN(n5651) );
  AND2_X1 U17516 ( .A1(n21219), .A2(n5653), .ZN(n5655) );
  NAND2_X1 U17517 ( .A1(n2456), .A2(n6476), .ZN(n5653) );
  INV_X1 U17518 ( .A(n11640), .ZN(n9302) );
  NAND2_X1 U17519 ( .A1(n9509), .A2(n11660), .ZN(n5657) );
  NOR2_X1 U17520 ( .A1(n49127), .A2(n49112), .ZN(n49065) );
  INV_X1 U17521 ( .A(n5660), .ZN(n44797) );
  OAI21_X1 U17522 ( .B1(n7518), .B2(n49085), .A(n49057), .ZN(n5660) );
  NAND2_X1 U17526 ( .A1(n40438), .A2(n5664), .ZN(n40441) );
  INV_X1 U17527 ( .A(n51520), .ZN(n32074) );
  NOR2_X1 U17528 ( .A1(n51520), .A2(n5665), .ZN(n31285) );
  NAND2_X1 U17531 ( .A1(n46290), .A2(n45937), .ZN(n49138) );
  NAND2_X1 U17532 ( .A1(n46290), .A2(n51017), .ZN(n44730) );
  OAI21_X1 U17533 ( .B1(n43421), .B2(n49148), .A(n51017), .ZN(n45942) );
  NAND2_X1 U17534 ( .A1(n49150), .A2(n51016), .ZN(n46283) );
  NAND2_X1 U17535 ( .A1(n49142), .A2(n51016), .ZN(n49143) );
  XNOR2_X1 U17536 ( .A(n51668), .B(n5670), .ZN(n15355) );
  XNOR2_X1 U17537 ( .A(n18148), .B(n5670), .ZN(n17332) );
  XNOR2_X1 U17538 ( .A(n18414), .B(n5670), .ZN(n15468) );
  XNOR2_X1 U17539 ( .A(n16953), .B(n5670), .ZN(n15668) );
  XNOR2_X1 U17540 ( .A(n5670), .B(n18507), .ZN(n17236) );
  INV_X1 U17542 ( .A(n18040), .ZN(n5671) );
  NAND2_X1 U17543 ( .A1(n5674), .A2(n5673), .ZN(n6138) );
  NAND3_X1 U17544 ( .A1(n36285), .A2(n42042), .A3(n42049), .ZN(n5674) );
  XNOR2_X1 U17545 ( .A(n43954), .B(n4649), .ZN(n41859) );
  XNOR2_X1 U17546 ( .A(n43954), .B(n2185), .ZN(n46131) );
  XNOR2_X1 U17547 ( .A(n5677), .B(n5676), .ZN(n26306) );
  XNOR2_X1 U17548 ( .A(n27430), .B(n26283), .ZN(n5676) );
  XNOR2_X1 U17549 ( .A(n26278), .B(n26273), .ZN(n5679) );
  XNOR2_X1 U17550 ( .A(n34726), .B(n51662), .ZN(n34736) );
  NAND3_X1 U17551 ( .A1(n29607), .A2(n29608), .A3(n5681), .ZN(n5680) );
  NAND2_X1 U17552 ( .A1(n2462), .A2(n51744), .ZN(n5681) );
  NAND2_X1 U17553 ( .A1(n21714), .A2(n5683), .ZN(n19914) );
  NAND2_X1 U17554 ( .A1(n463), .A2(n5683), .ZN(n19916) );
  NOR2_X1 U17555 ( .A1(n21712), .A2(n5683), .ZN(n21711) );
  NAND2_X1 U17556 ( .A1(n22183), .A2(n5683), .ZN(n21110) );
  XNOR2_X1 U17557 ( .A(n35619), .B(n5686), .ZN(n35620) );
  XNOR2_X1 U17558 ( .A(n34759), .B(n5686), .ZN(n34769) );
  XNOR2_X1 U17559 ( .A(n34862), .B(n5686), .ZN(n34863) );
  XNOR2_X1 U17560 ( .A(n33705), .B(n5686), .ZN(n33706) );
  XNOR2_X1 U17561 ( .A(n5686), .B(n33616), .ZN(n33619) );
  OAI21_X1 U17562 ( .B1(n30221), .B2(n27937), .A(n29261), .ZN(n27939) );
  NAND2_X1 U17563 ( .A1(n12055), .A2(n7019), .ZN(n10355) );
  NAND2_X1 U17564 ( .A1(n12058), .A2(n5687), .ZN(n8712) );
  NAND2_X1 U17565 ( .A1(n10354), .A2(n5687), .ZN(n10358) );
  NOR2_X1 U17566 ( .A1(n8349), .A2(n5687), .ZN(n9219) );
  INV_X1 U17567 ( .A(n45641), .ZN(n5692) );
  AND2_X1 U17568 ( .A1(n5693), .A2(n28862), .ZN(n28962) );
  NAND2_X1 U17569 ( .A1(n28951), .A2(n5056), .ZN(n28505) );
  NAND2_X1 U17570 ( .A1(n28867), .A2(n5693), .ZN(n29789) );
  NAND2_X1 U17571 ( .A1(n28951), .A2(n5693), .ZN(n28501) );
  OAI21_X1 U17572 ( .B1(n28952), .B2(n52251), .A(n29790), .ZN(n28459) );
  NAND2_X1 U17574 ( .A1(n18877), .A2(n5694), .ZN(n18878) );
  INV_X1 U17575 ( .A(n29565), .ZN(n5696) );
  NAND2_X1 U17576 ( .A1(n5697), .A2(n29563), .ZN(n29565) );
  AND2_X1 U17577 ( .A1(n26197), .A2(n29550), .ZN(n5697) );
  NAND2_X1 U17578 ( .A1(n30085), .A2(n5698), .ZN(n29644) );
  OAI211_X1 U17579 ( .C1(n23667), .C2(n7494), .A(n23666), .B(n5701), .ZN(n5703) );
  NAND4_X2 U17580 ( .A1(n5702), .A2(n23678), .A3(n23676), .A4(n23677), .ZN(
        n28048) );
  NAND2_X1 U17581 ( .A1(n28601), .A2(n30143), .ZN(n5704) );
  NAND4_X2 U17582 ( .A1(n5707), .A2(n29582), .A3(n29580), .A4(n29581), .ZN(
        n37066) );
  NAND2_X1 U17583 ( .A1(n29576), .A2(n7978), .ZN(n5707) );
  AOI21_X1 U17584 ( .B1(n7084), .B2(n48915), .A(n5709), .ZN(n5708) );
  NAND2_X1 U17585 ( .A1(n48882), .A2(n48908), .ZN(n48887) );
  NAND2_X1 U17586 ( .A1(n36080), .A2(n5710), .ZN(n34982) );
  NAND2_X1 U17587 ( .A1(n37988), .A2(n36518), .ZN(n37981) );
  XNOR2_X1 U17588 ( .A(n25860), .B(n33407), .ZN(n25181) );
  XNOR2_X1 U17589 ( .A(n51523), .B(n51484), .ZN(n22400) );
  XNOR2_X1 U17590 ( .A(n51523), .B(n28343), .ZN(n28344) );
  NAND2_X1 U17592 ( .A1(n51723), .A2(n30788), .ZN(n30785) );
  NAND2_X1 U17593 ( .A1(n29892), .A2(n30790), .ZN(n23661) );
  NAND2_X1 U17594 ( .A1(n20317), .A2(n5716), .ZN(n20492) );
  XNOR2_X1 U17595 ( .A(n37080), .B(n7610), .ZN(n5717) );
  NAND2_X1 U17596 ( .A1(n31379), .A2(n3241), .ZN(n5721) );
  OR2_X1 U17597 ( .A1(n30528), .A2(n3241), .ZN(n5720) );
  OAI211_X1 U17598 ( .C1(n22210), .C2(n22209), .A(n23092), .B(n5723), .ZN(
        n22216) );
  XNOR2_X1 U17599 ( .A(n41569), .B(n5724), .ZN(n41570) );
  XNOR2_X1 U17600 ( .A(n51409), .B(n5724), .ZN(n41251) );
  XNOR2_X1 U17601 ( .A(n42517), .B(n52038), .ZN(n42518) );
  XNOR2_X1 U17602 ( .A(n5724), .B(n43524), .ZN(n42955) );
  XNOR2_X1 U17604 ( .A(n7351), .B(n5725), .ZN(n25091) );
  XNOR2_X1 U17605 ( .A(n7351), .B(n2542), .ZN(n17995) );
  INV_X1 U17606 ( .A(n7351), .ZN(n5726) );
  NAND4_X2 U17607 ( .A1(n5807), .A2(n5728), .A3(n37395), .A4(n5727), .ZN(
        n40785) );
  NAND2_X1 U17608 ( .A1(n37525), .A2(n37388), .ZN(n5727) );
  NOR2_X1 U17609 ( .A1(n2372), .A2(n5729), .ZN(n5728) );
  NAND2_X1 U17610 ( .A1(n37386), .A2(n37392), .ZN(n37525) );
  NAND2_X1 U17611 ( .A1(n10039), .A2(n2538), .ZN(n5731) );
  OAI21_X1 U17612 ( .B1(n13296), .B2(n13729), .A(n469), .ZN(n5734) );
  OAI21_X1 U17613 ( .B1(n5735), .B2(n17987), .A(n22907), .ZN(n17988) );
  INV_X1 U17614 ( .A(n6094), .ZN(n5735) );
  NAND2_X1 U17615 ( .A1(n5736), .A2(n5542), .ZN(n6094) );
  NOR2_X1 U17616 ( .A1(n5740), .A2(n5739), .ZN(n5738) );
  AOI21_X1 U17617 ( .B1(n35896), .B2(n35895), .A(n5741), .ZN(n5740) );
  NAND2_X1 U17618 ( .A1(n10554), .A2(n9830), .ZN(n9826) );
  NAND2_X1 U17619 ( .A1(n31197), .A2(n31198), .ZN(n5745) );
  INV_X1 U17620 ( .A(n5747), .ZN(n40872) );
  OAI21_X1 U17621 ( .B1(n40861), .B2(n40543), .A(n5747), .ZN(n39749) );
  NAND2_X1 U17622 ( .A1(n18246), .A2(n19891), .ZN(n5748) );
  OAI211_X1 U17623 ( .C1(n32492), .C2(n32491), .A(n32490), .B(n5752), .ZN(
        n5751) );
  AOI22_X1 U17624 ( .A1(n3664), .A2(n32489), .B1(n32487), .B2(n32488), .ZN(
        n5752) );
  AND3_X1 U17625 ( .A1(n5755), .A2(n32493), .A3(n5754), .ZN(n5753) );
  NAND2_X1 U17626 ( .A1(n32482), .A2(n32483), .ZN(n5754) );
  NAND3_X1 U17627 ( .A1(n32481), .A2(n5756), .A3(n32478), .ZN(n5755) );
  INV_X1 U17628 ( .A(n32480), .ZN(n5756) );
  NAND3_X1 U17629 ( .A1(n29855), .A2(n731), .A3(n30723), .ZN(n27590) );
  NAND4_X2 U17630 ( .A1(n5758), .A2(n46031), .A3(n5760), .A4(n5757), .ZN(
        n49899) );
  NAND2_X1 U17631 ( .A1(n5762), .A2(n49652), .ZN(n5757) );
  NAND3_X1 U17632 ( .A1(n5759), .A2(n51733), .A3(n46027), .ZN(n5758) );
  NAND2_X1 U17633 ( .A1(n49660), .A2(n49659), .ZN(n5759) );
  NOR2_X1 U17634 ( .A1(n2350), .A2(n5761), .ZN(n5760) );
  XNOR2_X1 U17635 ( .A(n52211), .B(n46028), .ZN(n5763) );
  NAND2_X1 U17636 ( .A1(n27563), .A2(n5769), .ZN(n5767) );
  NAND2_X1 U17637 ( .A1(n17456), .A2(n18374), .ZN(n20039) );
  INV_X1 U17638 ( .A(n5771), .ZN(n5770) );
  XNOR2_X1 U17640 ( .A(n49511), .B(n49510), .ZN(n5772) );
  NOR2_X1 U17641 ( .A1(n10848), .A2(n5773), .ZN(n6250) );
  OAI211_X1 U17642 ( .C1(n11467), .C2(n11628), .A(n10847), .B(n5774), .ZN(
        n5773) );
  NAND3_X1 U17643 ( .A1(n11464), .A2(n10852), .A3(n11460), .ZN(n5774) );
  NAND2_X1 U17644 ( .A1(n30768), .A2(n30757), .ZN(n27560) );
  XNOR2_X1 U17646 ( .A(n41656), .B(n52068), .ZN(n46109) );
  XNOR2_X1 U17647 ( .A(n5775), .B(n42340), .ZN(n42341) );
  XNOR2_X1 U17648 ( .A(n44007), .B(n5775), .ZN(n44008) );
  XNOR2_X1 U17649 ( .A(n5775), .B(n43124), .ZN(n43125) );
  XNOR2_X1 U17650 ( .A(n43551), .B(n52068), .ZN(n43557) );
  XNOR2_X1 U17651 ( .A(n42454), .B(n52068), .ZN(n42456) );
  NOR2_X1 U17653 ( .A1(n2348), .A2(n5776), .ZN(n12347) );
  XNOR2_X1 U17654 ( .A(n5777), .B(n35237), .ZN(n33989) );
  XNOR2_X1 U17655 ( .A(n5777), .B(n33217), .ZN(n33219) );
  XNOR2_X1 U17656 ( .A(n5777), .B(n35075), .ZN(n32934) );
  OR2_X1 U17657 ( .A1(n31950), .A2(n32409), .ZN(n5780) );
  NAND2_X1 U17658 ( .A1(n29157), .A2(n5781), .ZN(n29161) );
  NAND2_X1 U17659 ( .A1(n49273), .A2(n46199), .ZN(n45679) );
  NAND2_X1 U17660 ( .A1(n49274), .A2(n5783), .ZN(n46199) );
  NAND2_X1 U17661 ( .A1(n5784), .A2(n51418), .ZN(n37396) );
  XNOR2_X1 U17662 ( .A(n33603), .B(n51381), .ZN(n33650) );
  INV_X1 U17663 ( .A(n38722), .ZN(n38727) );
  XNOR2_X1 U17664 ( .A(n5785), .B(n4823), .ZN(n22452) );
  XNOR2_X1 U17665 ( .A(n5785), .B(n25869), .ZN(n25870) );
  XNOR2_X2 U17666 ( .A(n5785), .B(n26159), .ZN(n27242) );
  XNOR2_X1 U17667 ( .A(n25755), .B(n5785), .ZN(n25756) );
  NAND2_X1 U17669 ( .A1(n5787), .A2(n51302), .ZN(n47539) );
  INV_X1 U17670 ( .A(n47547), .ZN(n47571) );
  NAND4_X2 U17671 ( .A1(n5790), .A2(n5795), .A3(n5794), .A4(n5789), .ZN(n31608) );
  NAND2_X1 U17672 ( .A1(n29231), .A2(n29223), .ZN(n5789) );
  NAND2_X1 U17673 ( .A1(n29231), .A2(n29232), .ZN(n5791) );
  NAND2_X1 U17674 ( .A1(n29244), .A2(n29243), .ZN(n5793) );
  INV_X1 U17675 ( .A(n47110), .ZN(n46881) );
  NAND2_X1 U17676 ( .A1(n46881), .A2(n46720), .ZN(n46724) );
  INV_X1 U17677 ( .A(n5796), .ZN(n7475) );
  NAND2_X1 U17678 ( .A1(n27040), .A2(n2213), .ZN(n5796) );
  NOR2_X1 U17679 ( .A1(n5796), .A2(n6303), .ZN(n27037) );
  INV_X1 U17680 ( .A(n37659), .ZN(n38724) );
  NAND2_X1 U17681 ( .A1(n2436), .A2(n37659), .ZN(n38321) );
  NAND2_X1 U17682 ( .A1(n40526), .A2(n40869), .ZN(n40529) );
  NAND3_X1 U17683 ( .A1(n40526), .A2(n40869), .A3(n40525), .ZN(n40534) );
  OAI21_X1 U17684 ( .B1(n39747), .B2(n40868), .A(n40859), .ZN(n38357) );
  NAND3_X1 U17685 ( .A1(n5798), .A2(n5797), .A3(n50194), .ZN(n50202) );
  INV_X1 U17686 ( .A(n7201), .ZN(n5799) );
  NAND2_X1 U17687 ( .A1(n24043), .A2(n23394), .ZN(n5802) );
  NAND2_X1 U17689 ( .A1(n40785), .A2(n40778), .ZN(n40591) );
  NAND3_X1 U17691 ( .A1(n37390), .A2(n37391), .A3(n5808), .ZN(n5807) );
  NOR2_X1 U17692 ( .A1(n5812), .A2(n42054), .ZN(n8500) );
  OAI22_X1 U17693 ( .A1(n5813), .A2(n51208), .B1(n17496), .B2(n2166), .ZN(
        n6951) );
  NAND2_X1 U17695 ( .A1(n49619), .A2(n7798), .ZN(n5815) );
  NAND2_X1 U17696 ( .A1(n30633), .A2(n31368), .ZN(n5819) );
  NAND3_X1 U17697 ( .A1(n32294), .A2(n386), .A3(n32300), .ZN(n5820) );
  NAND2_X1 U17698 ( .A1(n27951), .A2(n29174), .ZN(n5822) );
  NAND3_X1 U17699 ( .A1(n27951), .A2(n29174), .A3(n5821), .ZN(n27959) );
  NAND2_X1 U17700 ( .A1(n5822), .A2(n29172), .ZN(n29176) );
  NAND2_X1 U17701 ( .A1(n5823), .A2(n42089), .ZN(n42088) );
  AND2_X1 U17702 ( .A1(n42086), .A2(n5824), .ZN(n5823) );
  NAND4_X1 U17703 ( .A1(n7647), .A2(n42089), .A3(n42093), .A4(n5824), .ZN(
        n42090) );
  NAND3_X1 U17704 ( .A1(n5825), .A2(n14223), .A3(n14233), .ZN(n12931) );
  NAND2_X1 U17705 ( .A1(n12922), .A2(n13970), .ZN(n5825) );
  OR2_X1 U17707 ( .A1(n27827), .A2(n26722), .ZN(n27024) );
  NOR2_X1 U17709 ( .A1(n11186), .A2(n11582), .ZN(n5827) );
  AND2_X1 U17710 ( .A1(n11186), .A2(n11530), .ZN(n12559) );
  AND2_X1 U17712 ( .A1(n39027), .A2(n467), .ZN(n7815) );
  XNOR2_X2 U17713 ( .A(n34786), .B(n34785), .ZN(n39464) );
  INV_X1 U17714 ( .A(n39028), .ZN(n34806) );
  NAND2_X1 U17715 ( .A1(n5829), .A2(n21958), .ZN(n21959) );
  NAND2_X1 U17717 ( .A1(n23147), .A2(n51123), .ZN(n5829) );
  NAND2_X1 U17718 ( .A1(n12923), .A2(n5540), .ZN(n5830) );
  NAND4_X2 U17719 ( .A1(n9778), .A2(n9776), .A3(n9777), .A4(n9775), .ZN(n13968) );
  OR2_X1 U17720 ( .A1(n21024), .A2(n975), .ZN(n17615) );
  INV_X1 U17721 ( .A(n21024), .ZN(n5833) );
  NAND2_X1 U17724 ( .A1(n5836), .A2(n50612), .ZN(n5835) );
  NAND2_X1 U17725 ( .A1(n50610), .A2(n50609), .ZN(n5836) );
  NAND2_X1 U17726 ( .A1(n30383), .A2(n30382), .ZN(n5840) );
  NAND2_X1 U17727 ( .A1(n5843), .A2(n30371), .ZN(n5842) );
  OAI211_X1 U17729 ( .C1(n46894), .C2(n43683), .A(n45158), .B(n47000), .ZN(
        n5850) );
  NAND2_X1 U17730 ( .A1(n43685), .A2(n47003), .ZN(n5851) );
  NAND3_X1 U17731 ( .A1(n44473), .A2(n45153), .A3(n47150), .ZN(n5852) );
  NAND2_X1 U17732 ( .A1(n19044), .A2(n20122), .ZN(n5854) );
  NAND3_X2 U17733 ( .A1(n7388), .A2(n39392), .A3(n39391), .ZN(n42006) );
  XNOR2_X1 U17734 ( .A(n23043), .B(n5855), .ZN(n7012) );
  XNOR2_X1 U17735 ( .A(n24526), .B(n5855), .ZN(n7801) );
  XNOR2_X1 U17736 ( .A(n5855), .B(n42769), .ZN(n25122) );
  XNOR2_X1 U17737 ( .A(n5855), .B(n27234), .ZN(n24263) );
  XNOR2_X1 U17738 ( .A(n5855), .B(n27362), .ZN(n25954) );
  XNOR2_X1 U17739 ( .A(n51056), .B(n5855), .ZN(n27482) );
  XNOR2_X2 U17740 ( .A(n24891), .B(n28038), .ZN(n5855) );
  INV_X1 U17741 ( .A(n18055), .ZN(n5856) );
  NAND2_X1 U17742 ( .A1(n5858), .A2(n47899), .ZN(n5857) );
  INV_X1 U17743 ( .A(n47925), .ZN(n5858) );
  OAI21_X1 U17744 ( .B1(n40732), .B2(n52215), .A(n40372), .ZN(n38607) );
  INV_X1 U17748 ( .A(n39192), .ZN(n39379) );
  NAND2_X1 U17749 ( .A1(n37031), .A2(n51102), .ZN(n39192) );
  NAND4_X2 U17750 ( .A1(n7395), .A2(n5863), .A3(n31551), .A4(n31552), .ZN(
        n35841) );
  NAND2_X1 U17751 ( .A1(n5868), .A2(n31538), .ZN(n31448) );
  NAND2_X1 U17752 ( .A1(n5866), .A2(n32665), .ZN(n31170) );
  NAND2_X1 U17753 ( .A1(n5867), .A2(n31452), .ZN(n5866) );
  NAND3_X1 U17754 ( .A1(n381), .A2(n31546), .A3(n5868), .ZN(n31179) );
  MUX2_X1 U17755 ( .A(n31441), .B(n31442), .S(n31452), .Z(n31460) );
  NAND2_X1 U17757 ( .A1(n18299), .A2(n19491), .ZN(n5869) );
  NAND2_X1 U17758 ( .A1(n18308), .A2(n18307), .ZN(n5870) );
  NAND3_X1 U17759 ( .A1(n20079), .A2(n20078), .A3(n20082), .ZN(n5871) );
  OR2_X2 U17760 ( .A1(n5872), .A2(n38006), .ZN(n6541) );
  INV_X1 U17761 ( .A(n32678), .ZN(n5872) );
  INV_X1 U17762 ( .A(n38006), .ZN(n38002) );
  INV_X2 U17763 ( .A(n41058), .ZN(n41065) );
  NAND2_X1 U17764 ( .A1(n41063), .A2(n41058), .ZN(n40493) );
  AND2_X2 U17765 ( .A1(n5873), .A2(n34978), .ZN(n41058) );
  XNOR2_X1 U17767 ( .A(n45415), .B(n5874), .ZN(n43028) );
  XNOR2_X1 U17768 ( .A(n42235), .B(n52145), .ZN(n42236) );
  XNOR2_X1 U17769 ( .A(n43710), .B(n5874), .ZN(n42578) );
  XNOR2_X1 U17770 ( .A(n45269), .B(n5874), .ZN(n45276) );
  XNOR2_X1 U17771 ( .A(n43027), .B(n52145), .ZN(n44529) );
  XNOR2_X1 U17772 ( .A(n42645), .B(n52145), .ZN(n43303) );
  INV_X1 U17775 ( .A(n20428), .ZN(n5875) );
  NAND2_X1 U17776 ( .A1(n20426), .A2(n6454), .ZN(n17859) );
  NAND2_X1 U17777 ( .A1(n20423), .A2(n6454), .ZN(n20347) );
  INV_X1 U17778 ( .A(n33648), .ZN(n5876) );
  INV_X1 U17781 ( .A(n44254), .ZN(n5877) );
  NAND2_X1 U17782 ( .A1(n23989), .A2(n24002), .ZN(n5878) );
  NAND2_X1 U17783 ( .A1(n23983), .A2(n22426), .ZN(n23989) );
  INV_X1 U17784 ( .A(n23989), .ZN(n22534) );
  NAND2_X1 U17785 ( .A1(n17050), .A2(n17458), .ZN(n5879) );
  NAND2_X1 U17786 ( .A1(n20046), .A2(n5881), .ZN(n5880) );
  NAND3_X1 U17788 ( .A1(n28142), .A2(n7888), .A3(n28511), .ZN(n5931) );
  NAND3_X1 U17790 ( .A1(n51348), .A2(n41065), .A3(n40500), .ZN(n5884) );
  OAI21_X1 U17791 ( .B1(n41046), .B2(n41057), .A(n5884), .ZN(n41050) );
  XNOR2_X2 U17792 ( .A(n5885), .B(n46077), .ZN(n46267) );
  XNOR2_X1 U17793 ( .A(n42796), .B(n42527), .ZN(n5885) );
  AND2_X1 U17795 ( .A1(n48884), .A2(n48876), .ZN(n5888) );
  NAND2_X1 U17797 ( .A1(n38767), .A2(n38766), .ZN(n5894) );
  INV_X1 U17798 ( .A(n44327), .ZN(n5891) );
  NOR2_X1 U17799 ( .A1(n5894), .A2(n5893), .ZN(n5892) );
  NOR2_X1 U17800 ( .A1(n38768), .A2(n2344), .ZN(n5895) );
  NAND2_X1 U17801 ( .A1(n7519), .A2(n5897), .ZN(n5896) );
  NAND3_X1 U17802 ( .A1(n23513), .A2(n52207), .A3(n24292), .ZN(n5898) );
  NAND4_X1 U17803 ( .A1(n40193), .A2(n40195), .A3(n40200), .A4(n40194), .ZN(
        n5901) );
  NAND2_X1 U17804 ( .A1(n40197), .A2(n5901), .ZN(n5900) );
  NAND2_X1 U17806 ( .A1(n17418), .A2(n23068), .ZN(n23595) );
  NAND2_X1 U17807 ( .A1(n5905), .A2(n13820), .ZN(n5903) );
  OAI22_X1 U17809 ( .A1(n11794), .A2(n14321), .B1(n13826), .B2(n13045), .ZN(
        n5905) );
  NAND2_X1 U17810 ( .A1(n11795), .A2(n14307), .ZN(n5907) );
  OAI21_X1 U17811 ( .B1(n11797), .B2(n13827), .A(n13600), .ZN(n5908) );
  NOR2_X1 U17813 ( .A1(n51126), .A2(n19047), .ZN(n16491) );
  XNOR2_X1 U17814 ( .A(n33343), .B(n34572), .ZN(n30887) );
  NAND2_X1 U17815 ( .A1(n6271), .A2(n31603), .ZN(n5914) );
  NAND2_X1 U17816 ( .A1(n11648), .A2(n9507), .ZN(n11651) );
  NAND2_X1 U17817 ( .A1(n5915), .A2(n11662), .ZN(n9513) );
  INV_X1 U17819 ( .A(n11649), .ZN(n5917) );
  NAND2_X1 U17821 ( .A1(n17984), .A2(n5922), .ZN(n5921) );
  NOR2_X1 U17822 ( .A1(n5924), .A2(n2199), .ZN(n49738) );
  NAND2_X1 U17823 ( .A1(n5924), .A2(n2198), .ZN(n50375) );
  XNOR2_X2 U17825 ( .A(n46057), .B(n46056), .ZN(n5924) );
  OR2_X1 U17826 ( .A1(n50034), .A2(n50386), .ZN(n47316) );
  NAND2_X1 U17827 ( .A1(n50034), .A2(n50386), .ZN(n49732) );
  AND2_X1 U17828 ( .A1(n5924), .A2(n49730), .ZN(n47015) );
  NAND2_X1 U17829 ( .A1(n49740), .A2(n5924), .ZN(n50389) );
  NAND4_X1 U17830 ( .A1(n50377), .A2(n50387), .A3(n51058), .A4(n5924), .ZN(
        n49734) );
  NAND2_X1 U17831 ( .A1(n5925), .A2(n51713), .ZN(n13367) );
  NAND3_X1 U17833 ( .A1(n10291), .A2(n10278), .A3(n5930), .ZN(n5929) );
  INV_X1 U17834 ( .A(n28947), .ZN(n28958) );
  NAND2_X1 U17835 ( .A1(n28867), .A2(n28862), .ZN(n28947) );
  NAND2_X1 U17836 ( .A1(n37806), .A2(n39472), .ZN(n36214) );
  NAND2_X1 U17837 ( .A1(n37806), .A2(n37802), .ZN(n34701) );
  NAND2_X1 U17838 ( .A1(n37806), .A2(n39474), .ZN(n7198) );
  NAND2_X1 U17839 ( .A1(n7197), .A2(n37806), .ZN(n7196) );
  NAND3_X1 U17841 ( .A1(n2475), .A2(n18933), .A3(n18932), .ZN(n18934) );
  NAND2_X1 U17842 ( .A1(n49522), .A2(n2192), .ZN(n45024) );
  OAI21_X1 U17843 ( .B1(n39065), .B2(n5943), .A(n41487), .ZN(n7417) );
  NOR2_X1 U17844 ( .A1(n6138), .A2(n5943), .ZN(n36290) );
  NAND3_X1 U17845 ( .A1(n5945), .A2(n29750), .A3(n29751), .ZN(n5944) );
  NAND3_X1 U17846 ( .A1(n30444), .A2(n30448), .A3(n29746), .ZN(n5945) );
  NAND2_X1 U17847 ( .A1(n12339), .A2(n12341), .ZN(n5946) );
  NAND2_X1 U17848 ( .A1(n10285), .A2(n5948), .ZN(n5947) );
  NAND3_X1 U17849 ( .A1(n10282), .A2(n9739), .A3(n12328), .ZN(n5948) );
  NAND4_X2 U17850 ( .A1(n5952), .A2(n23522), .A3(n7731), .A4(n5949), .ZN(
        n28352) );
  NAND2_X1 U17851 ( .A1(n23520), .A2(n5950), .ZN(n5949) );
  MUX2_X1 U17852 ( .A(n19093), .B(n19098), .S(n17076), .Z(n16313) );
  XNOR2_X1 U17854 ( .A(n23938), .B(n5955), .ZN(n5954) );
  XNOR2_X1 U17855 ( .A(n49938), .B(n5957), .ZN(Plaintext[137]) );
  NAND2_X1 U17856 ( .A1(n49935), .A2(n49926), .ZN(n5959) );
  XNOR2_X1 U17857 ( .A(n5961), .B(n671), .ZN(n43050) );
  XNOR2_X1 U17858 ( .A(n46068), .B(n44541), .ZN(n5961) );
  NAND2_X1 U17859 ( .A1(n652), .A2(n49916), .ZN(n7549) );
  XNOR2_X1 U17860 ( .A(n5965), .B(n47680), .ZN(Plaintext[16]) );
  NAND2_X1 U17861 ( .A1(n52041), .A2(n45844), .ZN(n5968) );
  NAND2_X1 U17862 ( .A1(n5971), .A2(n20110), .ZN(n5970) );
  NAND3_X1 U17864 ( .A1(n19545), .A2(n20110), .A3(n20123), .ZN(n5972) );
  NAND2_X1 U17865 ( .A1(n2426), .A2(n19543), .ZN(n5973) );
  NAND2_X1 U17866 ( .A1(n32919), .A2(n5975), .ZN(n28814) );
  NAND3_X1 U17867 ( .A1(n5980), .A2(n6735), .A3(n38545), .ZN(n5979) );
  INV_X1 U17868 ( .A(n19475), .ZN(n21250) );
  INV_X1 U17869 ( .A(n45848), .ZN(n46603) );
  NOR2_X1 U17870 ( .A1(n7703), .A2(n5981), .ZN(n7702) );
  AOI21_X1 U17871 ( .B1(n40650), .B2(n5982), .A(n39768), .ZN(n5981) );
  NAND2_X1 U17872 ( .A1(n41433), .A2(n41435), .ZN(n5982) );
  NAND2_X1 U17873 ( .A1(n5983), .A2(n41442), .ZN(n40650) );
  NAND2_X1 U17875 ( .A1(n5982), .A2(n40650), .ZN(n38916) );
  INV_X1 U17877 ( .A(n41435), .ZN(n5983) );
  XNOR2_X1 U17878 ( .A(n5985), .B(n27462), .ZN(n5984) );
  XNOR2_X1 U17879 ( .A(n27448), .B(n27449), .ZN(n5985) );
  XNOR2_X1 U17880 ( .A(n556), .B(n16142), .ZN(n14835) );
  XNOR2_X1 U17881 ( .A(n16372), .B(n557), .ZN(n16147) );
  XNOR2_X1 U17882 ( .A(n557), .B(n15516), .ZN(n15518) );
  OAI21_X1 U17883 ( .B1(n5986), .B2(n46569), .A(n46571), .ZN(n6585) );
  OAI211_X1 U17884 ( .C1(n5986), .C2(n47106), .A(n45142), .B(n45141), .ZN(
        n45143) );
  NAND2_X1 U17886 ( .A1(n37677), .A2(n5988), .ZN(n5987) );
  AND2_X1 U17887 ( .A1(n47507), .A2(n5991), .ZN(n5993) );
  OAI21_X1 U17888 ( .B1(n13970), .B2(n13219), .A(n16221), .ZN(n6642) );
  INV_X1 U17889 ( .A(n32784), .ZN(n5995) );
  NAND4_X2 U17890 ( .A1(n27520), .A2(n27522), .A3(n27521), .A4(n27519), .ZN(
        n32784) );
  XNOR2_X1 U17891 ( .A(n5996), .B(n15215), .ZN(n15216) );
  XNOR2_X1 U17892 ( .A(n5996), .B(n18425), .ZN(n18426) );
  XNOR2_X1 U17893 ( .A(n17803), .B(n5996), .ZN(n17806) );
  XNOR2_X1 U17894 ( .A(n5996), .B(n16532), .ZN(n16533) );
  INV_X1 U17895 ( .A(n35468), .ZN(n5997) );
  XNOR2_X1 U17896 ( .A(n35749), .B(n5998), .ZN(n36746) );
  XNOR2_X1 U17897 ( .A(n5999), .B(n33145), .ZN(n32583) );
  NAND2_X1 U17898 ( .A1(n23471), .A2(n23470), .ZN(n6002) );
  OAI22_X1 U17900 ( .A1(n10954), .A2(n10955), .B1(n6005), .B2(n10956), .ZN(
        n10958) );
  NAND2_X1 U17901 ( .A1(n10964), .A2(n6003), .ZN(n10128) );
  NOR2_X1 U17902 ( .A1(n6004), .A2(n9859), .ZN(n6003) );
  NAND4_X1 U17903 ( .A1(n9856), .A2(n10957), .A3(n10127), .A4(n6005), .ZN(
        n10129) );
  NOR2_X1 U17904 ( .A1(n6009), .A2(n6008), .ZN(n6007) );
  NAND2_X1 U17905 ( .A1(n6812), .A2(n6813), .ZN(n6008) );
  NAND2_X1 U17906 ( .A1(n42972), .A2(n6810), .ZN(n7793) );
  NAND2_X1 U17907 ( .A1(n45898), .A2(n49184), .ZN(n6810) );
  NAND2_X1 U17908 ( .A1(n32396), .A2(n32066), .ZN(n32394) );
  NAND2_X1 U17909 ( .A1(n23160), .A2(n21948), .ZN(n16688) );
  AND2_X1 U17911 ( .A1(n38277), .A2(n6011), .ZN(n35415) );
  XNOR2_X2 U17912 ( .A(n34523), .B(n34522), .ZN(n37624) );
  XNOR2_X2 U17913 ( .A(n33549), .B(n35482), .ZN(n36766) );
  XNOR2_X1 U17914 ( .A(n51409), .B(n6012), .ZN(n44202) );
  XNOR2_X1 U17915 ( .A(n43197), .B(n6012), .ZN(n38753) );
  XNOR2_X1 U17916 ( .A(n51439), .B(n6012), .ZN(n43812) );
  XNOR2_X1 U17917 ( .A(n46073), .B(n6012), .ZN(n44344) );
  XNOR2_X2 U17918 ( .A(n46059), .B(n44541), .ZN(n6012) );
  NAND2_X1 U17919 ( .A1(n37624), .A2(n38275), .ZN(n35866) );
  XNOR2_X2 U17920 ( .A(n6018), .B(n34490), .ZN(n38275) );
  NAND2_X1 U17922 ( .A1(n47899), .A2(n648), .ZN(n6020) );
  NAND2_X1 U17923 ( .A1(n6023), .A2(n20071), .ZN(n6021) );
  NAND2_X1 U17924 ( .A1(n16212), .A2(n19143), .ZN(n6022) );
  NAND2_X1 U17925 ( .A1(n19135), .A2(n19143), .ZN(n19500) );
  NAND2_X1 U17926 ( .A1(n45669), .A2(n6025), .ZN(n42401) );
  NAND2_X1 U17927 ( .A1(n49277), .A2(n6026), .ZN(n44780) );
  NAND2_X1 U17930 ( .A1(n42403), .A2(n42404), .ZN(n6030) );
  NAND2_X1 U17932 ( .A1(n41082), .A2(n41084), .ZN(n39706) );
  INV_X1 U17933 ( .A(n39706), .ZN(n6032) );
  NAND2_X1 U17934 ( .A1(n39144), .A2(n38878), .ZN(n6033) );
  OR2_X1 U17935 ( .A1(n41082), .A2(n8316), .ZN(n38878) );
  XNOR2_X1 U17936 ( .A(n18450), .B(n18617), .ZN(n14585) );
  NAND3_X1 U17940 ( .A1(n51699), .A2(n15437), .A3(n15434), .ZN(n6038) );
  NAND3_X1 U17942 ( .A1(n6980), .A2(n42205), .A3(n41932), .ZN(n6040) );
  NAND2_X1 U17944 ( .A1(n20827), .A2(n2335), .ZN(n19278) );
  AND2_X2 U17946 ( .A1(n6430), .A2(n19282), .ZN(n24001) );
  NOR2_X1 U17947 ( .A1(n19662), .A2(n19658), .ZN(n6044) );
  NAND2_X1 U17948 ( .A1(n7259), .A2(n19891), .ZN(n19884) );
  AND2_X1 U17950 ( .A1(n431), .A2(n40774), .ZN(n40767) );
  NAND2_X1 U17951 ( .A1(n6045), .A2(n40768), .ZN(n40771) );
  NAND3_X1 U17952 ( .A1(n432), .A2(n40774), .A3(n40775), .ZN(n6045) );
  INV_X1 U17953 ( .A(n40778), .ZN(n6046) );
  NAND2_X1 U17954 ( .A1(n12640), .A2(n12074), .ZN(n6572) );
  NOR2_X1 U17955 ( .A1(n6048), .A2(n30768), .ZN(n7984) );
  NOR2_X1 U17956 ( .A1(n6048), .A2(n30751), .ZN(n29922) );
  INV_X1 U17957 ( .A(n10037), .ZN(n9461) );
  OR2_X2 U17958 ( .A1(n43577), .A2(n50314), .ZN(n49993) );
  XNOR2_X2 U17959 ( .A(n7719), .B(n7720), .ZN(n50314) );
  NAND3_X1 U17960 ( .A1(n6051), .A2(n37520), .A3(n38501), .ZN(n6050) );
  INV_X1 U17961 ( .A(n35950), .ZN(n6051) );
  NAND2_X1 U17962 ( .A1(n37384), .A2(n38496), .ZN(n35950) );
  NAND2_X1 U17963 ( .A1(n22836), .A2(n6052), .ZN(n22838) );
  NAND2_X1 U17964 ( .A1(n22822), .A2(n6053), .ZN(n6052) );
  NAND4_X2 U17965 ( .A1(n10380), .A2(n6054), .A3(n10378), .A4(n10379), .ZN(
        n13797) );
  INV_X1 U17966 ( .A(n29868), .ZN(n29700) );
  OAI211_X1 U17967 ( .C1(n28735), .C2(n30430), .A(n6055), .B(n29862), .ZN(
        n28736) );
  NOR2_X1 U17968 ( .A1(n40123), .A2(n40124), .ZN(n7462) );
  NAND4_X1 U17969 ( .A1(n6058), .A2(n27797), .A3(n51747), .A4(n27800), .ZN(
        n6056) );
  INV_X1 U17970 ( .A(n26314), .ZN(n6057) );
  NAND2_X1 U17971 ( .A1(n20557), .A2(n17420), .ZN(n6063) );
  OAI211_X2 U17972 ( .C1(n31707), .C2(n6066), .A(n31717), .B(n6065), .ZN(
        n34169) );
  INV_X1 U17973 ( .A(n13362), .ZN(n6072) );
  INV_X1 U17974 ( .A(n14536), .ZN(n6070) );
  NAND4_X2 U17975 ( .A1(n12187), .A2(n6068), .A3(n12188), .A4(n6071), .ZN(
        n16294) );
  NAND2_X1 U17976 ( .A1(n14362), .A2(n6072), .ZN(n6071) );
  INV_X1 U17978 ( .A(n51380), .ZN(n28247) );
  XNOR2_X1 U17979 ( .A(n28248), .B(n6076), .ZN(n28263) );
  XNOR2_X1 U17980 ( .A(n51120), .B(n6077), .ZN(n6076) );
  INV_X1 U17981 ( .A(n28246), .ZN(n6077) );
  INV_X1 U17982 ( .A(n25840), .ZN(n6080) );
  XNOR2_X1 U17983 ( .A(n52075), .B(n52058), .ZN(n44287) );
  XNOR2_X1 U17984 ( .A(n52074), .B(n42077), .ZN(n42570) );
  XNOR2_X1 U17985 ( .A(n52074), .B(n44223), .ZN(n44224) );
  XNOR2_X2 U17986 ( .A(n32434), .B(n32433), .ZN(n38006) );
  XNOR2_X2 U17987 ( .A(n26432), .B(n6082), .ZN(n27290) );
  NOR2_X2 U17988 ( .A1(n21917), .A2(n21918), .ZN(n6082) );
  XNOR2_X1 U17989 ( .A(n25673), .B(n2545), .ZN(n23775) );
  XNOR2_X1 U17990 ( .A(n25673), .B(n2544), .ZN(n24944) );
  XNOR2_X1 U17991 ( .A(n6082), .B(n21944), .ZN(n24373) );
  NAND2_X1 U17992 ( .A1(n6083), .A2(n30171), .ZN(n30302) );
  INV_X1 U17993 ( .A(n739), .ZN(n6084) );
  AND2_X1 U17994 ( .A1(n39397), .A2(n38995), .ZN(n6090) );
  NAND3_X1 U17995 ( .A1(n26819), .A2(n26818), .A3(n6092), .ZN(n26820) );
  OR2_X1 U17996 ( .A1(n27691), .A2(n6092), .ZN(n6091) );
  NAND2_X1 U17997 ( .A1(n6093), .A2(n32491), .ZN(n32490) );
  NAND2_X1 U17998 ( .A1(n31205), .A2(n32485), .ZN(n6093) );
  INV_X2 U17999 ( .A(n32472), .ZN(n32025) );
  OAI21_X1 U18000 ( .B1(n41695), .B2(n41621), .A(n41704), .ZN(n41613) );
  OAI211_X1 U18001 ( .C1(n22898), .C2(n22899), .A(n22897), .B(n6094), .ZN(
        n22900) );
  XNOR2_X1 U18002 ( .A(n27420), .B(n2412), .ZN(n6095) );
  XNOR2_X1 U18003 ( .A(n6095), .B(n24402), .ZN(n24406) );
  OAI21_X1 U18004 ( .B1(n46374), .B2(n48550), .A(n6097), .ZN(n6096) );
  INV_X1 U18006 ( .A(n8403), .ZN(n6099) );
  NAND2_X1 U18007 ( .A1(n44844), .A2(n6888), .ZN(n6100) );
  NAND3_X1 U18008 ( .A1(n6104), .A2(n40797), .A3(n40801), .ZN(n38762) );
  INV_X1 U18009 ( .A(n38759), .ZN(n6104) );
  NAND3_X1 U18010 ( .A1(n31042), .A2(n31815), .A3(n6105), .ZN(n31044) );
  NAND2_X1 U18011 ( .A1(n6107), .A2(n31826), .ZN(n30572) );
  NAND2_X1 U18012 ( .A1(n31821), .A2(n6107), .ZN(n31823) );
  NAND4_X1 U18013 ( .A1(n6809), .A2(n31034), .A3(n50986), .A4(n6107), .ZN(
        n31036) );
  NAND3_X1 U18014 ( .A1(n30848), .A2(n31039), .A3(n6107), .ZN(n6324) );
  OAI21_X1 U18015 ( .B1(n6994), .B2(n6109), .A(n6108), .ZN(n6993) );
  NAND2_X1 U18017 ( .A1(n30830), .A2(n31303), .ZN(n6112) );
  NAND2_X2 U18018 ( .A1(n6113), .A2(n7312), .ZN(n31302) );
  NAND2_X1 U18019 ( .A1(n6115), .A2(n40499), .ZN(n6114) );
  NAND2_X1 U18020 ( .A1(n40493), .A2(n41064), .ZN(n6115) );
  NAND3_X1 U18021 ( .A1(n10605), .A2(n10619), .A3(n10606), .ZN(n9873) );
  NAND3_X1 U18023 ( .A1(n39665), .A2(n39666), .A3(n6121), .ZN(n6120) );
  NAND2_X1 U18024 ( .A1(n40000), .A2(n51297), .ZN(n6121) );
  XNOR2_X2 U18025 ( .A(n6123), .B(Key[33]), .ZN(n10552) );
  NAND2_X1 U18026 ( .A1(n39008), .A2(n39269), .ZN(n37198) );
  AND2_X1 U18027 ( .A1(n39258), .A2(n39019), .ZN(n39008) );
  NAND3_X1 U18029 ( .A1(n19681), .A2(n19687), .A3(n19680), .ZN(n19682) );
  NAND2_X2 U18030 ( .A1(n6125), .A2(n43451), .ZN(n49534) );
  NAND2_X1 U18031 ( .A1(n6127), .A2(n43447), .ZN(n6126) );
  NAND2_X1 U18032 ( .A1(n7168), .A2(n2505), .ZN(n6127) );
  MUX2_X1 U18033 ( .A(n26904), .B(n26737), .S(n27706), .Z(n8601) );
  NAND2_X1 U18034 ( .A1(n6130), .A2(n6129), .ZN(n8375) );
  NAND2_X1 U18036 ( .A1(n36448), .A2(n35210), .ZN(n6130) );
  INV_X1 U18037 ( .A(n20132), .ZN(n19066) );
  NOR2_X1 U18038 ( .A1(n20132), .A2(n51756), .ZN(n19075) );
  XNOR2_X1 U18039 ( .A(n6131), .B(n36844), .ZN(n33488) );
  XNOR2_X1 U18040 ( .A(n33472), .B(n34739), .ZN(n6131) );
  NAND2_X1 U18041 ( .A1(n17065), .A2(n51756), .ZN(n20143) );
  INV_X1 U18042 ( .A(n50280), .ZN(n50254) );
  NAND2_X1 U18043 ( .A1(n50269), .A2(n51372), .ZN(n50271) );
  INV_X1 U18044 ( .A(n44118), .ZN(n6132) );
  NAND2_X1 U18045 ( .A1(n23317), .A2(n23316), .ZN(n22249) );
  NAND2_X1 U18046 ( .A1(n29389), .A2(n29390), .ZN(n6135) );
  NAND2_X1 U18047 ( .A1(n51052), .A2(n6136), .ZN(n40031) );
  OR2_X1 U18049 ( .A1(n52134), .A2(n23246), .ZN(n21847) );
  NAND2_X1 U18051 ( .A1(n22340), .A2(n26891), .ZN(n6139) );
  NAND2_X1 U18052 ( .A1(n27641), .A2(n27730), .ZN(n6140) );
  XNOR2_X2 U18053 ( .A(n6141), .B(n19441), .ZN(n27618) );
  NAND2_X1 U18054 ( .A1(n8581), .A2(n29153), .ZN(n8579) );
  NAND2_X1 U18056 ( .A1(n30459), .A2(n51693), .ZN(n29734) );
  INV_X1 U18058 ( .A(n7761), .ZN(n6144) );
  XNOR2_X1 U18059 ( .A(n35805), .B(n35803), .ZN(n6146) );
  NAND2_X1 U18061 ( .A1(n6149), .A2(n38738), .ZN(n6148) );
  INV_X1 U18062 ( .A(n10420), .ZN(n12168) );
  NAND2_X1 U18064 ( .A1(n12167), .A2(n12171), .ZN(n6153) );
  INV_X1 U18065 ( .A(n20656), .ZN(n21656) );
  OAI21_X1 U18066 ( .B1(n20659), .B2(n20650), .A(n21648), .ZN(n20655) );
  NAND3_X2 U18067 ( .A1(n29878), .A2(n6154), .A3(n29879), .ZN(n32439) );
  AND2_X1 U18068 ( .A1(n29876), .A2(n29877), .ZN(n6154) );
  XNOR2_X1 U18069 ( .A(n33104), .B(n2549), .ZN(n35801) );
  NAND2_X1 U18070 ( .A1(n31961), .A2(n32359), .ZN(n6156) );
  INV_X1 U18071 ( .A(n31466), .ZN(n6157) );
  XNOR2_X1 U18072 ( .A(n2305), .B(n23015), .ZN(n6158) );
  NAND2_X1 U18073 ( .A1(n49714), .A2(n6161), .ZN(n6160) );
  NAND2_X1 U18074 ( .A1(n51094), .A2(n6162), .ZN(n6161) );
  NOR2_X1 U18075 ( .A1(n49710), .A2(n42990), .ZN(n6162) );
  NAND2_X1 U18077 ( .A1(n21532), .A2(n6165), .ZN(n6164) );
  INV_X1 U18078 ( .A(n29140), .ZN(n30304) );
  NAND2_X1 U18080 ( .A1(n17496), .A2(n6168), .ZN(n18292) );
  XNOR2_X1 U18081 ( .A(n35389), .B(n37309), .ZN(n6170) );
  NAND2_X1 U18082 ( .A1(n14605), .A2(n14011), .ZN(n10733) );
  NAND4_X2 U18083 ( .A1(n12587), .A2(n12588), .A3(n12585), .A4(n12586), .ZN(
        n17923) );
  XNOR2_X1 U18084 ( .A(n16927), .B(n8033), .ZN(n16928) );
  INV_X1 U18085 ( .A(n8775), .ZN(n7936) );
  XNOR2_X2 U18087 ( .A(n42374), .B(n51338), .ZN(n42788) );
  XNOR2_X2 U18088 ( .A(Key[132]), .B(Ciphertext[89]), .ZN(n11590) );
  AND3_X2 U18090 ( .A1(n11254), .A2(n11253), .A3(n11252), .ZN(n12961) );
  INV_X1 U18091 ( .A(n43401), .ZN(n45943) );
  XNOR2_X1 U18092 ( .A(n2103), .B(n42452), .ZN(n42454) );
  OR2_X2 U18094 ( .A1(n352), .A2(n13683), .ZN(n15106) );
  NAND2_X1 U18096 ( .A1(n45809), .A2(n46740), .ZN(n7867) );
  OAI21_X1 U18097 ( .B1(n50901), .B2(n8294), .A(n50903), .ZN(n50944) );
  INV_X1 U18098 ( .A(n8241), .ZN(n30857) );
  XNOR2_X2 U18099 ( .A(n34219), .B(n37067), .ZN(n34143) );
  XNOR2_X1 U18100 ( .A(n42748), .B(n43297), .ZN(n6846) );
  NAND4_X2 U18101 ( .A1(n14375), .A2(n14376), .A3(n14374), .A4(n14373), .ZN(
        n18739) );
  NAND3_X2 U18102 ( .A1(n27851), .A2(n7996), .A3(n27850), .ZN(n31422) );
  INV_X1 U18104 ( .A(n22087), .ZN(n20405) );
  INV_X1 U18106 ( .A(n30696), .ZN(n6253) );
  NAND4_X2 U18107 ( .A1(n12686), .A2(n12685), .A3(n12688), .A4(n12687), .ZN(
        n14911) );
  NAND4_X2 U18111 ( .A1(n12827), .A2(n12826), .A3(n12829), .A4(n12828), .ZN(
        n14803) );
  INV_X1 U18112 ( .A(n27234), .ZN(n7557) );
  XNOR2_X1 U18113 ( .A(n26303), .B(n7557), .ZN(n7182) );
  INV_X1 U18115 ( .A(n39195), .ZN(n37031) );
  INV_X1 U18116 ( .A(n10338), .ZN(n7530) );
  NOR2_X1 U18117 ( .A1(n8428), .A2(n8427), .ZN(n9250) );
  NAND4_X2 U18118 ( .A1(n10212), .A2(n10211), .A3(n10210), .A4(n10209), .ZN(
        n19248) );
  OAI211_X1 U18120 ( .C1(n39233), .C2(n39240), .A(n39242), .B(n2536), .ZN(
        n6848) );
  XNOR2_X1 U18124 ( .A(n8270), .B(n8269), .ZN(n8268) );
  AND2_X2 U18126 ( .A1(n20314), .A2(n21473), .ZN(n21460) );
  XNOR2_X1 U18127 ( .A(n28081), .B(n7899), .ZN(n7898) );
  XNOR2_X1 U18128 ( .A(n36974), .B(n2431), .ZN(n7385) );
  INV_X1 U18130 ( .A(n40477), .ZN(n37171) );
  OR2_X2 U18131 ( .A1(n46446), .A2(n46412), .ZN(n48463) );
  INV_X2 U18132 ( .A(n25789), .ZN(n28669) );
  NOR2_X1 U18133 ( .A1(n41430), .A2(n39767), .ZN(n7703) );
  NOR2_X1 U18134 ( .A1(n12223), .A2(n6073), .ZN(n13419) );
  OAI22_X1 U18135 ( .A1(n39751), .A2(n8199), .B1(n39938), .B2(n39937), .ZN(
        n8200) );
  INV_X2 U18136 ( .A(n36771), .ZN(n39262) );
  NAND4_X2 U18137 ( .A1(n14988), .A2(n14987), .A3(n14986), .A4(n14985), .ZN(
        n18831) );
  INV_X1 U18138 ( .A(n18897), .ZN(n7431) );
  NOR2_X1 U18139 ( .A1(n18245), .A2(n8630), .ZN(n8629) );
  XNOR2_X2 U18141 ( .A(n28245), .B(n28367), .ZN(n29764) );
  BUF_X2 U18142 ( .A(n8849), .Z(n10031) );
  INV_X1 U18143 ( .A(n9067), .ZN(n11797) );
  NAND2_X1 U18144 ( .A1(n767), .A2(n6180), .ZN(n6179) );
  NAND2_X1 U18145 ( .A1(n6182), .A2(n11282), .ZN(n6181) );
  OAI21_X1 U18146 ( .B1(n11668), .B2(n11676), .A(n6183), .ZN(n6182) );
  NAND2_X1 U18147 ( .A1(n11670), .A2(n11669), .ZN(n6183) );
  AND2_X2 U18148 ( .A1(n11685), .A2(n11270), .ZN(n11676) );
  NAND3_X1 U18149 ( .A1(n6186), .A2(n40204), .A3(n6185), .ZN(n38383) );
  NAND3_X1 U18152 ( .A1(n31169), .A2(n5867), .A3(n381), .ZN(n6189) );
  NAND2_X1 U18153 ( .A1(n6189), .A2(n6187), .ZN(n30802) );
  NAND2_X1 U18154 ( .A1(n31455), .A2(n31454), .ZN(n6187) );
  OAI21_X1 U18155 ( .B1(n30755), .B2(n51697), .A(n6191), .ZN(n6190) );
  INV_X1 U18156 ( .A(n16036), .ZN(n6193) );
  NAND2_X1 U18157 ( .A1(n6193), .A2(n6192), .ZN(n13040) );
  NOR2_X1 U18158 ( .A1(n13040), .A2(n13384), .ZN(n12810) );
  NAND2_X1 U18159 ( .A1(n6197), .A2(n33004), .ZN(n6196) );
  NAND3_X1 U18160 ( .A1(n31012), .A2(n31013), .A3(n6196), .ZN(n6195) );
  OAI21_X1 U18161 ( .B1(n40151), .B2(n6202), .A(n37470), .ZN(n6201) );
  NAND2_X1 U18162 ( .A1(n4950), .A2(n40556), .ZN(n6202) );
  INV_X1 U18163 ( .A(n23142), .ZN(n6207) );
  XNOR2_X1 U18164 ( .A(n24802), .B(n24801), .ZN(n6208) );
  XNOR2_X1 U18165 ( .A(n24815), .B(n25182), .ZN(n6209) );
  XNOR2_X1 U18166 ( .A(n45396), .B(n6210), .ZN(n45397) );
  XNOR2_X1 U18167 ( .A(n45395), .B(n45394), .ZN(n6210) );
  NAND2_X1 U18168 ( .A1(n11688), .A2(n10591), .ZN(n11681) );
  INV_X1 U18170 ( .A(n8997), .ZN(n6214) );
  NAND3_X1 U18171 ( .A1(n6219), .A2(n34992), .A3(n6216), .ZN(n6215) );
  NOR2_X1 U18172 ( .A1(n36542), .A2(n6218), .ZN(n6217) );
  INV_X1 U18173 ( .A(n37968), .ZN(n6219) );
  NAND3_X1 U18174 ( .A1(n29264), .A2(n28662), .A3(n28658), .ZN(n6220) );
  NAND2_X1 U18175 ( .A1(n35914), .A2(n36251), .ZN(n6221) );
  NAND2_X1 U18176 ( .A1(n19524), .A2(n21177), .ZN(n19528) );
  NAND2_X1 U18177 ( .A1(n19530), .A2(n19529), .ZN(n6225) );
  NAND2_X1 U18179 ( .A1(n6227), .A2(n598), .ZN(n21224) );
  INV_X1 U18180 ( .A(n17309), .ZN(n6227) );
  NAND2_X1 U18181 ( .A1(n19514), .A2(n19504), .ZN(n17309) );
  XNOR2_X2 U18182 ( .A(n6228), .B(n16654), .ZN(n19514) );
  XNOR2_X1 U18183 ( .A(n8408), .B(n17976), .ZN(n6228) );
  NAND2_X1 U18184 ( .A1(n47514), .A2(n46793), .ZN(n6231) );
  AOI22_X1 U18185 ( .A1(n46790), .A2(n47502), .B1(n46780), .B2(n47543), .ZN(
        n6232) );
  INV_X1 U18186 ( .A(n46795), .ZN(n6233) );
  NAND2_X1 U18187 ( .A1(n19438), .A2(n6237), .ZN(n19439) );
  NAND2_X1 U18188 ( .A1(n19437), .A2(n6238), .ZN(n6237) );
  INV_X1 U18189 ( .A(n22846), .ZN(n6238) );
  NAND2_X1 U18190 ( .A1(n4413), .A2(n22861), .ZN(n22846) );
  XNOR2_X1 U18191 ( .A(n24319), .B(n23941), .ZN(n28295) );
  AOI21_X1 U18193 ( .B1(n28158), .B2(n28872), .A(n6245), .ZN(n6244) );
  AND2_X1 U18194 ( .A1(n29033), .A2(n28874), .ZN(n6245) );
  NAND2_X1 U18195 ( .A1(n50034), .A2(n49731), .ZN(n47309) );
  NAND3_X1 U18196 ( .A1(n23154), .A2(n23157), .A3(n6247), .ZN(n19591) );
  NAND2_X1 U18197 ( .A1(n6010), .A2(n23473), .ZN(n6247) );
  INV_X1 U18198 ( .A(n32447), .ZN(n32445) );
  NAND2_X1 U18199 ( .A1(n31954), .A2(n32356), .ZN(n32447) );
  XNOR2_X1 U18201 ( .A(n46118), .B(n45049), .ZN(n45062) );
  NAND4_X4 U18202 ( .A1(n7240), .A2(n7237), .A3(n7238), .A4(n36096), .ZN(
        n44240) );
  NAND2_X1 U18203 ( .A1(n6254), .A2(n6252), .ZN(n28760) );
  NAND2_X1 U18204 ( .A1(n6253), .A2(n30392), .ZN(n6252) );
  NAND2_X1 U18205 ( .A1(n28757), .A2(n51257), .ZN(n6254) );
  NAND2_X1 U18206 ( .A1(n6255), .A2(n2479), .ZN(n30697) );
  NAND2_X1 U18207 ( .A1(n28757), .A2(n6256), .ZN(n6255) );
  NAND2_X1 U18208 ( .A1(n6257), .A2(n2438), .ZN(n30700) );
  NAND2_X1 U18209 ( .A1(n28757), .A2(n30393), .ZN(n6257) );
  NAND3_X1 U18210 ( .A1(n2523), .A2(n21712), .A3(n6260), .ZN(n6258) );
  NOR2_X1 U18212 ( .A1(n2141), .A2(n37649), .ZN(n36406) );
  NOR2_X1 U18213 ( .A1(n34630), .A2(n6262), .ZN(n34637) );
  NAND2_X1 U18214 ( .A1(n6264), .A2(n2141), .ZN(n6263) );
  XNOR2_X1 U18215 ( .A(n6265), .B(n4940), .ZN(n23122) );
  XNOR2_X1 U18216 ( .A(n6265), .B(n23682), .ZN(n23683) );
  XNOR2_X1 U18217 ( .A(n6265), .B(n24223), .ZN(n24224) );
  XNOR2_X1 U18218 ( .A(n7971), .B(n6265), .ZN(n25466) );
  NAND2_X2 U18219 ( .A1(n6266), .A2(n22872), .ZN(n6265) );
  NAND2_X1 U18220 ( .A1(n30821), .A2(n32906), .ZN(n6268) );
  NAND2_X1 U18221 ( .A1(n32896), .A2(n32906), .ZN(n6271) );
  NAND2_X1 U18222 ( .A1(n32540), .A2(n32634), .ZN(n32906) );
  XNOR2_X1 U18224 ( .A(n39125), .B(n51362), .ZN(n39154) );
  NAND2_X1 U18227 ( .A1(n14672), .A2(n14666), .ZN(n6274) );
  NAND3_X1 U18228 ( .A1(n7755), .A2(n51347), .A3(n785), .ZN(n6275) );
  NAND4_X2 U18229 ( .A1(n9398), .A2(n9399), .A3(n9397), .A4(n9396), .ZN(n14666) );
  INV_X1 U18230 ( .A(n36604), .ZN(n6276) );
  NAND2_X1 U18231 ( .A1(n6277), .A2(n22386), .ZN(n22388) );
  XNOR2_X1 U18232 ( .A(n15504), .B(n17976), .ZN(n15505) );
  XNOR2_X2 U18233 ( .A(n19261), .B(n16754), .ZN(n18750) );
  NAND2_X2 U18234 ( .A1(n15084), .A2(n15083), .ZN(n19261) );
  NAND2_X1 U18236 ( .A1(n15550), .A2(n15549), .ZN(n6280) );
  NAND2_X1 U18238 ( .A1(n8338), .A2(n27679), .ZN(n6284) );
  NAND4_X2 U18239 ( .A1(n6286), .A2(n34094), .A3(n8010), .A4(n8008), .ZN(
        n39857) );
  NAND2_X1 U18240 ( .A1(n32107), .A2(n32560), .ZN(n32087) );
  NAND2_X1 U18242 ( .A1(n29318), .A2(n29317), .ZN(n6288) );
  NAND2_X1 U18243 ( .A1(n29332), .A2(n29333), .ZN(n6289) );
  NAND2_X1 U18244 ( .A1(n46511), .A2(n48166), .ZN(n48421) );
  NAND2_X1 U18245 ( .A1(n15766), .A2(n2189), .ZN(n15061) );
  NAND2_X1 U18246 ( .A1(n52177), .A2(n29326), .ZN(n29328) );
  NAND4_X1 U18247 ( .A1(n6296), .A2(n6297), .A3(n6298), .A4(n7128), .ZN(n10210) );
  NAND2_X1 U18248 ( .A1(n14179), .A2(n12907), .ZN(n7128) );
  NAND2_X1 U18249 ( .A1(n13135), .A2(n13148), .ZN(n13150) );
  NAND2_X1 U18250 ( .A1(n6295), .A2(n13148), .ZN(n6297) );
  INV_X1 U18251 ( .A(n12213), .ZN(n6299) );
  NAND3_X1 U18252 ( .A1(n27831), .A2(n27832), .A3(n6602), .ZN(n6301) );
  NAND2_X1 U18253 ( .A1(n27869), .A2(n6307), .ZN(n6305) );
  NAND2_X1 U18255 ( .A1(n6305), .A2(n27873), .ZN(n6304) );
  OR2_X1 U18256 ( .A1(n27870), .A2(n29990), .ZN(n6307) );
  XNOR2_X1 U18257 ( .A(n28340), .B(n26425), .ZN(n6308) );
  NAND2_X1 U18258 ( .A1(n22413), .A2(n22414), .ZN(n24810) );
  NAND3_X1 U18259 ( .A1(n6312), .A2(n7131), .A3(n17059), .ZN(n16767) );
  NAND3_X1 U18261 ( .A1(n17603), .A2(n6312), .A3(n16788), .ZN(n17498) );
  NAND2_X1 U18262 ( .A1(n18314), .A2(n18313), .ZN(n6314) );
  NAND2_X1 U18263 ( .A1(n18323), .A2(n20093), .ZN(n6315) );
  INV_X1 U18264 ( .A(n38464), .ZN(n6317) );
  INV_X1 U18265 ( .A(n35103), .ZN(n37414) );
  NAND2_X1 U18266 ( .A1(n10532), .A2(n6319), .ZN(n8856) );
  NAND2_X1 U18267 ( .A1(n14572), .A2(n6320), .ZN(n10878) );
  NAND3_X1 U18268 ( .A1(n6323), .A2(n30851), .A3(n30850), .ZN(n6322) );
  NAND3_X1 U18269 ( .A1(n6324), .A2(n31034), .A3(n30849), .ZN(n6323) );
  NAND2_X1 U18270 ( .A1(n9221), .A2(n12055), .ZN(n6329) );
  NAND2_X1 U18271 ( .A1(n6329), .A2(n12062), .ZN(n6328) );
  NAND2_X1 U18273 ( .A1(n8378), .A2(n6333), .ZN(n17474) );
  NAND2_X1 U18274 ( .A1(n6331), .A2(n6330), .ZN(n18036) );
  NAND2_X1 U18275 ( .A1(n6333), .A2(n18041), .ZN(n6330) );
  NAND2_X1 U18277 ( .A1(n2222), .A2(n6333), .ZN(n18046) );
  INV_X1 U18278 ( .A(n15398), .ZN(n6333) );
  NAND2_X2 U18279 ( .A1(n6334), .A2(n39254), .ZN(n41685) );
  INV_X1 U18280 ( .A(n41238), .ZN(n41671) );
  NAND2_X1 U18281 ( .A1(n40211), .A2(n40210), .ZN(n40217) );
  NAND3_X1 U18282 ( .A1(n1555), .A2(n15421), .A3(n15425), .ZN(n13259) );
  OR2_X1 U18285 ( .A1(n27697), .A2(n6338), .ZN(n6340) );
  NAND2_X1 U18286 ( .A1(n5267), .A2(n6339), .ZN(n6338) );
  NAND2_X1 U18287 ( .A1(n23623), .A2(n6341), .ZN(n23630) );
  NAND2_X1 U18288 ( .A1(n23622), .A2(n754), .ZN(n6341) );
  NAND3_X1 U18289 ( .A1(n30168), .A2(n30167), .A3(n28021), .ZN(n30174) );
  NAND2_X1 U18290 ( .A1(n30174), .A2(n6342), .ZN(n28030) );
  NAND3_X1 U18291 ( .A1(n39233), .A2(n39232), .A3(n39234), .ZN(n39238) );
  NAND2_X1 U18292 ( .A1(n38706), .A2(n38704), .ZN(n39234) );
  XNOR2_X1 U18293 ( .A(n6345), .B(n43168), .ZN(n42529) );
  NAND2_X1 U18294 ( .A1(n6350), .A2(n6348), .ZN(n6347) );
  NAND2_X1 U18295 ( .A1(n6349), .A2(n14595), .ZN(n6348) );
  NAND2_X1 U18296 ( .A1(n8038), .A2(n12995), .ZN(n6349) );
  INV_X1 U18297 ( .A(n48068), .ZN(n6355) );
  NAND2_X1 U18298 ( .A1(n48059), .A2(n6353), .ZN(n48004) );
  INV_X1 U18299 ( .A(n48074), .ZN(n6353) );
  NAND2_X1 U18300 ( .A1(n6355), .A2(n48074), .ZN(n6354) );
  OAI211_X1 U18301 ( .C1(n20506), .C2(n8001), .A(n17587), .B(n20519), .ZN(
        n6356) );
  INV_X1 U18302 ( .A(n21925), .ZN(n21026) );
  NAND2_X1 U18303 ( .A1(n17606), .A2(n17605), .ZN(n6359) );
  OAI21_X1 U18304 ( .B1(n17601), .B2(n17602), .A(n20105), .ZN(n6360) );
  NAND2_X1 U18306 ( .A1(n6363), .A2(n590), .ZN(n18285) );
  OAI21_X1 U18307 ( .B1(n17523), .B2(n18287), .A(n6364), .ZN(n17528) );
  NAND2_X1 U18308 ( .A1(n18287), .A2(n20012), .ZN(n6364) );
  AND2_X1 U18309 ( .A1(n35167), .A2(n35164), .ZN(n6365) );
  NAND3_X2 U18310 ( .A1(n6365), .A2(n35165), .A3(n35166), .ZN(n41275) );
  NAND4_X2 U18311 ( .A1(n26491), .A2(n26492), .A3(n26490), .A4(n27959), .ZN(
        n31383) );
  NAND2_X1 U18312 ( .A1(n13621), .A2(n6366), .ZN(n12835) );
  INV_X1 U18313 ( .A(n14664), .ZN(n6366) );
  NAND2_X1 U18314 ( .A1(n21018), .A2(n21934), .ZN(n21020) );
  INV_X1 U18315 ( .A(n38132), .ZN(n6367) );
  XNOR2_X1 U18317 ( .A(n26055), .B(n26054), .ZN(n6368) );
  OR2_X2 U18319 ( .A1(n6371), .A2(n38826), .ZN(n45426) );
  NAND2_X1 U18320 ( .A1(n353), .A2(n22375), .ZN(n22729) );
  NAND2_X1 U18321 ( .A1(n15389), .A2(n14806), .ZN(n14488) );
  AND2_X1 U18322 ( .A1(n15380), .A2(n15384), .ZN(n15364) );
  INV_X1 U18323 ( .A(n15367), .ZN(n6378) );
  NAND2_X1 U18324 ( .A1(n787), .A2(n15380), .ZN(n15375) );
  AND3_X1 U18325 ( .A1(n11458), .A2(n11456), .A3(n11457), .ZN(n6379) );
  NOR2_X1 U18326 ( .A1(n8153), .A2(n23922), .ZN(n6381) );
  NAND2_X1 U18327 ( .A1(n14123), .A2(n6384), .ZN(n13458) );
  OR2_X1 U18328 ( .A1(n15161), .A2(n6384), .ZN(n13462) );
  NAND2_X1 U18329 ( .A1(n14574), .A2(n7715), .ZN(n10870) );
  XNOR2_X1 U18330 ( .A(n15163), .B(n6384), .ZN(n14581) );
  NAND3_X1 U18331 ( .A1(n10873), .A2(n15173), .A3(n7715), .ZN(n10874) );
  AOI21_X1 U18333 ( .B1(n48987), .B2(n6391), .A(n6386), .ZN(n46941) );
  NAND2_X1 U18334 ( .A1(n8472), .A2(n6387), .ZN(n48990) );
  NAND2_X1 U18335 ( .A1(n23), .A2(n49047), .ZN(n6387) );
  NOR2_X1 U18336 ( .A1(n6389), .A2(n52179), .ZN(n48988) );
  NAND2_X1 U18337 ( .A1(n51310), .A2(n6391), .ZN(n46936) );
  AND2_X1 U18338 ( .A1(n49030), .A2(n6391), .ZN(n49039) );
  NAND2_X1 U18339 ( .A1(n49034), .A2(n6391), .ZN(n49032) );
  NAND2_X1 U18340 ( .A1(n52179), .A2(n49019), .ZN(n6390) );
  INV_X1 U18341 ( .A(n40493), .ZN(n40501) );
  INV_X1 U18343 ( .A(n51106), .ZN(n7627) );
  NOR2_X1 U18344 ( .A1(n32608), .A2(n32620), .ZN(n31556) );
  NAND2_X1 U18345 ( .A1(n581), .A2(n21389), .ZN(n6395) );
  AND2_X1 U18346 ( .A1(n4246), .A2(n63), .ZN(n36491) );
  AOI22_X1 U18347 ( .A1(n7838), .A2(n31025), .B1(n31026), .B2(n51479), .ZN(
        n6400) );
  NAND3_X1 U18348 ( .A1(n31803), .A2(n31028), .A3(n31798), .ZN(n6402) );
  NOR2_X1 U18350 ( .A1(n30431), .A2(n6403), .ZN(n29859) );
  NOR2_X1 U18351 ( .A1(n487), .A2(n30425), .ZN(n6404) );
  NAND2_X1 U18352 ( .A1(n2394), .A2(n12541), .ZN(n6407) );
  INV_X1 U18353 ( .A(n9117), .ZN(n12541) );
  NAND2_X1 U18354 ( .A1(n12535), .A2(n442), .ZN(n6410) );
  XNOR2_X1 U18355 ( .A(n15185), .B(n6411), .ZN(n16897) );
  XNOR2_X1 U18356 ( .A(n17938), .B(n6412), .ZN(n6411) );
  NAND3_X1 U18357 ( .A1(n6414), .A2(n50015), .A3(n50016), .ZN(n6413) );
  NAND3_X1 U18358 ( .A1(n50011), .A2(n6416), .A3(n6415), .ZN(n6414) );
  NAND2_X1 U18359 ( .A1(n50329), .A2(n50009), .ZN(n6415) );
  NAND2_X1 U18360 ( .A1(n38950), .A2(n38953), .ZN(n39417) );
  NAND2_X1 U18361 ( .A1(n31379), .A2(n33002), .ZN(n6417) );
  OAI211_X1 U18362 ( .C1(n9175), .C2(n10449), .A(n10349), .B(n6423), .ZN(
        n10350) );
  INV_X1 U18363 ( .A(n25603), .ZN(n29252) );
  XNOR2_X1 U18365 ( .A(n43924), .B(n6425), .ZN(n43926) );
  NOR2_X1 U18366 ( .A1(n41588), .A2(n6426), .ZN(n6429) );
  NAND3_X1 U18367 ( .A1(n683), .A2(n42006), .A3(n6236), .ZN(n6426) );
  NAND3_X1 U18368 ( .A1(n41585), .A2(n6428), .A3(n41584), .ZN(n6427) );
  NAND2_X1 U18369 ( .A1(n6429), .A2(n42011), .ZN(n6428) );
  NOR2_X1 U18370 ( .A1(n41588), .A2(n41587), .ZN(n41580) );
  NAND3_X1 U18371 ( .A1(n19278), .A2(n19279), .A3(n19967), .ZN(n6431) );
  INV_X1 U18372 ( .A(n21155), .ZN(n6433) );
  NAND4_X2 U18373 ( .A1(n2271), .A2(n8320), .A3(n17072), .A4(n17073), .ZN(
        n21155) );
  NAND2_X1 U18374 ( .A1(n4987), .A2(n22849), .ZN(n19610) );
  INV_X1 U18375 ( .A(n33174), .ZN(n38027) );
  NAND2_X1 U18376 ( .A1(n35159), .A2(n35155), .ZN(n36373) );
  XNOR2_X1 U18377 ( .A(n25385), .B(n6434), .ZN(n16856) );
  XNOR2_X1 U18378 ( .A(n24461), .B(n6434), .ZN(n24462) );
  XNOR2_X1 U18379 ( .A(n6434), .B(n25224), .ZN(n25225) );
  NAND4_X2 U18380 ( .A1(n16135), .A2(n16133), .A3(n16132), .A4(n16134), .ZN(
        n6434) );
  XNOR2_X1 U18381 ( .A(n17802), .B(n19244), .ZN(n17807) );
  XNOR2_X2 U18382 ( .A(n8670), .B(n9170), .ZN(n19244) );
  NAND3_X2 U18383 ( .A1(n36388), .A2(n6440), .A3(n6436), .ZN(n40651) );
  NAND2_X1 U18384 ( .A1(n6439), .A2(n6438), .ZN(n6437) );
  AOI21_X1 U18385 ( .B1(n36380), .B2(n38034), .A(n36381), .ZN(n6438) );
  NAND2_X1 U18386 ( .A1(n36379), .A2(n38043), .ZN(n6439) );
  INV_X1 U18387 ( .A(n40651), .ZN(n39157) );
  NAND2_X1 U18388 ( .A1(n36377), .A2(n36376), .ZN(n6441) );
  NAND2_X1 U18389 ( .A1(n36369), .A2(n36370), .ZN(n6442) );
  NAND2_X1 U18390 ( .A1(n14307), .A2(n13826), .ZN(n11796) );
  NAND2_X1 U18391 ( .A1(n9024), .A2(n9787), .ZN(n6446) );
  XNOR2_X1 U18392 ( .A(n24450), .B(n24449), .ZN(n6448) );
  NAND2_X1 U18393 ( .A1(n36578), .A2(n36577), .ZN(n6451) );
  NAND2_X1 U18394 ( .A1(n6452), .A2(n17838), .ZN(n20434) );
  NAND3_X1 U18395 ( .A1(n6452), .A2(n17838), .A3(n6454), .ZN(n6453) );
  NAND2_X1 U18396 ( .A1(n6455), .A2(n6453), .ZN(n19325) );
  INV_X1 U18397 ( .A(n20432), .ZN(n6454) );
  NAND2_X1 U18398 ( .A1(n19323), .A2(n20432), .ZN(n6455) );
  INV_X1 U18400 ( .A(n37224), .ZN(n6456) );
  INV_X1 U18401 ( .A(n37228), .ZN(n6457) );
  NAND2_X1 U18402 ( .A1(n31093), .A2(n29387), .ZN(n6458) );
  NAND2_X1 U18403 ( .A1(n29392), .A2(n31094), .ZN(n6459) );
  NAND2_X1 U18404 ( .A1(n29386), .A2(n31087), .ZN(n6460) );
  INV_X1 U18405 ( .A(n6462), .ZN(n21314) );
  NOR2_X1 U18406 ( .A1(n23185), .A2(n6462), .ZN(n22670) );
  INV_X1 U18407 ( .A(n26944), .ZN(n27662) );
  NOR2_X1 U18408 ( .A1(n5307), .A2(n12052), .ZN(n6464) );
  OAI211_X1 U18409 ( .C1(n21618), .C2(n21637), .A(n21626), .B(n6467), .ZN(
        n6466) );
  INV_X1 U18410 ( .A(n21626), .ZN(n20255) );
  NAND2_X1 U18411 ( .A1(n6466), .A2(n21639), .ZN(n20263) );
  OR2_X1 U18412 ( .A1(n20254), .A2(n21630), .ZN(n6467) );
  INV_X1 U18415 ( .A(n41348), .ZN(n6471) );
  OAI21_X1 U18416 ( .B1(n6473), .B2(n8278), .A(n6472), .ZN(n6701) );
  NAND2_X1 U18417 ( .A1(n52107), .A2(n49450), .ZN(n6473) );
  NAND2_X1 U18419 ( .A1(n38747), .A2(n38746), .ZN(n6474) );
  INV_X1 U18420 ( .A(n21196), .ZN(n6476) );
  INV_X1 U18421 ( .A(n11419), .ZN(n6477) );
  NAND2_X1 U18422 ( .A1(n14096), .A2(n14453), .ZN(n6494) );
  INV_X1 U18423 ( .A(n6479), .ZN(n12372) );
  XNOR2_X1 U18424 ( .A(n42326), .B(n52084), .ZN(n42335) );
  NAND2_X1 U18425 ( .A1(n39529), .A2(n39530), .ZN(n6480) );
  NAND2_X1 U18426 ( .A1(n14453), .A2(n6481), .ZN(n12972) );
  NAND3_X1 U18427 ( .A1(n14442), .A2(n6481), .A3(n640), .ZN(n14443) );
  NOR2_X1 U18428 ( .A1(n14453), .A2(n6481), .ZN(n11432) );
  AOI21_X1 U18429 ( .B1(n14450), .B2(n6481), .A(n14455), .ZN(n14451) );
  INV_X1 U18430 ( .A(n47174), .ZN(n6482) );
  NAND3_X1 U18431 ( .A1(n50773), .A2(n50787), .A3(n50798), .ZN(n47174) );
  OAI211_X1 U18432 ( .C1(n51353), .C2(n50808), .A(n6482), .B(n50738), .ZN(
        n50758) );
  OR2_X1 U18433 ( .A1(n52147), .A2(n6483), .ZN(n29240) );
  NAND2_X1 U18434 ( .A1(n27918), .A2(n30256), .ZN(n6483) );
  NAND2_X1 U18435 ( .A1(n29235), .A2(n6488), .ZN(n27971) );
  OAI21_X1 U18436 ( .B1(n52147), .B2(n2158), .A(n6484), .ZN(n30262) );
  NAND2_X1 U18437 ( .A1(n2158), .A2(n6485), .ZN(n6484) );
  OR2_X1 U18438 ( .A1(n52147), .A2(n6486), .ZN(n6485) );
  OAI21_X1 U18439 ( .B1(n29235), .B2(n6488), .A(n30263), .ZN(n6487) );
  XNOR2_X2 U18440 ( .A(n8984), .B(Key[158]), .ZN(n10742) );
  OAI21_X1 U18441 ( .B1(n585), .B2(n19865), .A(n6489), .ZN(n19031) );
  NAND2_X1 U18442 ( .A1(n19871), .A2(n19853), .ZN(n6489) );
  INV_X1 U18443 ( .A(n16986), .ZN(n19649) );
  OAI22_X1 U18444 ( .A1(n32202), .A2(n32210), .B1(n6969), .B2(n32194), .ZN(
        n29105) );
  NAND2_X1 U18445 ( .A1(n6969), .A2(n32194), .ZN(n32202) );
  AOI22_X1 U18446 ( .A1(n6493), .A2(n14097), .B1(n51384), .B2(n6491), .ZN(
        n6495) );
  NAND2_X1 U18447 ( .A1(n14097), .A2(n6492), .ZN(n14436) );
  NOR2_X1 U18448 ( .A1(n6494), .A2(n14444), .ZN(n6493) );
  NAND2_X1 U18449 ( .A1(n19011), .A2(n19005), .ZN(n6497) );
  NAND2_X1 U18450 ( .A1(n19012), .A2(n6499), .ZN(n6498) );
  NAND2_X1 U18451 ( .A1(n41533), .A2(n6505), .ZN(n6504) );
  OAI21_X1 U18452 ( .B1(n39696), .B2(n51455), .A(n6507), .ZN(n6509) );
  NAND2_X1 U18453 ( .A1(n6509), .A2(n39697), .ZN(n6508) );
  XNOR2_X2 U18454 ( .A(n28396), .B(n25909), .ZN(n26053) );
  NAND2_X1 U18455 ( .A1(n6515), .A2(n20044), .ZN(n17044) );
  NAND2_X1 U18456 ( .A1(n6516), .A2(n8704), .ZN(n15403) );
  NAND2_X1 U18457 ( .A1(n32602), .A2(n32988), .ZN(n6517) );
  INV_X1 U18458 ( .A(n32589), .ZN(n6522) );
  NAND2_X1 U18459 ( .A1(n32604), .A2(n6520), .ZN(n6519) );
  NAND2_X1 U18463 ( .A1(n40873), .A2(n40876), .ZN(n39966) );
  INV_X1 U18465 ( .A(n45747), .ZN(n6526) );
  NAND2_X1 U18466 ( .A1(n45211), .A2(n49170), .ZN(n6527) );
  NAND2_X1 U18467 ( .A1(n45210), .A2(n49161), .ZN(n6528) );
  NAND2_X1 U18468 ( .A1(n19426), .A2(n6529), .ZN(n19428) );
  NAND3_X1 U18469 ( .A1(n6530), .A2(n19435), .A3(n21885), .ZN(n22334) );
  NAND2_X1 U18470 ( .A1(n8111), .A2(n45575), .ZN(n6531) );
  OAI21_X1 U18471 ( .B1(n48176), .B2(n48175), .A(n6531), .ZN(n48185) );
  NAND2_X1 U18472 ( .A1(n7289), .A2(n6531), .ZN(n45586) );
  NAND3_X1 U18473 ( .A1(n6532), .A2(n45213), .A3(n48808), .ZN(n48806) );
  NAND3_X1 U18474 ( .A1(n37833), .A2(n39830), .A3(n40384), .ZN(n6534) );
  NAND2_X1 U18475 ( .A1(n1931), .A2(n40381), .ZN(n40384) );
  NAND2_X1 U18476 ( .A1(n40380), .A2(n38622), .ZN(n37833) );
  NAND2_X1 U18477 ( .A1(n37837), .A2(n40385), .ZN(n6535) );
  NAND3_X1 U18478 ( .A1(n39487), .A2(n37798), .A3(n39472), .ZN(n37799) );
  NAND2_X1 U18479 ( .A1(n46255), .A2(n664), .ZN(n6536) );
  AOI22_X1 U18480 ( .A1(n9675), .A2(n12097), .B1(n9676), .B2(n11351), .ZN(
        n6537) );
  NAND4_X1 U18481 ( .A1(n9681), .A2(n9683), .A3(n9682), .A4(n6537), .ZN(n11732) );
  NAND2_X1 U18482 ( .A1(n30073), .A2(n29591), .ZN(n31122) );
  AND4_X2 U18483 ( .A1(n26897), .A2(n26896), .A3(n26895), .A4(n26894), .ZN(
        n30073) );
  INV_X1 U18484 ( .A(n38543), .ZN(n6538) );
  NAND2_X1 U18485 ( .A1(n6541), .A2(n34971), .ZN(n34976) );
  NOR2_X1 U18486 ( .A1(n6541), .A2(n38019), .ZN(n32679) );
  NAND2_X1 U18487 ( .A1(n38177), .A2(n6541), .ZN(n38180) );
  OAI22_X1 U18488 ( .A1(n38013), .A2(n38012), .B1(n38014), .B2(n6541), .ZN(
        n38022) );
  OAI211_X1 U18489 ( .C1(n35027), .C2(n6541), .A(n38015), .B(n38189), .ZN(
        n34977) );
  OAI22_X1 U18490 ( .A1(n35025), .A2(n6541), .B1(n38190), .B2(n38015), .ZN(
        n7070) );
  NAND2_X1 U18491 ( .A1(n35024), .A2(n6541), .ZN(n35030) );
  NAND4_X2 U18492 ( .A1(n11990), .A2(n11991), .A3(n11989), .A4(n11988), .ZN(
        n15324) );
  NAND3_X1 U18493 ( .A1(n41940), .A2(n41942), .A3(n41941), .ZN(n6545) );
  INV_X1 U18494 ( .A(n11979), .ZN(n12663) );
  INV_X1 U18495 ( .A(n12660), .ZN(n12648) );
  OAI211_X1 U18496 ( .C1(n11979), .C2(n12661), .A(n11977), .B(n11971), .ZN(
        n11972) );
  NAND2_X1 U18497 ( .A1(n10338), .A2(n11986), .ZN(n11971) );
  INV_X1 U18499 ( .A(n41147), .ZN(n38617) );
  NAND2_X1 U18500 ( .A1(n52083), .A2(n40388), .ZN(n41147) );
  INV_X1 U18501 ( .A(n39453), .ZN(n6553) );
  INV_X1 U18502 ( .A(n39450), .ZN(n34800) );
  NOR2_X1 U18503 ( .A1(n45179), .A2(n51292), .ZN(n47078) );
  INV_X1 U18504 ( .A(n46816), .ZN(n47074) );
  INV_X1 U18505 ( .A(n6558), .ZN(n6556) );
  NAND2_X1 U18506 ( .A1(n26638), .A2(n26635), .ZN(n6558) );
  OAI21_X1 U18507 ( .B1(n30533), .B2(n3241), .A(n30529), .ZN(n6562) );
  NAND3_X1 U18508 ( .A1(n6760), .A2(n6556), .A3(n6560), .ZN(n6555) );
  NAND2_X1 U18509 ( .A1(n6560), .A2(n6557), .ZN(n7550) );
  XNOR2_X2 U18510 ( .A(n8557), .B(n17176), .ZN(n21185) );
  XNOR2_X2 U18511 ( .A(n14378), .B(n6563), .ZN(n17546) );
  OAI21_X1 U18513 ( .B1(n6570), .B2(n6567), .A(n6569), .ZN(n6566) );
  NAND2_X1 U18514 ( .A1(n6570), .A2(n6569), .ZN(n6568) );
  NAND3_X1 U18515 ( .A1(n6571), .A2(n12619), .A3(n10462), .ZN(n10323) );
  NAND2_X1 U18516 ( .A1(n6572), .A2(n12620), .ZN(n9211) );
  XNOR2_X1 U18517 ( .A(n6573), .B(n47401), .ZN(n43216) );
  XNOR2_X1 U18518 ( .A(n6573), .B(n42560), .ZN(n42561) );
  XNOR2_X1 U18520 ( .A(n6573), .B(n42350), .ZN(n42351) );
  NAND4_X2 U18521 ( .A1(n41625), .A2(n41627), .A3(n41628), .A4(n41626), .ZN(
        n6573) );
  INV_X2 U18522 ( .A(n50744), .ZN(n50798) );
  NAND2_X1 U18523 ( .A1(n39484), .A2(n36216), .ZN(n38981) );
  NOR2_X1 U18526 ( .A1(n32486), .A2(n32025), .ZN(n29625) );
  NAND2_X1 U18527 ( .A1(n32791), .A2(n32784), .ZN(n6577) );
  INV_X1 U18528 ( .A(n680), .ZN(n6578) );
  OAI211_X1 U18529 ( .C1(n6579), .C2(n42205), .A(n41925), .B(n41926), .ZN(
        n41929) );
  NAND2_X1 U18530 ( .A1(n6617), .A2(n41938), .ZN(n6579) );
  OR2_X1 U18531 ( .A1(n40248), .A2(n6580), .ZN(n38923) );
  NAND3_X1 U18533 ( .A1(n27685), .A2(n27582), .A3(n26955), .ZN(n24468) );
  XNOR2_X1 U18534 ( .A(n33941), .B(n33927), .ZN(n6582) );
  XNOR2_X1 U18535 ( .A(n6583), .B(n2200), .ZN(n15689) );
  XNOR2_X1 U18536 ( .A(n17666), .B(n52205), .ZN(n17670) );
  XNOR2_X1 U18537 ( .A(n6583), .B(n17794), .ZN(n17795) );
  XNOR2_X1 U18538 ( .A(n13865), .B(n52205), .ZN(n13866) );
  XNOR2_X1 U18539 ( .A(n52205), .B(n15800), .ZN(n16234) );
  NAND2_X1 U18540 ( .A1(n6584), .A2(n10513), .ZN(n10515) );
  OAI22_X1 U18541 ( .A1(n9836), .A2(n8438), .B1(n10526), .B2(n6584), .ZN(n6608) );
  INV_X1 U18542 ( .A(n6585), .ZN(n6589) );
  NOR2_X1 U18544 ( .A1(n22721), .A2(n22470), .ZN(n6591) );
  OAI21_X1 U18545 ( .B1(n22716), .B2(n22488), .A(n22709), .ZN(n6592) );
  NAND2_X1 U18546 ( .A1(n2083), .A2(n22464), .ZN(n22709) );
  NOR2_X1 U18548 ( .A1(n30290), .A2(n27113), .ZN(n27115) );
  NAND2_X1 U18549 ( .A1(n34653), .A2(n36425), .ZN(n36060) );
  AND4_X2 U18550 ( .A1(n2246), .A2(n18911), .A3(n18912), .A4(n2525), .ZN(
        n21873) );
  NAND2_X1 U18551 ( .A1(n609), .A2(n38763), .ZN(n43334) );
  INV_X1 U18552 ( .A(n38763), .ZN(n39613) );
  INV_X1 U18553 ( .A(n43334), .ZN(n41006) );
  AND2_X1 U18555 ( .A1(n41083), .A2(n41085), .ZN(n38868) );
  NAND2_X1 U18556 ( .A1(n19869), .A2(n374), .ZN(n19867) );
  XNOR2_X1 U18557 ( .A(n17225), .B(n16958), .ZN(n6599) );
  INV_X1 U18558 ( .A(n33562), .ZN(n35573) );
  INV_X1 U18559 ( .A(n38491), .ZN(n37524) );
  XNOR2_X1 U18560 ( .A(n42278), .B(n6600), .ZN(n40467) );
  INV_X1 U18561 ( .A(n45285), .ZN(n6600) );
  NAND2_X1 U18562 ( .A1(n22908), .A2(n22367), .ZN(n22914) );
  NAND2_X1 U18564 ( .A1(n17618), .A2(n20503), .ZN(n22357) );
  XNOR2_X1 U18565 ( .A(n6603), .B(n32802), .ZN(n32803) );
  XNOR2_X1 U18566 ( .A(n6603), .B(n35790), .ZN(n36680) );
  XNOR2_X1 U18567 ( .A(n6603), .B(n34739), .ZN(n35360) );
  XNOR2_X1 U18568 ( .A(n33082), .B(n51361), .ZN(n34230) );
  NOR2_X1 U18569 ( .A1(n47613), .A2(n47586), .ZN(n6604) );
  NAND3_X1 U18570 ( .A1(n29354), .A2(n7817), .A3(n29353), .ZN(n6607) );
  MUX2_X1 U18571 ( .A(n17412), .B(n19520), .S(n598), .Z(n16684) );
  OAI22_X1 U18572 ( .A1(n16674), .A2(n765), .B1(n7050), .B2(n21234), .ZN(
        n16675) );
  NAND2_X1 U18573 ( .A1(n6608), .A2(n10520), .ZN(n9489) );
  INV_X1 U18574 ( .A(n13136), .ZN(n6609) );
  NOR2_X1 U18575 ( .A1(n14184), .A2(n14183), .ZN(n6610) );
  NAND2_X1 U18576 ( .A1(n13135), .A2(n13152), .ZN(n13138) );
  NAND2_X1 U18577 ( .A1(n14182), .A2(n14181), .ZN(n6611) );
  NAND3_X1 U18578 ( .A1(n13135), .A2(n13152), .A3(n6609), .ZN(n14181) );
  NAND2_X1 U18579 ( .A1(n6612), .A2(n38337), .ZN(n35410) );
  OAI21_X1 U18583 ( .B1(n31087), .B2(n31086), .A(n31088), .ZN(n8333) );
  NAND2_X1 U18584 ( .A1(n50675), .A2(n50721), .ZN(n6620) );
  NAND2_X1 U18585 ( .A1(n6618), .A2(n50677), .ZN(n50690) );
  NAND2_X1 U18586 ( .A1(n50729), .A2(n6620), .ZN(n7748) );
  NAND2_X1 U18587 ( .A1(n23151), .A2(n23152), .ZN(n6621) );
  NAND2_X1 U18588 ( .A1(n6624), .A2(n23467), .ZN(n6623) );
  AND3_X1 U18589 ( .A1(n23153), .A2(n6010), .A3(n23157), .ZN(n6624) );
  NAND3_X1 U18590 ( .A1(n23467), .A2(n23465), .A3(n23160), .ZN(n7043) );
  NAND2_X1 U18592 ( .A1(n6628), .A2(n21649), .ZN(n6626) );
  NAND2_X1 U18593 ( .A1(n19401), .A2(n764), .ZN(n6631) );
  INV_X1 U18594 ( .A(n37516), .ZN(n37527) );
  NAND3_X1 U18595 ( .A1(n6633), .A2(n37526), .A3(n6632), .ZN(n35948) );
  OR2_X1 U18596 ( .A1(n37516), .A2(n37386), .ZN(n6632) );
  AOI21_X1 U18597 ( .B1(n37517), .B2(n38501), .A(n38494), .ZN(n6633) );
  NAND2_X1 U18598 ( .A1(n13104), .A2(n11821), .ZN(n6634) );
  NAND2_X2 U18599 ( .A1(n8710), .A2(n29145), .ZN(n32407) );
  NAND3_X1 U18600 ( .A1(n7430), .A2(n6635), .A3(n32407), .ZN(n32414) );
  NAND2_X1 U18601 ( .A1(n25418), .A2(n6636), .ZN(n29227) );
  AND2_X1 U18602 ( .A1(n52102), .A2(n25107), .ZN(n6636) );
  NAND2_X1 U18603 ( .A1(n6638), .A2(n37637), .ZN(n36004) );
  NOR2_X1 U18604 ( .A1(n6639), .A2(n46533), .ZN(n46534) );
  NAND2_X1 U18605 ( .A1(n6642), .A2(n6641), .ZN(n6640) );
  NAND2_X1 U18606 ( .A1(n30125), .A2(n31873), .ZN(n28490) );
  INV_X1 U18607 ( .A(n39912), .ZN(n6645) );
  NAND2_X1 U18608 ( .A1(n6647), .A2(n36396), .ZN(n6646) );
  INV_X1 U18609 ( .A(n48481), .ZN(n48488) );
  XNOR2_X2 U18610 ( .A(n44379), .B(n44378), .ZN(n48248) );
  NAND2_X1 U18611 ( .A1(n19046), .A2(n19045), .ZN(n6651) );
  INV_X1 U18612 ( .A(n19053), .ZN(n6652) );
  INV_X1 U18613 ( .A(n43629), .ZN(n6653) );
  NAND2_X1 U18616 ( .A1(n41573), .A2(n4943), .ZN(n42003) );
  NAND2_X1 U18617 ( .A1(n41588), .A2(n41997), .ZN(n41573) );
  XNOR2_X1 U18619 ( .A(n26147), .B(n6656), .ZN(n25715) );
  XNOR2_X1 U18620 ( .A(n6656), .B(n51415), .ZN(n27221) );
  XNOR2_X2 U18621 ( .A(n26375), .B(n6656), .ZN(n26556) );
  XNOR2_X1 U18622 ( .A(n6656), .B(n26378), .ZN(n27362) );
  INV_X1 U18623 ( .A(n37489), .ZN(n37437) );
  OR2_X2 U18625 ( .A1(n38540), .A2(n38539), .ZN(n41328) );
  NAND2_X1 U18626 ( .A1(n6661), .A2(n11346), .ZN(n12250) );
  AOI21_X1 U18627 ( .B1(n7286), .B2(n6661), .A(n7285), .ZN(n9643) );
  OAI211_X1 U18628 ( .C1(n9423), .C2(n6661), .A(n9422), .B(n9421), .ZN(n9424)
         );
  OAI21_X1 U18629 ( .B1(n10745), .B2(n10744), .A(n6661), .ZN(n10751) );
  NAND2_X1 U18630 ( .A1(n23631), .A2(n6662), .ZN(n23649) );
  INV_X1 U18631 ( .A(n20847), .ZN(n6662) );
  XNOR2_X1 U18632 ( .A(n44209), .B(n6663), .ZN(n42739) );
  XNOR2_X1 U18633 ( .A(n42561), .B(n6663), .ZN(n42567) );
  XNOR2_X1 U18634 ( .A(n2103), .B(n6663), .ZN(n40722) );
  XNOR2_X1 U18635 ( .A(n45389), .B(n6663), .ZN(n42455) );
  XNOR2_X1 U18636 ( .A(n42670), .B(n6663), .ZN(n43661) );
  XNOR2_X1 U18637 ( .A(n45042), .B(n6663), .ZN(n45044) );
  XNOR2_X2 U18638 ( .A(n44017), .B(n44217), .ZN(n6663) );
  NAND2_X1 U18639 ( .A1(n6664), .A2(n52091), .ZN(n45741) );
  NAND2_X1 U18640 ( .A1(n51328), .A2(n45711), .ZN(n48821) );
  NAND2_X1 U18642 ( .A1(n24033), .A2(n22107), .ZN(n23393) );
  NAND4_X2 U18643 ( .A1(n6666), .A2(n14236), .A3(n14237), .A4(n14235), .ZN(
        n17973) );
  NAND2_X1 U18644 ( .A1(n14233), .A2(n14232), .ZN(n6667) );
  NAND2_X1 U18645 ( .A1(n13208), .A2(n13207), .ZN(n13209) );
  NAND2_X1 U18646 ( .A1(n47291), .A2(n6669), .ZN(n44613) );
  NAND2_X1 U18647 ( .A1(n6669), .A2(n50351), .ZN(n49962) );
  AOI22_X1 U18648 ( .A1(n49961), .A2(n50347), .B1(n44608), .B2(n6669), .ZN(
        n49970) );
  MUX2_X1 U18649 ( .A(n47286), .B(n47287), .S(n44607), .Z(n47297) );
  NAND2_X1 U18650 ( .A1(n51026), .A2(n50344), .ZN(n44607) );
  XNOR2_X2 U18651 ( .A(n6670), .B(n18471), .ZN(n18495) );
  NAND2_X1 U18653 ( .A1(n9914), .A2(n10068), .ZN(n6672) );
  NAND2_X1 U18654 ( .A1(n48269), .A2(n6673), .ZN(n44430) );
  NOR2_X1 U18655 ( .A1(n48433), .A2(n48273), .ZN(n6673) );
  OAI21_X1 U18656 ( .B1(n48429), .B2(n6674), .A(n48433), .ZN(n44669) );
  NAND2_X1 U18657 ( .A1(n9636), .A2(n11359), .ZN(n11373) );
  NOR2_X1 U18658 ( .A1(n12111), .A2(n6675), .ZN(n9633) );
  INV_X1 U18659 ( .A(n9636), .ZN(n6675) );
  INV_X1 U18660 ( .A(n47858), .ZN(n47803) );
  AOI21_X1 U18661 ( .B1(n47817), .B2(n47803), .A(n6679), .ZN(n47822) );
  NAND3_X1 U18662 ( .A1(n598), .A2(n19503), .A3(n52065), .ZN(n21231) );
  NAND2_X1 U18664 ( .A1(n26068), .A2(n27830), .ZN(n6681) );
  NAND3_X1 U18667 ( .A1(n35146), .A2(n38567), .A3(n688), .ZN(n6777) );
  NAND2_X1 U18668 ( .A1(n29698), .A2(n29703), .ZN(n30430) );
  NAND3_X1 U18669 ( .A1(n8024), .A2(n12514), .A3(n12518), .ZN(n8915) );
  NAND2_X1 U18670 ( .A1(n10826), .A2(n6683), .ZN(n9157) );
  NOR2_X1 U18671 ( .A1(n11255), .A2(n6684), .ZN(n6683) );
  NAND3_X1 U18672 ( .A1(n6685), .A2(n49228), .A3(n49376), .ZN(n49285) );
  OR2_X1 U18673 ( .A1(n6687), .A2(n15108), .ZN(n6686) );
  INV_X1 U18675 ( .A(n15108), .ZN(n14974) );
  OAI211_X1 U18676 ( .C1(n14242), .C2(n14245), .A(n8977), .B(n6686), .ZN(n8978) );
  NAND2_X1 U18677 ( .A1(n352), .A2(n14982), .ZN(n6687) );
  NAND2_X2 U18678 ( .A1(n49681), .A2(n6688), .ZN(n49850) );
  INV_X1 U18679 ( .A(n49820), .ZN(n6689) );
  NAND2_X1 U18680 ( .A1(n49766), .A2(n49782), .ZN(n49820) );
  NAND3_X1 U18681 ( .A1(n6692), .A2(n23480), .A3(n6691), .ZN(n6690) );
  NAND3_X1 U18682 ( .A1(n23478), .A2(n23489), .A3(n23479), .ZN(n6691) );
  NAND2_X1 U18683 ( .A1(n23486), .A2(n23477), .ZN(n6692) );
  NAND2_X1 U18684 ( .A1(n6694), .A2(n23485), .ZN(n6693) );
  OAI22_X1 U18685 ( .A1(n23484), .A2(n23483), .B1(n23482), .B2(n23481), .ZN(
        n6694) );
  OAI211_X1 U18686 ( .C1(n6698), .C2(n6697), .A(n6696), .B(n6695), .ZN(
        Plaintext[109]) );
  NAND2_X1 U18687 ( .A1(n6698), .A2(n47205), .ZN(n6695) );
  NAND4_X1 U18688 ( .A1(n47204), .A2(n6700), .A3(n47202), .A4(n6699), .ZN(
        n6698) );
  NAND2_X1 U18689 ( .A1(n49417), .A2(n6703), .ZN(n6699) );
  NAND3_X1 U18690 ( .A1(n49459), .A2(n49461), .A3(n6702), .ZN(n6700) );
  AND2_X1 U18691 ( .A1(n51091), .A2(n49445), .ZN(n6702) );
  AND2_X1 U18692 ( .A1(n47201), .A2(n49443), .ZN(n6703) );
  NAND2_X1 U18693 ( .A1(n49721), .A2(n51094), .ZN(n46001) );
  XNOR2_X1 U18694 ( .A(n32803), .B(n32758), .ZN(n6707) );
  OAI21_X1 U18695 ( .B1(n29151), .B2(n6709), .A(n29150), .ZN(n29165) );
  NAND2_X1 U18696 ( .A1(n14199), .A2(n51671), .ZN(n14082) );
  NAND3_X1 U18697 ( .A1(n12388), .A2(n12386), .A3(n12387), .ZN(n6710) );
  MUX2_X1 U18698 ( .A(n16815), .B(n16816), .S(n18374), .Z(n16817) );
  NAND2_X1 U18699 ( .A1(n10683), .A2(n6712), .ZN(n10685) );
  NAND2_X1 U18703 ( .A1(n40338), .A2(n39855), .ZN(n39647) );
  NAND2_X1 U18704 ( .A1(n6716), .A2(n28520), .ZN(n6715) );
  NAND2_X1 U18705 ( .A1(n11353), .A2(n6786), .ZN(n12371) );
  INV_X1 U18706 ( .A(n23755), .ZN(n24191) );
  XNOR2_X1 U18707 ( .A(n25915), .B(n6720), .ZN(n6719) );
  XNOR2_X2 U18708 ( .A(n26509), .B(n20174), .ZN(n25915) );
  NAND2_X1 U18709 ( .A1(n20890), .A2(n23411), .ZN(n22317) );
  NAND2_X1 U18710 ( .A1(n20091), .A2(n20090), .ZN(n6722) );
  NAND2_X1 U18712 ( .A1(n6725), .A2(n6724), .ZN(n13739) );
  NAND2_X1 U18713 ( .A1(n13738), .A2(n6726), .ZN(n6725) );
  NAND2_X1 U18714 ( .A1(n6728), .A2(n21629), .ZN(n6727) );
  NAND2_X1 U18715 ( .A1(n35000), .A2(n2532), .ZN(n35004) );
  NAND3_X1 U18716 ( .A1(n40751), .A2(n41348), .A3(n41360), .ZN(n40746) );
  NAND2_X1 U18717 ( .A1(n778), .A2(n18313), .ZN(n17056) );
  INV_X1 U18718 ( .A(n18313), .ZN(n20104) );
  NAND2_X1 U18719 ( .A1(n14712), .A2(n14720), .ZN(n13338) );
  NAND2_X1 U18720 ( .A1(n38528), .A2(n38529), .ZN(n38531) );
  XNOR2_X1 U18722 ( .A(n37137), .B(n52164), .ZN(n35464) );
  XNOR2_X1 U18723 ( .A(n7544), .B(n52164), .ZN(n34519) );
  NAND2_X1 U18724 ( .A1(n6730), .A2(n5417), .ZN(n27146) );
  NOR2_X1 U18725 ( .A1(n51726), .A2(n6730), .ZN(n6970) );
  NAND2_X1 U18726 ( .A1(n27951), .A2(n51726), .ZN(n27961) );
  AOI21_X1 U18727 ( .B1(n29146), .B2(n6730), .A(n30245), .ZN(n29151) );
  XNOR2_X1 U18728 ( .A(n23881), .B(n6731), .ZN(n6732) );
  XNOR2_X1 U18729 ( .A(n28067), .B(n2293), .ZN(n6731) );
  NOR2_X1 U18731 ( .A1(n38557), .A2(n6734), .ZN(n38218) );
  OAI21_X1 U18733 ( .B1(n38548), .B2(n38547), .A(n6735), .ZN(n7660) );
  NAND2_X1 U18734 ( .A1(n40002), .A2(n40011), .ZN(n40018) );
  NAND2_X1 U18735 ( .A1(n6743), .A2(n6742), .ZN(n45762) );
  NAND2_X1 U18736 ( .A1(n45760), .A2(n46637), .ZN(n6743) );
  NAND3_X1 U18739 ( .A1(n38721), .A2(n5593), .A3(n2436), .ZN(n6749) );
  OAI21_X1 U18741 ( .B1(n6757), .B2(n44417), .A(n6750), .ZN(n6751) );
  OR2_X2 U18742 ( .A1(n6752), .A2(n6751), .ZN(n48074) );
  NAND2_X1 U18743 ( .A1(n46628), .A2(n6754), .ZN(n6753) );
  INV_X1 U18744 ( .A(n44421), .ZN(n6754) );
  NAND2_X1 U18746 ( .A1(n8645), .A2(n8646), .ZN(n6757) );
  NAND2_X1 U18747 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  NAND2_X1 U18748 ( .A1(n33016), .A2(n26634), .ZN(n6759) );
  NAND2_X1 U18750 ( .A1(n28530), .A2(n28874), .ZN(n6764) );
  NAND2_X1 U18751 ( .A1(n28875), .A2(n28883), .ZN(n6765) );
  INV_X1 U18752 ( .A(n41641), .ZN(n41643) );
  NAND2_X2 U18753 ( .A1(n6766), .A2(n6767), .ZN(n41647) );
  NAND3_X1 U18754 ( .A1(n34689), .A2(n34687), .A3(n34688), .ZN(n6767) );
  NOR2_X1 U18755 ( .A1(n30429), .A2(n30433), .ZN(n6768) );
  AOI22_X1 U18756 ( .A1(n728), .A2(n6768), .B1(n6771), .B2(n6770), .ZN(n6769)
         );
  INV_X1 U18757 ( .A(n30424), .ZN(n30427) );
  NAND2_X1 U18758 ( .A1(n29867), .A2(n51746), .ZN(n30424) );
  XNOR2_X1 U18760 ( .A(n6773), .B(n25646), .ZN(n24963) );
  XNOR2_X1 U18761 ( .A(n24303), .B(n6773), .ZN(n24304) );
  XNOR2_X1 U18762 ( .A(n26106), .B(n6773), .ZN(n26107) );
  XNOR2_X1 U18763 ( .A(n27452), .B(n6773), .ZN(n25638) );
  XNOR2_X1 U18764 ( .A(n25425), .B(n6773), .ZN(n25917) );
  NAND3_X1 U18765 ( .A1(n8577), .A2(n8578), .A3(n38196), .ZN(n6774) );
  NAND3_X1 U18766 ( .A1(n689), .A2(n38204), .A3(n38576), .ZN(n6778) );
  NAND2_X1 U18767 ( .A1(n35146), .A2(n6781), .ZN(n6780) );
  NAND2_X1 U18768 ( .A1(n38573), .A2(n36098), .ZN(n6784) );
  NAND2_X1 U18769 ( .A1(n32672), .A2(n32671), .ZN(n6785) );
  INV_X1 U18770 ( .A(n21186), .ZN(n21178) );
  NAND2_X1 U18772 ( .A1(n48649), .A2(n6787), .ZN(n48561) );
  NAND2_X1 U18773 ( .A1(n48638), .A2(n48581), .ZN(n6787) );
  NAND2_X1 U18774 ( .A1(n6788), .A2(n48647), .ZN(n48581) );
  NAND2_X1 U18775 ( .A1(n31546), .A2(n31538), .ZN(n31443) );
  NAND4_X2 U18776 ( .A1(n6792), .A2(n6791), .A3(n6790), .A4(n6789), .ZN(n31538) );
  NAND2_X1 U18777 ( .A1(n30787), .A2(n26829), .ZN(n6790) );
  AND3_X1 U18778 ( .A1(n13853), .A2(n6793), .A3(n14473), .ZN(n13561) );
  NAND3_X1 U18779 ( .A1(n11735), .A2(n11734), .A3(n6794), .ZN(n11748) );
  NAND2_X1 U18780 ( .A1(n36467), .A2(n38332), .ZN(n6795) );
  NAND2_X1 U18781 ( .A1(n6798), .A2(n6797), .ZN(n13392) );
  NAND3_X1 U18782 ( .A1(n5099), .A2(n14527), .A3(n6192), .ZN(n6797) );
  NAND2_X1 U18783 ( .A1(n13392), .A2(n13035), .ZN(n13043) );
  INV_X1 U18784 ( .A(n14520), .ZN(n14528) );
  INV_X1 U18785 ( .A(n13034), .ZN(n6799) );
  XNOR2_X1 U18787 ( .A(n6801), .B(n48614), .ZN(Plaintext[57]) );
  NAND4_X1 U18788 ( .A1(n6806), .A2(n48610), .A3(n6805), .A4(n6802), .ZN(n6801) );
  NAND2_X1 U18789 ( .A1(n48622), .A2(n52042), .ZN(n6803) );
  OR2_X1 U18790 ( .A1(n48622), .A2(n48612), .ZN(n6804) );
  XNOR2_X1 U18791 ( .A(n25649), .B(n25639), .ZN(n6808) );
  NAND2_X1 U18793 ( .A1(n31827), .A2(n6809), .ZN(n26709) );
  XNOR2_X2 U18794 ( .A(n45344), .B(n45345), .ZN(n48531) );
  NAND2_X1 U18795 ( .A1(n46984), .A2(n50363), .ZN(n50360) );
  AND2_X1 U18796 ( .A1(n49599), .A2(n49598), .ZN(n6814) );
  NAND2_X1 U18797 ( .A1(n6816), .A2(n50888), .ZN(n6815) );
  NAND2_X1 U18798 ( .A1(n50851), .A2(n6818), .ZN(n6816) );
  NOR2_X1 U18799 ( .A1(n21458), .A2(n21474), .ZN(n6819) );
  NAND2_X1 U18800 ( .A1(n41319), .A2(n40730), .ZN(n41320) );
  AND3_X2 U18801 ( .A1(n6821), .A2(n38579), .A3(n6820), .ZN(n40730) );
  NAND2_X1 U18802 ( .A1(n38574), .A2(n38573), .ZN(n6821) );
  NAND2_X1 U18803 ( .A1(n31548), .A2(n31549), .ZN(n7393) );
  NAND2_X1 U18804 ( .A1(n13971), .A2(n5540), .ZN(n13215) );
  XNOR2_X1 U18805 ( .A(n26448), .B(n24936), .ZN(n24144) );
  NOR2_X2 U18806 ( .A1(n22309), .A2(n6822), .ZN(n24936) );
  NAND2_X1 U18807 ( .A1(n46877), .A2(n6823), .ZN(n46879) );
  NAND2_X1 U18808 ( .A1(n47089), .A2(n2159), .ZN(n6823) );
  XNOR2_X1 U18809 ( .A(n6826), .B(n37292), .ZN(n34043) );
  XNOR2_X1 U18810 ( .A(n34434), .B(n6826), .ZN(n34435) );
  XNOR2_X1 U18811 ( .A(n34855), .B(n6826), .ZN(n34857) );
  XNOR2_X1 U18812 ( .A(n34856), .B(n6826), .ZN(n37091) );
  XNOR2_X1 U18813 ( .A(n6826), .B(n36983), .ZN(n35546) );
  XNOR2_X1 U18814 ( .A(n6826), .B(n33526), .ZN(n34350) );
  INV_X1 U18816 ( .A(n6828), .ZN(n6827) );
  AOI21_X1 U18817 ( .B1(n40442), .B2(n2854), .A(n6830), .ZN(n6829) );
  NOR2_X1 U18818 ( .A1(n6851), .A2(n40402), .ZN(n6830) );
  INV_X1 U18819 ( .A(n47617), .ZN(n6831) );
  XNOR2_X1 U18820 ( .A(n35351), .B(n35350), .ZN(n6832) );
  NAND2_X1 U18821 ( .A1(n13764), .A2(n14145), .ZN(n6834) );
  NAND2_X1 U18822 ( .A1(n7475), .A2(n26724), .ZN(n6836) );
  NAND2_X1 U18823 ( .A1(n26720), .A2(n29441), .ZN(n6838) );
  NAND2_X1 U18824 ( .A1(n10197), .A2(n10196), .ZN(n6841) );
  NOR2_X1 U18825 ( .A1(n51403), .A2(n20144), .ZN(n19062) );
  NAND4_X2 U18826 ( .A1(n17307), .A2(n6843), .A3(n17306), .A4(n17308), .ZN(
        n22639) );
  NAND3_X1 U18827 ( .A1(n19782), .A2(n19783), .A3(n2182), .ZN(n6843) );
  NAND2_X1 U18828 ( .A1(n20156), .A2(n19535), .ZN(n17090) );
  NAND2_X1 U18829 ( .A1(n6848), .A2(n51508), .ZN(n6847) );
  INV_X1 U18830 ( .A(n8909), .ZN(n6849) );
  NAND2_X1 U18831 ( .A1(n6849), .A2(n12464), .ZN(n12451) );
  XNOR2_X2 U18832 ( .A(n8897), .B(Key[133]), .ZN(n12464) );
  INV_X1 U18833 ( .A(n6852), .ZN(n6850) );
  NAND3_X2 U18834 ( .A1(n7210), .A2(n7213), .A3(n44782), .ZN(n49112) );
  INV_X1 U18835 ( .A(n25198), .ZN(n25199) );
  INV_X1 U18836 ( .A(n30178), .ZN(n6853) );
  NAND2_X1 U18837 ( .A1(n29616), .A2(n29618), .ZN(n28607) );
  NAND2_X1 U18838 ( .A1(n28030), .A2(n30164), .ZN(n6854) );
  NAND2_X1 U18839 ( .A1(n28029), .A2(n30167), .ZN(n6855) );
  XNOR2_X1 U18840 ( .A(n34454), .B(n34453), .ZN(n6856) );
  NAND2_X1 U18841 ( .A1(n40009), .A2(n39094), .ZN(n6859) );
  NOR2_X1 U18842 ( .A1(n38416), .A2(n6861), .ZN(n6860) );
  INV_X1 U18843 ( .A(n39995), .ZN(n6861) );
  NAND2_X1 U18844 ( .A1(n12667), .A2(n11874), .ZN(n12674) );
  OR2_X1 U18845 ( .A1(n35422), .A2(n37629), .ZN(n6862) );
  NAND2_X1 U18846 ( .A1(n38276), .A2(n38272), .ZN(n35424) );
  OAI211_X1 U18848 ( .C1(n20415), .C2(n5923), .A(n6864), .B(n21397), .ZN(
        n20377) );
  NAND2_X1 U18849 ( .A1(n20376), .A2(n581), .ZN(n6865) );
  NAND2_X1 U18850 ( .A1(n724), .A2(n31300), .ZN(n31312) );
  NAND3_X1 U18851 ( .A1(n24778), .A2(n24777), .A3(n6867), .ZN(n6866) );
  NAND3_X1 U18852 ( .A1(n19782), .A2(n6868), .A3(n19783), .ZN(n19790) );
  NAND2_X1 U18854 ( .A1(n8441), .A2(n19023), .ZN(n21283) );
  INV_X1 U18855 ( .A(n36105), .ZN(n6869) );
  NOR2_X1 U18856 ( .A1(n11853), .A2(n14485), .ZN(n7733) );
  NAND2_X1 U18857 ( .A1(n41088), .A2(n39700), .ZN(n39701) );
  NAND2_X1 U18858 ( .A1(n41083), .A2(n39704), .ZN(n6870) );
  OAI21_X1 U18859 ( .B1(n51396), .B2(n41469), .A(n6871), .ZN(n41478) );
  NAND4_X1 U18860 ( .A1(n41410), .A2(n44845), .A3(n51317), .A4(n46583), .ZN(
        n6871) );
  NAND2_X1 U18861 ( .A1(n6874), .A2(n6873), .ZN(n6872) );
  NAND3_X1 U18862 ( .A1(n27894), .A2(n29329), .A3(n27893), .ZN(n6874) );
  NAND2_X1 U18863 ( .A1(n21953), .A2(n51250), .ZN(n21167) );
  NAND2_X1 U18866 ( .A1(n33427), .A2(n36189), .ZN(n33453) );
  NAND2_X1 U18867 ( .A1(n39335), .A2(n33461), .ZN(n33427) );
  NAND2_X1 U18868 ( .A1(n46276), .A2(n6879), .ZN(n45693) );
  INV_X1 U18869 ( .A(n45237), .ZN(n6879) );
  INV_X1 U18870 ( .A(n45237), .ZN(n46354) );
  XNOR2_X2 U18871 ( .A(n42573), .B(n42574), .ZN(n45237) );
  XNOR2_X2 U18872 ( .A(n8563), .B(Key[60]), .ZN(n12301) );
  NOR2_X1 U18873 ( .A1(n6882), .A2(n6880), .ZN(n35439) );
  NAND2_X1 U18875 ( .A1(n6885), .A2(n6884), .ZN(n6883) );
  NAND2_X1 U18876 ( .A1(n38428), .A2(n40014), .ZN(n6886) );
  INV_X1 U18877 ( .A(n31088), .ZN(n6892) );
  NAND2_X1 U18878 ( .A1(n29688), .A2(n6892), .ZN(n6890) );
  NAND2_X1 U18879 ( .A1(n30912), .A2(n30593), .ZN(n6895) );
  NAND2_X1 U18880 ( .A1(n31086), .A2(n6894), .ZN(n6893) );
  NAND2_X1 U18881 ( .A1(n30910), .A2(n6895), .ZN(n6894) );
  NAND2_X1 U18882 ( .A1(n6897), .A2(n21733), .ZN(n6896) );
  NAND2_X1 U18883 ( .A1(n20865), .A2(n22261), .ZN(n6897) );
  NAND2_X1 U18884 ( .A1(n6899), .A2(n23342), .ZN(n6898) );
  INV_X1 U18885 ( .A(n21140), .ZN(n6899) );
  XNOR2_X1 U18886 ( .A(n35032), .B(n6900), .ZN(n34187) );
  XNOR2_X1 U18887 ( .A(n6901), .B(n34000), .ZN(n6900) );
  XNOR2_X1 U18888 ( .A(n33186), .B(n6902), .ZN(n6901) );
  INV_X1 U18889 ( .A(n20613), .ZN(n6903) );
  XNOR2_X2 U18890 ( .A(n16077), .B(n16076), .ZN(n16125) );
  NAND4_X2 U18891 ( .A1(n38099), .A2(n38100), .A3(n38097), .A4(n38098), .ZN(
        n40081) );
  NAND2_X1 U18894 ( .A1(n10438), .A2(n11943), .ZN(n6910) );
  NAND2_X1 U18895 ( .A1(n11943), .A2(n6912), .ZN(n6911) );
  NAND3_X1 U18896 ( .A1(n6914), .A2(n441), .A3(n21873), .ZN(n6915) );
  NAND2_X1 U18897 ( .A1(n22964), .A2(n756), .ZN(n6913) );
  INV_X1 U18898 ( .A(n6915), .ZN(n22255) );
  NAND2_X1 U18899 ( .A1(n441), .A2(n21873), .ZN(n21863) );
  NOR2_X1 U18900 ( .A1(n6916), .A2(n51746), .ZN(n29707) );
  NAND2_X1 U18901 ( .A1(n6916), .A2(n486), .ZN(n27514) );
  AND2_X1 U18902 ( .A1(n30436), .A2(n6916), .ZN(n30437) );
  MUX2_X1 U18903 ( .A(n30436), .B(n29703), .S(n6916), .Z(n29702) );
  NOR2_X1 U18904 ( .A1(n29863), .A2(n6916), .ZN(n29875) );
  OAI22_X1 U18905 ( .A1(n28328), .A2(n29866), .B1(n28332), .B2(n6916), .ZN(
        n28331) );
  NAND2_X1 U18906 ( .A1(n23536), .A2(n3816), .ZN(n23537) );
  XNOR2_X2 U18907 ( .A(n44505), .B(n6918), .ZN(n50280) );
  XNOR2_X1 U18908 ( .A(n41969), .B(n51420), .ZN(n43936) );
  NAND2_X1 U18909 ( .A1(n18875), .A2(n20671), .ZN(n20669) );
  NAND3_X1 U18910 ( .A1(n18875), .A2(n20671), .A3(n20228), .ZN(n6919) );
  XNOR2_X1 U18912 ( .A(n7556), .B(n6921), .ZN(n32273) );
  XNOR2_X1 U18913 ( .A(n6921), .B(n35237), .ZN(n34759) );
  XNOR2_X1 U18914 ( .A(n34331), .B(n6921), .ZN(n34336) );
  XNOR2_X1 U18915 ( .A(n30337), .B(n6921), .ZN(n30501) );
  XNOR2_X1 U18916 ( .A(n33210), .B(n6921), .ZN(n33211) );
  XNOR2_X1 U18917 ( .A(n6922), .B(n25429), .ZN(n22695) );
  NAND2_X1 U18918 ( .A1(n20287), .A2(n43702), .ZN(n6923) );
  NAND2_X1 U18919 ( .A1(n20288), .A2(n43702), .ZN(n6924) );
  XNOR2_X1 U18920 ( .A(n26092), .B(n6926), .ZN(n28302) );
  XNOR2_X1 U18921 ( .A(n26092), .B(n6927), .ZN(n28439) );
  NAND4_X2 U18922 ( .A1(n31653), .A2(n8546), .A3(n31652), .A4(n8545), .ZN(
        n36747) );
  INV_X1 U18923 ( .A(n24244), .ZN(n21822) );
  NAND4_X2 U18924 ( .A1(n20206), .A2(n20205), .A3(n20203), .A4(n20204), .ZN(
        n21820) );
  NAND3_X2 U18925 ( .A1(n25852), .A2(n25851), .A3(n25854), .ZN(n31873) );
  NAND4_X2 U18926 ( .A1(n25517), .A2(n25519), .A3(n7683), .A4(n25518), .ZN(
        n31876) );
  XNOR2_X2 U18927 ( .A(n25221), .B(n25220), .ZN(n27987) );
  NAND3_X1 U18929 ( .A1(n21319), .A2(n19549), .A3(n20903), .ZN(n22003) );
  OR2_X2 U18930 ( .A1(n19502), .A2(n19501), .ZN(n22586) );
  NAND2_X1 U18931 ( .A1(n19515), .A2(n19514), .ZN(n6931) );
  NAND2_X1 U18932 ( .A1(n19516), .A2(n52065), .ZN(n6932) );
  XNOR2_X2 U18933 ( .A(n18534), .B(n17213), .ZN(n18394) );
  NAND2_X1 U18935 ( .A1(n14307), .A2(n14311), .ZN(n14310) );
  NAND3_X1 U18936 ( .A1(n14307), .A2(n14311), .A3(n14320), .ZN(n14314) );
  NAND2_X1 U18937 ( .A1(n31645), .A2(n32724), .ZN(n8548) );
  NAND3_X1 U18938 ( .A1(n16128), .A2(n16863), .A3(n6936), .ZN(n6934) );
  NAND2_X1 U18939 ( .A1(n21527), .A2(n7160), .ZN(n16865) );
  NAND3_X1 U18941 ( .A1(n21528), .A2(n21525), .A3(n18895), .ZN(n6936) );
  NAND3_X1 U18942 ( .A1(n28745), .A2(n30425), .A3(n30433), .ZN(n29691) );
  INV_X1 U18943 ( .A(n30431), .ZN(n30433) );
  INV_X1 U18945 ( .A(n15196), .ZN(n15200) );
  XNOR2_X1 U18947 ( .A(n33171), .B(n33170), .ZN(n6937) );
  INV_X1 U18949 ( .A(n30833), .ZN(n30649) );
  NAND2_X1 U18950 ( .A1(n31306), .A2(n31300), .ZN(n30833) );
  NAND2_X1 U18951 ( .A1(n41642), .A2(n41650), .ZN(n41104) );
  OAI21_X1 U18952 ( .B1(n6942), .B2(n45927), .A(n49277), .ZN(n45935) );
  XNOR2_X1 U18953 ( .A(n6944), .B(n51441), .ZN(n6943) );
  INV_X1 U18954 ( .A(n10742), .ZN(n10734) );
  NAND2_X1 U18955 ( .A1(n8994), .A2(n11341), .ZN(n12245) );
  NAND2_X1 U18956 ( .A1(n6946), .A2(n633), .ZN(n6954) );
  NAND3_X1 U18957 ( .A1(n18292), .A2(n20020), .A3(n6947), .ZN(n6946) );
  NAND2_X1 U18958 ( .A1(n2166), .A2(n16797), .ZN(n6947) );
  NOR2_X1 U18959 ( .A1(n17516), .A2(n633), .ZN(n6948) );
  AOI21_X1 U18960 ( .B1(n17529), .B2(n6951), .A(n6950), .ZN(n6955) );
  NAND2_X1 U18961 ( .A1(n20010), .A2(n16801), .ZN(n6950) );
  NAND2_X1 U18962 ( .A1(n48974), .A2(n48954), .ZN(n48929) );
  NAND2_X2 U18963 ( .A1(n6958), .A2(n6956), .ZN(n50483) );
  NAND2_X1 U18964 ( .A1(n50362), .A2(n6957), .ZN(n6956) );
  NAND2_X1 U18965 ( .A1(n46971), .A2(n47144), .ZN(n50359) );
  NAND3_X1 U18966 ( .A1(n39095), .A2(n6962), .A3(n39099), .ZN(n38423) );
  NAND2_X1 U18967 ( .A1(n40011), .A2(n6963), .ZN(n38426) );
  NOR2_X1 U18968 ( .A1(n6965), .A2(n39667), .ZN(n6963) );
  NAND2_X1 U18970 ( .A1(n32204), .A2(n6969), .ZN(n30889) );
  OAI21_X1 U18971 ( .B1(n29158), .B2(n29156), .A(n26486), .ZN(n24990) );
  NAND2_X1 U18972 ( .A1(n5821), .A2(n6970), .ZN(n26486) );
  XNOR2_X2 U18974 ( .A(n18824), .B(n6972), .ZN(n21351) );
  XNOR2_X1 U18975 ( .A(n6973), .B(n18699), .ZN(n6972) );
  XNOR2_X1 U18976 ( .A(n18700), .B(n18698), .ZN(n6973) );
  XNOR2_X1 U18978 ( .A(n6975), .B(n35229), .ZN(n6974) );
  XNOR2_X1 U18979 ( .A(n6976), .B(n35228), .ZN(n6975) );
  XNOR2_X1 U18980 ( .A(n37077), .B(n36986), .ZN(n6976) );
  OAI22_X1 U18981 ( .A1(n38640), .A2(n38257), .B1(n37224), .B2(n6977), .ZN(
        n6978) );
  NAND2_X1 U18982 ( .A1(n37688), .A2(n2188), .ZN(n6977) );
  INV_X1 U18983 ( .A(n37224), .ZN(n38264) );
  OAI21_X1 U18984 ( .B1(n38632), .B2(n5989), .A(n6978), .ZN(n35302) );
  NAND2_X1 U18985 ( .A1(n6979), .A2(n11598), .ZN(n11602) );
  NAND2_X1 U18986 ( .A1(n11591), .A2(n11613), .ZN(n6979) );
  INV_X1 U18987 ( .A(n11608), .ZN(n9278) );
  INV_X1 U18988 ( .A(n30241), .ZN(n30240) );
  NAND2_X1 U18989 ( .A1(n29038), .A2(n29039), .ZN(n29040) );
  NAND2_X1 U18990 ( .A1(n35940), .A2(n36186), .ZN(n6981) );
  NAND3_X1 U18991 ( .A1(n6983), .A2(n33035), .A3(n32883), .ZN(n31527) );
  NAND2_X1 U18992 ( .A1(n32885), .A2(n6984), .ZN(n6983) );
  NAND2_X1 U18993 ( .A1(n33041), .A2(n32879), .ZN(n32885) );
  INV_X1 U18995 ( .A(n49635), .ZN(n50292) );
  NAND2_X1 U18996 ( .A1(n52172), .A2(n6986), .ZN(n48332) );
  NAND3_X1 U18997 ( .A1(n6987), .A2(n51728), .A3(n48381), .ZN(n48281) );
  NAND2_X1 U18998 ( .A1(n8104), .A2(n6987), .ZN(n48296) );
  NAND2_X1 U18999 ( .A1(n51087), .A2(n6987), .ZN(n48376) );
  INV_X1 U19000 ( .A(n32645), .ZN(n31533) );
  NAND2_X1 U19001 ( .A1(n44680), .A2(n6988), .ZN(n44683) );
  NOR2_X1 U19002 ( .A1(n46458), .A2(n604), .ZN(n6988) );
  INV_X1 U19003 ( .A(n44678), .ZN(n48247) );
  NAND2_X1 U19005 ( .A1(n40794), .A2(n51358), .ZN(n6998) );
  NAND2_X1 U19006 ( .A1(n7000), .A2(n51357), .ZN(n6999) );
  INV_X1 U19007 ( .A(n7282), .ZN(n7003) );
  AOI21_X1 U19008 ( .B1(n38495), .B2(n7004), .A(n38494), .ZN(n38497) );
  AND2_X1 U19009 ( .A1(n35953), .A2(n38492), .ZN(n35571) );
  NAND2_X1 U19010 ( .A1(n37392), .A2(n7004), .ZN(n37393) );
  NOR2_X1 U19011 ( .A1(n35950), .A2(n7004), .ZN(n35576) );
  XNOR2_X1 U19012 ( .A(n43520), .B(n43518), .ZN(n7005) );
  NAND2_X1 U19013 ( .A1(n23657), .A2(n23656), .ZN(n7008) );
  NAND2_X1 U19014 ( .A1(n7010), .A2(n21397), .ZN(n7009) );
  OAI22_X1 U19015 ( .A1(n21393), .A2(n21374), .B1(n20794), .B2(n1860), .ZN(
        n7010) );
  NAND2_X1 U19017 ( .A1(n37554), .A2(n2364), .ZN(n35929) );
  XNOR2_X1 U19018 ( .A(n51057), .B(n7012), .ZN(n23286) );
  NAND2_X1 U19020 ( .A1(n27570), .A2(n7013), .ZN(n29896) );
  AND2_X1 U19021 ( .A1(n26828), .A2(n7014), .ZN(n7013) );
  INV_X1 U19022 ( .A(n27566), .ZN(n7014) );
  OR2_X1 U19023 ( .A1(n681), .A2(n7015), .ZN(n7860) );
  NAND2_X1 U19024 ( .A1(n6046), .A2(n40785), .ZN(n7015) );
  OAI21_X1 U19025 ( .B1(n7018), .B2(n7016), .A(n2192), .ZN(n43493) );
  NAND2_X1 U19026 ( .A1(n49506), .A2(n7017), .ZN(n7016) );
  NOR2_X1 U19027 ( .A1(n43491), .A2(n49534), .ZN(n7018) );
  OR2_X1 U19028 ( .A1(n5335), .A2(n10722), .ZN(n7081) );
  NOR2_X1 U19029 ( .A1(n12285), .A2(n5335), .ZN(n10720) );
  NAND2_X1 U19030 ( .A1(n12291), .A2(n5335), .ZN(n10226) );
  NAND2_X1 U19031 ( .A1(n8480), .A2(n551), .ZN(n39281) );
  OAI21_X1 U19032 ( .B1(n39283), .B2(n39282), .A(n39281), .ZN(n7022) );
  INV_X1 U19033 ( .A(n39369), .ZN(n7026) );
  INV_X1 U19035 ( .A(n7034), .ZN(n41674) );
  NAND2_X1 U19036 ( .A1(n41678), .A2(n7034), .ZN(n7031) );
  NAND2_X1 U19037 ( .A1(n41677), .A2(n41676), .ZN(n7029) );
  OAI21_X1 U19038 ( .B1(n41668), .B2(n41669), .A(n6335), .ZN(n7032) );
  NAND2_X1 U19039 ( .A1(n41684), .A2(n41685), .ZN(n7033) );
  XNOR2_X2 U19040 ( .A(n43107), .B(n7035), .ZN(n49990) );
  INV_X1 U19041 ( .A(n19076), .ZN(n19064) );
  NAND3_X1 U19042 ( .A1(n19075), .A2(n19064), .A3(n7845), .ZN(n7037) );
  NAND4_X1 U19043 ( .A1(n41423), .A2(n41422), .A3(n41421), .A4(n7039), .ZN(
        n41758) );
  MUX2_X1 U19044 ( .A(n41411), .B(n42000), .S(n41580), .Z(n7039) );
  NAND2_X1 U19045 ( .A1(n13827), .A2(n13819), .ZN(n13817) );
  NAND2_X1 U19046 ( .A1(n435), .A2(n31746), .ZN(n7040) );
  NAND2_X1 U19047 ( .A1(n7226), .A2(n28918), .ZN(n7042) );
  NAND2_X1 U19048 ( .A1(n28989), .A2(n7042), .ZN(n29025) );
  NOR2_X1 U19049 ( .A1(n7043), .A2(n23153), .ZN(n21960) );
  OR2_X1 U19050 ( .A1(n7044), .A2(n2159), .ZN(n47108) );
  INV_X1 U19051 ( .A(n46869), .ZN(n7044) );
  NAND2_X1 U19052 ( .A1(n5953), .A2(n7045), .ZN(n20778) );
  XNOR2_X2 U19053 ( .A(n8787), .B(Key[79]), .ZN(n8796) );
  INV_X1 U19054 ( .A(n44109), .ZN(n7046) );
  INV_X1 U19055 ( .A(n44109), .ZN(n7047) );
  INV_X1 U19056 ( .A(n44458), .ZN(n46781) );
  INV_X1 U19057 ( .A(n19514), .ZN(n7050) );
  NAND2_X1 U19058 ( .A1(n16677), .A2(n6226), .ZN(n19513) );
  NAND2_X1 U19059 ( .A1(n17039), .A2(n19503), .ZN(n7049) );
  OAI21_X1 U19060 ( .B1(n29271), .B2(n29282), .A(n8424), .ZN(n7051) );
  INV_X1 U19061 ( .A(n28710), .ZN(n7052) );
  XNOR2_X2 U19062 ( .A(Key[91]), .B(Ciphertext[42]), .ZN(n12690) );
  INV_X2 U19063 ( .A(n12205), .ZN(n12198) );
  NAND2_X1 U19064 ( .A1(n14280), .A2(n14294), .ZN(n13013) );
  INV_X1 U19066 ( .A(n8793), .ZN(n7054) );
  NAND3_X1 U19067 ( .A1(n8798), .A2(n8797), .A3(n12367), .ZN(n7055) );
  NAND2_X1 U19068 ( .A1(n32175), .A2(n32957), .ZN(n32964) );
  OR2_X2 U19069 ( .A1(n28209), .A2(n28210), .ZN(n32957) );
  NAND2_X2 U19070 ( .A1(n7061), .A2(n46527), .ZN(n48702) );
  NAND2_X1 U19071 ( .A1(n48169), .A2(n46521), .ZN(n7062) );
  NAND2_X1 U19072 ( .A1(n46520), .A2(n1752), .ZN(n7063) );
  NAND2_X1 U19073 ( .A1(n40899), .A2(n40276), .ZN(n39582) );
  NAND3_X1 U19074 ( .A1(n2224), .A2(n40269), .A3(n40903), .ZN(n40276) );
  NAND2_X2 U19076 ( .A1(n7065), .A2(n30239), .ZN(n32608) );
  NAND2_X1 U19079 ( .A1(n35027), .A2(n35026), .ZN(n7068) );
  NAND2_X1 U19080 ( .A1(n7070), .A2(n38192), .ZN(n7069) );
  NOR2_X1 U19081 ( .A1(n24157), .A2(n1942), .ZN(n7077) );
  NAND4_X2 U19082 ( .A1(n32833), .A2(n32834), .A3(n32835), .A4(n7078), .ZN(
        n36991) );
  NAND2_X1 U19083 ( .A1(n32831), .A2(n32832), .ZN(n7078) );
  XNOR2_X2 U19084 ( .A(n42507), .B(n42506), .ZN(n48461) );
  NAND4_X2 U19085 ( .A1(n9448), .A2(n9449), .A3(n9446), .A4(n9447), .ZN(n7079)
         );
  XNOR2_X1 U19086 ( .A(n16701), .B(n7079), .ZN(n16534) );
  XNOR2_X1 U19087 ( .A(n7079), .B(n19248), .ZN(n17802) );
  XNOR2_X1 U19088 ( .A(n17938), .B(n7079), .ZN(n17651) );
  XNOR2_X1 U19089 ( .A(n7079), .B(n17365), .ZN(n14510) );
  NAND2_X1 U19090 ( .A1(n8353), .A2(n22765), .ZN(n22767) );
  NAND3_X1 U19092 ( .A1(n29229), .A2(n29230), .A3(n30256), .ZN(n7082) );
  INV_X1 U19093 ( .A(n8796), .ZN(n12350) );
  NAND2_X1 U19094 ( .A1(n12358), .A2(n12359), .ZN(n10985) );
  INV_X1 U19096 ( .A(n7607), .ZN(n48873) );
  NOR2_X1 U19097 ( .A1(n48905), .A2(n7085), .ZN(n7084) );
  NAND2_X1 U19098 ( .A1(n48913), .A2(n48862), .ZN(n7085) );
  NAND2_X1 U19099 ( .A1(n30267), .A2(n52147), .ZN(n29226) );
  INV_X1 U19100 ( .A(n19009), .ZN(n21197) );
  NAND2_X1 U19102 ( .A1(n29592), .A2(n7089), .ZN(n30062) );
  INV_X1 U19103 ( .A(n29588), .ZN(n7088) );
  NAND4_X1 U19104 ( .A1(n7092), .A2(n7090), .A3(n30062), .A4(n7087), .ZN(n7091) );
  NAND2_X1 U19105 ( .A1(n30946), .A2(n7088), .ZN(n7087) );
  AND2_X1 U19106 ( .A1(n362), .A2(n29591), .ZN(n7089) );
  NAND2_X1 U19107 ( .A1(n30946), .A2(n29592), .ZN(n7090) );
  NAND2_X1 U19108 ( .A1(n31115), .A2(n7093), .ZN(n7092) );
  XNOR2_X1 U19109 ( .A(n15018), .B(n2375), .ZN(n17966) );
  XNOR2_X1 U19110 ( .A(n15018), .B(n2355), .ZN(n15504) );
  NAND2_X1 U19111 ( .A1(n766), .A2(n5388), .ZN(n21294) );
  NAND2_X1 U19112 ( .A1(n19720), .A2(n19796), .ZN(n7100) );
  INV_X1 U19113 ( .A(n7102), .ZN(n37876) );
  XNOR2_X2 U19114 ( .A(n43696), .B(n41302), .ZN(n7102) );
  XNOR2_X1 U19115 ( .A(n37876), .B(n7101), .ZN(n45265) );
  XNOR2_X1 U19116 ( .A(n7102), .B(n45250), .ZN(n42449) );
  NAND2_X1 U19118 ( .A1(n22175), .A2(n21712), .ZN(n7104) );
  OAI21_X1 U19119 ( .B1(n40599), .B2(n40600), .A(n7105), .ZN(n7107) );
  INV_X1 U19120 ( .A(n52202), .ZN(n7110) );
  XNOR2_X2 U19121 ( .A(n44187), .B(n44186), .ZN(n46471) );
  NAND4_X1 U19122 ( .A1(n19564), .A2(n22140), .A3(n22144), .A4(n51660), .ZN(
        n7111) );
  NAND2_X1 U19123 ( .A1(n50466), .A2(n50485), .ZN(n7112) );
  XNOR2_X1 U19125 ( .A(n7115), .B(n51436), .ZN(n15658) );
  XNOR2_X1 U19126 ( .A(n637), .B(n7115), .ZN(n16270) );
  XNOR2_X1 U19127 ( .A(n7115), .B(n15821), .ZN(n15822) );
  XNOR2_X1 U19128 ( .A(n16730), .B(n7115), .ZN(n16200) );
  XNOR2_X1 U19129 ( .A(n7115), .B(n16963), .ZN(n18161) );
  NOR2_X1 U19130 ( .A1(n7435), .A2(n7434), .ZN(n7116) );
  OAI21_X1 U19131 ( .B1(n39857), .B2(n40329), .A(n39643), .ZN(n37864) );
  NAND2_X1 U19132 ( .A1(n19917), .A2(n7119), .ZN(n20564) );
  NAND2_X1 U19133 ( .A1(n7120), .A2(n40874), .ZN(n40875) );
  MUX2_X1 U19134 ( .A(n40546), .B(n40547), .S(n39968), .Z(n40548) );
  XNOR2_X1 U19135 ( .A(n7121), .B(n46137), .ZN(n43516) );
  XNOR2_X1 U19136 ( .A(n7121), .B(n42758), .ZN(n42759) );
  XNOR2_X1 U19137 ( .A(n7121), .B(n46143), .ZN(n46152) );
  NOR2_X1 U19138 ( .A1(n52147), .A2(n7124), .ZN(n7123) );
  NAND2_X1 U19139 ( .A1(n25107), .A2(n27918), .ZN(n7124) );
  XNOR2_X1 U19140 ( .A(n15541), .B(n15540), .ZN(n7125) );
  AND2_X1 U19141 ( .A1(n20503), .A2(n18085), .ZN(n17589) );
  NAND2_X1 U19144 ( .A1(n13481), .A2(n15045), .ZN(n13482) );
  NAND2_X1 U19145 ( .A1(n7128), .A2(n13136), .ZN(n14188) );
  NAND3_X1 U19146 ( .A1(n7130), .A2(n20087), .A3(n7131), .ZN(n7129) );
  NAND3_X1 U19147 ( .A1(n17603), .A2(n20086), .A3(n17503), .ZN(n7130) );
  NAND2_X1 U19148 ( .A1(n31781), .A2(n31778), .ZN(n31777) );
  XNOR2_X1 U19149 ( .A(n36677), .B(n34838), .ZN(n7132) );
  NAND2_X1 U19150 ( .A1(n20865), .A2(n22262), .ZN(n7134) );
  NAND2_X1 U19151 ( .A1(n49409), .A2(n47192), .ZN(n47196) );
  OR2_X2 U19152 ( .A1(n49400), .A2(n45926), .ZN(n49465) );
  XNOR2_X2 U19153 ( .A(n33225), .B(n33224), .ZN(n36632) );
  NAND2_X1 U19154 ( .A1(n19140), .A2(n20075), .ZN(n16211) );
  XNOR2_X2 U19155 ( .A(n16198), .B(n7136), .ZN(n20075) );
  NAND2_X1 U19156 ( .A1(n41693), .A2(n41690), .ZN(n7137) );
  AOI21_X1 U19157 ( .B1(n544), .B2(n50486), .A(n50465), .ZN(n7138) );
  OR2_X1 U19158 ( .A1(n7139), .A2(n7138), .ZN(n50373) );
  NAND2_X1 U19160 ( .A1(n7142), .A2(n7141), .ZN(n50291) );
  NAND2_X1 U19161 ( .A1(n50288), .A2(n50287), .ZN(n7142) );
  NAND2_X1 U19162 ( .A1(n39240), .A2(n51063), .ZN(n39219) );
  NAND2_X1 U19164 ( .A1(n24119), .A2(n24117), .ZN(n7144) );
  NAND3_X1 U19165 ( .A1(n28011), .A2(n28010), .A3(n7145), .ZN(n7335) );
  NAND2_X1 U19166 ( .A1(n28604), .A2(n7147), .ZN(n28613) );
  INV_X1 U19167 ( .A(n9239), .ZN(n7148) );
  NAND2_X1 U19168 ( .A1(n9236), .A2(n12169), .ZN(n7149) );
  NAND2_X1 U19169 ( .A1(n40141), .A2(n7488), .ZN(n7153) );
  NAND2_X1 U19170 ( .A1(n40138), .A2(n40139), .ZN(n7154) );
  NAND2_X1 U19171 ( .A1(n40142), .A2(n40143), .ZN(n7155) );
  NAND2_X1 U19172 ( .A1(n11835), .A2(n14223), .ZN(n7157) );
  NAND3_X1 U19173 ( .A1(n40293), .A2(n40295), .A3(n42044), .ZN(n7158) );
  NOR2_X1 U19174 ( .A1(n49047), .A2(n7161), .ZN(n49003) );
  NAND3_X1 U19175 ( .A1(n29149), .A2(n29147), .A3(n29148), .ZN(n29150) );
  NAND2_X1 U19176 ( .A1(n29156), .A2(n7532), .ZN(n29149) );
  AND2_X1 U19180 ( .A1(n29178), .A2(n29177), .ZN(n7165) );
  AND2_X1 U19181 ( .A1(n7430), .A2(n32398), .ZN(n29214) );
  NAND2_X1 U19182 ( .A1(n32080), .A2(n32402), .ZN(n32398) );
  XNOR2_X1 U19183 ( .A(n7166), .B(n51758), .ZN(n17146) );
  XNOR2_X1 U19184 ( .A(n7166), .B(n17906), .ZN(n17907) );
  XNOR2_X1 U19185 ( .A(n462), .B(n7166), .ZN(n14506) );
  NOR2_X2 U19186 ( .A1(n14244), .A2(n13029), .ZN(n7166) );
  NAND2_X1 U19187 ( .A1(n11903), .A2(n11899), .ZN(n11066) );
  NOR2_X1 U19188 ( .A1(n49669), .A2(n50020), .ZN(n7168) );
  NAND3_X1 U19190 ( .A1(n22555), .A2(n19757), .A3(n7170), .ZN(n19766) );
  NAND2_X1 U19191 ( .A1(n22977), .A2(n22434), .ZN(n7170) );
  NAND3_X1 U19193 ( .A1(n35991), .A2(n35990), .A3(n7172), .ZN(n7171) );
  NAND2_X1 U19194 ( .A1(n31624), .A2(n30854), .ZN(n31584) );
  INV_X1 U19195 ( .A(n47282), .ZN(n7175) );
  NAND3_X1 U19196 ( .A1(n7179), .A2(n10963), .A3(n9857), .ZN(n7178) );
  OR2_X1 U19197 ( .A1(n29641), .A2(n31509), .ZN(n7183) );
  AND2_X1 U19198 ( .A1(n22979), .A2(n22434), .ZN(n22558) );
  NAND2_X1 U19199 ( .A1(n19018), .A2(n19782), .ZN(n7186) );
  AND2_X1 U19200 ( .A1(n40768), .A2(n40778), .ZN(n40786) );
  XNOR2_X1 U19201 ( .A(n17691), .B(n7191), .ZN(n17692) );
  XNOR2_X1 U19202 ( .A(n17972), .B(n7191), .ZN(n15990) );
  XNOR2_X1 U19203 ( .A(n15738), .B(n7191), .ZN(n15498) );
  XNOR2_X1 U19204 ( .A(n17381), .B(n7191), .ZN(n18139) );
  XNOR2_X1 U19205 ( .A(n18713), .B(n7191), .ZN(n18715) );
  NAND3_X1 U19206 ( .A1(n10811), .A2(n11593), .A3(n11591), .ZN(n10812) );
  INV_X1 U19207 ( .A(n11611), .ZN(n10815) );
  NAND2_X1 U19208 ( .A1(n51526), .A2(n52143), .ZN(n47368) );
  NOR2_X1 U19209 ( .A1(n20375), .A2(n358), .ZN(n7193) );
  NAND2_X1 U19210 ( .A1(n17981), .A2(n7193), .ZN(n8052) );
  INV_X1 U19211 ( .A(n30663), .ZN(n23859) );
  INV_X1 U19213 ( .A(n26859), .ZN(n23806) );
  NAND2_X1 U19214 ( .A1(n23859), .A2(n30670), .ZN(n26859) );
  XNOR2_X2 U19215 ( .A(n17829), .B(n14239), .ZN(n17381) );
  NAND3_X1 U19216 ( .A1(n10761), .A2(n10762), .A3(n10760), .ZN(n7195) );
  OAI21_X1 U19217 ( .B1(n38974), .B2(n39471), .A(n7196), .ZN(n38975) );
  NOR2_X1 U19218 ( .A1(n38973), .A2(n37809), .ZN(n7197) );
  OAI21_X1 U19219 ( .B1(n39477), .B2(n39476), .A(n7198), .ZN(n39491) );
  XNOR2_X1 U19220 ( .A(n7199), .B(n37324), .ZN(n34153) );
  XNOR2_X1 U19221 ( .A(n7199), .B(n34896), .ZN(n34063) );
  XNOR2_X1 U19222 ( .A(n31811), .B(n7199), .ZN(n31812) );
  INV_X1 U19223 ( .A(n50192), .ZN(n7201) );
  NAND4_X1 U19224 ( .A1(n7203), .A2(n47308), .A3(n47302), .A4(n7202), .ZN(
        n7206) );
  NAND3_X1 U19225 ( .A1(n50299), .A2(n50307), .A3(n7724), .ZN(n7202) );
  NAND2_X1 U19228 ( .A1(n47305), .A2(n47304), .ZN(n7205) );
  NAND2_X1 U19229 ( .A1(n41693), .A2(n41692), .ZN(n41617) );
  NOR2_X1 U19230 ( .A1(n37892), .A2(n2139), .ZN(n34907) );
  NAND2_X1 U19231 ( .A1(n36389), .A2(n38912), .ZN(n7208) );
  INV_X1 U19232 ( .A(n7208), .ZN(n41432) );
  NOR2_X1 U19233 ( .A1(n7209), .A2(n49525), .ZN(n49548) );
  NAND3_X1 U19234 ( .A1(n45929), .A2(n44776), .A3(n7212), .ZN(n7211) );
  NAND2_X1 U19236 ( .A1(n44775), .A2(n49275), .ZN(n45929) );
  INV_X1 U19237 ( .A(n49977), .ZN(n47355) );
  NAND3_X1 U19239 ( .A1(n21407), .A2(n21403), .A3(n20600), .ZN(n20603) );
  OAI211_X1 U19240 ( .C1(n41280), .C2(n52192), .A(n7217), .B(n41285), .ZN(
        n40415) );
  NAND2_X1 U19241 ( .A1(n7218), .A2(n41029), .ZN(n41274) );
  INV_X1 U19242 ( .A(n20604), .ZN(n7219) );
  NAND3_X1 U19243 ( .A1(n38184), .A2(n36365), .A3(n36364), .ZN(n7225) );
  AND2_X1 U19244 ( .A1(n12606), .A2(n12607), .ZN(n7227) );
  XNOR2_X1 U19245 ( .A(n28111), .B(n28112), .ZN(n7229) );
  OAI21_X1 U19246 ( .B1(n32381), .B2(n7230), .A(n32374), .ZN(n32375) );
  NAND2_X1 U19247 ( .A1(n32386), .A2(n30484), .ZN(n32381) );
  NAND2_X1 U19248 ( .A1(n32385), .A2(n32840), .ZN(n7230) );
  NAND3_X1 U19249 ( .A1(n7232), .A2(n32879), .A3(n32867), .ZN(n7231) );
  NAND2_X1 U19251 ( .A1(n19171), .A2(n19332), .ZN(n7233) );
  NAND2_X1 U19252 ( .A1(n19172), .A2(n20434), .ZN(n7234) );
  AOI22_X1 U19253 ( .A1(n12599), .A2(n12598), .B1(n7236), .B2(n12597), .ZN(
        n12608) );
  NAND2_X1 U19254 ( .A1(n3692), .A2(n7235), .ZN(n11917) );
  NAND2_X1 U19255 ( .A1(n11137), .A2(n2395), .ZN(n7235) );
  INV_X1 U19256 ( .A(n11137), .ZN(n7236) );
  NAND3_X1 U19257 ( .A1(n40120), .A2(n36085), .A3(n7239), .ZN(n7238) );
  NAND2_X1 U19258 ( .A1(n36084), .A2(n38769), .ZN(n7241) );
  XNOR2_X1 U19259 ( .A(n7556), .B(n33989), .ZN(n34026) );
  NAND2_X1 U19260 ( .A1(n7243), .A2(n15424), .ZN(n15427) );
  NAND2_X1 U19261 ( .A1(n51023), .A2(n1556), .ZN(n7243) );
  NAND3_X1 U19262 ( .A1(n7246), .A2(n9270), .A3(n13256), .ZN(n9271) );
  OAI21_X1 U19263 ( .B1(n12028), .B2(n14872), .A(n7244), .ZN(n12030) );
  NOR2_X1 U19264 ( .A1(n51023), .A2(n1555), .ZN(n7244) );
  AOI21_X1 U19265 ( .B1(n7246), .B2(n13880), .A(n50966), .ZN(n13884) );
  INV_X1 U19266 ( .A(n51023), .ZN(n7246) );
  NAND2_X1 U19267 ( .A1(n17856), .A2(n20359), .ZN(n19170) );
  XNOR2_X2 U19268 ( .A(n17851), .B(n2318), .ZN(n20359) );
  NAND2_X1 U19269 ( .A1(n27126), .A2(n27131), .ZN(n27986) );
  NAND2_X1 U19270 ( .A1(n7248), .A2(n7247), .ZN(n7523) );
  NAND2_X1 U19271 ( .A1(n20986), .A2(n7249), .ZN(n7248) );
  NAND2_X1 U19272 ( .A1(n20984), .A2(n755), .ZN(n7249) );
  NAND2_X1 U19274 ( .A1(n31224), .A2(n31223), .ZN(n7252) );
  NAND2_X1 U19275 ( .A1(n7253), .A2(n51023), .ZN(n13872) );
  NAND2_X1 U19276 ( .A1(n7259), .A2(n19662), .ZN(n19659) );
  NAND2_X1 U19277 ( .A1(n19664), .A2(n7949), .ZN(n19665) );
  NAND3_X1 U19278 ( .A1(n793), .A2(n51141), .A3(n11411), .ZN(n11398) );
  XNOR2_X1 U19279 ( .A(n7254), .B(n24629), .ZN(n24630) );
  XNOR2_X1 U19280 ( .A(n7254), .B(n26060), .ZN(n26061) );
  XNOR2_X1 U19281 ( .A(n7254), .B(n23401), .ZN(n23402) );
  XNOR2_X1 U19282 ( .A(n7254), .B(n24317), .ZN(n24318) );
  XNOR2_X1 U19283 ( .A(n7351), .B(n7254), .ZN(n25542) );
  NAND4_X1 U19284 ( .A1(n7256), .A2(n19899), .A3(n19888), .A4(n7255), .ZN(
        n7257) );
  NAND2_X1 U19285 ( .A1(n2475), .A2(n19666), .ZN(n7255) );
  NAND2_X1 U19286 ( .A1(n6043), .A2(n15630), .ZN(n19886) );
  OAI21_X1 U19287 ( .B1(n19898), .B2(n19897), .A(n7261), .ZN(n7260) );
  XNOR2_X2 U19288 ( .A(n33924), .B(n33923), .ZN(n37976) );
  OAI21_X1 U19289 ( .B1(n27106), .B2(n28881), .A(n7262), .ZN(n27108) );
  NAND2_X1 U19290 ( .A1(n7263), .A2(n29030), .ZN(n7262) );
  NAND2_X1 U19291 ( .A1(n28882), .A2(n28155), .ZN(n7263) );
  NAND2_X1 U19292 ( .A1(n40649), .A2(n39766), .ZN(n39771) );
  AND2_X1 U19293 ( .A1(n52179), .A2(n49020), .ZN(n49016) );
  NAND4_X2 U19294 ( .A1(n46263), .A2(n46261), .A3(n46260), .A4(n46262), .ZN(
        n49020) );
  XNOR2_X1 U19295 ( .A(n33890), .B(n7271), .ZN(n33999) );
  NAND2_X1 U19296 ( .A1(n7274), .A2(n7272), .ZN(n42516) );
  NAND2_X1 U19297 ( .A1(n48448), .A2(n46448), .ZN(n7273) );
  NAND2_X1 U19298 ( .A1(n7276), .A2(n7275), .ZN(n7274) );
  INV_X2 U19299 ( .A(n48461), .ZN(n7275) );
  NAND3_X1 U19300 ( .A1(n45618), .A2(n46449), .A3(n42489), .ZN(n7276) );
  NAND2_X1 U19301 ( .A1(n7278), .A2(n47480), .ZN(n7277) );
  NAND2_X1 U19302 ( .A1(n47475), .A2(n7279), .ZN(n7278) );
  INV_X1 U19303 ( .A(n3198), .ZN(n7279) );
  AOI21_X1 U19304 ( .B1(n11395), .B2(n2494), .A(n10361), .ZN(n7282) );
  NAND2_X1 U19306 ( .A1(n10734), .A2(n9425), .ZN(n10747) );
  NAND2_X1 U19307 ( .A1(n37985), .A2(n36351), .ZN(n36521) );
  OAI21_X1 U19308 ( .B1(n36534), .B2(n37985), .A(n7287), .ZN(n36536) );
  NOR2_X1 U19309 ( .A1(n7290), .A2(n46514), .ZN(n46515) );
  OR2_X1 U19310 ( .A1(n45576), .A2(n7290), .ZN(n7289) );
  XNOR2_X1 U19311 ( .A(n33617), .B(n7291), .ZN(n32929) );
  NAND2_X1 U19312 ( .A1(n18330), .A2(n18059), .ZN(n7294) );
  XNOR2_X1 U19313 ( .A(n25753), .B(n25751), .ZN(n7295) );
  OAI21_X1 U19314 ( .B1(n38330), .B2(n38329), .A(n35407), .ZN(n38331) );
  OAI21_X1 U19315 ( .B1(n35390), .B2(n37673), .A(n35407), .ZN(n35414) );
  XNOR2_X1 U19318 ( .A(n33133), .B(n36951), .ZN(n34719) );
  XNOR2_X1 U19319 ( .A(n7297), .B(n34719), .ZN(n35599) );
  XNOR2_X1 U19320 ( .A(n7298), .B(n35586), .ZN(n7297) );
  INV_X1 U19321 ( .A(n34719), .ZN(n35587) );
  OAI211_X1 U19322 ( .C1(n42885), .C2(n49233), .A(n49241), .B(n42884), .ZN(
        n7302) );
  NAND3_X1 U19323 ( .A1(n49242), .A2(n49397), .A3(n49689), .ZN(n49241) );
  NAND2_X1 U19324 ( .A1(n42902), .A2(n49230), .ZN(n7300) );
  NAND2_X1 U19325 ( .A1(n7302), .A2(n588), .ZN(n7301) );
  INV_X1 U19326 ( .A(n24287), .ZN(n7303) );
  NAND2_X1 U19327 ( .A1(n7303), .A2(n24292), .ZN(n24289) );
  NAND2_X1 U19328 ( .A1(n14304), .A2(n9067), .ZN(n13599) );
  NAND2_X1 U19329 ( .A1(n7304), .A2(n13822), .ZN(n9067) );
  NAND2_X1 U19332 ( .A1(n7305), .A2(n42201), .ZN(n38924) );
  AND2_X1 U19333 ( .A1(n40806), .A2(n43323), .ZN(n38754) );
  NAND2_X1 U19334 ( .A1(n7314), .A2(n2420), .ZN(n7313) );
  NAND2_X1 U19335 ( .A1(n29411), .A2(n26905), .ZN(n7315) );
  NAND2_X1 U19336 ( .A1(n27717), .A2(n27706), .ZN(n7316) );
  XNOR2_X1 U19337 ( .A(n8482), .B(n33145), .ZN(n34883) );
  XNOR2_X1 U19338 ( .A(n7317), .B(n34883), .ZN(n7318) );
  XNOR2_X1 U19339 ( .A(n26575), .B(n7319), .ZN(n24593) );
  XNOR2_X1 U19340 ( .A(n24616), .B(n51648), .ZN(n22281) );
  INV_X1 U19341 ( .A(n47389), .ZN(n7324) );
  NAND2_X1 U19342 ( .A1(n47389), .A2(n7322), .ZN(n50956) );
  NAND2_X1 U19343 ( .A1(n50934), .A2(n7323), .ZN(n7322) );
  XNOR2_X1 U19344 ( .A(n7325), .B(n16181), .ZN(n16185) );
  XNOR2_X1 U19345 ( .A(n563), .B(n16176), .ZN(n7325) );
  NAND2_X1 U19346 ( .A1(n10923), .A2(n10922), .ZN(n7326) );
  AND2_X1 U19347 ( .A1(n7328), .A2(n10917), .ZN(n7327) );
  NAND3_X1 U19348 ( .A1(n10220), .A2(n10218), .A3(n10219), .ZN(n7328) );
  INV_X1 U19349 ( .A(n41172), .ZN(n41610) );
  XNOR2_X1 U19350 ( .A(n17726), .B(n17725), .ZN(n17840) );
  XNOR2_X1 U19351 ( .A(n17727), .B(n17840), .ZN(n7329) );
  OAI211_X1 U19352 ( .C1(n7331), .C2(n47108), .A(n45145), .B(n7330), .ZN(
        n45146) );
  NAND2_X1 U19353 ( .A1(n46881), .A2(n7332), .ZN(n7330) );
  NAND2_X1 U19354 ( .A1(n7332), .A2(n46721), .ZN(n7331) );
  NAND3_X1 U19355 ( .A1(n29321), .A2(n27890), .A3(n29323), .ZN(n27901) );
  NAND2_X1 U19356 ( .A1(n29622), .A2(n29616), .ZN(n32981) );
  NAND2_X1 U19357 ( .A1(n28157), .A2(n28879), .ZN(n7334) );
  XNOR2_X1 U19358 ( .A(n23206), .B(n7338), .ZN(n23015) );
  XNOR2_X1 U19359 ( .A(n26300), .B(n842), .ZN(n7338) );
  XNOR2_X1 U19361 ( .A(n7339), .B(n43079), .ZN(n43080) );
  XNOR2_X1 U19362 ( .A(n41464), .B(n7339), .ZN(n41465) );
  XNOR2_X1 U19363 ( .A(n42981), .B(n7339), .ZN(n42982) );
  NAND2_X1 U19364 ( .A1(n11525), .A2(n7341), .ZN(n11529) );
  XNOR2_X1 U19365 ( .A(n42964), .B(n43819), .ZN(n42965) );
  XNOR2_X2 U19366 ( .A(n41754), .B(n46137), .ZN(n43819) );
  NAND3_X1 U19367 ( .A1(n7343), .A2(n39544), .A3(n7342), .ZN(n7344) );
  NAND2_X1 U19368 ( .A1(n41932), .A2(n40251), .ZN(n7342) );
  NAND2_X1 U19369 ( .A1(n41942), .A2(n40251), .ZN(n7343) );
  NAND2_X1 U19370 ( .A1(n26309), .A2(n2528), .ZN(n26344) );
  XNOR2_X2 U19371 ( .A(Key[188]), .B(Ciphertext[97]), .ZN(n11276) );
  NAND2_X1 U19372 ( .A1(n21969), .A2(n23479), .ZN(n20992) );
  NAND2_X1 U19373 ( .A1(n50997), .A2(n11869), .ZN(n7355) );
  XNOR2_X1 U19374 ( .A(n37051), .B(n7359), .ZN(n7358) );
  XNOR2_X1 U19375 ( .A(n35247), .B(n7360), .ZN(n7359) );
  NAND2_X1 U19377 ( .A1(n29428), .A2(n7362), .ZN(n27715) );
  NAND2_X1 U19378 ( .A1(n33018), .A2(n31375), .ZN(n26635) );
  INV_X1 U19379 ( .A(n33803), .ZN(n7364) );
  XNOR2_X1 U19380 ( .A(n33729), .B(n7365), .ZN(n33803) );
  INV_X1 U19381 ( .A(n34082), .ZN(n7365) );
  XNOR2_X2 U19382 ( .A(n8204), .B(n46120), .ZN(n45415) );
  NOR2_X1 U19384 ( .A1(n29269), .A2(n8422), .ZN(n7368) );
  NOR2_X1 U19385 ( .A1(n7370), .A2(n29269), .ZN(n7369) );
  NAND3_X1 U19386 ( .A1(n14668), .A2(n14669), .A3(n14667), .ZN(n7371) );
  NAND2_X2 U19387 ( .A1(n7372), .A2(n37725), .ZN(n42154) );
  NAND2_X1 U19388 ( .A1(n48834), .A2(n48792), .ZN(n45754) );
  AND3_X2 U19389 ( .A1(n7376), .A2(n45374), .A3(n45375), .ZN(n48792) );
  AOI21_X1 U19390 ( .B1(n34683), .B2(n37548), .A(n3164), .ZN(n7378) );
  XNOR2_X1 U19391 ( .A(n18129), .B(n18123), .ZN(n7379) );
  XNOR2_X1 U19392 ( .A(n18122), .B(n7379), .ZN(n7381) );
  XNOR2_X2 U19393 ( .A(n7380), .B(n18130), .ZN(n19796) );
  INV_X1 U19394 ( .A(n32299), .ZN(n7383) );
  NAND2_X1 U19395 ( .A1(n27926), .A2(n2247), .ZN(n7382) );
  NAND3_X1 U19396 ( .A1(n21528), .A2(n20608), .A3(n20611), .ZN(n18905) );
  NAND2_X1 U19397 ( .A1(n39375), .A2(n37881), .ZN(n37033) );
  NOR2_X1 U19398 ( .A1(n10726), .A2(n10724), .ZN(n7386) );
  XNOR2_X1 U19399 ( .A(n7387), .B(n42961), .ZN(n42696) );
  XNOR2_X1 U19400 ( .A(n7387), .B(n51398), .ZN(n43118) );
  XNOR2_X1 U19401 ( .A(n45090), .B(n7387), .ZN(n45092) );
  NAND4_X1 U19403 ( .A1(n13764), .A2(n13124), .A3(n14155), .A4(n10766), .ZN(
        n10767) );
  NAND2_X1 U19404 ( .A1(n4907), .A2(n30854), .ZN(n30549) );
  OAI21_X1 U19405 ( .B1(n49719), .B2(n49721), .A(n45910), .ZN(n45911) );
  NAND3_X1 U19406 ( .A1(n7400), .A2(n36167), .A3(n38050), .ZN(n7396) );
  NAND2_X1 U19407 ( .A1(n36336), .A2(n7402), .ZN(n7401) );
  NAND2_X1 U19408 ( .A1(n36335), .A2(n36338), .ZN(n7403) );
  XNOR2_X1 U19409 ( .A(n41706), .B(n41690), .ZN(n41696) );
  NAND3_X1 U19410 ( .A1(n39000), .A2(n7407), .A3(n39001), .ZN(n7404) );
  NAND3_X1 U19411 ( .A1(n39005), .A2(n39003), .A3(n39004), .ZN(n7405) );
  NAND2_X1 U19412 ( .A1(n32823), .A2(n7408), .ZN(n31399) );
  NAND2_X1 U19413 ( .A1(n7409), .A2(n31904), .ZN(n32429) );
  XNOR2_X2 U19415 ( .A(n18825), .B(n17964), .ZN(n21389) );
  NAND2_X1 U19416 ( .A1(n29882), .A2(n742), .ZN(n7410) );
  NAND2_X1 U19417 ( .A1(n30360), .A2(n30733), .ZN(n28765) );
  NAND2_X1 U19418 ( .A1(n7412), .A2(n14342), .ZN(n7411) );
  OAI21_X1 U19419 ( .B1(n41429), .B2(n40651), .A(n7414), .ZN(n41452) );
  NAND2_X1 U19420 ( .A1(n41452), .A2(n40652), .ZN(n40645) );
  NAND2_X1 U19421 ( .A1(n10527), .A2(n10096), .ZN(n10100) );
  XNOR2_X2 U19422 ( .A(n7415), .B(Key[0]), .ZN(n10096) );
  XNOR2_X2 U19423 ( .A(n7416), .B(n33294), .ZN(n36248) );
  XNOR2_X1 U19424 ( .A(n33293), .B(n33584), .ZN(n7416) );
  NAND2_X1 U19427 ( .A1(n47937), .A2(n47989), .ZN(n47941) );
  NAND2_X1 U19429 ( .A1(n46701), .A2(n46703), .ZN(n7419) );
  INV_X1 U19431 ( .A(n21530), .ZN(n7421) );
  OAI21_X1 U19433 ( .B1(n36898), .B2(n37720), .A(n2362), .ZN(n7422) );
  NAND3_X1 U19434 ( .A1(n42149), .A2(n52092), .A3(n42136), .ZN(n41766) );
  OAI211_X1 U19435 ( .C1(n42145), .C2(n51375), .A(n687), .B(n7424), .ZN(n7423)
         );
  OR2_X1 U19436 ( .A1(n11542), .A2(n12501), .ZN(n7425) );
  NAND2_X1 U19437 ( .A1(n667), .A2(n7426), .ZN(n46971) );
  INV_X1 U19438 ( .A(n6811), .ZN(n7426) );
  NAND2_X1 U19440 ( .A1(n47144), .A2(n7426), .ZN(n46802) );
  NAND2_X1 U19441 ( .A1(n7427), .A2(n623), .ZN(n29597) );
  OR2_X2 U19444 ( .A1(n7919), .A2(n2104), .ZN(n47109) );
  NAND3_X1 U19445 ( .A1(n21527), .A2(n20188), .A3(n21525), .ZN(n20187) );
  XNOR2_X1 U19446 ( .A(n7432), .B(n34110), .ZN(n34112) );
  XNOR2_X1 U19447 ( .A(n33343), .B(n34753), .ZN(n7432) );
  INV_X1 U19448 ( .A(n7432), .ZN(n34109) );
  INV_X1 U19449 ( .A(n51708), .ZN(n12518) );
  OR2_X1 U19451 ( .A1(n51709), .A2(n12512), .ZN(n11538) );
  NOR2_X1 U19452 ( .A1(n7433), .A2(n51709), .ZN(n11540) );
  NAND2_X1 U19453 ( .A1(n9153), .A2(n12514), .ZN(n7433) );
  NAND2_X1 U19455 ( .A1(n36471), .A2(n35315), .ZN(n7437) );
  XNOR2_X2 U19456 ( .A(n7751), .B(Key[182]), .ZN(n10262) );
  NAND2_X1 U19457 ( .A1(n10261), .A2(n12356), .ZN(n9783) );
  INV_X1 U19458 ( .A(n26944), .ZN(n7438) );
  INV_X2 U19459 ( .A(n22823), .ZN(n22830) );
  NAND2_X1 U19460 ( .A1(n22823), .A2(n22506), .ZN(n22494) );
  INV_X1 U19461 ( .A(n20192), .ZN(n7440) );
  NAND2_X1 U19462 ( .A1(n50787), .A2(n7441), .ZN(n47182) );
  AOI21_X1 U19463 ( .B1(n12224), .B2(n13417), .A(n13419), .ZN(n7442) );
  NAND3_X2 U19464 ( .A1(n7443), .A2(n10600), .A3(n10599), .ZN(n14341) );
  OAI211_X1 U19465 ( .C1(n10596), .C2(n11686), .A(n7445), .B(n10595), .ZN(
        n7444) );
  XNOR2_X1 U19466 ( .A(n30810), .B(n30809), .ZN(n31358) );
  INV_X1 U19467 ( .A(n38226), .ZN(n38541) );
  INV_X1 U19468 ( .A(n38552), .ZN(n38544) );
  NAND2_X1 U19469 ( .A1(n46721), .A2(n2104), .ZN(n47095) );
  AND2_X1 U19470 ( .A1(n46565), .A2(n7449), .ZN(n8334) );
  NAND2_X1 U19471 ( .A1(n46872), .A2(n2104), .ZN(n46719) );
  OAI21_X1 U19472 ( .B1(n44578), .B2(n2104), .A(n7919), .ZN(n44576) );
  NAND2_X1 U19473 ( .A1(n22857), .A2(n22849), .ZN(n22844) );
  NAND2_X1 U19475 ( .A1(n19325), .A2(n19326), .ZN(n7450) );
  OAI211_X1 U19477 ( .C1(n7460), .C2(n7455), .A(n7454), .B(n50684), .ZN(n7458)
         );
  INV_X1 U19478 ( .A(n50690), .ZN(n7454) );
  OR2_X1 U19479 ( .A1(n50718), .A2(n50708), .ZN(n7455) );
  AOI21_X1 U19480 ( .B1(n50718), .B2(n50705), .A(n1224), .ZN(n7456) );
  NOR2_X1 U19482 ( .A1(n50710), .A2(n50723), .ZN(n7460) );
  NAND2_X1 U19483 ( .A1(n24105), .A2(n23129), .ZN(n24116) );
  XNOR2_X1 U19484 ( .A(n28372), .B(n28371), .ZN(n28373) );
  NAND2_X1 U19486 ( .A1(n13853), .A2(n13854), .ZN(n7466) );
  OAI22_X1 U19487 ( .A1(n11743), .A2(n13853), .B1(n7466), .B2(n13844), .ZN(
        n11744) );
  NAND2_X1 U19488 ( .A1(n14481), .A2(n7466), .ZN(n14886) );
  AND2_X1 U19489 ( .A1(n50530), .A2(n50529), .ZN(n7467) );
  OR2_X1 U19490 ( .A1(n50501), .A2(n50502), .ZN(n7472) );
  NAND2_X1 U19491 ( .A1(n50551), .A2(n50526), .ZN(n50494) );
  NAND3_X1 U19492 ( .A1(n27040), .A2(n2213), .A3(n26069), .ZN(n27030) );
  OAI22_X1 U19493 ( .A1(n50434), .A2(n50458), .B1(n50482), .B2(n50469), .ZN(
        n7476) );
  NAND2_X1 U19494 ( .A1(n29993), .A2(n2450), .ZN(n7477) );
  NAND2_X1 U19495 ( .A1(n29996), .A2(n31150), .ZN(n7480) );
  NAND2_X1 U19496 ( .A1(n4150), .A2(n11630), .ZN(n11462) );
  INV_X1 U19497 ( .A(n34629), .ZN(n7483) );
  NAND2_X1 U19498 ( .A1(n24157), .A2(n23821), .ZN(n23271) );
  NAND2_X1 U19499 ( .A1(n7484), .A2(n20638), .ZN(n20624) );
  OAI21_X1 U19500 ( .B1(n20623), .B2(n7484), .A(n20638), .ZN(n20198) );
  OAI21_X1 U19501 ( .B1(n21548), .B2(n21547), .A(n7484), .ZN(n21550) );
  OAI22_X1 U19503 ( .A1(n20749), .A2(n7484), .B1(n20746), .B2(n21547), .ZN(
        n18496) );
  NAND2_X1 U19505 ( .A1(n9096), .A2(n11224), .ZN(n7485) );
  NAND2_X1 U19506 ( .A1(n14641), .A2(n14644), .ZN(n13664) );
  INV_X1 U19508 ( .A(n40838), .ZN(n7488) );
  INV_X1 U19509 ( .A(n24026), .ZN(n7494) );
  NAND2_X1 U19510 ( .A1(n44578), .A2(n7495), .ZN(n47103) );
  NAND2_X1 U19511 ( .A1(n47089), .A2(n44578), .ZN(n45145) );
  NOR2_X2 U19512 ( .A1(n13780), .A2(n788), .ZN(n13178) );
  OAI211_X1 U19513 ( .C1(n41246), .C2(n41245), .A(n41685), .B(n41244), .ZN(
        n7499) );
  INV_X1 U19514 ( .A(n41244), .ZN(n40716) );
  NOR2_X1 U19515 ( .A1(n46012), .A2(n7501), .ZN(n7500) );
  NAND3_X1 U19516 ( .A1(n46007), .A2(n46010), .A3(n46011), .ZN(n7501) );
  XNOR2_X1 U19518 ( .A(n37023), .B(n34411), .ZN(n7508) );
  OR2_X1 U19519 ( .A1(n24280), .A2(n7509), .ZN(n7510) );
  NAND2_X1 U19520 ( .A1(n24289), .A2(n23513), .ZN(n7509) );
  INV_X1 U19521 ( .A(n24280), .ZN(n23506) );
  AOI22_X1 U19522 ( .A1(n31219), .A2(n31217), .B1(n7512), .B2(n31216), .ZN(
        n31228) );
  INV_X1 U19523 ( .A(n31214), .ZN(n7512) );
  NAND2_X1 U19524 ( .A1(n716), .A2(n50981), .ZN(n31214) );
  NAND2_X1 U19526 ( .A1(n13525), .A2(n51066), .ZN(n13527) );
  XNOR2_X2 U19527 ( .A(n25180), .B(n25179), .ZN(n30178) );
  XNOR2_X2 U19528 ( .A(n9173), .B(Key[68]), .ZN(n11979) );
  NAND2_X1 U19529 ( .A1(n7518), .A2(n7517), .ZN(n49123) );
  OR2_X1 U19530 ( .A1(n44772), .A2(n49126), .ZN(n7517) );
  NAND4_X2 U19532 ( .A1(n7525), .A2(n7522), .A3(n7523), .A4(n7521), .ZN(n26285) );
  NAND2_X1 U19534 ( .A1(n20983), .A2(n7527), .ZN(n7526) );
  NAND2_X1 U19535 ( .A1(n20985), .A2(n24292), .ZN(n20983) );
  AOI21_X1 U19536 ( .B1(n20990), .B2(n23478), .A(n23485), .ZN(n7528) );
  AOI22_X1 U19537 ( .A1(n7530), .A2(n12649), .B1(n12647), .B2(n2227), .ZN(
        n12656) );
  AOI21_X1 U19538 ( .B1(n9192), .B2(n7530), .A(n12659), .ZN(n9194) );
  NOR2_X1 U19539 ( .A1(n8082), .A2(n7532), .ZN(n8581) );
  AOI21_X1 U19540 ( .B1(n27961), .B2(n7532), .A(n29158), .ZN(n27962) );
  AOI21_X1 U19541 ( .B1(n29149), .B2(n29147), .A(n7531), .ZN(n27955) );
  NAND2_X1 U19542 ( .A1(n8582), .A2(n7532), .ZN(n8580) );
  NAND3_X2 U19543 ( .A1(n16795), .A2(n16794), .A3(n16796), .ZN(n21975) );
  OAI21_X1 U19544 ( .B1(n21991), .B2(n21975), .A(n7533), .ZN(n16854) );
  NAND2_X1 U19545 ( .A1(n21991), .A2(n7534), .ZN(n7533) );
  NAND2_X1 U19546 ( .A1(n23489), .A2(n7535), .ZN(n7534) );
  OAI21_X1 U19547 ( .B1(n9184), .B2(n9185), .A(n9183), .ZN(n7536) );
  NAND2_X1 U19548 ( .A1(n7539), .A2(n7537), .ZN(n13886) );
  NAND2_X1 U19549 ( .A1(n7538), .A2(n9196), .ZN(n7537) );
  NAND3_X1 U19550 ( .A1(n7541), .A2(n9196), .A3(n7540), .ZN(n7539) );
  NAND3_X1 U19551 ( .A1(n13886), .A2(n14870), .A3(n50966), .ZN(n15422) );
  NAND3_X1 U19552 ( .A1(n33014), .A2(n7542), .A3(n33013), .ZN(n33015) );
  AND2_X1 U19553 ( .A1(n31383), .A2(n33002), .ZN(n33019) );
  AOI21_X1 U19554 ( .B1(n49905), .B2(n49923), .A(n49878), .ZN(n49880) );
  NAND2_X1 U19555 ( .A1(n20727), .A2(n20721), .ZN(n7545) );
  NAND2_X1 U19556 ( .A1(n23563), .A2(n23547), .ZN(n20727) );
  XNOR2_X1 U19557 ( .A(n16623), .B(n17327), .ZN(n19112) );
  INV_X1 U19558 ( .A(n38593), .ZN(n38166) );
  XNOR2_X2 U19559 ( .A(n35665), .B(n35664), .ZN(n38593) );
  NAND2_X1 U19562 ( .A1(n720), .A2(n31383), .ZN(n30543) );
  NAND3_X1 U19563 ( .A1(n29148), .A2(n29174), .A3(n29152), .ZN(n7548) );
  NAND2_X1 U19564 ( .A1(n7549), .A2(n49923), .ZN(n49924) );
  XNOR2_X1 U19565 ( .A(n376), .B(n7550), .ZN(n26717) );
  XNOR2_X1 U19566 ( .A(n35829), .B(n7550), .ZN(n33820) );
  XNOR2_X1 U19567 ( .A(n37046), .B(n7550), .ZN(n37048) );
  XNOR2_X1 U19568 ( .A(n32742), .B(n7550), .ZN(n35033) );
  NAND3_X1 U19569 ( .A1(n38949), .A2(n39410), .A3(n39208), .ZN(n38947) );
  XNOR2_X1 U19570 ( .A(n7553), .B(n7552), .ZN(n7551) );
  XNOR2_X1 U19571 ( .A(n26520), .B(n24982), .ZN(n7552) );
  NAND2_X1 U19572 ( .A1(n11896), .A2(n11895), .ZN(n7554) );
  INV_X1 U19573 ( .A(n14769), .ZN(n15240) );
  INV_X2 U19574 ( .A(n41540), .ZN(n41554) );
  NAND2_X1 U19575 ( .A1(n41544), .A2(n41540), .ZN(n40981) );
  XNOR2_X1 U19577 ( .A(n32935), .B(n7556), .ZN(n35065) );
  XNOR2_X1 U19578 ( .A(n7556), .B(n35237), .ZN(n33382) );
  XNOR2_X1 U19579 ( .A(n7556), .B(n33988), .ZN(n33990) );
  XNOR2_X1 U19580 ( .A(n7556), .B(n36970), .ZN(n36973) );
  XNOR2_X1 U19581 ( .A(n25953), .B(n445), .ZN(n25955) );
  XNOR2_X1 U19582 ( .A(n28276), .B(n445), .ZN(n25461) );
  XNOR2_X1 U19583 ( .A(n444), .B(n26555), .ZN(n26558) );
  XNOR2_X1 U19584 ( .A(n24435), .B(n444), .ZN(n24440) );
  XNOR2_X1 U19585 ( .A(n26142), .B(n444), .ZN(n28280) );
  NAND2_X1 U19586 ( .A1(n29319), .A2(n52216), .ZN(n27890) );
  XNOR2_X1 U19588 ( .A(n25964), .B(n25963), .ZN(n7560) );
  NAND4_X1 U19589 ( .A1(n13823), .A2(n13824), .A3(n14318), .A4(n13822), .ZN(
        n13830) );
  AND2_X1 U19590 ( .A1(n10296), .A2(n10302), .ZN(n10293) );
  XNOR2_X2 U19591 ( .A(n7563), .B(Key[149]), .ZN(n10302) );
  NAND3_X1 U19592 ( .A1(n7725), .A2(n50288), .A3(n7567), .ZN(n7566) );
  NAND2_X1 U19593 ( .A1(n7724), .A2(n46037), .ZN(n7569) );
  NAND2_X1 U19594 ( .A1(n41374), .A2(n38885), .ZN(n40240) );
  XNOR2_X1 U19595 ( .A(n33101), .B(n37091), .ZN(n32338) );
  NAND4_X2 U19596 ( .A1(n30865), .A2(n30864), .A3(n30862), .A4(n30863), .ZN(
        n35632) );
  INV_X2 U19597 ( .A(n14929), .ZN(n15766) );
  NAND2_X1 U19598 ( .A1(n1672), .A2(n31624), .ZN(n31583) );
  NAND2_X1 U19599 ( .A1(n28663), .A2(n28664), .ZN(n7573) );
  NAND2_X1 U19600 ( .A1(n7576), .A2(n49695), .ZN(n7577) );
  INV_X1 U19601 ( .A(n42886), .ZN(n7576) );
  NAND2_X1 U19602 ( .A1(n18378), .A2(n20035), .ZN(n7581) );
  NAND2_X1 U19603 ( .A1(n7583), .A2(n771), .ZN(n7582) );
  NAND2_X1 U19604 ( .A1(n18383), .A2(n18382), .ZN(n7583) );
  NAND2_X1 U19606 ( .A1(n18375), .A2(n7585), .ZN(n7584) );
  NAND2_X1 U19607 ( .A1(n11000), .A2(n7588), .ZN(n7587) );
  NAND2_X1 U19610 ( .A1(n12884), .A2(n7591), .ZN(n12885) );
  XNOR2_X1 U19611 ( .A(n51362), .B(n41743), .ZN(n41744) );
  XNOR2_X1 U19612 ( .A(n51362), .B(n43363), .ZN(n43364) );
  XNOR2_X1 U19613 ( .A(n52085), .B(n51362), .ZN(n42533) );
  XNOR2_X1 U19614 ( .A(n43048), .B(n51362), .ZN(n45368) );
  NAND2_X1 U19615 ( .A1(n7593), .A2(n23157), .ZN(n23159) );
  INV_X1 U19616 ( .A(n36586), .ZN(n35881) );
  OAI21_X1 U19617 ( .B1(n24776), .B2(n3765), .A(n2642), .ZN(n26939) );
  NOR2_X1 U19618 ( .A1(n27067), .A2(n24776), .ZN(n27659) );
  NAND2_X1 U19619 ( .A1(n27660), .A2(n24776), .ZN(n26878) );
  OAI21_X1 U19620 ( .B1(n7597), .B2(n7596), .A(n36459), .ZN(n7595) );
  NAND2_X1 U19621 ( .A1(n34410), .A2(n36044), .ZN(n7596) );
  NAND2_X1 U19622 ( .A1(n36584), .A2(n35878), .ZN(n7597) );
  NAND2_X1 U19623 ( .A1(n7598), .A2(n31684), .ZN(n30014) );
  NAND2_X1 U19624 ( .A1(n49081), .A2(n49070), .ZN(n7600) );
  NAND3_X1 U19625 ( .A1(n49081), .A2(n49070), .A3(n2460), .ZN(n7599) );
  AOI21_X1 U19626 ( .B1(n44799), .B2(n49107), .A(n7600), .ZN(n44806) );
  NAND2_X1 U19628 ( .A1(n2484), .A2(n7602), .ZN(n7601) );
  NAND2_X1 U19630 ( .A1(n28551), .A2(n26501), .ZN(n7605) );
  AND2_X1 U19631 ( .A1(n7606), .A2(n48893), .ZN(n45704) );
  INV_X1 U19633 ( .A(n46349), .ZN(n46269) );
  NAND2_X1 U19634 ( .A1(n45238), .A2(n46356), .ZN(n46349) );
  NOR2_X1 U19635 ( .A1(n45690), .A2(n7615), .ZN(n45691) );
  OAI21_X1 U19636 ( .B1(n46266), .B2(n46349), .A(n45689), .ZN(n7615) );
  INV_X1 U19637 ( .A(n38704), .ZN(n39225) );
  AND2_X1 U19638 ( .A1(n6172), .A2(n52143), .ZN(n46008) );
  NAND2_X1 U19640 ( .A1(n50010), .A2(n52143), .ZN(n49995) );
  OAI22_X1 U19641 ( .A1(n50318), .A2(n52224), .B1(n50316), .B2(n7616), .ZN(
        n50319) );
  NAND2_X1 U19642 ( .A1(n46006), .A2(n52143), .ZN(n46007) );
  OAI21_X1 U19643 ( .B1(n31931), .B2(n31934), .A(n31347), .ZN(n29607) );
  XNOR2_X1 U19644 ( .A(n36851), .B(n36679), .ZN(n7620) );
  NAND2_X1 U19645 ( .A1(n11809), .A2(n7621), .ZN(n11810) );
  INV_X1 U19646 ( .A(n12977), .ZN(n7621) );
  NAND4_X2 U19647 ( .A1(n31478), .A2(n31479), .A3(n31480), .A4(n31477), .ZN(
        n7624) );
  XNOR2_X1 U19648 ( .A(n7624), .B(n33838), .ZN(n33839) );
  XNOR2_X1 U19649 ( .A(n37066), .B(n7624), .ZN(n33194) );
  XNOR2_X1 U19650 ( .A(n7624), .B(n35523), .ZN(n35524) );
  XNOR2_X1 U19651 ( .A(n34013), .B(n7624), .ZN(n34019) );
  NAND2_X1 U19654 ( .A1(n19837), .A2(n19834), .ZN(n19831) );
  NAND2_X1 U19655 ( .A1(n7630), .A2(n7629), .ZN(n40489) );
  NAND2_X1 U19656 ( .A1(n40488), .A2(n41110), .ZN(n7629) );
  NAND2_X1 U19658 ( .A1(n41256), .A2(n41112), .ZN(n40486) );
  INV_X1 U19661 ( .A(n37735), .ZN(n39005) );
  NAND2_X1 U19662 ( .A1(n7634), .A2(n39003), .ZN(n36917) );
  NAND3_X1 U19663 ( .A1(n7634), .A2(n39004), .A3(n7632), .ZN(n7635) );
  NOR2_X1 U19664 ( .A1(n37735), .A2(n39400), .ZN(n7632) );
  NAND4_X2 U19665 ( .A1(n7635), .A2(n36925), .A3(n36924), .A4(n36923), .ZN(
        n41735) );
  NAND2_X1 U19666 ( .A1(n7639), .A2(n49987), .ZN(n46014) );
  XNOR2_X1 U19667 ( .A(n16250), .B(n7643), .ZN(n7642) );
  NAND2_X1 U19668 ( .A1(n34907), .A2(n37890), .ZN(n7644) );
  NAND2_X1 U19669 ( .A1(n30721), .A2(n29851), .ZN(n29848) );
  AND2_X1 U19670 ( .A1(n42086), .A2(n42092), .ZN(n7647) );
  INV_X1 U19673 ( .A(n23425), .ZN(n22313) );
  NAND2_X1 U19674 ( .A1(n23425), .A2(n23412), .ZN(n7651) );
  AOI21_X1 U19675 ( .B1(n20156), .B2(n20158), .A(n20155), .ZN(n7653) );
  OAI21_X1 U19676 ( .B1(n20156), .B2(n4081), .A(n7652), .ZN(n20111) );
  INV_X1 U19677 ( .A(n25740), .ZN(n24965) );
  NAND2_X1 U19678 ( .A1(n15031), .A2(n13806), .ZN(n13807) );
  NAND2_X1 U19679 ( .A1(n13797), .A2(n69), .ZN(n13806) );
  NAND2_X1 U19680 ( .A1(n27609), .A2(n23861), .ZN(n30673) );
  NAND2_X1 U19681 ( .A1(n11974), .A2(n10451), .ZN(n10345) );
  INV_X1 U19683 ( .A(n46288), .ZN(n7657) );
  NAND2_X1 U19684 ( .A1(n49147), .A2(n7656), .ZN(n46289) );
  NAND2_X1 U19685 ( .A1(n7657), .A2(n49137), .ZN(n49147) );
  INV_X1 U19686 ( .A(n29591), .ZN(n7659) );
  INV_X1 U19687 ( .A(n31110), .ZN(n29584) );
  NAND4_X4 U19688 ( .A1(n38351), .A2(n38349), .A3(n38348), .A4(n38350), .ZN(
        n40862) );
  XNOR2_X1 U19690 ( .A(n8736), .B(n25144), .ZN(n7664) );
  OAI211_X1 U19691 ( .C1(n47255), .C2(n7671), .A(n7669), .B(n7668), .ZN(
        Plaintext[63]) );
  NAND2_X1 U19692 ( .A1(n47255), .A2(n34420), .ZN(n7668) );
  INV_X1 U19693 ( .A(n7675), .ZN(n7670) );
  NAND2_X1 U19694 ( .A1(n7673), .A2(n7672), .ZN(n7671) );
  NAND2_X1 U19695 ( .A1(n48698), .A2(n7676), .ZN(n7672) );
  NAND2_X1 U19696 ( .A1(n47246), .A2(n655), .ZN(n7675) );
  NAND2_X1 U19697 ( .A1(n47245), .A2(n47404), .ZN(n7676) );
  NAND2_X1 U19698 ( .A1(n21885), .A2(n22861), .ZN(n19609) );
  NAND2_X1 U19699 ( .A1(n30982), .A2(n30983), .ZN(n30974) );
  NAND2_X1 U19700 ( .A1(n29279), .A2(n27924), .ZN(n7683) );
  NAND2_X1 U19701 ( .A1(n34090), .A2(n36027), .ZN(n37956) );
  INV_X1 U19702 ( .A(n50344), .ZN(n7684) );
  XNOR2_X2 U19703 ( .A(n43877), .B(n44361), .ZN(n50344) );
  NAND2_X1 U19704 ( .A1(n39714), .A2(n7685), .ZN(n39715) );
  NAND2_X1 U19705 ( .A1(n41084), .A2(n39709), .ZN(n34668) );
  XNOR2_X1 U19706 ( .A(n19208), .B(n19209), .ZN(n7686) );
  AND2_X1 U19707 ( .A1(n8856), .A2(n8857), .ZN(n7687) );
  INV_X1 U19708 ( .A(n13590), .ZN(n7688) );
  XNOR2_X1 U19709 ( .A(n26294), .B(n8596), .ZN(n24675) );
  NAND3_X1 U19710 ( .A1(n19455), .A2(n21269), .A3(n19774), .ZN(n19453) );
  OR2_X1 U19711 ( .A1(n2182), .A2(n19016), .ZN(n19774) );
  NAND2_X1 U19712 ( .A1(n23442), .A2(n7689), .ZN(n22585) );
  AND4_X2 U19713 ( .A1(n7690), .A2(n28794), .A3(n28795), .A4(n7691), .ZN(
        n32633) );
  INV_X1 U19715 ( .A(n7694), .ZN(n10830) );
  OR2_X1 U19716 ( .A1(n7694), .A2(n51709), .ZN(n11256) );
  NAND2_X1 U19717 ( .A1(n11263), .A2(n7693), .ZN(n11264) );
  XNOR2_X1 U19718 ( .A(n42269), .B(n42268), .ZN(n42872) );
  INV_X1 U19719 ( .A(n43365), .ZN(n7695) );
  XNOR2_X1 U19720 ( .A(n7695), .B(n42872), .ZN(n7696) );
  OAI21_X1 U19721 ( .B1(n45844), .B2(n46915), .A(n7700), .ZN(n7698) );
  NAND3_X1 U19722 ( .A1(n46694), .A2(n46607), .A3(n46692), .ZN(n7699) );
  AND2_X1 U19723 ( .A1(n31577), .A2(n30853), .ZN(n7705) );
  INV_X1 U19724 ( .A(n38543), .ZN(n38558) );
  INV_X1 U19725 ( .A(n38221), .ZN(n38217) );
  NAND2_X1 U19726 ( .A1(n3817), .A2(n6538), .ZN(n38221) );
  OAI21_X1 U19727 ( .B1(n24280), .B2(n24279), .A(n7706), .ZN(n24281) );
  NOR2_X1 U19728 ( .A1(n24283), .A2(n7707), .ZN(n24277) );
  XNOR2_X2 U19729 ( .A(n7708), .B(Key[144]), .ZN(n12285) );
  NAND2_X1 U19732 ( .A1(n13530), .A2(n12767), .ZN(n7717) );
  XNOR2_X1 U19735 ( .A(n25350), .B(n25349), .ZN(n27093) );
  INV_X1 U19736 ( .A(n30210), .ZN(n30207) );
  XNOR2_X2 U19737 ( .A(n8960), .B(Key[119]), .ZN(n12705) );
  XNOR2_X2 U19738 ( .A(n37056), .B(n37057), .ZN(n37924) );
  NAND2_X1 U19739 ( .A1(n30484), .A2(n7723), .ZN(n32379) );
  INV_X1 U19740 ( .A(n47307), .ZN(n7724) );
  NAND2_X1 U19741 ( .A1(n49641), .A2(n50287), .ZN(n7725) );
  NAND3_X1 U19742 ( .A1(n9297), .A2(n10609), .A3(n10618), .ZN(n7726) );
  NAND2_X1 U19743 ( .A1(n9914), .A2(n10618), .ZN(n7727) );
  NAND3_X1 U19744 ( .A1(n41345), .A2(n41349), .A3(n40358), .ZN(n40738) );
  XNOR2_X1 U19746 ( .A(n26254), .B(n24926), .ZN(n25491) );
  NAND2_X1 U19747 ( .A1(n13526), .A2(n11841), .ZN(n13513) );
  INV_X1 U19748 ( .A(n8002), .ZN(n13497) );
  NAND2_X1 U19749 ( .A1(n39169), .A2(n38667), .ZN(n39183) );
  INV_X1 U19750 ( .A(n419), .ZN(n37158) );
  NAND2_X1 U19751 ( .A1(n34428), .A2(n36051), .ZN(n7730) );
  NAND2_X1 U19752 ( .A1(n24067), .A2(n23736), .ZN(n7731) );
  INV_X1 U19753 ( .A(n36454), .ZN(n36047) );
  NAND3_X1 U19754 ( .A1(n14489), .A2(n7735), .A3(n787), .ZN(n13925) );
  OAI211_X1 U19755 ( .C1(n15362), .C2(n7735), .A(n14823), .B(n14822), .ZN(
        n14824) );
  OR2_X1 U19756 ( .A1(n14817), .A2(n7735), .ZN(n7734) );
  NAND2_X1 U19758 ( .A1(n31426), .A2(n31428), .ZN(n7736) );
  NAND2_X1 U19759 ( .A1(n50728), .A2(n50723), .ZN(n7746) );
  OAI211_X1 U19760 ( .C1(n7742), .C2(n7740), .A(n7738), .B(n7737), .ZN(
        Plaintext[173]) );
  OAI21_X1 U19761 ( .B1(n7739), .B2(n50737), .A(n7747), .ZN(n7738) );
  NAND2_X1 U19762 ( .A1(n7746), .A2(n7741), .ZN(n7740) );
  INV_X1 U19763 ( .A(n50737), .ZN(n7741) );
  NAND2_X1 U19764 ( .A1(n50725), .A2(n50724), .ZN(n7745) );
  XNOR2_X1 U19765 ( .A(n16953), .B(n16412), .ZN(n17768) );
  XNOR2_X1 U19766 ( .A(n17768), .B(n13268), .ZN(n13572) );
  NAND3_X1 U19767 ( .A1(n7756), .A2(n12950), .A3(n7754), .ZN(n11321) );
  NAND2_X1 U19768 ( .A1(n14673), .A2(n7757), .ZN(n13627) );
  OAI21_X1 U19769 ( .B1(n35150), .B2(n7760), .A(n7758), .ZN(n36104) );
  NAND2_X1 U19770 ( .A1(n38562), .A2(n7759), .ZN(n7758) );
  NAND2_X1 U19771 ( .A1(n38572), .A2(n36098), .ZN(n7760) );
  NAND2_X1 U19772 ( .A1(n43180), .A2(n49990), .ZN(n47356) );
  NAND2_X1 U19773 ( .A1(n40034), .A2(n40185), .ZN(n7763) );
  NAND2_X1 U19774 ( .A1(n7765), .A2(n48162), .ZN(n7764) );
  NAND2_X1 U19775 ( .A1(n48151), .A2(n48154), .ZN(n7765) );
  INV_X1 U19776 ( .A(n48103), .ZN(n48151) );
  NAND4_X2 U19777 ( .A1(n7769), .A2(n7770), .A3(n7768), .A4(n11807), .ZN(
        n16435) );
  NAND2_X1 U19778 ( .A1(n11802), .A2(n11801), .ZN(n7768) );
  NAND2_X1 U19779 ( .A1(n11803), .A2(n13487), .ZN(n7770) );
  INV_X1 U19780 ( .A(n7771), .ZN(n34051) );
  XNOR2_X2 U19781 ( .A(n34841), .B(n8135), .ZN(n7771) );
  XNOR2_X1 U19782 ( .A(n34572), .B(n7771), .ZN(n36796) );
  XNOR2_X1 U19783 ( .A(n515), .B(n7771), .ZN(n33860) );
  XNOR2_X1 U19784 ( .A(n33724), .B(n7771), .ZN(n33725) );
  XNOR2_X1 U19785 ( .A(n36986), .B(n7771), .ZN(n36987) );
  XNOR2_X1 U19786 ( .A(n34574), .B(n7771), .ZN(n35549) );
  NAND4_X2 U19787 ( .A1(n7773), .A2(n23618), .A3(n51789), .A4(n23619), .ZN(
        n27309) );
  NAND2_X1 U19788 ( .A1(n389), .A2(n2178), .ZN(n47161) );
  NOR2_X1 U19789 ( .A1(n663), .A2(n2178), .ZN(n46889) );
  NAND2_X1 U19790 ( .A1(n47155), .A2(n7776), .ZN(n47157) );
  OR2_X1 U19791 ( .A1(n47159), .A2(n2178), .ZN(n7776) );
  OAI21_X1 U19792 ( .B1(n44470), .B2(n2178), .A(n47149), .ZN(n44475) );
  OAI21_X1 U19793 ( .B1(n38406), .B2(n39674), .A(n7779), .ZN(n7778) );
  NAND3_X1 U19795 ( .A1(n12441), .A2(n12440), .A3(n12709), .ZN(n12689) );
  XNOR2_X1 U19796 ( .A(n16720), .B(n16952), .ZN(n16721) );
  NAND2_X1 U19797 ( .A1(n27669), .A2(n26747), .ZN(n7783) );
  XNOR2_X1 U19798 ( .A(n35085), .B(n7787), .ZN(n34041) );
  XNOR2_X1 U19799 ( .A(n7787), .B(n35532), .ZN(n35533) );
  XNOR2_X1 U19800 ( .A(n35536), .B(n7787), .ZN(n32996) );
  XNOR2_X1 U19801 ( .A(n7787), .B(n35644), .ZN(n35646) );
  NAND4_X2 U19802 ( .A1(n29570), .A2(n7788), .A3(n29572), .A4(n29571), .ZN(
        n31512) );
  NAND2_X1 U19803 ( .A1(n7791), .A2(n7790), .ZN(n7789) );
  NAND2_X1 U19804 ( .A1(n51676), .A2(n21155), .ZN(n7790) );
  NAND2_X1 U19805 ( .A1(n23547), .A2(n23568), .ZN(n7791) );
  OR2_X2 U19806 ( .A1(n7792), .A2(n8035), .ZN(n23068) );
  NAND2_X1 U19807 ( .A1(n15770), .A2(n14929), .ZN(n15304) );
  NOR2_X1 U19808 ( .A1(n42988), .A2(n7793), .ZN(n7795) );
  NAND2_X1 U19809 ( .A1(n31447), .A2(n31455), .ZN(n31540) );
  XNOR2_X1 U19810 ( .A(n7799), .B(n26155), .ZN(n23721) );
  XNOR2_X1 U19811 ( .A(n7800), .B(n7801), .ZN(n7799) );
  XNOR2_X1 U19812 ( .A(n23718), .B(n23717), .ZN(n7800) );
  INV_X1 U19813 ( .A(n14983), .ZN(n15119) );
  OAI21_X1 U19814 ( .B1(n14246), .B2(n14984), .A(n7803), .ZN(n14243) );
  NAND3_X1 U19815 ( .A1(n14980), .A2(n15117), .A3(n14247), .ZN(n7803) );
  NAND2_X1 U19816 ( .A1(n30677), .A2(n30676), .ZN(n7804) );
  INV_X1 U19817 ( .A(n24687), .ZN(n26864) );
  INV_X1 U19818 ( .A(n30677), .ZN(n27599) );
  NAND2_X1 U19819 ( .A1(n24687), .A2(n26909), .ZN(n30677) );
  INV_X1 U19820 ( .A(n30664), .ZN(n7805) );
  AND2_X1 U19821 ( .A1(n51434), .A2(n21185), .ZN(n19529) );
  INV_X1 U19822 ( .A(n23094), .ZN(n7806) );
  INV_X1 U19823 ( .A(n7808), .ZN(n23097) );
  NAND2_X1 U19824 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  OAI21_X1 U19825 ( .B1(n23099), .B2(n23098), .A(n7808), .ZN(n23295) );
  OAI21_X1 U19826 ( .B1(n14018), .B2(n14036), .A(n13737), .ZN(n11047) );
  NAND2_X1 U19827 ( .A1(n41999), .A2(n42000), .ZN(n42005) );
  INV_X1 U19828 ( .A(n37790), .ZN(n39375) );
  OAI21_X1 U19829 ( .B1(n7812), .B2(n11466), .A(n11635), .ZN(n9102) );
  OAI21_X1 U19830 ( .B1(n11628), .B2(n7812), .A(n10852), .ZN(n9327) );
  XNOR2_X1 U19831 ( .A(n7813), .B(n15850), .ZN(n15871) );
  XNOR2_X1 U19832 ( .A(n19210), .B(n16732), .ZN(n7813) );
  INV_X1 U19833 ( .A(n7815), .ZN(n7814) );
  NAND3_X1 U19834 ( .A1(n7814), .A2(n51737), .A3(n39035), .ZN(n36255) );
  NAND3_X1 U19835 ( .A1(n29340), .A2(n29339), .A3(n2537), .ZN(n7816) );
  XNOR2_X1 U19836 ( .A(n27425), .B(n52170), .ZN(n27426) );
  XNOR2_X1 U19837 ( .A(n25805), .B(n7819), .ZN(n27218) );
  XNOR2_X1 U19838 ( .A(n28246), .B(n52170), .ZN(n26010) );
  XNOR2_X1 U19839 ( .A(n25137), .B(n52170), .ZN(n25138) );
  XNOR2_X1 U19840 ( .A(n25934), .B(n7819), .ZN(n8178) );
  NAND3_X1 U19841 ( .A1(n23625), .A2(n23638), .A3(n7820), .ZN(n23091) );
  NOR2_X1 U19842 ( .A1(n7823), .A2(n12286), .ZN(n10225) );
  NAND3_X1 U19843 ( .A1(n7823), .A2(n12276), .A3(n12294), .ZN(n12281) );
  NOR2_X1 U19844 ( .A1(n10715), .A2(n7823), .ZN(n9003) );
  NAND2_X1 U19845 ( .A1(n7822), .A2(n7821), .ZN(n8606) );
  NAND2_X1 U19846 ( .A1(n12292), .A2(n7823), .ZN(n7821) );
  NAND2_X1 U19847 ( .A1(n12293), .A2(n7823), .ZN(n12295) );
  NAND3_X1 U19848 ( .A1(n50275), .A2(n50276), .A3(n7824), .ZN(n50285) );
  NAND2_X1 U19849 ( .A1(n29438), .A2(n29447), .ZN(n7826) );
  INV_X1 U19851 ( .A(n18357), .ZN(n18346) );
  XNOR2_X1 U19852 ( .A(n7828), .B(n34078), .ZN(n35120) );
  NAND4_X2 U19853 ( .A1(n31757), .A2(n7829), .A3(n31756), .A4(n31758), .ZN(
        n37304) );
  OAI21_X1 U19856 ( .B1(n36562), .B2(n36489), .A(n34640), .ZN(n7837) );
  OAI21_X1 U19857 ( .B1(n35314), .B2(n7837), .A(n36015), .ZN(n34645) );
  NAND3_X1 U19858 ( .A1(n36492), .A2(n36473), .A3(n4246), .ZN(n36489) );
  NOR2_X1 U19859 ( .A1(n36576), .A2(n2086), .ZN(n35314) );
  NAND2_X1 U19860 ( .A1(n18352), .A2(n18346), .ZN(n19065) );
  NAND2_X1 U19862 ( .A1(n46286), .A2(n7840), .ZN(n43402) );
  NAND2_X1 U19863 ( .A1(n7841), .A2(n44730), .ZN(n7840) );
  NAND2_X1 U19864 ( .A1(n43401), .A2(n7842), .ZN(n7841) );
  NAND2_X1 U19865 ( .A1(n10218), .A2(n10137), .ZN(n10935) );
  NAND2_X1 U19866 ( .A1(n18346), .A2(n7844), .ZN(n7843) );
  INV_X1 U19867 ( .A(n20144), .ZN(n7845) );
  NAND2_X1 U19868 ( .A1(n23211), .A2(n8732), .ZN(n7846) );
  INV_X1 U19869 ( .A(n40572), .ZN(n7848) );
  XNOR2_X1 U19870 ( .A(n43106), .B(n43105), .ZN(n7849) );
  XNOR2_X1 U19871 ( .A(n18669), .B(n2407), .ZN(n16505) );
  NAND2_X1 U19872 ( .A1(n13119), .A2(n13118), .ZN(n7853) );
  OR2_X1 U19873 ( .A1(n38493), .A2(n5364), .ZN(n37526) );
  NAND2_X1 U19874 ( .A1(n7856), .A2(n7855), .ZN(n7854) );
  NAND2_X1 U19875 ( .A1(n20208), .A2(n20207), .ZN(n7855) );
  INV_X1 U19876 ( .A(n40591), .ZN(n40059) );
  XNOR2_X1 U19877 ( .A(n15666), .B(n7863), .ZN(n7862) );
  XNOR2_X2 U19878 ( .A(n7862), .B(n51407), .ZN(n20211) );
  NAND2_X1 U19880 ( .A1(n7868), .A2(n435), .ZN(n32294) );
  INV_X1 U19881 ( .A(n31749), .ZN(n7868) );
  INV_X1 U19882 ( .A(n32294), .ZN(n31843) );
  AOI21_X1 U19883 ( .B1(n38484), .B2(n38478), .A(n37416), .ZN(n38126) );
  NAND2_X1 U19884 ( .A1(n38484), .A2(n38478), .ZN(n37425) );
  NAND2_X1 U19885 ( .A1(n36120), .A2(n38483), .ZN(n7869) );
  INV_X1 U19886 ( .A(n9335), .ZN(n11272) );
  INV_X1 U19887 ( .A(n37591), .ZN(n35458) );
  XNOR2_X2 U19888 ( .A(n33743), .B(n8336), .ZN(n37591) );
  XNOR2_X1 U19890 ( .A(n44039), .B(n44038), .ZN(n7872) );
  NAND2_X1 U19891 ( .A1(n28487), .A2(n31886), .ZN(n30118) );
  NAND2_X1 U19892 ( .A1(n7875), .A2(n7874), .ZN(n7873) );
  INV_X1 U19893 ( .A(n10244), .ZN(n9031) );
  NAND2_X1 U19894 ( .A1(n10244), .A2(n10195), .ZN(n9753) );
  XNOR2_X1 U19895 ( .A(n395), .B(n28423), .ZN(n26049) );
  XNOR2_X1 U19896 ( .A(n395), .B(n749), .ZN(n24721) );
  XNOR2_X1 U19897 ( .A(n27447), .B(n396), .ZN(n23843) );
  XNOR2_X1 U19898 ( .A(n395), .B(n24732), .ZN(n24637) );
  XNOR2_X1 U19899 ( .A(n25737), .B(n396), .ZN(n8335) );
  XNOR2_X1 U19900 ( .A(n27445), .B(n396), .ZN(n23369) );
  XNOR2_X1 U19901 ( .A(n8621), .B(n396), .ZN(n26513) );
  XNOR2_X1 U19902 ( .A(n25423), .B(n396), .ZN(n27463) );
  XNOR2_X1 U19903 ( .A(n24966), .B(n396), .ZN(n26216) );
  AND2_X1 U19905 ( .A1(n13977), .A2(n13982), .ZN(n7878) );
  NAND2_X1 U19906 ( .A1(n31882), .A2(n31879), .ZN(n31877) );
  INV_X1 U19908 ( .A(n50329), .ZN(n7883) );
  NAND2_X1 U19909 ( .A1(n46968), .A2(n50329), .ZN(n7881) );
  OR2_X1 U19910 ( .A1(n14099), .A2(n51383), .ZN(n7886) );
  INV_X1 U19911 ( .A(n28137), .ZN(n7888) );
  XNOR2_X1 U19912 ( .A(n42453), .B(n44300), .ZN(n41630) );
  NOR2_X2 U19913 ( .A1(n7889), .A2(n40721), .ZN(n44904) );
  INV_X1 U19915 ( .A(n12087), .ZN(n12093) );
  NAND2_X1 U19916 ( .A1(n12380), .A2(n11352), .ZN(n12385) );
  NAND2_X1 U19917 ( .A1(n12085), .A2(n11353), .ZN(n7894) );
  NAND2_X1 U19918 ( .A1(n8643), .A2(n12087), .ZN(n12101) );
  NAND2_X1 U19919 ( .A1(n27885), .A2(n30208), .ZN(n7896) );
  NAND2_X1 U19920 ( .A1(n38982), .A2(n38983), .ZN(n38984) );
  NAND2_X1 U19921 ( .A1(n39483), .A2(n7159), .ZN(n38983) );
  NOR2_X1 U19922 ( .A1(n7901), .A2(n28504), .ZN(n28514) );
  OAI21_X1 U19923 ( .B1(n7901), .B2(n28958), .A(n28957), .ZN(n28959) );
  NAND2_X1 U19924 ( .A1(n28503), .A2(n7902), .ZN(n7901) );
  NAND2_X1 U19925 ( .A1(n38004), .A2(n2377), .ZN(n7903) );
  OAI21_X1 U19926 ( .B1(n10221), .B2(n10218), .A(n7904), .ZN(n10139) );
  XNOR2_X2 U19927 ( .A(n8899), .B(Key[161]), .ZN(n11884) );
  NAND4_X2 U19928 ( .A1(n11506), .A2(n11504), .A3(n11507), .A4(n11505), .ZN(
        n15384) );
  NAND2_X1 U19929 ( .A1(n7906), .A2(n15384), .ZN(n15367) );
  INV_X1 U19930 ( .A(n15358), .ZN(n15365) );
  NAND2_X1 U19931 ( .A1(n22978), .A2(n22977), .ZN(n23002) );
  INV_X2 U19933 ( .A(n37774), .ZN(n37782) );
  OR2_X1 U19934 ( .A1(n2120), .A2(n38275), .ZN(n7914) );
  NAND2_X1 U19935 ( .A1(n38291), .A2(n37623), .ZN(n7915) );
  NAND3_X1 U19936 ( .A1(n7917), .A2(n36631), .A3(n36630), .ZN(n36637) );
  NAND2_X1 U19937 ( .A1(n36640), .A2(n38071), .ZN(n7917) );
  INV_X1 U19939 ( .A(n7922), .ZN(n40141) );
  NAND2_X1 U19940 ( .A1(n40815), .A2(n40835), .ZN(n7922) );
  NAND3_X1 U19941 ( .A1(n37710), .A2(n39691), .A3(n7921), .ZN(n37715) );
  NAND2_X1 U19942 ( .A1(n7922), .A2(n40828), .ZN(n7921) );
  NAND2_X1 U19943 ( .A1(n27775), .A2(n31088), .ZN(n30605) );
  AND2_X2 U19944 ( .A1(n7924), .A2(n7923), .ZN(n24283) );
  NAND2_X1 U19945 ( .A1(n7950), .A2(n18873), .ZN(n7924) );
  OR2_X2 U19946 ( .A1(n7925), .A2(n27587), .ZN(n32472) );
  NAND2_X1 U19948 ( .A1(n12235), .A2(n7928), .ZN(n7927) );
  NAND2_X1 U19949 ( .A1(n12235), .A2(n12232), .ZN(n14152) );
  INV_X1 U19950 ( .A(n51641), .ZN(n12401) );
  NAND2_X1 U19951 ( .A1(n12236), .A2(n14145), .ZN(n7929) );
  NAND3_X1 U19952 ( .A1(n38550), .A2(n38212), .A3(n6734), .ZN(n7931) );
  NAND2_X1 U19953 ( .A1(n38213), .A2(n36141), .ZN(n7932) );
  INV_X1 U19954 ( .A(n31603), .ZN(n32636) );
  XNOR2_X1 U19955 ( .A(n24438), .B(n7935), .ZN(n7934) );
  XNOR2_X1 U19956 ( .A(n25071), .B(n25727), .ZN(n7935) );
  NAND2_X1 U19957 ( .A1(n21310), .A2(n7937), .ZN(n21311) );
  INV_X1 U19958 ( .A(n24279), .ZN(n7938) );
  XNOR2_X1 U19960 ( .A(n7939), .B(n43728), .ZN(n27267) );
  XNOR2_X1 U19961 ( .A(n7939), .B(n28076), .ZN(n28077) );
  XNOR2_X1 U19962 ( .A(n25365), .B(n7939), .ZN(n25366) );
  NAND3_X2 U19963 ( .A1(n22173), .A2(n22174), .A3(n7940), .ZN(n7939) );
  NAND3_X1 U19966 ( .A1(n30710), .A2(n30712), .A3(n29854), .ZN(n7943) );
  NAND2_X1 U19967 ( .A1(n20669), .A2(n7951), .ZN(n7950) );
  INV_X1 U19968 ( .A(n10256), .ZN(n7952) );
  NAND2_X1 U19969 ( .A1(n10248), .A2(n10249), .ZN(n7953) );
  NAND3_X1 U19972 ( .A1(n13324), .A2(n14607), .A3(n14605), .ZN(n13325) );
  AND2_X1 U19973 ( .A1(n14610), .A2(n14601), .ZN(n14607) );
  NAND2_X1 U19974 ( .A1(n30058), .A2(n7957), .ZN(n29588) );
  NAND2_X1 U19975 ( .A1(n18887), .A2(n19794), .ZN(n7958) );
  XNOR2_X1 U19976 ( .A(n35468), .B(n34779), .ZN(n34780) );
  NAND2_X1 U19977 ( .A1(n7962), .A2(n31641), .ZN(n7959) );
  NAND2_X1 U19978 ( .A1(n7963), .A2(n31632), .ZN(n7960) );
  AOI21_X1 U19979 ( .B1(n31639), .B2(n7961), .A(n706), .ZN(n7962) );
  OAI21_X1 U19980 ( .B1(n31630), .B2(n31631), .A(n31629), .ZN(n7963) );
  INV_X1 U19981 ( .A(n7964), .ZN(n7969) );
  NAND2_X1 U19982 ( .A1(n7970), .A2(n11631), .ZN(n7965) );
  NAND2_X1 U19983 ( .A1(n7969), .A2(n7968), .ZN(n7967) );
  OAI22_X1 U19984 ( .A1(n11628), .A2(n11629), .B1(n11630), .B2(n11632), .ZN(
        n7970) );
  INV_X1 U19985 ( .A(n11461), .ZN(n11632) );
  XNOR2_X1 U19987 ( .A(n22926), .B(n7971), .ZN(n22927) );
  XNOR2_X1 U19988 ( .A(n23122), .B(n7971), .ZN(n24705) );
  XNOR2_X1 U19989 ( .A(n25563), .B(n7971), .ZN(n26009) );
  NAND2_X1 U19990 ( .A1(n732), .A2(n7972), .ZN(n8649) );
  OR2_X2 U19991 ( .A1(n7973), .A2(n29462), .ZN(n27015) );
  NAND2_X1 U19995 ( .A1(n7977), .A2(n40388), .ZN(n39835) );
  NAND2_X1 U19996 ( .A1(n33270), .A2(n36317), .ZN(n7976) );
  OAI211_X1 U19997 ( .C1(n31517), .C2(n31518), .A(n7978), .B(n31516), .ZN(
        n31520) );
  INV_X1 U19998 ( .A(n30936), .ZN(n7978) );
  NAND4_X1 U19999 ( .A1(n7979), .A2(n38838), .A3(n39943), .A4(n39754), .ZN(
        n38834) );
  NAND3_X1 U20000 ( .A1(n39762), .A2(n7979), .A3(n38839), .ZN(n38840) );
  NAND2_X1 U20002 ( .A1(n11824), .A2(n11823), .ZN(n7981) );
  NOR2_X1 U20004 ( .A1(n7986), .A2(n7985), .ZN(n37951) );
  NAND2_X1 U20005 ( .A1(n41539), .A2(n40943), .ZN(n8754) );
  NAND2_X1 U20006 ( .A1(n23473), .A2(n21947), .ZN(n23464) );
  NAND2_X1 U20007 ( .A1(n38284), .A2(n38272), .ZN(n38286) );
  INV_X1 U20008 ( .A(n20116), .ZN(n20120) );
  AND2_X1 U20010 ( .A1(n22386), .A2(n50977), .ZN(n22376) );
  NAND2_X1 U20011 ( .A1(n19710), .A2(n19709), .ZN(n7988) );
  NAND3_X1 U20012 ( .A1(n19634), .A2(n19635), .A3(n19633), .ZN(n19707) );
  NAND2_X2 U20014 ( .A1(n7991), .A2(n26651), .ZN(n29308) );
  INV_X1 U20015 ( .A(n28695), .ZN(n7991) );
  XNOR2_X2 U20016 ( .A(n25698), .B(n25699), .ZN(n28695) );
  AND2_X1 U20017 ( .A1(n11234), .A2(n7992), .ZN(n11627) );
  NAND2_X1 U20018 ( .A1(n20317), .A2(n2403), .ZN(n7995) );
  NAND2_X1 U20019 ( .A1(n31891), .A2(n31422), .ZN(n31144) );
  NAND3_X1 U20020 ( .A1(n27848), .A2(n29306), .A3(n27847), .ZN(n7996) );
  OR2_X2 U20021 ( .A1(n40939), .A2(n40940), .ZN(n41544) );
  NAND2_X1 U20022 ( .A1(n7998), .A2(n39378), .ZN(n39200) );
  XNOR2_X1 U20025 ( .A(n8003), .B(n36934), .ZN(n36936) );
  XNOR2_X1 U20026 ( .A(n8004), .B(n36933), .ZN(n8003) );
  XNOR2_X1 U20027 ( .A(n36930), .B(n8005), .ZN(n8004) );
  XNOR2_X1 U20028 ( .A(n36931), .B(n36929), .ZN(n8005) );
  NAND2_X1 U20029 ( .A1(n50541), .A2(n50555), .ZN(n50518) );
  NAND2_X1 U20030 ( .A1(n50553), .A2(n50552), .ZN(n50541) );
  NAND2_X1 U20031 ( .A1(n47041), .A2(n50266), .ZN(n8007) );
  NAND2_X1 U20032 ( .A1(n8014), .A2(n34086), .ZN(n8008) );
  NAND2_X1 U20033 ( .A1(n19070), .A2(n16807), .ZN(n18354) );
  MUX2_X1 U20034 ( .A(n16809), .B(n16810), .S(n19070), .Z(n16811) );
  INV_X1 U20035 ( .A(n50638), .ZN(n50642) );
  INV_X1 U20036 ( .A(n52081), .ZN(n8018) );
  NOR2_X1 U20037 ( .A1(n8019), .A2(n30798), .ZN(n29904) );
  NAND2_X1 U20038 ( .A1(n29907), .A2(n29905), .ZN(n30798) );
  NAND3_X1 U20039 ( .A1(n29907), .A2(n2524), .A3(n29905), .ZN(n23657) );
  INV_X1 U20040 ( .A(n30789), .ZN(n8019) );
  NAND2_X1 U20042 ( .A1(n51709), .A2(n642), .ZN(n12525) );
  NAND2_X1 U20043 ( .A1(n47150), .A2(n44471), .ZN(n45158) );
  XNOR2_X1 U20046 ( .A(n8027), .B(n16497), .ZN(n8026) );
  XNOR2_X1 U20047 ( .A(n16507), .B(n2317), .ZN(n8027) );
  INV_X1 U20048 ( .A(n18152), .ZN(n8029) );
  INV_X1 U20050 ( .A(n39854), .ZN(n8032) );
  NOR2_X1 U20051 ( .A1(n21204), .A2(n8036), .ZN(n8035) );
  XNOR2_X1 U20052 ( .A(n34294), .B(n35278), .ZN(n8037) );
  OAI21_X1 U20053 ( .B1(n32149), .B2(n8041), .A(n31864), .ZN(n31865) );
  OR2_X1 U20055 ( .A1(n32784), .A2(n32785), .ZN(n8042) );
  NAND2_X1 U20056 ( .A1(n32785), .A2(n32788), .ZN(n8043) );
  NAND2_X1 U20057 ( .A1(n10368), .A2(n9632), .ZN(n10694) );
  NOR2_X2 U20058 ( .A1(n9406), .A2(n9405), .ZN(n9632) );
  XNOR2_X1 U20060 ( .A(n52103), .B(n41888), .ZN(n8046) );
  NAND2_X1 U20061 ( .A1(n8047), .A2(n39168), .ZN(n39170) );
  NAND2_X1 U20062 ( .A1(n39167), .A2(n419), .ZN(n8048) );
  NOR2_X1 U20063 ( .A1(n38675), .A2(n51496), .ZN(n39166) );
  NAND2_X1 U20064 ( .A1(n10383), .A2(n8050), .ZN(n9602) );
  OAI21_X1 U20065 ( .B1(n8052), .B2(n21393), .A(n17982), .ZN(n8051) );
  NAND2_X1 U20066 ( .A1(n22916), .A2(n22367), .ZN(n22164) );
  AND2_X1 U20067 ( .A1(n8053), .A2(n26807), .ZN(n8054) );
  NAND2_X1 U20068 ( .A1(n27641), .A2(n8055), .ZN(n8053) );
  NAND3_X2 U20069 ( .A1(n26809), .A2(n8054), .A3(n26808), .ZN(n31490) );
  NAND2_X1 U20070 ( .A1(n48125), .A2(n48124), .ZN(n48126) );
  NAND2_X1 U20071 ( .A1(n2742), .A2(n8056), .ZN(n45578) );
  NOR2_X1 U20072 ( .A1(n48416), .A2(n48404), .ZN(n8056) );
  OAI21_X1 U20073 ( .B1(n48402), .B2(n8057), .A(n2447), .ZN(n48407) );
  NOR2_X1 U20074 ( .A1(n8060), .A2(n48116), .ZN(n8059) );
  NAND2_X1 U20075 ( .A1(n46547), .A2(n48112), .ZN(n8060) );
  NAND3_X1 U20076 ( .A1(n45609), .A2(n45610), .A3(n8067), .ZN(n8066) );
  NAND2_X1 U20078 ( .A1(n8072), .A2(n39760), .ZN(n8071) );
  AOI21_X1 U20080 ( .B1(n8073), .B2(n12683), .A(n12461), .ZN(n8246) );
  AND2_X1 U20081 ( .A1(n8906), .A2(n7354), .ZN(n12683) );
  INV_X1 U20082 ( .A(n14252), .ZN(n8075) );
  AND2_X1 U20084 ( .A1(n8077), .A2(n2436), .ZN(n38718) );
  NOR2_X2 U20085 ( .A1(n41355), .A2(n40740), .ZN(n40751) );
  AOI22_X1 U20086 ( .A1(n29169), .A2(n29172), .B1(n29152), .B2(n8082), .ZN(
        n26485) );
  OR2_X1 U20087 ( .A1(n27955), .A2(n8082), .ZN(n8136) );
  XNOR2_X2 U20088 ( .A(Key[20]), .B(Ciphertext[73]), .ZN(n11581) );
  XNOR2_X1 U20089 ( .A(n15720), .B(n17284), .ZN(n15722) );
  INV_X1 U20090 ( .A(n15719), .ZN(n17186) );
  NAND2_X1 U20092 ( .A1(n50262), .A2(n8084), .ZN(n47067) );
  NAND3_X1 U20093 ( .A1(n47040), .A2(n8451), .A3(n8085), .ZN(n47041) );
  NAND2_X1 U20094 ( .A1(n31697), .A2(n8086), .ZN(n8087) );
  XNOR2_X1 U20095 ( .A(n8087), .B(n35293), .ZN(n35294) );
  XNOR2_X1 U20096 ( .A(n37137), .B(n8087), .ZN(n35383) );
  NAND2_X1 U20098 ( .A1(n27166), .A2(n8091), .ZN(n27541) );
  INV_X1 U20099 ( .A(n29848), .ZN(n8091) );
  NAND4_X1 U20100 ( .A1(n8092), .A2(n26757), .A3(n26758), .A4(n26759), .ZN(
        n26770) );
  OR2_X1 U20101 ( .A1(n26753), .A2(n51111), .ZN(n8093) );
  NAND4_X1 U20102 ( .A1(n20228), .A2(n20682), .A3(n51090), .A4(n20232), .ZN(
        n8095) );
  NAND2_X1 U20103 ( .A1(n48488), .A2(n48248), .ZN(n8097) );
  NAND2_X1 U20104 ( .A1(n11065), .A2(n2211), .ZN(n8098) );
  NAND3_X1 U20105 ( .A1(n48398), .A2(n48399), .A3(n8100), .ZN(n48401) );
  NAND3_X1 U20106 ( .A1(n8101), .A2(n48389), .A3(n48390), .ZN(n8100) );
  NAND2_X1 U20107 ( .A1(n13277), .A2(n14763), .ZN(n13282) );
  NAND2_X1 U20108 ( .A1(n26197), .A2(n29568), .ZN(n29554) );
  NAND2_X1 U20111 ( .A1(n48392), .A2(n8104), .ZN(n48395) );
  NAND2_X1 U20112 ( .A1(n48380), .A2(n8104), .ZN(n48360) );
  NAND2_X1 U20113 ( .A1(n48329), .A2(n8104), .ZN(n48299) );
  NAND3_X1 U20114 ( .A1(n48341), .A2(n8104), .A3(n52172), .ZN(n48342) );
  NAND3_X1 U20115 ( .A1(n48387), .A2(n8104), .A3(n48388), .ZN(n48389) );
  XNOR2_X1 U20116 ( .A(n16920), .B(n2216), .ZN(n15125) );
  NAND4_X2 U20117 ( .A1(n34672), .A2(n34673), .A3(n8110), .A4(n34671), .ZN(
        n8204) );
  INV_X1 U20118 ( .A(n46337), .ZN(n48411) );
  NOR2_X1 U20119 ( .A1(n48173), .A2(n46337), .ZN(n8111) );
  NOR2_X1 U20120 ( .A1(n8113), .A2(n8112), .ZN(n30970) );
  INV_X1 U20121 ( .A(n33032), .ZN(n8112) );
  NAND2_X1 U20123 ( .A1(n47360), .A2(n8115), .ZN(n8114) );
  NAND3_X1 U20124 ( .A1(n49976), .A2(n49975), .A3(n8116), .ZN(n8115) );
  OR2_X1 U20125 ( .A1(n49977), .A2(n49978), .ZN(n8116) );
  XNOR2_X1 U20126 ( .A(n8120), .B(n26609), .ZN(n8119) );
  NAND3_X1 U20127 ( .A1(n2470), .A2(n12753), .A3(n8121), .ZN(n11306) );
  OR2_X1 U20128 ( .A1(n38740), .A2(n41355), .ZN(n41347) );
  INV_X1 U20129 ( .A(n10398), .ZN(n9429) );
  XNOR2_X1 U20130 ( .A(n45091), .B(n43363), .ZN(n42264) );
  NAND4_X2 U20131 ( .A1(n8124), .A2(n39318), .A3(n41242), .A4(n39317), .ZN(
        n43943) );
  OAI21_X1 U20133 ( .B1(n14634), .B2(n14633), .A(n14632), .ZN(n8126) );
  INV_X1 U20134 ( .A(n14642), .ZN(n8128) );
  NOR2_X1 U20135 ( .A1(n46311), .A2(n8130), .ZN(n8132) );
  XNOR2_X1 U20136 ( .A(n8132), .B(n4639), .ZN(Plaintext[90]) );
  OR2_X1 U20137 ( .A1(n49002), .A2(n46279), .ZN(n8133) );
  OAI21_X1 U20138 ( .B1(n39174), .B2(n38667), .A(n8134), .ZN(n38668) );
  NAND2_X1 U20139 ( .A1(n32214), .A2(n32210), .ZN(n31764) );
  XNOR2_X2 U20140 ( .A(Key[123]), .B(Ciphertext[74]), .ZN(n11530) );
  NAND3_X1 U20141 ( .A1(n11581), .A2(n12574), .A3(n11530), .ZN(n11191) );
  INV_X1 U20142 ( .A(n11186), .ZN(n12574) );
  XNOR2_X2 U20143 ( .A(n42270), .B(n8138), .ZN(n49170) );
  NAND2_X1 U20144 ( .A1(n15440), .A2(n8140), .ZN(n14831) );
  NAND2_X1 U20145 ( .A1(n15325), .A2(n15440), .ZN(n15338) );
  NOR2_X1 U20146 ( .A1(n40921), .A2(n8142), .ZN(n40965) );
  NAND2_X1 U20147 ( .A1(n40959), .A2(n8143), .ZN(n8142) );
  AND2_X1 U20148 ( .A1(n41375), .A2(n41374), .ZN(n8143) );
  INV_X1 U20149 ( .A(n45751), .ZN(n8144) );
  NOR2_X1 U20150 ( .A1(n45713), .A2(n45754), .ZN(n45747) );
  NAND2_X1 U20151 ( .A1(n13723), .A2(n15285), .ZN(n8146) );
  NAND2_X1 U20152 ( .A1(n15273), .A2(n15279), .ZN(n8147) );
  INV_X1 U20153 ( .A(n15285), .ZN(n14057) );
  NAND2_X1 U20154 ( .A1(n18590), .A2(n21435), .ZN(n8148) );
  NAND2_X1 U20155 ( .A1(n20321), .A2(n21438), .ZN(n19166) );
  NAND3_X1 U20156 ( .A1(n23926), .A2(n8149), .A3(n23911), .ZN(n21502) );
  INV_X1 U20159 ( .A(n39943), .ZN(n8150) );
  NOR2_X1 U20160 ( .A1(n8153), .A2(n8152), .ZN(n8151) );
  NAND2_X1 U20161 ( .A1(n23144), .A2(n23145), .ZN(n8152) );
  AOI21_X1 U20162 ( .B1(n12497), .B2(n8154), .A(n642), .ZN(n12499) );
  INV_X1 U20163 ( .A(n8154), .ZN(n12495) );
  NAND3_X1 U20164 ( .A1(n47665), .A2(n47664), .A3(n47666), .ZN(n8155) );
  NAND4_X2 U20165 ( .A1(n8158), .A2(n45767), .A3(n45769), .A4(n8156), .ZN(
        n47689) );
  NAND3_X1 U20166 ( .A1(n8157), .A2(n45765), .A3(n47909), .ZN(n8156) );
  NAND2_X1 U20167 ( .A1(n23336), .A2(n21755), .ZN(n21757) );
  OAI21_X1 U20169 ( .B1(n10706), .B2(n8161), .A(n10705), .ZN(n10707) );
  NAND2_X1 U20171 ( .A1(n31358), .A2(n38558), .ZN(n35179) );
  NAND2_X1 U20172 ( .A1(n41446), .A2(n41442), .ZN(n38909) );
  OR2_X2 U20173 ( .A1(n36310), .A2(n36311), .ZN(n41442) );
  AND2_X1 U20174 ( .A1(n45752), .A2(n8168), .ZN(n8166) );
  AOI22_X1 U20175 ( .A1(n8166), .A2(n48806), .B1(n48799), .B2(n48816), .ZN(
        n8164) );
  OAI211_X1 U20176 ( .C1(n48799), .C2(n45711), .A(n52091), .B(n48793), .ZN(
        n8165) );
  NAND2_X1 U20177 ( .A1(n45712), .A2(n48798), .ZN(n8167) );
  NOR2_X1 U20178 ( .A1(n48792), .A2(n48834), .ZN(n8168) );
  NAND3_X1 U20179 ( .A1(n8169), .A2(n10875), .A3(n10874), .ZN(n10876) );
  NAND2_X1 U20180 ( .A1(n8170), .A2(n15171), .ZN(n8169) );
  NAND2_X1 U20181 ( .A1(n29908), .A2(n30780), .ZN(n8171) );
  NAND2_X1 U20182 ( .A1(n30782), .A2(n30795), .ZN(n8172) );
  NAND2_X1 U20183 ( .A1(n43329), .A2(n37605), .ZN(n37609) );
  OR2_X1 U20184 ( .A1(n39393), .A2(n38998), .ZN(n34904) );
  NAND3_X1 U20185 ( .A1(n8173), .A2(n39003), .A3(n38995), .ZN(n38996) );
  INV_X1 U20186 ( .A(n39393), .ZN(n8173) );
  NAND2_X1 U20187 ( .A1(n17546), .A2(n18331), .ZN(n18070) );
  OAI21_X1 U20188 ( .B1(n9906), .B2(n9477), .A(n8174), .ZN(n9478) );
  XNOR2_X1 U20190 ( .A(n8179), .B(n8178), .ZN(n26355) );
  AOI21_X1 U20191 ( .B1(n8182), .B2(n30709), .A(n8181), .ZN(n8180) );
  NOR2_X1 U20192 ( .A1(n30710), .A2(n30709), .ZN(n8181) );
  NAND2_X1 U20193 ( .A1(n30708), .A2(n30721), .ZN(n8183) );
  NAND2_X1 U20194 ( .A1(n28915), .A2(n29006), .ZN(n28922) );
  NAND2_X1 U20195 ( .A1(n28020), .A2(n29013), .ZN(n8184) );
  INV_X1 U20197 ( .A(n13088), .ZN(n12915) );
  NAND2_X1 U20199 ( .A1(n39877), .A2(n41170), .ZN(n8193) );
  INV_X2 U20200 ( .A(n50189), .ZN(n50222) );
  NOR2_X1 U20201 ( .A1(n39754), .A2(n39937), .ZN(n8199) );
  NAND2_X1 U20202 ( .A1(n8201), .A2(n48156), .ZN(n48118) );
  NAND2_X1 U20203 ( .A1(n48155), .A2(n48140), .ZN(n48115) );
  INV_X1 U20204 ( .A(n31495), .ZN(n8203) );
  XNOR2_X1 U20205 ( .A(n8515), .B(n8204), .ZN(n41858) );
  XNOR2_X1 U20206 ( .A(n52096), .B(n8204), .ZN(n40881) );
  XNOR2_X1 U20207 ( .A(n8204), .B(n46113), .ZN(n46114) );
  XNOR2_X1 U20208 ( .A(n8204), .B(n43622), .ZN(n43624) );
  XNOR2_X1 U20209 ( .A(n8204), .B(n46111), .ZN(n44880) );
  NAND2_X1 U20210 ( .A1(n27677), .A2(n27690), .ZN(n26815) );
  NAND3_X1 U20211 ( .A1(n20721), .A2(n22275), .A3(n23570), .ZN(n20723) );
  NAND2_X1 U20212 ( .A1(n52108), .A2(n39144), .ZN(n34667) );
  NAND2_X1 U20213 ( .A1(n41088), .A2(n8206), .ZN(n38361) );
  AND2_X1 U20214 ( .A1(n52108), .A2(n39713), .ZN(n8206) );
  XNOR2_X1 U20215 ( .A(n38870), .B(n38869), .ZN(n34669) );
  NAND2_X1 U20216 ( .A1(n41078), .A2(n52108), .ZN(n41081) );
  AND2_X2 U20217 ( .A1(n8207), .A2(n46380), .ZN(n46501) );
  INV_X1 U20218 ( .A(n45661), .ZN(n46493) );
  INV_X1 U20219 ( .A(n45661), .ZN(n8207) );
  XNOR2_X1 U20220 ( .A(n25886), .B(n8208), .ZN(n25887) );
  XNOR2_X1 U20221 ( .A(n27467), .B(n8208), .ZN(n24494) );
  XNOR2_X1 U20222 ( .A(n8208), .B(n24757), .ZN(n26190) );
  XNOR2_X1 U20223 ( .A(n22282), .B(n8208), .ZN(n25289) );
  XNOR2_X1 U20224 ( .A(n26034), .B(n8208), .ZN(n26036) );
  XNOR2_X2 U20225 ( .A(n22281), .B(n28353), .ZN(n8208) );
  AND2_X1 U20226 ( .A1(n41690), .A2(n41706), .ZN(n41164) );
  NAND3_X1 U20227 ( .A1(n48148), .A2(n48149), .A3(n2397), .ZN(Plaintext[45])
         );
  NAND3_X1 U20229 ( .A1(n46476), .A2(n46477), .A3(n8210), .ZN(n46481) );
  INV_X1 U20230 ( .A(n8212), .ZN(n14847) );
  XNOR2_X1 U20231 ( .A(n52200), .B(n8212), .ZN(n14050) );
  XNOR2_X1 U20232 ( .A(n18579), .B(n8212), .ZN(n17647) );
  INV_X1 U20233 ( .A(n18795), .ZN(n8211) );
  XNOR2_X1 U20234 ( .A(n8212), .B(n16542), .ZN(n16543) );
  NAND2_X1 U20235 ( .A1(n8217), .A2(n23174), .ZN(n8216) );
  NAND2_X1 U20237 ( .A1(n41081), .A2(n8218), .ZN(n41091) );
  NAND2_X1 U20238 ( .A1(n38868), .A2(n39140), .ZN(n8219) );
  XNOR2_X1 U20239 ( .A(n16176), .B(n8221), .ZN(n16290) );
  NAND2_X1 U20240 ( .A1(n13091), .A2(n641), .ZN(n8225) );
  OR2_X1 U20241 ( .A1(n14317), .A2(n8226), .ZN(n11798) );
  NAND2_X1 U20242 ( .A1(n8227), .A2(n13819), .ZN(n14315) );
  AOI21_X1 U20243 ( .B1(n14307), .B2(n8227), .A(n13819), .ZN(n13609) );
  NAND3_X1 U20244 ( .A1(n13827), .A2(n8227), .A3(n13826), .ZN(n13828) );
  AOI21_X1 U20245 ( .B1(n14304), .B2(n14305), .A(n8227), .ZN(n14329) );
  NAND3_X1 U20246 ( .A1(n8228), .A2(n32896), .A3(n32909), .ZN(n32545) );
  NAND2_X1 U20247 ( .A1(n36425), .A2(n36616), .ZN(n34924) );
  NAND3_X1 U20248 ( .A1(n20403), .A2(n8230), .A3(n22748), .ZN(n22937) );
  NAND2_X1 U20249 ( .A1(n22075), .A2(n8229), .ZN(n22076) );
  OAI211_X1 U20250 ( .C1(n39111), .C2(n39938), .A(n8231), .B(n38830), .ZN(
        n36504) );
  OR3_X1 U20251 ( .A1(n684), .A2(n39754), .A3(n39751), .ZN(n8231) );
  NAND2_X1 U20252 ( .A1(n20384), .A2(n20383), .ZN(n20385) );
  XNOR2_X1 U20253 ( .A(n26393), .B(n25430), .ZN(n25431) );
  NAND3_X1 U20254 ( .A1(n8234), .A2(n41332), .A3(n41330), .ZN(n41335) );
  XNOR2_X1 U20255 ( .A(n8235), .B(n41328), .ZN(n8234) );
  NAND2_X1 U20256 ( .A1(n38559), .A2(n8285), .ZN(n8236) );
  NAND2_X1 U20257 ( .A1(n30853), .A2(n31637), .ZN(n8241) );
  NAND3_X1 U20258 ( .A1(n31581), .A2(n30854), .A3(n31636), .ZN(n8238) );
  NAND2_X1 U20259 ( .A1(n31638), .A2(n30855), .ZN(n31581) );
  OAI211_X1 U20261 ( .C1(n50473), .C2(n50458), .A(n8244), .B(n8243), .ZN(n8245) );
  NAND2_X1 U20262 ( .A1(n50458), .A2(n50457), .ZN(n50477) );
  OAI21_X1 U20263 ( .B1(n19749), .B2(n22736), .A(n5371), .ZN(n19748) );
  NAND3_X1 U20264 ( .A1(n8251), .A2(n714), .A3(n32395), .ZN(n8252) );
  OAI21_X1 U20265 ( .B1(n32394), .B2(n7430), .A(n51640), .ZN(n8251) );
  INV_X1 U20266 ( .A(n32414), .ZN(n8253) );
  XNOR2_X1 U20267 ( .A(n26053), .B(n28129), .ZN(n26222) );
  XNOR2_X2 U20268 ( .A(n25825), .B(n25903), .ZN(n28129) );
  AND2_X1 U20269 ( .A1(n23769), .A2(n23768), .ZN(n8255) );
  XNOR2_X1 U20270 ( .A(n24948), .B(n27242), .ZN(n25270) );
  INV_X1 U20271 ( .A(n25270), .ZN(n24950) );
  NAND3_X1 U20272 ( .A1(n678), .A2(n40860), .A3(n2490), .ZN(n38355) );
  AND3_X2 U20273 ( .A1(n8259), .A2(n8258), .A3(n8257), .ZN(n48353) );
  NAND2_X1 U20274 ( .A1(n48264), .A2(n48265), .ZN(n8257) );
  NAND2_X1 U20275 ( .A1(n48266), .A2(n48433), .ZN(n8258) );
  NAND3_X2 U20278 ( .A1(n8261), .A2(n19974), .A3(n19975), .ZN(n24041) );
  NAND2_X1 U20279 ( .A1(n19973), .A2(n20827), .ZN(n8262) );
  NAND2_X1 U20280 ( .A1(n19971), .A2(n19972), .ZN(n8263) );
  NAND2_X1 U20281 ( .A1(n22129), .A2(n52134), .ZN(n23237) );
  XNOR2_X1 U20282 ( .A(n25832), .B(n8267), .ZN(n25228) );
  XNOR2_X1 U20283 ( .A(n22810), .B(n25831), .ZN(n8267) );
  XNOR2_X1 U20284 ( .A(n27506), .B(n22747), .ZN(n25832) );
  XNOR2_X1 U20285 ( .A(n42638), .B(n8268), .ZN(n42639) );
  XNOR2_X1 U20286 ( .A(n44567), .B(n45304), .ZN(n8270) );
  XNOR2_X1 U20287 ( .A(n43352), .B(n44971), .ZN(n43039) );
  NAND3_X1 U20290 ( .A1(n47195), .A2(n49442), .A3(n51453), .ZN(n8278) );
  NAND3_X1 U20291 ( .A1(n37782), .A2(n36191), .A3(n39335), .ZN(n36195) );
  INV_X1 U20292 ( .A(n39335), .ZN(n33464) );
  NAND4_X1 U20293 ( .A1(n13103), .A2(n13092), .A3(n641), .A4(n13086), .ZN(
        n8279) );
  NAND3_X1 U20294 ( .A1(n11163), .A2(n11164), .A3(n8279), .ZN(n11165) );
  XNOR2_X1 U20295 ( .A(n8283), .B(n36940), .ZN(n33889) );
  INV_X1 U20297 ( .A(n18360), .ZN(n18345) );
  NAND2_X1 U20298 ( .A1(n51756), .A2(n20132), .ZN(n18360) );
  NAND2_X1 U20300 ( .A1(n8286), .A2(n10174), .ZN(n9456) );
  NOR2_X1 U20301 ( .A1(n10187), .A2(n8286), .ZN(n10188) );
  AOI22_X1 U20302 ( .A1(n8287), .A2(n21945), .B1(n23153), .B2(n16688), .ZN(
        n16694) );
  OAI21_X1 U20303 ( .B1(n27065), .B2(n736), .A(n8331), .ZN(n8289) );
  NAND2_X1 U20304 ( .A1(n50945), .A2(n50944), .ZN(n50963) );
  NAND2_X1 U20305 ( .A1(n8297), .A2(n9328), .ZN(n8295) );
  NAND2_X1 U20306 ( .A1(n11625), .A2(n11477), .ZN(n8297) );
  NAND3_X1 U20307 ( .A1(n18864), .A2(n8300), .A3(n8299), .ZN(n8298) );
  NAND2_X1 U20308 ( .A1(n18105), .A2(n20228), .ZN(n8299) );
  NAND2_X1 U20309 ( .A1(n1597), .A2(n8302), .ZN(n8301) );
  NAND3_X1 U20310 ( .A1(n8402), .A2(n23316), .A3(n23310), .ZN(n8304) );
  NAND2_X1 U20311 ( .A1(n8304), .A2(n8303), .ZN(n21005) );
  NOR2_X1 U20312 ( .A1(n27820), .A2(n27808), .ZN(n26324) );
  OAI211_X1 U20313 ( .C1(n7766), .C2(n8307), .A(n48156), .B(n8305), .ZN(n8308)
         );
  INV_X1 U20314 ( .A(n48154), .ZN(n8306) );
  NAND2_X1 U20315 ( .A1(n48093), .A2(n48094), .ZN(n8307) );
  INV_X1 U20316 ( .A(n22375), .ZN(n8310) );
  NAND2_X1 U20317 ( .A1(n12691), .A2(n12692), .ZN(n8312) );
  NAND2_X1 U20319 ( .A1(n41085), .A2(n8316), .ZN(n8317) );
  NAND2_X1 U20320 ( .A1(n39708), .A2(n8317), .ZN(n38872) );
  INV_X1 U20321 ( .A(n19210), .ZN(n8319) );
  XNOR2_X2 U20322 ( .A(n8318), .B(n17143), .ZN(n21186) );
  XNOR2_X1 U20323 ( .A(n17144), .B(n8319), .ZN(n8318) );
  NAND2_X1 U20324 ( .A1(n17071), .A2(n51756), .ZN(n8320) );
  XNOR2_X1 U20325 ( .A(n8323), .B(n24591), .ZN(n8596) );
  NAND2_X1 U20326 ( .A1(n9349), .A2(n11709), .ZN(n8325) );
  NAND2_X1 U20327 ( .A1(n9350), .A2(n11200), .ZN(n8326) );
  XNOR2_X2 U20328 ( .A(n35544), .B(n37086), .ZN(n34754) );
  NAND2_X1 U20329 ( .A1(n31942), .A2(n31941), .ZN(n8330) );
  NAND2_X1 U20330 ( .A1(n31332), .A2(n31331), .ZN(n31942) );
  INV_X2 U20331 ( .A(n30037), .ZN(n31931) );
  NAND2_X1 U20332 ( .A1(n30037), .A2(n31340), .ZN(n31334) );
  NAND2_X1 U20333 ( .A1(n7044), .A2(n8334), .ZN(n44573) );
  XNOR2_X1 U20334 ( .A(n35474), .B(n33537), .ZN(n8336) );
  XNOR2_X1 U20335 ( .A(n44146), .B(n43751), .ZN(n43149) );
  NAND2_X1 U20336 ( .A1(n39612), .A2(n41007), .ZN(n8337) );
  XNOR2_X1 U20337 ( .A(n16920), .B(n16527), .ZN(n17356) );
  XNOR2_X2 U20338 ( .A(n17264), .B(n14803), .ZN(n16527) );
  NAND4_X2 U20339 ( .A1(n14800), .A2(n14801), .A3(n8341), .A4(n14802), .ZN(
        n17264) );
  NOR2_X1 U20340 ( .A1(n8342), .A2(n14792), .ZN(n8341) );
  NOR2_X1 U20341 ( .A1(n32486), .A2(n32478), .ZN(n8343) );
  NAND4_X1 U20342 ( .A1(n8345), .A2(n32483), .A3(n8343), .A4(n8344), .ZN(
        n32023) );
  XNOR2_X2 U20344 ( .A(n43275), .B(n43274), .ZN(n49667) );
  NAND2_X1 U20345 ( .A1(n32424), .A2(n32428), .ZN(n31260) );
  INV_X1 U20346 ( .A(n12059), .ZN(n8347) );
  NAND2_X1 U20347 ( .A1(n8347), .A2(n12052), .ZN(n10660) );
  NOR2_X1 U20348 ( .A1(n12059), .A2(n8349), .ZN(n8348) );
  NOR2_X1 U20349 ( .A1(n51347), .A2(n12950), .ZN(n8350) );
  INV_X1 U20350 ( .A(n12950), .ZN(n14674) );
  XNOR2_X1 U20351 ( .A(n35760), .B(n34627), .ZN(n8352) );
  XNOR2_X2 U20352 ( .A(n8352), .B(n8351), .ZN(n37646) );
  INV_X1 U20353 ( .A(n22207), .ZN(n22766) );
  XNOR2_X1 U20354 ( .A(n8357), .B(n2215), .ZN(n8356) );
  XNOR2_X1 U20355 ( .A(n15653), .B(n16098), .ZN(n8357) );
  NOR2_X1 U20356 ( .A1(n32473), .A2(n8361), .ZN(n8360) );
  INV_X1 U20358 ( .A(n28870), .ZN(n8364) );
  INV_X1 U20359 ( .A(n14365), .ZN(n14366) );
  XNOR2_X2 U20360 ( .A(n15996), .B(n19272), .ZN(n21620) );
  NAND2_X1 U20361 ( .A1(n32684), .A2(n31660), .ZN(n31659) );
  INV_X1 U20363 ( .A(n19612), .ZN(n8370) );
  XNOR2_X1 U20364 ( .A(n42504), .B(n52103), .ZN(n43892) );
  XNOR2_X2 U20365 ( .A(n44154), .B(n44156), .ZN(n42504) );
  NAND4_X2 U20366 ( .A1(n8373), .A2(n40019), .A3(n40020), .A4(n8372), .ZN(
        n44156) );
  NAND2_X1 U20367 ( .A1(n40006), .A2(n40007), .ZN(n8373) );
  NOR2_X1 U20368 ( .A1(n8375), .A2(n35207), .ZN(n8374) );
  NOR2_X2 U20369 ( .A1(n40014), .A2(n39103), .ZN(n39099) );
  NAND4_X2 U20371 ( .A1(n48471), .A2(n8379), .A3(n8380), .A4(n48472), .ZN(
        n48652) );
  NAND3_X1 U20372 ( .A1(n36459), .A2(n696), .A3(n36050), .ZN(n8381) );
  INV_X1 U20373 ( .A(n36045), .ZN(n35879) );
  INV_X1 U20374 ( .A(n36052), .ZN(n36589) );
  OAI21_X1 U20375 ( .B1(n15134), .B2(n8388), .A(n15137), .ZN(n8387) );
  AND2_X1 U20376 ( .A1(n15136), .A2(n15138), .ZN(n8388) );
  OAI21_X1 U20377 ( .B1(n41239), .B2(n41240), .A(n41238), .ZN(n8392) );
  INV_X1 U20378 ( .A(n21504), .ZN(n8394) );
  NAND2_X1 U20379 ( .A1(n23895), .A2(n22521), .ZN(n22524) );
  NAND2_X1 U20381 ( .A1(n20488), .A2(n19359), .ZN(n21451) );
  XNOR2_X2 U20382 ( .A(n8396), .B(Key[87]), .ZN(n12161) );
  NAND2_X1 U20384 ( .A1(n13575), .A2(n13576), .ZN(n14276) );
  XNOR2_X1 U20386 ( .A(n15666), .B(n8399), .ZN(n8398) );
  XNOR2_X1 U20387 ( .A(n8400), .B(n19198), .ZN(n8399) );
  XNOR2_X1 U20388 ( .A(n14908), .B(n16320), .ZN(n8400) );
  NAND2_X1 U20389 ( .A1(n17532), .A2(n20015), .ZN(n8401) );
  NAND3_X1 U20390 ( .A1(n8639), .A2(n2197), .A3(n10008), .ZN(n8820) );
  XNOR2_X1 U20392 ( .A(n19196), .B(n8403), .ZN(n17766) );
  XNOR2_X1 U20393 ( .A(n18407), .B(n8403), .ZN(n16729) );
  XNOR2_X1 U20394 ( .A(n16624), .B(n8403), .ZN(n15321) );
  XNOR2_X1 U20395 ( .A(n17888), .B(n8403), .ZN(n17890) );
  NAND2_X1 U20396 ( .A1(n30081), .A2(n30082), .ZN(n30927) );
  NAND2_X1 U20397 ( .A1(n32334), .A2(n32335), .ZN(n8404) );
  XNOR2_X1 U20398 ( .A(n28083), .B(n8406), .ZN(n8405) );
  NAND3_X1 U20399 ( .A1(n39400), .A2(n38995), .A3(n3735), .ZN(n38993) );
  NAND2_X1 U20400 ( .A1(n8639), .A2(n8407), .ZN(n11021) );
  NAND2_X1 U20402 ( .A1(n30772), .A2(n29921), .ZN(n30752) );
  INV_X1 U20403 ( .A(n17037), .ZN(n8411) );
  XNOR2_X2 U20404 ( .A(n8413), .B(n37025), .ZN(n39369) );
  XNOR2_X1 U20405 ( .A(n8414), .B(n37019), .ZN(n8413) );
  XNOR2_X1 U20406 ( .A(n37022), .B(n37018), .ZN(n8414) );
  NAND2_X1 U20407 ( .A1(n14711), .A2(n14709), .ZN(n14200) );
  NAND2_X1 U20409 ( .A1(n28712), .A2(n29282), .ZN(n8417) );
  INV_X1 U20411 ( .A(n9249), .ZN(n8428) );
  NAND3_X2 U20412 ( .A1(n22069), .A2(n8433), .A3(n8430), .ZN(n25495) );
  NAND2_X1 U20413 ( .A1(n22060), .A2(n22059), .ZN(n8433) );
  NAND2_X1 U20414 ( .A1(n29304), .A2(n8436), .ZN(n8435) );
  OR2_X1 U20415 ( .A1(n51517), .A2(n28695), .ZN(n8436) );
  NOR2_X1 U20416 ( .A1(n28688), .A2(n26651), .ZN(n29304) );
  NAND2_X1 U20417 ( .A1(n8438), .A2(n10529), .ZN(n10634) );
  NAND4_X2 U20418 ( .A1(n13109), .A2(n13108), .A3(n13107), .A4(n8439), .ZN(
        n14427) );
  NAND2_X1 U20419 ( .A1(n13101), .A2(n13100), .ZN(n8440) );
  INV_X1 U20420 ( .A(n19119), .ZN(n8441) );
  XNOR2_X1 U20421 ( .A(n8442), .B(n8443), .ZN(n23938) );
  NAND3_X2 U20422 ( .A1(n21288), .A2(n21289), .A3(n8445), .ZN(n23175) );
  NAND4_X1 U20423 ( .A1(n8447), .A2(n47605), .A3(n47600), .A4(n47601), .ZN(
        n47602) );
  NAND2_X1 U20424 ( .A1(n47622), .A2(n47595), .ZN(n8447) );
  NAND3_X1 U20425 ( .A1(n43966), .A2(n43965), .A3(n8451), .ZN(n43984) );
  OAI21_X1 U20426 ( .B1(n47343), .B2(n47342), .A(n8452), .ZN(n47344) );
  NAND2_X1 U20427 ( .A1(n50252), .A2(n44001), .ZN(n8452) );
  INV_X1 U20428 ( .A(n29542), .ZN(n8454) );
  NAND2_X1 U20429 ( .A1(n10582), .A2(n10583), .ZN(n8456) );
  NAND2_X1 U20430 ( .A1(n18731), .A2(n21637), .ZN(n15999) );
  XNOR2_X1 U20431 ( .A(n35618), .B(n8460), .ZN(n34337) );
  NAND2_X1 U20432 ( .A1(n8462), .A2(n8461), .ZN(n39024) );
  OAI21_X1 U20433 ( .B1(n14827), .B2(n15435), .A(n15437), .ZN(n8463) );
  XNOR2_X1 U20434 ( .A(n593), .B(n26556), .ZN(n8464) );
  INV_X1 U20435 ( .A(n32105), .ZN(n32096) );
  NAND2_X1 U20436 ( .A1(n8466), .A2(n32088), .ZN(n32101) );
  NAND2_X1 U20437 ( .A1(n32565), .A2(n32087), .ZN(n8466) );
  NAND2_X1 U20438 ( .A1(n32103), .A2(n8467), .ZN(n32565) );
  NOR2_X1 U20439 ( .A1(n32105), .A2(n8468), .ZN(n8467) );
  INV_X1 U20440 ( .A(n32558), .ZN(n8468) );
  NAND2_X1 U20441 ( .A1(n8471), .A2(n46494), .ZN(n46407) );
  NAND3_X1 U20442 ( .A1(n8471), .A2(n46387), .A3(n46503), .ZN(n46188) );
  INV_X1 U20443 ( .A(n46386), .ZN(n8471) );
  AND2_X1 U20444 ( .A1(n49029), .A2(n49020), .ZN(n8472) );
  NAND2_X1 U20445 ( .A1(n37826), .A2(n37825), .ZN(n42212) );
  NOR2_X1 U20446 ( .A1(n8477), .A2(n2405), .ZN(n8476) );
  NAND2_X1 U20447 ( .A1(n37829), .A2(n37830), .ZN(n8477) );
  NAND3_X1 U20448 ( .A1(n39258), .A2(n8429), .A3(n8480), .ZN(n8478) );
  NAND2_X1 U20449 ( .A1(n11409), .A2(n12145), .ZN(n11402) );
  INV_X1 U20450 ( .A(n25813), .ZN(n23977) );
  XNOR2_X2 U20451 ( .A(n6563), .B(n8488), .ZN(n18942) );
  NAND2_X1 U20453 ( .A1(n20760), .A2(n8490), .ZN(n19288) );
  NAND2_X1 U20454 ( .A1(n21600), .A2(n21358), .ZN(n18685) );
  INV_X1 U20455 ( .A(n21360), .ZN(n8489) );
  NAND2_X1 U20457 ( .A1(n18723), .A2(n21609), .ZN(n8493) );
  NAND2_X1 U20460 ( .A1(n40293), .A2(n40049), .ZN(n41483) );
  XNOR2_X1 U20461 ( .A(n16701), .B(n47401), .ZN(n8501) );
  NAND2_X1 U20462 ( .A1(n51127), .A2(n19892), .ZN(n18938) );
  XNOR2_X2 U20463 ( .A(n40631), .B(n40630), .ZN(n44873) );
  NAND3_X1 U20464 ( .A1(n13599), .A2(n14318), .A3(n13598), .ZN(n8505) );
  NAND2_X1 U20465 ( .A1(n16882), .A2(n18932), .ZN(n8506) );
  NAND2_X1 U20466 ( .A1(n24283), .A2(n24287), .ZN(n21905) );
  INV_X1 U20467 ( .A(n51643), .ZN(n8508) );
  XNOR2_X1 U20468 ( .A(n34275), .B(n35810), .ZN(n35077) );
  XNOR2_X2 U20469 ( .A(n51739), .B(n51445), .ZN(n35810) );
  INV_X1 U20470 ( .A(n23001), .ZN(n22981) );
  NAND2_X1 U20471 ( .A1(n22983), .A2(n22434), .ZN(n23001) );
  INV_X1 U20473 ( .A(n38483), .ZN(n8509) );
  INV_X1 U20474 ( .A(n10498), .ZN(n8510) );
  NAND2_X1 U20476 ( .A1(n8514), .A2(n14999), .ZN(n13708) );
  NAND2_X1 U20477 ( .A1(n26905), .A2(n51351), .ZN(n29410) );
  XNOR2_X1 U20478 ( .A(n8515), .B(n4645), .ZN(n43245) );
  XNOR2_X1 U20479 ( .A(n40814), .B(n8515), .ZN(n42729) );
  NAND2_X1 U20481 ( .A1(n19620), .A2(n23485), .ZN(n8520) );
  NAND2_X1 U20482 ( .A1(n19624), .A2(n23483), .ZN(n8521) );
  NAND3_X1 U20483 ( .A1(n24036), .A2(n23671), .A3(n8524), .ZN(n23672) );
  INV_X1 U20484 ( .A(n354), .ZN(n8524) );
  NAND2_X1 U20485 ( .A1(n23675), .A2(n8525), .ZN(n22110) );
  NOR2_X1 U20486 ( .A1(n8526), .A2(n354), .ZN(n8525) );
  NAND2_X1 U20487 ( .A1(n9916), .A2(n9917), .ZN(n8527) );
  OR2_X2 U20488 ( .A1(n8529), .A2(n8530), .ZN(n50533) );
  NAND3_X1 U20489 ( .A1(n49744), .A2(n8533), .A3(n8531), .ZN(n8530) );
  NAND2_X1 U20490 ( .A1(n47015), .A2(n47309), .ZN(n8532) );
  NAND2_X1 U20492 ( .A1(n30470), .A2(n8536), .ZN(n8535) );
  NAND2_X1 U20493 ( .A1(n30469), .A2(n32417), .ZN(n8538) );
  NAND4_X1 U20494 ( .A1(n15302), .A2(n1486), .A3(n14929), .A4(n15304), .ZN(
        n12744) );
  AND2_X1 U20495 ( .A1(n38764), .A2(n41004), .ZN(n43335) );
  NAND2_X1 U20496 ( .A1(n32821), .A2(n32825), .ZN(n32415) );
  NAND4_X2 U20499 ( .A1(n8543), .A2(n32262), .A3(n32261), .A4(n32260), .ZN(
        n33973) );
  INV_X1 U20500 ( .A(n32238), .ZN(n8543) );
  INV_X1 U20502 ( .A(n14550), .ZN(n14534) );
  AND2_X1 U20504 ( .A1(n31654), .A2(n8547), .ZN(n8546) );
  NAND2_X1 U20505 ( .A1(n31646), .A2(n32463), .ZN(n8547) );
  NAND2_X1 U20506 ( .A1(n16878), .A2(n16877), .ZN(n8549) );
  NAND2_X1 U20507 ( .A1(n8551), .A2(n16876), .ZN(n8550) );
  NAND2_X1 U20508 ( .A1(n16874), .A2(n8552), .ZN(n8551) );
  NAND2_X1 U20512 ( .A1(n39386), .A2(n39192), .ZN(n39383) );
  NAND3_X1 U20513 ( .A1(n39386), .A2(n39192), .A3(n39376), .ZN(n38959) );
  NAND3_X1 U20514 ( .A1(n18933), .A2(n15636), .A3(n19886), .ZN(n8556) );
  INV_X1 U20515 ( .A(n15617), .ZN(n8557) );
  AOI22_X1 U20516 ( .A1(n21158), .A2(n22274), .B1(n23559), .B2(n21157), .ZN(
        n21159) );
  INV_X1 U20517 ( .A(n18086), .ZN(n18080) );
  NAND2_X1 U20518 ( .A1(n18086), .A2(n20504), .ZN(n8558) );
  NAND2_X1 U20519 ( .A1(n18087), .A2(n20504), .ZN(n8560) );
  NAND3_X1 U20520 ( .A1(n22361), .A2(n22912), .A3(n22360), .ZN(n22366) );
  NAND2_X1 U20521 ( .A1(n29462), .A2(n29459), .ZN(n29472) );
  NAND2_X1 U20522 ( .A1(n804), .A2(n12301), .ZN(n10938) );
  XNOR2_X1 U20523 ( .A(n488), .B(n593), .ZN(n21680) );
  OAI211_X1 U20524 ( .C1(n8565), .C2(n49605), .A(n49606), .B(n45720), .ZN(
        n8564) );
  INV_X1 U20525 ( .A(n49605), .ZN(n49554) );
  NOR2_X1 U20527 ( .A1(n45719), .A2(n49580), .ZN(n8565) );
  NAND2_X1 U20528 ( .A1(n13509), .A2(n13530), .ZN(n12932) );
  AND2_X2 U20529 ( .A1(n9300), .A2(n8566), .ZN(n13526) );
  NAND2_X1 U20530 ( .A1(n9298), .A2(n9299), .ZN(n8567) );
  NAND2_X1 U20531 ( .A1(n45614), .A2(n48456), .ZN(n8570) );
  XNOR2_X2 U20532 ( .A(n42432), .B(n42431), .ZN(n46444) );
  XNOR2_X1 U20534 ( .A(n17879), .B(n16628), .ZN(n8571) );
  XNOR2_X1 U20535 ( .A(n16720), .B(n8571), .ZN(n16400) );
  NAND2_X1 U20536 ( .A1(n18223), .A2(n19793), .ZN(n8573) );
  XNOR2_X1 U20537 ( .A(n44911), .B(n43000), .ZN(n41298) );
  NAND3_X2 U20538 ( .A1(n8583), .A2(n41297), .A3(n41296), .ZN(n44911) );
  OAI22_X1 U20539 ( .A1(n10775), .A2(n14160), .B1(n14150), .B2(n13122), .ZN(
        n8584) );
  NAND2_X1 U20540 ( .A1(n46441), .A2(n46449), .ZN(n46443) );
  XNOR2_X1 U20541 ( .A(n25220), .B(n24971), .ZN(n24984) );
  NAND2_X1 U20542 ( .A1(n14323), .A2(n8587), .ZN(n14324) );
  NAND3_X1 U20543 ( .A1(n14321), .A2(n14322), .A3(n14320), .ZN(n8587) );
  NAND2_X1 U20544 ( .A1(n8589), .A2(n20466), .ZN(n8588) );
  NAND2_X1 U20545 ( .A1(n20476), .A2(n20471), .ZN(n8593) );
  AND2_X1 U20546 ( .A1(n20481), .A2(n20482), .ZN(n8594) );
  NAND2_X1 U20548 ( .A1(n8597), .A2(n40910), .ZN(n40271) );
  NAND3_X1 U20549 ( .A1(n8599), .A2(n26733), .A3(n2420), .ZN(n8598) );
  INV_X1 U20550 ( .A(n8600), .ZN(n8599) );
  OAI21_X1 U20551 ( .B1(n24674), .B2(n51679), .A(n26989), .ZN(n8600) );
  INV_X1 U20552 ( .A(n50128), .ZN(n8603) );
  OAI211_X1 U20553 ( .C1(n50116), .C2(n50142), .A(n50099), .B(n8602), .ZN(
        n50100) );
  NAND2_X1 U20555 ( .A1(n12324), .A2(n9667), .ZN(n12341) );
  NAND2_X1 U20556 ( .A1(n17565), .A2(n17566), .ZN(n8604) );
  NAND2_X1 U20557 ( .A1(n19398), .A2(n17576), .ZN(n17579) );
  NAND2_X1 U20558 ( .A1(n8606), .A2(n10723), .ZN(n9017) );
  NAND3_X1 U20560 ( .A1(n40340), .A2(n40327), .A3(n8608), .ZN(n8607) );
  OR2_X1 U20561 ( .A1(n39855), .A2(n39857), .ZN(n39644) );
  XNOR2_X1 U20562 ( .A(n33359), .B(n8609), .ZN(n8611) );
  NOR2_X1 U20564 ( .A1(n13598), .A2(n14320), .ZN(n8612) );
  NAND2_X1 U20565 ( .A1(n8614), .A2(n8613), .ZN(n40431) );
  NAND2_X1 U20566 ( .A1(n41280), .A2(n41025), .ZN(n8614) );
  NAND2_X1 U20567 ( .A1(n50632), .A2(n50633), .ZN(n50635) );
  NAND4_X1 U20569 ( .A1(n20952), .A2(n22154), .A3(n21027), .A4(n8617), .ZN(
        n21920) );
  NOR2_X1 U20570 ( .A1(n22144), .A2(n21026), .ZN(n8617) );
  NAND2_X1 U20572 ( .A1(n38035), .A2(n35155), .ZN(n34207) );
  XNOR2_X1 U20573 ( .A(n43763), .B(n43775), .ZN(n8620) );
  XNOR2_X2 U20574 ( .A(n46095), .B(n8620), .ZN(n43798) );
  INV_X1 U20575 ( .A(n20094), .ZN(n8624) );
  NAND2_X1 U20577 ( .A1(n10101), .A2(n10109), .ZN(n10526) );
  XNOR2_X2 U20578 ( .A(n8626), .B(Key[89]), .ZN(n10109) );
  NAND2_X1 U20579 ( .A1(n26619), .A2(n28155), .ZN(n28529) );
  NAND2_X1 U20580 ( .A1(n47138), .A2(n47137), .ZN(n8628) );
  NAND2_X1 U20581 ( .A1(n22491), .A2(n20298), .ZN(n22837) );
  NAND3_X1 U20583 ( .A1(n18249), .A2(n18248), .A3(n8631), .ZN(n8630) );
  NAND2_X1 U20584 ( .A1(n19632), .A2(n19885), .ZN(n8631) );
  NAND2_X1 U20585 ( .A1(n39378), .A2(n39367), .ZN(n38966) );
  NOR2_X1 U20587 ( .A1(n37881), .A2(n37790), .ZN(n39378) );
  NAND2_X1 U20588 ( .A1(n31600), .A2(n32907), .ZN(n8634) );
  NAND2_X1 U20589 ( .A1(n31601), .A2(n32547), .ZN(n8635) );
  INV_X1 U20590 ( .A(n37034), .ZN(n37168) );
  INV_X1 U20592 ( .A(n30346), .ZN(n29061) );
  INV_X1 U20594 ( .A(n14643), .ZN(n9162) );
  INV_X1 U20595 ( .A(n30788), .ZN(n8640) );
  OAI22_X1 U20596 ( .A1(n20375), .A2(n20408), .B1(n1860), .B2(n20805), .ZN(
        n20409) );
  NAND2_X1 U20597 ( .A1(n8642), .A2(n21388), .ZN(n21390) );
  NAND2_X1 U20598 ( .A1(n20805), .A2(n5923), .ZN(n8642) );
  INV_X1 U20599 ( .A(n41110), .ZN(n39598) );
  INV_X1 U20600 ( .A(n46626), .ZN(n8645) );
  XNOR2_X2 U20601 ( .A(n8647), .B(n25699), .ZN(n29462) );
  XNOR2_X1 U20602 ( .A(n24517), .B(n2401), .ZN(n8647) );
  XNOR2_X1 U20605 ( .A(n34860), .B(n34849), .ZN(n8650) );
  NAND2_X1 U20606 ( .A1(n8652), .A2(n10391), .ZN(n8651) );
  NAND3_X1 U20607 ( .A1(n8654), .A2(n9431), .A3(n9244), .ZN(n8652) );
  OR2_X1 U20608 ( .A1(n11402), .A2(n11407), .ZN(n8654) );
  INV_X1 U20609 ( .A(n46996), .ZN(n47162) );
  INV_X1 U20610 ( .A(n43687), .ZN(n8655) );
  OR2_X2 U20611 ( .A1(n8655), .A2(n46996), .ZN(n47154) );
  XNOR2_X1 U20612 ( .A(n26548), .B(n8657), .ZN(n27481) );
  XNOR2_X1 U20613 ( .A(n26372), .B(n8657), .ZN(n26373) );
  XNOR2_X1 U20614 ( .A(n8657), .B(n27234), .ZN(n25962) );
  INV_X1 U20615 ( .A(n14831), .ZN(n8661) );
  NAND4_X1 U20616 ( .A1(n8660), .A2(n8662), .A3(n15433), .A4(n8659), .ZN(n8658) );
  NAND2_X1 U20617 ( .A1(n15444), .A2(n15437), .ZN(n8659) );
  NAND2_X1 U20618 ( .A1(n8661), .A2(n15437), .ZN(n8660) );
  NAND3_X1 U20619 ( .A1(n15326), .A2(n15437), .A3(n15431), .ZN(n8662) );
  NAND2_X1 U20621 ( .A1(n8390), .A2(n32175), .ZN(n32763) );
  AND2_X1 U20622 ( .A1(n11895), .A2(n510), .ZN(n11894) );
  NAND2_X1 U20623 ( .A1(n11894), .A2(n12474), .ZN(n8664) );
  NAND3_X1 U20624 ( .A1(n11896), .A2(n12488), .A3(n11895), .ZN(n8665) );
  NAND2_X1 U20625 ( .A1(n11908), .A2(n12486), .ZN(n8666) );
  INV_X1 U20626 ( .A(n11066), .ZN(n8667) );
  XNOR2_X1 U20627 ( .A(n18427), .B(n8670), .ZN(n16140) );
  XNOR2_X1 U20628 ( .A(n17936), .B(n8670), .ZN(n16469) );
  XNOR2_X1 U20629 ( .A(n17803), .B(n8670), .ZN(n16238) );
  XNOR2_X1 U20630 ( .A(n13985), .B(n8670), .ZN(n15511) );
  XNOR2_X1 U20631 ( .A(n18582), .B(n8670), .ZN(n18648) );
  NAND2_X1 U20632 ( .A1(n22991), .A2(n2477), .ZN(n8674) );
  NAND2_X1 U20633 ( .A1(n39376), .A2(n39375), .ZN(n39384) );
  NAND2_X1 U20634 ( .A1(n725), .A2(n29992), .ZN(n31140) );
  NAND2_X1 U20636 ( .A1(n29655), .A2(n31899), .ZN(n29989) );
  OR2_X1 U20637 ( .A1(n29655), .A2(n31899), .ZN(n8677) );
  XNOR2_X1 U20638 ( .A(n8678), .B(n36993), .ZN(n37004) );
  XNOR2_X1 U20639 ( .A(n37002), .B(n37126), .ZN(n8678) );
  AOI21_X1 U20640 ( .B1(n51137), .B2(n8796), .A(n8795), .ZN(n8679) );
  NAND2_X1 U20641 ( .A1(n12364), .A2(n8679), .ZN(n9025) );
  NOR2_X1 U20642 ( .A1(n32895), .A2(n8681), .ZN(n8682) );
  AND2_X1 U20643 ( .A1(n6270), .A2(n8682), .ZN(n32898) );
  NAND2_X1 U20644 ( .A1(n50578), .A2(n50641), .ZN(n44113) );
  XNOR2_X1 U20646 ( .A(n17225), .B(n17226), .ZN(n8683) );
  NAND2_X1 U20647 ( .A1(n15552), .A2(n8688), .ZN(n15558) );
  NOR3_X1 U20648 ( .A1(n48100), .A2(n48112), .A3(n8689), .ZN(n8690) );
  NAND4_X1 U20651 ( .A1(n38218), .A2(n35175), .A3(n38558), .A4(n51738), .ZN(
        n38220) );
  OR2_X1 U20652 ( .A1(n47745), .A2(n47763), .ZN(n47792) );
  AND2_X1 U20653 ( .A1(n46637), .A2(n46635), .ZN(n44868) );
  OR2_X1 U20654 ( .A1(n39449), .A2(n39448), .ZN(n39457) );
  INV_X1 U20655 ( .A(n49105), .ZN(n49106) );
  NAND4_X1 U20657 ( .A1(n48447), .A2(n48446), .A3(n48445), .A4(n48444), .ZN(
        n48567) );
  AND2_X1 U20658 ( .A1(n47874), .A2(n47803), .ZN(n47804) );
  OR2_X1 U20659 ( .A1(n50935), .A2(n50950), .ZN(n47389) );
  NOR2_X1 U20660 ( .A1(n47689), .A2(n47686), .ZN(n45859) );
  NAND4_X1 U20661 ( .A1(n38463), .A2(n38462), .A3(n38461), .A4(n38460), .ZN(
        n41820) );
  AND3_X1 U20662 ( .A1(n49544), .A2(n49543), .A3(n49542), .ZN(n49545) );
  NAND4_X2 U20663 ( .A1(n40891), .A2(n40889), .A3(n40888), .A4(n40890), .ZN(
        n44237) );
  OR2_X1 U20664 ( .A1(n37653), .A2(n37632), .ZN(n35739) );
  OAI21_X1 U20666 ( .B1(n45871), .B2(n45870), .A(n52149), .ZN(n45882) );
  INV_X1 U20667 ( .A(n47528), .ZN(n47579) );
  NAND4_X2 U20668 ( .A1(n40930), .A2(n40927), .A3(n40928), .A4(n40929), .ZN(
        n44030) );
  NAND4_X2 U20669 ( .A1(n40914), .A2(n40915), .A3(n40913), .A4(n40912), .ZN(
        n43619) );
  NOR2_X1 U20670 ( .A1(n44113), .A2(n50638), .ZN(n50575) );
  NAND4_X2 U20671 ( .A1(n49634), .A2(n49633), .A3(n49632), .A4(n49631), .ZN(
        n49853) );
  OR2_X1 U20672 ( .A1(n40357), .A2(n41342), .ZN(n39892) );
  INV_X1 U20674 ( .A(n50784), .ZN(n50773) );
  AND3_X1 U20676 ( .A1(n36230), .A2(n36229), .A3(n36228), .ZN(n36238) );
  NAND4_X1 U20677 ( .A1(n47365), .A2(n47364), .A3(n47363), .A4(n47362), .ZN(
        n47381) );
  AND2_X1 U20678 ( .A1(n43493), .A2(n49543), .ZN(n43494) );
  AND2_X1 U20679 ( .A1(n40277), .A2(n40276), .ZN(n40278) );
  NAND4_X2 U20680 ( .A1(n41295), .A2(n39123), .A3(n39122), .A4(n39124), .ZN(
        n42961) );
  INV_X1 U20681 ( .A(n47785), .ZN(n47787) );
  OR2_X1 U20682 ( .A1(n50387), .A2(n47315), .ZN(n47320) );
  INV_X1 U20683 ( .A(n47928), .ZN(n47986) );
  NAND4_X2 U20685 ( .A1(n50355), .A2(n50356), .A3(n50354), .A4(n50353), .ZN(
        n50452) );
  XNOR2_X2 U20686 ( .A(n42734), .B(n37354), .ZN(n48273) );
  XNOR2_X1 U20687 ( .A(n51525), .B(n43682), .ZN(n43687) );
  OR2_X1 U20688 ( .A1(n39902), .A2(n37356), .ZN(n39560) );
  XNOR2_X2 U20689 ( .A(n43209), .B(n41518), .ZN(n45099) );
  NAND4_X2 U20690 ( .A1(n41517), .A2(n41516), .A3(n41515), .A4(n41514), .ZN(
        n43209) );
  OAI211_X2 U20691 ( .C1(n39460), .C2(n39041), .A(n39040), .B(n39039), .ZN(
        n41691) );
  OR2_X1 U20692 ( .A1(n46772), .A2(n51304), .ZN(n45173) );
  XNOR2_X1 U20693 ( .A(n43379), .B(n43149), .ZN(n43162) );
  NAND4_X2 U20694 ( .A1(n36324), .A2(n36323), .A3(n36633), .A4(n36322), .ZN(
        n41435) );
  NAND4_X4 U20696 ( .A1(n44468), .A2(n44467), .A3(n44466), .A4(n44465), .ZN(
        n50721) );
  CLKBUF_X1 U20697 ( .A(n34629), .Z(n36414) );
  OAI211_X2 U20698 ( .C1(n14881), .C2(n14880), .A(n14879), .B(n15416), .ZN(
        n17213) );
  OR2_X1 U20699 ( .A1(n48521), .A2(n48518), .ZN(n45563) );
  OR2_X1 U20700 ( .A1(n22434), .A2(n22983), .ZN(n22436) );
  NAND4_X2 U20701 ( .A1(n12747), .A2(n12746), .A3(n12745), .A4(n12744), .ZN(
        n18438) );
  OAI222_X1 U20702 ( .A1(n50542), .A2(n50554), .B1(n50520), .B2(n50534), .C1(
        n47051), .C2(n50490), .ZN(n47052) );
  XNOR2_X1 U20703 ( .A(n27372), .B(n24703), .ZN(n24704) );
  NOR2_X1 U20704 ( .A1(n40972), .A2(n41380), .ZN(n40958) );
  NAND4_X2 U20705 ( .A1(n29965), .A2(n29964), .A3(n29963), .A4(n29962), .ZN(
        n37325) );
  NAND4_X2 U20706 ( .A1(n31128), .A2(n31127), .A3(n31126), .A4(n31125), .ZN(
        n34163) );
  AND2_X1 U20707 ( .A1(n14863), .A2(n15438), .ZN(n8697) );
  AND3_X1 U20708 ( .A1(n11279), .A2(n9973), .A3(n11276), .ZN(n8698) );
  NAND3_X1 U20709 ( .A1(n11729), .A2(n11728), .A3(n11727), .ZN(n8699) );
  XOR2_X1 U20710 ( .A(n52180), .B(n16458), .Z(n8700) );
  OR2_X1 U20711 ( .A1(n13143), .A2(n13142), .ZN(n8701) );
  OR2_X1 U20712 ( .A1(n13298), .A2(n13306), .ZN(n8702) );
  AND4_X1 U20713 ( .A1(n17482), .A2(n17483), .A3(n17481), .A4(n17480), .ZN(
        n8703) );
  AND2_X1 U20714 ( .A1(n51374), .A2(n19425), .ZN(n8704) );
  AND2_X1 U20715 ( .A1(n51432), .A2(n12619), .ZN(n8705) );
  AND2_X1 U20716 ( .A1(n19675), .A2(n19671), .ZN(n8707) );
  AND2_X1 U20717 ( .A1(n40893), .A2(n40901), .ZN(n8708) );
  AND2_X1 U20718 ( .A1(n14220), .A2(n13964), .ZN(n8709) );
  OR2_X1 U20720 ( .A1(n31622), .A2(n31584), .ZN(n8713) );
  AND2_X1 U20721 ( .A1(n28192), .A2(n28191), .ZN(n8714) );
  XOR2_X1 U20722 ( .A(n18430), .B(n18429), .Z(n8715) );
  AND4_X1 U20723 ( .A1(n15168), .A2(n15179), .A3(n15167), .A4(n15177), .ZN(
        n8716) );
  OR2_X1 U20724 ( .A1(n17486), .A2(n17485), .ZN(n8717) );
  AND2_X1 U20725 ( .A1(n12620), .A2(n10462), .ZN(n8718) );
  OR2_X1 U20726 ( .A1(n2089), .A2(n37782), .ZN(n8719) );
  OR2_X1 U20727 ( .A1(n39702), .A2(n38366), .ZN(n8721) );
  INV_X1 U20728 ( .A(n4121), .ZN(n42452) );
  OR2_X1 U20729 ( .A1(n12351), .A2(n12350), .ZN(n8724) );
  AND2_X1 U20730 ( .A1(n11707), .A2(n11704), .ZN(n8725) );
  AND3_X1 U20731 ( .A1(n11653), .A2(n11652), .A3(n11651), .ZN(n8726) );
  AND4_X1 U20732 ( .A1(n21397), .A2(n20789), .A3(n20790), .A4(n21369), .ZN(
        n8727) );
  XOR2_X1 U20733 ( .A(n14624), .B(n14623), .Z(n8728) );
  XOR2_X1 U20734 ( .A(n16605), .B(n16604), .Z(n8729) );
  AND2_X1 U20735 ( .A1(n23247), .A2(n23257), .ZN(n8730) );
  XOR2_X1 U20736 ( .A(n16430), .B(n16429), .Z(n8731) );
  XOR2_X1 U20737 ( .A(n23523), .B(n27325), .Z(n8733) );
  XOR2_X1 U20738 ( .A(n26453), .B(n26452), .Z(n8734) );
  AND2_X1 U20739 ( .A1(n29536), .A2(n29535), .ZN(n8735) );
  OR2_X1 U20740 ( .A1(n29461), .A2(n29456), .ZN(n8739) );
  NAND2_X1 U20741 ( .A1(n29505), .A2(n29504), .ZN(n8740) );
  AND3_X1 U20742 ( .A1(n32580), .A2(n32581), .A3(n32579), .ZN(n8741) );
  OR2_X1 U20743 ( .A1(n29013), .A2(n28926), .ZN(n8742) );
  AND2_X1 U20745 ( .A1(n2143), .A2(n30458), .ZN(n8747) );
  XOR2_X1 U20746 ( .A(n33619), .B(n34264), .Z(n8748) );
  AND2_X1 U20747 ( .A1(n30410), .A2(n30409), .ZN(n8750) );
  XOR2_X1 U20748 ( .A(n34606), .B(n36817), .Z(n8751) );
  NAND2_X1 U20749 ( .A1(n36218), .A2(n36214), .ZN(n8753) );
  AND3_X1 U20750 ( .A1(n39894), .A2(n39893), .A3(n39892), .ZN(n8755) );
  AND2_X1 U20751 ( .A1(n41231), .A2(n41228), .ZN(n8756) );
  XOR2_X1 U20752 ( .A(n41882), .B(n44170), .Z(n8757) );
  OR2_X1 U20753 ( .A1(n41481), .A2(n480), .ZN(n8758) );
  AND2_X1 U20754 ( .A1(n39767), .A2(n41433), .ZN(n8759) );
  XOR2_X1 U20755 ( .A(n41906), .B(n46082), .Z(n8760) );
  XOR2_X1 U20756 ( .A(n43322), .B(n41129), .Z(n8762) );
  AND4_X1 U20757 ( .A1(n50285), .A2(n50284), .A3(n50283), .A4(n50282), .ZN(
        n8763) );
  AND3_X1 U20758 ( .A1(n50548), .A2(n50550), .A3(n50552), .ZN(n8764) );
  OR2_X1 U20759 ( .A1(n45987), .A2(n49717), .ZN(n8765) );
  AND4_X1 U20760 ( .A1(n47102), .A2(n47101), .A3(n47100), .A4(n47099), .ZN(
        n8766) );
  AND2_X1 U20761 ( .A1(n45198), .A2(n50910), .ZN(n8767) );
  AND3_X1 U20762 ( .A1(n49125), .A2(n49124), .A3(n49102), .ZN(n8768) );
  AND2_X1 U20763 ( .A1(n42196), .A2(n47872), .ZN(n8769) );
  OR2_X1 U20764 ( .A1(n10633), .A2(n9482), .ZN(n10507) );
  OR2_X1 U20765 ( .A1(n51004), .A2(n12333), .ZN(n12326) );
  XNOR2_X1 U20766 ( .A(n9197), .B(Key[54]), .ZN(n9204) );
  INV_X1 U20767 ( .A(Ciphertext[155]), .ZN(n8785) );
  AND2_X1 U20768 ( .A1(n9057), .A2(n12314), .ZN(n12310) );
  OR2_X1 U20769 ( .A1(n9915), .A2(n9476), .ZN(n9918) );
  BUF_X1 U20771 ( .A(n8839), .Z(n10142) );
  OR2_X1 U20772 ( .A1(n12286), .A2(n10724), .ZN(n9700) );
  INV_X1 U20773 ( .A(n12310), .ZN(n9652) );
  INV_X1 U20774 ( .A(n10251), .ZN(n10201) );
  BUF_X1 U20776 ( .A(n8773), .Z(n10250) );
  OR3_X1 U20777 ( .A1(n10667), .A2(n10288), .A3(n51004), .ZN(n10278) );
  OR3_X1 U20778 ( .A1(n12674), .A2(n11875), .A3(n11884), .ZN(n11876) );
  NOR2_X1 U20779 ( .A1(n12620), .A2(n8705), .ZN(n12621) );
  XNOR2_X1 U20780 ( .A(Key[78]), .B(Ciphertext[191]), .ZN(n9407) );
  INV_X1 U20781 ( .A(n9417), .ZN(n8987) );
  XNOR2_X1 U20782 ( .A(Key[170]), .B(Ciphertext[67]), .ZN(n9153) );
  INV_X1 U20783 ( .A(n10695), .ZN(n10368) );
  INV_X1 U20784 ( .A(n12144), .ZN(n11417) );
  AND2_X1 U20785 ( .A1(n9981), .A2(n10589), .ZN(n11671) );
  AND2_X1 U20786 ( .A1(n10863), .A2(n12557), .ZN(n11519) );
  INV_X1 U20787 ( .A(n13430), .ZN(n13431) );
  INV_X1 U20788 ( .A(n9280), .ZN(n11612) );
  NOR2_X1 U20789 ( .A1(n11676), .A2(n8698), .ZN(n9979) );
  INV_X1 U20790 ( .A(n9700), .ZN(n9703) );
  AND2_X1 U20791 ( .A1(n10418), .A2(n11329), .ZN(n12151) );
  INV_X1 U20792 ( .A(n11620), .ZN(n10852) );
  AND2_X1 U20793 ( .A1(n10018), .A2(n11639), .ZN(n9508) );
  AOI211_X1 U20794 ( .C1(n9936), .C2(n11216), .A(n9935), .B(n8725), .ZN(n9937)
         );
  NOR2_X1 U20795 ( .A1(n14703), .A2(n14720), .ZN(n13742) );
  INV_X1 U20796 ( .A(n14199), .ZN(n14701) );
  INV_X1 U20797 ( .A(n12031), .ZN(n12028) );
  NAND4_X1 U20798 ( .A1(n10461), .A2(n10460), .A3(n10459), .A4(n10458), .ZN(
        n10499) );
  NAND4_X1 U20799 ( .A1(n11143), .A2(n11142), .A3(n11141), .A4(n11140), .ZN(
        n11144) );
  AND2_X1 U20800 ( .A1(n14484), .A2(n787), .ZN(n15372) );
  OR2_X1 U20801 ( .A1(n11715), .A2(n9146), .ZN(n9150) );
  AND2_X1 U20803 ( .A1(n10817), .A2(n11600), .ZN(n10818) );
  INV_X1 U20804 ( .A(n10719), .ZN(n9717) );
  NAND4_X1 U20805 ( .A1(n9664), .A2(n9663), .A3(n9662), .A4(n9661), .ZN(n9721)
         );
  INV_X1 U20806 ( .A(n13965), .ZN(n13966) );
  OR2_X1 U20807 ( .A1(n13082), .A2(n13091), .ZN(n13083) );
  OAI21_X1 U20808 ( .B1(n14036), .B2(n8702), .A(n12406), .ZN(n12407) );
  INV_X1 U20812 ( .A(n15334), .ZN(n14827) );
  NAND4_X1 U20813 ( .A1(n12646), .A2(n12645), .A3(n12644), .A4(n12643), .ZN(
        n12740) );
  NOR2_X1 U20814 ( .A1(n14473), .A2(n13856), .ZN(n13560) );
  INV_X1 U20815 ( .A(n15199), .ZN(n15242) );
  INV_X1 U20816 ( .A(n13628), .ZN(n9437) );
  INV_X1 U20817 ( .A(n18175), .ZN(n15640) );
  XNOR2_X1 U20818 ( .A(n15153), .B(n4487), .ZN(n15155) );
  NOR3_X1 U20819 ( .A1(n8709), .A2(n13967), .A3(n13966), .ZN(n16223) );
  AND2_X1 U20820 ( .A1(n13144), .A2(n8701), .ZN(n13156) );
  AND2_X1 U20821 ( .A1(n12853), .A2(n14439), .ZN(n12859) );
  INV_X1 U20822 ( .A(n13385), .ZN(n13035) );
  INV_X1 U20824 ( .A(n15034), .ZN(n15048) );
  INV_X1 U20825 ( .A(n16711), .ZN(n18448) );
  XNOR2_X1 U20826 ( .A(n18394), .B(n18393), .ZN(n18395) );
  XNOR2_X1 U20827 ( .A(n18437), .B(n15155), .ZN(n16593) );
  INV_X1 U20828 ( .A(n13033), .ZN(n13044) );
  AND2_X1 U20829 ( .A1(n13322), .A2(n14612), .ZN(n14003) );
  XNOR2_X1 U20830 ( .A(n15593), .B(n18546), .ZN(n15594) );
  INV_X1 U20831 ( .A(n19404), .ZN(n19405) );
  NAND4_X1 U20832 ( .A1(n15348), .A2(n15347), .A3(n15346), .A4(n15345), .ZN(
        n16201) );
  XNOR2_X1 U20833 ( .A(n16765), .B(n15990), .ZN(n14699) );
  XNOR2_X1 U20834 ( .A(n15594), .B(n15595), .ZN(n15599) );
  XNOR2_X1 U20835 ( .A(n15272), .B(n15271), .ZN(n15398) );
  XNOR2_X1 U20836 ( .A(n17910), .B(n17909), .ZN(n17911) );
  OR2_X1 U20838 ( .A1(n574), .A2(n20132), .ZN(n16808) );
  OR2_X1 U20839 ( .A1(n21361), .A2(n21359), .ZN(n18684) );
  OR2_X1 U20840 ( .A1(n18327), .A2(n18326), .ZN(n18328) );
  XNOR2_X1 U20841 ( .A(n16545), .B(n16544), .ZN(n16546) );
  XNOR2_X1 U20842 ( .A(n18632), .B(n18631), .ZN(n18635) );
  INV_X1 U20844 ( .A(n18903), .ZN(n18899) );
  AND3_X1 U20845 ( .A1(n21243), .A2(n21249), .A3(n17083), .ZN(n18968) );
  INV_X1 U20846 ( .A(n19675), .ZN(n19688) );
  INV_X1 U20847 ( .A(n18232), .ZN(n19674) );
  OR2_X1 U20848 ( .A1(n19793), .A2(n19801), .ZN(n18219) );
  INV_X1 U20849 ( .A(n20792), .ZN(n21370) );
  XNOR2_X1 U20850 ( .A(n18589), .B(n18588), .ZN(n18610) );
  INV_X1 U20851 ( .A(n20063), .ZN(n19136) );
  XNOR2_X1 U20852 ( .A(n17842), .B(n18568), .ZN(n17851) );
  XNOR2_X1 U20853 ( .A(n15709), .B(n15710), .ZN(n15723) );
  XNOR2_X1 U20854 ( .A(n18719), .B(n18718), .ZN(n18726) );
  NAND2_X1 U20855 ( .A1(n19418), .A2(n19412), .ZN(n15402) );
  XNOR2_X1 U20856 ( .A(n11183), .B(n18604), .ZN(n16392) );
  XNOR2_X1 U20857 ( .A(n15985), .B(n15984), .ZN(n15997) );
  XNOR2_X1 U20859 ( .A(n15574), .B(n15575), .ZN(n15631) );
  NAND4_X1 U20860 ( .A1(n20220), .A2(n19672), .A3(n19671), .A4(n51006), .ZN(
        n20214) );
  INV_X1 U20861 ( .A(n19377), .ZN(n14740) );
  XNOR2_X1 U20862 ( .A(n15320), .B(n15319), .ZN(n15399) );
  OR2_X1 U20863 ( .A1(n18963), .A2(n18962), .ZN(n19097) );
  XNOR2_X1 U20864 ( .A(n17373), .B(n17372), .ZN(n17405) );
  OR2_X1 U20865 ( .A1(n19837), .A2(n21185), .ZN(n19838) );
  BUF_X1 U20866 ( .A(n19966), .Z(n21483) );
  INV_X1 U20867 ( .A(n20072), .ZN(n19491) );
  OR2_X1 U20868 ( .A1(n20316), .A2(n21468), .ZN(n17747) );
  OAI21_X1 U20869 ( .B1(n20208), .B2(n18239), .A(n18238), .ZN(n18240) );
  AND3_X1 U20870 ( .A1(n20703), .A2(n20702), .A3(n20701), .ZN(n20704) );
  INV_X1 U20871 ( .A(n21836), .ZN(n21838) );
  NOR2_X1 U20872 ( .A1(n8727), .A2(n20793), .ZN(n20804) );
  AOI21_X1 U20873 ( .B1(n20483), .B2(n14741), .A(n14740), .ZN(n14748) );
  AND2_X1 U20874 ( .A1(n21218), .A2(n19807), .ZN(n18114) );
  AOI21_X1 U20875 ( .B1(n19130), .B2(n19129), .A(n19128), .ZN(n19149) );
  XNOR2_X1 U20876 ( .A(n15741), .B(n15740), .ZN(n15742) );
  OR2_X1 U20877 ( .A1(n23763), .A2(n2210), .ZN(n23193) );
  NOR2_X1 U20878 ( .A1(n22363), .A2(n22918), .ZN(n22368) );
  NAND4_X1 U20880 ( .A1(n20154), .A2(n20153), .A3(n20152), .A4(n20151), .ZN(
        n20161) );
  OR2_X1 U20881 ( .A1(n21196), .A2(n21214), .ZN(n19808) );
  OR2_X1 U20882 ( .A1(n23763), .A2(n24187), .ZN(n22606) );
  INV_X1 U20883 ( .A(n22994), .ZN(n22997) );
  INV_X1 U20884 ( .A(n22368), .ZN(n21040) );
  INV_X1 U20885 ( .A(n22920), .ZN(n22899) );
  NAND4_X1 U20886 ( .A1(n21241), .A2(n21240), .A3(n21239), .A4(n21238), .ZN(
        n22061) );
  OAI21_X1 U20887 ( .B1(n19811), .B2(n19810), .A(n19809), .ZN(n19825) );
  INV_X1 U20888 ( .A(n21723), .ZN(n20311) );
  NAND4_X1 U20889 ( .A1(n20756), .A2(n20755), .A3(n20754), .A4(n20753), .ZN(
        n20787) );
  AND2_X1 U20890 ( .A1(n23535), .A2(n23374), .ZN(n24324) );
  AND4_X1 U20891 ( .A1(n21573), .A2(n21572), .A3(n21571), .A4(n21570), .ZN(
        n21589) );
  INV_X1 U20892 ( .A(n22436), .ZN(n19758) );
  AND2_X1 U20893 ( .A1(n24194), .A2(n24193), .ZN(n24195) );
  INV_X1 U20894 ( .A(n22175), .ZN(n21717) );
  INV_X1 U20895 ( .A(n22223), .ZN(n24254) );
  NOR2_X1 U20896 ( .A1(n23835), .A2(n24146), .ZN(n21801) );
  INV_X1 U20897 ( .A(n22555), .ZN(n22567) );
  AND2_X1 U20898 ( .A1(n21707), .A2(n20566), .ZN(n20569) );
  OR2_X1 U20900 ( .A1(n25057), .A2(n25056), .ZN(n22768) );
  OR2_X1 U20902 ( .A1(n23343), .A2(n21150), .ZN(n20870) );
  OR2_X1 U20903 ( .A1(n22768), .A2(n22213), .ZN(n22214) );
  INV_X1 U20904 ( .A(n22574), .ZN(n22581) );
  XNOR2_X1 U20905 ( .A(n25802), .B(n25801), .ZN(n25804) );
  XNOR2_X1 U20907 ( .A(n24382), .B(n24381), .ZN(n24451) );
  INV_X1 U20908 ( .A(n27806), .ZN(n27807) );
  INV_X1 U20909 ( .A(n25965), .ZN(n25966) );
  BUF_X1 U20910 ( .A(n25002), .Z(n25533) );
  XNOR2_X1 U20911 ( .A(n24490), .B(n24491), .ZN(n24563) );
  XNOR2_X1 U20912 ( .A(n23743), .B(n25103), .ZN(n23744) );
  XNOR2_X1 U20913 ( .A(n26271), .B(n26270), .ZN(n26288) );
  INV_X1 U20914 ( .A(n29881), .ZN(n28773) );
  INV_X1 U20915 ( .A(n29867), .ZN(n28745) );
  XNOR2_X1 U20916 ( .A(n23190), .B(n23189), .ZN(n23301) );
  XNOR2_X1 U20917 ( .A(n25392), .B(n25391), .ZN(n25393) );
  AND3_X1 U20919 ( .A1(n25202), .A2(n25201), .A3(n25200), .ZN(n25203) );
  XNOR2_X1 U20920 ( .A(n22696), .B(n27183), .ZN(n27158) );
  XNOR2_X1 U20921 ( .A(n27360), .B(n27359), .ZN(n28764) );
  INV_X1 U20923 ( .A(n27821), .ZN(n27809) );
  INV_X1 U20925 ( .A(n29063), .ZN(n29069) );
  OR2_X1 U20926 ( .A1(n27717), .A2(n29413), .ZN(n26732) );
  XNOR2_X1 U20927 ( .A(n24607), .B(n24606), .ZN(n24649) );
  INV_X1 U20928 ( .A(n31420), .ZN(n27868) );
  XNOR2_X1 U20929 ( .A(n26454), .B(n8734), .ZN(n26455) );
  AND2_X1 U20930 ( .A1(n29446), .A2(n2213), .ZN(n26643) );
  INV_X1 U20931 ( .A(n29332), .ZN(n28644) );
  AND2_X1 U20933 ( .A1(n28679), .A2(n28678), .ZN(n28680) );
  OAI21_X1 U20934 ( .B1(n29460), .B2(n24561), .A(n8739), .ZN(n26690) );
  AND2_X1 U20935 ( .A1(n28205), .A2(n28204), .ZN(n28206) );
  OAI21_X1 U20936 ( .B1(n28984), .B2(n29714), .A(n28983), .ZN(n28985) );
  INV_X1 U20937 ( .A(n29220), .ZN(n27919) );
  OR2_X1 U20938 ( .A1(n32726), .A2(n32725), .ZN(n32727) );
  INV_X1 U20939 ( .A(n29714), .ZN(n28175) );
  OR2_X1 U20940 ( .A1(n30365), .A2(n1121), .ZN(n29890) );
  INV_X1 U20941 ( .A(n31987), .ZN(n31192) );
  OR2_X1 U20942 ( .A1(n31443), .A2(n31454), .ZN(n31444) );
  OR2_X1 U20943 ( .A1(n32822), .A2(n32420), .ZN(n31402) );
  OR2_X1 U20944 ( .A1(n31236), .A2(n29372), .ZN(n29374) );
  NAND4_X1 U20945 ( .A1(n27003), .A2(n27002), .A3(n27001), .A4(n27000), .ZN(
        n27023) );
  INV_X1 U20946 ( .A(n30930), .ZN(n29642) );
  OR2_X1 U20947 ( .A1(n32429), .A2(n31249), .ZN(n31250) );
  INV_X1 U20948 ( .A(n27075), .ZN(n27064) );
  AOI21_X1 U20949 ( .B1(n28576), .B2(n29007), .A(n28575), .ZN(n28597) );
  AND3_X1 U20951 ( .A1(n30728), .A2(n30729), .A3(n30727), .ZN(n30730) );
  OR2_X1 U20953 ( .A1(n32923), .A2(n32922), .ZN(n32924) );
  INV_X1 U20954 ( .A(n32409), .ZN(n33154) );
  INV_X1 U20955 ( .A(n32684), .ZN(n30143) );
  NAND4_X1 U20956 ( .A1(n30158), .A2(n30157), .A3(n30156), .A4(n30155), .ZN(
        n31967) );
  INV_X1 U20957 ( .A(n32661), .ZN(n31182) );
  NAND4_X1 U20958 ( .A1(n32713), .A2(n32712), .A3(n32711), .A4(n32710), .ZN(
        n33419) );
  AND2_X1 U20959 ( .A1(n32065), .A2(n8711), .ZN(n32086) );
  OR2_X1 U20960 ( .A1(n32987), .A2(n32976), .ZN(n32978) );
  NAND4_X1 U20961 ( .A1(n31984), .A2(n31983), .A3(n31982), .A4(n31981), .ZN(
        n33703) );
  INV_X1 U20962 ( .A(n31645), .ZN(n32731) );
  AND2_X1 U20963 ( .A1(n32720), .A2(n29753), .ZN(n32714) );
  NAND4_X1 U20964 ( .A1(n32308), .A2(n32307), .A3(n32306), .A4(n32305), .ZN(
        n32952) );
  XNOR2_X1 U20965 ( .A(n35522), .B(n37065), .ZN(n35048) );
  INV_X1 U20968 ( .A(n35630), .ZN(n35078) );
  OR2_X1 U20970 ( .A1(n38270), .A2(n2123), .ZN(n35416) );
  XNOR2_X1 U20971 ( .A(n33135), .B(n33134), .ZN(n34210) );
  XNOR2_X1 U20972 ( .A(n35349), .B(n33727), .ZN(n33778) );
  XNOR2_X1 U20973 ( .A(n33304), .B(n33537), .ZN(n33305) );
  INV_X1 U20974 ( .A(n34528), .ZN(n38273) );
  XNOR2_X1 U20975 ( .A(n36677), .B(n36678), .ZN(n36679) );
  XNOR2_X1 U20976 ( .A(n34437), .B(n34438), .ZN(n34569) );
  XNOR2_X1 U20977 ( .A(n37311), .B(n37310), .ZN(n37312) );
  INV_X1 U20978 ( .A(n36269), .ZN(n33678) );
  OR2_X1 U20979 ( .A1(n38160), .A2(n37448), .ZN(n35695) );
  XNOR2_X1 U20980 ( .A(n36845), .B(n36846), .ZN(n36853) );
  OR2_X1 U20981 ( .A1(n34908), .A2(n39395), .ZN(n34909) );
  XNOR2_X1 U20982 ( .A(n35245), .B(n35244), .ZN(n35304) );
  INV_X1 U20983 ( .A(n33649), .ZN(n34676) );
  AND2_X1 U20984 ( .A1(n36325), .A2(n31621), .ZN(n36326) );
  INV_X1 U20985 ( .A(n36233), .ZN(n37586) );
  INV_X1 U20986 ( .A(n39182), .ZN(n38676) );
  XNOR2_X1 U20987 ( .A(n34600), .B(n34599), .ZN(n34629) );
  INV_X1 U20988 ( .A(n35230), .ZN(n34448) );
  OR2_X1 U20989 ( .A1(n37680), .A2(n38641), .ZN(n37683) );
  XNOR2_X1 U20990 ( .A(n37310), .B(n33305), .ZN(n33310) );
  INV_X1 U20993 ( .A(n37618), .ZN(n38277) );
  INV_X1 U20994 ( .A(n38494), .ZN(n37384) );
  INV_X1 U20995 ( .A(n34569), .ZN(n34583) );
  INV_X1 U20996 ( .A(n37405), .ZN(n33674) );
  AND2_X1 U20997 ( .A1(n37579), .A2(n35695), .ZN(n35696) );
  NOR2_X1 U20998 ( .A1(n40404), .A2(n40453), .ZN(n38373) );
  AND2_X1 U20999 ( .A1(n37368), .A2(n35453), .ZN(n35454) );
  XNOR2_X1 U21000 ( .A(n34828), .B(n34827), .ZN(n34908) );
  XNOR2_X1 U21001 ( .A(n31762), .B(n34522), .ZN(n35017) );
  NOR2_X1 U21002 ( .A1(n41004), .A2(n43323), .ZN(n38760) );
  INV_X1 U21003 ( .A(n37633), .ZN(n37648) );
  INV_X1 U21005 ( .A(n38093), .ZN(n36642) );
  AND2_X1 U21006 ( .A1(n34699), .A2(n39486), .ZN(n38979) );
  OR2_X1 U21007 ( .A1(n37751), .A2(n37762), .ZN(n35924) );
  INV_X1 U21008 ( .A(n38760), .ZN(n37604) );
  AND2_X1 U21009 ( .A1(n39361), .A2(n39195), .ZN(n39374) );
  OAI21_X1 U21010 ( .B1(n33782), .B2(n37590), .A(n37588), .ZN(n33786) );
  INV_X1 U21011 ( .A(n42044), .ZN(n42045) );
  OR2_X1 U21012 ( .A1(n681), .A2(n432), .ZN(n39527) );
  OR2_X1 U21013 ( .A1(n37153), .A2(n51496), .ZN(n37154) );
  OR2_X1 U21014 ( .A1(n39856), .A2(n39644), .ZN(n38848) );
  NAND4_X1 U21015 ( .A1(n37234), .A2(n37233), .A3(n37232), .A4(n37231), .ZN(
        n37345) );
  OR2_X1 U21016 ( .A1(n5060), .A2(n8752), .ZN(n36179) );
  AND2_X1 U21017 ( .A1(n2086), .A2(n36491), .ZN(n36498) );
  AOI21_X1 U21018 ( .B1(n39374), .B2(n39381), .A(n39373), .ZN(n39391) );
  AND3_X1 U21019 ( .A1(n36646), .A2(n36645), .A3(n36644), .ZN(n36647) );
  INV_X1 U21020 ( .A(n40231), .ZN(n40229) );
  AND2_X1 U21021 ( .A1(n35856), .A2(n35855), .ZN(n35859) );
  OR2_X1 U21022 ( .A1(n39220), .A2(n39233), .ZN(n39257) );
  AND2_X1 U21023 ( .A1(n8753), .A2(n33877), .ZN(n33878) );
  INV_X1 U21024 ( .A(n40287), .ZN(n40290) );
  INV_X1 U21025 ( .A(n40869), .ZN(n39962) );
  OR2_X1 U21026 ( .A1(n40570), .A2(n40569), .ZN(n40575) );
  INV_X1 U21027 ( .A(n41850), .ZN(n43225) );
  NOR2_X1 U21028 ( .A1(n38410), .A2(n39674), .ZN(n40690) );
  AND2_X1 U21029 ( .A1(n39906), .A2(n39912), .ZN(n39562) );
  INV_X1 U21030 ( .A(n41981), .ZN(n41982) );
  INV_X1 U21031 ( .A(n40830), .ZN(n40833) );
  OAI21_X1 U21032 ( .B1(n36392), .B2(n39157), .A(n39774), .ZN(n36393) );
  AND2_X1 U21033 ( .A1(n40867), .A2(n40866), .ZN(n40879) );
  INV_X1 U21034 ( .A(n41098), .ZN(n41983) );
  AND2_X1 U21035 ( .A1(n37360), .A2(n37361), .ZN(n37362) );
  INV_X1 U21037 ( .A(n43236), .ZN(n40814) );
  OR2_X1 U21038 ( .A1(n40738), .A2(n6469), .ZN(n39637) );
  OR2_X1 U21039 ( .A1(n39593), .A2(n40486), .ZN(n39596) );
  XNOR2_X1 U21040 ( .A(n46150), .B(n43111), .ZN(n43112) );
  OR2_X1 U21041 ( .A1(n39666), .A2(n39100), .ZN(n39107) );
  OR2_X1 U21042 ( .A1(n39965), .A2(n39964), .ZN(n39975) );
  XNOR2_X1 U21043 ( .A(n43344), .B(n44153), .ZN(n44964) );
  XNOR2_X1 U21044 ( .A(n51371), .B(n45258), .ZN(n44299) );
  XNOR2_X1 U21045 ( .A(n42665), .B(n42664), .ZN(n42667) );
  NOR2_X1 U21046 ( .A1(n46392), .A2(n46489), .ZN(n46393) );
  XNOR2_X1 U21047 ( .A(n42238), .B(n42237), .ZN(n42271) );
  XNOR2_X1 U21048 ( .A(n42667), .B(n42666), .ZN(n42673) );
  AND2_X1 U21049 ( .A1(n45589), .A2(n48259), .ZN(n48423) );
  NOR2_X1 U21050 ( .A1(n45828), .A2(n45827), .ZN(n44280) );
  XNOR2_X1 U21051 ( .A(n41907), .B(n8760), .ZN(n41912) );
  XNOR2_X1 U21053 ( .A(n45301), .B(n45302), .ZN(n45628) );
  XNOR2_X1 U21054 ( .A(n42970), .B(n42969), .ZN(n42971) );
  XNOR2_X1 U21055 ( .A(n42655), .B(n44532), .ZN(n42685) );
  INV_X1 U21056 ( .A(n45095), .ZN(n43366) );
  XNOR2_X1 U21057 ( .A(n42956), .B(n45439), .ZN(n45995) );
  XNOR2_X1 U21058 ( .A(n43160), .B(n43159), .ZN(n43161) );
  INV_X1 U21059 ( .A(n50387), .ZN(n47327) );
  XNOR2_X1 U21060 ( .A(n43932), .B(n43760), .ZN(n43761) );
  AND2_X1 U21061 ( .A1(n46971), .A2(n46984), .ZN(n46798) );
  OR2_X1 U21062 ( .A1(n46824), .A2(n47074), .ZN(n46812) );
  XNOR2_X1 U21064 ( .A(n42120), .B(n42119), .ZN(n42177) );
  XNOR2_X1 U21065 ( .A(n45476), .B(n45477), .ZN(n45495) );
  XNOR2_X1 U21066 ( .A(n42547), .B(n42546), .ZN(n42605) );
  XNOR2_X1 U21067 ( .A(n42830), .B(n44949), .ZN(n42883) );
  XNOR2_X1 U21068 ( .A(n42843), .B(n45136), .ZN(n43479) );
  XNOR2_X1 U21070 ( .A(n46096), .B(n46095), .ZN(n47013) );
  XNOR2_X1 U21071 ( .A(n45136), .B(n45135), .ZN(n46648) );
  XNOR2_X1 U21073 ( .A(n45473), .B(n43743), .ZN(n46978) );
  OR2_X1 U21075 ( .A1(n44998), .A2(n44997), .ZN(n44999) );
  OR2_X1 U21076 ( .A1(n45552), .A2(n48219), .ZN(n45553) );
  OR2_X1 U21077 ( .A1(n45548), .A2(n48204), .ZN(n48211) );
  OAI21_X1 U21078 ( .B1(n46351), .B2(n46350), .A(n46269), .ZN(n46365) );
  NOR2_X1 U21079 ( .A1(n42617), .A2(n42616), .ZN(n42810) );
  OAI211_X1 U21080 ( .C1(n45899), .C2(n45898), .A(n8765), .B(n45897), .ZN(
        n45906) );
  NOR2_X1 U21081 ( .A1(n49146), .A2(n49137), .ZN(n49142) );
  OR2_X1 U21082 ( .A1(n45922), .A2(n49231), .ZN(n49696) );
  AND3_X1 U21083 ( .A1(n49746), .A2(n49745), .A3(n49744), .ZN(n49747) );
  BUF_X1 U21084 ( .A(n46034), .Z(n50296) );
  INV_X1 U21085 ( .A(n47335), .ZN(n50266) );
  AND4_X1 U21086 ( .A1(n44616), .A2(n44615), .A3(n47294), .A4(n44614), .ZN(
        n44617) );
  AND4_X1 U21087 ( .A1(n45030), .A2(n46910), .A3(n45029), .A4(n45028), .ZN(
        n45038) );
  AND3_X1 U21088 ( .A1(n45174), .A2(n45175), .A3(n45173), .ZN(n45182) );
  OR2_X1 U21089 ( .A1(n48941), .A2(n51510), .ZN(n48942) );
  INV_X1 U21091 ( .A(n47786), .ZN(n47728) );
  INV_X1 U21092 ( .A(n48020), .ZN(n48054) );
  AND2_X1 U21093 ( .A1(n45554), .A2(n45553), .ZN(n45555) );
  OR2_X1 U21094 ( .A1(n48160), .A2(n48159), .ZN(n48161) );
  AND2_X1 U21096 ( .A1(n44803), .A2(n44802), .ZN(n44804) );
  NAND4_X1 U21097 ( .A1(n46171), .A2(n46172), .A3(n46170), .A4(n46169), .ZN(
        n46173) );
  NAND4_X1 U21098 ( .A1(n47299), .A2(n47298), .A3(n47297), .A4(n47296), .ZN(
        n47382) );
  NAND4_X1 U21100 ( .A1(n45038), .A2(n45037), .A3(n45036), .A4(n45035), .ZN(
        n45192) );
  AOI211_X1 U21101 ( .C1(n48730), .C2(n48751), .A(n48722), .B(n48734), .ZN(
        n46422) );
  INV_X1 U21103 ( .A(n49793), .ZN(n49844) );
  NOR2_X1 U21104 ( .A1(n50198), .A2(n50180), .ZN(n47385) );
  AND3_X1 U21105 ( .A1(n42194), .A2(n47834), .A3(n42193), .ZN(n42197) );
  AND2_X1 U21107 ( .A1(n44445), .A2(n44444), .ZN(n44446) );
  AND3_X1 U21108 ( .A1(n44438), .A2(n44437), .A3(n44436), .ZN(n44449) );
  AND3_X1 U21109 ( .A1(n44796), .A2(n44797), .A3(n44795), .ZN(n44808) );
  AND2_X1 U21111 ( .A1(n44627), .A2(n44626), .ZN(n44636) );
  NAND4_X1 U21112 ( .A1(n44449), .A2(n44448), .A3(n44447), .A4(n44446), .ZN(
        n44451) );
  INV_X1 U21113 ( .A(Ciphertext[145]), .ZN(n8770) );
  XNOR2_X1 U21114 ( .A(n8770), .B(Key[140]), .ZN(n8773) );
  INV_X1 U21115 ( .A(Ciphertext[148]), .ZN(n8771) );
  INV_X1 U21116 ( .A(Ciphertext[149]), .ZN(n8772) );
  XNOR2_X1 U21117 ( .A(Key[37]), .B(Ciphertext[144]), .ZN(n8775) );
  XNOR2_X1 U21119 ( .A(Key[51]), .B(Ciphertext[146]), .ZN(n10252) );
  INV_X1 U21120 ( .A(n10252), .ZN(n9744) );
  INV_X1 U21121 ( .A(n11004), .ZN(n9029) );
  INV_X1 U21122 ( .A(n10199), .ZN(n8776) );
  INV_X1 U21124 ( .A(n9026), .ZN(n9751) );
  NAND2_X1 U21125 ( .A1(n9030), .A2(n9748), .ZN(n8774) );
  OAI21_X1 U21126 ( .B1(n9751), .B2(n9748), .A(n8774), .ZN(n8780) );
  XOR2_X1 U21127 ( .A(Ciphertext[147]), .B(Ciphertext[144]), .Z(n8778) );
  XNOR2_X1 U21128 ( .A(n4613), .B(n4754), .ZN(n8777) );
  XNOR2_X1 U21129 ( .A(n8778), .B(n8777), .ZN(n9752) );
  INV_X1 U21130 ( .A(n9752), .ZN(n10194) );
  INV_X1 U21131 ( .A(n10245), .ZN(n9033) );
  NAND2_X1 U21133 ( .A1(n11003), .A2(n10192), .ZN(n8779) );
  OAI21_X1 U21137 ( .B1(n10240), .B2(n11015), .A(n10192), .ZN(n9750) );
  NAND3_X1 U21138 ( .A1(n8782), .A2(n9748), .A3(n9750), .ZN(n8783) );
  AND2_X1 U21139 ( .A1(n10252), .A2(n51762), .ZN(n11006) );
  MUX2_X1 U21140 ( .A(n8784), .B(n8783), .S(n11006), .Z(n13582) );
  INV_X1 U21141 ( .A(Ciphertext[152]), .ZN(n8786) );
  INV_X1 U21143 ( .A(n10268), .ZN(n10261) );
  AND2_X1 U21144 ( .A1(n9022), .A2(n10261), .ZN(n10992) );
  INV_X1 U21145 ( .A(n10992), .ZN(n8789) );
  NAND2_X1 U21146 ( .A1(n10268), .A2(n9786), .ZN(n12351) );
  NOR2_X1 U21147 ( .A1(n12351), .A2(n12356), .ZN(n9020) );
  INV_X1 U21148 ( .A(n9020), .ZN(n10982) );
  INV_X1 U21149 ( .A(Ciphertext[150]), .ZN(n8787) );
  XNOR2_X1 U21150 ( .A(Key[4]), .B(Ciphertext[153]), .ZN(n8795) );
  INV_X1 U21151 ( .A(Ciphertext[154]), .ZN(n8788) );
  XNOR2_X1 U21152 ( .A(n8788), .B(Key[107]), .ZN(n8790) );
  NAND2_X1 U21153 ( .A1(n8791), .A2(n10267), .ZN(n10981) );
  NAND2_X1 U21154 ( .A1(n12356), .A2(n8795), .ZN(n10986) );
  AOI22_X1 U21155 ( .A1(n8789), .A2(n10982), .B1(n10981), .B2(n10986), .ZN(
        n8794) );
  NAND2_X1 U21157 ( .A1(n10262), .A2(n9782), .ZN(n10990) );
  NOR2_X1 U21158 ( .A1(n10990), .A2(n8791), .ZN(n10258) );
  AND2_X1 U21159 ( .A1(n10268), .A2(n9022), .ZN(n10988) );
  NAND2_X1 U21160 ( .A1(n10988), .A2(n10262), .ZN(n8792) );
  OAI22_X1 U21163 ( .A1(n10258), .A2(n8792), .B1(n12363), .B2(n52008), .ZN(
        n8793) );
  INV_X1 U21164 ( .A(n12351), .ZN(n12358) );
  INV_X1 U21165 ( .A(n10990), .ZN(n12354) );
  NAND3_X1 U21166 ( .A1(n8796), .A2(n10268), .A3(n10272), .ZN(n8797) );
  INV_X1 U21167 ( .A(Ciphertext[132]), .ZN(n8799) );
  NAND2_X1 U21169 ( .A1(n10054), .A2(n10121), .ZN(n9851) );
  INV_X1 U21170 ( .A(Ciphertext[135]), .ZN(n8800) );
  INV_X1 U21171 ( .A(n8803), .ZN(n10961) );
  INV_X1 U21172 ( .A(Ciphertext[137]), .ZN(n8801) );
  NAND2_X1 U21173 ( .A1(n10955), .A2(n10968), .ZN(n8802) );
  AOI21_X1 U21174 ( .B1(n9851), .B2(n10956), .A(n8802), .ZN(n8806) );
  INV_X1 U21175 ( .A(n10955), .ZN(n9850) );
  INV_X1 U21176 ( .A(n10968), .ZN(n10052) );
  NAND3_X1 U21177 ( .A1(n10054), .A2(n9850), .A3(n10052), .ZN(n8804) );
  INV_X1 U21178 ( .A(n10954), .ZN(n10963) );
  NOR2_X1 U21179 ( .A1(n8806), .A2(n8805), .ZN(n8816) );
  NAND2_X1 U21180 ( .A1(n10956), .A2(n10052), .ZN(n10971) );
  INV_X1 U21181 ( .A(Ciphertext[134]), .ZN(n8807) );
  XNOR2_X1 U21182 ( .A(n8807), .B(Key[159]), .ZN(n9855) );
  INV_X1 U21183 ( .A(n9855), .ZN(n10124) );
  AND2_X1 U21184 ( .A1(n10968), .A2(n10124), .ZN(n10957) );
  INV_X1 U21185 ( .A(n10957), .ZN(n8808) );
  NAND3_X1 U21186 ( .A1(n10971), .A2(n10121), .A3(n8808), .ZN(n8810) );
  INV_X1 U21187 ( .A(n10964), .ZN(n8809) );
  MUX2_X1 U21188 ( .A(n9863), .B(n8810), .S(n8809), .Z(n8815) );
  NAND3_X1 U21189 ( .A1(n10960), .A2(n10122), .A3(n10955), .ZN(n8813) );
  NAND3_X1 U21190 ( .A1(n10964), .A2(n10122), .A3(n10970), .ZN(n8812) );
  INV_X1 U21191 ( .A(n9856), .ZN(n13233) );
  NAND3_X1 U21192 ( .A1(n10957), .A2(n13233), .A3(n10122), .ZN(n8811) );
  NAND2_X1 U21194 ( .A1(n12198), .A2(n13590), .ZN(n14289) );
  INV_X1 U21196 ( .A(Ciphertext[127]), .ZN(n8817) );
  XNOR2_X1 U21198 ( .A(Key[28]), .B(Ciphertext[129]), .ZN(n10004) );
  INV_X1 U21199 ( .A(n10004), .ZN(n10008) );
  INV_X1 U21200 ( .A(Ciphertext[126]), .ZN(n8819) );
  MUX2_X1 U21201 ( .A(n8820), .B(n10003), .S(n11035), .Z(n8831) );
  INV_X1 U21202 ( .A(Ciphertext[131]), .ZN(n8821) );
  INV_X1 U21203 ( .A(Ciphertext[128]), .ZN(n8822) );
  INV_X1 U21204 ( .A(n10579), .ZN(n8824) );
  NOR2_X1 U21205 ( .A1(n11023), .A2(n10578), .ZN(n8823) );
  NAND2_X1 U21206 ( .A1(n10162), .A2(n10579), .ZN(n11036) );
  INV_X1 U21207 ( .A(n11036), .ZN(n10000) );
  INV_X1 U21209 ( .A(n10169), .ZN(n10159) );
  NAND3_X1 U21210 ( .A1(n11032), .A2(n10159), .A3(n11037), .ZN(n8829) );
  NAND2_X1 U21211 ( .A1(n790), .A2(n8639), .ZN(n8827) );
  NAND2_X1 U21212 ( .A1(n8639), .A2(n10004), .ZN(n10581) );
  INV_X1 U21213 ( .A(n10581), .ZN(n8825) );
  NAND2_X1 U21214 ( .A1(n8825), .A2(n11027), .ZN(n8826) );
  NAND4_X1 U21215 ( .A1(n10170), .A2(n8827), .A3(n10575), .A4(n8826), .ZN(
        n8828) );
  NAND2_X1 U21216 ( .A1(n14280), .A2(n12204), .ZN(n14290) );
  OAI21_X1 U21218 ( .B1(n14290), .B2(n13583), .A(n14285), .ZN(n8862) );
  INV_X1 U21219 ( .A(Ciphertext[142]), .ZN(n8832) );
  INV_X1 U21220 ( .A(Ciphertext[139]), .ZN(n8833) );
  INV_X1 U21222 ( .A(Ciphertext[138]), .ZN(n8834) );
  INV_X1 U21223 ( .A(n10134), .ZN(n10924) );
  INV_X1 U21224 ( .A(n10919), .ZN(n8839) );
  NAND2_X1 U21225 ( .A1(n10142), .A2(n10925), .ZN(n8835) );
  NAND2_X1 U21226 ( .A1(n10914), .A2(n8835), .ZN(n8837) );
  INV_X1 U21227 ( .A(Ciphertext[140]), .ZN(n8836) );
  XNOR2_X1 U21228 ( .A(n8836), .B(Key[9]), .ZN(n10138) );
  INV_X1 U21229 ( .A(n10931), .ZN(n10217) );
  INV_X1 U21230 ( .A(n10148), .ZN(n9806) );
  INV_X1 U21231 ( .A(n10218), .ZN(n8838) );
  INV_X1 U21232 ( .A(n10138), .ZN(n10221) );
  NAND2_X1 U21233 ( .A1(n10148), .A2(n52188), .ZN(n10137) );
  NAND2_X1 U21234 ( .A1(n10137), .A2(n10147), .ZN(n10144) );
  INV_X1 U21235 ( .A(n10144), .ZN(n8841) );
  OAI21_X1 U21236 ( .B1(n10147), .B2(n10919), .A(n10143), .ZN(n8842) );
  NAND2_X1 U21237 ( .A1(n10932), .A2(n8842), .ZN(n8845) );
  OAI21_X1 U21238 ( .B1(n10921), .B2(n10142), .A(n10217), .ZN(n8843) );
  NAND3_X1 U21239 ( .A1(n8843), .A2(n10219), .A3(n10137), .ZN(n8844) );
  INV_X1 U21240 ( .A(n10526), .ZN(n10532) );
  XNOR2_X1 U21241 ( .A(Key[61]), .B(Ciphertext[120]), .ZN(n8849) );
  INV_X1 U21242 ( .A(Ciphertext[122]), .ZN(n8847) );
  NAND3_X1 U21243 ( .A1(n10532), .A2(n10529), .A3(n9482), .ZN(n9842) );
  INV_X1 U21244 ( .A(n10101), .ZN(n8853) );
  NAND2_X1 U21245 ( .A1(n10529), .A2(n10519), .ZN(n10097) );
  NAND2_X1 U21246 ( .A1(n9484), .A2(n10097), .ZN(n8848) );
  AND2_X1 U21247 ( .A1(n9842), .A2(n8848), .ZN(n8859) );
  INV_X1 U21248 ( .A(n10519), .ZN(n10525) );
  INV_X1 U21249 ( .A(n10508), .ZN(n9836) );
  AND2_X1 U21250 ( .A1(n10101), .A2(n10026), .ZN(n10509) );
  INV_X1 U21251 ( .A(n10509), .ZN(n10105) );
  OAI21_X1 U21252 ( .B1(n9836), .B2(n10105), .A(n10522), .ZN(n8852) );
  OAI21_X1 U21253 ( .B1(n10522), .B2(n10096), .A(n10514), .ZN(n8851) );
  NAND3_X1 U21254 ( .A1(n10508), .A2(n10514), .A3(n9482), .ZN(n8850) );
  NAND4_X1 U21255 ( .A1(n8852), .A2(n8851), .A3(n10633), .A4(n8850), .ZN(n8858) );
  NAND3_X1 U21256 ( .A1(n10109), .A2(n10525), .A3(n10101), .ZN(n8854) );
  OAI211_X1 U21257 ( .C1(n8853), .C2(n1210), .A(n10508), .B(n8854), .ZN(n8855)
         );
  NAND2_X1 U21258 ( .A1(n8855), .A2(n10520), .ZN(n8857) );
  NOR2_X1 U21259 ( .A1(n14287), .A2(n14294), .ZN(n14286) );
  NAND2_X1 U21260 ( .A1(n14286), .A2(n13590), .ZN(n8860) );
  NAND4_X1 U21263 ( .A1(n14285), .A2(n13588), .A3(n14287), .A4(n12204), .ZN(
        n13978) );
  NAND4_X1 U21265 ( .A1(n5411), .A2(n13573), .A3(n12204), .A4(n13583), .ZN(
        n8863) );
  AND2_X1 U21266 ( .A1(n13978), .A2(n8863), .ZN(n8865) );
  NAND2_X1 U21267 ( .A1(n13588), .A2(n12204), .ZN(n14288) );
  NAND2_X1 U21268 ( .A1(n14288), .A2(n784), .ZN(n8864) );
  AND2_X1 U21270 ( .A1(n14285), .A2(n13979), .ZN(n12197) );
  NAND2_X1 U21271 ( .A1(n13013), .A2(n13583), .ZN(n13018) );
  OAI211_X1 U21272 ( .C1(n12198), .C2(n14287), .A(n12197), .B(n13018), .ZN(
        n13982) );
  INV_X1 U21273 ( .A(Ciphertext[59]), .ZN(n8866) );
  INV_X1 U21274 ( .A(Ciphertext[57]), .ZN(n8867) );
  INV_X1 U21275 ( .A(n11900), .ZN(n11903) );
  NOR2_X1 U21276 ( .A1(n8667), .A2(n12483), .ZN(n8868) );
  XNOR2_X1 U21277 ( .A(Key[11]), .B(Ciphertext[58]), .ZN(n10790) );
  INV_X1 U21278 ( .A(n10790), .ZN(n12488) );
  OAI211_X1 U21279 ( .C1(n11894), .C2(n8868), .A(n12488), .B(n11065), .ZN(
        n8876) );
  XNOR2_X1 U21280 ( .A(Key[86]), .B(Ciphertext[55]), .ZN(n8871) );
  NOR2_X1 U21281 ( .A1(n11488), .A2(n2116), .ZN(n8869) );
  NAND2_X1 U21282 ( .A1(n11900), .A2(n11899), .ZN(n12486) );
  NAND2_X1 U21283 ( .A1(n800), .A2(n11903), .ZN(n12471) );
  INV_X1 U21284 ( .A(n12471), .ZN(n10791) );
  AOI22_X1 U21285 ( .A1(n8869), .A2(n12486), .B1(n10791), .B2(n12470), .ZN(
        n8875) );
  NOR2_X1 U21287 ( .A1(n12488), .A2(n12481), .ZN(n8870) );
  AND2_X1 U21288 ( .A1(n11485), .A2(n12470), .ZN(n12487) );
  AOI21_X1 U21289 ( .B1(n10791), .B2(n8870), .A(n12487), .ZN(n8874) );
  INV_X1 U21290 ( .A(n12475), .ZN(n11902) );
  NOR2_X1 U21291 ( .A1(n11485), .A2(n510), .ZN(n8872) );
  INV_X1 U21292 ( .A(n8871), .ZN(n11489) );
  OAI211_X1 U21293 ( .C1(n11902), .C2(n8872), .A(n11908), .B(n11065), .ZN(
        n8873) );
  INV_X1 U21294 ( .A(n13683), .ZN(n8976) );
  INV_X1 U21295 ( .A(Ciphertext[40]), .ZN(n8877) );
  XNOR2_X1 U21296 ( .A(n8877), .B(Key[77]), .ZN(n12725) );
  INV_X1 U21297 ( .A(n8880), .ZN(n11942) );
  INV_X1 U21298 ( .A(Ciphertext[41]), .ZN(n8878) );
  NAND2_X1 U21299 ( .A1(n11942), .A2(n12728), .ZN(n12722) );
  INV_X1 U21300 ( .A(Ciphertext[36]), .ZN(n8879) );
  XNOR2_X1 U21301 ( .A(n8879), .B(Key[49]), .ZN(n8886) );
  NAND3_X1 U21302 ( .A1(n11941), .A2(n8882), .A3(n12720), .ZN(n11950) );
  INV_X1 U21303 ( .A(n12725), .ZN(n11954) );
  AND2_X1 U21304 ( .A1(n11107), .A2(n11954), .ZN(n10422) );
  NAND2_X1 U21305 ( .A1(n10422), .A2(n11108), .ZN(n8883) );
  OAI211_X1 U21306 ( .C1(n11112), .C2(n12722), .A(n11950), .B(n8883), .ZN(
        n8884) );
  INV_X1 U21307 ( .A(n8884), .ZN(n8895) );
  INV_X1 U21308 ( .A(n8885), .ZN(n10428) );
  NAND2_X1 U21309 ( .A1(n10438), .A2(n10431), .ZN(n11951) );
  NAND2_X1 U21310 ( .A1(n11951), .A2(n12720), .ZN(n8889) );
  OR2_X1 U21311 ( .A1(n11108), .A2(n12728), .ZN(n10437) );
  INV_X1 U21313 ( .A(n8886), .ZN(n10423) );
  NAND2_X1 U21314 ( .A1(n10423), .A2(n8885), .ZN(n11957) );
  NAND3_X1 U21315 ( .A1(n10438), .A2(n11964), .A3(n11957), .ZN(n8887) );
  OAI21_X1 U21316 ( .B1(n10437), .B2(n11109), .A(n8887), .ZN(n8888) );
  NAND2_X1 U21317 ( .A1(n8889), .A2(n8888), .ZN(n8894) );
  NOR2_X1 U21318 ( .A1(n11107), .A2(n5484), .ZN(n8890) );
  INV_X1 U21319 ( .A(n12722), .ZN(n10439) );
  OAI21_X1 U21320 ( .B1(n10431), .B2(n8890), .A(n10439), .ZN(n8892) );
  AND2_X1 U21321 ( .A1(n12728), .A2(n12720), .ZN(n11956) );
  NAND3_X1 U21322 ( .A1(n10438), .A2(n11956), .A3(n11957), .ZN(n8891) );
  NAND3_X1 U21323 ( .A1(n11955), .A2(n11958), .A3(n11956), .ZN(n8893) );
  NOR2_X1 U21324 ( .A1(n8976), .A2(n14252), .ZN(n15118) );
  INV_X1 U21325 ( .A(n15118), .ZN(n8958) );
  INV_X1 U21326 ( .A(Ciphertext[51]), .ZN(n8896) );
  INV_X1 U21327 ( .A(Ciphertext[48]), .ZN(n8897) );
  INV_X1 U21328 ( .A(Ciphertext[53]), .ZN(n8898) );
  INV_X1 U21329 ( .A(Ciphertext[52]), .ZN(n8899) );
  INV_X1 U21330 ( .A(Ciphertext[49]), .ZN(n8900) );
  INV_X1 U21331 ( .A(n11501), .ZN(n11077) );
  AND2_X1 U21332 ( .A1(n8909), .A2(n12464), .ZN(n11869) );
  NAND2_X1 U21333 ( .A1(n11869), .A2(n12673), .ZN(n11499) );
  NAND3_X1 U21334 ( .A1(n12675), .A2(n12464), .A3(n592), .ZN(n11079) );
  OAI211_X1 U21335 ( .C1(n11890), .C2(n8901), .A(n11499), .B(n11079), .ZN(
        n8905) );
  AND2_X1 U21336 ( .A1(n12458), .A2(n11874), .ZN(n11498) );
  INV_X1 U21337 ( .A(n11498), .ZN(n8903) );
  INV_X1 U21338 ( .A(n11869), .ZN(n12667) );
  NAND2_X1 U21339 ( .A1(n11083), .A2(n12667), .ZN(n8902) );
  INV_X1 U21340 ( .A(n8901), .ZN(n11870) );
  OAI21_X1 U21341 ( .B1(n8903), .B2(n8902), .A(n12450), .ZN(n8904) );
  NOR2_X1 U21342 ( .A1(n8905), .A2(n8904), .ZN(n8911) );
  NAND2_X1 U21343 ( .A1(n12675), .A2(n11077), .ZN(n12679) );
  NAND4_X1 U21344 ( .A1(n11501), .A2(n8909), .A3(n12458), .A4(n12680), .ZN(
        n8906) );
  INV_X1 U21345 ( .A(n12454), .ZN(n12462) );
  NAND2_X1 U21346 ( .A1(n8907), .A2(n592), .ZN(n8910) );
  INV_X1 U21347 ( .A(Ciphertext[71]), .ZN(n8912) );
  INV_X1 U21348 ( .A(n8915), .ZN(n8918) );
  INV_X1 U21349 ( .A(Ciphertext[69]), .ZN(n8914) );
  XNOR2_X1 U21350 ( .A(n8914), .B(Key[184]), .ZN(n8916) );
  INV_X1 U21351 ( .A(n8916), .ZN(n12502) );
  INV_X1 U21352 ( .A(n11550), .ZN(n11258) );
  INV_X1 U21353 ( .A(n9153), .ZN(n12512) );
  NAND2_X1 U21354 ( .A1(n12514), .A2(n12512), .ZN(n12523) );
  NAND2_X1 U21355 ( .A1(n8915), .A2(n12523), .ZN(n8917) );
  OAI211_X1 U21356 ( .C1(n8918), .C2(n11258), .A(n8917), .B(n11539), .ZN(n8929) );
  NAND2_X1 U21357 ( .A1(n642), .A2(n51653), .ZN(n11548) );
  INV_X1 U21358 ( .A(n11548), .ZN(n8919) );
  OAI21_X1 U21359 ( .B1(n8919), .B2(n11539), .A(n12506), .ZN(n8920) );
  NAND2_X1 U21360 ( .A1(n8920), .A2(n11255), .ZN(n8921) );
  AND2_X1 U21361 ( .A1(n51709), .A2(n12512), .ZN(n12500) );
  NAND2_X1 U21362 ( .A1(n8921), .A2(n12500), .ZN(n8928) );
  AND2_X1 U21363 ( .A1(n10831), .A2(n12512), .ZN(n11537) );
  NAND3_X1 U21364 ( .A1(n11537), .A2(n51653), .A3(n12502), .ZN(n8925) );
  INV_X1 U21365 ( .A(n11538), .ZN(n8922) );
  NAND3_X1 U21366 ( .A1(n8922), .A2(n12502), .A3(n8024), .ZN(n8924) );
  NAND3_X1 U21367 ( .A1(n51709), .A2(n10831), .A3(n8024), .ZN(n8923) );
  AND3_X1 U21368 ( .A1(n8925), .A2(n8924), .A3(n8923), .ZN(n8926) );
  NAND2_X1 U21369 ( .A1(n15103), .A2(n14983), .ZN(n13026) );
  XNOR2_X1 U21370 ( .A(Key[142]), .B(Ciphertext[63]), .ZN(n11091) );
  INV_X1 U21371 ( .A(n11091), .ZN(n10781) );
  XNOR2_X1 U21372 ( .A(Key[25]), .B(Ciphertext[60]), .ZN(n8949) );
  INV_X1 U21373 ( .A(Ciphertext[65]), .ZN(n8930) );
  XNOR2_X1 U21376 ( .A(Key[128]), .B(Ciphertext[61]), .ZN(n8945) );
  INV_X1 U21377 ( .A(n8945), .ZN(n12536) );
  INV_X1 U21378 ( .A(Ciphertext[64]), .ZN(n8931) );
  INV_X1 U21379 ( .A(n12549), .ZN(n10782) );
  INV_X1 U21380 ( .A(Ciphertext[62]), .ZN(n8932) );
  XOR2_X1 U21381 ( .A(Ciphertext[63]), .B(Ciphertext[60]), .Z(n8934) );
  XNOR2_X1 U21382 ( .A(Key[25]), .B(Key[142]), .ZN(n8933) );
  XNOR2_X1 U21383 ( .A(n8934), .B(n8933), .ZN(n12543) );
  INV_X1 U21384 ( .A(n12542), .ZN(n8941) );
  NAND3_X1 U21385 ( .A1(n12543), .A2(n12541), .A3(n8941), .ZN(n8935) );
  OAI21_X1 U21386 ( .B1(n8936), .B2(n11096), .A(n8935), .ZN(n8940) );
  AND2_X1 U21387 ( .A1(n8949), .A2(n11091), .ZN(n10780) );
  NAND3_X1 U21388 ( .A1(n12549), .A2(n12541), .A3(n10780), .ZN(n8938) );
  INV_X1 U21390 ( .A(n10780), .ZN(n9118) );
  NOR2_X1 U21392 ( .A1(n8940), .A2(n8939), .ZN(n8957) );
  INV_X1 U21393 ( .A(n11089), .ZN(n11100) );
  NAND2_X1 U21394 ( .A1(n11447), .A2(n9118), .ZN(n8944) );
  NOR2_X1 U21395 ( .A1(n11443), .A2(n11091), .ZN(n12547) );
  NAND2_X1 U21396 ( .A1(n12537), .A2(n6409), .ZN(n8950) );
  INV_X1 U21397 ( .A(n10778), .ZN(n9110) );
  OAI21_X1 U21398 ( .B1(n12547), .B2(n8950), .A(n9110), .ZN(n8942) );
  INV_X1 U21399 ( .A(n11449), .ZN(n8947) );
  INV_X1 U21400 ( .A(n11445), .ZN(n12533) );
  NOR2_X1 U21401 ( .A1(n12533), .A2(n10781), .ZN(n8946) );
  OAI21_X1 U21402 ( .B1(n8947), .B2(n8946), .A(n11447), .ZN(n8955) );
  OAI21_X1 U21403 ( .B1(n12533), .B2(n51673), .A(n8948), .ZN(n8953) );
  NOR2_X1 U21405 ( .A1(n12546), .A2(n12538), .ZN(n8952) );
  INV_X1 U21406 ( .A(n8950), .ZN(n8951) );
  OAI21_X1 U21407 ( .B1(n8953), .B2(n8952), .A(n8951), .ZN(n8954) );
  INV_X1 U21408 ( .A(n352), .ZN(n15117) );
  AOI21_X1 U21409 ( .B1(n8958), .B2(n13026), .A(n15117), .ZN(n14250) );
  INV_X1 U21410 ( .A(n15100), .ZN(n8974) );
  INV_X1 U21411 ( .A(Ciphertext[43]), .ZN(n8959) );
  XNOR2_X1 U21412 ( .A(n8959), .B(Key[2]), .ZN(n8961) );
  INV_X1 U21413 ( .A(Ciphertext[46]), .ZN(n8960) );
  AND2_X1 U21414 ( .A1(n12705), .A2(n8961), .ZN(n12441) );
  NAND2_X1 U21415 ( .A1(n12441), .A2(n12690), .ZN(n11928) );
  INV_X1 U21416 ( .A(n8961), .ZN(n11931) );
  INV_X1 U21417 ( .A(Ciphertext[45]), .ZN(n8962) );
  XNOR2_X1 U21418 ( .A(n8962), .B(Key[16]), .ZN(n8968) );
  NAND2_X1 U21419 ( .A1(n12696), .A2(n7780), .ZN(n8963) );
  INV_X1 U21420 ( .A(n8968), .ZN(n12695) );
  INV_X1 U21421 ( .A(Ciphertext[47]), .ZN(n8964) );
  AOI21_X1 U21422 ( .B1(n8965), .B2(n11937), .A(n2156), .ZN(n8973) );
  INV_X1 U21423 ( .A(Ciphertext[44]), .ZN(n8966) );
  OR2_X1 U21424 ( .A1(n8967), .A2(n12700), .ZN(n8972) );
  AND2_X1 U21425 ( .A1(n8968), .A2(n12690), .ZN(n12692) );
  AOI22_X1 U21426 ( .A1(n12696), .A2(n11125), .B1(n12692), .B2(n12435), .ZN(
        n8970) );
  INV_X1 U21427 ( .A(n12700), .ZN(n11933) );
  NAND2_X1 U21428 ( .A1(n10487), .A2(n11123), .ZN(n12703) );
  NAND2_X1 U21429 ( .A1(n11931), .A2(n11933), .ZN(n11122) );
  INV_X1 U21430 ( .A(n12440), .ZN(n12443) );
  OAI211_X1 U21431 ( .C1(n12696), .C2(n2156), .A(n11122), .B(n12443), .ZN(
        n8969) );
  OAI211_X1 U21432 ( .C1(n8970), .C2(n12711), .A(n12703), .B(n8969), .ZN(n8971) );
  INV_X1 U21433 ( .A(n14982), .ZN(n14251) );
  OAI211_X1 U21434 ( .C1(n14250), .C2(n8974), .A(n15106), .B(n14251), .ZN(
        n8982) );
  NAND2_X1 U21435 ( .A1(n352), .A2(n13683), .ZN(n14977) );
  NAND2_X1 U21436 ( .A1(n8975), .A2(n14984), .ZN(n8981) );
  OR2_X1 U21437 ( .A1(n14982), .A2(n15119), .ZN(n14245) );
  AND2_X1 U21438 ( .A1(n8976), .A2(n14252), .ZN(n14242) );
  NAND2_X1 U21439 ( .A1(n15118), .A2(n14983), .ZN(n8977) );
  INV_X1 U21440 ( .A(n8978), .ZN(n8980) );
  NOR2_X1 U21441 ( .A1(n14977), .A2(n8075), .ZN(n13022) );
  NAND2_X1 U21442 ( .A1(n13022), .A2(n780), .ZN(n8979) );
  INV_X1 U21443 ( .A(Ciphertext[178]), .ZN(n8983) );
  INV_X1 U21444 ( .A(Ciphertext[175]), .ZN(n8984) );
  INV_X1 U21445 ( .A(Ciphertext[174]), .ZN(n8985) );
  XNOR2_X1 U21446 ( .A(n8985), .B(Key[55]), .ZN(n8988) );
  INV_X1 U21447 ( .A(Ciphertext[177]), .ZN(n8986) );
  AND2_X1 U21448 ( .A1(n12266), .A2(n11341), .ZN(n12256) );
  INV_X1 U21449 ( .A(n12266), .ZN(n9419) );
  INV_X1 U21450 ( .A(n12258), .ZN(n12268) );
  INV_X1 U21451 ( .A(Ciphertext[179]), .ZN(n8989) );
  INV_X1 U21453 ( .A(Ciphertext[176]), .ZN(n8990) );
  XNOR2_X1 U21454 ( .A(n8990), .B(Key[69]), .ZN(n12255) );
  AND2_X1 U21455 ( .A1(n9647), .A2(n12255), .ZN(n12260) );
  NAND2_X1 U21456 ( .A1(n8994), .A2(n12242), .ZN(n10746) );
  AND2_X1 U21457 ( .A1(n12255), .A2(n12263), .ZN(n12269) );
  OAI211_X1 U21458 ( .C1(n11341), .C2(n10742), .A(n10746), .B(n12269), .ZN(
        n8991) );
  INV_X1 U21459 ( .A(n12260), .ZN(n10743) );
  NOR2_X1 U21460 ( .A1(n12256), .A2(n10743), .ZN(n8996) );
  NAND2_X1 U21461 ( .A1(n9417), .A2(n11341), .ZN(n10748) );
  INV_X1 U21462 ( .A(n12255), .ZN(n9425) );
  NAND2_X1 U21463 ( .A1(n12263), .A2(n9425), .ZN(n12246) );
  MUX2_X1 U21464 ( .A(n8996), .B(n8995), .S(n12267), .Z(n8997) );
  INV_X1 U21465 ( .A(Ciphertext[169]), .ZN(n8998) );
  INV_X1 U21466 ( .A(Ciphertext[172]), .ZN(n8999) );
  XNOR2_X1 U21467 ( .A(n8999), .B(Key[41]), .ZN(n9001) );
  INV_X1 U21468 ( .A(n9001), .ZN(n9698) );
  INV_X1 U21470 ( .A(Ciphertext[168]), .ZN(n9000) );
  INV_X1 U21471 ( .A(Ciphertext[170]), .ZN(n9002) );
  XNOR2_X1 U21472 ( .A(n9002), .B(Key[27]), .ZN(n9004) );
  INV_X1 U21473 ( .A(n9004), .ZN(n12294) );
  AND2_X1 U21475 ( .A1(n12278), .A2(n9015), .ZN(n9014) );
  INV_X1 U21476 ( .A(n9014), .ZN(n12290) );
  OAI21_X1 U21477 ( .B1(n12290), .B2(n12277), .A(n12291), .ZN(n9006) );
  NOR2_X1 U21478 ( .A1(n10234), .A2(n12294), .ZN(n9005) );
  OAI21_X1 U21479 ( .B1(n9006), .B2(n9005), .A(n10725), .ZN(n9012) );
  NAND3_X1 U21480 ( .A1(n9007), .A2(n10716), .A3(n9698), .ZN(n9009) );
  NAND3_X1 U21481 ( .A1(n12292), .A2(n10716), .A3(n4797), .ZN(n9008) );
  AND2_X1 U21482 ( .A1(n9009), .A2(n9008), .ZN(n9011) );
  NOR2_X1 U21483 ( .A1(n12276), .A2(n12277), .ZN(n10233) );
  NAND3_X1 U21484 ( .A1(n10233), .A2(n12292), .A3(n12291), .ZN(n9010) );
  OAI22_X1 U21486 ( .A1(n4797), .A2(n12286), .B1(n10715), .B2(n3445), .ZN(
        n9016) );
  NAND2_X1 U21487 ( .A1(n13820), .A2(n14311), .ZN(n13604) );
  AND2_X1 U21488 ( .A1(n8796), .A2(n805), .ZN(n9787) );
  INV_X1 U21489 ( .A(n10991), .ZN(n9024) );
  AND3_X1 U21490 ( .A1(n12350), .A2(n10267), .A3(n9022), .ZN(n9023) );
  NOR2_X1 U21491 ( .A1(n9780), .A2(n12352), .ZN(n12364) );
  INV_X1 U21492 ( .A(n12352), .ZN(n10976) );
  NOR2_X1 U21493 ( .A1(n13604), .A2(n13826), .ZN(n14303) );
  NAND3_X1 U21494 ( .A1(n11004), .A2(n7936), .A3(n10252), .ZN(n9747) );
  OAI21_X1 U21495 ( .B1(n9030), .B2(n9029), .A(n9028), .ZN(n10198) );
  NAND2_X1 U21496 ( .A1(n9031), .A2(n10195), .ZN(n10998) );
  NAND2_X1 U21497 ( .A1(n10198), .A2(n10998), .ZN(n9040) );
  NAND2_X1 U21498 ( .A1(n10251), .A2(n7936), .ZN(n9754) );
  INV_X1 U21499 ( .A(n9754), .ZN(n9035) );
  AOI21_X1 U21500 ( .B1(n9754), .B2(n9033), .A(n9032), .ZN(n9034) );
  OAI21_X1 U21501 ( .B1(n9752), .B2(n9035), .A(n9034), .ZN(n9039) );
  OAI21_X1 U21502 ( .B1(n11008), .B2(n10199), .A(n10240), .ZN(n9036) );
  AOI22_X1 U21503 ( .A1(n11004), .A2(n11001), .B1(n9037), .B2(n9036), .ZN(
        n9038) );
  NOR2_X1 U21504 ( .A1(n51064), .A2(n14311), .ZN(n13046) );
  INV_X1 U21505 ( .A(Ciphertext[167]), .ZN(n9042) );
  AND2_X1 U21506 ( .A1(n12340), .A2(n12325), .ZN(n10672) );
  NAND3_X1 U21507 ( .A1(n10672), .A2(n10288), .A3(n12338), .ZN(n10668) );
  INV_X1 U21508 ( .A(n9049), .ZN(n12323) );
  INV_X1 U21509 ( .A(Ciphertext[163]), .ZN(n9043) );
  XNOR2_X1 U21510 ( .A(n9043), .B(Key[74]), .ZN(n9045) );
  INV_X1 U21511 ( .A(n12340), .ZN(n12336) );
  NAND4_X1 U21512 ( .A1(n10673), .A2(n51462), .A3(n12336), .A4(n9044), .ZN(
        n9047) );
  INV_X1 U21513 ( .A(n9045), .ZN(n9668) );
  NAND2_X1 U21514 ( .A1(n9668), .A2(n9049), .ZN(n10279) );
  NAND3_X1 U21515 ( .A1(n10671), .A2(n51004), .A3(n12328), .ZN(n9046) );
  OAI211_X1 U21516 ( .C1(n10668), .C2(n12323), .A(n9047), .B(n9046), .ZN(n9053) );
  OAI21_X1 U21518 ( .B1(n12341), .B2(n9049), .A(n9048), .ZN(n9050) );
  NAND2_X1 U21519 ( .A1(n9050), .A2(n12340), .ZN(n9052) );
  OAI21_X1 U21520 ( .B1(n12332), .B2(n12340), .A(n9668), .ZN(n9051) );
  OR2_X1 U21521 ( .A1(n13046), .A2(n14317), .ZN(n13832) );
  INV_X1 U21522 ( .A(Ciphertext[157]), .ZN(n9054) );
  XNOR2_X1 U21523 ( .A(n9054), .B(Key[32]), .ZN(n9056) );
  INV_X1 U21524 ( .A(Ciphertext[159]), .ZN(n9055) );
  AND2_X1 U21525 ( .A1(n9057), .A2(n12315), .ZN(n10948) );
  AND2_X1 U21526 ( .A1(n12303), .A2(n12313), .ZN(n10940) );
  NAND2_X1 U21527 ( .A1(n10948), .A2(n10940), .ZN(n10950) );
  AND2_X1 U21528 ( .A1(n12313), .A2(n12314), .ZN(n9773) );
  NAND2_X1 U21529 ( .A1(n9772), .A2(n9773), .ZN(n9060) );
  INV_X1 U21530 ( .A(n10293), .ZN(n10947) );
  NAND3_X1 U21531 ( .A1(n10947), .A2(n12299), .A3(n10945), .ZN(n9059) );
  INV_X1 U21532 ( .A(n10948), .ZN(n10951) );
  NAND2_X1 U21533 ( .A1(n10296), .A2(n12313), .ZN(n9657) );
  NAND3_X1 U21534 ( .A1(n10951), .A2(n12314), .A3(n9657), .ZN(n9058) );
  NAND4_X1 U21535 ( .A1(n9060), .A2(n9059), .A3(n9058), .A4(n12301), .ZN(n9061) );
  NAND2_X1 U21536 ( .A1(n9656), .A2(n12313), .ZN(n9755) );
  OAI22_X1 U21537 ( .A1(n9755), .A2(n10939), .B1(n12303), .B2(n9762), .ZN(
        n9062) );
  NAND2_X1 U21538 ( .A1(n9062), .A2(n9767), .ZN(n9063) );
  NAND2_X1 U21539 ( .A1(n14307), .A2(n14317), .ZN(n13610) );
  OR3_X1 U21540 ( .A1(n11796), .A2(n14320), .A3(n13827), .ZN(n9065) );
  NAND2_X1 U21542 ( .A1(n14319), .A2(n14315), .ZN(n9064) );
  OAI211_X1 U21543 ( .C1(n13819), .C2(n13610), .A(n9065), .B(n9064), .ZN(n9066) );
  AOI21_X1 U21545 ( .B1(n14321), .B2(n9067), .A(n13045), .ZN(n9068) );
  NAND2_X1 U21546 ( .A1(n9068), .A2(n13599), .ZN(n9069) );
  INV_X1 U21548 ( .A(Ciphertext[84]), .ZN(n9071) );
  XNOR2_X1 U21549 ( .A(n9071), .B(Key[1]), .ZN(n9074) );
  XNOR2_X1 U21550 ( .A(Key[118]), .B(Ciphertext[87]), .ZN(n9073) );
  NOR2_X1 U21551 ( .A1(n3250), .A2(n11588), .ZN(n10810) );
  INV_X1 U21552 ( .A(Ciphertext[88]), .ZN(n9072) );
  NAND2_X1 U21553 ( .A1(n10810), .A2(n9279), .ZN(n11596) );
  NAND2_X1 U21555 ( .A1(n9083), .A2(n11590), .ZN(n11615) );
  INV_X1 U21556 ( .A(n9073), .ZN(n10816) );
  NOR2_X1 U21557 ( .A1(n11598), .A2(n10816), .ZN(n9896) );
  INV_X1 U21558 ( .A(n11615), .ZN(n10809) );
  NAND2_X1 U21559 ( .A1(n9896), .A2(n10809), .ZN(n9077) );
  NAND2_X1 U21560 ( .A1(n9278), .A2(n11590), .ZN(n11242) );
  INV_X1 U21561 ( .A(n11242), .ZN(n9075) );
  NAND3_X1 U21562 ( .A1(n9075), .A2(n11613), .A3(n10815), .ZN(n9076) );
  OAI211_X1 U21563 ( .C1(n11596), .C2(n11615), .A(n9077), .B(n9076), .ZN(n9082) );
  INV_X1 U21564 ( .A(n11604), .ZN(n9893) );
  AOI21_X1 U21566 ( .B1(n9893), .B2(n9083), .A(n11601), .ZN(n9080) );
  NAND3_X1 U21567 ( .A1(n11591), .A2(n10809), .A3(n11604), .ZN(n9079) );
  INV_X1 U21568 ( .A(n11598), .ZN(n9888) );
  NAND4_X1 U21569 ( .A1(n11592), .A2(n9888), .A3(n9895), .A4(n11590), .ZN(
        n9078) );
  XNOR2_X1 U21572 ( .A(Key[1]), .B(Key[118]), .ZN(n9085) );
  XNOR2_X1 U21573 ( .A(Ciphertext[84]), .B(Ciphertext[87]), .ZN(n9084) );
  XNOR2_X1 U21574 ( .A(n9085), .B(n9084), .ZN(n11250) );
  INV_X1 U21575 ( .A(n11250), .ZN(n10814) );
  NAND3_X1 U21576 ( .A1(n10814), .A2(n9280), .A3(n10815), .ZN(n9086) );
  AND2_X1 U21577 ( .A1(n10805), .A2(n9086), .ZN(n9092) );
  INV_X1 U21578 ( .A(n10806), .ZN(n9088) );
  NAND2_X1 U21580 ( .A1(n9279), .A2(n11604), .ZN(n9890) );
  OAI21_X1 U21581 ( .B1(n9088), .B2(n9087), .A(n9890), .ZN(n9091) );
  NAND2_X1 U21582 ( .A1(n11613), .A2(n11588), .ZN(n11610) );
  OAI211_X1 U21583 ( .C1(n11247), .C2(n10816), .A(n9089), .B(n9895), .ZN(n9090) );
  INV_X1 U21584 ( .A(Ciphertext[80]), .ZN(n9094) );
  XNOR2_X1 U21585 ( .A(Key[151]), .B(Ciphertext[78]), .ZN(n9103) );
  INV_X1 U21586 ( .A(Ciphertext[79]), .ZN(n9095) );
  OAI22_X1 U21587 ( .A1(n11633), .A2(n11470), .B1(n454), .B2(n11467), .ZN(
        n9096) );
  XNOR2_X1 U21588 ( .A(Key[179]), .B(Ciphertext[82]), .ZN(n9098) );
  NAND2_X1 U21589 ( .A1(n454), .A2(n11226), .ZN(n11224) );
  INV_X1 U21590 ( .A(n11634), .ZN(n11466) );
  AND2_X1 U21591 ( .A1(n11621), .A2(n11466), .ZN(n11631) );
  INV_X1 U21592 ( .A(Ciphertext[81]), .ZN(n9097) );
  INV_X1 U21593 ( .A(n9104), .ZN(n11624) );
  NAND4_X1 U21594 ( .A1(n11631), .A2(n11630), .A3(n11468), .A4(n11460), .ZN(
        n9101) );
  OAI21_X1 U21595 ( .B1(n11468), .B2(n11467), .A(n454), .ZN(n9099) );
  NAND2_X1 U21596 ( .A1(n11477), .A2(n9099), .ZN(n9100) );
  AND2_X2 U21598 ( .A1(n11468), .A2(n454), .ZN(n11620) );
  NAND2_X1 U21599 ( .A1(n11467), .A2(n11620), .ZN(n9323) );
  INV_X1 U21600 ( .A(n9323), .ZN(n10851) );
  NAND2_X1 U21601 ( .A1(n10851), .A2(n9102), .ZN(n9107) );
  NAND2_X1 U21602 ( .A1(n9104), .A2(n9103), .ZN(n11629) );
  NAND2_X1 U21603 ( .A1(n11629), .A2(n11224), .ZN(n11474) );
  INV_X1 U21604 ( .A(n11474), .ZN(n9105) );
  INV_X1 U21605 ( .A(n453), .ZN(n11229) );
  NAND3_X1 U21606 ( .A1(n9105), .A2(n51239), .A3(n11466), .ZN(n9106) );
  INV_X1 U21607 ( .A(n14635), .ZN(n9135) );
  NAND2_X1 U21608 ( .A1(n10786), .A2(n12543), .ZN(n9112) );
  NAND3_X1 U21609 ( .A1(n11446), .A2(n9109), .A3(n9110), .ZN(n9111) );
  NAND2_X1 U21610 ( .A1(n9112), .A2(n9111), .ZN(n9116) );
  MUX2_X1 U21611 ( .A(n12533), .B(n11089), .S(n12546), .Z(n9114) );
  INV_X1 U21612 ( .A(n10787), .ZN(n11092) );
  NAND3_X1 U21613 ( .A1(n11092), .A2(n9109), .A3(n442), .ZN(n9113) );
  NAND3_X1 U21614 ( .A1(n11446), .A2(n11445), .A3(n9118), .ZN(n11095) );
  INV_X1 U21617 ( .A(Ciphertext[72]), .ZN(n9122) );
  XNOR2_X1 U21618 ( .A(n9122), .B(Key[109]), .ZN(n9124) );
  INV_X1 U21619 ( .A(n9124), .ZN(n12573) );
  INV_X1 U21620 ( .A(Ciphertext[75]), .ZN(n9123) );
  XNOR2_X1 U21621 ( .A(n9123), .B(Key[34]), .ZN(n9129) );
  INV_X1 U21622 ( .A(n9129), .ZN(n11514) );
  NAND2_X1 U21623 ( .A1(n11566), .A2(n11567), .ZN(n9134) );
  NAND2_X1 U21624 ( .A1(n11582), .A2(n9129), .ZN(n11569) );
  NAND2_X1 U21625 ( .A1(n11569), .A2(n12555), .ZN(n12565) );
  NAND2_X1 U21626 ( .A1(n11582), .A2(n11514), .ZN(n11570) );
  NAND2_X1 U21627 ( .A1(n11570), .A2(n11581), .ZN(n9125) );
  OAI211_X1 U21628 ( .C1(n12565), .C2(n11567), .A(n12570), .B(n9125), .ZN(
        n9128) );
  INV_X1 U21629 ( .A(n11568), .ZN(n10863) );
  INV_X1 U21630 ( .A(n12556), .ZN(n9132) );
  INV_X1 U21631 ( .A(n11510), .ZN(n9131) );
  NAND2_X1 U21632 ( .A1(n11189), .A2(n12572), .ZN(n9130) );
  OR2_X1 U21633 ( .A1(n11570), .A2(n12574), .ZN(n11532) );
  INV_X1 U21634 ( .A(n11532), .ZN(n11193) );
  INV_X1 U21635 ( .A(n10859), .ZN(n10860) );
  NAND2_X1 U21636 ( .A1(n9132), .A2(n7340), .ZN(n12569) );
  OAI211_X1 U21637 ( .C1(n11193), .C2(n10860), .A(n51491), .B(n12569), .ZN(
        n9133) );
  NAND3_X1 U21638 ( .A1(n9135), .A2(n14633), .A3(n8121), .ZN(n9161) );
  XNOR2_X1 U21639 ( .A(Key[174]), .B(Ciphertext[95]), .ZN(n9148) );
  AND2_X1 U21640 ( .A1(n9491), .A2(n9926), .ZN(n11199) );
  INV_X1 U21641 ( .A(Ciphertext[93]), .ZN(n9136) );
  XNOR2_X1 U21642 ( .A(n9136), .B(Key[160]), .ZN(n9139) );
  INV_X1 U21643 ( .A(Ciphertext[90]), .ZN(n9137) );
  XNOR2_X1 U21644 ( .A(n9137), .B(Key[43]), .ZN(n9140) );
  INV_X1 U21646 ( .A(Ciphertext[94]), .ZN(n9138) );
  INV_X1 U21647 ( .A(n51649), .ZN(n9142) );
  INV_X1 U21648 ( .A(n9139), .ZN(n9495) );
  INV_X1 U21649 ( .A(Ciphertext[91]), .ZN(n9141) );
  XNOR2_X1 U21650 ( .A(n9141), .B(Key[146]), .ZN(n9147) );
  MUX2_X1 U21651 ( .A(n9143), .B(n11697), .S(n9500), .Z(n9152) );
  AND2_X1 U21652 ( .A1(n9144), .A2(n9932), .ZN(n9145) );
  AND2_X1 U21653 ( .A1(n643), .A2(n9491), .ZN(n11709) );
  OAI21_X1 U21654 ( .B1(n9145), .B2(n9499), .A(n11709), .ZN(n9151) );
  INV_X1 U21656 ( .A(n11707), .ZN(n9146) );
  INV_X1 U21657 ( .A(n11203), .ZN(n11212) );
  INV_X1 U21658 ( .A(n9147), .ZN(n11695) );
  OAI22_X1 U21659 ( .A1(n11212), .A2(n11210), .B1(n9146), .B2(n11209), .ZN(
        n9149) );
  AND2_X1 U21660 ( .A1(n11209), .A2(n9499), .ZN(n11198) );
  INV_X1 U21661 ( .A(n9500), .ZN(n11211) );
  AND2_X1 U21663 ( .A1(n643), .A2(n11705), .ZN(n11204) );
  NAND2_X1 U21664 ( .A1(n14644), .A2(n12756), .ZN(n12943) );
  NAND2_X1 U21665 ( .A1(n12943), .A2(n13669), .ZN(n9159) );
  OAI211_X1 U21666 ( .C1(n10832), .C2(n642), .A(n11258), .B(n11538), .ZN(n9155) );
  NAND2_X1 U21667 ( .A1(n51653), .A2(n9153), .ZN(n12498) );
  INV_X1 U21668 ( .A(n12498), .ZN(n10833) );
  NAND4_X1 U21669 ( .A1(n11550), .A2(n10833), .A3(n51709), .A4(n8024), .ZN(
        n9154) );
  AND2_X1 U21670 ( .A1(n9155), .A2(n9154), .ZN(n9158) );
  INV_X1 U21671 ( .A(n11537), .ZN(n10826) );
  INV_X1 U21672 ( .A(n11539), .ZN(n10836) );
  NAND2_X1 U21673 ( .A1(n10838), .A2(n10836), .ZN(n9156) );
  NAND4_X1 U21674 ( .A1(n9159), .A2(n9162), .A3(n13667), .A4(n13664), .ZN(
        n9160) );
  AND2_X1 U21675 ( .A1(n9161), .A2(n9160), .ZN(n14564) );
  AOI21_X1 U21676 ( .B1(n9162), .B2(n12756), .A(n14641), .ZN(n9165) );
  OAI21_X1 U21677 ( .B1(n9162), .B2(n12756), .A(n3254), .ZN(n9164) );
  OAI21_X1 U21678 ( .B1(n13659), .B2(n14642), .A(n14644), .ZN(n9163) );
  OAI21_X1 U21679 ( .B1(n9165), .B2(n9164), .A(n9163), .ZN(n14563) );
  NAND2_X1 U21680 ( .A1(n13669), .A2(n12755), .ZN(n9166) );
  NOR2_X1 U21681 ( .A1(n14632), .A2(n9166), .ZN(n14562) );
  NAND2_X1 U21682 ( .A1(n14562), .A2(n2114), .ZN(n9169) );
  INV_X1 U21683 ( .A(n12753), .ZN(n9167) );
  NAND2_X1 U21684 ( .A1(n14561), .A2(n2114), .ZN(n9168) );
  NAND4_X1 U21685 ( .A1(n14564), .A2(n14563), .A3(n9169), .A4(n9168), .ZN(
        n9170) );
  INV_X1 U21686 ( .A(Ciphertext[27]), .ZN(n9171) );
  XNOR2_X1 U21687 ( .A(n9171), .B(Key[82]), .ZN(n9178) );
  INV_X1 U21688 ( .A(n11986), .ZN(n9180) );
  INV_X1 U21689 ( .A(Ciphertext[29]), .ZN(n9172) );
  AOI21_X1 U21690 ( .B1(n9180), .B2(n10456), .A(n12659), .ZN(n9177) );
  INV_X1 U21691 ( .A(Ciphertext[25]), .ZN(n9173) );
  INV_X1 U21692 ( .A(Ciphertext[28]), .ZN(n9174) );
  AND2_X1 U21694 ( .A1(n11986), .A2(n10456), .ZN(n11982) );
  INV_X1 U21695 ( .A(n11982), .ZN(n9176) );
  AND2_X1 U21696 ( .A1(n11979), .A2(n797), .ZN(n11974) );
  INV_X1 U21697 ( .A(n11974), .ZN(n9175) );
  OAI22_X1 U21698 ( .A1(n9177), .A2(n11973), .B1(n9176), .B2(n9175), .ZN(n9185) );
  OAI211_X1 U21699 ( .C1(n12657), .C2(n11986), .A(n9179), .B(n10455), .ZN(
        n9184) );
  OAI21_X1 U21701 ( .B1(n794), .B2(n10449), .A(n9181), .ZN(n9182) );
  NAND2_X1 U21702 ( .A1(n9182), .A2(n11973), .ZN(n9183) );
  NOR2_X1 U21703 ( .A1(n2227), .A2(n11984), .ZN(n9187) );
  OAI21_X1 U21704 ( .B1(n10451), .B2(n9187), .A(n11979), .ZN(n9190) );
  NAND2_X1 U21705 ( .A1(n10456), .A2(n12648), .ZN(n9191) );
  NAND4_X1 U21706 ( .A1(n10457), .A2(n12660), .A3(n9188), .A4(n2227), .ZN(
        n9189) );
  NAND3_X1 U21707 ( .A1(n9190), .A2(n9191), .A3(n9189), .ZN(n9195) );
  INV_X1 U21708 ( .A(n9191), .ZN(n9192) );
  INV_X1 U21709 ( .A(Ciphertext[23]), .ZN(n9197) );
  INV_X1 U21710 ( .A(Ciphertext[20]), .ZN(n9198) );
  INV_X1 U21711 ( .A(n12635), .ZN(n12619) );
  INV_X1 U21712 ( .A(Ciphertext[22]), .ZN(n9199) );
  INV_X1 U21713 ( .A(n9203), .ZN(n12068) );
  NOR2_X1 U21714 ( .A1(n12637), .A2(n12068), .ZN(n9206) );
  INV_X1 U21715 ( .A(Ciphertext[21]), .ZN(n9200) );
  XNOR2_X1 U21716 ( .A(n9200), .B(Key[40]), .ZN(n9210) );
  AOI22_X1 U21717 ( .A1(n9206), .A2(n12069), .B1(n12628), .B2(n9201), .ZN(
        n9213) );
  INV_X1 U21718 ( .A(Ciphertext[19]), .ZN(n9202) );
  NAND2_X1 U21719 ( .A1(n9207), .A2(n9203), .ZN(n12071) );
  NOR2_X1 U21720 ( .A1(n12071), .A2(n10465), .ZN(n10464) );
  INV_X1 U21721 ( .A(n9204), .ZN(n9208) );
  OAI21_X1 U21722 ( .B1(n3347), .B2(n9208), .A(n12631), .ZN(n9205) );
  INV_X1 U21724 ( .A(n12616), .ZN(n10463) );
  INV_X1 U21725 ( .A(n9207), .ZN(n12066) );
  INV_X1 U21726 ( .A(n12620), .ZN(n9564) );
  NAND2_X1 U21727 ( .A1(n10465), .A2(n12066), .ZN(n9209) );
  OAI211_X1 U21728 ( .C1(n12069), .C2(n12618), .A(n9564), .B(n9209), .ZN(n9212) );
  INV_X1 U21729 ( .A(Ciphertext[0]), .ZN(n9214) );
  INV_X1 U21730 ( .A(n9380), .ZN(n12046) );
  INV_X1 U21731 ( .A(Ciphertext[4]), .ZN(n9215) );
  XNOR2_X2 U21732 ( .A(n9215), .B(Key[17]), .ZN(n11393) );
  XNOR2_X1 U21733 ( .A(Key[92]), .B(Ciphertext[1]), .ZN(n9384) );
  INV_X1 U21734 ( .A(n9384), .ZN(n10361) );
  AND2_X1 U21735 ( .A1(n11393), .A2(n10361), .ZN(n10354) );
  INV_X1 U21736 ( .A(n10354), .ZN(n11390) );
  NOR2_X1 U21737 ( .A1(n12046), .A2(n11390), .ZN(n9220) );
  INV_X1 U21738 ( .A(Ciphertext[5]), .ZN(n9216) );
  XNOR2_X1 U21739 ( .A(n9216), .B(Key[120]), .ZN(n9218) );
  INV_X1 U21740 ( .A(Ciphertext[2]), .ZN(n9217) );
  INV_X1 U21741 ( .A(n10360), .ZN(n9221) );
  INV_X1 U21742 ( .A(n11393), .ZN(n12052) );
  INV_X1 U21743 ( .A(n12045), .ZN(n12043) );
  NAND3_X1 U21744 ( .A1(n10362), .A2(n12057), .A3(n9221), .ZN(n9222) );
  AND2_X1 U21745 ( .A1(n9386), .A2(n9222), .ZN(n12050) );
  INV_X1 U21746 ( .A(n10362), .ZN(n12054) );
  INV_X1 U21747 ( .A(n10666), .ZN(n9224) );
  MUX2_X1 U21748 ( .A(n10362), .B(n10664), .S(n12051), .Z(n9223) );
  NOR2_X1 U21749 ( .A1(n9224), .A2(n9223), .ZN(n9228) );
  XOR2_X1 U21750 ( .A(Ciphertext[3]), .B(Ciphertext[0]), .Z(n9226) );
  XNOR2_X1 U21751 ( .A(Key[106]), .B(Key[181]), .ZN(n9225) );
  XNOR2_X1 U21752 ( .A(n9226), .B(n9225), .ZN(n12053) );
  NAND3_X1 U21753 ( .A1(n12053), .A2(n12047), .A3(n12045), .ZN(n9227) );
  INV_X1 U21754 ( .A(Ciphertext[13]), .ZN(n9229) );
  XNOR2_X1 U21755 ( .A(n9229), .B(Key[176]), .ZN(n9589) );
  INV_X1 U21756 ( .A(Ciphertext[16]), .ZN(n9230) );
  XNOR2_X1 U21757 ( .A(n9230), .B(Key[101]), .ZN(n10333) );
  AND2_X1 U21758 ( .A1(n9589), .A2(n10333), .ZN(n12160) );
  INV_X1 U21759 ( .A(Ciphertext[12]), .ZN(n9231) );
  XNOR2_X1 U21760 ( .A(Key[190]), .B(Ciphertext[15]), .ZN(n11329) );
  NAND2_X1 U21762 ( .A1(n12160), .A2(n10417), .ZN(n12153) );
  INV_X1 U21763 ( .A(n11328), .ZN(n11325) );
  INV_X1 U21764 ( .A(n9589), .ZN(n9235) );
  INV_X1 U21765 ( .A(n10333), .ZN(n12166) );
  NAND3_X1 U21766 ( .A1(n11325), .A2(n12171), .A3(n12169), .ZN(n9584) );
  INV_X1 U21768 ( .A(n11330), .ZN(n9232) );
  NAND3_X1 U21769 ( .A1(n9232), .A2(n11328), .A3(n12169), .ZN(n9233) );
  AND3_X1 U21770 ( .A1(n12153), .A2(n9584), .A3(n9233), .ZN(n9241) );
  NOR2_X1 U21771 ( .A1(n11324), .A2(n10413), .ZN(n12158) );
  OAI211_X1 U21772 ( .C1(n12158), .C2(n10418), .A(n548), .B(n12175), .ZN(n9240) );
  NAND2_X1 U21773 ( .A1(n10418), .A2(n9585), .ZN(n10412) );
  NAND2_X1 U21774 ( .A1(n12152), .A2(n10412), .ZN(n9236) );
  INV_X1 U21775 ( .A(n12178), .ZN(n9591) );
  NAND2_X1 U21777 ( .A1(n10413), .A2(n11329), .ZN(n12177) );
  INV_X1 U21778 ( .A(n12177), .ZN(n12174) );
  OAI211_X1 U21779 ( .C1(n9591), .C2(n10413), .A(n9238), .B(n9237), .ZN(n9239)
         );
  INV_X1 U21780 ( .A(n12133), .ZN(n12143) );
  INV_X1 U21781 ( .A(Ciphertext[6]), .ZN(n9242) );
  NAND2_X1 U21782 ( .A1(n12143), .A2(n12129), .ZN(n9252) );
  INV_X1 U21783 ( .A(Ciphertext[8]), .ZN(n9243) );
  INV_X1 U21785 ( .A(n11403), .ZN(n9605) );
  NAND2_X1 U21786 ( .A1(n51141), .A2(n9605), .ZN(n9604) );
  INV_X1 U21787 ( .A(n9604), .ZN(n11407) );
  NAND2_X1 U21788 ( .A1(n11410), .A2(n12139), .ZN(n9244) );
  INV_X1 U21789 ( .A(n12130), .ZN(n9431) );
  INV_X1 U21790 ( .A(Ciphertext[9]), .ZN(n9245) );
  INV_X1 U21791 ( .A(n9433), .ZN(n9598) );
  INV_X1 U21792 ( .A(n12141), .ZN(n10391) );
  NAND2_X1 U21793 ( .A1(n11410), .A2(n11411), .ZN(n12140) );
  INV_X1 U21794 ( .A(n12140), .ZN(n9247) );
  INV_X1 U21796 ( .A(n12137), .ZN(n10385) );
  AND2_X1 U21797 ( .A1(n11403), .A2(n51141), .ZN(n10392) );
  INV_X1 U21798 ( .A(n10392), .ZN(n9246) );
  AOI22_X1 U21799 ( .A1(n9247), .A2(n10385), .B1(n12130), .B2(n9246), .ZN(
        n9251) );
  NAND2_X1 U21800 ( .A1(n10398), .A2(n9433), .ZN(n12134) );
  INV_X1 U21801 ( .A(n12134), .ZN(n11408) );
  NOR2_X1 U21802 ( .A1(n11410), .A2(n9598), .ZN(n9248) );
  OAI21_X1 U21803 ( .B1(n11408), .B2(n9248), .A(n10383), .ZN(n9249) );
  OR2_X1 U21804 ( .A1(n15422), .A2(n13888), .ZN(n15412) );
  INV_X1 U21805 ( .A(Ciphertext[35]), .ZN(n9253) );
  AND2_X1 U21806 ( .A1(n12595), .A2(n9547), .ZN(n11920) );
  XNOR2_X1 U21808 ( .A(Key[124]), .B(Ciphertext[33]), .ZN(n11914) );
  INV_X1 U21810 ( .A(n12594), .ZN(n9258) );
  INV_X1 U21811 ( .A(Ciphertext[30]), .ZN(n9255) );
  INV_X1 U21812 ( .A(n11136), .ZN(n11921) );
  OAI21_X1 U21813 ( .B1(n10480), .B2(n11921), .A(n3377), .ZN(n9257) );
  NOR2_X1 U21814 ( .A1(n9548), .A2(n9539), .ZN(n9551) );
  INV_X1 U21815 ( .A(n9551), .ZN(n9256) );
  OAI211_X1 U21816 ( .C1(n51140), .C2(n9258), .A(n9257), .B(n9256), .ZN(n9266)
         );
  INV_X1 U21817 ( .A(n12589), .ZN(n12596) );
  NAND2_X1 U21818 ( .A1(n9542), .A2(n12596), .ZN(n11129) );
  NAND2_X1 U21819 ( .A1(n9537), .A2(n11129), .ZN(n9261) );
  NOR2_X1 U21820 ( .A1(n12601), .A2(n52140), .ZN(n9262) );
  NAND2_X1 U21821 ( .A1(n9262), .A2(n10480), .ZN(n9552) );
  NAND2_X1 U21822 ( .A1(n10474), .A2(n52140), .ZN(n12600) );
  AND2_X1 U21823 ( .A1(n9547), .A2(n11137), .ZN(n12592) );
  NAND2_X1 U21824 ( .A1(n9262), .A2(n12592), .ZN(n9260) );
  NAND4_X1 U21825 ( .A1(n9261), .A2(n9552), .A3(n11130), .A4(n9260), .ZN(n9265) );
  INV_X1 U21826 ( .A(n9262), .ZN(n11919) );
  NOR2_X1 U21827 ( .A1(n12597), .A2(n357), .ZN(n9264) );
  NAND2_X1 U21828 ( .A1(n50966), .A2(n13874), .ZN(n13261) );
  INV_X1 U21829 ( .A(n9267), .ZN(n9269) );
  OAI211_X1 U21830 ( .C1(n13875), .C2(n13874), .A(n9269), .B(n9268), .ZN(n9272) );
  OAI21_X1 U21831 ( .B1(n11613), .B2(n11590), .A(n9888), .ZN(n9276) );
  NAND2_X1 U21832 ( .A1(n11589), .A2(n10809), .ZN(n9275) );
  MUX2_X1 U21833 ( .A(n9276), .B(n9275), .S(n11588), .Z(n9285) );
  INV_X1 U21834 ( .A(n11593), .ZN(n11249) );
  INV_X1 U21835 ( .A(n11610), .ZN(n9277) );
  NAND2_X1 U21836 ( .A1(n11598), .A2(n11590), .ZN(n11614) );
  NAND2_X1 U21837 ( .A1(n9279), .A2(n3250), .ZN(n9283) );
  INV_X1 U21841 ( .A(Ciphertext[110]), .ZN(n9286) );
  INV_X1 U21842 ( .A(Ciphertext[113]), .ZN(n9287) );
  NAND2_X1 U21843 ( .A1(n10072), .A2(n10068), .ZN(n10070) );
  INV_X1 U21844 ( .A(Ciphertext[108]), .ZN(n9288) );
  XNOR2_X1 U21845 ( .A(Key[94]), .B(Ciphertext[111]), .ZN(n9289) );
  XNOR2_X1 U21847 ( .A(Key[5]), .B(Ciphertext[112]), .ZN(n9292) );
  INV_X1 U21848 ( .A(n9292), .ZN(n9476) );
  OAI211_X1 U21850 ( .C1(n10605), .C2(n10610), .A(n9908), .B(n10618), .ZN(
        n9290) );
  AND2_X1 U21851 ( .A1(n9290), .A2(n9873), .ZN(n9300) );
  AND2_X1 U21852 ( .A1(n10617), .A2(n10072), .ZN(n10609) );
  AND2_X1 U21853 ( .A1(n10072), .A2(n10065), .ZN(n10611) );
  INV_X1 U21854 ( .A(n10611), .ZN(n9297) );
  NAND2_X1 U21855 ( .A1(n10617), .A2(n9476), .ZN(n9874) );
  INV_X1 U21856 ( .A(n10072), .ZN(n9914) );
  OAI21_X1 U21857 ( .B1(n9915), .B2(n10070), .A(n10610), .ZN(n9294) );
  INV_X1 U21858 ( .A(n10616), .ZN(n9293) );
  NAND2_X1 U21859 ( .A1(n9294), .A2(n9293), .ZN(n9299) );
  NAND2_X1 U21860 ( .A1(n10072), .A2(n9476), .ZN(n9295) );
  OAI211_X1 U21861 ( .C1(n10064), .C2(n10074), .A(n9295), .B(n9297), .ZN(n9296) );
  OAI211_X1 U21862 ( .C1(n52185), .C2(n9297), .A(n9296), .B(n10617), .ZN(n9298) );
  INV_X1 U21863 ( .A(Ciphertext[106]), .ZN(n9301) );
  XNOR2_X1 U21864 ( .A(n9301), .B(Key[155]), .ZN(n9306) );
  INV_X1 U21866 ( .A(n11639), .ZN(n9510) );
  NAND2_X1 U21867 ( .A1(n9302), .A2(n10562), .ZN(n11650) );
  INV_X1 U21868 ( .A(Ciphertext[104]), .ZN(n9303) );
  XNOR2_X1 U21869 ( .A(n9303), .B(Key[141]), .ZN(n9308) );
  INV_X1 U21870 ( .A(Ciphertext[107]), .ZN(n9304) );
  INV_X1 U21872 ( .A(n11640), .ZN(n10572) );
  INV_X1 U21873 ( .A(n10562), .ZN(n9305) );
  INV_X1 U21874 ( .A(n9306), .ZN(n9939) );
  NAND3_X1 U21875 ( .A1(n10013), .A2(n11658), .A3(n11662), .ZN(n9311) );
  INV_X1 U21876 ( .A(n11644), .ZN(n9307) );
  NAND3_X1 U21877 ( .A1(n9307), .A2(n11654), .A3(n9317), .ZN(n9310) );
  NAND3_X1 U21878 ( .A1(n11649), .A2(n11658), .A3(n11641), .ZN(n9309) );
  INV_X1 U21879 ( .A(n11663), .ZN(n9944) );
  NAND2_X1 U21880 ( .A1(n11641), .A2(n3079), .ZN(n10570) );
  INV_X1 U21881 ( .A(n10570), .ZN(n9316) );
  AOI22_X1 U21882 ( .A1(n9318), .A2(n11648), .B1(n10563), .B2(n11658), .ZN(
        n9320) );
  NAND3_X1 U21884 ( .A1(n11464), .A2(n11461), .A3(n11460), .ZN(n9326) );
  AND2_X1 U21885 ( .A1(n9325), .A2(n9326), .ZN(n9330) );
  INV_X1 U21886 ( .A(n11234), .ZN(n11628) );
  NAND3_X1 U21887 ( .A1(n9327), .A2(n11631), .A3(n11460), .ZN(n9329) );
  NAND2_X1 U21888 ( .A1(n11635), .A2(n11224), .ZN(n9328) );
  NOR2_X1 U21889 ( .A1(n51682), .A2(n51066), .ZN(n10884) );
  INV_X1 U21890 ( .A(Ciphertext[96]), .ZN(n9331) );
  XNOR2_X1 U21891 ( .A(n9331), .B(Key[85]), .ZN(n9335) );
  INV_X1 U21892 ( .A(Ciphertext[99]), .ZN(n9332) );
  INV_X1 U21893 ( .A(Ciphertext[100]), .ZN(n9333) );
  XNOR2_X1 U21894 ( .A(n9333), .B(Key[113]), .ZN(n9519) );
  INV_X1 U21895 ( .A(n11276), .ZN(n10590) );
  INV_X1 U21896 ( .A(n11270), .ZN(n11679) );
  INV_X1 U21897 ( .A(Ciphertext[101]), .ZN(n9334) );
  XNOR2_X1 U21898 ( .A(n9334), .B(Key[24]), .ZN(n9336) );
  MUX2_X1 U21899 ( .A(n10589), .B(n11679), .S(n9341), .Z(n9347) );
  XNOR2_X1 U21902 ( .A(Key[99]), .B(Ciphertext[98]), .ZN(n9337) );
  AND2_X1 U21903 ( .A1(n9340), .A2(n9337), .ZN(n11688) );
  INV_X1 U21904 ( .A(n11688), .ZN(n9970) );
  INV_X1 U21905 ( .A(n9337), .ZN(n10594) );
  OAI22_X1 U21906 ( .A1(n11686), .A2(n9970), .B1(n9969), .B2(n11280), .ZN(
        n9338) );
  NAND2_X1 U21907 ( .A1(n9338), .A2(n10589), .ZN(n9346) );
  NAND2_X1 U21908 ( .A1(n11272), .A2(n9339), .ZN(n9981) );
  INV_X1 U21909 ( .A(n11671), .ZN(n9344) );
  NAND2_X1 U21910 ( .A1(n9337), .A2(n11276), .ZN(n9522) );
  INV_X1 U21911 ( .A(n11279), .ZN(n9520) );
  OAI21_X1 U21912 ( .B1(n9520), .B2(n9340), .A(n11276), .ZN(n9343) );
  NAND3_X1 U21913 ( .A1(n11270), .A2(n9973), .A3(n9974), .ZN(n9342) );
  OAI211_X1 U21914 ( .C1(n11279), .C2(n9347), .A(n9346), .B(n9345), .ZN(n10881) );
  NAND2_X1 U21916 ( .A1(n11696), .A2(n11695), .ZN(n9497) );
  INV_X1 U21917 ( .A(n9497), .ZN(n11200) );
  INV_X1 U21918 ( .A(n11714), .ZN(n9498) );
  OAI22_X1 U21919 ( .A1(n9498), .A2(n11203), .B1(n11697), .B2(n11705), .ZN(
        n9350) );
  NAND2_X1 U21920 ( .A1(n11697), .A2(n11695), .ZN(n9348) );
  OAI21_X1 U21921 ( .B1(n51650), .B2(n11697), .A(n9348), .ZN(n9349) );
  NOR2_X1 U21922 ( .A1(n11710), .A2(n11705), .ZN(n11208) );
  INV_X1 U21923 ( .A(n11204), .ZN(n9351) );
  OAI21_X1 U21924 ( .B1(n11211), .B2(n9491), .A(n9351), .ZN(n9352) );
  NAND2_X1 U21925 ( .A1(n11198), .A2(n11707), .ZN(n9494) );
  NAND2_X1 U21926 ( .A1(n11705), .A2(n11695), .ZN(n11699) );
  OAI21_X1 U21927 ( .B1(n11711), .B2(n11705), .A(n11699), .ZN(n9354) );
  NAND3_X1 U21928 ( .A1(n11711), .A2(n11696), .A3(n9926), .ZN(n9353) );
  OAI211_X1 U21929 ( .C1(n9500), .C2(n11711), .A(n9354), .B(n9353), .ZN(n9355)
         );
  INV_X1 U21930 ( .A(n13514), .ZN(n13521) );
  INV_X1 U21931 ( .A(n10881), .ZN(n13502) );
  NOR2_X1 U21932 ( .A1(n13502), .A2(n51683), .ZN(n12768) );
  INV_X1 U21933 ( .A(n12768), .ZN(n9356) );
  OAI211_X1 U21934 ( .C1(n13497), .C2(n12769), .A(n13521), .B(n9356), .ZN(
        n9359) );
  OAI211_X1 U21935 ( .C1(n13501), .C2(n11841), .A(n13525), .B(n13500), .ZN(
        n12936) );
  AOI21_X1 U21936 ( .B1(n11841), .B2(n51067), .A(n13514), .ZN(n9358) );
  XNOR2_X1 U21937 ( .A(n15677), .B(n17804), .ZN(n9450) );
  INV_X1 U21938 ( .A(Ciphertext[180]), .ZN(n9360) );
  XNOR2_X1 U21939 ( .A(Key[22]), .B(Ciphertext[183]), .ZN(n11354) );
  INV_X1 U21940 ( .A(Ciphertext[185]), .ZN(n9361) );
  INV_X1 U21941 ( .A(Ciphertext[182]), .ZN(n9362) );
  INV_X1 U21942 ( .A(Ciphertext[184]), .ZN(n9363) );
  XNOR2_X1 U21943 ( .A(n9363), .B(Key[125]), .ZN(n9365) );
  INV_X1 U21944 ( .A(n9365), .ZN(n12381) );
  NAND2_X1 U21945 ( .A1(n12373), .A2(n12381), .ZN(n9367) );
  INV_X1 U21946 ( .A(Ciphertext[181]), .ZN(n9364) );
  NAND3_X1 U21947 ( .A1(n51138), .A2(n12373), .A3(n10686), .ZN(n9366) );
  OAI211_X1 U21948 ( .C1(n10683), .C2(n9367), .A(n12092), .B(n9366), .ZN(n9368) );
  INV_X1 U21949 ( .A(n9368), .ZN(n9375) );
  INV_X1 U21950 ( .A(n11353), .ZN(n11352) );
  NAND2_X1 U21951 ( .A1(n12381), .A2(n11353), .ZN(n12391) );
  INV_X1 U21952 ( .A(n12084), .ZN(n12384) );
  NAND3_X1 U21953 ( .A1(n12389), .A2(n12373), .A3(n11352), .ZN(n9370) );
  INV_X1 U21954 ( .A(n12391), .ZN(n12376) );
  NAND2_X1 U21955 ( .A1(n12376), .A2(n51138), .ZN(n9687) );
  INV_X1 U21956 ( .A(n9687), .ZN(n9371) );
  AND2_X1 U21957 ( .A1(n12379), .A2(n10686), .ZN(n9680) );
  OAI21_X1 U21958 ( .B1(n9371), .B2(n12087), .A(n9680), .ZN(n9374) );
  NOR2_X1 U21959 ( .A1(n12088), .A2(n12383), .ZN(n9372) );
  OAI21_X1 U21961 ( .B1(n11351), .B2(n9372), .A(n12097), .ZN(n9373) );
  INV_X1 U21962 ( .A(n2149), .ZN(n13632) );
  AND2_X1 U21963 ( .A1(n12059), .A2(n10354), .ZN(n10661) );
  INV_X1 U21964 ( .A(n10665), .ZN(n12060) );
  NAND2_X1 U21965 ( .A1(n12060), .A2(n10355), .ZN(n9377) );
  NOR2_X1 U21966 ( .A1(n11393), .A2(n799), .ZN(n9376) );
  INV_X1 U21967 ( .A(n9378), .ZN(n9383) );
  AND2_X1 U21968 ( .A1(n9221), .A2(n799), .ZN(n9379) );
  AOI21_X1 U21969 ( .B1(n9379), .B2(n11388), .A(n12043), .ZN(n9382) );
  NAND2_X1 U21970 ( .A1(n9380), .A2(n10360), .ZN(n9381) );
  NAND3_X1 U21971 ( .A1(n11393), .A2(n10662), .A3(n12058), .ZN(n9385) );
  NAND2_X1 U21972 ( .A1(n9387), .A2(n11387), .ZN(n9391) );
  NAND3_X1 U21973 ( .A1(n10664), .A2(n12057), .A3(n799), .ZN(n9388) );
  OAI22_X1 U21974 ( .A1(n4797), .A2(n10715), .B1(n10722), .B2(n10724), .ZN(
        n9393) );
  OAI21_X1 U21975 ( .B1(n9704), .B2(n9393), .A(n10723), .ZN(n9398) );
  NAND2_X1 U21976 ( .A1(n10724), .A2(n12282), .ZN(n10224) );
  AND3_X1 U21977 ( .A1(n10234), .A2(n10224), .A3(n12294), .ZN(n9395) );
  OAI21_X1 U21978 ( .B1(n12285), .B2(n12282), .A(n12280), .ZN(n12284) );
  INV_X1 U21979 ( .A(n12284), .ZN(n9394) );
  INV_X1 U21980 ( .A(n12286), .ZN(n10235) );
  AOI22_X1 U21981 ( .A1(n9395), .A2(n9394), .B1(n10235), .B2(n12276), .ZN(
        n9397) );
  INV_X1 U21982 ( .A(n12276), .ZN(n12283) );
  OAI211_X1 U21983 ( .C1(n12283), .C2(n9699), .A(n10725), .B(n10716), .ZN(
        n9396) );
  INV_X1 U21984 ( .A(Ciphertext[186]), .ZN(n9400) );
  BUF_X2 U21985 ( .A(n9406), .Z(n11359) );
  INV_X1 U21986 ( .A(Ciphertext[189]), .ZN(n9401) );
  INV_X1 U21987 ( .A(n12107), .ZN(n9408) );
  INV_X1 U21988 ( .A(Ciphertext[190]), .ZN(n9402) );
  INV_X1 U21989 ( .A(n11361), .ZN(n11367) );
  INV_X1 U21990 ( .A(Ciphertext[187]), .ZN(n9403) );
  INV_X1 U21991 ( .A(n9407), .ZN(n10702) );
  NAND2_X1 U21992 ( .A1(n10702), .A2(n12117), .ZN(n9404) );
  AND2_X1 U21993 ( .A1(n12110), .A2(n9404), .ZN(n9416) );
  AND2_X1 U21995 ( .A1(n51256), .A2(n11375), .ZN(n9410) );
  XNOR2_X1 U21996 ( .A(n51391), .B(n12112), .ZN(n9409) );
  AOI22_X1 U21997 ( .A1(n9410), .A2(n12114), .B1(n9409), .B2(n9408), .ZN(n9415) );
  OAI211_X1 U21998 ( .C1(n11375), .C2(n12125), .A(n10702), .B(n51391), .ZN(
        n9411) );
  INV_X1 U21999 ( .A(n9411), .ZN(n9412) );
  INV_X1 U22000 ( .A(n12111), .ZN(n11370) );
  OAI211_X1 U22001 ( .C1(n11377), .C2(n11368), .A(n9412), .B(n11370), .ZN(
        n9414) );
  NOR2_X1 U22002 ( .A1(n10695), .A2(n10702), .ZN(n12121) );
  NAND3_X1 U22003 ( .A1(n12121), .A2(n11377), .A3(n11370), .ZN(n9413) );
  AND2_X1 U22004 ( .A1(n14666), .A2(n11315), .ZN(n13623) );
  NAND2_X1 U22005 ( .A1(n13622), .A2(n13623), .ZN(n13628) );
  INV_X1 U22006 ( .A(n12269), .ZN(n10735) );
  INV_X1 U22007 ( .A(n9417), .ZN(n11345) );
  INV_X1 U22008 ( .A(n12254), .ZN(n12264) );
  NOR2_X1 U22009 ( .A1(n10735), .A2(n12264), .ZN(n9418) );
  NOR2_X1 U22010 ( .A1(n9647), .A2(n9419), .ZN(n9420) );
  OAI21_X1 U22011 ( .B1(n12256), .B2(n9420), .A(n12243), .ZN(n9422) );
  NAND2_X1 U22012 ( .A1(n12257), .A2(n10741), .ZN(n9421) );
  INV_X1 U22013 ( .A(n9424), .ZN(n9428) );
  OAI21_X1 U22014 ( .B1(n10743), .B2(n10734), .A(n12241), .ZN(n9426) );
  OAI211_X1 U22015 ( .C1(n6267), .C2(n12243), .A(n9426), .B(n10747), .ZN(n9427) );
  NAND3_X1 U22016 ( .A1(n11406), .A2(n9602), .A3(n9430), .ZN(n9432) );
  OAI211_X1 U22017 ( .C1(n9433), .C2(n51141), .A(n11403), .B(n9429), .ZN(n9434) );
  AOI21_X1 U22018 ( .B1(n51141), .B2(n9598), .A(n438), .ZN(n9435) );
  OAI21_X1 U22019 ( .B1(n9435), .B2(n10385), .A(n12132), .ZN(n9436) );
  MUX2_X1 U22020 ( .A(n14664), .B(n12834), .S(n2150), .Z(n13630) );
  AOI22_X1 U22021 ( .A1(n9437), .A2(n783), .B1(n14672), .B2(n13630), .ZN(n9449) );
  NAND2_X1 U22022 ( .A1(n14665), .A2(n783), .ZN(n9441) );
  NAND2_X1 U22023 ( .A1(n14664), .A2(n2150), .ZN(n11311) );
  NAND2_X1 U22024 ( .A1(n783), .A2(n785), .ZN(n9438) );
  OAI22_X1 U22025 ( .A1(n9441), .A2(n12950), .B1(n11311), .B2(n9438), .ZN(
        n9440) );
  NOR2_X1 U22026 ( .A1(n12948), .A2(n6366), .ZN(n9439) );
  NOR2_X1 U22027 ( .A1(n9440), .A2(n9439), .ZN(n9448) );
  AND2_X1 U22028 ( .A1(n12834), .A2(n14666), .ZN(n9442) );
  OAI211_X1 U22029 ( .C1(n9442), .C2(n7755), .A(n9441), .B(n785), .ZN(n9444)
         );
  INV_X1 U22030 ( .A(n9442), .ZN(n13639) );
  OAI21_X1 U22031 ( .B1(n13639), .B2(n12950), .A(n13633), .ZN(n9443) );
  NAND2_X1 U22032 ( .A1(n9444), .A2(n9443), .ZN(n9447) );
  NOR2_X1 U22033 ( .A1(n14664), .A2(n14666), .ZN(n12840) );
  MUX2_X1 U22034 ( .A(n12840), .B(n14664), .S(n11315), .Z(n9445) );
  NAND2_X1 U22035 ( .A1(n9445), .A2(n13632), .ZN(n9446) );
  XNOR2_X1 U22036 ( .A(Key[136]), .B(Ciphertext[117]), .ZN(n9465) );
  INV_X1 U22037 ( .A(Ciphertext[114]), .ZN(n9451) );
  INV_X1 U22038 ( .A(Ciphertext[118]), .ZN(n9452) );
  AND2_X1 U22039 ( .A1(n10554), .A2(n10045), .ZN(n9951) );
  INV_X1 U22040 ( .A(n9459), .ZN(n10556) );
  NAND2_X1 U22041 ( .A1(n10556), .A2(n10552), .ZN(n9954) );
  INV_X1 U22042 ( .A(Ciphertext[115]), .ZN(n9453) );
  NOR2_X1 U22043 ( .A1(n9954), .A2(n10536), .ZN(n9961) );
  NAND2_X1 U22044 ( .A1(n9951), .A2(n9961), .ZN(n9964) );
  NAND3_X1 U22045 ( .A1(n10184), .A2(n10174), .A3(n9465), .ZN(n9458) );
  XOR2_X1 U22046 ( .A(Ciphertext[114]), .B(Ciphertext[117]), .Z(n9455) );
  XNOR2_X1 U22047 ( .A(Key[136]), .B(Key[19]), .ZN(n9454) );
  XNOR2_X1 U22048 ( .A(n9455), .B(n9454), .ZN(n10551) );
  INV_X1 U22049 ( .A(n10547), .ZN(n10179) );
  INV_X1 U22050 ( .A(n10554), .ZN(n10546) );
  NAND2_X1 U22051 ( .A1(n10541), .A2(n10179), .ZN(n9463) );
  NAND2_X1 U22052 ( .A1(n10536), .A2(n10540), .ZN(n9460) );
  NAND3_X1 U22053 ( .A1(n9826), .A2(n3850), .A3(n9460), .ZN(n9462) );
  MUX2_X1 U22054 ( .A(n9463), .B(n9462), .S(n10178), .Z(n9469) );
  OAI22_X1 U22055 ( .A1(n2093), .A2(n9464), .B1(n10555), .B2(n9826), .ZN(n9466) );
  AND2_X1 U22056 ( .A1(n10540), .A2(n51761), .ZN(n9953) );
  INV_X1 U22058 ( .A(n9952), .ZN(n10173) );
  NOR2_X1 U22059 ( .A1(n52185), .A2(n10607), .ZN(n9471) );
  AOI22_X1 U22060 ( .A1(n10605), .A2(n9471), .B1(n51212), .B2(n10065), .ZN(
        n9475) );
  INV_X1 U22061 ( .A(n9915), .ZN(n10608) );
  INV_X1 U22062 ( .A(n10610), .ZN(n9907) );
  INV_X1 U22063 ( .A(n9908), .ZN(n9906) );
  NAND3_X1 U22065 ( .A1(n10619), .A2(n9914), .A3(n10618), .ZN(n9472) );
  NAND4_X1 U22066 ( .A1(n9475), .A2(n9474), .A3(n9473), .A4(n9472), .ZN(n9479)
         );
  NOR2_X1 U22067 ( .A1(n10610), .A2(n51212), .ZN(n10603) );
  INV_X1 U22068 ( .A(n10603), .ZN(n9477) );
  NAND2_X1 U22069 ( .A1(n10525), .A2(n10031), .ZN(n10110) );
  NAND3_X1 U22070 ( .A1(n10513), .A2(n10520), .A3(n10110), .ZN(n10511) );
  AOI21_X1 U22071 ( .B1(n10525), .B2(n10026), .A(n10101), .ZN(n9480) );
  AND2_X1 U22072 ( .A1(n10527), .A2(n10530), .ZN(n10104) );
  AND2_X1 U22074 ( .A1(n9481), .A2(n10511), .ZN(n9490) );
  NAND2_X1 U22075 ( .A1(n10519), .A2(n9482), .ZN(n9483) );
  OAI21_X1 U22076 ( .B1(n10031), .B2(n10026), .A(n9483), .ZN(n9485) );
  NAND2_X1 U22077 ( .A1(n10097), .A2(n10110), .ZN(n10033) );
  INV_X1 U22078 ( .A(n10033), .ZN(n9486) );
  NAND2_X1 U22079 ( .A1(n9486), .A2(n10513), .ZN(n9487) );
  NAND2_X1 U22080 ( .A1(n9494), .A2(n9926), .ZN(n9493) );
  OAI21_X1 U22081 ( .B1(n11210), .B2(n11209), .A(n9146), .ZN(n9492) );
  NAND4_X1 U22082 ( .A1(n9493), .A2(n9492), .A3(n9491), .A4(n11203), .ZN(n9506) );
  INV_X1 U22083 ( .A(n9494), .ZN(n11214) );
  OAI22_X1 U22084 ( .A1(n11210), .A2(n9495), .B1(n51182), .B2(n11704), .ZN(
        n9496) );
  NOR2_X1 U22085 ( .A1(n9498), .A2(n9497), .ZN(n9936) );
  NAND2_X1 U22086 ( .A1(n9936), .A2(n11715), .ZN(n9504) );
  NAND2_X1 U22087 ( .A1(n9499), .A2(n9926), .ZN(n9933) );
  NOR2_X1 U22088 ( .A1(n13092), .A2(n13088), .ZN(n12823) );
  INV_X1 U22089 ( .A(n11650), .ZN(n9507) );
  NAND2_X1 U22090 ( .A1(n9507), .A2(n11658), .ZN(n10571) );
  INV_X1 U22091 ( .A(n10571), .ZN(n9509) );
  OAI211_X1 U22092 ( .C1(n9939), .C2(n11650), .A(n9511), .B(n11641), .ZN(n9512) );
  NAND2_X1 U22093 ( .A1(n9512), .A2(n11644), .ZN(n9514) );
  AND2_X1 U22094 ( .A1(n10563), .A2(n11639), .ZN(n9943) );
  NAND2_X1 U22095 ( .A1(n9939), .A2(n11662), .ZN(n11643) );
  NAND3_X1 U22096 ( .A1(n9943), .A2(n11644), .A3(n11643), .ZN(n9517) );
  AND2_X1 U22097 ( .A1(n11657), .A2(n9517), .ZN(n9518) );
  INV_X1 U22098 ( .A(n9519), .ZN(n11687) );
  INV_X1 U22099 ( .A(n11683), .ZN(n10587) );
  OAI21_X1 U22100 ( .B1(n11274), .B2(n10587), .A(n9520), .ZN(n9521) );
  INV_X1 U22101 ( .A(n11669), .ZN(n9980) );
  NOR2_X1 U22102 ( .A1(n9974), .A2(n9980), .ZN(n9524) );
  NOR2_X1 U22103 ( .A1(n11672), .A2(n9524), .ZN(n9528) );
  NAND3_X1 U22104 ( .A1(n11688), .A2(n11670), .A3(n11683), .ZN(n9527) );
  NOR2_X1 U22105 ( .A1(n11687), .A2(n11275), .ZN(n9525) );
  NAND2_X1 U22106 ( .A1(n10590), .A2(n9969), .ZN(n11668) );
  OAI211_X1 U22107 ( .C1(n11270), .C2(n9525), .A(n9341), .B(n11668), .ZN(n9526) );
  INV_X1 U22108 ( .A(n12914), .ZN(n11160) );
  NAND2_X1 U22109 ( .A1(n9529), .A2(n11160), .ZN(n9533) );
  OR2_X1 U22110 ( .A1(n13086), .A2(n12915), .ZN(n13100) );
  AND2_X1 U22111 ( .A1(n12914), .A2(n1244), .ZN(n11824) );
  NAND2_X1 U22112 ( .A1(n11824), .A2(n13090), .ZN(n11168) );
  NAND2_X1 U22113 ( .A1(n11160), .A2(n13086), .ZN(n13082) );
  NOR2_X1 U22114 ( .A1(n13091), .A2(n13089), .ZN(n13076) );
  NOR2_X1 U22115 ( .A1(n13086), .A2(n13088), .ZN(n13105) );
  NAND2_X1 U22116 ( .A1(n13086), .A2(n13088), .ZN(n9530) );
  NOR2_X1 U22117 ( .A1(n13091), .A2(n9530), .ZN(n9531) );
  XNOR2_X1 U22118 ( .A(n4817), .B(n4568), .ZN(n25744) );
  XNOR2_X1 U22119 ( .A(n25744), .B(n4647), .ZN(n17243) );
  XNOR2_X1 U22120 ( .A(n47737), .B(n4589), .ZN(n27174) );
  XNOR2_X1 U22121 ( .A(n17243), .B(n27174), .ZN(n9534) );
  XNOR2_X2 U22122 ( .A(n47401), .B(n4800), .ZN(n43691) );
  XNOR2_X1 U22123 ( .A(n48597), .B(n4121), .ZN(n37288) );
  XNOR2_X1 U22124 ( .A(n43691), .B(n37288), .ZN(n28303) );
  XNOR2_X1 U22125 ( .A(n9534), .B(n28303), .ZN(n44909) );
  XNOR2_X1 U22126 ( .A(Key[2]), .B(Key[170]), .ZN(n18636) );
  XNOR2_X1 U22127 ( .A(n4641), .B(n4353), .ZN(n9535) );
  XNOR2_X1 U22128 ( .A(n18636), .B(n9535), .ZN(n34113) );
  XNOR2_X1 U22129 ( .A(n44909), .B(n34113), .ZN(n9536) );
  XNOR2_X1 U22130 ( .A(n16904), .B(n9536), .ZN(n9631) );
  NOR2_X1 U22131 ( .A1(n12600), .A2(n9538), .ZN(n11139) );
  NAND2_X1 U22132 ( .A1(n11139), .A2(n3377), .ZN(n9541) );
  NOR2_X1 U22133 ( .A1(n51140), .A2(n52140), .ZN(n9543) );
  NOR2_X1 U22135 ( .A1(n10471), .A2(n12590), .ZN(n11128) );
  NAND3_X1 U22136 ( .A1(n11132), .A2(n9539), .A3(n9548), .ZN(n9550) );
  NAND2_X1 U22137 ( .A1(n11920), .A2(n51140), .ZN(n9549) );
  AND2_X1 U22138 ( .A1(n9550), .A2(n9549), .ZN(n9554) );
  NAND2_X1 U22139 ( .A1(n9551), .A2(n795), .ZN(n9553) );
  AND2_X1 U22142 ( .A1(n12659), .A2(n12663), .ZN(n12647) );
  INV_X1 U22143 ( .A(n12647), .ZN(n9557) );
  NAND3_X1 U22144 ( .A1(n10445), .A2(n10451), .A3(n12649), .ZN(n9560) );
  NAND2_X1 U22145 ( .A1(n11979), .A2(n12649), .ZN(n11985) );
  NAND3_X1 U22146 ( .A1(n10451), .A2(n794), .A3(n11985), .ZN(n9559) );
  NAND2_X1 U22147 ( .A1(n9560), .A2(n9559), .ZN(n9561) );
  NAND2_X1 U22148 ( .A1(n10338), .A2(n10449), .ZN(n9563) );
  AND2_X1 U22149 ( .A1(n11978), .A2(n11984), .ZN(n12658) );
  NAND2_X1 U22150 ( .A1(n12658), .A2(n11979), .ZN(n9562) );
  MUX2_X1 U22151 ( .A(n9563), .B(n9562), .S(n10456), .Z(n9615) );
  AND2_X1 U22152 ( .A1(n15259), .A2(n14784), .ZN(n14134) );
  INV_X1 U22153 ( .A(n14134), .ZN(n9626) );
  INV_X1 U22155 ( .A(n12071), .ZN(n12640) );
  NAND3_X1 U22156 ( .A1(n10463), .A2(n10462), .A3(n9208), .ZN(n9565) );
  NOR2_X1 U22157 ( .A1(n12637), .A2(n12627), .ZN(n12624) );
  NOR2_X1 U22158 ( .A1(n12073), .A2(n10465), .ZN(n9567) );
  AOI22_X1 U22159 ( .A1(n12624), .A2(n12632), .B1(n9567), .B2(n12069), .ZN(
        n9572) );
  NOR2_X1 U22160 ( .A1(n12073), .A2(n51432), .ZN(n10319) );
  OAI21_X1 U22161 ( .B1(n12631), .B2(n12619), .A(n12618), .ZN(n9568) );
  OAI211_X1 U22162 ( .C1(n10319), .C2(n9568), .A(n10465), .B(n12617), .ZN(
        n9571) );
  NAND2_X1 U22163 ( .A1(n12616), .A2(n12631), .ZN(n9569) );
  OAI211_X1 U22164 ( .C1(n12616), .C2(n12068), .A(n9569), .B(n12620), .ZN(
        n9570) );
  INV_X1 U22165 ( .A(n11108), .ZN(n12729) );
  NAND2_X1 U22166 ( .A1(n12729), .A2(n12722), .ZN(n11111) );
  INV_X1 U22167 ( .A(n11111), .ZN(n9574) );
  INV_X1 U22168 ( .A(n11943), .ZN(n11105) );
  NAND2_X1 U22169 ( .A1(n8881), .A2(n5484), .ZN(n9575) );
  NAND2_X1 U22170 ( .A1(n11961), .A2(n9575), .ZN(n9577) );
  NAND2_X1 U22171 ( .A1(n12720), .A2(n8881), .ZN(n11948) );
  INV_X1 U22172 ( .A(n11948), .ZN(n9576) );
  NAND2_X1 U22173 ( .A1(n9576), .A2(n8885), .ZN(n9578) );
  NAND2_X1 U22174 ( .A1(n9577), .A2(n9578), .ZN(n9580) );
  AOI21_X1 U22175 ( .B1(n9578), .B2(n12720), .A(n12728), .ZN(n9579) );
  NAND2_X1 U22176 ( .A1(n9580), .A2(n9579), .ZN(n9583) );
  OAI21_X1 U22177 ( .B1(n10431), .B2(n12722), .A(n11108), .ZN(n9581) );
  INV_X1 U22179 ( .A(n12160), .ZN(n12179) );
  OAI21_X1 U22180 ( .B1(n11322), .B2(n12179), .A(n9584), .ZN(n9586) );
  NAND4_X1 U22181 ( .A1(n548), .A2(n52132), .A3(n10413), .A4(n12166), .ZN(
        n9587) );
  OAI21_X1 U22182 ( .B1(n9591), .B2(n10328), .A(n9587), .ZN(n9588) );
  INV_X1 U22183 ( .A(n9588), .ZN(n9596) );
  INV_X1 U22184 ( .A(n10418), .ZN(n12156) );
  NAND2_X1 U22185 ( .A1(n548), .A2(n9589), .ZN(n9590) );
  OAI211_X1 U22186 ( .C1(n12156), .C2(n12173), .A(n9591), .B(n9590), .ZN(n9592) );
  NAND2_X1 U22187 ( .A1(n9592), .A2(n11328), .ZN(n9595) );
  OAI21_X1 U22188 ( .B1(n9626), .B2(n13069), .A(n13065), .ZN(n9597) );
  INV_X1 U22189 ( .A(n9597), .ZN(n9630) );
  NOR2_X1 U22191 ( .A1(n793), .A2(n12132), .ZN(n9600) );
  NAND2_X1 U22192 ( .A1(n11423), .A2(n9598), .ZN(n11401) );
  OAI21_X1 U22193 ( .B1(n11401), .B2(n11402), .A(n12133), .ZN(n9599) );
  OAI21_X1 U22194 ( .B1(n9601), .B2(n9600), .A(n9599), .ZN(n9613) );
  OAI211_X1 U22195 ( .C1(n12139), .C2(n12129), .A(n11399), .B(n9602), .ZN(
        n9603) );
  NAND2_X1 U22196 ( .A1(n9603), .A2(n12130), .ZN(n9612) );
  INV_X1 U22198 ( .A(n12138), .ZN(n11422) );
  OAI211_X1 U22199 ( .C1(n11422), .C2(n12129), .A(n9607), .B(n9606), .ZN(n9608) );
  INV_X1 U22200 ( .A(n9608), .ZN(n9611) );
  INV_X1 U22201 ( .A(n11416), .ZN(n9609) );
  NAND2_X1 U22202 ( .A1(n9609), .A2(n51141), .ZN(n9610) );
  NAND2_X1 U22203 ( .A1(n14784), .A2(n15256), .ZN(n14791) );
  NAND2_X1 U22204 ( .A1(n14791), .A2(n51685), .ZN(n9614) );
  OAI211_X1 U22205 ( .C1(n15264), .C2(n13061), .A(n9614), .B(n15260), .ZN(
        n9625) );
  INV_X1 U22206 ( .A(n9615), .ZN(n9618) );
  INV_X1 U22207 ( .A(n9616), .ZN(n9617) );
  INV_X1 U22208 ( .A(n13061), .ZN(n14790) );
  OAI21_X1 U22209 ( .B1(n9618), .B2(n9617), .A(n14790), .ZN(n9619) );
  AOI22_X1 U22211 ( .A1(n15257), .A2(n9619), .B1(n14790), .B2(n15263), .ZN(
        n9620) );
  AND2_X1 U22212 ( .A1(n15259), .A2(n14783), .ZN(n14794) );
  NAND2_X1 U22213 ( .A1(n9620), .A2(n14794), .ZN(n9624) );
  NOR2_X1 U22214 ( .A1(n13057), .A2(n13069), .ZN(n9622) );
  NAND2_X1 U22215 ( .A1(n14784), .A2(n13061), .ZN(n14797) );
  INV_X1 U22216 ( .A(n14797), .ZN(n9621) );
  NAND2_X1 U22217 ( .A1(n15256), .A2(n14783), .ZN(n13058) );
  AOI22_X1 U22218 ( .A1(n9622), .A2(n51685), .B1(n9621), .B2(n13058), .ZN(
        n9623) );
  NAND2_X1 U22219 ( .A1(n9626), .A2(n14790), .ZN(n9628) );
  NOR2_X1 U22220 ( .A1(n14783), .A2(n15256), .ZN(n9627) );
  NAND2_X1 U22221 ( .A1(n9628), .A2(n9627), .ZN(n9629) );
  XNOR2_X1 U22222 ( .A(n9631), .B(n17125), .ZN(n9803) );
  NAND2_X1 U22224 ( .A1(n9636), .A2(n12107), .ZN(n10372) );
  NOR2_X1 U22225 ( .A1(n9407), .A2(n11375), .ZN(n10374) );
  OAI21_X1 U22226 ( .B1(n10373), .B2(n9633), .A(n10374), .ZN(n9634) );
  AND2_X1 U22227 ( .A1(n9635), .A2(n9634), .ZN(n9694) );
  INV_X1 U22228 ( .A(n10374), .ZN(n12118) );
  AND2_X1 U22229 ( .A1(n11377), .A2(n12112), .ZN(n12105) );
  NAND2_X1 U22230 ( .A1(n11359), .A2(n12117), .ZN(n10709) );
  NAND2_X1 U22231 ( .A1(n10709), .A2(n12117), .ZN(n9637) );
  NAND3_X1 U22232 ( .A1(n11365), .A2(n12105), .A3(n9637), .ZN(n9638) );
  NAND2_X1 U22233 ( .A1(n11375), .A2(n12117), .ZN(n12106) );
  NAND2_X1 U22234 ( .A1(n12112), .A2(n10375), .ZN(n9639) );
  AND2_X1 U22235 ( .A1(n12112), .A2(n11375), .ZN(n10704) );
  NAND2_X1 U22238 ( .A1(n12250), .A2(n12253), .ZN(n9642) );
  AOI21_X1 U22239 ( .B1(n9643), .B2(n9642), .A(n11345), .ZN(n9651) );
  INV_X1 U22240 ( .A(n12256), .ZN(n9644) );
  NAND2_X1 U22241 ( .A1(n12257), .A2(n9644), .ZN(n9645) );
  AOI21_X1 U22242 ( .B1(n9646), .B2(n10735), .A(n9645), .ZN(n9650) );
  AOI21_X1 U22243 ( .B1(n6267), .B2(n11345), .A(n10734), .ZN(n9648) );
  OAI22_X1 U22244 ( .A1(n9648), .A2(n11346), .B1(n10742), .B2(n12263), .ZN(
        n9649) );
  NAND2_X1 U22245 ( .A1(n13841), .A2(n13849), .ZN(n13839) );
  NAND4_X1 U22246 ( .A1(n9653), .A2(n10302), .A3(n12317), .A4(n9652), .ZN(
        n9664) );
  NOR2_X1 U22249 ( .A1(n2313), .A2(n9655), .ZN(n9663) );
  NAND4_X1 U22250 ( .A1(n9758), .A2(n12301), .A3(n10296), .A4(n9656), .ZN(
        n9660) );
  AND2_X1 U22251 ( .A1(n12301), .A2(n12314), .ZN(n10303) );
  INV_X1 U22252 ( .A(n10939), .ZN(n10300) );
  INV_X1 U22253 ( .A(n9657), .ZN(n9658) );
  NAND4_X1 U22254 ( .A1(n10303), .A2(n10300), .A3(n9658), .A4(n9656), .ZN(
        n9659) );
  AND2_X1 U22255 ( .A1(n9660), .A2(n9659), .ZN(n9662) );
  INV_X1 U22256 ( .A(n12328), .ZN(n9737) );
  NAND3_X1 U22257 ( .A1(n9737), .A2(n10672), .A3(n12344), .ZN(n9666) );
  NAND2_X1 U22258 ( .A1(n10277), .A2(n10671), .ZN(n9665) );
  AND2_X1 U22259 ( .A1(n9666), .A2(n9665), .ZN(n9674) );
  AND2_X1 U22260 ( .A1(n51004), .A2(n9667), .ZN(n9669) );
  OAI21_X1 U22261 ( .B1(n10672), .B2(n9669), .A(n9668), .ZN(n9670) );
  NAND2_X1 U22262 ( .A1(n10279), .A2(n12336), .ZN(n12322) );
  NAND3_X1 U22263 ( .A1(n9670), .A2(n12341), .A3(n12322), .ZN(n9673) );
  AOI22_X1 U22264 ( .A1(n10673), .A2(n3649), .B1(n10676), .B2(n12333), .ZN(
        n9672) );
  NAND3_X1 U22266 ( .A1(n12334), .A2(n12332), .A3(n12344), .ZN(n9671) );
  AND2_X1 U22267 ( .A1(n13855), .A2(n13845), .ZN(n13552) );
  INV_X1 U22268 ( .A(n13841), .ZN(n13844) );
  AND3_X1 U22269 ( .A1(n13849), .A2(n13855), .A3(n13845), .ZN(n9690) );
  NAND2_X1 U22270 ( .A1(n11353), .A2(n10687), .ZN(n12094) );
  NOR2_X1 U22271 ( .A1(n12094), .A2(n12373), .ZN(n9676) );
  OAI21_X1 U22272 ( .B1(n12088), .B2(n12380), .A(n12383), .ZN(n9675) );
  AND2_X1 U22273 ( .A1(n12373), .A2(n10686), .ZN(n12085) );
  NAND3_X1 U22274 ( .A1(n12085), .A2(n12094), .A3(n12088), .ZN(n9678) );
  AND2_X1 U22275 ( .A1(n9678), .A2(n9677), .ZN(n9683) );
  INV_X1 U22276 ( .A(n12094), .ZN(n12370) );
  NAND3_X1 U22277 ( .A1(n9680), .A2(n12370), .A3(n9679), .ZN(n9681) );
  NAND2_X1 U22278 ( .A1(n12088), .A2(n12383), .ZN(n12095) );
  NAND2_X1 U22279 ( .A1(n12380), .A2(n12383), .ZN(n9684) );
  AND2_X1 U22280 ( .A1(n12092), .A2(n9684), .ZN(n9686) );
  NAND3_X1 U22281 ( .A1(n12087), .A2(n7895), .A3(n12383), .ZN(n9685) );
  OAI211_X1 U22282 ( .C1(n12095), .C2(n12391), .A(n9686), .B(n9685), .ZN(n9689) );
  AND2_X1 U22283 ( .A1(n9689), .A2(n9688), .ZN(n11730) );
  NOR2_X1 U22284 ( .A1(n13855), .A2(n13845), .ZN(n11780) );
  INV_X1 U22287 ( .A(n9694), .ZN(n9712) );
  INV_X1 U22288 ( .A(n9695), .ZN(n9697) );
  NAND3_X1 U22289 ( .A1(n9697), .A2(n9696), .A3(n304), .ZN(n9711) );
  AOI21_X1 U22290 ( .B1(n9700), .B2(n10722), .A(n12291), .ZN(n9701) );
  OAI21_X1 U22291 ( .B1(n9703), .B2(n9702), .A(n9701), .ZN(n9709) );
  NAND3_X1 U22292 ( .A1(n12283), .A2(n10725), .A3(n12291), .ZN(n9707) );
  NAND2_X1 U22293 ( .A1(n10225), .A2(n12291), .ZN(n9706) );
  INV_X1 U22294 ( .A(n9704), .ZN(n9705) );
  INV_X1 U22295 ( .A(n9720), .ZN(n9710) );
  OAI21_X1 U22296 ( .B1(n9712), .B2(n9711), .A(n9710), .ZN(n11738) );
  NAND2_X1 U22297 ( .A1(n10715), .A2(n12291), .ZN(n10719) );
  INV_X1 U22298 ( .A(n10716), .ZN(n9713) );
  NAND2_X1 U22299 ( .A1(n12276), .A2(n12282), .ZN(n9714) );
  OAI21_X1 U22300 ( .B1(n12280), .B2(n12276), .A(n9714), .ZN(n9715) );
  NAND2_X1 U22301 ( .A1(n9715), .A2(n10726), .ZN(n9716) );
  NOR2_X1 U22304 ( .A1(n14482), .A2(n13854), .ZN(n13559) );
  NAND2_X1 U22305 ( .A1(n14473), .A2(n13854), .ZN(n13547) );
  INV_X1 U22306 ( .A(n13547), .ZN(n9723) );
  OAI211_X1 U22307 ( .C1(n13841), .C2(n13845), .A(n13854), .B(n13856), .ZN(
        n9722) );
  OAI211_X1 U22308 ( .C1(n9723), .C2(n13856), .A(n9722), .B(n14482), .ZN(n9726) );
  NAND2_X1 U22309 ( .A1(n14473), .A2(n13849), .ZN(n13550) );
  OAI21_X1 U22310 ( .B1(n13550), .B2(n13853), .A(n9724), .ZN(n11741) );
  NAND2_X1 U22311 ( .A1(n11741), .A2(n14472), .ZN(n9725) );
  NAND2_X1 U22312 ( .A1(n10924), .A2(n9807), .ZN(n9729) );
  NAND2_X1 U22313 ( .A1(n10144), .A2(n9729), .ZN(n9731) );
  AOI22_X1 U22314 ( .A1(n10219), .A2(n8840), .B1(n10222), .B2(n10148), .ZN(
        n9730) );
  OR2_X1 U22315 ( .A1(n10217), .A2(n10143), .ZN(n10933) );
  NAND2_X1 U22317 ( .A1(n10221), .A2(n10925), .ZN(n9732) );
  OAI211_X1 U22318 ( .C1(n10222), .C2(n10142), .A(n9732), .B(n10921), .ZN(
        n9734) );
  NAND2_X1 U22319 ( .A1(n10926), .A2(n10143), .ZN(n9733) );
  AND2_X1 U22320 ( .A1(n51004), .A2(n12336), .ZN(n10282) );
  NAND2_X1 U22321 ( .A1(n12337), .A2(n12323), .ZN(n9739) );
  INV_X1 U22323 ( .A(n12339), .ZN(n10285) );
  OAI22_X1 U22324 ( .A1(n9737), .A2(n51194), .B1(n10277), .B2(n10285), .ZN(
        n9738) );
  AND2_X1 U22325 ( .A1(n10671), .A2(n10288), .ZN(n10678) );
  AOI21_X1 U22326 ( .B1(n9739), .B2(n12333), .A(n52199), .ZN(n9740) );
  OR2_X1 U22328 ( .A1(n9740), .A2(n12321), .ZN(n9741) );
  XNOR2_X1 U22329 ( .A(n14234), .B(n14228), .ZN(n9779) );
  INV_X1 U22330 ( .A(n11005), .ZN(n10247) );
  NAND2_X1 U22331 ( .A1(n9744), .A2(n11015), .ZN(n11012) );
  INV_X1 U22332 ( .A(n11012), .ZN(n9749) );
  INV_X1 U22333 ( .A(n9755), .ZN(n9757) );
  OAI21_X1 U22334 ( .B1(n10296), .B2(n12314), .A(n12317), .ZN(n9756) );
  OAI211_X1 U22335 ( .C1(n10300), .C2(n12317), .A(n9757), .B(n9756), .ZN(n9761) );
  NAND3_X1 U22336 ( .A1(n9758), .A2(n12301), .A3(n9772), .ZN(n9760) );
  INV_X1 U22337 ( .A(n10938), .ZN(n12304) );
  NAND2_X1 U22338 ( .A1(n10945), .A2(n12304), .ZN(n9759) );
  AND3_X1 U22339 ( .A1(n9761), .A2(n9760), .A3(n9759), .ZN(n9778) );
  NOR2_X1 U22340 ( .A1(n9758), .A2(n9772), .ZN(n9766) );
  NOR2_X1 U22341 ( .A1(n9763), .A2(n12314), .ZN(n9764) );
  AOI22_X1 U22342 ( .A1(n9766), .A2(n12304), .B1(n9765), .B2(n9764), .ZN(n9777) );
  INV_X1 U22343 ( .A(n9767), .ZN(n12307) );
  AND2_X1 U22344 ( .A1(n10302), .A2(n12315), .ZN(n10292) );
  AND2_X1 U22345 ( .A1(n10302), .A2(n12314), .ZN(n12302) );
  NAND3_X1 U22346 ( .A1(n9767), .A2(n12302), .A3(n12312), .ZN(n9768) );
  OAI211_X1 U22347 ( .C1(n9770), .C2(n12307), .A(n9769), .B(n9768), .ZN(n9771)
         );
  INV_X1 U22348 ( .A(n9771), .ZN(n9776) );
  OAI21_X1 U22349 ( .B1(n9774), .B2(n12301), .A(n9773), .ZN(n9775) );
  NAND3_X1 U22350 ( .A1(n9779), .A2(n13971), .A3(n13968), .ZN(n13225) );
  INV_X1 U22351 ( .A(n9780), .ZN(n10978) );
  NAND2_X1 U22352 ( .A1(n10259), .A2(n8791), .ZN(n9791) );
  NAND2_X1 U22353 ( .A1(n9786), .A2(n12356), .ZN(n10265) );
  OAI21_X1 U22354 ( .B1(n10267), .B2(n10272), .A(n10262), .ZN(n9784) );
  NAND2_X1 U22355 ( .A1(n9785), .A2(n9784), .ZN(n9790) );
  NOR2_X1 U22356 ( .A1(n9786), .A2(n12350), .ZN(n9788) );
  INV_X1 U22357 ( .A(n9787), .ZN(n12357) );
  OAI211_X1 U22358 ( .C1(n10988), .C2(n9788), .A(n10983), .B(n12357), .ZN(
        n9789) );
  NAND4_X1 U22359 ( .A1(n9791), .A2(n10265), .A3(n9790), .A4(n9789), .ZN(n9792) );
  NOR2_X1 U22360 ( .A1(n10954), .A2(n3316), .ZN(n9793) );
  NAND2_X1 U22361 ( .A1(n10960), .A2(n9856), .ZN(n9849) );
  OR2_X1 U22362 ( .A1(n9849), .A2(n10956), .ZN(n10060) );
  INV_X1 U22363 ( .A(n10054), .ZN(n9860) );
  OAI21_X1 U22364 ( .B1(n9859), .B2(n10954), .A(n6004), .ZN(n9794) );
  NAND2_X1 U22365 ( .A1(n9794), .A2(n10957), .ZN(n9796) );
  NAND2_X1 U22366 ( .A1(n10051), .A2(n10124), .ZN(n13231) );
  INV_X1 U22367 ( .A(n10119), .ZN(n13230) );
  NAND3_X1 U22368 ( .A1(n13231), .A2(n13230), .A3(n9856), .ZN(n9797) );
  INV_X1 U22369 ( .A(n14224), .ZN(n13226) );
  NOR2_X1 U22370 ( .A1(n13221), .A2(n14224), .ZN(n9798) );
  NOR2_X1 U22371 ( .A1(n13968), .A2(n14220), .ZN(n13958) );
  AND2_X1 U22372 ( .A1(n14220), .A2(n14234), .ZN(n13216) );
  NAND2_X1 U22374 ( .A1(n14224), .A2(n14220), .ZN(n12923) );
  OAI21_X1 U22375 ( .B1(n13960), .B2(n14234), .A(n13221), .ZN(n9799) );
  AND2_X1 U22376 ( .A1(n14220), .A2(n13968), .ZN(n13222) );
  NAND2_X1 U22377 ( .A1(n9799), .A2(n13222), .ZN(n9800) );
  NAND2_X1 U22378 ( .A1(n10134), .A2(n10216), .ZN(n10918) );
  AND2_X1 U22379 ( .A1(n8840), .A2(n10925), .ZN(n9804) );
  NOR2_X1 U22380 ( .A1(n10217), .A2(n9804), .ZN(n9805) );
  AOI22_X1 U22381 ( .A1(n10918), .A2(n9805), .B1(n10935), .B2(n10219), .ZN(
        n9817) );
  INV_X1 U22382 ( .A(n9808), .ZN(n9810) );
  INV_X1 U22383 ( .A(n10922), .ZN(n10214) );
  AND2_X1 U22384 ( .A1(n10221), .A2(n10919), .ZN(n10140) );
  OAI211_X1 U22385 ( .C1(n9810), .C2(n10920), .A(n9809), .B(n10140), .ZN(n9816) );
  NAND2_X1 U22386 ( .A1(n10219), .A2(n10134), .ZN(n9811) );
  NAND4_X1 U22387 ( .A1(n9811), .A2(n10147), .A3(n10926), .A4(n10218), .ZN(
        n9815) );
  INV_X1 U22388 ( .A(n10137), .ZN(n10215) );
  INV_X1 U22389 ( .A(n10926), .ZN(n9812) );
  OAI21_X1 U22390 ( .B1(n10215), .B2(n9812), .A(n10921), .ZN(n9813) );
  NAND2_X1 U22391 ( .A1(n9813), .A2(n10216), .ZN(n9814) );
  NOR2_X1 U22392 ( .A1(n11036), .A2(n580), .ZN(n10586) );
  OAI21_X1 U22393 ( .B1(n11032), .B2(n10162), .A(n8639), .ZN(n9819) );
  NAND3_X1 U22394 ( .A1(n8410), .A2(n11027), .A3(n10578), .ZN(n9818) );
  AND2_X1 U22395 ( .A1(n9819), .A2(n9818), .ZN(n9824) );
  NOR2_X1 U22396 ( .A1(n10169), .A2(n580), .ZN(n9821) );
  NOR2_X1 U22397 ( .A1(n2197), .A2(n10584), .ZN(n9820) );
  AOI22_X1 U22398 ( .A1(n9821), .A2(n11025), .B1(n11032), .B2(n9820), .ZN(
        n9823) );
  NOR2_X1 U22399 ( .A1(n2173), .A2(n51657), .ZN(n13200) );
  NAND2_X1 U22400 ( .A1(n803), .A2(n10540), .ZN(n10177) );
  OAI22_X1 U22401 ( .A1(n10177), .A2(n9464), .B1(n9826), .B2(n10037), .ZN(
        n9827) );
  NOR2_X1 U22402 ( .A1(n9827), .A2(n9961), .ZN(n9834) );
  OAI22_X1 U22403 ( .A1(n2093), .A2(n9952), .B1(n9464), .B2(n10539), .ZN(n9828) );
  NAND2_X1 U22404 ( .A1(n9828), .A2(n10179), .ZN(n9833) );
  NAND2_X1 U22405 ( .A1(n9829), .A2(n10174), .ZN(n9832) );
  NAND2_X1 U22406 ( .A1(n9464), .A2(n10540), .ZN(n10038) );
  OAI211_X1 U22407 ( .C1(n9830), .C2(n10552), .A(n10038), .B(n10555), .ZN(
        n9831) );
  MUX2_X1 U22408 ( .A(n51657), .B(n13200), .S(n13207), .Z(n9870) );
  OAI21_X1 U22409 ( .B1(n10633), .B2(n10530), .A(n9835), .ZN(n10107) );
  INV_X1 U22410 ( .A(n10107), .ZN(n9838) );
  NAND3_X1 U22411 ( .A1(n10532), .A2(n10096), .A3(n10110), .ZN(n9837) );
  OAI211_X1 U22414 ( .C1(n9838), .C2(n10105), .A(n9837), .B(n10632), .ZN(n9847) );
  NAND3_X1 U22415 ( .A1(n10508), .A2(n10026), .A3(n10633), .ZN(n10516) );
  OAI21_X1 U22416 ( .B1(n8853), .B2(n10095), .A(n10516), .ZN(n9839) );
  NAND2_X1 U22417 ( .A1(n9839), .A2(n10104), .ZN(n9845) );
  NOR2_X1 U22418 ( .A1(n10100), .A2(n10031), .ZN(n10521) );
  INV_X1 U22419 ( .A(n10521), .ZN(n9844) );
  NAND2_X1 U22420 ( .A1(n10529), .A2(n10096), .ZN(n9840) );
  OAI21_X1 U22421 ( .B1(n10110), .B2(n10096), .A(n9840), .ZN(n9841) );
  NAND2_X1 U22422 ( .A1(n9841), .A2(n9484), .ZN(n9843) );
  NAND4_X1 U22423 ( .A1(n9845), .A2(n9844), .A3(n9843), .A4(n9842), .ZN(n9846)
         );
  OAI21_X1 U22425 ( .B1(n9849), .B2(n10962), .A(n9848), .ZN(n9854) );
  AOI21_X1 U22426 ( .B1(n9852), .B2(n9851), .A(n9858), .ZN(n9853) );
  NAND3_X1 U22428 ( .A1(n10962), .A2(n10960), .A3(n10955), .ZN(n10058) );
  NAND2_X1 U22429 ( .A1(n9856), .A2(n9855), .ZN(n9857) );
  OAI22_X1 U22430 ( .A1(n13233), .A2(n9860), .B1(n10956), .B2(n10055), .ZN(
        n9861) );
  NAND2_X1 U22432 ( .A1(n13233), .A2(n10962), .ZN(n10050) );
  NAND2_X1 U22433 ( .A1(n9864), .A2(n10957), .ZN(n9865) );
  NAND2_X1 U22434 ( .A1(n13933), .A2(n13947), .ZN(n9869) );
  NAND2_X1 U22436 ( .A1(n2173), .A2(n51656), .ZN(n13932) );
  NAND2_X1 U22437 ( .A1(n52185), .A2(n9914), .ZN(n9871) );
  NOR2_X1 U22438 ( .A1(n9921), .A2(n9871), .ZN(n10624) );
  INV_X1 U22439 ( .A(n10624), .ZN(n9872) );
  NOR2_X1 U22440 ( .A1(n9874), .A2(n10065), .ZN(n10078) );
  INV_X1 U22441 ( .A(n10078), .ZN(n9875) );
  OAI22_X1 U22442 ( .A1(n9875), .A2(n10601), .B1(n10610), .B2(n9921), .ZN(
        n9876) );
  NAND2_X1 U22443 ( .A1(n9876), .A2(n10072), .ZN(n9882) );
  INV_X1 U22444 ( .A(n10064), .ZN(n10604) );
  NAND3_X1 U22445 ( .A1(n10605), .A2(n52185), .A3(n10604), .ZN(n9877) );
  AND2_X1 U22446 ( .A1(n10615), .A2(n9877), .ZN(n9881) );
  OAI21_X1 U22447 ( .B1(n9918), .B2(n10069), .A(n9906), .ZN(n9879) );
  NAND2_X1 U22448 ( .A1(n9879), .A2(n9878), .ZN(n9880) );
  NAND2_X1 U22449 ( .A1(n638), .A2(n13930), .ZN(n11759) );
  AOI22_X1 U22450 ( .A1(n9883), .A2(n13206), .B1(n13941), .B2(n11759), .ZN(
        n14836) );
  INV_X1 U22451 ( .A(n51655), .ZN(n13949) );
  NAND4_X1 U22452 ( .A1(n13934), .A2(n13207), .A3(n13947), .A4(n2173), .ZN(
        n9887) );
  NAND3_X1 U22453 ( .A1(n11865), .A2(n6668), .A3(n11862), .ZN(n9886) );
  NAND3_X1 U22454 ( .A1(n13941), .A2(n13947), .A3(n13948), .ZN(n9885) );
  NAND3_X1 U22455 ( .A1(n11862), .A2(n13206), .A3(n13947), .ZN(n9884) );
  NAND2_X1 U22456 ( .A1(n11610), .A2(n11591), .ZN(n10819) );
  NAND3_X1 U22457 ( .A1(n9888), .A2(n11613), .A3(n9895), .ZN(n9889) );
  OAI211_X1 U22458 ( .C1(n9890), .C2(n11612), .A(n10819), .B(n9889), .ZN(n9891) );
  INV_X1 U22459 ( .A(n9891), .ZN(n9904) );
  OAI211_X1 U22460 ( .C1(n9893), .C2(n11598), .A(n11596), .B(n9892), .ZN(n9894) );
  NAND2_X1 U22461 ( .A1(n9894), .A2(n11593), .ZN(n9903) );
  NAND2_X1 U22462 ( .A1(n11596), .A2(n9895), .ZN(n9899) );
  INV_X1 U22463 ( .A(n9896), .ZN(n9897) );
  NAND2_X1 U22464 ( .A1(n9897), .A2(n11244), .ZN(n9898) );
  NAND4_X1 U22465 ( .A1(n9899), .A2(n11590), .A3(n9898), .A4(n11604), .ZN(
        n9902) );
  NAND2_X1 U22466 ( .A1(n10814), .A2(n9900), .ZN(n9901) );
  NAND4_X2 U22467 ( .A1(n9903), .A2(n9904), .A3(n9902), .A4(n9901), .ZN(n12893) );
  INV_X1 U22468 ( .A(n10618), .ZN(n9905) );
  NAND2_X1 U22469 ( .A1(n9908), .A2(n9905), .ZN(n9913) );
  NAND2_X1 U22470 ( .A1(n10068), .A2(n10077), .ZN(n10073) );
  OAI22_X1 U22471 ( .A1(n10601), .A2(n10070), .B1(n9906), .B2(n10073), .ZN(
        n9912) );
  AND2_X1 U22472 ( .A1(n9914), .A2(n10617), .ZN(n9922) );
  NAND2_X1 U22473 ( .A1(n9910), .A2(n9909), .ZN(n9911) );
  AOI21_X1 U22474 ( .B1(n9913), .B2(n9912), .A(n9911), .ZN(n9925) );
  NOR2_X1 U22475 ( .A1(n10064), .A2(n10617), .ZN(n10602) );
  INV_X1 U22476 ( .A(n10602), .ZN(n9917) );
  OAI22_X1 U22477 ( .A1(n10601), .A2(n10616), .B1(n9921), .B2(n10074), .ZN(
        n9919) );
  NAND2_X1 U22479 ( .A1(n11709), .A2(n11200), .ZN(n9931) );
  NAND2_X1 U22480 ( .A1(n11705), .A2(n11704), .ZN(n11701) );
  INV_X1 U22481 ( .A(n11701), .ZN(n9928) );
  OAI21_X1 U22482 ( .B1(n9928), .B2(n9927), .A(n9926), .ZN(n9929) );
  OAI21_X1 U22483 ( .B1(n11705), .B2(n791), .A(n9929), .ZN(n9930) );
  MUX2_X1 U22484 ( .A(n9931), .B(n9930), .S(n11697), .Z(n9938) );
  NAND2_X1 U22487 ( .A1(n9938), .A2(n9937), .ZN(n12788) );
  NAND2_X1 U22488 ( .A1(n11655), .A2(n7185), .ZN(n9940) );
  AOI21_X1 U22489 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(n9950) );
  OAI21_X1 U22490 ( .B1(n10572), .B2(n11662), .A(n11650), .ZN(n9942) );
  INV_X1 U22491 ( .A(n9943), .ZN(n9947) );
  NAND3_X1 U22492 ( .A1(n11654), .A2(n11644), .A3(n11662), .ZN(n9945) );
  NAND4_X1 U22493 ( .A1(n9948), .A2(n9947), .A3(n9946), .A4(n9945), .ZN(n9949)
         );
  AND2_X1 U22494 ( .A1(n12894), .A2(n12790), .ZN(n13995) );
  INV_X1 U22495 ( .A(n12788), .ZN(n12794) );
  INV_X1 U22496 ( .A(n9954), .ZN(n9955) );
  NAND3_X1 U22497 ( .A1(n10184), .A2(n9955), .A3(n10178), .ZN(n9957) );
  NAND3_X1 U22498 ( .A1(n10548), .A2(n10037), .A3(n10540), .ZN(n9956) );
  NOR2_X1 U22500 ( .A1(n9959), .A2(n9958), .ZN(n9967) );
  NOR2_X1 U22501 ( .A1(n9960), .A2(n10554), .ZN(n9962) );
  INV_X1 U22502 ( .A(n10551), .ZN(n10041) );
  AOI22_X1 U22503 ( .A1(n9962), .A2(n9961), .B1(n10041), .B2(n10541), .ZN(
        n9966) );
  INV_X1 U22504 ( .A(n10174), .ZN(n10036) );
  NOR2_X1 U22505 ( .A1(n10036), .A2(n10536), .ZN(n9963) );
  NAND2_X1 U22506 ( .A1(n10042), .A2(n9963), .ZN(n9965) );
  NOR2_X1 U22507 ( .A1(n12794), .A2(n483), .ZN(n14655) );
  INV_X1 U22508 ( .A(n14655), .ZN(n13440) );
  NOR2_X1 U22509 ( .A1(n12894), .A2(n13432), .ZN(n12888) );
  INV_X1 U22510 ( .A(n12888), .ZN(n9968) );
  NAND2_X1 U22511 ( .A1(n13440), .A2(n9968), .ZN(n9989) );
  INV_X1 U22512 ( .A(n9974), .ZN(n11685) );
  NAND3_X1 U22513 ( .A1(n11669), .A2(n9969), .A3(n9337), .ZN(n10595) );
  INV_X1 U22514 ( .A(n10595), .ZN(n9972) );
  NOR2_X1 U22515 ( .A1(n11272), .A2(n9341), .ZN(n9971) );
  OAI22_X1 U22516 ( .A1(n9972), .A2(n9971), .B1(n11673), .B2(n9970), .ZN(n9978) );
  NAND3_X1 U22517 ( .A1(n11682), .A2(n11687), .A3(n9974), .ZN(n9977) );
  INV_X1 U22518 ( .A(n11681), .ZN(n9975) );
  NAND2_X1 U22519 ( .A1(n9975), .A2(n11683), .ZN(n9976) );
  NAND4_X1 U22520 ( .A1(n9979), .A2(n9978), .A3(n9977), .A4(n9976), .ZN(n9988)
         );
  OAI22_X1 U22521 ( .A1(n10590), .A2(n11280), .B1(n9980), .B2(n9341), .ZN(
        n9982) );
  NAND2_X1 U22522 ( .A1(n9982), .A2(n9981), .ZN(n9986) );
  INV_X1 U22523 ( .A(n11673), .ZN(n9983) );
  NAND2_X1 U22524 ( .A1(n9983), .A2(n11279), .ZN(n9984) );
  OAI211_X1 U22525 ( .C1(n11670), .C2(n11683), .A(n9984), .B(n9341), .ZN(n9985) );
  AOI22_X1 U22526 ( .A1(n13996), .A2(n13995), .B1(n9989), .B2(n13450), .ZN(
        n9995) );
  INV_X1 U22528 ( .A(n13994), .ZN(n9994) );
  AND2_X1 U22529 ( .A1(n12794), .A2(n12893), .ZN(n13434) );
  NOR2_X1 U22530 ( .A1(n12787), .A2(n12893), .ZN(n12792) );
  AND2_X1 U22531 ( .A1(n13449), .A2(n12787), .ZN(n11752) );
  NAND3_X1 U22532 ( .A1(n11752), .A2(n12894), .A3(n483), .ZN(n9990) );
  AND2_X1 U22533 ( .A1(n9991), .A2(n9990), .ZN(n13998) );
  NAND2_X1 U22534 ( .A1(n2072), .A2(n13449), .ZN(n13438) );
  NAND2_X1 U22535 ( .A1(n4383), .A2(n12894), .ZN(n12037) );
  OAI211_X1 U22536 ( .C1(n13434), .C2(n13432), .A(n13436), .B(n12037), .ZN(
        n9992) );
  NAND2_X1 U22537 ( .A1(n9992), .A2(n483), .ZN(n14000) );
  OAI211_X1 U22538 ( .C1(n9995), .C2(n9994), .A(n9993), .B(n14000), .ZN(n9996)
         );
  NAND2_X1 U22539 ( .A1(n11035), .A2(n10004), .ZN(n10005) );
  NAND2_X1 U22540 ( .A1(n9997), .A2(n10003), .ZN(n9999) );
  INV_X1 U22541 ( .A(n10005), .ZN(n11022) );
  NAND3_X1 U22542 ( .A1(n11022), .A2(n11037), .A3(n10579), .ZN(n10001) );
  OR2_X1 U22543 ( .A1(n10003), .A2(n10002), .ZN(n11033) );
  NAND2_X1 U22545 ( .A1(n10007), .A2(n10159), .ZN(n10088) );
  OR2_X1 U22546 ( .A1(n10578), .A2(n10162), .ZN(n10157) );
  NAND4_X1 U22548 ( .A1(n580), .A2(n10008), .A3(n8639), .A4(n10580), .ZN(
        n10009) );
  OAI211_X1 U22549 ( .C1(n10157), .C2(n11030), .A(n10010), .B(n10009), .ZN(
        n10011) );
  OAI21_X1 U22550 ( .B1(n10566), .B2(n7185), .A(n11647), .ZN(n10014) );
  AOI22_X1 U22551 ( .A1(n10014), .A2(n11655), .B1(n11648), .B2(n11650), .ZN(
        n10025) );
  OAI21_X1 U22552 ( .B1(n10562), .B2(n11660), .A(n11641), .ZN(n10017) );
  NAND2_X1 U22553 ( .A1(n7185), .A2(n11662), .ZN(n10016) );
  OAI211_X1 U22554 ( .C1(n9507), .C2(n10017), .A(n11654), .B(n10016), .ZN(
        n10023) );
  INV_X1 U22555 ( .A(n10018), .ZN(n10019) );
  NAND3_X1 U22556 ( .A1(n11647), .A2(n10019), .A3(n11662), .ZN(n10021) );
  INV_X1 U22557 ( .A(n11655), .ZN(n10020) );
  NAND4_X1 U22558 ( .A1(n10021), .A2(n10020), .A3(n11663), .A4(n5917), .ZN(
        n10022) );
  AOI21_X1 U22559 ( .B1(n10096), .B2(n10026), .A(n10101), .ZN(n10029) );
  NAND3_X1 U22560 ( .A1(n10520), .A2(n10109), .A3(n10031), .ZN(n10028) );
  NAND3_X1 U22561 ( .A1(n10532), .A2(n9482), .A3(n10110), .ZN(n10027) );
  OAI211_X1 U22562 ( .C1(n10029), .C2(n10097), .A(n10028), .B(n10027), .ZN(
        n10030) );
  NAND2_X1 U22563 ( .A1(n10031), .A2(n9482), .ZN(n10531) );
  MUX2_X1 U22564 ( .A(n10032), .B(n8853), .S(n10096), .Z(n10035) );
  NAND3_X1 U22565 ( .A1(n10033), .A2(n10109), .A3(n10111), .ZN(n10034) );
  NAND2_X1 U22566 ( .A1(n10174), .A2(n10546), .ZN(n10040) );
  NAND4_X1 U22567 ( .A1(n10038), .A2(n10037), .A3(n10036), .A4(n10547), .ZN(
        n10039) );
  INV_X1 U22568 ( .A(n10555), .ZN(n10549) );
  NAND3_X1 U22569 ( .A1(n10047), .A2(n10955), .A3(n10127), .ZN(n10049) );
  NAND3_X1 U22570 ( .A1(n10960), .A2(n10054), .A3(n10961), .ZN(n10048) );
  NAND4_X1 U22571 ( .A1(n10051), .A2(n10050), .A3(n10049), .A4(n10048), .ZN(
        n10062) );
  AND2_X1 U22572 ( .A1(n10122), .A2(n10124), .ZN(n10966) );
  AND2_X1 U22573 ( .A1(n10052), .A2(n10967), .ZN(n10053) );
  OAI21_X1 U22574 ( .B1(n10055), .B2(n10122), .A(n3316), .ZN(n10056) );
  OAI21_X1 U22575 ( .B1(n10962), .B2(n10056), .A(n10964), .ZN(n10057) );
  NAND4_X1 U22576 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n10061) );
  XNOR2_X1 U22578 ( .A(n10905), .B(n13780), .ZN(n10063) );
  AND2_X1 U22579 ( .A1(n13782), .A2(n10901), .ZN(n10082) );
  NOR2_X1 U22580 ( .A1(n10610), .A2(n10064), .ZN(n10067) );
  OAI21_X1 U22581 ( .B1(n10617), .B2(n10065), .A(n10070), .ZN(n10066) );
  AOI22_X1 U22582 ( .A1(n10067), .A2(n10609), .B1(n10066), .B2(n10610), .ZN(
        n10081) );
  NAND4_X1 U22583 ( .A1(n10068), .A2(n10074), .A3(n10607), .A4(n10077), .ZN(
        n10071) );
  MUX2_X1 U22584 ( .A(n10071), .B(n10070), .S(n10069), .Z(n10080) );
  NAND3_X1 U22585 ( .A1(n10619), .A2(n10072), .A3(n10610), .ZN(n10076) );
  NAND3_X1 U22586 ( .A1(n10619), .A2(n10074), .A3(n10073), .ZN(n10075) );
  NAND2_X1 U22587 ( .A1(n10078), .A2(n10077), .ZN(n10079) );
  OAI21_X1 U22588 ( .B1(n10083), .B2(n10082), .A(n13779), .ZN(n10092) );
  NAND2_X1 U22589 ( .A1(n12419), .A2(n13173), .ZN(n12017) );
  NAND2_X1 U22590 ( .A1(n10905), .A2(n13779), .ZN(n13773) );
  OAI21_X1 U22591 ( .B1(n10905), .B2(n12017), .A(n13773), .ZN(n10085) );
  OAI21_X1 U22592 ( .B1(n13172), .B2(n13173), .A(n13174), .ZN(n10084) );
  NOR2_X1 U22593 ( .A1(n10085), .A2(n10084), .ZN(n10087) );
  OR2_X1 U22594 ( .A1(n13782), .A2(n13172), .ZN(n12424) );
  NAND2_X1 U22595 ( .A1(n13172), .A2(n13779), .ZN(n10906) );
  INV_X1 U22596 ( .A(n10906), .ZN(n10086) );
  AOI22_X1 U22597 ( .A1(n10087), .A2(n12424), .B1(n13161), .B2(n10086), .ZN(
        n10091) );
  AOI21_X1 U22598 ( .B1(n10899), .B2(n10898), .A(n13170), .ZN(n13179) );
  INV_X1 U22599 ( .A(n13179), .ZN(n12013) );
  INV_X1 U22600 ( .A(n13774), .ZN(n13169) );
  INV_X1 U22601 ( .A(n13178), .ZN(n10089) );
  OR2_X1 U22602 ( .A1(n12416), .A2(n10089), .ZN(n13187) );
  INV_X1 U22603 ( .A(n17648), .ZN(n10093) );
  XNOR2_X1 U22604 ( .A(n10094), .B(n10093), .ZN(n10658) );
  INV_X1 U22605 ( .A(n10097), .ZN(n10095) );
  NAND2_X1 U22606 ( .A1(n10097), .A2(n10096), .ZN(n10098) );
  NAND2_X1 U22608 ( .A1(n10101), .A2(n9482), .ZN(n10102) );
  NAND2_X1 U22609 ( .A1(n10103), .A2(n10102), .ZN(n10117) );
  NAND2_X1 U22610 ( .A1(n10107), .A2(n10106), .ZN(n10115) );
  NAND2_X1 U22611 ( .A1(n10108), .A2(n10530), .ZN(n10114) );
  OAI22_X1 U22612 ( .A1(n10526), .A2(n10508), .B1(n10110), .B2(n10109), .ZN(
        n10112) );
  OAI21_X1 U22613 ( .B1(n10968), .B2(n10122), .A(n6004), .ZN(n10118) );
  AND2_X1 U22614 ( .A1(n10119), .A2(n10118), .ZN(n10133) );
  NOR2_X1 U22615 ( .A1(n10121), .A2(n10120), .ZN(n10123) );
  AOI22_X1 U22616 ( .A1(n10960), .A2(n10123), .B1(n10968), .B2(n10122), .ZN(
        n10131) );
  NAND3_X1 U22617 ( .A1(n10125), .A2(n10124), .A3(n10955), .ZN(n10130) );
  AND2_X1 U22618 ( .A1(n13135), .A2(n51136), .ZN(n10172) );
  NAND2_X1 U22619 ( .A1(n10222), .A2(n10134), .ZN(n10136) );
  NAND2_X1 U22620 ( .A1(n10219), .A2(n10142), .ZN(n10146) );
  NAND3_X1 U22621 ( .A1(n10144), .A2(n10931), .A3(n10143), .ZN(n10145) );
  MUX2_X1 U22622 ( .A(n10146), .B(n10145), .S(n10218), .Z(n10155) );
  NOR2_X1 U22623 ( .A1(n10215), .A2(n10147), .ZN(n10150) );
  NOR2_X1 U22624 ( .A1(n10217), .A2(n10148), .ZN(n10149) );
  INV_X1 U22625 ( .A(n10219), .ZN(n10151) );
  MUX2_X1 U22626 ( .A(n10924), .B(n10218), .S(n10151), .Z(n10152) );
  NAND2_X1 U22627 ( .A1(n10152), .A2(n10926), .ZN(n10153) );
  NAND2_X1 U22629 ( .A1(n10575), .A2(n8639), .ZN(n10158) );
  OAI21_X1 U22630 ( .B1(n2197), .B2(n10575), .A(n10158), .ZN(n10160) );
  NAND2_X1 U22631 ( .A1(n10160), .A2(n10159), .ZN(n10168) );
  OAI21_X1 U22632 ( .B1(n11036), .B2(n10161), .A(n11030), .ZN(n10164) );
  NOR2_X1 U22633 ( .A1(n11031), .A2(n11035), .ZN(n10163) );
  OAI211_X1 U22634 ( .C1(n10164), .C2(n10163), .A(n10162), .B(n10578), .ZN(
        n10167) );
  NAND2_X1 U22635 ( .A1(n10165), .A2(n11037), .ZN(n10166) );
  NAND3_X1 U22636 ( .A1(n10172), .A2(n6609), .A3(n13148), .ZN(n10191) );
  NAND2_X1 U22637 ( .A1(n10172), .A2(n13136), .ZN(n10190) );
  NAND3_X1 U22638 ( .A1(n10551), .A2(n10173), .A3(n10179), .ZN(n10176) );
  NAND3_X1 U22639 ( .A1(n10541), .A2(n10174), .A3(n10178), .ZN(n10175) );
  NAND4_X1 U22640 ( .A1(n10177), .A2(n10184), .A3(n3850), .A4(n10178), .ZN(
        n10181) );
  NAND3_X1 U22641 ( .A1(n10541), .A2(n10179), .A3(n10178), .ZN(n10180) );
  INV_X1 U22642 ( .A(n10182), .ZN(n10185) );
  NOR2_X1 U22643 ( .A1(n10552), .A2(n9461), .ZN(n10183) );
  AOI22_X1 U22644 ( .A1(n10185), .A2(n10555), .B1(n10184), .B2(n10183), .ZN(
        n10189) );
  NOR3_X1 U22645 ( .A1(n10186), .A2(n10540), .A3(n9461), .ZN(n10187) );
  MUX2_X1 U22646 ( .A(n10191), .B(n10190), .S(n13142), .Z(n10212) );
  NAND2_X1 U22647 ( .A1(n10247), .A2(n10192), .ZN(n10197) );
  AND2_X1 U22648 ( .A1(n10240), .A2(n11015), .ZN(n10193) );
  NOR2_X1 U22649 ( .A1(n11008), .A2(n10193), .ZN(n10196) );
  AND2_X1 U22650 ( .A1(n10199), .A2(n11015), .ZN(n10241) );
  NOR2_X1 U22652 ( .A1(n10201), .A2(n7936), .ZN(n11002) );
  OAI21_X1 U22653 ( .B1(n11002), .B2(n11014), .A(n2704), .ZN(n10202) );
  NAND2_X1 U22654 ( .A1(n12907), .A2(n13142), .ZN(n14183) );
  NAND2_X1 U22655 ( .A1(n12907), .A2(n51136), .ZN(n13143) );
  OAI22_X1 U22656 ( .A1(n14178), .A2(n14183), .B1(n13143), .B2(n10204), .ZN(
        n10207) );
  OAI21_X1 U22657 ( .B1(n51136), .B2(n12907), .A(n14179), .ZN(n10205) );
  NAND2_X1 U22658 ( .A1(n13136), .A2(n14178), .ZN(n11172) );
  NOR2_X1 U22659 ( .A1(n10205), .A2(n11172), .ZN(n10206) );
  NOR2_X1 U22660 ( .A1(n10207), .A2(n10206), .ZN(n10211) );
  AND2_X1 U22661 ( .A1(n14178), .A2(n12907), .ZN(n12217) );
  INV_X1 U22662 ( .A(n12217), .ZN(n13130) );
  AND2_X1 U22663 ( .A1(n51136), .A2(n14186), .ZN(n12213) );
  NAND3_X1 U22665 ( .A1(n13139), .A2(n13152), .A3(n14179), .ZN(n10209) );
  NAND2_X1 U22666 ( .A1(n10926), .A2(n52188), .ZN(n10929) );
  OAI211_X1 U22667 ( .C1(n10926), .C2(n10920), .A(n10222), .B(n10218), .ZN(
        n10213) );
  NAND2_X1 U22668 ( .A1(n10217), .A2(n10223), .ZN(n10220) );
  NAND3_X1 U22669 ( .A1(n10222), .A2(n52188), .A3(n10221), .ZN(n10917) );
  INV_X1 U22670 ( .A(n10223), .ZN(n10923) );
  INV_X1 U22671 ( .A(n10225), .ZN(n10228) );
  NAND2_X1 U22672 ( .A1(n12294), .A2(n12282), .ZN(n10718) );
  OAI22_X1 U22673 ( .A1(n12276), .A2(n12286), .B1(n10718), .B2(n10226), .ZN(
        n10227) );
  AOI21_X1 U22674 ( .B1(n10229), .B2(n10228), .A(n10227), .ZN(n10238) );
  INV_X1 U22675 ( .A(n10715), .ZN(n12293) );
  NAND3_X1 U22676 ( .A1(n10723), .A2(n12293), .A3(n10234), .ZN(n10237) );
  NAND3_X1 U22677 ( .A1(n10723), .A2(n10235), .A3(n12290), .ZN(n10236) );
  AND3_X1 U22678 ( .A1(n11011), .A2(n10240), .A3(n51762), .ZN(n10243) );
  INV_X1 U22679 ( .A(n10241), .ZN(n10242) );
  AOI22_X1 U22680 ( .A1(n10244), .A2(n11004), .B1(n10243), .B2(n10242), .ZN(
        n10249) );
  NAND3_X1 U22681 ( .A1(n10247), .A2(n10246), .A3(n10245), .ZN(n10248) );
  NAND2_X1 U22682 ( .A1(n10251), .A2(n10250), .ZN(n10254) );
  AND2_X1 U22683 ( .A1(n10252), .A2(n11015), .ZN(n10253) );
  AOI21_X1 U22684 ( .B1(n10255), .B2(n10254), .A(n10253), .ZN(n10256) );
  INV_X1 U22685 ( .A(n10984), .ZN(n10257) );
  AOI22_X1 U22686 ( .A1(n10258), .A2(n10272), .B1(n10257), .B2(n10976), .ZN(
        n10276) );
  NAND2_X1 U22687 ( .A1(n10259), .A2(n8796), .ZN(n12353) );
  NAND3_X1 U22688 ( .A1(n12363), .A2(n10988), .A3(n9782), .ZN(n10260) );
  OAI21_X1 U22689 ( .B1(n10262), .B2(n10261), .A(n51137), .ZN(n10263) );
  OAI211_X1 U22690 ( .C1(n10976), .C2(n51137), .A(n10263), .B(n10272), .ZN(
        n10271) );
  INV_X1 U22691 ( .A(n10989), .ZN(n10270) );
  INV_X1 U22692 ( .A(n10265), .ZN(n10266) );
  OAI211_X1 U22693 ( .C1(n10268), .C2(n10267), .A(n10266), .B(n8791), .ZN(
        n10269) );
  AND3_X1 U22694 ( .A1(n10271), .A2(n10270), .A3(n10269), .ZN(n10275) );
  OAI21_X1 U22695 ( .B1(n10990), .B2(n10272), .A(n12351), .ZN(n10273) );
  NAND2_X1 U22696 ( .A1(n10273), .A2(n8796), .ZN(n10274) );
  INV_X1 U22698 ( .A(n12344), .ZN(n10667) );
  INV_X1 U22699 ( .A(n10281), .ZN(n10284) );
  OAI21_X1 U22700 ( .B1(n51194), .B2(n12337), .A(n10285), .ZN(n10283) );
  OAI22_X1 U22701 ( .A1(n10286), .A2(n10285), .B1(n10279), .B2(n12337), .ZN(
        n10287) );
  INV_X1 U22703 ( .A(n12331), .ZN(n10290) );
  OAI21_X1 U22704 ( .B1(n10290), .B2(n10289), .A(n10672), .ZN(n10291) );
  INV_X1 U22705 ( .A(n10292), .ZN(n10295) );
  NAND2_X1 U22706 ( .A1(n10293), .A2(n9656), .ZN(n10294) );
  OAI211_X1 U22707 ( .C1(n10938), .C2(n10295), .A(n10294), .B(n12301), .ZN(
        n10301) );
  INV_X1 U22708 ( .A(n9758), .ZN(n10298) );
  AND2_X1 U22709 ( .A1(n10296), .A2(n12315), .ZN(n10297) );
  OAI21_X1 U22710 ( .B1(n10298), .B2(n10297), .A(n12317), .ZN(n10299) );
  NAND3_X1 U22711 ( .A1(n10301), .A2(n10300), .A3(n10299), .ZN(n10309) );
  AOI21_X1 U22712 ( .B1(n12301), .B2(n12313), .A(n12314), .ZN(n10306) );
  INV_X1 U22713 ( .A(n12299), .ZN(n10942) );
  NAND3_X1 U22714 ( .A1(n10942), .A2(n10951), .A3(n10302), .ZN(n10305) );
  INV_X1 U22715 ( .A(n10303), .ZN(n10304) );
  OAI211_X1 U22716 ( .C1(n10306), .C2(n12300), .A(n10305), .B(n10304), .ZN(
        n10307) );
  INV_X1 U22717 ( .A(n10307), .ZN(n10308) );
  NAND2_X1 U22718 ( .A1(n10309), .A2(n10308), .ZN(n13761) );
  NAND2_X1 U22719 ( .A1(n14149), .A2(n51175), .ZN(n14967) );
  INV_X1 U22720 ( .A(n14145), .ZN(n13114) );
  INV_X1 U22722 ( .A(n13762), .ZN(n10775) );
  NAND3_X1 U22723 ( .A1(n10775), .A2(n14160), .A3(n13761), .ZN(n10310) );
  XNOR2_X1 U22724 ( .A(n4461), .B(n14160), .ZN(n10312) );
  NAND3_X1 U22725 ( .A1(n10313), .A2(n14159), .A3(n14966), .ZN(n10314) );
  MUX2_X1 U22726 ( .A(n12617), .B(n12638), .S(n12071), .Z(n12080) );
  NAND2_X1 U22727 ( .A1(n12080), .A2(n12628), .ZN(n10318) );
  NOR2_X1 U22728 ( .A1(n12071), .A2(n12638), .ZN(n12075) );
  AOI21_X1 U22729 ( .B1(n12617), .B2(n12616), .A(n3347), .ZN(n10316) );
  OAI21_X1 U22730 ( .B1(n12075), .B2(n10316), .A(n10465), .ZN(n10317) );
  OAI22_X1 U22731 ( .A1(n12618), .A2(n12617), .B1(n12616), .B2(n12066), .ZN(
        n10320) );
  OAI211_X1 U22732 ( .C1(n10320), .C2(n10319), .A(n9208), .B(n12619), .ZN(
        n10325) );
  OAI21_X1 U22733 ( .B1(n12638), .B2(n12619), .A(n9208), .ZN(n10321) );
  NAND2_X1 U22734 ( .A1(n10321), .A2(n10462), .ZN(n10324) );
  INV_X1 U22735 ( .A(n12618), .ZN(n10467) );
  OAI211_X1 U22737 ( .C1(n548), .C2(n10328), .A(n11325), .B(n12179), .ZN(
        n10332) );
  NAND3_X1 U22738 ( .A1(n12178), .A2(n10333), .A3(n10413), .ZN(n10331) );
  NAND3_X1 U22739 ( .A1(n10418), .A2(n12173), .A3(n12175), .ZN(n10330) );
  NAND2_X1 U22740 ( .A1(n548), .A2(n10328), .ZN(n10329) );
  NAND4_X1 U22741 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10337) );
  NAND2_X1 U22742 ( .A1(n11328), .A2(n12173), .ZN(n12159) );
  NAND3_X1 U22743 ( .A1(n12159), .A2(n12160), .A3(n12169), .ZN(n10335) );
  AND2_X1 U22744 ( .A1(n10333), .A2(n12173), .ZN(n11323) );
  NAND3_X1 U22745 ( .A1(n11323), .A2(n548), .A3(n12177), .ZN(n10334) );
  AOI21_X1 U22746 ( .B1(n10335), .B2(n10334), .A(n10417), .ZN(n10336) );
  OR2_X1 U22747 ( .A1(n10337), .A2(n10336), .ZN(n13804) );
  NAND2_X1 U22749 ( .A1(n10445), .A2(n10449), .ZN(n10340) );
  NAND2_X1 U22750 ( .A1(n11974), .A2(n10444), .ZN(n10339) );
  NAND2_X1 U22751 ( .A1(n10340), .A2(n10455), .ZN(n10341) );
  NAND2_X1 U22752 ( .A1(n2227), .A2(n12648), .ZN(n10343) );
  NOR2_X1 U22753 ( .A1(n11973), .A2(n10343), .ZN(n10344) );
  NAND2_X1 U22754 ( .A1(n10344), .A2(n12649), .ZN(n10352) );
  NAND2_X1 U22755 ( .A1(n10449), .A2(n11978), .ZN(n10347) );
  OAI21_X1 U22756 ( .B1(n10347), .B2(n10346), .A(n10345), .ZN(n10348) );
  INV_X1 U22757 ( .A(n10348), .ZN(n10351) );
  NAND2_X1 U22758 ( .A1(n11984), .A2(n12663), .ZN(n10349) );
  NAND2_X1 U22759 ( .A1(n10665), .A2(n10361), .ZN(n10359) );
  NAND3_X1 U22760 ( .A1(n10362), .A2(n10356), .A3(n10355), .ZN(n10357) );
  OAI22_X1 U22761 ( .A1(n10362), .A2(n12055), .B1(n10361), .B2(n10360), .ZN(
        n10363) );
  MUX2_X1 U22762 ( .A(n10364), .B(n10363), .S(n12051), .Z(n10365) );
  NAND2_X1 U22763 ( .A1(n13801), .A2(n13804), .ZN(n10381) );
  NAND2_X1 U22764 ( .A1(n10702), .A2(n11375), .ZN(n10367) );
  NOR2_X1 U22765 ( .A1(n9632), .A2(n12123), .ZN(n10369) );
  NOR2_X1 U22766 ( .A1(n10367), .A2(n9632), .ZN(n12120) );
  NAND3_X1 U22768 ( .A1(n12114), .A2(n11359), .A3(n11375), .ZN(n10371) );
  AND2_X1 U22769 ( .A1(n10372), .A2(n10371), .ZN(n10379) );
  NAND2_X1 U22770 ( .A1(n11372), .A2(n11375), .ZN(n10377) );
  NAND2_X1 U22771 ( .A1(n10699), .A2(n10695), .ZN(n10376) );
  NAND4_X1 U22772 ( .A1(n10377), .A2(n12112), .A3(n10376), .A4(n11368), .ZN(
        n10378) );
  NAND2_X1 U22773 ( .A1(n10381), .A2(n13797), .ZN(n10382) );
  OAI211_X1 U22774 ( .C1(n13798), .C2(n13801), .A(n13483), .B(n10382), .ZN(
        n10405) );
  XNOR2_X1 U22775 ( .A(n13801), .B(n13800), .ZN(n10402) );
  NAND3_X1 U22776 ( .A1(n12146), .A2(n11403), .A3(n10390), .ZN(n10389) );
  AND2_X1 U22777 ( .A1(n12137), .A2(n11410), .ZN(n10384) );
  NAND2_X1 U22778 ( .A1(n10384), .A2(n10383), .ZN(n10388) );
  NAND2_X1 U22779 ( .A1(n10384), .A2(n10392), .ZN(n10387) );
  NAND3_X1 U22780 ( .A1(n11400), .A2(n10385), .A3(n11423), .ZN(n10386) );
  NAND4_X1 U22781 ( .A1(n10389), .A2(n10388), .A3(n10387), .A4(n10386), .ZN(
        n10397) );
  NAND3_X1 U22782 ( .A1(n11400), .A2(n2105), .A3(n11410), .ZN(n10395) );
  NAND3_X1 U22783 ( .A1(n12141), .A2(n10390), .A3(n51141), .ZN(n10394) );
  OAI21_X1 U22787 ( .B1(n12138), .B2(n11410), .A(n2105), .ZN(n10399) );
  MUX2_X1 U22788 ( .A(n11398), .B(n10399), .S(n11417), .Z(n10400) );
  NAND3_X1 U22789 ( .A1(n10402), .A2(n15044), .A3(n15034), .ZN(n10404) );
  INV_X1 U22790 ( .A(n13804), .ZN(n15047) );
  NAND3_X1 U22791 ( .A1(n13475), .A2(n15047), .A3(n15044), .ZN(n10403) );
  OR2_X1 U22792 ( .A1(n13797), .A2(n15047), .ZN(n12773) );
  NOR2_X1 U22793 ( .A1(n12773), .A2(n69), .ZN(n15039) );
  INV_X1 U22794 ( .A(n15039), .ZN(n10411) );
  NAND2_X1 U22795 ( .A1(n15046), .A2(n13483), .ZN(n13805) );
  INV_X1 U22796 ( .A(n13805), .ZN(n13487) );
  NAND3_X1 U22797 ( .A1(n13487), .A2(n15048), .A3(n15030), .ZN(n10410) );
  NAND2_X1 U22798 ( .A1(n15045), .A2(n13487), .ZN(n10409) );
  NAND2_X1 U22799 ( .A1(n10407), .A2(n13798), .ZN(n10408) );
  XNOR2_X1 U22800 ( .A(n4909), .B(n4208), .ZN(n25426) );
  XNOR2_X1 U22801 ( .A(n25426), .B(n4650), .ZN(n33862) );
  XNOR2_X1 U22802 ( .A(n17118), .B(n33862), .ZN(n16029) );
  XNOR2_X1 U22803 ( .A(n16372), .B(n16029), .ZN(n10656) );
  OAI21_X1 U22804 ( .B1(n10414), .B2(n10417), .A(n12178), .ZN(n10416) );
  AND2_X1 U22805 ( .A1(n12177), .A2(n548), .ZN(n12167) );
  NAND3_X1 U22806 ( .A1(n12167), .A2(n12160), .A3(n12173), .ZN(n10415) );
  NAND2_X1 U22807 ( .A1(n12170), .A2(n12173), .ZN(n10420) );
  NOR2_X1 U22808 ( .A1(n12174), .A2(n548), .ZN(n10421) );
  NAND2_X1 U22809 ( .A1(n12728), .A2(n8881), .ZN(n12730) );
  NAND2_X1 U22810 ( .A1(n12724), .A2(n12730), .ZN(n10426) );
  AND2_X1 U22811 ( .A1(n12728), .A2(n11954), .ZN(n11946) );
  INV_X1 U22812 ( .A(n10422), .ZN(n10427) );
  OAI22_X1 U22813 ( .A1(n11943), .A2(n11109), .B1(n10427), .B2(n5484), .ZN(
        n10425) );
  AOI22_X1 U22814 ( .A1(n10426), .A2(n11946), .B1(n10425), .B2(n10424), .ZN(
        n10443) );
  AND2_X1 U22815 ( .A1(n11942), .A2(n11964), .ZN(n12718) );
  INV_X1 U22816 ( .A(n10431), .ZN(n10429) );
  INV_X1 U22817 ( .A(n11957), .ZN(n10432) );
  OAI222_X1 U22818 ( .A1(n12727), .A2(n10429), .B1(n11109), .B2(n5473), .C1(
        n10427), .C2(n10432), .ZN(n10436) );
  NAND2_X1 U22819 ( .A1(n11957), .A2(n11942), .ZN(n10430) );
  NAND3_X1 U22821 ( .A1(n10438), .A2(n12728), .A3(n10432), .ZN(n10433) );
  AOI21_X1 U22823 ( .B1(n12718), .B2(n10436), .A(n10435), .ZN(n10442) );
  INV_X1 U22824 ( .A(n10437), .ZN(n11960) );
  MUX2_X1 U22825 ( .A(n11957), .B(n11943), .S(n10438), .Z(n10440) );
  NAND2_X1 U22826 ( .A1(n10440), .A2(n10439), .ZN(n10441) );
  NOR2_X1 U22827 ( .A1(n15136), .A2(n15133), .ZN(n15139) );
  NAND2_X1 U22828 ( .A1(n10457), .A2(n9188), .ZN(n12661) );
  NAND2_X1 U22829 ( .A1(n12661), .A2(n11979), .ZN(n10446) );
  NAND4_X1 U22830 ( .A1(n10446), .A2(n12659), .A3(n10449), .A4(n11973), .ZN(
        n10448) );
  NAND4_X1 U22831 ( .A1(n12652), .A2(n10456), .A3(n12663), .A4(n12649), .ZN(
        n10447) );
  AND3_X1 U22832 ( .A1(n11977), .A2(n10448), .A3(n10447), .ZN(n10461) );
  NOR2_X1 U22833 ( .A1(n11973), .A2(n12659), .ZN(n12654) );
  NOR2_X1 U22834 ( .A1(n10449), .A2(n12659), .ZN(n10450) );
  AOI22_X1 U22835 ( .A1(n12654), .A2(n10451), .B1(n10450), .B2(n11974), .ZN(
        n10460) );
  AND3_X1 U22836 ( .A1(n10456), .A2(n9188), .A3(n12649), .ZN(n10454) );
  NOR2_X1 U22837 ( .A1(n11986), .A2(n12649), .ZN(n10453) );
  INV_X1 U22838 ( .A(n11973), .ZN(n10452) );
  AOI21_X1 U22840 ( .B1(n10465), .B2(n51433), .A(n12630), .ZN(n10466) );
  AOI22_X1 U22841 ( .A1(n10467), .A2(n10466), .B1(n12628), .B2(n12631), .ZN(
        n10470) );
  NAND3_X1 U22843 ( .A1(n10472), .A2(n10474), .A3(n9539), .ZN(n10484) );
  OAI21_X1 U22844 ( .B1(n10474), .B2(n3377), .A(n12602), .ZN(n10475) );
  NAND2_X1 U22845 ( .A1(n51140), .A2(n52140), .ZN(n10476) );
  AND3_X1 U22846 ( .A1(n10478), .A2(n10477), .A3(n10476), .ZN(n10483) );
  NAND2_X1 U22847 ( .A1(n12596), .A2(n357), .ZN(n10479) );
  NAND3_X1 U22848 ( .A1(n11922), .A2(n11137), .A3(n10479), .ZN(n10482) );
  AND2_X1 U22849 ( .A1(n52140), .A2(n357), .ZN(n11912) );
  NAND2_X1 U22850 ( .A1(n10480), .A2(n11912), .ZN(n10481) );
  NAND3_X1 U22851 ( .A1(n10487), .A2(n12696), .A3(n12710), .ZN(n12439) );
  NAND4_X1 U22852 ( .A1(n12435), .A2(n11933), .A3(n12695), .A4(n12709), .ZN(
        n10486) );
  AND2_X1 U22853 ( .A1(n12700), .A2(n11931), .ZN(n11930) );
  NAND3_X1 U22854 ( .A1(n11930), .A2(n802), .A3(n12709), .ZN(n10485) );
  AND3_X1 U22855 ( .A1(n10486), .A2(n12439), .A3(n10485), .ZN(n10497) );
  INV_X1 U22856 ( .A(n10487), .ZN(n12713) );
  NOR2_X1 U22857 ( .A1(n12713), .A2(n12690), .ZN(n12436) );
  OAI21_X1 U22858 ( .B1(n12436), .B2(n12701), .A(n12441), .ZN(n10496) );
  NOR2_X1 U22859 ( .A1(n12713), .A2(n802), .ZN(n11926) );
  INV_X1 U22860 ( .A(n12699), .ZN(n10488) );
  OAI21_X1 U22861 ( .B1(n11926), .B2(n12440), .A(n10488), .ZN(n10495) );
  NAND2_X1 U22862 ( .A1(n11123), .A2(n12700), .ZN(n10490) );
  OAI21_X1 U22863 ( .B1(n12700), .B2(n12702), .A(n10490), .ZN(n10489) );
  INV_X1 U22864 ( .A(n12692), .ZN(n12704) );
  NAND3_X1 U22865 ( .A1(n10489), .A2(n12704), .A3(n12709), .ZN(n10493) );
  INV_X1 U22866 ( .A(n10490), .ZN(n10491) );
  NAND3_X1 U22867 ( .A1(n10491), .A2(n12699), .A3(n12709), .ZN(n10492) );
  AND2_X1 U22868 ( .A1(n10493), .A2(n10492), .ZN(n10494) );
  NAND4_X2 U22869 ( .A1(n10497), .A2(n10496), .A3(n10494), .A4(n10495), .ZN(
        n15131) );
  OAI211_X1 U22870 ( .C1(n15136), .C2(n14260), .A(n13708), .B(n15126), .ZN(
        n10498) );
  AND2_X1 U22871 ( .A1(n15133), .A2(n14257), .ZN(n14995) );
  INV_X1 U22872 ( .A(n10499), .ZN(n15138) );
  AND2_X1 U22873 ( .A1(n15133), .A2(n15138), .ZN(n14268) );
  NAND2_X1 U22874 ( .A1(n13696), .A2(n14268), .ZN(n10505) );
  NAND2_X1 U22875 ( .A1(n13709), .A2(n15132), .ZN(n13698) );
  AOI22_X1 U22876 ( .A1(n10500), .A2(n15131), .B1(n13698), .B2(n13697), .ZN(
        n10504) );
  AND2_X1 U22877 ( .A1(n15133), .A2(n15126), .ZN(n13703) );
  INV_X1 U22878 ( .A(n10501), .ZN(n14270) );
  NAND2_X1 U22879 ( .A1(n13703), .A2(n14270), .ZN(n10503) );
  INV_X1 U22880 ( .A(n14257), .ZN(n14271) );
  NAND3_X1 U22881 ( .A1(n13711), .A2(n14271), .A3(n15136), .ZN(n10502) );
  XNOR2_X1 U22883 ( .A(n4939), .B(n4746), .ZN(n26042) );
  XNOR2_X1 U22884 ( .A(n26042), .B(n4624), .ZN(n33387) );
  XNOR2_X1 U22885 ( .A(n17117), .B(n33387), .ZN(n10655) );
  OAI211_X1 U22886 ( .C1(n10527), .C2(n10508), .A(n10507), .B(n10530), .ZN(
        n10510) );
  NAND2_X1 U22887 ( .A1(n10510), .A2(n10509), .ZN(n10512) );
  NAND2_X1 U22888 ( .A1(n10512), .A2(n10511), .ZN(n10518) );
  AOI21_X1 U22889 ( .B1(n10516), .B2(n10515), .A(n10514), .ZN(n10517) );
  NOR2_X1 U22890 ( .A1(n10518), .A2(n10517), .ZN(n10649) );
  MUX2_X1 U22891 ( .A(n10524), .B(n10523), .S(n10522), .Z(n10647) );
  NAND2_X1 U22892 ( .A1(n10649), .A2(n10647), .ZN(n10628) );
  OAI211_X1 U22895 ( .C1(n9484), .C2(n9482), .A(n10634), .B(n10633), .ZN(
        n10533) );
  OAI21_X1 U22896 ( .B1(n10532), .B2(n10531), .A(n10530), .ZN(n10648) );
  AOI21_X1 U22897 ( .B1(n10534), .B2(n10533), .A(n10648), .ZN(n10535) );
  NAND2_X1 U22898 ( .A1(n10537), .A2(n10536), .ZN(n10561) );
  NAND2_X1 U22899 ( .A1(n10555), .A2(n51761), .ZN(n10542) );
  NAND4_X1 U22900 ( .A1(n10542), .A2(n10541), .A3(n10540), .A4(n10539), .ZN(
        n10543) );
  OAI21_X1 U22901 ( .B1(n10544), .B2(n10552), .A(n10543), .ZN(n10545) );
  INV_X1 U22902 ( .A(n10545), .ZN(n10560) );
  NOR2_X1 U22903 ( .A1(n10547), .A2(n10546), .ZN(n10550) );
  AOI22_X1 U22904 ( .A1(n10551), .A2(n10550), .B1(n10549), .B2(n10548), .ZN(
        n10559) );
  NAND3_X1 U22905 ( .A1(n10554), .A2(n10552), .A3(n9461), .ZN(n10553) );
  OAI21_X1 U22906 ( .B1(n10555), .B2(n10554), .A(n10553), .ZN(n10557) );
  NAND2_X1 U22907 ( .A1(n10557), .A2(n10556), .ZN(n10558) );
  AOI21_X1 U22908 ( .B1(n10563), .B2(n7185), .A(n10562), .ZN(n10564) );
  AOI22_X1 U22909 ( .A1(n11654), .A2(n10564), .B1(n11655), .B2(n10566), .ZN(
        n10568) );
  OAI211_X1 U22910 ( .C1(n10566), .C2(n11641), .A(n10565), .B(n11650), .ZN(
        n10567) );
  OAI211_X1 U22911 ( .C1(n10569), .C2(n11644), .A(n10568), .B(n10567), .ZN(
        n10574) );
  NAND2_X1 U22912 ( .A1(n14339), .A2(n13417), .ZN(n14330) );
  NAND3_X1 U22913 ( .A1(n11025), .A2(n10575), .A3(n10578), .ZN(n10576) );
  NAND3_X1 U22914 ( .A1(n10579), .A2(n8639), .A3(n11035), .ZN(n10583) );
  NAND3_X1 U22915 ( .A1(n10581), .A2(n11027), .A3(n10580), .ZN(n10582) );
  NOR2_X1 U22916 ( .A1(n10587), .A2(n11272), .ZN(n10588) );
  OAI21_X1 U22917 ( .B1(n11676), .B2(n10588), .A(n11269), .ZN(n10600) );
  OAI211_X1 U22918 ( .C1(n10590), .C2(n11275), .A(n10589), .B(n9341), .ZN(
        n10592) );
  NOR2_X1 U22919 ( .A1(n10592), .A2(n10591), .ZN(n10593) );
  OAI21_X1 U22920 ( .B1(n11676), .B2(n10594), .A(n10593), .ZN(n10599) );
  NAND2_X1 U22921 ( .A1(n11688), .A2(n11683), .ZN(n10596) );
  NAND3_X1 U22922 ( .A1(n11269), .A2(n11669), .A3(n11268), .ZN(n10598) );
  NAND3_X1 U22923 ( .A1(n11270), .A2(n11688), .A3(n11268), .ZN(n10597) );
  NAND2_X1 U22924 ( .A1(n14331), .A2(n14341), .ZN(n13008) );
  AOI22_X1 U22925 ( .A1(n10604), .A2(n10603), .B1(n10602), .B2(n10601), .ZN(
        n10627) );
  NAND2_X1 U22926 ( .A1(n10605), .A2(n52185), .ZN(n10614) );
  NAND4_X1 U22927 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10613) );
  NAND3_X1 U22928 ( .A1(n10611), .A2(n10610), .A3(n10617), .ZN(n10612) );
  AND4_X1 U22929 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(
        n10626) );
  OAI21_X1 U22930 ( .B1(n10616), .B2(n10618), .A(n10617), .ZN(n10623) );
  OAI21_X1 U22933 ( .B1(n10624), .B2(n10623), .A(n10622), .ZN(n10625) );
  INV_X1 U22934 ( .A(n10628), .ZN(n10646) );
  INV_X1 U22935 ( .A(n10648), .ZN(n10637) );
  NAND2_X1 U22937 ( .A1(n9484), .A2(n10633), .ZN(n10630) );
  NAND3_X1 U22938 ( .A1(n10632), .A2(n51782), .A3(n10630), .ZN(n10636) );
  AND2_X1 U22939 ( .A1(n10634), .A2(n10633), .ZN(n10635) );
  MUX2_X1 U22940 ( .A(n10636), .B(n10635), .S(n9482), .Z(n10644) );
  OAI21_X1 U22941 ( .B1(n14339), .B2(n6073), .A(n13425), .ZN(n10638) );
  AND2_X1 U22943 ( .A1(n13418), .A2(n14342), .ZN(n10640) );
  AOI21_X1 U22944 ( .B1(n10640), .B2(n14346), .A(n14344), .ZN(n10643) );
  NAND2_X1 U22945 ( .A1(n14342), .A2(n6073), .ZN(n13402) );
  NAND2_X1 U22946 ( .A1(n13425), .A2(n13402), .ZN(n10642) );
  NAND2_X1 U22947 ( .A1(n13417), .A2(n14345), .ZN(n12223) );
  INV_X1 U22948 ( .A(n12223), .ZN(n10641) );
  NAND2_X1 U22949 ( .A1(n14339), .A2(n14341), .ZN(n13003) );
  AOI22_X1 U22950 ( .A1(n10643), .A2(n10642), .B1(n10641), .B2(n13003), .ZN(
        n10654) );
  INV_X1 U22951 ( .A(n10644), .ZN(n10645) );
  NAND3_X1 U22952 ( .A1(n10649), .A2(n10648), .A3(n10647), .ZN(n10650) );
  NAND2_X1 U22953 ( .A1(n14353), .A2(n14331), .ZN(n10652) );
  NAND3_X1 U22954 ( .A1(n10652), .A2(n6073), .A3(n13412), .ZN(n10653) );
  XNOR2_X1 U22955 ( .A(n10655), .B(n18791), .ZN(n14112) );
  XNOR2_X1 U22956 ( .A(n10656), .B(n14112), .ZN(n10657) );
  NAND3_X1 U22957 ( .A1(n12045), .A2(n9221), .A3(n10662), .ZN(n10663) );
  OR2_X1 U22958 ( .A1(n10668), .A2(n10667), .ZN(n10682) );
  AOI22_X1 U22959 ( .A1(n10671), .A2(n10670), .B1(n12339), .B2(n12341), .ZN(
        n10681) );
  INV_X1 U22960 ( .A(n10672), .ZN(n12342) );
  NAND3_X1 U22961 ( .A1(n51462), .A2(n12342), .A3(n12325), .ZN(n10675) );
  INV_X1 U22962 ( .A(n10676), .ZN(n10674) );
  NAND4_X1 U22963 ( .A1(n10675), .A2(n10674), .A3(n10673), .A4(n10288), .ZN(
        n10680) );
  OAI21_X1 U22964 ( .B1(n10678), .B2(n10677), .A(n10676), .ZN(n10679) );
  INV_X1 U22965 ( .A(n13317), .ZN(n10692) );
  NOR2_X1 U22966 ( .A1(n12369), .A2(n12389), .ZN(n10684) );
  MUX2_X1 U22967 ( .A(n10685), .B(n10684), .S(n12094), .Z(n10691) );
  AND2_X1 U22968 ( .A1(n10686), .A2(n12380), .ZN(n12098) );
  NAND3_X1 U22970 ( .A1(n12087), .A2(n12380), .A3(n12379), .ZN(n10688) );
  OAI211_X1 U22971 ( .C1(n11353), .C2(n12383), .A(n10689), .B(n10688), .ZN(
        n10690) );
  NAND2_X1 U22972 ( .A1(n10692), .A2(n13316), .ZN(n10732) );
  INV_X1 U22973 ( .A(n10704), .ZN(n10693) );
  OAI22_X1 U22974 ( .A1(n10694), .A2(n12112), .B1(n11373), .B2(n10693), .ZN(
        n10698) );
  NAND2_X1 U22975 ( .A1(n10695), .A2(n11368), .ZN(n10696) );
  NOR2_X1 U22976 ( .A1(n10698), .A2(n10697), .ZN(n10714) );
  INV_X1 U22977 ( .A(n10699), .ZN(n10700) );
  NOR2_X1 U22978 ( .A1(n6677), .A2(n11375), .ZN(n10703) );
  OAI21_X1 U22979 ( .B1(n10703), .B2(n10702), .A(n10701), .ZN(n10708) );
  NAND3_X1 U22980 ( .A1(n12114), .A2(n11379), .A3(n10704), .ZN(n10705) );
  AOI21_X1 U22981 ( .B1(n12107), .B2(n51391), .A(n11377), .ZN(n10711) );
  NAND2_X1 U22982 ( .A1(n12107), .A2(n10709), .ZN(n10710) );
  OAI211_X1 U22983 ( .C1(n12121), .C2(n12113), .A(n10711), .B(n10710), .ZN(
        n10712) );
  NAND2_X1 U22984 ( .A1(n14170), .A2(n14605), .ZN(n10731) );
  NAND2_X1 U22985 ( .A1(n10717), .A2(n10716), .ZN(n10730) );
  AND2_X1 U22986 ( .A1(n12276), .A2(n10718), .ZN(n10721) );
  OAI21_X1 U22987 ( .B1(n10721), .B2(n10720), .A(n10719), .ZN(n10729) );
  AOI22_X1 U22988 ( .A1(n12292), .A2(n10724), .B1(n10723), .B2(n10722), .ZN(
        n10728) );
  NAND3_X1 U22989 ( .A1(n12283), .A2(n10726), .A3(n10725), .ZN(n10727) );
  MUX2_X1 U22990 ( .A(n10732), .B(n10731), .S(n13322), .Z(n10762) );
  INV_X1 U22991 ( .A(n14605), .ZN(n14611) );
  OAI21_X1 U22992 ( .B1(n14611), .B2(n14170), .A(n10733), .ZN(n10755) );
  INV_X1 U22993 ( .A(n12271), .ZN(n11343) );
  OAI21_X1 U22994 ( .B1(n10743), .B2(n10741), .A(n11343), .ZN(n10739) );
  NAND2_X1 U22995 ( .A1(n11346), .A2(n10734), .ZN(n10736) );
  AOI21_X1 U22996 ( .B1(n10737), .B2(n10736), .A(n10735), .ZN(n10738) );
  NAND2_X1 U22997 ( .A1(n10740), .A2(n12254), .ZN(n10752) );
  NOR2_X1 U22998 ( .A1(n10743), .A2(n10742), .ZN(n10744) );
  INV_X1 U22999 ( .A(n10746), .ZN(n10749) );
  NOR2_X1 U23000 ( .A1(n10748), .A2(n10747), .ZN(n11334) );
  OAI21_X1 U23001 ( .B1(n10749), .B2(n11334), .A(n12263), .ZN(n10750) );
  INV_X1 U23003 ( .A(n14612), .ZN(n10754) );
  NAND3_X1 U23004 ( .A1(n10755), .A2(n14006), .A3(n10754), .ZN(n10761) );
  NOR2_X1 U23005 ( .A1(n13316), .A2(n13322), .ZN(n14166) );
  INV_X1 U23006 ( .A(n14166), .ZN(n10758) );
  NOR2_X1 U23007 ( .A1(n51534), .A2(n14605), .ZN(n14169) );
  INV_X1 U23008 ( .A(n14169), .ZN(n10757) );
  OAI21_X1 U23009 ( .B1(n10758), .B2(n14600), .A(n10757), .ZN(n10759) );
  NAND2_X1 U23010 ( .A1(n10759), .A2(n14607), .ZN(n10760) );
  XNOR2_X1 U23011 ( .A(n13316), .B(n14601), .ZN(n10763) );
  NAND2_X1 U23012 ( .A1(n10763), .A2(n14010), .ZN(n10764) );
  NAND2_X1 U23013 ( .A1(n14006), .A2(n13323), .ZN(n14009) );
  INV_X1 U23014 ( .A(n14009), .ZN(n14171) );
  AND2_X1 U23015 ( .A1(n14160), .A2(n14149), .ZN(n12238) );
  NAND3_X1 U23016 ( .A1(n12238), .A2(n14150), .A3(n14159), .ZN(n10768) );
  AND2_X1 U23017 ( .A1(n10768), .A2(n10767), .ZN(n10777) );
  AND2_X1 U23018 ( .A1(n14155), .A2(n13122), .ZN(n10769) );
  OAI21_X1 U23019 ( .B1(n10769), .B2(n12231), .A(n14966), .ZN(n10774) );
  AOI21_X1 U23020 ( .B1(n13122), .B2(n51175), .A(n14966), .ZN(n10770) );
  OAI21_X1 U23021 ( .B1(n10770), .B2(n14156), .A(n14159), .ZN(n10773) );
  OAI21_X1 U23022 ( .B1(n14164), .B2(n14155), .A(n14156), .ZN(n10772) );
  AND2_X1 U23024 ( .A1(n14155), .A2(n14164), .ZN(n13117) );
  INV_X1 U23025 ( .A(n12546), .ZN(n12540) );
  NOR2_X1 U23026 ( .A1(n10778), .A2(n12545), .ZN(n10779) );
  AOI22_X1 U23027 ( .A1(n10786), .A2(n10780), .B1(n12540), .B2(n10779), .ZN(
        n11458) );
  INV_X1 U23028 ( .A(n51674), .ZN(n10785) );
  NAND2_X1 U23029 ( .A1(n10781), .A2(n12537), .ZN(n10783) );
  OAI22_X1 U23030 ( .A1(n10783), .A2(n12533), .B1(n10782), .B2(n9109), .ZN(
        n10784) );
  AOI22_X1 U23031 ( .A1(n12547), .A2(n11445), .B1(n11446), .B2(n12536), .ZN(
        n10789) );
  AND2_X1 U23035 ( .A1(n11489), .A2(n12480), .ZN(n12474) );
  NAND2_X1 U23036 ( .A1(n10791), .A2(n12474), .ZN(n11893) );
  NAND2_X1 U23037 ( .A1(n11070), .A2(n11893), .ZN(n10804) );
  NAND2_X1 U23038 ( .A1(n12491), .A2(n2211), .ZN(n10793) );
  NAND3_X1 U23041 ( .A1(n11485), .A2(n11489), .A3(n2211), .ZN(n10794) );
  INV_X1 U23042 ( .A(n12474), .ZN(n11898) );
  OAI21_X1 U23043 ( .B1(n8099), .B2(n10794), .A(n11898), .ZN(n10798) );
  AND2_X1 U23044 ( .A1(n11066), .A2(n12475), .ZN(n10797) );
  AND2_X1 U23045 ( .A1(n510), .A2(n2211), .ZN(n10795) );
  NOR2_X1 U23046 ( .A1(n11488), .A2(n10795), .ZN(n10796) );
  AOI22_X1 U23047 ( .A1(n11893), .A2(n10798), .B1(n10797), .B2(n10796), .ZN(
        n10802) );
  INV_X1 U23048 ( .A(n12491), .ZN(n10800) );
  NOR2_X1 U23049 ( .A1(n12478), .A2(n510), .ZN(n10799) );
  OAI21_X1 U23050 ( .B1(n10800), .B2(n10799), .A(n11895), .ZN(n10801) );
  NAND4_X1 U23051 ( .A1(n10804), .A2(n10803), .A3(n10802), .A4(n10801), .ZN(
        n10858) );
  OAI21_X1 U23054 ( .B1(n10806), .B2(n11598), .A(n10805), .ZN(n10807) );
  INV_X1 U23055 ( .A(n10807), .ZN(n10824) );
  NAND2_X1 U23056 ( .A1(n3250), .A2(n11608), .ZN(n10808) );
  OAI211_X1 U23057 ( .C1(n11600), .C2(n11611), .A(n10809), .B(n10808), .ZN(
        n10813) );
  INV_X1 U23058 ( .A(n10810), .ZN(n10811) );
  AND2_X1 U23059 ( .A1(n10813), .A2(n10812), .ZN(n10823) );
  OR2_X1 U23060 ( .A1(n10814), .A2(n11244), .ZN(n10822) );
  NAND2_X1 U23061 ( .A1(n11599), .A2(n11601), .ZN(n10820) );
  AOI21_X1 U23062 ( .B1(n10816), .B2(n10815), .A(n9083), .ZN(n10817) );
  NAND3_X1 U23063 ( .A1(n10820), .A2(n10819), .A3(n10818), .ZN(n10821) );
  INV_X1 U23064 ( .A(n10832), .ZN(n10825) );
  OAI21_X1 U23065 ( .B1(n10826), .B2(n12514), .A(n10825), .ZN(n10828) );
  INV_X1 U23066 ( .A(n12506), .ZN(n11261) );
  NAND2_X1 U23067 ( .A1(n8024), .A2(n51653), .ZN(n10835) );
  NOR2_X1 U23068 ( .A1(n11261), .A2(n10835), .ZN(n10827) );
  INV_X1 U23069 ( .A(n11549), .ZN(n12503) );
  NAND3_X1 U23070 ( .A1(n12503), .A2(n11258), .A3(n8024), .ZN(n10829) );
  AND2_X1 U23071 ( .A1(n10830), .A2(n10829), .ZN(n10840) );
  NAND3_X1 U23072 ( .A1(n11550), .A2(n10833), .A3(n8024), .ZN(n10834) );
  INV_X1 U23073 ( .A(n12504), .ZN(n12524) );
  NOR2_X1 U23074 ( .A1(n10835), .A2(n12516), .ZN(n10837) );
  OR2_X1 U23075 ( .A1(n15165), .A2(n14577), .ZN(n13456) );
  XNOR2_X1 U23076 ( .A(n11229), .B(n11460), .ZN(n10842) );
  NAND2_X1 U23077 ( .A1(n10842), .A2(n11634), .ZN(n10844) );
  NAND3_X1 U23078 ( .A1(n11630), .A2(n11468), .A3(n11634), .ZN(n10843) );
  NAND2_X1 U23079 ( .A1(n11634), .A2(n11624), .ZN(n10846) );
  NOR2_X1 U23080 ( .A1(n11625), .A2(n10846), .ZN(n10848) );
  NAND3_X1 U23081 ( .A1(n4150), .A2(n11470), .A3(n11467), .ZN(n10847) );
  NOR2_X1 U23082 ( .A1(n11635), .A2(n11634), .ZN(n10850) );
  NOR2_X1 U23083 ( .A1(n10852), .A2(n11633), .ZN(n10849) );
  AOI22_X1 U23084 ( .A1(n10851), .A2(n10850), .B1(n10849), .B2(n11629), .ZN(
        n10856) );
  AOI21_X1 U23085 ( .B1(n11629), .B2(n11635), .A(n11468), .ZN(n10854) );
  NOR2_X1 U23086 ( .A1(n10852), .A2(n11460), .ZN(n10853) );
  OAI21_X1 U23087 ( .B1(n10854), .B2(n10853), .A(n11631), .ZN(n10855) );
  INV_X1 U23088 ( .A(n10858), .ZN(n14579) );
  OAI21_X1 U23089 ( .B1(n10860), .B2(n51760), .A(n12572), .ZN(n10861) );
  INV_X1 U23090 ( .A(n11570), .ZN(n12578) );
  NAND2_X1 U23091 ( .A1(n12574), .A2(n11581), .ZN(n11512) );
  OAI21_X1 U23092 ( .B1(n12556), .B2(n11189), .A(n11530), .ZN(n10862) );
  XNOR2_X1 U23093 ( .A(n12573), .B(n11514), .ZN(n12558) );
  INV_X1 U23094 ( .A(n12558), .ZN(n11565) );
  NAND2_X1 U23095 ( .A1(n15163), .A2(n15177), .ZN(n15164) );
  OAI211_X1 U23096 ( .C1(n15174), .C2(n15167), .A(n15171), .B(n15164), .ZN(
        n10868) );
  NAND2_X1 U23097 ( .A1(n15161), .A2(n15177), .ZN(n10865) );
  NAND2_X1 U23098 ( .A1(n10866), .A2(n15178), .ZN(n10867) );
  INV_X1 U23099 ( .A(n10877), .ZN(n14574) );
  NAND2_X1 U23100 ( .A1(n15161), .A2(n15173), .ZN(n15158) );
  INV_X1 U23101 ( .A(n15158), .ZN(n10869) );
  AOI21_X1 U23102 ( .B1(n10870), .B2(n10869), .A(n14128), .ZN(n10871) );
  INV_X1 U23103 ( .A(n10871), .ZN(n10872) );
  NAND2_X1 U23104 ( .A1(n15161), .A2(n15167), .ZN(n10875) );
  OR2_X1 U23105 ( .A1(n15177), .A2(n51370), .ZN(n13464) );
  INV_X1 U23106 ( .A(n13464), .ZN(n10873) );
  NOR2_X1 U23107 ( .A1(n15163), .A2(n15177), .ZN(n14575) );
  AND2_X1 U23108 ( .A1(n51370), .A2(n15167), .ZN(n13457) );
  OAI21_X1 U23110 ( .B1(n13512), .B2(n10882), .A(n13524), .ZN(n12934) );
  NAND2_X1 U23111 ( .A1(n11840), .A2(n13525), .ZN(n10883) );
  NAND2_X1 U23112 ( .A1(n12934), .A2(n10883), .ZN(n10896) );
  NOR2_X1 U23113 ( .A1(n11843), .A2(n13502), .ZN(n13498) );
  NOR2_X1 U23114 ( .A1(n13512), .A2(n13526), .ZN(n10886) );
  NAND2_X1 U23115 ( .A1(n10884), .A2(n13514), .ZN(n10885) );
  OAI211_X1 U23116 ( .C1(n13498), .C2(n13514), .A(n10886), .B(n10885), .ZN(
        n10895) );
  OR2_X1 U23117 ( .A1(n13525), .A2(n13526), .ZN(n10888) );
  NAND2_X1 U23118 ( .A1(n51683), .A2(n13526), .ZN(n10887) );
  OAI22_X1 U23119 ( .A1(n11840), .A2(n10888), .B1(n11841), .B2(n10887), .ZN(
        n10891) );
  NOR2_X1 U23120 ( .A1(n10889), .A2(n11845), .ZN(n10890) );
  NOR2_X1 U23121 ( .A1(n10891), .A2(n10890), .ZN(n10894) );
  NOR2_X1 U23122 ( .A1(n13506), .A2(n13525), .ZN(n10892) );
  OAI211_X1 U23123 ( .C1(n13499), .C2(n10892), .A(n13500), .B(n51066), .ZN(
        n10893) );
  NAND4_X2 U23124 ( .A1(n10896), .A2(n10895), .A3(n10894), .A4(n10893), .ZN(
        n17690) );
  AND2_X1 U23125 ( .A1(n13780), .A2(n13173), .ZN(n10907) );
  NAND2_X1 U23126 ( .A1(n10905), .A2(n12419), .ZN(n10897) );
  NAND4_X1 U23127 ( .A1(n10907), .A2(n10899), .A3(n10898), .A4(n10897), .ZN(
        n10900) );
  MUX2_X1 U23128 ( .A(n10900), .B(n10906), .S(n13169), .Z(n10912) );
  AND2_X1 U23129 ( .A1(n13782), .A2(n13780), .ZN(n10902) );
  AOI22_X1 U23130 ( .A1(n10905), .A2(n12423), .B1(n10902), .B2(n10901), .ZN(
        n10911) );
  NOR2_X1 U23131 ( .A1(n13787), .A2(n12419), .ZN(n10903) );
  OAI21_X1 U23132 ( .B1(n10904), .B2(n10903), .A(n13178), .ZN(n10910) );
  NAND2_X1 U23133 ( .A1(n13780), .A2(n788), .ZN(n13166) );
  OAI21_X1 U23135 ( .B1(n13161), .B2(n10906), .A(n13778), .ZN(n10908) );
  OAI21_X1 U23136 ( .B1(n10908), .B2(n13772), .A(n13170), .ZN(n10909) );
  NAND4_X1 U23137 ( .A1(n52189), .A2(n10920), .A3(n9807), .A4(n10925), .ZN(
        n10916) );
  NAND4_X1 U23138 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(
        n10937) );
  NAND2_X1 U23139 ( .A1(n10931), .A2(n9807), .ZN(n10934) );
  OAI21_X1 U23140 ( .B1(n10939), .B2(n10938), .A(n12300), .ZN(n10941) );
  NAND2_X1 U23141 ( .A1(n10941), .A2(n10940), .ZN(n10944) );
  NAND3_X1 U23142 ( .A1(n10942), .A2(n12317), .A3(n12312), .ZN(n10943) );
  OAI21_X1 U23143 ( .B1(n10945), .B2(n12303), .A(n804), .ZN(n10946) );
  OAI21_X1 U23144 ( .B1(n10948), .B2(n10947), .A(n10946), .ZN(n10949) );
  NAND2_X1 U23145 ( .A1(n10952), .A2(n12302), .ZN(n10953) );
  NAND2_X1 U23146 ( .A1(n10958), .A2(n10957), .ZN(n10975) );
  AOI22_X1 U23147 ( .A1(n10962), .A2(n10961), .B1(n10960), .B2(n10959), .ZN(
        n10974) );
  NAND3_X1 U23148 ( .A1(n10965), .A2(n10964), .A3(n10963), .ZN(n10973) );
  OAI21_X1 U23149 ( .B1(n10968), .B2(n10967), .A(n10966), .ZN(n10969) );
  NAND3_X1 U23150 ( .A1(n10971), .A2(n10970), .A3(n10969), .ZN(n10972) );
  INV_X1 U23151 ( .A(n10988), .ZN(n10977) );
  NAND2_X1 U23152 ( .A1(n10992), .A2(n12357), .ZN(n12362) );
  OAI211_X1 U23153 ( .C1(n10987), .C2(n10977), .A(n12362), .B(n10976), .ZN(
        n10980) );
  OAI22_X1 U23156 ( .A1(n10990), .A2(n12350), .B1(n51137), .B2(n12356), .ZN(
        n10994) );
  NOR2_X1 U23157 ( .A1(n10991), .A2(n8791), .ZN(n10993) );
  INV_X1 U23159 ( .A(n10998), .ZN(n10999) );
  OAI21_X1 U23160 ( .B1(n11001), .B2(n11000), .A(n10999), .ZN(n11020) );
  OAI21_X1 U23161 ( .B1(n11003), .B2(n11002), .A(n11011), .ZN(n11019) );
  NAND3_X1 U23162 ( .A1(n11005), .A2(n11004), .A3(n11008), .ZN(n11010) );
  INV_X1 U23163 ( .A(n11006), .ZN(n11007) );
  NAND3_X1 U23164 ( .A1(n11008), .A2(n11015), .A3(n11007), .ZN(n11009) );
  AND2_X1 U23165 ( .A1(n11010), .A2(n11009), .ZN(n11018) );
  NAND2_X1 U23166 ( .A1(n11012), .A2(n11011), .ZN(n11013) );
  OAI211_X1 U23167 ( .C1(n11016), .C2(n11015), .A(n11014), .B(n11013), .ZN(
        n11017) );
  NAND4_X2 U23168 ( .A1(n11020), .A2(n11018), .A3(n11019), .A4(n11017), .ZN(
        n14022) );
  OAI22_X1 U23169 ( .A1(n13296), .A2(n469), .B1(n14036), .B2(n14033), .ZN(
        n11042) );
  INV_X1 U23170 ( .A(n13291), .ZN(n13306) );
  INV_X1 U23171 ( .A(n11021), .ZN(n11026) );
  OAI211_X1 U23172 ( .C1(n11026), .C2(n11025), .A(n11024), .B(n11036), .ZN(
        n11039) );
  NAND2_X1 U23173 ( .A1(n580), .A2(n11027), .ZN(n11029) );
  OAI22_X1 U23174 ( .A1(n11032), .A2(n11031), .B1(n11030), .B2(n11029), .ZN(
        n11034) );
  AND2_X1 U23175 ( .A1(n13729), .A2(n12410), .ZN(n11041) );
  NAND2_X1 U23176 ( .A1(n11042), .A2(n11041), .ZN(n11054) );
  INV_X1 U23177 ( .A(n13736), .ZN(n14024) );
  NAND3_X1 U23178 ( .A1(n14024), .A2(n469), .A3(n14022), .ZN(n11046) );
  NAND2_X1 U23179 ( .A1(n14032), .A2(n14022), .ZN(n14028) );
  INV_X1 U23180 ( .A(n14028), .ZN(n11043) );
  OAI21_X1 U23181 ( .B1(n11043), .B2(n13291), .A(n14030), .ZN(n11045) );
  MUX2_X1 U23183 ( .A(n11046), .B(n11045), .S(n47), .Z(n11053) );
  INV_X1 U23184 ( .A(n14029), .ZN(n13303) );
  OR2_X1 U23185 ( .A1(n14033), .A2(n13303), .ZN(n14018) );
  NOR2_X1 U23186 ( .A1(n14032), .A2(n14030), .ZN(n14019) );
  INV_X1 U23187 ( .A(n14022), .ZN(n13297) );
  NAND2_X1 U23188 ( .A1(n11049), .A2(n11048), .ZN(n11051) );
  AND2_X1 U23189 ( .A1(n13291), .A2(n469), .ZN(n14023) );
  NOR2_X1 U23190 ( .A1(n13291), .A2(n469), .ZN(n11050) );
  AND2_X1 U23191 ( .A1(n14030), .A2(n11050), .ZN(n14035) );
  AOI21_X1 U23192 ( .B1(n11051), .B2(n14023), .A(n14035), .ZN(n11052) );
  XNOR2_X1 U23193 ( .A(n16653), .B(n16485), .ZN(n11183) );
  NOR2_X1 U23194 ( .A1(n13061), .A2(n14139), .ZN(n13064) );
  NOR2_X1 U23195 ( .A1(n15259), .A2(n13064), .ZN(n11058) );
  NAND2_X1 U23196 ( .A1(n13061), .A2(n14139), .ZN(n15255) );
  OAI211_X1 U23197 ( .C1(n11058), .C2(n14137), .A(n15255), .B(n15266), .ZN(
        n11057) );
  NAND2_X1 U23198 ( .A1(n14784), .A2(n13069), .ZN(n13060) );
  INV_X1 U23199 ( .A(n13060), .ZN(n11056) );
  INV_X1 U23200 ( .A(n14791), .ZN(n15265) );
  OR2_X1 U23201 ( .A1(n13061), .A2(n13069), .ZN(n14796) );
  NAND3_X1 U23202 ( .A1(n11058), .A2(n15265), .A3(n14796), .ZN(n11061) );
  INV_X1 U23203 ( .A(n14784), .ZN(n15250) );
  NAND4_X1 U23204 ( .A1(n51685), .A2(n15250), .A3(n14139), .A4(n13061), .ZN(
        n14787) );
  INV_X1 U23205 ( .A(n15254), .ZN(n13071) );
  NAND2_X1 U23206 ( .A1(n13071), .A2(n15257), .ZN(n14143) );
  INV_X1 U23207 ( .A(n14143), .ZN(n11059) );
  NAND2_X1 U23208 ( .A1(n11059), .A2(n15259), .ZN(n11060) );
  NAND3_X1 U23210 ( .A1(n12491), .A2(n11063), .A3(n11062), .ZN(n11064) );
  NOR2_X1 U23211 ( .A1(n11067), .A2(n12478), .ZN(n11068) );
  NOR2_X1 U23212 ( .A1(n11069), .A2(n11068), .ZN(n11076) );
  INV_X1 U23213 ( .A(n11070), .ZN(n11075) );
  OAI22_X1 U23214 ( .A1(n11488), .A2(n12486), .B1(n11898), .B2(n510), .ZN(
        n11073) );
  NOR2_X1 U23215 ( .A1(n11071), .A2(n12471), .ZN(n11072) );
  OAI211_X1 U23216 ( .C1(n11073), .C2(n11072), .A(n2211), .B(n12481), .ZN(
        n11074) );
  AND2_X1 U23217 ( .A1(n11884), .A2(n12679), .ZN(n11088) );
  OAI21_X1 U23218 ( .B1(n592), .B2(n12676), .A(n12672), .ZN(n11087) );
  OAI21_X1 U23219 ( .B1(n12672), .B2(n592), .A(n11874), .ZN(n11078) );
  NAND2_X1 U23220 ( .A1(n11078), .A2(n50997), .ZN(n11081) );
  NAND2_X1 U23221 ( .A1(n12667), .A2(n11884), .ZN(n12459) );
  INV_X1 U23222 ( .A(n12459), .ZN(n11080) );
  NAND4_X1 U23223 ( .A1(n11081), .A2(n11080), .A3(n11501), .A4(n11079), .ZN(
        n11086) );
  OAI211_X1 U23224 ( .C1(n11879), .C2(n592), .A(n11084), .B(n12676), .ZN(
        n11085) );
  NOR2_X1 U23225 ( .A1(n51673), .A2(n11089), .ZN(n11455) );
  OAI21_X1 U23226 ( .B1(n11455), .B2(n12538), .A(n11443), .ZN(n11090) );
  NAND2_X1 U23227 ( .A1(n11090), .A2(n11447), .ZN(n11104) );
  NAND4_X1 U23228 ( .A1(n51673), .A2(n442), .A3(n12537), .A4(n6409), .ZN(
        n11094) );
  NAND3_X1 U23229 ( .A1(n11092), .A2(n12537), .A3(n11091), .ZN(n11093) );
  AND3_X1 U23230 ( .A1(n11095), .A2(n11094), .A3(n11093), .ZN(n11103) );
  INV_X1 U23231 ( .A(n11096), .ZN(n11098) );
  INV_X1 U23232 ( .A(n12543), .ZN(n11097) );
  AOI22_X1 U23233 ( .A1(n11098), .A2(n51674), .B1(n12549), .B2(n11097), .ZN(
        n11102) );
  INV_X1 U23234 ( .A(n11446), .ZN(n11099) );
  OAI21_X1 U23235 ( .B1(n12535), .B2(n12540), .A(n11100), .ZN(n11101) );
  INV_X1 U23237 ( .A(n15189), .ZN(n15234) );
  INV_X1 U23238 ( .A(n15235), .ZN(n11150) );
  OR2_X1 U23240 ( .A1(n11108), .A2(n11107), .ZN(n12732) );
  NAND2_X1 U23241 ( .A1(n11109), .A2(n11964), .ZN(n11110) );
  NAND4_X1 U23242 ( .A1(n11111), .A2(n12732), .A3(n11948), .A4(n11110), .ZN(
        n11116) );
  OAI21_X1 U23243 ( .B1(n8882), .B2(n11964), .A(n11113), .ZN(n11115) );
  NAND3_X1 U23244 ( .A1(n11960), .A2(n11942), .A3(n11958), .ZN(n11114) );
  NAND2_X1 U23245 ( .A1(n15244), .A2(n14767), .ZN(n11118) );
  NAND3_X1 U23246 ( .A1(n11150), .A2(n15234), .A3(n11118), .ZN(n11119) );
  OAI21_X1 U23247 ( .B1(n14769), .B2(n15234), .A(n11119), .ZN(n11146) );
  INV_X1 U23248 ( .A(n12696), .ZN(n12442) );
  INV_X1 U23249 ( .A(n11930), .ZN(n11120) );
  OAI211_X1 U23250 ( .C1(n12699), .C2(n12690), .A(n12442), .B(n11120), .ZN(
        n11121) );
  OAI22_X1 U23251 ( .A1(n12701), .A2(n12705), .B1(n11123), .B2(n12440), .ZN(
        n11124) );
  AND2_X1 U23252 ( .A1(n12700), .A2(n12709), .ZN(n12444) );
  NAND2_X1 U23253 ( .A1(n11124), .A2(n12444), .ZN(n11127) );
  INV_X1 U23254 ( .A(n12436), .ZN(n11126) );
  NAND2_X1 U23255 ( .A1(n11125), .A2(n12441), .ZN(n12698) );
  NAND2_X1 U23256 ( .A1(n11128), .A2(n11920), .ZN(n11143) );
  NAND3_X1 U23257 ( .A1(n12597), .A2(n795), .A3(n9539), .ZN(n11135) );
  NAND3_X1 U23258 ( .A1(n11132), .A2(n1307), .A3(n52140), .ZN(n11134) );
  NAND3_X1 U23259 ( .A1(n3692), .A2(n1307), .A3(n357), .ZN(n11133) );
  AND3_X1 U23260 ( .A1(n11135), .A2(n11134), .A3(n11133), .ZN(n11141) );
  INV_X1 U23263 ( .A(n11144), .ZN(n15243) );
  OR2_X1 U23264 ( .A1(n13277), .A2(n15243), .ZN(n15237) );
  INV_X1 U23265 ( .A(n15237), .ZN(n15203) );
  NAND2_X1 U23266 ( .A1(n14769), .A2(n15196), .ZN(n11145) );
  NAND3_X1 U23267 ( .A1(n11146), .A2(n15203), .A3(n11145), .ZN(n11156) );
  INV_X1 U23268 ( .A(n15236), .ZN(n14120) );
  NOR2_X1 U23269 ( .A1(n14120), .A2(n14763), .ZN(n11147) );
  AND2_X1 U23270 ( .A1(n15189), .A2(n15204), .ZN(n15197) );
  AOI22_X1 U23271 ( .A1(n11147), .A2(n15205), .B1(n14769), .B2(n15197), .ZN(
        n11155) );
  INV_X1 U23272 ( .A(n14767), .ZN(n14759) );
  NAND2_X1 U23273 ( .A1(n14759), .A2(n15204), .ZN(n13271) );
  INV_X1 U23274 ( .A(n13271), .ZN(n11148) );
  AND2_X1 U23275 ( .A1(n15189), .A2(n15233), .ZN(n14762) );
  OAI21_X1 U23276 ( .B1(n15245), .B2(n11148), .A(n14762), .ZN(n11154) );
  NAND2_X1 U23277 ( .A1(n15188), .A2(n15243), .ZN(n11151) );
  AND2_X1 U23278 ( .A1(n14767), .A2(n15204), .ZN(n15194) );
  NAND4_X1 U23279 ( .A1(n13277), .A2(n15243), .A3(n15194), .A4(n15189), .ZN(
        n11149) );
  OAI21_X1 U23280 ( .B1(n11151), .B2(n11150), .A(n11149), .ZN(n11152) );
  INV_X1 U23281 ( .A(n11152), .ZN(n11153) );
  NAND2_X1 U23282 ( .A1(n13102), .A2(n12914), .ZN(n13075) );
  NOR2_X1 U23283 ( .A1(n13091), .A2(n11160), .ZN(n12913) );
  INV_X1 U23284 ( .A(n12913), .ZN(n11158) );
  NOR2_X1 U23285 ( .A1(n12915), .A2(n13092), .ZN(n13077) );
  NAND2_X1 U23286 ( .A1(n11158), .A2(n13077), .ZN(n11159) );
  INV_X1 U23287 ( .A(n12820), .ZN(n11166) );
  NAND3_X1 U23288 ( .A1(n13091), .A2(n11160), .A3(n13102), .ZN(n11164) );
  INV_X1 U23289 ( .A(n11161), .ZN(n11162) );
  NAND3_X1 U23290 ( .A1(n11162), .A2(n13086), .A3(n13092), .ZN(n11163) );
  NOR2_X1 U23291 ( .A1(n11166), .A2(n11165), .ZN(n11171) );
  INV_X1 U23292 ( .A(n13100), .ZN(n11167) );
  OAI211_X1 U23293 ( .C1(n11167), .C2(n13092), .A(n13091), .B(n13089), .ZN(
        n11170) );
  INV_X1 U23294 ( .A(n11168), .ZN(n11169) );
  INV_X1 U23295 ( .A(n12907), .ZN(n13137) );
  MUX2_X1 U23296 ( .A(n14181), .B(n11172), .S(n13137), .Z(n11182) );
  NAND3_X1 U23297 ( .A1(n12900), .A2(n14178), .A3(n13148), .ZN(n13144) );
  INV_X1 U23298 ( .A(n13144), .ZN(n11174) );
  NAND2_X1 U23299 ( .A1(n13148), .A2(n14186), .ZN(n14190) );
  NOR2_X1 U23300 ( .A1(n3679), .A2(n14178), .ZN(n12905) );
  NOR2_X1 U23301 ( .A1(n12907), .A2(n13152), .ZN(n12216) );
  INV_X1 U23302 ( .A(n12216), .ZN(n11173) );
  OAI22_X1 U23303 ( .A1(n11174), .A2(n12899), .B1(n12905), .B2(n11173), .ZN(
        n11181) );
  NAND2_X1 U23304 ( .A1(n12907), .A2(n14186), .ZN(n14177) );
  NAND4_X1 U23305 ( .A1(n12907), .A2(n13135), .A3(n13152), .A4(n14186), .ZN(
        n11175) );
  OAI211_X1 U23306 ( .C1(n13153), .C2(n14177), .A(n11176), .B(n11175), .ZN(
        n11177) );
  AND2_X1 U23307 ( .A1(n11178), .A2(n13148), .ZN(n12906) );
  OAI21_X1 U23308 ( .B1(n6609), .B2(n13137), .A(n14187), .ZN(n11179) );
  NAND2_X1 U23309 ( .A1(n12906), .A2(n11179), .ZN(n11180) );
  XNOR2_X1 U23310 ( .A(n18704), .B(n560), .ZN(n18604) );
  AND2_X1 U23311 ( .A1(n11581), .A2(n11514), .ZN(n12553) );
  NAND2_X1 U23312 ( .A1(n12553), .A2(n11530), .ZN(n11185) );
  INV_X1 U23315 ( .A(n11508), .ZN(n11187) );
  NOR2_X1 U23316 ( .A1(n11187), .A2(n11186), .ZN(n12566) );
  OAI21_X1 U23317 ( .B1(n11569), .B2(n11189), .A(n11188), .ZN(n11190) );
  NOR2_X1 U23318 ( .A1(n12566), .A2(n11190), .ZN(n11196) );
  INV_X1 U23319 ( .A(n11191), .ZN(n11192) );
  NAND3_X1 U23320 ( .A1(n11192), .A2(n12556), .A3(n51491), .ZN(n11195) );
  NOR2_X1 U23321 ( .A1(n12572), .A2(n51760), .ZN(n11520) );
  NAND2_X1 U23322 ( .A1(n11193), .A2(n11520), .ZN(n11194) );
  NAND3_X1 U23323 ( .A1(n11715), .A2(n11714), .A3(n11696), .ZN(n11207) );
  INV_X1 U23324 ( .A(n11709), .ZN(n11202) );
  INV_X1 U23325 ( .A(n11198), .ZN(n11706) );
  NAND2_X1 U23326 ( .A1(n11706), .A2(n11199), .ZN(n11201) );
  OAI211_X1 U23327 ( .C1(n11212), .C2(n11202), .A(n11201), .B(n11200), .ZN(
        n11206) );
  NAND3_X1 U23328 ( .A1(n11204), .A2(n9146), .A3(n11203), .ZN(n11205) );
  AND3_X1 U23329 ( .A1(n11206), .A2(n11207), .A3(n11205), .ZN(n11223) );
  INV_X1 U23330 ( .A(n11711), .ZN(n11216) );
  NAND2_X1 U23331 ( .A1(n11208), .A2(n11216), .ZN(n11222) );
  OAI22_X1 U23332 ( .A1(n11212), .A2(n11211), .B1(n11210), .B2(n11209), .ZN(
        n11213) );
  OAI21_X1 U23333 ( .B1(n11214), .B2(n11213), .A(n11709), .ZN(n11221) );
  XNOR2_X1 U23334 ( .A(n9933), .B(n11705), .ZN(n11219) );
  AOI21_X1 U23335 ( .B1(n51970), .B2(n11215), .A(n11695), .ZN(n11218) );
  OAI21_X1 U23336 ( .B1(n11216), .B2(n11696), .A(n9933), .ZN(n11217) );
  NAND3_X1 U23337 ( .A1(n11219), .A2(n11218), .A3(n11217), .ZN(n11220) );
  NAND2_X1 U23339 ( .A1(n11635), .A2(n453), .ZN(n11225) );
  AND2_X1 U23340 ( .A1(n11634), .A2(n11467), .ZN(n11476) );
  OAI211_X1 U23341 ( .C1(n11635), .C2(n11226), .A(n11225), .B(n11476), .ZN(
        n11227) );
  INV_X1 U23342 ( .A(n11627), .ZN(n11240) );
  AND2_X1 U23343 ( .A1(n453), .A2(n11467), .ZN(n11469) );
  INV_X1 U23344 ( .A(n11469), .ZN(n11228) );
  NOR2_X1 U23345 ( .A1(n11228), .A2(n11468), .ZN(n11232) );
  NAND2_X1 U23346 ( .A1(n11624), .A2(n11229), .ZN(n11230) );
  NAND2_X1 U23347 ( .A1(n11230), .A2(n11619), .ZN(n11231) );
  AOI22_X1 U23348 ( .A1(n11232), .A2(n3024), .B1(n11464), .B2(n11231), .ZN(
        n11236) );
  INV_X1 U23349 ( .A(n11460), .ZN(n11233) );
  NAND3_X1 U23350 ( .A1(n11631), .A2(n11234), .A3(n11233), .ZN(n11235) );
  AND2_X1 U23352 ( .A1(n11244), .A2(n11242), .ZN(n11246) );
  NAND2_X1 U23353 ( .A1(n9083), .A2(n3250), .ZN(n11243) );
  OAI21_X1 U23354 ( .B1(n11244), .B2(n11243), .A(n11610), .ZN(n11245) );
  OAI21_X1 U23355 ( .B1(n11247), .B2(n11246), .A(n11245), .ZN(n11254) );
  NOR2_X1 U23356 ( .A1(n11598), .A2(n9083), .ZN(n11248) );
  AOI22_X1 U23357 ( .A1(n11248), .A2(n11600), .B1(n11601), .B2(n11608), .ZN(
        n11253) );
  OAI22_X1 U23358 ( .A1(n11250), .A2(n11612), .B1(n11249), .B2(n11613), .ZN(
        n11251) );
  NAND2_X1 U23359 ( .A1(n11251), .A2(n11611), .ZN(n11252) );
  INV_X1 U23360 ( .A(n12961), .ZN(n14072) );
  NAND2_X1 U23361 ( .A1(n12963), .A2(n3512), .ZN(n14407) );
  NAND2_X1 U23362 ( .A1(n11257), .A2(n11256), .ZN(n11267) );
  NAND3_X1 U23363 ( .A1(n11258), .A2(n12512), .A3(n51653), .ZN(n11259) );
  AND2_X1 U23366 ( .A1(n642), .A2(n12518), .ZN(n12507) );
  NAND3_X1 U23367 ( .A1(n11262), .A2(n12507), .A3(n12504), .ZN(n11265) );
  NAND2_X1 U23368 ( .A1(n12515), .A2(n12514), .ZN(n12511) );
  INV_X1 U23369 ( .A(n14410), .ZN(n12965) );
  NOR2_X1 U23370 ( .A1(n14407), .A2(n12965), .ZN(n14074) );
  INV_X1 U23371 ( .A(n14074), .ZN(n11287) );
  NAND2_X1 U23372 ( .A1(n11269), .A2(n11268), .ZN(n11680) );
  INV_X1 U23373 ( .A(n11680), .ZN(n11271) );
  AOI22_X1 U23374 ( .A1(n11271), .A2(n11669), .B1(n11686), .B2(n11270), .ZN(
        n11286) );
  AND2_X1 U23375 ( .A1(n11272), .A2(n11276), .ZN(n11273) );
  NOR2_X1 U23376 ( .A1(n11274), .A2(n11273), .ZN(n11277) );
  NAND2_X1 U23377 ( .A1(n9337), .A2(n9341), .ZN(n11684) );
  INV_X1 U23378 ( .A(n11684), .ZN(n11282) );
  NAND2_X1 U23379 ( .A1(n11276), .A2(n11275), .ZN(n11674) );
  OAI21_X1 U23380 ( .B1(n11685), .B2(n11280), .A(n11279), .ZN(n11281) );
  NAND2_X1 U23381 ( .A1(n11281), .A2(n11673), .ZN(n11284) );
  OAI21_X1 U23382 ( .B1(n11672), .B2(n11282), .A(n11671), .ZN(n11283) );
  MUX2_X1 U23383 ( .A(n14065), .B(n11287), .S(n14393), .Z(n11302) );
  AND2_X1 U23384 ( .A1(n12961), .A2(n14410), .ZN(n11998) );
  INV_X1 U23385 ( .A(n11998), .ZN(n11288) );
  NAND2_X1 U23386 ( .A1(n14412), .A2(n12963), .ZN(n11297) );
  AND2_X1 U23387 ( .A1(n12961), .A2(n14070), .ZN(n11289) );
  INV_X1 U23388 ( .A(n14412), .ZN(n12871) );
  NAND3_X1 U23389 ( .A1(n11289), .A2(n12871), .A3(n14393), .ZN(n12863) );
  OAI21_X1 U23390 ( .B1(n11288), .B2(n11297), .A(n12863), .ZN(n11292) );
  AND2_X1 U23391 ( .A1(n14070), .A2(n14072), .ZN(n11290) );
  NAND4_X1 U23392 ( .A1(n12871), .A2(n11290), .A3(n12963), .A4(n14410), .ZN(
        n11291) );
  INV_X1 U23393 ( .A(n11293), .ZN(n14411) );
  OR2_X1 U23394 ( .A1(n14394), .A2(n14408), .ZN(n12867) );
  OAI21_X1 U23395 ( .B1(n12867), .B2(n14410), .A(n14072), .ZN(n11295) );
  NAND2_X1 U23397 ( .A1(n11295), .A2(n11294), .ZN(n11300) );
  INV_X1 U23398 ( .A(n12869), .ZN(n11999) );
  INV_X1 U23399 ( .A(n11297), .ZN(n11298) );
  NAND2_X1 U23400 ( .A1(n14071), .A2(n11298), .ZN(n11299) );
  XNOR2_X1 U23401 ( .A(n15883), .B(n4855), .ZN(n16758) );
  NAND2_X1 U23402 ( .A1(n12756), .A2(n13669), .ZN(n14640) );
  NAND3_X1 U23403 ( .A1(n12757), .A2(n14641), .A3(n12756), .ZN(n11305) );
  NAND2_X1 U23404 ( .A1(n11306), .A2(n11305), .ZN(n11307) );
  NOR2_X1 U23405 ( .A1(n14639), .A2(n11307), .ZN(n11309) );
  AOI22_X1 U23407 ( .A1(n12754), .A2(n14631), .B1(n13653), .B2(n13667), .ZN(
        n11308) );
  INV_X1 U23408 ( .A(n14673), .ZN(n11310) );
  NAND2_X1 U23409 ( .A1(n13632), .A2(n785), .ZN(n14663) );
  OR2_X1 U23411 ( .A1(n14666), .A2(n7755), .ZN(n12949) );
  NAND4_X1 U23414 ( .A1(n13632), .A2(n14665), .A3(n11315), .A4(n783), .ZN(
        n13640) );
  INV_X1 U23415 ( .A(n13640), .ZN(n11316) );
  OAI21_X1 U23416 ( .B1(n14671), .B2(n11316), .A(n785), .ZN(n11320) );
  OAI21_X1 U23417 ( .B1(n2150), .B2(n14664), .A(n13620), .ZN(n11318) );
  NAND2_X1 U23418 ( .A1(n14666), .A2(n785), .ZN(n12831) );
  INV_X1 U23419 ( .A(n12831), .ZN(n11317) );
  NAND2_X1 U23420 ( .A1(n11318), .A2(n11317), .ZN(n11319) );
  XNOR2_X1 U23421 ( .A(n15454), .B(n16758), .ZN(n15609) );
  OAI211_X1 U23422 ( .C1(n11330), .C2(n11322), .A(n12161), .B(n12169), .ZN(
        n11327) );
  NAND3_X1 U23423 ( .A1(n11323), .A2(n12169), .A3(n12175), .ZN(n11326) );
  OAI211_X1 U23424 ( .C1(n12178), .C2(n11328), .A(n12160), .B(n12175), .ZN(
        n11332) );
  NAND4_X1 U23425 ( .A1(n12171), .A2(n11330), .A3(n11329), .A4(n12169), .ZN(
        n11331) );
  INV_X1 U23426 ( .A(n11334), .ZN(n11336) );
  OAI21_X1 U23427 ( .B1(n11344), .B2(n11339), .A(n11338), .ZN(n11340) );
  NAND3_X1 U23428 ( .A1(n12260), .A2(n11341), .A3(n12254), .ZN(n11342) );
  NOR2_X1 U23429 ( .A1(n11346), .A2(n11345), .ZN(n11347) );
  OAI21_X1 U23430 ( .B1(n11348), .B2(n11347), .A(n12269), .ZN(n11349) );
  OAI21_X1 U23431 ( .B1(n12379), .B2(n12383), .A(n12380), .ZN(n11350) );
  OAI211_X1 U23432 ( .C1(n11351), .C2(n12380), .A(n12097), .B(n11350), .ZN(
        n11356) );
  OAI22_X1 U23433 ( .A1(n51138), .A2(n12094), .B1(n12093), .B2(n11354), .ZN(
        n11355) );
  XNOR2_X1 U23434 ( .A(Key[153]), .B(Key[78]), .ZN(n11358) );
  XNOR2_X1 U23435 ( .A(Ciphertext[191]), .B(Ciphertext[188]), .ZN(n11357) );
  XNOR2_X1 U23436 ( .A(n11358), .B(n11357), .ZN(n11360) );
  NAND2_X1 U23437 ( .A1(n11360), .A2(n11359), .ZN(n11362) );
  OAI21_X1 U23438 ( .B1(n51391), .B2(n11368), .A(n11362), .ZN(n11364) );
  NAND2_X1 U23439 ( .A1(n11362), .A2(n12106), .ZN(n11363) );
  NAND3_X1 U23440 ( .A1(n11364), .A2(n12108), .A3(n11363), .ZN(n11386) );
  NAND2_X1 U23441 ( .A1(n11366), .A2(n12112), .ZN(n11385) );
  AND2_X1 U23442 ( .A1(n11367), .A2(n12112), .ZN(n11369) );
  NAND4_X1 U23443 ( .A1(n11370), .A2(n11369), .A3(n11368), .A4(n11377), .ZN(
        n11371) );
  AND2_X1 U23444 ( .A1(n11371), .A2(n11372), .ZN(n11384) );
  INV_X1 U23445 ( .A(n11373), .ZN(n11382) );
  OAI21_X1 U23446 ( .B1(n4167), .B2(n11375), .A(n11374), .ZN(n11381) );
  NAND4_X1 U23447 ( .A1(n12107), .A2(n11377), .A3(n12112), .A4(n12117), .ZN(
        n11378) );
  OAI21_X1 U23449 ( .B1(n11382), .B2(n11381), .A(n11380), .ZN(n11383) );
  NAND2_X1 U23450 ( .A1(n11388), .A2(n11387), .ZN(n11392) );
  NAND2_X1 U23451 ( .A1(n11389), .A2(n12055), .ZN(n11391) );
  MUX2_X1 U23452 ( .A(n11392), .B(n11391), .S(n11390), .Z(n11397) );
  AND3_X1 U23453 ( .A1(n11393), .A2(n12055), .A3(n9221), .ZN(n11394) );
  NAND2_X1 U23454 ( .A1(n11399), .A2(n11398), .ZN(n11405) );
  OAI22_X1 U23455 ( .A1(n793), .A2(n5507), .B1(n11402), .B2(n11401), .ZN(
        n11404) );
  OAI21_X1 U23456 ( .B1(n11405), .B2(n11404), .A(n11403), .ZN(n11427) );
  NAND3_X1 U23457 ( .A1(n11408), .A2(n11407), .A3(n11411), .ZN(n11413) );
  AND2_X1 U23458 ( .A1(n11410), .A2(n51141), .ZN(n12136) );
  NAND2_X1 U23459 ( .A1(n12136), .A2(n11411), .ZN(n11412) );
  NAND2_X1 U23460 ( .A1(n11413), .A2(n11412), .ZN(n11414) );
  AOI21_X1 U23461 ( .B1(n11415), .B2(n12130), .A(n11414), .ZN(n11426) );
  OAI21_X1 U23462 ( .B1(n11418), .B2(n11417), .A(n11416), .ZN(n11419) );
  NOR2_X1 U23463 ( .A1(n438), .A2(n12129), .ZN(n11420) );
  OAI211_X1 U23464 ( .C1(n12141), .C2(n11420), .A(n12139), .B(n12132), .ZN(
        n11421) );
  OAI21_X1 U23465 ( .B1(n11422), .B2(n12137), .A(n11421), .ZN(n11424) );
  NAND2_X1 U23466 ( .A1(n11424), .A2(n11423), .ZN(n11425) );
  AND2_X1 U23467 ( .A1(n12976), .A2(n14455), .ZN(n11811) );
  OAI211_X1 U23470 ( .C1(n52312), .C2(n2253), .A(n14096), .B(n51383), .ZN(
        n11431) );
  NAND4_X1 U23471 ( .A1(n14097), .A2(n14096), .A3(n14453), .A4(n14454), .ZN(
        n11429) );
  AND3_X1 U23472 ( .A1(n11431), .A2(n11430), .A3(n11429), .ZN(n11437) );
  NOR2_X1 U23473 ( .A1(n12972), .A2(n14103), .ZN(n14452) );
  INV_X1 U23474 ( .A(n14099), .ZN(n14104) );
  OAI21_X1 U23475 ( .B1(n14452), .B2(n11432), .A(n14104), .ZN(n11436) );
  NOR2_X1 U23476 ( .A1(n14107), .A2(n51383), .ZN(n14458) );
  NAND2_X1 U23477 ( .A1(n14458), .A2(n14434), .ZN(n11434) );
  AND2_X1 U23478 ( .A1(n12848), .A2(n11434), .ZN(n11435) );
  XNOR2_X1 U23479 ( .A(n4691), .B(n4916), .ZN(n25013) );
  XNOR2_X1 U23480 ( .A(n4712), .B(n4754), .ZN(n11439) );
  XNOR2_X1 U23481 ( .A(n25013), .B(n11439), .ZN(n34710) );
  INV_X1 U23482 ( .A(n4247), .ZN(n47459) );
  XNOR2_X1 U23483 ( .A(n47459), .B(n4818), .ZN(n41740) );
  INV_X1 U23484 ( .A(n41740), .ZN(n28070) );
  XNOR2_X1 U23485 ( .A(n28070), .B(n4721), .ZN(n33897) );
  XNOR2_X1 U23486 ( .A(n34710), .B(n33897), .ZN(n11440) );
  XNOR2_X1 U23487 ( .A(n4923), .B(n4865), .ZN(n26178) );
  XNOR2_X1 U23488 ( .A(n26178), .B(n4897), .ZN(n34711) );
  XNOR2_X1 U23489 ( .A(n11440), .B(n34711), .ZN(n11441) );
  INV_X1 U23490 ( .A(n45463), .ZN(n24928) );
  XNOR2_X1 U23491 ( .A(n49790), .B(n4788), .ZN(n28071) );
  XNOR2_X1 U23492 ( .A(n24928), .B(n28071), .ZN(n42539) );
  XNOR2_X1 U23493 ( .A(n4934), .B(n4930), .ZN(n34709) );
  XNOR2_X1 U23494 ( .A(n42327), .B(n34709), .ZN(n25284) );
  XNOR2_X1 U23495 ( .A(n42539), .B(n25284), .ZN(n33899) );
  XNOR2_X1 U23496 ( .A(n11441), .B(n33899), .ZN(n11442) );
  XNOR2_X1 U23497 ( .A(n16064), .B(n11442), .ZN(n11563) );
  NOR2_X1 U23498 ( .A1(n12532), .A2(n11443), .ZN(n11444) );
  AOI22_X1 U23499 ( .A1(n9109), .A2(n11446), .B1(n11445), .B2(n11444), .ZN(
        n11451) );
  NAND3_X1 U23500 ( .A1(n12543), .A2(n11447), .A3(n8941), .ZN(n11450) );
  NAND3_X1 U23501 ( .A1(n12546), .A2(n11447), .A3(n12538), .ZN(n11448) );
  AND4_X1 U23502 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(
        n11459) );
  OAI21_X1 U23503 ( .B1(n12536), .B2(n6409), .A(n12533), .ZN(n11453) );
  OAI21_X1 U23504 ( .B1(n11454), .B2(n11453), .A(n11452), .ZN(n11457) );
  NAND2_X1 U23505 ( .A1(n11455), .A2(n12537), .ZN(n11456) );
  NAND2_X1 U23506 ( .A1(n11620), .A2(n11629), .ZN(n11478) );
  NAND2_X1 U23508 ( .A1(n11465), .A2(n11464), .ZN(n11483) );
  OAI211_X1 U23509 ( .C1(n11468), .C2(n11624), .A(n11467), .B(n11466), .ZN(
        n11473) );
  NAND2_X1 U23510 ( .A1(n11476), .A2(n11470), .ZN(n11471) );
  OAI211_X1 U23511 ( .C1(n11474), .C2(n11473), .A(n11472), .B(n11471), .ZN(
        n11475) );
  INV_X1 U23512 ( .A(n11475), .ZN(n11482) );
  AOI22_X1 U23513 ( .A1(n11477), .A2(n4150), .B1(n11620), .B2(n11476), .ZN(
        n11481) );
  INV_X1 U23514 ( .A(n11478), .ZN(n11479) );
  NAND2_X1 U23515 ( .A1(n11479), .A2(n11635), .ZN(n11480) );
  INV_X1 U23516 ( .A(n15363), .ZN(n14492) );
  NOR2_X1 U23517 ( .A1(n11485), .A2(n11903), .ZN(n11486) );
  NAND2_X1 U23518 ( .A1(n5251), .A2(n11488), .ZN(n12473) );
  OAI211_X1 U23519 ( .C1(n2116), .C2(n11489), .A(n12473), .B(n12471), .ZN(
        n11490) );
  NAND2_X1 U23520 ( .A1(n12454), .A2(n11874), .ZN(n12669) );
  OAI211_X1 U23521 ( .C1(n12680), .C2(n8901), .A(n11499), .B(n12669), .ZN(
        n11491) );
  NAND2_X1 U23522 ( .A1(n12673), .A2(n50997), .ZN(n11494) );
  NAND2_X1 U23523 ( .A1(n11874), .A2(n592), .ZN(n11888) );
  NAND2_X1 U23524 ( .A1(n12671), .A2(n12451), .ZN(n11492) );
  NAND2_X1 U23527 ( .A1(n50997), .A2(n592), .ZN(n11875) );
  NAND4_X1 U23528 ( .A1(n11498), .A2(n11497), .A3(n12667), .A4(n12676), .ZN(
        n11505) );
  INV_X1 U23529 ( .A(n11499), .ZN(n11873) );
  OAI211_X1 U23530 ( .C1(n11501), .C2(n11500), .A(n11884), .B(n7354), .ZN(
        n11502) );
  OAI21_X1 U23531 ( .B1(n11873), .B2(n12675), .A(n11503), .ZN(n11504) );
  NAND2_X1 U23532 ( .A1(n14492), .A2(n14484), .ZN(n11554) );
  OR2_X1 U23533 ( .A1(n15385), .A2(n15358), .ZN(n14809) );
  NAND2_X1 U23534 ( .A1(n11508), .A2(n51760), .ZN(n11509) );
  NOR2_X1 U23535 ( .A1(n11510), .A2(n11509), .ZN(n12561) );
  NOR2_X1 U23536 ( .A1(n11573), .A2(n12557), .ZN(n11511) );
  NOR2_X1 U23537 ( .A1(n12561), .A2(n11511), .ZN(n11524) );
  OAI21_X1 U23538 ( .B1(n12558), .B2(n11568), .A(n11512), .ZN(n11513) );
  NAND2_X1 U23539 ( .A1(n11513), .A2(n51491), .ZN(n11523) );
  NAND3_X1 U23540 ( .A1(n51760), .A2(n11581), .A3(n11514), .ZN(n11516) );
  OAI21_X1 U23541 ( .B1(n11567), .B2(n11581), .A(n11516), .ZN(n11518) );
  NAND2_X1 U23542 ( .A1(n11516), .A2(n51760), .ZN(n11517) );
  NAND3_X1 U23543 ( .A1(n11518), .A2(n12570), .A3(n11517), .ZN(n11522) );
  AND2_X1 U23544 ( .A1(n12555), .A2(n11530), .ZN(n11580) );
  NAND3_X1 U23545 ( .A1(n11525), .A2(n11580), .A3(n11581), .ZN(n11527) );
  NAND3_X1 U23546 ( .A1(n12577), .A2(n11582), .A3(n12559), .ZN(n11526) );
  OAI211_X1 U23547 ( .C1(n11529), .C2(n11528), .A(n11527), .B(n11526), .ZN(
        n11535) );
  NAND2_X1 U23548 ( .A1(n12557), .A2(n11530), .ZN(n11533) );
  NAND3_X1 U23549 ( .A1(n11579), .A2(n12556), .A3(n12559), .ZN(n11531) );
  OAI21_X1 U23550 ( .B1(n11533), .B2(n11532), .A(n11531), .ZN(n11534) );
  MUX2_X1 U23551 ( .A(n11554), .B(n14809), .S(n51984), .Z(n11562) );
  OAI21_X1 U23552 ( .B1(n11537), .B2(n12500), .A(n8024), .ZN(n11542) );
  NAND2_X1 U23553 ( .A1(n12506), .A2(n12514), .ZN(n12501) );
  AOI22_X1 U23554 ( .A1(n11540), .A2(n11539), .B1(n642), .B2(n12516), .ZN(
        n11541) );
  INV_X1 U23555 ( .A(n12501), .ZN(n11547) );
  NAND3_X1 U23557 ( .A1(n11549), .A2(n11548), .A3(n12498), .ZN(n11551) );
  NAND2_X1 U23558 ( .A1(n11551), .A2(n11550), .ZN(n14812) );
  INV_X1 U23559 ( .A(n15384), .ZN(n15381) );
  INV_X1 U23560 ( .A(n13914), .ZN(n11552) );
  NAND2_X1 U23561 ( .A1(n11853), .A2(n15380), .ZN(n11555) );
  OAI211_X1 U23562 ( .C1(n13916), .C2(n15381), .A(n14806), .B(n11555), .ZN(
        n11553) );
  INV_X1 U23563 ( .A(n11554), .ZN(n11557) );
  INV_X1 U23564 ( .A(n11555), .ZN(n11556) );
  AND2_X1 U23565 ( .A1(n15386), .A2(n15381), .ZN(n14489) );
  OAI21_X1 U23566 ( .B1(n11557), .B2(n11556), .A(n14489), .ZN(n11560) );
  OAI21_X1 U23567 ( .B1(n15382), .B2(n15378), .A(n14488), .ZN(n11559) );
  NAND4_X2 U23568 ( .A1(n11562), .A2(n11560), .A3(n11561), .A4(n11559), .ZN(
        n17831) );
  XNOR2_X1 U23569 ( .A(n11563), .B(n17831), .ZN(n11564) );
  XNOR2_X1 U23570 ( .A(n15609), .B(n11564), .ZN(n11773) );
  NAND2_X1 U23571 ( .A1(n11566), .A2(n11565), .ZN(n11578) );
  INV_X1 U23572 ( .A(n12557), .ZN(n12568) );
  NAND2_X1 U23573 ( .A1(n11569), .A2(n11568), .ZN(n11571) );
  AOI22_X1 U23574 ( .A1(n11572), .A2(n11571), .B1(n12577), .B2(n11570), .ZN(
        n11577) );
  INV_X1 U23575 ( .A(n11573), .ZN(n11574) );
  NAND2_X1 U23576 ( .A1(n11574), .A2(n11579), .ZN(n12563) );
  NAND4_X1 U23577 ( .A1(n11578), .A2(n11577), .A3(n12563), .A4(n11576), .ZN(
        n11587) );
  NAND2_X1 U23578 ( .A1(n11579), .A2(n12578), .ZN(n11585) );
  INV_X1 U23579 ( .A(n11580), .ZN(n11583) );
  NAND3_X1 U23580 ( .A1(n11583), .A2(n11582), .A3(n11581), .ZN(n11584) );
  AOI21_X1 U23581 ( .B1(n11585), .B2(n12570), .A(n11584), .ZN(n11586) );
  INV_X1 U23582 ( .A(n11723), .ZN(n14519) );
  NAND3_X1 U23583 ( .A1(n11589), .A2(n11590), .A3(n11588), .ZN(n11597) );
  NAND3_X1 U23584 ( .A1(n11600), .A2(n11593), .A3(n11608), .ZN(n11594) );
  NAND4_X1 U23585 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11607) );
  NAND3_X1 U23586 ( .A1(n11602), .A2(n11601), .A3(n11600), .ZN(n11603) );
  OAI21_X1 U23587 ( .B1(n11605), .B2(n11604), .A(n11603), .ZN(n11606) );
  NAND2_X1 U23588 ( .A1(n11610), .A2(n11608), .ZN(n11609) );
  OAI21_X1 U23589 ( .B1(n11611), .B2(n11610), .A(n11609), .ZN(n11617) );
  AND3_X1 U23590 ( .A1(n11614), .A2(n11613), .A3(n11612), .ZN(n11616) );
  MUX2_X1 U23591 ( .A(n11617), .B(n11616), .S(n11615), .Z(n11618) );
  NAND2_X1 U23592 ( .A1(n11620), .A2(n11619), .ZN(n11623) );
  NAND3_X1 U23593 ( .A1(n11635), .A2(n11621), .A3(n454), .ZN(n11622) );
  OAI211_X1 U23594 ( .C1(n11625), .C2(n11624), .A(n11623), .B(n11622), .ZN(
        n11626) );
  INV_X1 U23595 ( .A(n11626), .ZN(n11638) );
  NAND2_X1 U23596 ( .A1(n11627), .A2(n11634), .ZN(n11637) );
  NAND4_X1 U23597 ( .A1(n11644), .A2(n11643), .A3(n11642), .A4(n11660), .ZN(
        n11645) );
  AND2_X1 U23598 ( .A1(n11645), .A2(n11646), .ZN(n11666) );
  NAND3_X1 U23599 ( .A1(n11648), .A2(n11655), .A3(n11647), .ZN(n11653) );
  NAND2_X1 U23600 ( .A1(n11663), .A2(n11649), .ZN(n11652) );
  NAND3_X1 U23601 ( .A1(n11655), .A2(n11654), .A3(n5917), .ZN(n11656) );
  AND2_X1 U23602 ( .A1(n11657), .A2(n11656), .ZN(n11665) );
  INV_X1 U23603 ( .A(n11658), .ZN(n11659) );
  OAI211_X1 U23604 ( .C1(n11663), .C2(n11662), .A(n11661), .B(n11660), .ZN(
        n11664) );
  NAND2_X1 U23605 ( .A1(n13384), .A2(n14515), .ZN(n11667) );
  NOR2_X1 U23606 ( .A1(n13034), .A2(n11667), .ZN(n13376) );
  AOI22_X1 U23607 ( .A1(n11673), .A2(n11682), .B1(n11672), .B2(n11671), .ZN(
        n11678) );
  NOR2_X1 U23608 ( .A1(n11674), .A2(n11687), .ZN(n11675) );
  OAI21_X1 U23609 ( .B1(n11676), .B2(n11675), .A(n9973), .ZN(n11677) );
  MUX2_X1 U23610 ( .A(n11681), .B(n11680), .S(n11679), .Z(n11692) );
  INV_X1 U23611 ( .A(n11686), .ZN(n11689) );
  NAND3_X1 U23612 ( .A1(n11689), .A2(n11688), .A3(n11687), .ZN(n11690) );
  NAND2_X1 U23615 ( .A1(n51650), .A2(n643), .ZN(n11700) );
  OAI21_X1 U23616 ( .B1(n11701), .B2(n11700), .A(n11699), .ZN(n11702) );
  NOR2_X1 U23617 ( .A1(n11703), .A2(n11702), .ZN(n11719) );
  NOR2_X1 U23618 ( .A1(n11705), .A2(n11704), .ZN(n11708) );
  OAI211_X1 U23619 ( .C1(n11709), .C2(n11708), .A(n11707), .B(n11706), .ZN(
        n11718) );
  NAND2_X1 U23620 ( .A1(n11712), .A2(n11711), .ZN(n11717) );
  NAND3_X1 U23621 ( .A1(n11715), .A2(n11714), .A3(n51650), .ZN(n11716) );
  OAI211_X1 U23622 ( .C1(n51019), .C2(n13384), .A(n14515), .B(n16036), .ZN(
        n11720) );
  NAND2_X1 U23623 ( .A1(n13033), .A2(n11720), .ZN(n11729) );
  AND2_X1 U23624 ( .A1(n16049), .A2(n13377), .ZN(n13387) );
  INV_X1 U23625 ( .A(n13387), .ZN(n11722) );
  AND2_X1 U23626 ( .A1(n14519), .A2(n51714), .ZN(n12813) );
  INV_X1 U23627 ( .A(n12813), .ZN(n11721) );
  AOI21_X1 U23628 ( .B1(n13372), .B2(n11722), .A(n11721), .ZN(n11726) );
  INV_X1 U23630 ( .A(n16045), .ZN(n11724) );
  AND2_X1 U23631 ( .A1(n13377), .A2(n51713), .ZN(n16043) );
  INV_X1 U23632 ( .A(n16043), .ZN(n16048) );
  OAI22_X1 U23633 ( .A1(n14516), .A2(n11724), .B1(n13040), .B2(n16048), .ZN(
        n11725) );
  NOR2_X1 U23634 ( .A1(n11726), .A2(n11725), .ZN(n11728) );
  OAI21_X1 U23635 ( .B1(n13384), .B2(n51714), .A(n51019), .ZN(n16038) );
  NOR2_X1 U23636 ( .A1(n16039), .A2(n14515), .ZN(n13370) );
  MUX2_X1 U23637 ( .A(n16038), .B(n13371), .S(n13370), .Z(n11727) );
  INV_X1 U23638 ( .A(n11730), .ZN(n11731) );
  NAND2_X1 U23639 ( .A1(n14472), .A2(n11731), .ZN(n11733) );
  NOR2_X1 U23640 ( .A1(n11733), .A2(n11732), .ZN(n14884) );
  INV_X1 U23641 ( .A(n14884), .ZN(n14471) );
  OR2_X1 U23642 ( .A1(n14482), .A2(n14473), .ZN(n14478) );
  INV_X1 U23643 ( .A(n14478), .ZN(n11734) );
  NAND2_X1 U23644 ( .A1(n13849), .A2(n14472), .ZN(n11736) );
  NOR2_X1 U23645 ( .A1(n11736), .A2(n13855), .ZN(n11739) );
  OR2_X1 U23646 ( .A1(n11738), .A2(n11737), .ZN(n13548) );
  INV_X1 U23647 ( .A(n13548), .ZN(n11781) );
  OAI21_X1 U23648 ( .B1(n13560), .B2(n11739), .A(n11781), .ZN(n11747) );
  NAND2_X1 U23649 ( .A1(n11741), .A2(n14883), .ZN(n11746) );
  NOR2_X1 U23650 ( .A1(n14473), .A2(n13849), .ZN(n11742) );
  AOI21_X1 U23651 ( .B1(n11742), .B2(n13841), .A(n13845), .ZN(n11743) );
  NAND2_X1 U23652 ( .A1(n13841), .A2(n13845), .ZN(n13551) );
  NAND2_X1 U23653 ( .A1(n11744), .A2(n13551), .ZN(n11745) );
  NAND4_X1 U23654 ( .A1(n11748), .A2(n11747), .A3(n11746), .A4(n11745), .ZN(
        n16559) );
  XNOR2_X1 U23655 ( .A(n8699), .B(n16559), .ZN(n16063) );
  NAND2_X1 U23656 ( .A1(n12894), .A2(n13432), .ZN(n12042) );
  INV_X1 U23657 ( .A(n12042), .ZN(n11749) );
  NAND2_X1 U23658 ( .A1(n12799), .A2(n11749), .ZN(n11751) );
  NAND2_X1 U23659 ( .A1(n12794), .A2(n13449), .ZN(n11750) );
  INV_X1 U23660 ( .A(n13445), .ZN(n11753) );
  NAND3_X1 U23661 ( .A1(n12786), .A2(n13450), .A3(n12791), .ZN(n11755) );
  AND2_X1 U23662 ( .A1(n13450), .A2(n483), .ZN(n12039) );
  NAND3_X1 U23663 ( .A1(n12039), .A2(n13995), .A3(n4383), .ZN(n11754) );
  AND2_X1 U23664 ( .A1(n11755), .A2(n11754), .ZN(n11758) );
  AND2_X1 U23665 ( .A1(n12787), .A2(n12893), .ZN(n14656) );
  OAI21_X1 U23666 ( .B1(n12888), .B2(n14657), .A(n786), .ZN(n11756) );
  INV_X1 U23667 ( .A(n11756), .ZN(n11757) );
  NOR2_X1 U23668 ( .A1(n13949), .A2(n13948), .ZN(n13197) );
  NAND2_X1 U23669 ( .A1(n13197), .A2(n6668), .ZN(n12880) );
  INV_X1 U23670 ( .A(n11759), .ZN(n11760) );
  NAND2_X1 U23671 ( .A1(n11760), .A2(n13941), .ZN(n11761) );
  NAND2_X1 U23672 ( .A1(n13948), .A2(n51656), .ZN(n13189) );
  NAND2_X1 U23673 ( .A1(n13947), .A2(n13207), .ZN(n11762) );
  NAND2_X1 U23674 ( .A1(n13947), .A2(n2173), .ZN(n12886) );
  NOR3_X1 U23675 ( .A1(n12886), .A2(n13933), .A3(n13930), .ZN(n11764) );
  NOR2_X1 U23678 ( .A1(n11764), .A2(n13946), .ZN(n11770) );
  INV_X1 U23679 ( .A(n13204), .ZN(n11768) );
  INV_X1 U23680 ( .A(n11865), .ZN(n13193) );
  NOR2_X1 U23681 ( .A1(n12882), .A2(n13193), .ZN(n11767) );
  NAND2_X1 U23682 ( .A1(n11765), .A2(n2173), .ZN(n11766) );
  XNOR2_X1 U23683 ( .A(n15876), .B(n16063), .ZN(n11772) );
  XNOR2_X1 U23684 ( .A(n11773), .B(n11772), .ZN(n11774) );
  XNOR2_X1 U23685 ( .A(n16392), .B(n11774), .ZN(n13540) );
  AOI22_X1 U23686 ( .A1(n13853), .A2(n11781), .B1(n14477), .B2(n13855), .ZN(
        n11785) );
  NOR2_X1 U23687 ( .A1(n13841), .A2(n14482), .ZN(n13851) );
  INV_X1 U23688 ( .A(n13851), .ZN(n11777) );
  OR2_X1 U23689 ( .A1(n13841), .A2(n13845), .ZN(n14479) );
  NAND2_X1 U23690 ( .A1(n13856), .A2(n13849), .ZN(n14474) );
  INV_X1 U23691 ( .A(n13560), .ZN(n11775) );
  OAI21_X1 U23692 ( .B1(n14479), .B2(n14474), .A(n11775), .ZN(n11776) );
  AOI21_X1 U23693 ( .B1(n11778), .B2(n11777), .A(n11776), .ZN(n11784) );
  AND2_X1 U23694 ( .A1(n13841), .A2(n13855), .ZN(n13850) );
  AND2_X1 U23695 ( .A1(n14482), .A2(n13854), .ZN(n11779) );
  AOI22_X1 U23696 ( .A1(n11781), .A2(n11780), .B1(n13850), .B2(n11779), .ZN(
        n11783) );
  NOR2_X1 U23697 ( .A1(n13841), .A2(n14473), .ZN(n14885) );
  INV_X1 U23698 ( .A(n14885), .ZN(n14480) );
  NOR2_X1 U23699 ( .A1(n14480), .A2(n13845), .ZN(n14889) );
  NAND2_X1 U23700 ( .A1(n14889), .A2(n14883), .ZN(n11782) );
  NAND4_X2 U23701 ( .A1(n11785), .A2(n11784), .A3(n11783), .A4(n11782), .ZN(
        n18827) );
  NAND2_X1 U23702 ( .A1(n14285), .A2(n14287), .ZN(n14296) );
  NAND2_X1 U23703 ( .A1(n13583), .A2(n14294), .ZN(n14277) );
  NAND2_X1 U23704 ( .A1(n14296), .A2(n14277), .ZN(n13011) );
  INV_X1 U23705 ( .A(n14290), .ZN(n11786) );
  NAND2_X1 U23706 ( .A1(n13011), .A2(n11786), .ZN(n11793) );
  INV_X1 U23707 ( .A(n14288), .ZN(n11788) );
  INV_X1 U23708 ( .A(n14289), .ZN(n14298) );
  OAI21_X1 U23709 ( .B1(n11788), .B2(n13576), .A(n14298), .ZN(n11792) );
  NOR2_X1 U23713 ( .A1(n14315), .A2(n14320), .ZN(n11795) );
  NOR2_X1 U23714 ( .A1(n11796), .A2(n14320), .ZN(n13831) );
  NAND2_X1 U23715 ( .A1(n13831), .A2(n13819), .ZN(n11800) );
  AND2_X1 U23716 ( .A1(n14318), .A2(n14307), .ZN(n13600) );
  NOR2_X1 U23717 ( .A1(n11798), .A2(n14311), .ZN(n14308) );
  OAI21_X1 U23718 ( .B1(n14318), .B2(n14307), .A(n14308), .ZN(n11799) );
  XNOR2_X1 U23719 ( .A(n563), .B(n19186), .ZN(n16345) );
  INV_X1 U23720 ( .A(n13488), .ZN(n11802) );
  INV_X1 U23721 ( .A(n15033), .ZN(n11801) );
  INV_X1 U23722 ( .A(n13797), .ZN(n15035) );
  NOR2_X1 U23723 ( .A1(n15035), .A2(n15034), .ZN(n12777) );
  INV_X1 U23724 ( .A(n13806), .ZN(n11803) );
  NOR2_X1 U23725 ( .A1(n15046), .A2(n13483), .ZN(n13481) );
  AND2_X1 U23726 ( .A1(n13797), .A2(n13801), .ZN(n12780) );
  NAND3_X1 U23727 ( .A1(n13798), .A2(n277), .A3(n13483), .ZN(n11808) );
  NOR2_X1 U23728 ( .A1(n15046), .A2(n13800), .ZN(n15038) );
  NAND2_X1 U23729 ( .A1(n15033), .A2(n15046), .ZN(n11805) );
  OAI211_X1 U23730 ( .C1(n15038), .C2(n15048), .A(n11806), .B(n11805), .ZN(
        n11807) );
  OR2_X1 U23731 ( .A1(n14103), .A2(n14444), .ZN(n14448) );
  INV_X1 U23732 ( .A(n14448), .ZN(n11809) );
  AND2_X1 U23733 ( .A1(n12848), .A2(n11810), .ZN(n11818) );
  INV_X1 U23734 ( .A(n11811), .ZN(n11812) );
  NAND3_X1 U23735 ( .A1(n11812), .A2(n51383), .A3(n14102), .ZN(n11817) );
  NAND2_X1 U23736 ( .A1(n11813), .A2(n14455), .ZN(n12856) );
  OR2_X1 U23737 ( .A1(n51383), .A2(n14444), .ZN(n14101) );
  INV_X1 U23738 ( .A(n14101), .ZN(n11814) );
  OAI21_X1 U23739 ( .B1(n12856), .B2(n11814), .A(n52312), .ZN(n11816) );
  OAI21_X1 U23740 ( .B1(n14434), .B2(n14097), .A(n14095), .ZN(n11815) );
  XNOR2_X1 U23741 ( .A(n16435), .B(n51703), .ZN(n15711) );
  OAI21_X1 U23742 ( .B1(n13091), .B2(n13104), .A(n11820), .ZN(n11822) );
  NAND2_X1 U23743 ( .A1(n11822), .A2(n11821), .ZN(n11828) );
  NOR2_X1 U23744 ( .A1(n13086), .A2(n13089), .ZN(n11823) );
  NOR2_X1 U23745 ( .A1(n13089), .A2(n12914), .ZN(n13093) );
  NAND2_X1 U23746 ( .A1(n13093), .A2(n13092), .ZN(n12818) );
  OAI22_X1 U23747 ( .A1(n13104), .A2(n13088), .B1(n13092), .B2(n11825), .ZN(
        n11826) );
  NAND2_X1 U23748 ( .A1(n11826), .A2(n13086), .ZN(n11827) );
  XNOR2_X1 U23749 ( .A(n4048), .B(n4845), .ZN(n26586) );
  XNOR2_X1 U23750 ( .A(n42889), .B(n26586), .ZN(n17950) );
  XNOR2_X1 U23751 ( .A(n17950), .B(n4026), .ZN(n33467) );
  XNOR2_X1 U23752 ( .A(n48814), .B(n4737), .ZN(n21828) );
  XNOR2_X1 U23753 ( .A(n6031), .B(n4864), .ZN(n25183) );
  XNOR2_X1 U23754 ( .A(n21828), .B(n25183), .ZN(n24127) );
  XNOR2_X1 U23755 ( .A(n4526), .B(n47679), .ZN(n28085) );
  XNOR2_X1 U23756 ( .A(n24127), .B(n28085), .ZN(n35604) );
  XNOR2_X1 U23757 ( .A(n33467), .B(n35604), .ZN(n11829) );
  XNOR2_X1 U23758 ( .A(n4585), .B(n4733), .ZN(n44952) );
  XNOR2_X1 U23759 ( .A(n4628), .B(n4599), .ZN(n43263) );
  XNOR2_X1 U23760 ( .A(n44952), .B(n2601), .ZN(n34377) );
  XNOR2_X1 U23761 ( .A(n4835), .B(n4317), .ZN(n27297) );
  XNOR2_X1 U23762 ( .A(n27297), .B(n4471), .ZN(n16777) );
  XNOR2_X1 U23763 ( .A(n34377), .B(n16777), .ZN(n40107) );
  XNOR2_X1 U23764 ( .A(n11829), .B(n40107), .ZN(n11830) );
  XNOR2_X1 U23765 ( .A(n18690), .B(n11830), .ZN(n11831) );
  XNOR2_X1 U23766 ( .A(n15711), .B(n11831), .ZN(n11832) );
  XNOR2_X1 U23767 ( .A(n16345), .B(n11832), .ZN(n12006) );
  AND2_X1 U23768 ( .A1(n13221), .A2(n14224), .ZN(n14223) );
  INV_X1 U23769 ( .A(n13220), .ZN(n11835) );
  INV_X1 U23770 ( .A(n13222), .ZN(n11834) );
  NAND2_X1 U23771 ( .A1(n14224), .A2(n13970), .ZN(n11833) );
  INV_X1 U23772 ( .A(n13960), .ZN(n13247) );
  OAI211_X1 U23773 ( .C1(n13247), .C2(n13970), .A(n13971), .B(n14234), .ZN(
        n11839) );
  OR2_X1 U23774 ( .A1(n13971), .A2(n14234), .ZN(n13244) );
  AND2_X1 U23775 ( .A1(n13219), .A2(n14234), .ZN(n12922) );
  NAND2_X1 U23776 ( .A1(n12922), .A2(n14224), .ZN(n14230) );
  NAND3_X1 U23777 ( .A1(n13226), .A2(n14234), .A3(n639), .ZN(n11836) );
  NAND2_X1 U23778 ( .A1(n14230), .A2(n11836), .ZN(n11837) );
  NAND2_X1 U23779 ( .A1(n11837), .A2(n13971), .ZN(n11838) );
  NAND2_X1 U23780 ( .A1(n12765), .A2(n12767), .ZN(n11850) );
  INV_X1 U23781 ( .A(n13513), .ZN(n13511) );
  AOI22_X1 U23782 ( .A1(n13515), .A2(n13511), .B1(n13509), .B2(n12938), .ZN(
        n11849) );
  NOR2_X1 U23783 ( .A1(n11841), .A2(n13526), .ZN(n13522) );
  NAND2_X1 U23784 ( .A1(n13514), .A2(n51683), .ZN(n11842) );
  AND2_X1 U23785 ( .A1(n51066), .A2(n11842), .ZN(n13496) );
  OAI21_X1 U23786 ( .B1(n13505), .B2(n13522), .A(n13496), .ZN(n11848) );
  INV_X1 U23787 ( .A(n11843), .ZN(n11846) );
  NOR2_X1 U23788 ( .A1(n13514), .A2(n13526), .ZN(n11844) );
  NAND3_X1 U23789 ( .A1(n955), .A2(n13501), .A3(n51683), .ZN(n12766) );
  OAI211_X1 U23790 ( .C1(n11846), .C2(n11845), .A(n11844), .B(n12766), .ZN(
        n11847) );
  XNOR2_X1 U23791 ( .A(n16571), .B(n17730), .ZN(n11858) );
  AOI21_X1 U23792 ( .B1(n11853), .B2(n15367), .A(n15363), .ZN(n11851) );
  AND2_X1 U23793 ( .A1(n11853), .A2(n15386), .ZN(n15374) );
  NAND3_X1 U23794 ( .A1(n15374), .A2(n787), .A3(n15358), .ZN(n11857) );
  NAND2_X1 U23795 ( .A1(n15386), .A2(n15384), .ZN(n14808) );
  NAND3_X1 U23796 ( .A1(n14808), .A2(n14492), .A3(n14484), .ZN(n11856) );
  OAI21_X1 U23797 ( .B1(n14485), .B2(n15385), .A(n11853), .ZN(n11854) );
  NAND2_X1 U23798 ( .A1(n11854), .A2(n15384), .ZN(n11855) );
  XNOR2_X1 U23799 ( .A(n11858), .B(n17947), .ZN(n17841) );
  INV_X1 U23800 ( .A(n13208), .ZN(n11859) );
  NOR2_X1 U23801 ( .A1(n13946), .A2(n11861), .ZN(n11868) );
  INV_X1 U23802 ( .A(n11862), .ZN(n11863) );
  OAI211_X1 U23803 ( .C1(n13206), .C2(n11863), .A(n13190), .B(n13197), .ZN(
        n11867) );
  INV_X1 U23804 ( .A(n12881), .ZN(n11864) );
  OAI21_X1 U23805 ( .B1(n781), .B2(n11865), .A(n11864), .ZN(n11866) );
  OAI21_X1 U23806 ( .B1(n11871), .B2(n592), .A(n11870), .ZN(n13895) );
  NAND2_X1 U23808 ( .A1(n12455), .A2(n11879), .ZN(n12687) );
  NAND3_X1 U23810 ( .A1(n12671), .A2(n12675), .A3(n11874), .ZN(n11877) );
  NAND4_X1 U23811 ( .A1(n12687), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(
        n13897) );
  INV_X1 U23812 ( .A(n13897), .ZN(n11892) );
  NAND2_X1 U23814 ( .A1(n11883), .A2(n11882), .ZN(n11887) );
  NAND3_X1 U23815 ( .A1(n11884), .A2(n11500), .A3(n12676), .ZN(n11885) );
  AOI21_X1 U23816 ( .B1(n11885), .B2(n12675), .A(n592), .ZN(n11886) );
  NAND2_X1 U23817 ( .A1(n11887), .A2(n11886), .ZN(n13894) );
  INV_X1 U23818 ( .A(n11888), .ZN(n11889) );
  NAND2_X1 U23819 ( .A1(n11889), .A2(n12675), .ZN(n11891) );
  MUX2_X1 U23820 ( .A(n11891), .B(n11890), .S(n12673), .Z(n13896) );
  AND2_X1 U23821 ( .A1(n12491), .A2(n11893), .ZN(n11911) );
  OAI21_X1 U23822 ( .B1(n11900), .B2(n12470), .A(n510), .ZN(n11901) );
  NAND2_X1 U23823 ( .A1(n11902), .A2(n11901), .ZN(n11910) );
  INV_X1 U23824 ( .A(n12486), .ZN(n11905) );
  AOI21_X1 U23825 ( .B1(n11903), .B2(n12470), .A(n2116), .ZN(n11904) );
  OAI21_X1 U23826 ( .B1(n11905), .B2(n12480), .A(n11904), .ZN(n11906) );
  OAI211_X1 U23827 ( .C1(n11908), .C2(n2211), .A(n11906), .B(n12481), .ZN(
        n11909) );
  INV_X1 U23828 ( .A(n11912), .ZN(n11913) );
  NAND3_X1 U23829 ( .A1(n795), .A2(n11915), .A3(n11920), .ZN(n11916) );
  NAND4_X1 U23830 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11925) );
  NAND2_X1 U23831 ( .A1(n12589), .A2(n11920), .ZN(n12609) );
  INV_X1 U23832 ( .A(n11922), .ZN(n11923) );
  OAI22_X1 U23833 ( .A1(n12609), .A2(n12605), .B1(n11923), .B2(n1307), .ZN(
        n11924) );
  NOR2_X1 U23834 ( .A1(n12701), .A2(n12711), .ZN(n12437) );
  INV_X1 U23835 ( .A(n12444), .ZN(n11927) );
  OAI21_X1 U23836 ( .B1(n11928), .B2(n11927), .A(n12689), .ZN(n11939) );
  NOR2_X1 U23837 ( .A1(n12705), .A2(n12709), .ZN(n11929) );
  OAI21_X1 U23838 ( .B1(n11930), .B2(n11929), .A(n12440), .ZN(n11936) );
  NAND2_X1 U23839 ( .A1(n2156), .A2(n11931), .ZN(n11935) );
  NAND3_X1 U23840 ( .A1(n12696), .A2(n11933), .A3(n12704), .ZN(n11934) );
  NAND4_X1 U23841 ( .A1(n11937), .A2(n11936), .A3(n11935), .A4(n11934), .ZN(
        n11938) );
  AND2_X1 U23843 ( .A1(n11943), .A2(n11941), .ZN(n12721) );
  INV_X1 U23844 ( .A(n12721), .ZN(n11945) );
  AND2_X1 U23845 ( .A1(n11942), .A2(n8881), .ZN(n11962) );
  NAND2_X1 U23846 ( .A1(n11962), .A2(n11943), .ZN(n11944) );
  AOI21_X1 U23847 ( .B1(n11945), .B2(n11944), .A(n11964), .ZN(n11953) );
  INV_X1 U23848 ( .A(n11946), .ZN(n11947) );
  NAND2_X1 U23849 ( .A1(n12722), .A2(n11947), .ZN(n11949) );
  NOR2_X1 U23850 ( .A1(n11953), .A2(n11952), .ZN(n11970) );
  NAND3_X1 U23851 ( .A1(n11955), .A2(n12718), .A3(n11954), .ZN(n11969) );
  INV_X1 U23852 ( .A(n11956), .ZN(n12723) );
  NOR2_X1 U23853 ( .A1(n12723), .A2(n11957), .ZN(n11959) );
  OAI21_X1 U23854 ( .B1(n11960), .B2(n11959), .A(n11958), .ZN(n11968) );
  INV_X1 U23855 ( .A(n11961), .ZN(n11966) );
  INV_X1 U23856 ( .A(n11962), .ZN(n11963) );
  NOR2_X1 U23857 ( .A1(n12729), .A2(n11963), .ZN(n11965) );
  OAI21_X1 U23858 ( .B1(n11966), .B2(n11965), .A(n11964), .ZN(n11967) );
  NAND4_X2 U23859 ( .A1(n11970), .A2(n11969), .A3(n11967), .A4(n11968), .ZN(
        n15438) );
  NOR2_X1 U23860 ( .A1(n12657), .A2(n11973), .ZN(n11975) );
  AOI22_X1 U23861 ( .A1(n11976), .A2(n11975), .B1(n11974), .B2(n12652), .ZN(
        n11990) );
  INV_X1 U23862 ( .A(n11977), .ZN(n11983) );
  OAI211_X1 U23863 ( .C1(n11979), .C2(n12648), .A(n11978), .B(n12649), .ZN(
        n11980) );
  INV_X1 U23864 ( .A(n11980), .ZN(n11981) );
  OAI21_X1 U23865 ( .B1(n11983), .B2(n11982), .A(n11981), .ZN(n11989) );
  OAI21_X1 U23866 ( .B1(n9188), .B2(n11984), .A(n794), .ZN(n11987) );
  NAND4_X1 U23867 ( .A1(n11987), .A2(n2227), .A3(n11986), .A4(n11985), .ZN(
        n11988) );
  NAND2_X1 U23869 ( .A1(n15434), .A2(n15341), .ZN(n15334) );
  NAND2_X1 U23870 ( .A1(n15435), .A2(n15440), .ZN(n14828) );
  NAND2_X1 U23871 ( .A1(n15325), .A2(n15448), .ZN(n11992) );
  OAI22_X1 U23872 ( .A1(n15438), .A2(n14828), .B1(n11992), .B2(n15437), .ZN(
        n11993) );
  NOR2_X1 U23873 ( .A1(n14408), .A2(n14412), .ZN(n14073) );
  NAND3_X1 U23874 ( .A1(n14073), .A2(n12961), .A3(n11999), .ZN(n11995) );
  INV_X1 U23875 ( .A(n14393), .ZN(n12865) );
  NAND2_X1 U23876 ( .A1(n12865), .A2(n14070), .ZN(n12966) );
  INV_X1 U23877 ( .A(n12966), .ZN(n14417) );
  AND2_X1 U23878 ( .A1(n14412), .A2(n14072), .ZN(n14415) );
  NAND2_X1 U23879 ( .A1(n14417), .A2(n14415), .ZN(n11994) );
  AND2_X1 U23880 ( .A1(n11995), .A2(n11994), .ZN(n12004) );
  NAND2_X1 U23881 ( .A1(n14393), .A2(n14070), .ZN(n14066) );
  INV_X1 U23882 ( .A(n14066), .ZN(n11997) );
  NOR2_X1 U23883 ( .A1(n12963), .A2(n14410), .ZN(n11996) );
  AOI22_X1 U23884 ( .A1(n12872), .A2(n11998), .B1(n11997), .B2(n11996), .ZN(
        n12003) );
  OAI21_X1 U23885 ( .B1(n14068), .B2(n12871), .A(n12872), .ZN(n12002) );
  OAI21_X1 U23886 ( .B1(n11999), .B2(n14408), .A(n14412), .ZN(n12000) );
  NAND2_X1 U23887 ( .A1(n12000), .A2(n14410), .ZN(n12001) );
  XNOR2_X1 U23888 ( .A(n17389), .B(n4676), .ZN(n15536) );
  XNOR2_X1 U23889 ( .A(n18480), .B(n15536), .ZN(n12005) );
  XNOR2_X1 U23890 ( .A(n12005), .B(n17841), .ZN(n16948) );
  XNOR2_X1 U23891 ( .A(n16948), .B(n12006), .ZN(n12195) );
  NAND2_X1 U23892 ( .A1(n14346), .A2(n13003), .ZN(n12229) );
  AOI21_X1 U23893 ( .B1(n14341), .B2(n13417), .A(n14339), .ZN(n12008) );
  AND2_X1 U23894 ( .A1(n14345), .A2(n13410), .ZN(n14338) );
  OAI21_X1 U23895 ( .B1(n12229), .B2(n12008), .A(n14338), .ZN(n12011) );
  NAND2_X1 U23896 ( .A1(n14344), .A2(n14341), .ZN(n14333) );
  NAND2_X1 U23897 ( .A1(n14353), .A2(n14333), .ZN(n12009) );
  INV_X1 U23898 ( .A(n13418), .ZN(n13400) );
  NAND2_X1 U23899 ( .A1(n12009), .A2(n13400), .ZN(n12010) );
  MUX2_X1 U23900 ( .A(n13161), .B(n13774), .S(n13166), .Z(n12015) );
  OR2_X1 U23901 ( .A1(n12013), .A2(n13773), .ZN(n12014) );
  OAI211_X1 U23902 ( .C1(n13161), .C2(n13174), .A(n12018), .B(n12017), .ZN(
        n12019) );
  OAI21_X1 U23903 ( .B1(n12417), .B2(n12019), .A(n13178), .ZN(n12020) );
  INV_X1 U23904 ( .A(n14023), .ZN(n12021) );
  NOR2_X1 U23905 ( .A1(n12021), .A2(n13729), .ZN(n14025) );
  AND2_X1 U23906 ( .A1(n14030), .A2(n14022), .ZN(n14021) );
  NAND2_X1 U23907 ( .A1(n13306), .A2(n469), .ZN(n13304) );
  INV_X1 U23908 ( .A(n13304), .ZN(n12022) );
  AOI22_X1 U23909 ( .A1(n14033), .A2(n14025), .B1(n14021), .B2(n12022), .ZN(
        n12026) );
  NOR2_X1 U23910 ( .A1(n13737), .A2(n469), .ZN(n12412) );
  INV_X1 U23911 ( .A(n14030), .ZN(n13308) );
  OAI21_X1 U23912 ( .B1(n12412), .B2(n13308), .A(n13729), .ZN(n12025) );
  OAI21_X1 U23913 ( .B1(n13308), .B2(n12023), .A(n6726), .ZN(n12024) );
  XNOR2_X1 U23914 ( .A(n12027), .B(n16661), .ZN(n12194) );
  NAND2_X1 U23916 ( .A1(n14870), .A2(n13874), .ZN(n12032) );
  NOR2_X1 U23917 ( .A1(n13262), .A2(n12032), .ZN(n12033) );
  NOR3_X1 U23918 ( .A1(n14871), .A2(n15425), .A3(n14870), .ZN(n12034) );
  AND2_X1 U23919 ( .A1(n13886), .A2(n13885), .ZN(n13252) );
  AOI21_X1 U23920 ( .B1(n12034), .B2(n13262), .A(n13252), .ZN(n12035) );
  INV_X1 U23921 ( .A(n13434), .ZN(n12038) );
  NAND4_X1 U23922 ( .A1(n12038), .A2(n12037), .A3(n13449), .A4(n12042), .ZN(
        n12040) );
  AND2_X1 U23923 ( .A1(n12040), .A2(n12039), .ZN(n14650) );
  INV_X1 U23924 ( .A(n14656), .ZN(n12041) );
  OR2_X1 U23925 ( .A1(n12042), .A2(n13449), .ZN(n14651) );
  NAND2_X1 U23926 ( .A1(n12044), .A2(n799), .ZN(n12049) );
  NAND3_X1 U23927 ( .A1(n12047), .A2(n12046), .A3(n12045), .ZN(n12048) );
  NAND3_X1 U23928 ( .A1(n12050), .A2(n12049), .A3(n12048), .ZN(n12065) );
  AOI22_X1 U23929 ( .A1(n12053), .A2(n12052), .B1(n12051), .B2(n12058), .ZN(
        n12063) );
  NAND3_X1 U23930 ( .A1(n12056), .A2(n12055), .A3(n12059), .ZN(n12061) );
  OAI211_X1 U23931 ( .C1(n12063), .C2(n12062), .A(n12061), .B(n2435), .ZN(
        n12064) );
  AOI21_X1 U23932 ( .B1(n12066), .B2(n12630), .A(n12635), .ZN(n12067) );
  NAND2_X1 U23933 ( .A1(n12631), .A2(n12630), .ZN(n12070) );
  NAND3_X1 U23934 ( .A1(n12628), .A2(n4041), .A3(n12074), .ZN(n12077) );
  INV_X1 U23935 ( .A(n12075), .ZN(n12076) );
  NAND2_X1 U23936 ( .A1(n4041), .A2(n12616), .ZN(n12642) );
  NAND2_X1 U23937 ( .A1(n12079), .A2(n12642), .ZN(n12082) );
  NAND3_X1 U23938 ( .A1(n12080), .A2(n12628), .A3(n3347), .ZN(n12081) );
  NAND2_X1 U23939 ( .A1(n12097), .A2(n51138), .ZN(n12086) );
  INV_X1 U23940 ( .A(n12085), .ZN(n12090) );
  NAND2_X1 U23942 ( .A1(n12087), .A2(n12088), .ZN(n12378) );
  NAND3_X1 U23943 ( .A1(n12370), .A2(n12098), .A3(n12088), .ZN(n12089) );
  INV_X1 U23944 ( .A(n12092), .ZN(n12096) );
  NAND3_X1 U23945 ( .A1(n12099), .A2(n12098), .A3(n12097), .ZN(n12102) );
  NAND2_X1 U23946 ( .A1(n12376), .A2(n12389), .ZN(n12100) );
  NOR2_X1 U23947 ( .A1(n14368), .A2(n14370), .ZN(n12983) );
  INV_X1 U23948 ( .A(n12105), .ZN(n12109) );
  NAND2_X1 U23949 ( .A1(n12111), .A2(n12114), .ZN(n12116) );
  INV_X1 U23950 ( .A(n12120), .ZN(n12124) );
  INV_X1 U23951 ( .A(n12121), .ZN(n12122) );
  OAI21_X1 U23952 ( .B1(n12124), .B2(n12123), .A(n12122), .ZN(n12126) );
  NAND2_X1 U23953 ( .A1(n12126), .A2(n12125), .ZN(n12127) );
  NAND3_X1 U23954 ( .A1(n12130), .A2(n438), .A3(n12129), .ZN(n12131) );
  OAI21_X1 U23955 ( .B1(n12133), .B2(n12132), .A(n12131), .ZN(n12135) );
  NAND2_X1 U23956 ( .A1(n12135), .A2(n12134), .ZN(n12150) );
  AOI21_X1 U23957 ( .B1(n12138), .B2(n12137), .A(n12136), .ZN(n12149) );
  NAND2_X1 U23958 ( .A1(n12140), .A2(n12139), .ZN(n12142) );
  OAI21_X1 U23959 ( .B1(n12143), .B2(n12142), .A(n12141), .ZN(n12148) );
  NAND3_X1 U23960 ( .A1(n12146), .A2(n438), .A3(n12144), .ZN(n12147) );
  NAND2_X1 U23961 ( .A1(n3038), .A2(n1283), .ZN(n14367) );
  NOR2_X1 U23962 ( .A1(n12151), .A2(n12173), .ZN(n12155) );
  INV_X1 U23963 ( .A(n12158), .ZN(n12154) );
  NAND4_X1 U23964 ( .A1(n12155), .A2(n12154), .A3(n12153), .A4(n12152), .ZN(
        n12165) );
  NOR2_X1 U23965 ( .A1(n12156), .A2(n12175), .ZN(n12157) );
  OAI211_X1 U23967 ( .C1(n12161), .C2(n12160), .A(n12159), .B(n12169), .ZN(
        n12162) );
  NAND2_X1 U23969 ( .A1(n12165), .A2(n12164), .ZN(n12185) );
  NAND3_X1 U23970 ( .A1(n12168), .A2(n12167), .A3(n12166), .ZN(n12184) );
  NAND3_X1 U23971 ( .A1(n12170), .A2(n12173), .A3(n12169), .ZN(n12172) );
  OAI211_X1 U23972 ( .C1(n12174), .C2(n12173), .A(n12172), .B(n12171), .ZN(
        n12183) );
  NAND2_X1 U23973 ( .A1(n12176), .A2(n12175), .ZN(n12181) );
  NAND2_X1 U23974 ( .A1(n12178), .A2(n12177), .ZN(n12180) );
  MUX2_X1 U23975 ( .A(n12181), .B(n12180), .S(n12179), .Z(n12182) );
  NOR2_X1 U23977 ( .A1(n14367), .A2(n14542), .ZN(n14362) );
  AND2_X1 U23978 ( .A1(n14542), .A2(n14552), .ZN(n14548) );
  OR2_X1 U23979 ( .A1(n14550), .A2(n14533), .ZN(n14363) );
  INV_X1 U23980 ( .A(n14363), .ZN(n13353) );
  NOR2_X1 U23981 ( .A1(n14544), .A2(n14542), .ZN(n12430) );
  AOI21_X1 U23982 ( .B1(n14548), .B2(n13353), .A(n12430), .ZN(n12188) );
  NAND2_X1 U23983 ( .A1(n13362), .A2(n14370), .ZN(n12981) );
  NAND2_X1 U23986 ( .A1(n16039), .A2(n14515), .ZN(n12805) );
  NAND2_X1 U23987 ( .A1(n12810), .A2(n12805), .ZN(n12192) );
  AND2_X1 U23988 ( .A1(n13377), .A2(n16036), .ZN(n14522) );
  INV_X1 U23989 ( .A(n14522), .ZN(n12189) );
  OAI211_X1 U23991 ( .C1(n16044), .C2(n12189), .A(n13370), .B(n12811), .ZN(
        n12191) );
  OR2_X1 U23992 ( .A1(n51019), .A2(n11723), .ZN(n14529) );
  AND2_X1 U23993 ( .A1(n51019), .A2(n16036), .ZN(n13037) );
  NAND2_X1 U23994 ( .A1(n14515), .A2(n13377), .ZN(n14525) );
  INV_X1 U23995 ( .A(n14525), .ZN(n13380) );
  OAI21_X1 U23996 ( .B1(n6799), .B2(n13037), .A(n13380), .ZN(n12190) );
  XNOR2_X1 U23997 ( .A(n16782), .B(n16658), .ZN(n15628) );
  INV_X1 U23998 ( .A(n15628), .ZN(n12193) );
  XNOR2_X1 U23999 ( .A(n12194), .B(n12193), .ZN(n14213) );
  XNOR2_X1 U24000 ( .A(n14213), .B(n12195), .ZN(n17479) );
  NAND2_X1 U24001 ( .A1(n17569), .A2(n17479), .ZN(n19399) );
  INV_X1 U24002 ( .A(n13015), .ZN(n14278) );
  AOI22_X1 U24003 ( .A1(n14278), .A2(n13587), .B1(n12197), .B2(n12196), .ZN(
        n12210) );
  AOI21_X1 U24004 ( .B1(n13588), .B2(n14285), .A(n12199), .ZN(n12201) );
  AOI21_X1 U24006 ( .B1(n12201), .B2(n13015), .A(n12200), .ZN(n12209) );
  OAI21_X1 U24007 ( .B1(n13588), .B2(n14285), .A(n12202), .ZN(n12203) );
  NAND3_X1 U24008 ( .A1(n12203), .A2(n14280), .A3(n14277), .ZN(n12208) );
  OAI22_X1 U24009 ( .A1(n14285), .A2(n14297), .B1(n784), .B2(n13583), .ZN(
        n12206) );
  OR2_X1 U24010 ( .A1(n14280), .A2(n12204), .ZN(n13012) );
  INV_X1 U24011 ( .A(n13012), .ZN(n13584) );
  NAND2_X1 U24012 ( .A1(n12206), .A2(n13584), .ZN(n12207) );
  NAND2_X1 U24013 ( .A1(n12211), .A2(n51136), .ZN(n13145) );
  OAI211_X1 U24014 ( .C1(n12903), .C2(n14184), .A(n12212), .B(n12907), .ZN(
        n12221) );
  NOR3_X1 U24015 ( .A1(n12907), .A2(n13135), .A3(n14186), .ZN(n12215) );
  AND2_X1 U24016 ( .A1(n13148), .A2(n13136), .ZN(n12214) );
  AOI22_X1 U24017 ( .A1(n12215), .A2(n12214), .B1(n12213), .B2(n12907), .ZN(
        n12220) );
  OAI211_X1 U24018 ( .C1(n13139), .C2(n51136), .A(n14179), .B(n12217), .ZN(
        n12218) );
  XNOR2_X1 U24020 ( .A(n17793), .B(n18447), .ZN(n15149) );
  AND2_X1 U24021 ( .A1(n14346), .A2(n14331), .ZN(n14340) );
  NOR2_X1 U24022 ( .A1(n13410), .A2(n14341), .ZN(n13421) );
  NAND3_X1 U24023 ( .A1(n14340), .A2(n14339), .A3(n13421), .ZN(n12226) );
  NOR2_X1 U24024 ( .A1(n12227), .A2(n13417), .ZN(n12222) );
  NAND2_X1 U24025 ( .A1(n13425), .A2(n12222), .ZN(n14351) );
  OAI211_X1 U24026 ( .C1(n12224), .C2(n13424), .A(n13425), .B(n6073), .ZN(
        n12225) );
  INV_X1 U24027 ( .A(n12227), .ZN(n14343) );
  NAND2_X1 U24028 ( .A1(n14343), .A2(n14344), .ZN(n12230) );
  INV_X1 U24029 ( .A(n12228), .ZN(n13404) );
  NAND3_X1 U24030 ( .A1(n13005), .A2(n13404), .A3(n12229), .ZN(n13814) );
  AND2_X1 U24031 ( .A1(n13410), .A2(n14341), .ZN(n13422) );
  NAND3_X1 U24032 ( .A1(n13425), .A2(n14331), .A3(n13422), .ZN(n13815) );
  NAND4_X1 U24033 ( .A1(n13816), .A2(n12230), .A3(n13814), .A4(n13815), .ZN(
        n15913) );
  XNOR2_X1 U24034 ( .A(n15149), .B(n15913), .ZN(n12402) );
  OR2_X1 U24035 ( .A1(n14155), .A2(n13761), .ZN(n13765) );
  INV_X1 U24036 ( .A(n13765), .ZN(n12232) );
  INV_X1 U24037 ( .A(n12231), .ZN(n12235) );
  NAND3_X1 U24038 ( .A1(n13763), .A2(n13117), .A3(n13122), .ZN(n12233) );
  NOR2_X1 U24039 ( .A1(n14149), .A2(n13761), .ZN(n12234) );
  NOR3_X1 U24040 ( .A1(n12234), .A2(n14155), .A3(n14160), .ZN(n12236) );
  NOR2_X1 U24041 ( .A1(n14155), .A2(n14966), .ZN(n13113) );
  OAI21_X1 U24042 ( .B1(n12237), .B2(n13113), .A(n13759), .ZN(n12240) );
  OAI21_X1 U24043 ( .B1(n13117), .B2(n13761), .A(n12238), .ZN(n12239) );
  NAND2_X1 U24044 ( .A1(n12243), .A2(n12242), .ZN(n12244) );
  NAND2_X1 U24045 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  NAND2_X1 U24046 ( .A1(n12249), .A2(n12248), .ZN(n12275) );
  AOI22_X1 U24047 ( .A1(n12253), .A2(n12252), .B1(n12251), .B2(n12250), .ZN(
        n12274) );
  INV_X1 U24048 ( .A(n12257), .ZN(n12259) );
  NAND3_X1 U24049 ( .A1(n12260), .A2(n12259), .A3(n12258), .ZN(n12261) );
  OAI21_X1 U24052 ( .B1(n12271), .B2(n12270), .A(n12269), .ZN(n12272) );
  NAND2_X1 U24053 ( .A1(n12278), .A2(n12277), .ZN(n12279) );
  NAND4_X1 U24054 ( .A1(n12281), .A2(n12285), .A3(n12280), .A4(n12279), .ZN(
        n12289) );
  OAI21_X1 U24055 ( .B1(n12283), .B2(n12285), .A(n12282), .ZN(n12288) );
  OAI211_X1 U24056 ( .C1(n12286), .C2(n12285), .A(n12284), .B(n12283), .ZN(
        n12287) );
  AND3_X1 U24057 ( .A1(n12289), .A2(n12288), .A3(n12287), .ZN(n12298) );
  NAND3_X1 U24058 ( .A1(n12292), .A2(n12291), .A3(n12290), .ZN(n12296) );
  MUX2_X1 U24059 ( .A(n12296), .B(n12295), .S(n12294), .Z(n12297) );
  OAI211_X1 U24060 ( .C1(n12302), .C2(n12301), .A(n12300), .B(n12299), .ZN(
        n12306) );
  NAND2_X1 U24061 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  OAI21_X1 U24062 ( .B1(n12315), .B2(n12313), .A(n12309), .ZN(n12311) );
  NAND2_X1 U24063 ( .A1(n12311), .A2(n12310), .ZN(n12319) );
  NOR2_X1 U24064 ( .A1(n12313), .A2(n12312), .ZN(n12316) );
  OAI22_X1 U24065 ( .A1(n9758), .A2(n12316), .B1(n12315), .B2(n12314), .ZN(
        n12318) );
  MUX2_X1 U24066 ( .A(n12319), .B(n12318), .S(n12317), .Z(n12320) );
  NAND3_X1 U24067 ( .A1(n12333), .A2(n52199), .A3(n12323), .ZN(n12327) );
  NAND3_X1 U24068 ( .A1(n12327), .A2(n10279), .A3(n12326), .ZN(n12329) );
  NAND3_X1 U24069 ( .A1(n12329), .A2(n12340), .A3(n12328), .ZN(n12330) );
  NAND2_X1 U24071 ( .A1(n12335), .A2(n12334), .ZN(n12348) );
  OAI22_X1 U24072 ( .A1(n10288), .A2(n12342), .B1(n12341), .B2(n12340), .ZN(
        n12345) );
  NAND2_X1 U24073 ( .A1(n12345), .A2(n12344), .ZN(n12346) );
  NAND2_X1 U24074 ( .A1(n14719), .A2(n14716), .ZN(n13743) );
  AOI21_X1 U24075 ( .B1(n805), .B2(n12356), .A(n9782), .ZN(n12361) );
  NAND2_X1 U24076 ( .A1(n12358), .A2(n12357), .ZN(n12360) );
  NAND4_X1 U24077 ( .A1(n12362), .A2(n12361), .A3(n12360), .A4(n12359), .ZN(
        n12366) );
  AOI21_X1 U24078 ( .B1(n14717), .B2(n14709), .A(n14711), .ZN(n12393) );
  NAND2_X1 U24079 ( .A1(n12370), .A2(n12379), .ZN(n12390) );
  OAI21_X1 U24080 ( .B1(n12372), .B2(n12371), .A(n12390), .ZN(n12374) );
  AOI21_X1 U24081 ( .B1(n12376), .B2(n12375), .A(n12383), .ZN(n12377) );
  OAI21_X1 U24082 ( .B1(n12378), .B2(n12380), .A(n12377), .ZN(n12388) );
  INV_X1 U24083 ( .A(n12379), .ZN(n12382) );
  OAI211_X1 U24084 ( .C1(n12382), .C2(n12381), .A(n9369), .B(n12380), .ZN(
        n12387) );
  NAND3_X1 U24085 ( .A1(n12385), .A2(n12384), .A3(n12383), .ZN(n12386) );
  MUX2_X1 U24086 ( .A(n12391), .B(n12390), .S(n12389), .Z(n12392) );
  NAND3_X1 U24087 ( .A1(n12394), .A2(n14704), .A3(n14197), .ZN(n12399) );
  NOR2_X1 U24088 ( .A1(n14713), .A2(n14720), .ZN(n14205) );
  INV_X1 U24089 ( .A(n14711), .ZN(n14703) );
  NAND2_X1 U24090 ( .A1(n14205), .A2(n14703), .ZN(n13334) );
  NOR2_X1 U24091 ( .A1(n51669), .A2(n14716), .ZN(n13331) );
  NOR2_X1 U24092 ( .A1(n14719), .A2(n14716), .ZN(n12395) );
  AOI22_X1 U24093 ( .A1(n13742), .A2(n13331), .B1(n13337), .B2(n12395), .ZN(
        n12397) );
  NAND2_X1 U24094 ( .A1(n14088), .A2(n14704), .ZN(n14084) );
  NOR2_X1 U24095 ( .A1(n14711), .A2(n51670), .ZN(n14085) );
  OAI211_X1 U24096 ( .C1(n12395), .C2(n14088), .A(n14084), .B(n14085), .ZN(
        n12396) );
  AOI21_X2 U24097 ( .B1(n12400), .B2(n12399), .A(n12398), .ZN(n16913) );
  NAND2_X1 U24099 ( .A1(n12403), .A2(n469), .ZN(n12405) );
  NOR2_X1 U24100 ( .A1(n12405), .A2(n12404), .ZN(n13298) );
  NOR2_X1 U24101 ( .A1(n13729), .A2(n469), .ZN(n13734) );
  NAND2_X1 U24102 ( .A1(n13734), .A2(n14030), .ZN(n12409) );
  NAND3_X1 U24103 ( .A1(n14019), .A2(n13306), .A3(n14033), .ZN(n12408) );
  NAND3_X1 U24104 ( .A1(n13729), .A2(n14022), .A3(n13291), .ZN(n13288) );
  NOR2_X1 U24105 ( .A1(n14030), .A2(n13729), .ZN(n13300) );
  NAND2_X1 U24106 ( .A1(n12410), .A2(n469), .ZN(n12411) );
  OAI211_X1 U24107 ( .C1(n6726), .C2(n13299), .A(n13300), .B(n12411), .ZN(
        n12414) );
  NAND2_X1 U24108 ( .A1(n12412), .A2(n14022), .ZN(n12413) );
  MUX2_X1 U24109 ( .A(n13779), .B(n13160), .S(n13774), .Z(n12415) );
  OAI21_X1 U24110 ( .B1(n12416), .B2(n13173), .A(n12415), .ZN(n12422) );
  NOR2_X1 U24111 ( .A1(n13779), .A2(n13173), .ZN(n13171) );
  NAND3_X1 U24112 ( .A1(n12417), .A2(n13186), .A3(n13776), .ZN(n12418) );
  NAND3_X1 U24113 ( .A1(n13178), .A2(n12419), .A3(n13174), .ZN(n12420) );
  NAND2_X1 U24114 ( .A1(n13174), .A2(n13173), .ZN(n13783) );
  AND4_X1 U24115 ( .A1(n12420), .A2(n13166), .A3(n12424), .A4(n13783), .ZN(
        n12421) );
  INV_X1 U24116 ( .A(n14545), .ZN(n13354) );
  NAND3_X1 U24117 ( .A1(n13361), .A2(n14550), .A3(n14542), .ZN(n12428) );
  NAND2_X1 U24118 ( .A1(n14540), .A2(n14550), .ZN(n12427) );
  NAND4_X1 U24119 ( .A1(n14536), .A2(n14534), .A3(n14544), .A4(n14552), .ZN(
        n12426) );
  NOR2_X1 U24120 ( .A1(n13354), .A2(n14552), .ZN(n14537) );
  NAND4_X1 U24121 ( .A1(n14537), .A2(n14536), .A3(n14544), .A4(n14550), .ZN(
        n12425) );
  OAI21_X1 U24122 ( .B1(n13354), .B2(n14550), .A(n14535), .ZN(n12429) );
  NAND2_X1 U24123 ( .A1(n14534), .A2(n14542), .ZN(n14541) );
  INV_X1 U24124 ( .A(n14541), .ZN(n12431) );
  NOR2_X1 U24125 ( .A1(n14370), .A2(n14553), .ZN(n13347) );
  AND2_X1 U24126 ( .A1(n306), .A2(n12698), .ZN(n12447) );
  INV_X1 U24127 ( .A(n12441), .ZN(n12714) );
  NAND2_X1 U24129 ( .A1(n12445), .A2(n12444), .ZN(n12446) );
  NAND2_X1 U24130 ( .A1(n12676), .A2(n50997), .ZN(n12452) );
  OAI211_X1 U24131 ( .C1(n12454), .C2(n592), .A(n12452), .B(n12451), .ZN(
        n12457) );
  INV_X1 U24132 ( .A(n12455), .ZN(n12456) );
  AND2_X1 U24133 ( .A1(n12456), .A2(n12457), .ZN(n12468) );
  NOR2_X1 U24134 ( .A1(n12458), .A2(n7354), .ZN(n12460) );
  OAI21_X1 U24135 ( .B1(n12461), .B2(n12460), .A(n12459), .ZN(n12467) );
  INV_X1 U24136 ( .A(n12673), .ZN(n12463) );
  OAI22_X1 U24137 ( .A1(n12464), .A2(n12463), .B1(n12462), .B2(n11500), .ZN(
        n12465) );
  NAND2_X1 U24138 ( .A1(n12465), .A2(n7354), .ZN(n12466) );
  NOR2_X1 U24139 ( .A1(n14962), .A2(n14957), .ZN(n15274) );
  NAND2_X1 U24140 ( .A1(n12471), .A2(n12470), .ZN(n12482) );
  AND2_X1 U24141 ( .A1(n12472), .A2(n12482), .ZN(n12477) );
  OAI211_X1 U24142 ( .C1(n12474), .C2(n12483), .A(n12473), .B(n800), .ZN(
        n12476) );
  MUX2_X1 U24143 ( .A(n12477), .B(n12476), .S(n12475), .Z(n12494) );
  NAND4_X1 U24144 ( .A1(n12482), .A2(n5251), .A3(n12480), .A4(n12479), .ZN(
        n12492) );
  INV_X1 U24145 ( .A(n12483), .ZN(n12485) );
  NAND3_X1 U24146 ( .A1(n12485), .A2(n12484), .A3(n8099), .ZN(n12490) );
  OAI211_X1 U24147 ( .C1(n2116), .C2(n12488), .A(n12487), .B(n12486), .ZN(
        n12489) );
  AND4_X1 U24148 ( .A1(n12490), .A2(n12492), .A3(n12491), .A4(n12489), .ZN(
        n12493) );
  NAND2_X2 U24149 ( .A1(n12494), .A2(n12493), .ZN(n14950) );
  NOR2_X1 U24150 ( .A1(n14950), .A2(n51500), .ZN(n12531) );
  NAND2_X1 U24151 ( .A1(n12506), .A2(n12518), .ZN(n12497) );
  NAND3_X1 U24152 ( .A1(n12501), .A2(n12500), .A3(n12504), .ZN(n12510) );
  NAND4_X1 U24153 ( .A1(n12507), .A2(n12506), .A3(n51653), .A4(n12504), .ZN(
        n12508) );
  AND3_X1 U24154 ( .A1(n12509), .A2(n12510), .A3(n12508), .ZN(n12530) );
  INV_X1 U24155 ( .A(n12511), .ZN(n12513) );
  NAND4_X1 U24156 ( .A1(n12519), .A2(n8024), .A3(n12518), .A4(n12517), .ZN(
        n12529) );
  INV_X1 U24157 ( .A(n12523), .ZN(n12520) );
  OAI21_X1 U24158 ( .B1(n12522), .B2(n12521), .A(n12520), .ZN(n12527) );
  OAI21_X1 U24159 ( .B1(n12525), .B2(n12524), .A(n12523), .ZN(n12526) );
  NAND2_X1 U24160 ( .A1(n12527), .A2(n12526), .ZN(n12528) );
  OAI21_X1 U24161 ( .B1(n15274), .B2(n12531), .A(n15279), .ZN(n12582) );
  OAI21_X1 U24162 ( .B1(n442), .B2(n12537), .A(n12536), .ZN(n12539) );
  AOI22_X1 U24163 ( .A1(n12540), .A2(n12539), .B1(n12545), .B2(n12538), .ZN(
        n12552) );
  INV_X1 U24164 ( .A(n12547), .ZN(n12548) );
  NAND3_X1 U24165 ( .A1(n12550), .A2(n12549), .A3(n12548), .ZN(n12551) );
  NOR2_X1 U24166 ( .A1(n15278), .A2(n14957), .ZN(n14052) );
  INV_X1 U24167 ( .A(n12553), .ZN(n12554) );
  OAI21_X1 U24168 ( .B1(n12556), .B2(n12555), .A(n12554), .ZN(n12560) );
  AOI22_X1 U24169 ( .A1(n12560), .A2(n12559), .B1(n12558), .B2(n12557), .ZN(
        n12564) );
  INV_X1 U24170 ( .A(n12561), .ZN(n12562) );
  INV_X1 U24171 ( .A(n12565), .ZN(n12567) );
  NAND2_X1 U24172 ( .A1(n12567), .A2(n12566), .ZN(n12580) );
  INV_X1 U24174 ( .A(n12572), .ZN(n12576) );
  NOR2_X1 U24175 ( .A1(n12574), .A2(n12573), .ZN(n12575) );
  AOI22_X1 U24176 ( .A1(n12578), .A2(n12577), .B1(n12576), .B2(n12575), .ZN(
        n12579) );
  AOI21_X1 U24177 ( .B1(n14052), .B2(n14938), .A(n2151), .ZN(n12581) );
  INV_X1 U24178 ( .A(n14950), .ZN(n14959) );
  NAND2_X1 U24179 ( .A1(n14959), .A2(n15278), .ZN(n14955) );
  NAND2_X1 U24180 ( .A1(n51500), .A2(n15279), .ZN(n14946) );
  NOR2_X1 U24181 ( .A1(n14946), .A2(n14962), .ZN(n12583) );
  AOI22_X1 U24182 ( .A1(n12583), .A2(n14949), .B1(n15273), .B2(n14956), .ZN(
        n12587) );
  OAI211_X1 U24184 ( .C1(n14935), .C2(n15278), .A(n51724), .B(n51500), .ZN(
        n12586) );
  INV_X1 U24185 ( .A(n14962), .ZN(n14692) );
  NOR2_X1 U24186 ( .A1(n14692), .A2(n14950), .ZN(n12584) );
  OAI211_X1 U24187 ( .C1(n14059), .C2(n12584), .A(n2151), .B(n14938), .ZN(
        n12585) );
  XNOR2_X1 U24188 ( .A(n17923), .B(n16011), .ZN(n12748) );
  NOR2_X1 U24189 ( .A1(n12589), .A2(n12604), .ZN(n12593) );
  NOR2_X1 U24190 ( .A1(n12590), .A2(n12605), .ZN(n12591) );
  AND2_X1 U24191 ( .A1(n12596), .A2(n52140), .ZN(n12599) );
  OAI22_X1 U24192 ( .A1(n12602), .A2(n12601), .B1(n12600), .B2(n3377), .ZN(
        n12603) );
  OAI21_X1 U24193 ( .B1(n12611), .B2(n1307), .A(n12609), .ZN(n12614) );
  MUX2_X1 U24194 ( .A(n12614), .B(n12613), .S(n51140), .Z(n12615) );
  NOR2_X1 U24195 ( .A1(n12632), .A2(n12618), .ZN(n12622) );
  AOI22_X1 U24196 ( .A1(n12624), .A2(n12623), .B1(n12622), .B2(n12621), .ZN(
        n12646) );
  INV_X1 U24197 ( .A(n12625), .ZN(n12636) );
  NOR2_X1 U24198 ( .A1(n12627), .A2(n51433), .ZN(n12629) );
  OAI21_X1 U24199 ( .B1(n12636), .B2(n12629), .A(n12628), .ZN(n12645) );
  OAI211_X1 U24200 ( .C1(n12631), .C2(n12630), .A(n3347), .B(n9208), .ZN(
        n12633) );
  NOR2_X1 U24201 ( .A1(n12633), .A2(n12632), .ZN(n12634) );
  OAI21_X1 U24202 ( .B1(n12636), .B2(n12635), .A(n12634), .ZN(n12644) );
  INV_X1 U24203 ( .A(n12637), .ZN(n12639) );
  AND2_X1 U24205 ( .A1(n12641), .A2(n12642), .ZN(n12643) );
  INV_X1 U24206 ( .A(n12740), .ZN(n15067) );
  NAND3_X1 U24207 ( .A1(n2227), .A2(n12649), .A3(n12648), .ZN(n12650) );
  AND2_X1 U24208 ( .A1(n12652), .A2(n12650), .ZN(n12655) );
  NOR2_X1 U24209 ( .A1(n12652), .A2(n2227), .ZN(n12653) );
  OAI21_X1 U24210 ( .B1(n12658), .B2(n12659), .A(n12657), .ZN(n12665) );
  INV_X1 U24211 ( .A(n12658), .ZN(n12662) );
  NAND4_X1 U24212 ( .A1(n12662), .A2(n12661), .A3(n12660), .A4(n12659), .ZN(
        n12664) );
  MUX2_X1 U24213 ( .A(n12665), .B(n12664), .S(n12663), .Z(n12666) );
  NAND2_X1 U24214 ( .A1(n12671), .A2(n12667), .ZN(n12668) );
  AOI21_X1 U24216 ( .B1(n11500), .B2(n12676), .A(n12675), .ZN(n12677) );
  NAND2_X1 U24217 ( .A1(n12678), .A2(n12677), .ZN(n12684) );
  INV_X1 U24218 ( .A(n12679), .ZN(n12681) );
  NAND2_X1 U24219 ( .A1(n12681), .A2(n12680), .ZN(n12682) );
  NAND3_X1 U24220 ( .A1(n12684), .A2(n12683), .A3(n12682), .ZN(n12685) );
  NAND2_X1 U24222 ( .A1(n15767), .A2(n15063), .ZN(n12738) );
  NAND3_X1 U24223 ( .A1(n12692), .A2(n12696), .A3(n12709), .ZN(n12693) );
  NAND2_X1 U24224 ( .A1(n12696), .A2(n12695), .ZN(n12697) );
  INV_X1 U24225 ( .A(n12703), .ZN(n12706) );
  NAND3_X1 U24226 ( .A1(n12706), .A2(n12705), .A3(n12704), .ZN(n12707) );
  NOR2_X1 U24227 ( .A1(n12711), .A2(n12710), .ZN(n12716) );
  NOR2_X1 U24228 ( .A1(n12713), .A2(n12712), .ZN(n12715) );
  MUX2_X1 U24229 ( .A(n12716), .B(n12715), .S(n12714), .Z(n12717) );
  AOI22_X1 U24230 ( .A1(n12721), .A2(n12720), .B1(n12719), .B2(n12718), .ZN(
        n12736) );
  OAI22_X1 U24231 ( .A1(n12724), .A2(n12723), .B1(n8882), .B2(n12722), .ZN(
        n12726) );
  NAND2_X1 U24232 ( .A1(n12726), .A2(n6912), .ZN(n12735) );
  AND3_X1 U24233 ( .A1(n12732), .A2(n12731), .A3(n12730), .ZN(n12734) );
  NAND2_X1 U24234 ( .A1(n15068), .A2(n14914), .ZN(n12737) );
  OAI211_X1 U24235 ( .C1(n12738), .C2(n15077), .A(n13789), .B(n12737), .ZN(
        n12739) );
  INV_X1 U24236 ( .A(n12739), .ZN(n12747) );
  INV_X1 U24237 ( .A(n14911), .ZN(n15066) );
  NAND3_X1 U24238 ( .A1(n15767), .A2(n15066), .A3(n15073), .ZN(n12741) );
  AND2_X1 U24239 ( .A1(n15060), .A2(n14911), .ZN(n15769) );
  NAND2_X1 U24240 ( .A1(n15769), .A2(n15068), .ZN(n14930) );
  NAND3_X1 U24241 ( .A1(n12741), .A2(n14929), .A3(n14930), .ZN(n12743) );
  NAND3_X1 U24242 ( .A1(n15300), .A2(n14911), .A3(n15770), .ZN(n12742) );
  NAND2_X1 U24243 ( .A1(n12743), .A2(n15299), .ZN(n12746) );
  AND2_X1 U24244 ( .A1(n2189), .A2(n15770), .ZN(n15069) );
  NAND2_X1 U24245 ( .A1(n15069), .A2(n14911), .ZN(n15298) );
  AND2_X1 U24246 ( .A1(n15303), .A2(n15298), .ZN(n12745) );
  XNOR2_X1 U24247 ( .A(n18438), .B(n12748), .ZN(n12749) );
  XNOR2_X1 U24248 ( .A(n17798), .B(n12749), .ZN(n17268) );
  AOI21_X1 U24249 ( .B1(n14642), .B2(n14633), .A(n12755), .ZN(n12751) );
  NOR2_X1 U24250 ( .A1(n12751), .A2(n14634), .ZN(n12752) );
  NOR2_X1 U24251 ( .A1(n14639), .A2(n12752), .ZN(n12762) );
  NOR2_X1 U24252 ( .A1(n13669), .A2(n3254), .ZN(n13650) );
  NAND2_X1 U24253 ( .A1(n13653), .A2(n13669), .ZN(n12759) );
  NAND2_X1 U24254 ( .A1(n14636), .A2(n3254), .ZN(n13654) );
  NAND4_X1 U24255 ( .A1(n14635), .A2(n13658), .A3(n3254), .A4(n13659), .ZN(
        n12760) );
  NOR2_X1 U24256 ( .A1(n13506), .A2(n13514), .ZN(n12763) );
  OAI21_X1 U24257 ( .B1(n13512), .B2(n12763), .A(n13527), .ZN(n12764) );
  OAI211_X1 U24258 ( .C1(n12765), .C2(n12764), .A(n13500), .B(n12766), .ZN(
        n12772) );
  NAND3_X1 U24259 ( .A1(n12768), .A2(n13501), .A3(n13526), .ZN(n12771) );
  XNOR2_X1 U24261 ( .A(n16919), .B(n16923), .ZN(n12804) );
  OR2_X1 U24262 ( .A1(n13797), .A2(n13804), .ZN(n13486) );
  OAI211_X1 U24263 ( .C1(n15034), .C2(n15033), .A(n13805), .B(n13801), .ZN(
        n12774) );
  NOR2_X1 U24264 ( .A1(n12773), .A2(n15034), .ZN(n13492) );
  OAI22_X1 U24265 ( .A1(n12775), .A2(n12774), .B1(n13492), .B2(n13801), .ZN(
        n12784) );
  AND2_X1 U24266 ( .A1(n15034), .A2(n13800), .ZN(n15049) );
  NOR3_X1 U24267 ( .A1(n15044), .A2(n13797), .A3(n13801), .ZN(n12778) );
  NOR2_X1 U24268 ( .A1(n15046), .A2(n13801), .ZN(n12776) );
  AOI22_X1 U24269 ( .A1(n15049), .A2(n12778), .B1(n12777), .B2(n12776), .ZN(
        n12783) );
  OAI21_X1 U24270 ( .B1(n15034), .B2(n13483), .A(n15035), .ZN(n12779) );
  AND2_X1 U24271 ( .A1(n13801), .A2(n13804), .ZN(n13795) );
  OAI21_X1 U24272 ( .B1(n13481), .B2(n12779), .A(n13795), .ZN(n12782) );
  NAND2_X1 U24273 ( .A1(n15049), .A2(n12780), .ZN(n12781) );
  NOR2_X1 U24274 ( .A1(n483), .A2(n12787), .ZN(n13990) );
  AND2_X1 U24275 ( .A1(n12787), .A2(n12788), .ZN(n13429) );
  NAND2_X1 U24276 ( .A1(n13429), .A2(n483), .ZN(n12789) );
  NAND2_X1 U24277 ( .A1(n4949), .A2(n483), .ZN(n13430) );
  AND2_X1 U24278 ( .A1(n12799), .A2(n13430), .ZN(n13447) );
  AND2_X1 U24279 ( .A1(n12791), .A2(n12790), .ZN(n13446) );
  NAND2_X1 U24280 ( .A1(n13447), .A2(n13446), .ZN(n12802) );
  INV_X1 U24281 ( .A(n12792), .ZN(n13448) );
  NOR2_X1 U24282 ( .A1(n12793), .A2(n13448), .ZN(n12889) );
  NAND2_X1 U24283 ( .A1(n12889), .A2(n12794), .ZN(n12801) );
  AOI21_X1 U24284 ( .B1(n13439), .B2(n12894), .A(n786), .ZN(n12798) );
  NAND2_X1 U24285 ( .A1(n12794), .A2(n13432), .ZN(n13991) );
  INV_X1 U24286 ( .A(n13991), .ZN(n12796) );
  NAND2_X1 U24287 ( .A1(n13449), .A2(n12893), .ZN(n12795) );
  NAND2_X1 U24288 ( .A1(n12796), .A2(n12795), .ZN(n12797) );
  OAI211_X1 U24289 ( .C1(n13450), .C2(n12799), .A(n12798), .B(n12797), .ZN(
        n12800) );
  XNOR2_X1 U24290 ( .A(n16023), .B(n16016), .ZN(n12803) );
  XNOR2_X1 U24291 ( .A(n12804), .B(n12803), .ZN(n12830) );
  OR2_X1 U24292 ( .A1(n11723), .A2(n51714), .ZN(n13039) );
  OR2_X1 U24293 ( .A1(n51019), .A2(n51714), .ZN(n13386) );
  OAI22_X1 U24294 ( .A1(n13372), .A2(n13039), .B1(n14516), .B2(n13386), .ZN(
        n12807) );
  NOR2_X1 U24296 ( .A1(n12807), .A2(n12806), .ZN(n12817) );
  OAI21_X1 U24297 ( .B1(n16039), .B2(n13384), .A(n51713), .ZN(n12808) );
  NOR2_X1 U24298 ( .A1(n12809), .A2(n12808), .ZN(n12812) );
  AOI22_X1 U24299 ( .A1(n12812), .A2(n12811), .B1(n12810), .B2(n51713), .ZN(
        n12816) );
  NAND2_X1 U24300 ( .A1(n12813), .A2(n16036), .ZN(n13391) );
  OAI21_X1 U24301 ( .B1(n14519), .B2(n51019), .A(n16049), .ZN(n12814) );
  NAND2_X1 U24302 ( .A1(n13035), .A2(n12814), .ZN(n12815) );
  NAND4_X2 U24303 ( .A1(n12816), .A2(n12817), .A3(n13391), .A4(n12815), .ZN(
        n18432) );
  OR2_X1 U24304 ( .A1(n12818), .A2(n12915), .ZN(n12819) );
  AND2_X1 U24305 ( .A1(n12820), .A2(n12819), .ZN(n12829) );
  MUX2_X1 U24306 ( .A(n13088), .B(n13086), .S(n13091), .Z(n12822) );
  OAI211_X1 U24307 ( .C1(n12822), .C2(n12914), .A(n13092), .B(n13081), .ZN(
        n12827) );
  AOI21_X1 U24308 ( .B1(n13103), .B2(n12823), .A(n13086), .ZN(n12825) );
  OAI211_X1 U24309 ( .C1(n13102), .C2(n13093), .A(n12825), .B(n12824), .ZN(
        n12826) );
  XNOR2_X1 U24310 ( .A(n14803), .B(n18432), .ZN(n18550) );
  XNOR2_X1 U24311 ( .A(n12830), .B(n18550), .ZN(n12878) );
  NAND2_X1 U24312 ( .A1(n13633), .A2(n14666), .ZN(n12951) );
  NOR2_X1 U24313 ( .A1(n12951), .A2(n2150), .ZN(n14617) );
  INV_X1 U24314 ( .A(n14617), .ZN(n12842) );
  AOI21_X1 U24315 ( .B1(n12948), .B2(n12831), .A(n7755), .ZN(n12833) );
  NAND3_X1 U24316 ( .A1(n14665), .A2(n12834), .A3(n14664), .ZN(n14667) );
  NAND2_X1 U24317 ( .A1(n13633), .A2(n2150), .ZN(n14670) );
  NOR2_X1 U24318 ( .A1(n14667), .A2(n14670), .ZN(n12832) );
  NOR2_X1 U24319 ( .A1(n12833), .A2(n12832), .ZN(n12839) );
  NOR2_X1 U24320 ( .A1(n12834), .A2(n2150), .ZN(n12836) );
  OAI21_X1 U24321 ( .B1(n12952), .B2(n12836), .A(n12835), .ZN(n12837) );
  OAI21_X1 U24323 ( .B1(n7755), .B2(n785), .A(n12948), .ZN(n14618) );
  NAND2_X1 U24324 ( .A1(n14618), .A2(n12840), .ZN(n12841) );
  OAI211_X1 U24325 ( .C1(n12842), .C2(n14664), .A(n14619), .B(n12841), .ZN(
        n16017) );
  XNOR2_X1 U24326 ( .A(n4653), .B(n4826), .ZN(n26525) );
  XNOR2_X1 U24327 ( .A(n26525), .B(n4744), .ZN(n35816) );
  XNOR2_X1 U24328 ( .A(n35816), .B(n4694), .ZN(n43620) );
  XNOR2_X1 U24329 ( .A(n4487), .B(n46552), .ZN(n15521) );
  XNOR2_X1 U24330 ( .A(n43620), .B(n15521), .ZN(n33977) );
  XNOR2_X1 U24331 ( .A(n4720), .B(n4781), .ZN(n24861) );
  XNOR2_X1 U24332 ( .A(n24861), .B(n4177), .ZN(n42025) );
  XNOR2_X1 U24333 ( .A(n33977), .B(n42025), .ZN(n12844) );
  XNOR2_X1 U24334 ( .A(n4874), .B(n4645), .ZN(n27353) );
  XNOR2_X1 U24335 ( .A(n27353), .B(n2604), .ZN(n42721) );
  XNOR2_X1 U24336 ( .A(n42721), .B(n3481), .ZN(n28116) );
  XNOR2_X1 U24337 ( .A(n49937), .B(n4287), .ZN(n28390) );
  XNOR2_X1 U24338 ( .A(n7744), .B(n4535), .ZN(n34027) );
  XNOR2_X1 U24339 ( .A(n28390), .B(n34027), .ZN(n27186) );
  XNOR2_X1 U24340 ( .A(n27186), .B(n4612), .ZN(n12843) );
  XNOR2_X1 U24341 ( .A(n28116), .B(n12843), .ZN(n34762) );
  XNOR2_X1 U24342 ( .A(n12844), .B(n34762), .ZN(n12845) );
  XNOR2_X1 U24343 ( .A(n16017), .B(n12845), .ZN(n12876) );
  OAI21_X1 U24344 ( .B1(n14100), .B2(n14453), .A(n14096), .ZN(n14094) );
  INV_X1 U24345 ( .A(n14094), .ZN(n12847) );
  INV_X1 U24346 ( .A(n14097), .ZN(n12846) );
  NAND3_X1 U24347 ( .A1(n12847), .A2(n14106), .A3(n12846), .ZN(n12849) );
  AND2_X1 U24348 ( .A1(n12849), .A2(n12848), .ZN(n12860) );
  INV_X1 U24350 ( .A(n14450), .ZN(n12851) );
  NAND2_X1 U24351 ( .A1(n14107), .A2(n14453), .ZN(n12850) );
  OAI22_X1 U24352 ( .A1(n12851), .A2(n12850), .B1(n14107), .B2(n14099), .ZN(
        n12852) );
  INV_X1 U24353 ( .A(n12852), .ZN(n12853) );
  NAND2_X1 U24354 ( .A1(n2253), .A2(n51383), .ZN(n14439) );
  NOR2_X1 U24355 ( .A1(n51383), .A2(n14454), .ZN(n12855) );
  OAI21_X1 U24356 ( .B1(n14107), .B2(n640), .A(n14455), .ZN(n12854) );
  OAI211_X1 U24357 ( .C1(n52312), .C2(n14455), .A(n12855), .B(n12854), .ZN(
        n12858) );
  NAND3_X1 U24358 ( .A1(n12856), .A2(n14450), .A3(n12977), .ZN(n12857) );
  OR3_X1 U24359 ( .A1(n14394), .A2(n12961), .A3(n14070), .ZN(n12864) );
  NAND2_X1 U24360 ( .A1(n14410), .A2(n12865), .ZN(n12964) );
  NAND2_X1 U24361 ( .A1(n12861), .A2(n14072), .ZN(n14405) );
  NAND2_X1 U24362 ( .A1(n14397), .A2(n12865), .ZN(n14419) );
  OR2_X1 U24363 ( .A1(n14412), .A2(n3512), .ZN(n12967) );
  NOR2_X1 U24364 ( .A1(n14410), .A2(n14070), .ZN(n12870) );
  OAI21_X1 U24365 ( .B1(n12870), .B2(n12865), .A(n14412), .ZN(n12866) );
  NAND4_X1 U24366 ( .A1(n14419), .A2(n12867), .A3(n12967), .A4(n12866), .ZN(
        n12874) );
  NAND3_X1 U24367 ( .A1(n12869), .A2(n12868), .A3(n12965), .ZN(n12873) );
  XNOR2_X2 U24368 ( .A(n16228), .B(n17665), .ZN(n16920) );
  XNOR2_X1 U24369 ( .A(n12876), .B(n16920), .ZN(n12877) );
  XNOR2_X1 U24370 ( .A(n12878), .B(n12877), .ZN(n12879) );
  INV_X1 U24371 ( .A(n19388), .ZN(n18014) );
  INV_X1 U24372 ( .A(n17479), .ZN(n18009) );
  OR2_X1 U24373 ( .A1(n12880), .A2(n13190), .ZN(n13938) );
  INV_X1 U24374 ( .A(n13934), .ZN(n12884) );
  AND3_X1 U24375 ( .A1(n12884), .A2(n12881), .A3(n13193), .ZN(n12883) );
  AOI21_X1 U24376 ( .B1(n13938), .B2(n12883), .A(n12882), .ZN(n12887) );
  NAND2_X1 U24377 ( .A1(n12889), .A2(n12888), .ZN(n12896) );
  NAND2_X1 U24378 ( .A1(n12900), .A2(n51136), .ZN(n12901) );
  AND3_X1 U24379 ( .A1(n12902), .A2(n13144), .A3(n12901), .ZN(n12911) );
  INV_X1 U24380 ( .A(n12903), .ZN(n12904) );
  NOR2_X1 U24381 ( .A1(n14178), .A2(n12907), .ZN(n14191) );
  NAND4_X1 U24382 ( .A1(n14189), .A2(n13142), .A3(n14178), .A4(n51136), .ZN(
        n12908) );
  NAND3_X1 U24383 ( .A1(n12913), .A2(n12912), .A3(n13089), .ZN(n13099) );
  NOR3_X1 U24384 ( .A1(n12915), .A2(n13086), .A3(n12914), .ZN(n12916) );
  XNOR2_X1 U24386 ( .A(n2126), .B(n51032), .ZN(n12960) );
  AOI21_X1 U24387 ( .B1(n14224), .B2(n16221), .A(n13968), .ZN(n12925) );
  INV_X1 U24388 ( .A(n12923), .ZN(n12924) );
  AOI22_X1 U24389 ( .A1(n13214), .A2(n12925), .B1(n12924), .B2(n13968), .ZN(
        n12930) );
  NAND2_X1 U24390 ( .A1(n13226), .A2(n14228), .ZN(n13972) );
  INV_X1 U24391 ( .A(n13958), .ZN(n12926) );
  NAND3_X1 U24392 ( .A1(n13972), .A2(n16221), .A3(n12926), .ZN(n12929) );
  NAND3_X1 U24394 ( .A1(n13971), .A2(n14228), .A3(n14234), .ZN(n13963) );
  NAND2_X1 U24395 ( .A1(n13967), .A2(n14220), .ZN(n12928) );
  MUX2_X1 U24396 ( .A(n13530), .B(n12932), .S(n13505), .Z(n12942) );
  INV_X1 U24397 ( .A(n12936), .ZN(n12937) );
  NAND3_X1 U24398 ( .A1(n12937), .A2(n13499), .A3(n13506), .ZN(n12940) );
  OAI21_X1 U24399 ( .B1(n13511), .B2(n12938), .A(n13525), .ZN(n12939) );
  XNOR2_X1 U24400 ( .A(n17906), .B(n16743), .ZN(n12958) );
  NAND3_X1 U24401 ( .A1(n12943), .A2(n2114), .A3(n13669), .ZN(n12944) );
  INV_X1 U24402 ( .A(n14636), .ZN(n13668) );
  MUX2_X1 U24403 ( .A(n12944), .B(n13668), .S(n13667), .Z(n12947) );
  OR2_X1 U24404 ( .A1(n13651), .A2(n14634), .ZN(n12946) );
  NAND3_X1 U24405 ( .A1(n14635), .A2(n14644), .A3(n13662), .ZN(n12945) );
  INV_X1 U24406 ( .A(n12948), .ZN(n13641) );
  NOR2_X1 U24407 ( .A1(n12949), .A2(n14664), .ZN(n13634) );
  NAND3_X1 U24408 ( .A1(n13622), .A2(n783), .A3(n12951), .ZN(n12955) );
  NAND2_X1 U24409 ( .A1(n13629), .A2(n12951), .ZN(n12954) );
  INV_X1 U24410 ( .A(n12952), .ZN(n12953) );
  XNOR2_X1 U24411 ( .A(n12958), .B(n2215), .ZN(n12959) );
  XNOR2_X1 U24412 ( .A(n12959), .B(n12960), .ZN(n13002) );
  NAND2_X1 U24413 ( .A1(n12964), .A2(n12963), .ZN(n14420) );
  INV_X1 U24414 ( .A(n14073), .ZN(n14418) );
  OR2_X1 U24415 ( .A1(n14420), .A2(n14418), .ZN(n12970) );
  NAND2_X1 U24416 ( .A1(n12966), .A2(n12965), .ZN(n12968) );
  OAI211_X1 U24417 ( .C1(n14415), .C2(n14394), .A(n12968), .B(n12967), .ZN(
        n12969) );
  NAND2_X1 U24418 ( .A1(n12975), .A2(n14096), .ZN(n12980) );
  OAI211_X1 U24419 ( .C1(n14095), .C2(n51383), .A(n12977), .B(n12976), .ZN(
        n12979) );
  NAND2_X1 U24420 ( .A1(n14434), .A2(n51383), .ZN(n12978) );
  XNOR2_X1 U24421 ( .A(n16980), .B(n17218), .ZN(n15650) );
  NAND3_X1 U24422 ( .A1(n12981), .A2(n14536), .A3(n14540), .ZN(n12986) );
  NAND2_X1 U24423 ( .A1(n12983), .A2(n12982), .ZN(n12985) );
  NAND2_X1 U24424 ( .A1(n13362), .A2(n13361), .ZN(n14358) );
  NAND4_X2 U24425 ( .A1(n12986), .A2(n12985), .A3(n12984), .A4(n14358), .ZN(
        n17771) );
  XNOR2_X1 U24426 ( .A(n4755), .B(n4454), .ZN(n24894) );
  XNOR2_X1 U24427 ( .A(n4659), .B(n4515), .ZN(n16739) );
  XNOR2_X1 U24428 ( .A(n24894), .B(n16739), .ZN(n21089) );
  INV_X1 U24429 ( .A(n38626), .ZN(n25062) );
  XNOR2_X1 U24430 ( .A(n21089), .B(n25062), .ZN(n25791) );
  INV_X1 U24431 ( .A(n25791), .ZN(n25576) );
  XNOR2_X1 U24432 ( .A(Key[180]), .B(Key[12]), .ZN(n24828) );
  XNOR2_X1 U24433 ( .A(n24828), .B(n4482), .ZN(n42619) );
  XNOR2_X1 U24434 ( .A(n25576), .B(n42619), .ZN(n35673) );
  XNOR2_X1 U24435 ( .A(n4325), .B(Key[150]), .ZN(n36755) );
  XNOR2_X1 U24436 ( .A(n2605), .B(n4490), .ZN(n25718) );
  XNOR2_X1 U24437 ( .A(n25040), .B(n2947), .ZN(n12987) );
  XNOR2_X1 U24438 ( .A(n25718), .B(n12987), .ZN(n35270) );
  XNOR2_X1 U24439 ( .A(n4931), .B(n842), .ZN(n44330) );
  XNOR2_X1 U24440 ( .A(n44330), .B(n26541), .ZN(n33442) );
  XNOR2_X1 U24441 ( .A(n35270), .B(n33442), .ZN(n12988) );
  XNOR2_X1 U24442 ( .A(n35673), .B(n12988), .ZN(n12989) );
  XNOR2_X1 U24443 ( .A(n17771), .B(n12989), .ZN(n12990) );
  XNOR2_X1 U24444 ( .A(n15650), .B(n12990), .ZN(n13000) );
  INV_X1 U24445 ( .A(n15157), .ZN(n12991) );
  AOI21_X1 U24446 ( .B1(n15159), .B2(n14575), .A(n12991), .ZN(n12993) );
  OAI21_X1 U24447 ( .B1(n12993), .B2(n51452), .A(n12992), .ZN(n17322) );
  NOR2_X1 U24448 ( .A1(n14612), .A2(n14010), .ZN(n12994) );
  INV_X1 U24449 ( .A(n14167), .ZN(n14606) );
  OAI211_X1 U24450 ( .C1(n14170), .C2(n14171), .A(n12995), .B(n14606), .ZN(
        n12998) );
  NAND2_X1 U24451 ( .A1(n14172), .A2(n14600), .ZN(n12997) );
  NAND3_X1 U24452 ( .A1(n14603), .A2(n14607), .A3(n14167), .ZN(n12996) );
  XNOR2_X1 U24453 ( .A(n15649), .B(n17322), .ZN(n15486) );
  XNOR2_X1 U24454 ( .A(n13000), .B(n15486), .ZN(n13001) );
  XNOR2_X1 U24455 ( .A(n13002), .B(n13001), .ZN(n13056) );
  AOI21_X1 U24456 ( .B1(n6073), .B2(n13418), .A(n14338), .ZN(n13004) );
  INV_X1 U24457 ( .A(n13812), .ZN(n13007) );
  NAND2_X1 U24458 ( .A1(n13006), .A2(n13007), .ZN(n13010) );
  OAI21_X1 U24459 ( .B1(n14342), .B2(n14341), .A(n13007), .ZN(n13009) );
  NAND3_X1 U24460 ( .A1(n13011), .A2(n14294), .A3(n13015), .ZN(n13021) );
  NOR2_X1 U24461 ( .A1(n14297), .A2(n13012), .ZN(n13016) );
  NAND2_X1 U24462 ( .A1(n14290), .A2(n13013), .ZN(n13014) );
  NOR2_X1 U24463 ( .A1(n14285), .A2(n13979), .ZN(n14279) );
  INV_X1 U24464 ( .A(n13018), .ZN(n13592) );
  NAND2_X1 U24465 ( .A1(n14279), .A2(n13592), .ZN(n13019) );
  XNOR2_X2 U24466 ( .A(n17208), .B(n18773), .ZN(n16330) );
  INV_X1 U24467 ( .A(n16330), .ZN(n16099) );
  INV_X1 U24468 ( .A(n13022), .ZN(n13025) );
  AOI21_X1 U24469 ( .B1(n14982), .B2(n8075), .A(n14983), .ZN(n13023) );
  OAI21_X1 U24470 ( .B1(n13023), .B2(n14980), .A(n15106), .ZN(n13024) );
  NAND2_X1 U24471 ( .A1(n14982), .A2(n13683), .ZN(n15109) );
  OR2_X1 U24472 ( .A1(n14982), .A2(n14984), .ZN(n15114) );
  OAI21_X1 U24473 ( .B1(n15109), .B2(n15108), .A(n15114), .ZN(n13028) );
  AOI21_X1 U24474 ( .B1(n13026), .B2(n14252), .A(n352), .ZN(n13027) );
  AND2_X1 U24475 ( .A1(n13028), .A2(n13027), .ZN(n13029) );
  NAND3_X1 U24476 ( .A1(n13697), .A2(n13709), .A3(n15138), .ZN(n13030) );
  OR2_X1 U24477 ( .A1(n15133), .A2(n15132), .ZN(n14267) );
  INV_X1 U24478 ( .A(n14995), .ZN(n13031) );
  INV_X1 U24479 ( .A(n13696), .ZN(n13715) );
  AND2_X1 U24480 ( .A1(n15132), .A2(n15126), .ZN(n14994) );
  OAI22_X1 U24481 ( .A1(n13715), .A2(n15134), .B1(n14993), .B2(n14994), .ZN(
        n13032) );
  NOR2_X1 U24482 ( .A1(n13036), .A2(n51019), .ZN(n13038) );
  AOI22_X1 U24483 ( .A1(n13038), .A2(n13039), .B1(n13037), .B2(n14519), .ZN(
        n13042) );
  INV_X1 U24484 ( .A(n13039), .ZN(n14514) );
  OAI21_X1 U24485 ( .B1(n14514), .B2(n13380), .A(n13040), .ZN(n13041) );
  NAND4_X2 U24486 ( .A1(n13044), .A2(n13043), .A3(n13042), .A4(n13041), .ZN(
        n16162) );
  AND4_X1 U24487 ( .A1(n13826), .A2(n14318), .A3(n14307), .A4(n14317), .ZN(
        n13047) );
  AOI22_X1 U24488 ( .A1(n13047), .A2(n13046), .B1(n14322), .B2(n13819), .ZN(
        n13053) );
  AND2_X1 U24489 ( .A1(n13820), .A2(n51064), .ZN(n13048) );
  OAI21_X1 U24490 ( .B1(n13048), .B2(n13605), .A(n13824), .ZN(n13052) );
  INV_X1 U24491 ( .A(n13048), .ZN(n13050) );
  NAND3_X1 U24492 ( .A1(n13050), .A2(n13049), .A3(n13827), .ZN(n13051) );
  XNOR2_X1 U24494 ( .A(n16162), .B(n51758), .ZN(n13054) );
  XNOR2_X1 U24495 ( .A(n2180), .B(n13054), .ZN(n17211) );
  XNOR2_X1 U24496 ( .A(n17211), .B(n16099), .ZN(n16972) );
  INV_X1 U24497 ( .A(n16972), .ZN(n13055) );
  NOR2_X1 U24498 ( .A1(n14137), .A2(n13061), .ZN(n14788) );
  NAND2_X1 U24499 ( .A1(n15263), .A2(n14784), .ZN(n13059) );
  OAI22_X1 U24500 ( .A1(n15263), .A2(n13060), .B1(n13059), .B2(n14796), .ZN(
        n13063) );
  NAND2_X1 U24501 ( .A1(n13061), .A2(n14783), .ZN(n14780) );
  OAI21_X1 U24502 ( .B1(n13069), .B2(n14780), .A(n15259), .ZN(n13062) );
  NAND2_X1 U24503 ( .A1(n13064), .A2(n3564), .ZN(n15251) );
  NAND2_X1 U24505 ( .A1(n13066), .A2(n15256), .ZN(n13074) );
  OAI22_X1 U24506 ( .A1(n15264), .A2(n15257), .B1(n14137), .B2(n14780), .ZN(
        n13068) );
  NOR2_X1 U24507 ( .A1(n14791), .A2(n14790), .ZN(n13067) );
  NAND2_X1 U24508 ( .A1(n51686), .A2(n14141), .ZN(n13070) );
  OAI21_X1 U24509 ( .B1(n14137), .B2(n15264), .A(n13070), .ZN(n13072) );
  NAND2_X1 U24510 ( .A1(n13075), .A2(n13089), .ZN(n13080) );
  INV_X1 U24511 ( .A(n13076), .ZN(n13079) );
  NAND2_X1 U24512 ( .A1(n13077), .A2(n13090), .ZN(n13078) );
  NOR2_X1 U24513 ( .A1(n13087), .A2(n13086), .ZN(n13097) );
  OAI211_X1 U24514 ( .C1(n13090), .C2(n13089), .A(n13103), .B(n13088), .ZN(
        n13096) );
  NAND3_X1 U24515 ( .A1(n13093), .A2(n13092), .A3(n13091), .ZN(n13094) );
  OAI211_X1 U24516 ( .C1(n13097), .C2(n13096), .A(n13095), .B(n13094), .ZN(
        n13098) );
  INV_X1 U24517 ( .A(n13098), .ZN(n13108) );
  NAND2_X1 U24518 ( .A1(n13106), .A2(n13105), .ZN(n13107) );
  NAND4_X1 U24519 ( .A1(n13764), .A2(n14150), .A3(n13124), .A4(n51175), .ZN(
        n13766) );
  INV_X1 U24520 ( .A(n13766), .ZN(n13111) );
  NAND2_X1 U24521 ( .A1(n13111), .A2(n13110), .ZN(n13121) );
  INV_X1 U24522 ( .A(n13763), .ZN(n13112) );
  NAND2_X1 U24523 ( .A1(n13112), .A2(n14155), .ZN(n13115) );
  AOI22_X1 U24524 ( .A1(n13115), .A2(n13762), .B1(n13114), .B2(n13113), .ZN(
        n13120) );
  NAND3_X1 U24525 ( .A1(n13117), .A2(n14159), .A3(n14160), .ZN(n13118) );
  OR2_X1 U24526 ( .A1(n14164), .A2(n14160), .ZN(n14146) );
  NAND2_X1 U24527 ( .A1(n14160), .A2(n14966), .ZN(n13123) );
  MUX2_X1 U24528 ( .A(n14146), .B(n13123), .S(n13122), .Z(n13128) );
  MUX2_X1 U24529 ( .A(n14150), .B(n51175), .S(n13124), .Z(n13127) );
  OAI21_X1 U24531 ( .B1(n13128), .B2(n13127), .A(n13126), .ZN(n13129) );
  NAND4_X1 U24532 ( .A1(n13139), .A2(n14179), .A3(n51136), .A4(n13130), .ZN(
        n13134) );
  NAND3_X1 U24533 ( .A1(n14191), .A2(n13132), .A3(n14179), .ZN(n13133) );
  AND2_X1 U24534 ( .A1(n13134), .A2(n13133), .ZN(n13159) );
  NOR2_X1 U24535 ( .A1(n13139), .A2(n13135), .ZN(n13141) );
  NAND2_X1 U24536 ( .A1(n13137), .A2(n13148), .ZN(n14185) );
  NOR2_X1 U24537 ( .A1(n14185), .A2(n13138), .ZN(n13140) );
  AOI22_X1 U24538 ( .A1(n13141), .A2(n14188), .B1(n13140), .B2(n13139), .ZN(
        n13158) );
  INV_X1 U24539 ( .A(n13145), .ZN(n13146) );
  NAND2_X1 U24540 ( .A1(n13146), .A2(n14186), .ZN(n13147) );
  OAI21_X1 U24541 ( .B1(n14191), .B2(n14187), .A(n13147), .ZN(n13149) );
  NAND2_X1 U24542 ( .A1(n13149), .A2(n13148), .ZN(n13155) );
  INV_X1 U24543 ( .A(n14183), .ZN(n13151) );
  NAND4_X1 U24544 ( .A1(n13153), .A2(n13152), .A3(n13151), .A4(n13150), .ZN(
        n13154) );
  INV_X1 U24545 ( .A(n13160), .ZN(n13163) );
  NAND2_X1 U24546 ( .A1(n13779), .A2(n13173), .ZN(n13162) );
  OAI211_X1 U24547 ( .C1(n13163), .C2(n13173), .A(n13177), .B(n13162), .ZN(
        n13165) );
  NAND3_X1 U24548 ( .A1(n13782), .A2(n13776), .A3(n13163), .ZN(n13164) );
  OAI211_X1 U24549 ( .C1(n13165), .C2(n13782), .A(n13778), .B(n13164), .ZN(
        n13184) );
  INV_X1 U24550 ( .A(n13166), .ZN(n13168) );
  NAND4_X1 U24551 ( .A1(n13171), .A2(n13170), .A3(n13172), .A4(n13780), .ZN(
        n13176) );
  NAND3_X1 U24552 ( .A1(n13174), .A2(n13173), .A3(n13172), .ZN(n13175) );
  AND2_X1 U24553 ( .A1(n13176), .A2(n13175), .ZN(n13182) );
  NAND3_X1 U24554 ( .A1(n13179), .A2(n13780), .A3(n13773), .ZN(n13180) );
  INV_X1 U24555 ( .A(n13189), .ZN(n13191) );
  INV_X1 U24556 ( .A(n13190), .ZN(n13950) );
  NAND2_X1 U24557 ( .A1(n13191), .A2(n13950), .ZN(n13195) );
  MUX2_X1 U24558 ( .A(n13195), .B(n13194), .S(n2173), .Z(n13213) );
  AOI22_X1 U24559 ( .A1(n13198), .A2(n13934), .B1(n13197), .B2(n13196), .ZN(
        n13199) );
  INV_X1 U24560 ( .A(n13200), .ZN(n13201) );
  NAND3_X1 U24561 ( .A1(n781), .A2(n13207), .A3(n13948), .ZN(n13203) );
  NAND3_X1 U24562 ( .A1(n13205), .A2(n13204), .A3(n13203), .ZN(n13211) );
  OR2_X1 U24563 ( .A1(n13948), .A2(n638), .ZN(n13940) );
  NAND2_X1 U24564 ( .A1(n1580), .A2(n13930), .ZN(n13935) );
  OAI211_X1 U24565 ( .C1(n13940), .C2(n13944), .A(n13209), .B(n13935), .ZN(
        n13210) );
  INV_X1 U24566 ( .A(n13214), .ZN(n13957) );
  NOR2_X1 U24567 ( .A1(n14224), .A2(n14220), .ZN(n13969) );
  NAND4_X1 U24568 ( .A1(n13957), .A2(n13969), .A3(n13215), .A4(n14234), .ZN(
        n13218) );
  NAND3_X1 U24569 ( .A1(n14223), .A2(n13970), .A3(n14220), .ZN(n13217) );
  NAND2_X1 U24570 ( .A1(n13216), .A2(n14224), .ZN(n13965) );
  AND3_X1 U24571 ( .A1(n13218), .A2(n13217), .A3(n13965), .ZN(n13251) );
  NOR2_X1 U24572 ( .A1(n14224), .A2(n13219), .ZN(n14227) );
  NAND3_X1 U24573 ( .A1(n13222), .A2(n13221), .A3(n13220), .ZN(n13223) );
  AND2_X1 U24574 ( .A1(n13224), .A2(n13223), .ZN(n13250) );
  INV_X1 U24575 ( .A(n13225), .ZN(n13243) );
  NAND2_X1 U24576 ( .A1(n13963), .A2(n13226), .ZN(n13242) );
  INV_X1 U24577 ( .A(n13227), .ZN(n13228) );
  NOR3_X1 U24578 ( .A1(n13229), .A2(n2468), .A3(n13228), .ZN(n13240) );
  NAND2_X1 U24579 ( .A1(n13231), .A2(n13230), .ZN(n13235) );
  INV_X1 U24580 ( .A(n13232), .ZN(n13234) );
  AOI21_X1 U24581 ( .B1(n13235), .B2(n13234), .A(n13233), .ZN(n13236) );
  NOR2_X1 U24582 ( .A1(n14228), .A2(n13236), .ZN(n13239) );
  INV_X1 U24583 ( .A(n13237), .ZN(n13238) );
  NAND4_X1 U24584 ( .A1(n13240), .A2(n13239), .A3(n14220), .A4(n13238), .ZN(
        n14232) );
  NAND2_X1 U24585 ( .A1(n14232), .A2(n13960), .ZN(n13241) );
  AOI22_X1 U24586 ( .A1(n13243), .A2(n13242), .B1(n13241), .B2(n13970), .ZN(
        n13249) );
  INV_X1 U24587 ( .A(n13244), .ZN(n13246) );
  NAND2_X1 U24588 ( .A1(n13960), .A2(n14221), .ZN(n13245) );
  OAI211_X1 U24589 ( .C1(n13247), .C2(n13969), .A(n13246), .B(n13245), .ZN(
        n13248) );
  NAND4_X2 U24590 ( .A1(n13251), .A2(n13250), .A3(n13249), .A4(n13248), .ZN(
        n16624) );
  INV_X1 U24592 ( .A(n14877), .ZN(n13254) );
  NAND2_X1 U24593 ( .A1(n7245), .A2(n14880), .ZN(n13253) );
  OAI22_X1 U24594 ( .A1(n13254), .A2(n13253), .B1(n15422), .B2(n1556), .ZN(
        n13255) );
  NOR2_X1 U24595 ( .A1(n50966), .A2(n15421), .ZN(n15426) );
  NAND3_X1 U24596 ( .A1(n15426), .A2(n1556), .A3(n13886), .ZN(n13258) );
  NOR3_X1 U24597 ( .A1(n13259), .A2(n14876), .A3(n14880), .ZN(n13260) );
  OR2_X1 U24598 ( .A1(n13261), .A2(n15425), .ZN(n13263) );
  XNOR2_X1 U24599 ( .A(n18408), .B(n17232), .ZN(n13266) );
  XNOR2_X1 U24600 ( .A(n13267), .B(n13266), .ZN(n13268) );
  NAND3_X1 U24601 ( .A1(n14763), .A2(n14767), .A3(n15233), .ZN(n13269) );
  OAI22_X1 U24602 ( .A1(n13269), .A2(n13277), .B1(n15206), .B2(n15196), .ZN(
        n13270) );
  NOR2_X1 U24603 ( .A1(n15187), .A2(n13270), .ZN(n13287) );
  OR2_X1 U24604 ( .A1(n13277), .A2(n15189), .ZN(n15207) );
  NOR2_X1 U24605 ( .A1(n15207), .A2(n15196), .ZN(n15241) );
  OR2_X1 U24606 ( .A1(n13271), .A2(n15206), .ZN(n14114) );
  NOR2_X1 U24607 ( .A1(n13272), .A2(n14114), .ZN(n13273) );
  NAND2_X1 U24609 ( .A1(n15189), .A2(n14767), .ZN(n15199) );
  OAI21_X1 U24610 ( .B1(n15188), .B2(n15236), .A(n15199), .ZN(n13275) );
  NAND3_X1 U24611 ( .A1(n15235), .A2(n15188), .A3(n15236), .ZN(n13279) );
  NAND2_X1 U24612 ( .A1(n15189), .A2(n15244), .ZN(n13281) );
  NOR2_X1 U24613 ( .A1(n15233), .A2(n14759), .ZN(n13276) );
  NAND4_X1 U24614 ( .A1(n13277), .A2(n13281), .A3(n14763), .A4(n13276), .ZN(
        n13278) );
  AND3_X1 U24615 ( .A1(n13280), .A2(n13279), .A3(n13278), .ZN(n13285) );
  INV_X1 U24616 ( .A(n13281), .ZN(n13283) );
  NOR2_X1 U24617 ( .A1(n15233), .A2(n14767), .ZN(n15193) );
  OAI211_X1 U24618 ( .C1(n14761), .C2(n13283), .A(n15193), .B(n13282), .ZN(
        n13284) );
  AND2_X1 U24620 ( .A1(n13729), .A2(n14022), .ZN(n14034) );
  NAND2_X1 U24621 ( .A1(n13303), .A2(n13729), .ZN(n13295) );
  NAND3_X1 U24622 ( .A1(n13304), .A2(n14030), .A3(n14022), .ZN(n13293) );
  NAND4_X1 U24623 ( .A1(n14032), .A2(n13297), .A3(n13303), .A4(n13291), .ZN(
        n13292) );
  NOR2_X1 U24624 ( .A1(n13296), .A2(n13295), .ZN(n13728) );
  NOR2_X1 U24625 ( .A1(n13297), .A2(n14030), .ZN(n13733) );
  NAND3_X1 U24626 ( .A1(n13733), .A2(n14032), .A3(n13298), .ZN(n13301) );
  NAND3_X1 U24628 ( .A1(n6726), .A2(n13303), .A3(n14030), .ZN(n14038) );
  OAI22_X1 U24629 ( .A1(n14022), .A2(n13736), .B1(n13304), .B2(n14032), .ZN(
        n13305) );
  NAND3_X1 U24630 ( .A1(n13305), .A2(n14033), .A3(n14030), .ZN(n13310) );
  AND2_X1 U24631 ( .A1(n13729), .A2(n13306), .ZN(n13307) );
  NOR2_X1 U24632 ( .A1(n14018), .A2(n13307), .ZN(n13727) );
  NAND4_X1 U24633 ( .A1(n13727), .A2(n13308), .A3(n782), .A4(n14028), .ZN(
        n13309) );
  XNOR2_X1 U24634 ( .A(n17891), .B(n51435), .ZN(n13345) );
  AOI22_X1 U24635 ( .A1(n13313), .A2(n14170), .B1(n13316), .B2(n14606), .ZN(
        n13315) );
  INV_X1 U24636 ( .A(n14603), .ZN(n13314) );
  NOR2_X1 U24637 ( .A1(n13317), .A2(n13316), .ZN(n14602) );
  INV_X1 U24638 ( .A(n14602), .ZN(n13319) );
  NOR2_X1 U24639 ( .A1(n14006), .A2(n13322), .ZN(n14596) );
  NAND3_X1 U24640 ( .A1(n14612), .A2(n14596), .A3(n14605), .ZN(n13318) );
  XNOR2_X1 U24642 ( .A(n14006), .B(n14600), .ZN(n13321) );
  AND2_X1 U24643 ( .A1(n13322), .A2(n14600), .ZN(n14008) );
  OAI21_X1 U24644 ( .B1(n14175), .B2(n14611), .A(n14008), .ZN(n13327) );
  INV_X1 U24646 ( .A(n14001), .ZN(n14004) );
  NAND3_X1 U24647 ( .A1(n14597), .A2(n14175), .A3(n14004), .ZN(n13326) );
  NAND4_X1 U24648 ( .A1(n13328), .A2(n13327), .A3(n13326), .A4(n13325), .ZN(
        n13329) );
  INV_X1 U24649 ( .A(n13331), .ZN(n13335) );
  NAND4_X1 U24650 ( .A1(n13335), .A2(n13742), .A3(n14719), .A4(n13743), .ZN(
        n13332) );
  NOR2_X1 U24651 ( .A1(n14711), .A2(n14704), .ZN(n14700) );
  NAND3_X1 U24652 ( .A1(n14720), .A2(n14709), .A3(n14716), .ZN(n13336) );
  OAI211_X1 U24653 ( .C1(n14199), .C2(n14717), .A(n14704), .B(n13336), .ZN(
        n13341) );
  NAND2_X1 U24654 ( .A1(n13337), .A2(n14709), .ZN(n13340) );
  NAND2_X1 U24655 ( .A1(n13338), .A2(n14711), .ZN(n13339) );
  INV_X1 U24656 ( .A(n14205), .ZN(n13751) );
  NOR2_X1 U24657 ( .A1(n14720), .A2(n14709), .ZN(n14202) );
  OR3_X1 U24658 ( .A1(n14202), .A2(n13343), .A3(n14713), .ZN(n13344) );
  OAI211_X1 U24659 ( .C1(n13751), .C2(n14200), .A(n14080), .B(n13344), .ZN(
        n14893) );
  XNOR2_X1 U24660 ( .A(n13345), .B(n18148), .ZN(n13399) );
  OAI21_X1 U24661 ( .B1(n13347), .B2(n14550), .A(n14548), .ZN(n13349) );
  NAND3_X1 U24662 ( .A1(n13347), .A2(n3038), .A3(n14550), .ZN(n13348) );
  NAND3_X1 U24663 ( .A1(n13349), .A2(n14365), .A3(n13348), .ZN(n13350) );
  NAND2_X1 U24664 ( .A1(n14370), .A2(n14553), .ZN(n13351) );
  NAND4_X1 U24665 ( .A1(n13353), .A2(n14545), .A3(n14370), .A4(n14542), .ZN(
        n13359) );
  NAND2_X1 U24666 ( .A1(n14533), .A2(n14550), .ZN(n13356) );
  NOR2_X1 U24667 ( .A1(n13354), .A2(n14370), .ZN(n13355) );
  NAND4_X1 U24668 ( .A1(n14536), .A2(n13356), .A3(n13355), .A4(n14552), .ZN(
        n13357) );
  OAI21_X1 U24669 ( .B1(n13362), .B2(n14536), .A(n13361), .ZN(n13364) );
  NAND3_X1 U24670 ( .A1(n14362), .A2(n14544), .A3(n13362), .ZN(n13363) );
  XNOR2_X1 U24671 ( .A(n4883), .B(Key[57]), .ZN(n22814) );
  XNOR2_X1 U24672 ( .A(n22814), .B(n4579), .ZN(n37138) );
  INV_X1 U24673 ( .A(n37138), .ZN(n13366) );
  XNOR2_X1 U24674 ( .A(n16628), .B(n13366), .ZN(n13397) );
  INV_X1 U24675 ( .A(n13367), .ZN(n13369) );
  NOR2_X1 U24676 ( .A1(n14519), .A2(n16036), .ZN(n13368) );
  OAI211_X1 U24677 ( .C1(n13370), .C2(n13369), .A(n13372), .B(n13368), .ZN(
        n13375) );
  INV_X1 U24678 ( .A(n13372), .ZN(n13373) );
  INV_X1 U24679 ( .A(n13376), .ZN(n13383) );
  NOR2_X1 U24680 ( .A1(n16049), .A2(n13377), .ZN(n14512) );
  AND2_X1 U24681 ( .A1(n51714), .A2(n16036), .ZN(n13379) );
  OAI21_X1 U24682 ( .B1(n14512), .B2(n13379), .A(n16045), .ZN(n13382) );
  NAND4_X1 U24683 ( .A1(n14519), .A2(n13380), .A3(n14527), .A4(n51018), .ZN(
        n13381) );
  AND3_X1 U24684 ( .A1(n13383), .A2(n13382), .A3(n13381), .ZN(n13395) );
  INV_X1 U24685 ( .A(n14529), .ZN(n16040) );
  OR2_X1 U24686 ( .A1(n13385), .A2(n6192), .ZN(n16035) );
  INV_X1 U24687 ( .A(n13386), .ZN(n13388) );
  NAND4_X1 U24688 ( .A1(n13388), .A2(n16044), .A3(n13387), .A4(n16039), .ZN(
        n13389) );
  NAND2_X1 U24690 ( .A1(n13392), .A2(n14515), .ZN(n13393) );
  NAND4_X2 U24691 ( .A1(n13394), .A2(n13395), .A3(n13393), .A4(n13396), .ZN(
        n17758) );
  XNOR2_X1 U24692 ( .A(n17758), .B(n13397), .ZN(n15473) );
  INV_X1 U24693 ( .A(n15473), .ZN(n13398) );
  XNOR2_X1 U24694 ( .A(n13399), .B(n13398), .ZN(n13536) );
  NAND3_X1 U24695 ( .A1(n14346), .A2(n13400), .A3(n13422), .ZN(n13407) );
  INV_X1 U24696 ( .A(n13401), .ZN(n13406) );
  INV_X1 U24697 ( .A(n13402), .ZN(n13403) );
  NAND3_X1 U24698 ( .A1(n13404), .A2(n13403), .A3(n14344), .ZN(n13405) );
  NOR2_X1 U24699 ( .A1(n14339), .A2(n14344), .ZN(n13408) );
  AOI22_X1 U24700 ( .A1(n13408), .A2(n14342), .B1(n14339), .B2(n6073), .ZN(
        n13416) );
  INV_X1 U24701 ( .A(n14338), .ZN(n13409) );
  OAI21_X1 U24702 ( .B1(n14337), .B2(n13409), .A(n14346), .ZN(n13415) );
  NAND3_X1 U24703 ( .A1(n14342), .A2(n6073), .A3(n14331), .ZN(n13413) );
  NAND2_X1 U24704 ( .A1(n6073), .A2(n13410), .ZN(n13411) );
  NAND3_X1 U24705 ( .A1(n13413), .A2(n13412), .A3(n13411), .ZN(n13414) );
  OAI211_X1 U24706 ( .C1(n13416), .C2(n14346), .A(n13415), .B(n13414), .ZN(
        n13428) );
  AND3_X1 U24707 ( .A1(n13418), .A2(n14344), .A3(n13417), .ZN(n13420) );
  AOI21_X1 U24708 ( .B1(n13420), .B2(n14346), .A(n13419), .ZN(n13427) );
  INV_X1 U24709 ( .A(n13421), .ZN(n14352) );
  INV_X1 U24710 ( .A(n13422), .ZN(n13423) );
  INV_X1 U24711 ( .A(n13429), .ZN(n13433) );
  INV_X1 U24712 ( .A(n13437), .ZN(n13455) );
  OAI21_X1 U24713 ( .B1(n13438), .B2(n4383), .A(n14655), .ZN(n13444) );
  NOR2_X1 U24714 ( .A1(n13445), .A2(n13439), .ZN(n13443) );
  OAI21_X1 U24715 ( .B1(n13444), .B2(n13443), .A(n13442), .ZN(n13454) );
  OAI22_X1 U24716 ( .A1(n14660), .A2(n13450), .B1(n13449), .B2(n13448), .ZN(
        n13451) );
  NAND2_X1 U24717 ( .A1(n13451), .A2(n13995), .ZN(n13452) );
  XNOR2_X1 U24718 ( .A(n18668), .B(n637), .ZN(n13474) );
  INV_X1 U24719 ( .A(n51369), .ZN(n15179) );
  NAND2_X1 U24720 ( .A1(n15165), .A2(n14574), .ZN(n13461) );
  OAI21_X1 U24721 ( .B1(n15159), .B2(n14574), .A(n13461), .ZN(n13469) );
  INV_X1 U24722 ( .A(n13462), .ZN(n13465) );
  INV_X1 U24723 ( .A(n14572), .ZN(n13466) );
  AOI21_X1 U24724 ( .B1(n13466), .B2(n15167), .A(n15163), .ZN(n13467) );
  INV_X1 U24725 ( .A(n4587), .ZN(n45866) );
  XNOR2_X1 U24726 ( .A(n45866), .B(n4937), .ZN(n17757) );
  INV_X1 U24727 ( .A(n17757), .ZN(n34411) );
  XNOR2_X1 U24728 ( .A(Key[171]), .B(n4739), .ZN(n42101) );
  XNOR2_X1 U24729 ( .A(n34411), .B(n42101), .ZN(n24200) );
  XNOR2_X1 U24730 ( .A(n45107), .B(n4451), .ZN(n13568) );
  XNOR2_X1 U24731 ( .A(n24200), .B(n13568), .ZN(n24010) );
  XNOR2_X1 U24732 ( .A(n24010), .B(n4605), .ZN(n31135) );
  XNOR2_X1 U24733 ( .A(Key[69]), .B(Key[111]), .ZN(n33429) );
  XNOR2_X1 U24734 ( .A(n4940), .B(n4565), .ZN(n36738) );
  XNOR2_X1 U24735 ( .A(n43368), .B(n36738), .ZN(n13470) );
  XNOR2_X1 U24736 ( .A(n45105), .B(n13470), .ZN(n13471) );
  XNOR2_X1 U24737 ( .A(n31135), .B(n13471), .ZN(n13472) );
  XNOR2_X1 U24738 ( .A(n17707), .B(n13472), .ZN(n13473) );
  XNOR2_X1 U24739 ( .A(n13474), .B(n13473), .ZN(n13535) );
  NAND2_X1 U24740 ( .A1(n69), .A2(n13804), .ZN(n13479) );
  NOR2_X1 U24742 ( .A1(n15044), .A2(n15034), .ZN(n13476) );
  AOI22_X1 U24743 ( .A1(n13476), .A2(n15030), .B1(n13480), .B2(n15048), .ZN(
        n13477) );
  NAND2_X1 U24744 ( .A1(n13798), .A2(n15046), .ZN(n15029) );
  OAI211_X1 U24745 ( .C1(n15029), .C2(n13483), .A(n15040), .B(n13482), .ZN(
        n13484) );
  INV_X1 U24746 ( .A(n13484), .ZN(n13495) );
  NOR2_X1 U24747 ( .A1(n15034), .A2(n13800), .ZN(n13485) );
  XNOR2_X1 U24748 ( .A(n69), .B(n13485), .ZN(n13491) );
  INV_X1 U24749 ( .A(n13486), .ZN(n13490) );
  NAND2_X1 U24750 ( .A1(n13487), .A2(n15034), .ZN(n13489) );
  NAND2_X1 U24751 ( .A1(n15034), .A2(n13797), .ZN(n15041) );
  NOR2_X1 U24752 ( .A1(n15041), .A2(n13801), .ZN(n13493) );
  OAI21_X1 U24753 ( .B1(n13493), .B2(n13492), .A(n15038), .ZN(n13494) );
  NAND4_X1 U24754 ( .A1(n13529), .A2(n13502), .A3(n13501), .A4(n13500), .ZN(
        n13510) );
  NAND2_X1 U24755 ( .A1(n13503), .A2(n9357), .ZN(n13508) );
  NAND3_X1 U24756 ( .A1(n13506), .A2(n13505), .A3(n51067), .ZN(n13507) );
  OAI211_X1 U24757 ( .C1(n13510), .C2(n13509), .A(n13508), .B(n13507), .ZN(
        n13519) );
  NAND3_X1 U24758 ( .A1(n13515), .A2(n13514), .A3(n13513), .ZN(n13516) );
  NAND2_X1 U24759 ( .A1(n13517), .A2(n13516), .ZN(n13518) );
  NOR2_X1 U24760 ( .A1(n13519), .A2(n13518), .ZN(n13534) );
  NAND3_X1 U24761 ( .A1(n13522), .A2(n13521), .A3(n51683), .ZN(n13523) );
  AND2_X1 U24762 ( .A1(n13524), .A2(n13523), .ZN(n13533) );
  NAND2_X1 U24763 ( .A1(n13526), .A2(n13525), .ZN(n13528) );
  OAI21_X1 U24764 ( .B1(n13529), .B2(n13528), .A(n13527), .ZN(n13531) );
  NAND2_X1 U24765 ( .A1(n13531), .A2(n13530), .ZN(n13532) );
  MUX2_X1 U24766 ( .A(n18023), .B(n17484), .S(n17569), .Z(n13537) );
  AOI21_X1 U24767 ( .B1(n13537), .B2(n17568), .A(n19398), .ZN(n13538) );
  AOI21_X1 U24768 ( .B1(n13539), .B2(n17484), .A(n13538), .ZN(n13544) );
  NAND2_X1 U24769 ( .A1(n18022), .A2(n18013), .ZN(n13541) );
  INV_X1 U24770 ( .A(n13540), .ZN(n18010) );
  MUX2_X1 U24771 ( .A(n13542), .B(n13541), .S(n19395), .Z(n13543) );
  INV_X1 U24772 ( .A(n21780), .ZN(n21117) );
  INV_X1 U24773 ( .A(n14477), .ZN(n13546) );
  NAND4_X1 U24774 ( .A1(n7465), .A2(n14482), .A3(n14472), .A4(n13855), .ZN(
        n13545) );
  OAI211_X1 U24775 ( .C1(n13548), .C2(n13547), .A(n13546), .B(n13545), .ZN(
        n13549) );
  MUX2_X1 U24776 ( .A(n13549), .B(n13552), .S(n13853), .Z(n13567) );
  INV_X1 U24777 ( .A(n13843), .ZN(n14476) );
  AOI21_X1 U24778 ( .B1(n14476), .B2(n13551), .A(n14883), .ZN(n13565) );
  INV_X1 U24779 ( .A(n13552), .ZN(n13553) );
  OAI21_X1 U24780 ( .B1(n13841), .B2(n13553), .A(n14883), .ZN(n13555) );
  OR2_X1 U24781 ( .A1(n13855), .A2(n14472), .ZN(n13848) );
  NOR2_X1 U24782 ( .A1(n14474), .A2(n13848), .ZN(n13554) );
  NOR2_X1 U24783 ( .A1(n13555), .A2(n13554), .ZN(n13564) );
  INV_X1 U24784 ( .A(n13848), .ZN(n13558) );
  INV_X1 U24785 ( .A(n13850), .ZN(n13556) );
  OAI211_X1 U24786 ( .C1(n13558), .C2(n13849), .A(n13557), .B(n13843), .ZN(
        n13563) );
  AOI22_X1 U24787 ( .A1(n13851), .A2(n13561), .B1(n13560), .B2(n13559), .ZN(
        n13562) );
  OAI211_X1 U24788 ( .C1(n13565), .C2(n13564), .A(n13563), .B(n13562), .ZN(
        n13566) );
  XNOR2_X1 U24790 ( .A(n17879), .B(n4793), .ZN(n16323) );
  XNOR2_X1 U24791 ( .A(n45883), .B(n4501), .ZN(n44044) );
  XNOR2_X1 U24792 ( .A(n44044), .B(n45106), .ZN(n25470) );
  XNOR2_X1 U24793 ( .A(n25470), .B(n801), .ZN(n41183) );
  XNOR2_X1 U24794 ( .A(Key[153]), .B(n4565), .ZN(n44934) );
  XNOR2_X1 U24795 ( .A(n44934), .B(n4431), .ZN(n20856) );
  XNOR2_X1 U24796 ( .A(n41183), .B(n20856), .ZN(n24707) );
  XNOR2_X1 U24797 ( .A(n41155), .B(n4883), .ZN(n16112) );
  XNOR2_X1 U24798 ( .A(n24707), .B(n16112), .ZN(n37301) );
  XNOR2_X1 U24799 ( .A(n13568), .B(n1224), .ZN(n41161) );
  XNOR2_X1 U24800 ( .A(n41161), .B(n33049), .ZN(n13569) );
  XNOR2_X1 U24801 ( .A(n37301), .B(n13569), .ZN(n13570) );
  XNOR2_X1 U24802 ( .A(n16323), .B(n13570), .ZN(n13571) );
  XNOR2_X1 U24803 ( .A(n13572), .B(n13571), .ZN(n13720) );
  NAND3_X1 U24804 ( .A1(n5411), .A2(n13573), .A3(n13583), .ZN(n13980) );
  NAND2_X1 U24805 ( .A1(n14276), .A2(n13980), .ZN(n13581) );
  NAND2_X1 U24806 ( .A1(n5411), .A2(n13576), .ZN(n13578) );
  NAND3_X1 U24807 ( .A1(n13579), .A2(n13578), .A3(n13577), .ZN(n13580) );
  NOR2_X1 U24808 ( .A1(n13581), .A2(n13580), .ZN(n13597) );
  NAND2_X1 U24809 ( .A1(n14286), .A2(n13583), .ZN(n13585) );
  MUX2_X1 U24810 ( .A(n13586), .B(n13585), .S(n13584), .Z(n13596) );
  OAI21_X1 U24811 ( .B1(n13588), .B2(n13979), .A(n14280), .ZN(n13589) );
  NAND4_X1 U24812 ( .A1(n13591), .A2(n13590), .A3(n14285), .A4(n13589), .ZN(
        n13595) );
  INV_X1 U24813 ( .A(n14296), .ZN(n13593) );
  NAND3_X1 U24814 ( .A1(n13593), .A2(n13592), .A3(n14290), .ZN(n13594) );
  NAND4_X2 U24815 ( .A1(n13597), .A2(n13596), .A3(n13594), .A4(n13595), .ZN(
        n17138) );
  NAND2_X1 U24816 ( .A1(n51064), .A2(n14317), .ZN(n13823) );
  INV_X1 U24817 ( .A(n13823), .ZN(n13602) );
  NOR2_X1 U24818 ( .A1(n14318), .A2(n14311), .ZN(n13601) );
  AND2_X1 U24819 ( .A1(n14311), .A2(n13826), .ZN(n13825) );
  AOI22_X1 U24820 ( .A1(n13602), .A2(n13601), .B1(n13600), .B2(n13825), .ZN(
        n13619) );
  NAND2_X1 U24821 ( .A1(n13819), .A2(n13822), .ZN(n13603) );
  NOR2_X1 U24822 ( .A1(n13604), .A2(n13603), .ZN(n13607) );
  NOR2_X1 U24823 ( .A1(n13605), .A2(n14318), .ZN(n13606) );
  AOI22_X1 U24824 ( .A1(n13607), .A2(n14318), .B1(n13606), .B2(n14322), .ZN(
        n13618) );
  INV_X1 U24825 ( .A(n14308), .ZN(n13608) );
  NAND2_X1 U24826 ( .A1(n13827), .A2(n13826), .ZN(n13612) );
  NAND3_X1 U24827 ( .A1(n13820), .A2(n13826), .A3(n14320), .ZN(n13611) );
  NAND4_X1 U24828 ( .A1(n13612), .A2(n13611), .A3(n13610), .A4(n13819), .ZN(
        n13615) );
  NAND3_X1 U24829 ( .A1(n14321), .A2(n14310), .A3(n14318), .ZN(n13614) );
  NAND2_X1 U24830 ( .A1(n14319), .A2(n14320), .ZN(n13613) );
  INV_X1 U24832 ( .A(n13620), .ZN(n13621) );
  NAND4_X1 U24833 ( .A1(n13622), .A2(n51347), .A3(n13633), .A4(n13621), .ZN(
        n13626) );
  INV_X1 U24834 ( .A(n13623), .ZN(n13624) );
  OR2_X1 U24835 ( .A1(n13624), .A2(n13633), .ZN(n13625) );
  AND4_X1 U24836 ( .A1(n13628), .A2(n13627), .A3(n13626), .A4(n13625), .ZN(
        n13638) );
  NAND2_X1 U24837 ( .A1(n13631), .A2(n13630), .ZN(n13636) );
  NAND3_X1 U24838 ( .A1(n13634), .A2(n13633), .A3(n13632), .ZN(n13635) );
  NAND4_X1 U24839 ( .A1(n13638), .A2(n13637), .A3(n13636), .A4(n13635), .ZN(
        n13644) );
  NAND2_X1 U24840 ( .A1(n13640), .A2(n13639), .ZN(n13642) );
  MUX2_X1 U24841 ( .A(n13642), .B(n13641), .S(n14664), .Z(n13643) );
  OR2_X2 U24842 ( .A1(n13644), .A2(n13643), .ZN(n18147) );
  XNOR2_X1 U24843 ( .A(n15396), .B(n16730), .ZN(n15824) );
  XNOR2_X1 U24844 ( .A(n15824), .B(n51668), .ZN(n13719) );
  INV_X1 U24845 ( .A(n13645), .ZN(n13648) );
  NOR2_X1 U24846 ( .A1(n13658), .A2(n13646), .ZN(n13647) );
  MUX2_X1 U24847 ( .A(n13648), .B(n13647), .S(n14641), .Z(n13649) );
  INV_X1 U24848 ( .A(n13649), .ZN(n13675) );
  NOR2_X1 U24849 ( .A1(n14637), .A2(n13650), .ZN(n13652) );
  OAI22_X1 U24850 ( .A1(n13652), .A2(n13651), .B1(n2114), .B2(n14632), .ZN(
        n13657) );
  INV_X1 U24851 ( .A(n13653), .ZN(n13655) );
  OAI21_X1 U24852 ( .B1(n14640), .B2(n13655), .A(n13654), .ZN(n13656) );
  NOR2_X1 U24853 ( .A1(n13657), .A2(n13656), .ZN(n13674) );
  NAND3_X1 U24854 ( .A1(n14633), .A2(n14641), .A3(n2114), .ZN(n13660) );
  INV_X1 U24856 ( .A(n13662), .ZN(n13665) );
  OR2_X1 U24857 ( .A1(n14641), .A2(n13667), .ZN(n13663) );
  OAI21_X1 U24859 ( .B1(n13668), .B2(n8128), .A(n13666), .ZN(n13670) );
  NOR2_X1 U24861 ( .A1(n14252), .A2(n13683), .ZN(n13688) );
  AND2_X1 U24863 ( .A1(n13676), .A2(n13677), .ZN(n13694) );
  OR2_X1 U24864 ( .A1(n14982), .A2(n14983), .ZN(n14978) );
  NAND2_X1 U24865 ( .A1(n14984), .A2(n14252), .ZN(n13679) );
  NAND3_X1 U24866 ( .A1(n14978), .A2(n15103), .A3(n13683), .ZN(n13678) );
  OAI21_X1 U24867 ( .B1(n14978), .B2(n13679), .A(n13678), .ZN(n13680) );
  NAND2_X1 U24868 ( .A1(n13680), .A2(n352), .ZN(n13693) );
  NAND2_X1 U24869 ( .A1(n14252), .A2(n13683), .ZN(n15113) );
  INV_X1 U24870 ( .A(n15113), .ZN(n13681) );
  AND2_X1 U24872 ( .A1(n14982), .A2(n14983), .ZN(n15107) );
  INV_X1 U24873 ( .A(n15107), .ZN(n13685) );
  XNOR2_X1 U24874 ( .A(n15103), .B(n14252), .ZN(n13684) );
  NAND4_X1 U24875 ( .A1(n13685), .A2(n13684), .A3(n15117), .A4(n13683), .ZN(
        n13686) );
  AND2_X1 U24876 ( .A1(n13687), .A2(n13686), .ZN(n13692) );
  AND2_X1 U24877 ( .A1(n13688), .A2(n15103), .ZN(n13689) );
  NAND4_X1 U24878 ( .A1(n13690), .A2(n14245), .A3(n13689), .A4(n14247), .ZN(
        n13691) );
  INV_X1 U24880 ( .A(n14267), .ZN(n13695) );
  NOR2_X1 U24881 ( .A1(n13698), .A2(n15133), .ZN(n13699) );
  NOR2_X1 U24882 ( .A1(n13700), .A2(n13699), .ZN(n13706) );
  NAND4_X1 U24885 ( .A1(n13707), .A2(n13706), .A3(n13705), .A4(n13704), .ZN(
        n13718) );
  NAND2_X1 U24886 ( .A1(n14268), .A2(n13708), .ZN(n13716) );
  NOR2_X1 U24887 ( .A1(n14271), .A2(n15132), .ZN(n14262) );
  INV_X1 U24888 ( .A(n14992), .ZN(n13710) );
  NAND3_X1 U24889 ( .A1(n13711), .A2(n14262), .A3(n13710), .ZN(n13714) );
  NOR2_X1 U24890 ( .A1(n15133), .A2(n14271), .ZN(n13712) );
  INV_X1 U24891 ( .A(n14260), .ZN(n14272) );
  OAI21_X1 U24892 ( .B1(n13712), .B2(n14272), .A(n14994), .ZN(n13713) );
  OAI211_X1 U24893 ( .C1(n13716), .C2(n13715), .A(n13714), .B(n13713), .ZN(
        n13717) );
  XNOR2_X1 U24894 ( .A(n19210), .B(n13719), .ZN(n15575) );
  NOR2_X1 U24896 ( .A1(n14681), .A2(n14057), .ZN(n14686) );
  NAND2_X1 U24897 ( .A1(n14962), .A2(n51500), .ZN(n13721) );
  NOR2_X1 U24898 ( .A1(n15286), .A2(n13721), .ZN(n13722) );
  NOR2_X1 U24899 ( .A1(n14686), .A2(n13722), .ZN(n13726) );
  NAND2_X1 U24900 ( .A1(n14962), .A2(n2151), .ZN(n14951) );
  NAND2_X1 U24901 ( .A1(n2151), .A2(n14957), .ZN(n15280) );
  NAND2_X1 U24902 ( .A1(n14951), .A2(n15280), .ZN(n13723) );
  NAND4_X1 U24903 ( .A1(n51724), .A2(n14938), .A3(n51500), .A4(n14059), .ZN(
        n13725) );
  XNOR2_X1 U24904 ( .A(n461), .B(n51031), .ZN(n13754) );
  INV_X1 U24905 ( .A(n13727), .ZN(n13732) );
  INV_X1 U24906 ( .A(n13728), .ZN(n13731) );
  NAND2_X1 U24907 ( .A1(n14021), .A2(n13729), .ZN(n13730) );
  OAI211_X1 U24908 ( .C1(n13732), .C2(n14030), .A(n13731), .B(n13730), .ZN(
        n13740) );
  INV_X1 U24909 ( .A(n13733), .ZN(n13735) );
  INV_X1 U24910 ( .A(n14718), .ZN(n13741) );
  OAI21_X1 U24911 ( .B1(n13742), .B2(n14202), .A(n13741), .ZN(n13748) );
  NAND2_X1 U24912 ( .A1(n14721), .A2(n14711), .ZN(n14198) );
  INV_X1 U24913 ( .A(n13742), .ZN(n13745) );
  INV_X1 U24914 ( .A(n13743), .ZN(n13744) );
  AND2_X1 U24916 ( .A1(n14709), .A2(n14712), .ZN(n14722) );
  NAND3_X1 U24917 ( .A1(n14701), .A2(n14722), .A3(n14085), .ZN(n13746) );
  OR2_X1 U24919 ( .A1(n13749), .A2(n14718), .ZN(n13750) );
  OAI21_X1 U24920 ( .B1(n13751), .B2(n14200), .A(n13750), .ZN(n13752) );
  XNOR2_X1 U24921 ( .A(n17158), .B(n18175), .ZN(n15579) );
  INV_X1 U24922 ( .A(n15579), .ZN(n16428) );
  XNOR2_X1 U24923 ( .A(n13754), .B(n16428), .ZN(n16517) );
  XNOR2_X1 U24924 ( .A(Key[42]), .B(Key[66]), .ZN(n25114) );
  XNOR2_X1 U24925 ( .A(n25114), .B(n36755), .ZN(n26370) );
  XNOR2_X1 U24926 ( .A(Key[6]), .B(Key[30]), .ZN(n26297) );
  XNOR2_X1 U24927 ( .A(n26370), .B(n26297), .ZN(n16251) );
  INV_X1 U24928 ( .A(n16251), .ZN(n18171) );
  XNOR2_X1 U24929 ( .A(n18171), .B(n41567), .ZN(n16509) );
  INV_X1 U24930 ( .A(n16509), .ZN(n13755) );
  XNOR2_X1 U24931 ( .A(n4415), .B(Key[18]), .ZN(n27483) );
  XNOR2_X1 U24932 ( .A(n27483), .B(n1336), .ZN(n28270) );
  XNOR2_X1 U24933 ( .A(n13755), .B(n28270), .ZN(n35392) );
  XNOR2_X1 U24934 ( .A(n38626), .B(n4931), .ZN(n44193) );
  XNOR2_X1 U24935 ( .A(n44193), .B(n4536), .ZN(n13756) );
  XNOR2_X1 U24936 ( .A(n13756), .B(n42619), .ZN(n35479) );
  XNOR2_X1 U24937 ( .A(n35479), .B(n4847), .ZN(n13757) );
  XNOR2_X1 U24938 ( .A(n35392), .B(n13757), .ZN(n13758) );
  XNOR2_X1 U24939 ( .A(n15957), .B(n13758), .ZN(n13769) );
  AND2_X1 U24940 ( .A1(n14149), .A2(n13761), .ZN(n14154) );
  AOI22_X1 U24941 ( .A1(n13763), .A2(n13762), .B1(n14154), .B2(n14155), .ZN(
        n13767) );
  XNOR2_X1 U24942 ( .A(n17218), .B(n17901), .ZN(n13768) );
  XNOR2_X1 U24943 ( .A(n13769), .B(n13768), .ZN(n13770) );
  INV_X1 U24944 ( .A(n13773), .ZN(n13775) );
  OAI21_X1 U24945 ( .B1(n13776), .B2(n13775), .A(n13774), .ZN(n13777) );
  MUX2_X1 U24947 ( .A(n13784), .B(n13783), .S(n13782), .Z(n13785) );
  AOI21_X1 U24949 ( .B1(n15081), .B2(n2189), .A(n15766), .ZN(n13793) );
  NAND2_X1 U24950 ( .A1(n1486), .A2(n14911), .ZN(n14919) );
  NOR2_X1 U24951 ( .A1(n15300), .A2(n14911), .ZN(n15305) );
  OAI22_X1 U24952 ( .A1(n14919), .A2(n15068), .B1(n15305), .B2(n15770), .ZN(
        n13792) );
  INV_X1 U24953 ( .A(n15767), .ZN(n15306) );
  NAND2_X1 U24954 ( .A1(n15068), .A2(n15309), .ZN(n13788) );
  INV_X1 U24955 ( .A(n13794), .ZN(n13796) );
  NAND3_X1 U24956 ( .A1(n13796), .A2(n13800), .A3(n13795), .ZN(n13810) );
  NAND2_X1 U24957 ( .A1(n13798), .A2(n13797), .ZN(n13799) );
  AND2_X1 U24958 ( .A1(n15040), .A2(n13799), .ZN(n13809) );
  OAI21_X1 U24959 ( .B1(n13800), .B2(n13801), .A(n15035), .ZN(n13803) );
  NAND2_X1 U24960 ( .A1(n51966), .A2(n13801), .ZN(n13802) );
  OAI211_X1 U24961 ( .C1(n15034), .C2(n13804), .A(n13803), .B(n13802), .ZN(
        n13808) );
  NOR2_X1 U24962 ( .A1(n13805), .A2(n15034), .ZN(n15031) );
  XNOR2_X1 U24963 ( .A(n511), .B(n17145), .ZN(n19229) );
  XNOR2_X1 U24964 ( .A(n2121), .B(n17771), .ZN(n15812) );
  XNOR2_X1 U24965 ( .A(n2215), .B(n15812), .ZN(n16096) );
  XNOR2_X1 U24966 ( .A(n16096), .B(n19229), .ZN(n13811) );
  NAND2_X1 U24967 ( .A1(n13812), .A2(n14345), .ZN(n13813) );
  XNOR2_X1 U24968 ( .A(n17787), .B(n18447), .ZN(n13837) );
  NAND2_X1 U24969 ( .A1(n13821), .A2(n13820), .ZN(n13836) );
  NAND2_X1 U24970 ( .A1(n13825), .A2(n14321), .ZN(n13829) );
  NAND4_X1 U24971 ( .A1(n13830), .A2(n14307), .A3(n13829), .A4(n13828), .ZN(
        n13835) );
  NAND4_X1 U24972 ( .A1(n14312), .A2(n14321), .A3(n14320), .A4(n14311), .ZN(
        n13834) );
  NAND2_X1 U24973 ( .A1(n13832), .A2(n13831), .ZN(n13833) );
  XNOR2_X1 U24974 ( .A(n14803), .B(n51135), .ZN(n17788) );
  XNOR2_X1 U24975 ( .A(n13837), .B(n17788), .ZN(n13867) );
  NAND2_X1 U24976 ( .A1(n13856), .A2(n14472), .ZN(n13838) );
  NAND2_X1 U24977 ( .A1(n13839), .A2(n13838), .ZN(n13840) );
  NAND2_X1 U24978 ( .A1(n13840), .A2(n14482), .ZN(n13847) );
  NAND3_X1 U24979 ( .A1(n13841), .A2(n13856), .A3(n13855), .ZN(n13842) );
  OAI211_X1 U24980 ( .C1(n13845), .C2(n13844), .A(n13843), .B(n13842), .ZN(
        n13846) );
  NOR2_X1 U24981 ( .A1(n13853), .A2(n13848), .ZN(n13852) );
  AOI22_X1 U24982 ( .A1(n13852), .A2(n13851), .B1(n13850), .B2(n13849), .ZN(
        n13860) );
  NAND3_X1 U24983 ( .A1(n14885), .A2(n13853), .A3(n14482), .ZN(n13859) );
  OAI21_X1 U24984 ( .B1(n13856), .B2(n13855), .A(n13854), .ZN(n13857) );
  NAND2_X1 U24985 ( .A1(n14477), .A2(n13857), .ZN(n13858) );
  XNOR2_X1 U24986 ( .A(Key[131]), .B(Key[107]), .ZN(n45051) );
  XNOR2_X1 U24987 ( .A(n45051), .B(n4694), .ZN(n17254) );
  XNOR2_X1 U24988 ( .A(n17254), .B(n23943), .ZN(n13862) );
  XNOR2_X1 U24989 ( .A(n26525), .B(n34265), .ZN(n25897) );
  XNOR2_X1 U24990 ( .A(n13862), .B(n25897), .ZN(n43713) );
  XNOR2_X1 U24991 ( .A(n32856), .B(n4627), .ZN(n23722) );
  XNOR2_X1 U24992 ( .A(n43713), .B(n23722), .ZN(n33216) );
  XNOR2_X1 U24993 ( .A(n27353), .B(n48843), .ZN(n24314) );
  XNOR2_X1 U24994 ( .A(n24314), .B(n7744), .ZN(n42920) );
  XNOR2_X1 U24995 ( .A(n4781), .B(n4612), .ZN(n15142) );
  XNOR2_X1 U24996 ( .A(n15142), .B(n4287), .ZN(n13863) );
  XNOR2_X1 U24997 ( .A(n42920), .B(n13863), .ZN(n34866) );
  XNOR2_X1 U24998 ( .A(n33216), .B(n34866), .ZN(n13864) );
  XNOR2_X1 U24999 ( .A(n16016), .B(n13864), .ZN(n13865) );
  XNOR2_X1 U25000 ( .A(n13866), .B(n13867), .ZN(n13871) );
  XNOR2_X1 U25001 ( .A(n17665), .B(n16919), .ZN(n15950) );
  INV_X1 U25002 ( .A(n16228), .ZN(n13868) );
  XNOR2_X1 U25003 ( .A(n15950), .B(n13868), .ZN(n15593) );
  INV_X1 U25004 ( .A(n15593), .ZN(n13869) );
  XNOR2_X1 U25005 ( .A(n16454), .B(n13869), .ZN(n13870) );
  XNOR2_X1 U25006 ( .A(n13871), .B(n13870), .ZN(n13976) );
  INV_X1 U25007 ( .A(n16023), .ZN(n13893) );
  INV_X1 U25008 ( .A(n13873), .ZN(n13879) );
  NOR2_X1 U25009 ( .A1(n15425), .A2(n13874), .ZN(n13878) );
  INV_X1 U25010 ( .A(n13875), .ZN(n13877) );
  AND3_X1 U25011 ( .A1(n14880), .A2(n14871), .A3(n15425), .ZN(n13876) );
  AOI22_X1 U25012 ( .A1(n13879), .A2(n13878), .B1(n13877), .B2(n13876), .ZN(
        n13891) );
  AOI21_X1 U25013 ( .B1(n15421), .B2(n15425), .A(n14880), .ZN(n13880) );
  NAND2_X1 U25014 ( .A1(n13881), .A2(n50966), .ZN(n13882) );
  OAI211_X1 U25015 ( .C1(n14875), .C2(n14870), .A(n14873), .B(n13882), .ZN(
        n13883) );
  NAND3_X1 U25017 ( .A1(n13886), .A2(n13885), .A3(n1556), .ZN(n13887) );
  NAND2_X1 U25018 ( .A1(n15434), .A2(n15324), .ZN(n15436) );
  NAND3_X1 U25019 ( .A1(n13896), .A2(n13895), .A3(n13894), .ZN(n13898) );
  OAI211_X1 U25020 ( .C1(n13898), .C2(n13897), .A(n15335), .B(n15324), .ZN(
        n13899) );
  AND2_X1 U25021 ( .A1(n15436), .A2(n13899), .ZN(n13901) );
  NAND3_X1 U25022 ( .A1(n15343), .A2(n15332), .A3(n15325), .ZN(n13900) );
  INV_X1 U25023 ( .A(n15440), .ZN(n14861) );
  MUX2_X1 U25024 ( .A(n13901), .B(n13900), .S(n14861), .Z(n13912) );
  NOR2_X1 U25027 ( .A1(n15440), .A2(n15341), .ZN(n15431) );
  INV_X1 U25028 ( .A(n15431), .ZN(n13906) );
  NAND2_X1 U25029 ( .A1(n15435), .A2(n15434), .ZN(n15323) );
  INV_X1 U25030 ( .A(n15323), .ZN(n13904) );
  NAND2_X1 U25031 ( .A1(n13904), .A2(n15343), .ZN(n13905) );
  INV_X1 U25032 ( .A(n14863), .ZN(n15446) );
  OAI211_X1 U25033 ( .C1(n13907), .C2(n13906), .A(n13905), .B(n15446), .ZN(
        n13908) );
  NAND2_X1 U25034 ( .A1(n13908), .A2(n15438), .ZN(n13910) );
  INV_X1 U25035 ( .A(n14860), .ZN(n13909) );
  NAND4_X1 U25036 ( .A1(n13912), .A2(n13911), .A3(n13910), .A4(n13909), .ZN(
        n15688) );
  NOR2_X1 U25037 ( .A1(n15363), .A2(n15358), .ZN(n14818) );
  NAND2_X1 U25038 ( .A1(n15381), .A2(n14491), .ZN(n13913) );
  NOR2_X1 U25039 ( .A1(n15363), .A2(n13913), .ZN(n13915) );
  NOR2_X1 U25040 ( .A1(n13914), .A2(n15358), .ZN(n14490) );
  AOI22_X1 U25041 ( .A1(n14818), .A2(n15386), .B1(n13915), .B2(n14490), .ZN(
        n13928) );
  NAND4_X1 U25042 ( .A1(n13918), .A2(n15381), .A3(n13916), .A4(n14485), .ZN(
        n13922) );
  INV_X1 U25043 ( .A(n15380), .ZN(n15359) );
  NAND3_X1 U25044 ( .A1(n13917), .A2(n15359), .A3(n11853), .ZN(n13921) );
  INV_X1 U25045 ( .A(n13918), .ZN(n13919) );
  NAND2_X1 U25046 ( .A1(n13919), .A2(n15382), .ZN(n13920) );
  NAND4_X1 U25047 ( .A1(n13922), .A2(n13921), .A3(n13920), .A4(n15385), .ZN(
        n13927) );
  OAI21_X1 U25048 ( .B1(n15375), .B2(n14484), .A(n11853), .ZN(n13924) );
  NAND2_X1 U25049 ( .A1(n787), .A2(n15384), .ZN(n15357) );
  NAND2_X1 U25050 ( .A1(n13930), .A2(n51657), .ZN(n13931) );
  MUX2_X1 U25051 ( .A(n13932), .B(n13931), .S(n13947), .Z(n13939) );
  NAND3_X1 U25052 ( .A1(n13934), .A2(n6668), .A3(n13933), .ZN(n13936) );
  AND2_X1 U25053 ( .A1(n13936), .A2(n13935), .ZN(n13937) );
  INV_X1 U25054 ( .A(n13940), .ZN(n13943) );
  AOI22_X1 U25055 ( .A1(n13943), .A2(n13942), .B1(n13941), .B2(n13948), .ZN(
        n13954) );
  NAND4_X1 U25057 ( .A1(n13950), .A2(n13949), .A3(n13948), .A4(n13947), .ZN(
        n13951) );
  NAND4_X1 U25058 ( .A1(n13954), .A2(n13953), .A3(n13952), .A4(n13951), .ZN(
        n13955) );
  NOR2_X1 U25059 ( .A1(n13956), .A2(n13955), .ZN(n15154) );
  NAND2_X1 U25060 ( .A1(n14233), .A2(n13957), .ZN(n16220) );
  INV_X1 U25061 ( .A(n16220), .ZN(n13962) );
  NAND2_X1 U25062 ( .A1(n13970), .A2(n14228), .ZN(n13959) );
  AOI21_X1 U25063 ( .B1(n13960), .B2(n13959), .A(n13958), .ZN(n16219) );
  INV_X1 U25064 ( .A(n16219), .ZN(n13961) );
  NAND3_X1 U25065 ( .A1(n13962), .A2(n14234), .A3(n13961), .ZN(n15151) );
  INV_X1 U25066 ( .A(n13963), .ZN(n13964) );
  INV_X1 U25067 ( .A(n16223), .ZN(n15150) );
  NOR2_X1 U25068 ( .A1(n13969), .A2(n13968), .ZN(n13975) );
  INV_X1 U25069 ( .A(n14223), .ZN(n13974) );
  NOR2_X1 U25070 ( .A1(n13971), .A2(n13970), .ZN(n14231) );
  INV_X1 U25071 ( .A(n13972), .ZN(n13973) );
  OAI21_X1 U25074 ( .B1(n15151), .B2(n15150), .A(n836), .ZN(n15796) );
  XNOR2_X1 U25075 ( .A(n15154), .B(n15796), .ZN(n16158) );
  OAI211_X1 U25076 ( .C1(n13980), .C2(n13979), .A(n13978), .B(n13977), .ZN(
        n13981) );
  INV_X1 U25077 ( .A(n13981), .ZN(n13983) );
  NAND3_X1 U25078 ( .A1(n13984), .A2(n13983), .A3(n13982), .ZN(n13985) );
  XNOR2_X1 U25079 ( .A(n4909), .B(n4723), .ZN(n34575) );
  XNOR2_X1 U25080 ( .A(n34575), .B(n18636), .ZN(n46097) );
  XNOR2_X1 U25081 ( .A(n4353), .B(n3336), .ZN(n28307) );
  XNOR2_X1 U25082 ( .A(n46097), .B(n28307), .ZN(n15213) );
  XNOR2_X1 U25083 ( .A(n15213), .B(n2903), .ZN(n25145) );
  XNOR2_X1 U25084 ( .A(n43691), .B(n4121), .ZN(n33388) );
  XOR2_X1 U25085 ( .A(n4647), .B(n42668), .Z(n13986) );
  XNOR2_X1 U25086 ( .A(n33388), .B(n13986), .ZN(n13987) );
  XNOR2_X1 U25087 ( .A(n25145), .B(n13987), .ZN(n13988) );
  XNOR2_X1 U25088 ( .A(n15677), .B(n13988), .ZN(n13989) );
  XNOR2_X1 U25089 ( .A(n15511), .B(n13989), .ZN(n14017) );
  NAND3_X1 U25090 ( .A1(n13991), .A2(n13990), .A3(n13994), .ZN(n13992) );
  AND2_X1 U25091 ( .A1(n13993), .A2(n13992), .ZN(n13999) );
  NAND3_X1 U25092 ( .A1(n13996), .A2(n13995), .A3(n13994), .ZN(n13997) );
  NAND4_X1 U25093 ( .A1(n14000), .A2(n13999), .A3(n13998), .A4(n13997), .ZN(
        n18202) );
  XNOR2_X1 U25094 ( .A(n18202), .B(n16701), .ZN(n17368) );
  NAND2_X1 U25095 ( .A1(n14001), .A2(n14006), .ZN(n14002) );
  OAI21_X1 U25096 ( .B1(n14003), .B2(n14002), .A(n14172), .ZN(n14016) );
  NOR2_X1 U25097 ( .A1(n14006), .A2(n14600), .ZN(n14005) );
  AOI22_X1 U25098 ( .A1(n14597), .A2(n14005), .B1(n14004), .B2(n14601), .ZN(
        n14015) );
  INV_X1 U25099 ( .A(n14006), .ZN(n14610) );
  XNOR2_X1 U25100 ( .A(n14596), .B(n14170), .ZN(n14007) );
  OAI22_X1 U25101 ( .A1(n14010), .A2(n14009), .B1(n14008), .B2(n14170), .ZN(
        n14012) );
  NAND2_X1 U25102 ( .A1(n14012), .A2(n14011), .ZN(n14013) );
  XNOR2_X1 U25104 ( .A(n17938), .B(n17368), .ZN(n17816) );
  XNOR2_X1 U25105 ( .A(n17816), .B(n14017), .ZN(n14051) );
  INV_X1 U25106 ( .A(n14018), .ZN(n14020) );
  NAND2_X1 U25107 ( .A1(n14021), .A2(n14033), .ZN(n14027) );
  INV_X1 U25108 ( .A(n14025), .ZN(n14026) );
  OAI21_X1 U25109 ( .B1(n782), .B2(n6726), .A(n14028), .ZN(n14031) );
  AND2_X1 U25110 ( .A1(n14032), .A2(n14033), .ZN(n14037) );
  AOI22_X1 U25111 ( .A1(n14037), .A2(n14036), .B1(n14035), .B2(n14034), .ZN(
        n14039) );
  NAND3_X1 U25113 ( .A1(n15077), .A2(n1486), .A3(n15770), .ZN(n14042) );
  NAND2_X1 U25114 ( .A1(n14042), .A2(n14914), .ZN(n14044) );
  NAND4_X1 U25115 ( .A1(n15306), .A2(n15063), .A3(n15766), .A4(n2189), .ZN(
        n14043) );
  AND2_X1 U25116 ( .A1(n14044), .A2(n14043), .ZN(n15777) );
  NOR2_X1 U25117 ( .A1(n15068), .A2(n15073), .ZN(n14045) );
  AOI22_X1 U25118 ( .A1(n14045), .A2(n14929), .B1(n15067), .B2(n15769), .ZN(
        n14048) );
  AND2_X1 U25119 ( .A1(n2189), .A2(n15309), .ZN(n15062) );
  INV_X1 U25120 ( .A(n15062), .ZN(n15778) );
  AOI21_X1 U25121 ( .B1(n15766), .B2(n15770), .A(n15778), .ZN(n14046) );
  OAI21_X1 U25122 ( .B1(n15306), .B2(n15766), .A(n14046), .ZN(n14047) );
  XNOR2_X1 U25123 ( .A(n15300), .B(n14911), .ZN(n14912) );
  OAI211_X1 U25124 ( .C1(n14912), .C2(n2189), .A(n15307), .B(n15766), .ZN(
        n15773) );
  NAND4_X1 U25125 ( .A1(n15777), .A2(n14048), .A3(n14047), .A4(n15773), .ZN(
        n14049) );
  XNOR2_X2 U25126 ( .A(n18643), .B(n14049), .ZN(n17127) );
  XNOR2_X1 U25127 ( .A(n14050), .B(n17127), .ZN(n14569) );
  OAI211_X1 U25128 ( .C1(n51724), .C2(n14949), .A(n14957), .B(n14680), .ZN(
        n14056) );
  INV_X1 U25129 ( .A(n14052), .ZN(n14053) );
  NOR2_X1 U25130 ( .A1(n14053), .A2(n14956), .ZN(n14682) );
  INV_X1 U25131 ( .A(n14682), .ZN(n14055) );
  NAND3_X1 U25132 ( .A1(n14951), .A2(n51500), .A3(n14950), .ZN(n14054) );
  AOI21_X1 U25133 ( .B1(n14958), .B2(n14962), .A(n2151), .ZN(n14058) );
  OAI21_X1 U25134 ( .B1(n14059), .B2(n14957), .A(n14058), .ZN(n14062) );
  NAND2_X1 U25136 ( .A1(n14393), .A2(n14072), .ZN(n14067) );
  OAI22_X1 U25137 ( .A1(n14068), .A2(n14067), .B1(n14410), .B2(n14066), .ZN(
        n14069) );
  NOR2_X1 U25138 ( .A1(n14403), .A2(n14069), .ZN(n14078) );
  NOR2_X1 U25139 ( .A1(n14410), .A2(n14072), .ZN(n14395) );
  AOI22_X1 U25140 ( .A1(n14074), .A2(n14073), .B1(n14400), .B2(n14395), .ZN(
        n14076) );
  NAND3_X1 U25141 ( .A1(n14420), .A2(n14408), .A3(n14415), .ZN(n14075) );
  BUF_X2 U25142 ( .A(n14508), .Z(n17812) );
  XNOR2_X1 U25143 ( .A(n14079), .B(n17812), .ZN(n16535) );
  INV_X1 U25144 ( .A(n16535), .ZN(n14111) );
  OAI21_X1 U25145 ( .B1(n14721), .B2(n14720), .A(n14703), .ZN(n14081) );
  OAI211_X1 U25146 ( .C1(n14082), .C2(n14205), .A(n14081), .B(n14080), .ZN(
        n14083) );
  NAND2_X1 U25147 ( .A1(n14083), .A2(n14719), .ZN(n14093) );
  INV_X1 U25148 ( .A(n14084), .ZN(n14087) );
  INV_X1 U25149 ( .A(n14085), .ZN(n14086) );
  OAI22_X1 U25150 ( .A1(n14087), .A2(n14197), .B1(n14086), .B2(n14712), .ZN(
        n14091) );
  NOR2_X1 U25151 ( .A1(n14717), .A2(n14720), .ZN(n14710) );
  AOI21_X1 U25152 ( .B1(n14200), .B2(n14088), .A(n14704), .ZN(n14089) );
  AOI22_X1 U25153 ( .A1(n14713), .A2(n14091), .B1(n14090), .B2(n14089), .ZN(
        n14092) );
  AND2_X1 U25154 ( .A1(n14107), .A2(n14455), .ZN(n14446) );
  AND2_X1 U25155 ( .A1(n14103), .A2(n14455), .ZN(n14105) );
  INV_X1 U25156 ( .A(n17364), .ZN(n16237) );
  XNOR2_X1 U25157 ( .A(n16237), .B(n17365), .ZN(n14110) );
  XNOR2_X1 U25158 ( .A(n14111), .B(n14110), .ZN(n15607) );
  INV_X1 U25159 ( .A(n15607), .ZN(n14113) );
  XNOR2_X1 U25160 ( .A(n17125), .B(n43293), .ZN(n15682) );
  INV_X1 U25161 ( .A(n14114), .ZN(n14116) );
  NAND3_X1 U25162 ( .A1(n15235), .A2(n15233), .A3(n15196), .ZN(n14119) );
  NAND2_X1 U25163 ( .A1(n14117), .A2(n15196), .ZN(n14118) );
  NAND2_X1 U25164 ( .A1(n15235), .A2(n14120), .ZN(n14121) );
  NAND2_X1 U25165 ( .A1(n14574), .A2(n15177), .ZN(n15172) );
  INV_X1 U25166 ( .A(n15172), .ZN(n14127) );
  NOR2_X1 U25167 ( .A1(n15161), .A2(n51370), .ZN(n14126) );
  NAND2_X1 U25168 ( .A1(n15167), .A2(n15173), .ZN(n15176) );
  INV_X1 U25169 ( .A(n15176), .ZN(n14130) );
  INV_X1 U25170 ( .A(n14128), .ZN(n14129) );
  OAI21_X1 U25171 ( .B1(n14130), .B2(n14129), .A(n15168), .ZN(n14131) );
  INV_X1 U25172 ( .A(n18697), .ZN(n15743) );
  NAND2_X1 U25173 ( .A1(n14134), .A2(n15254), .ZN(n14136) );
  NAND2_X1 U25174 ( .A1(n15264), .A2(n15256), .ZN(n14135) );
  NAND2_X1 U25175 ( .A1(n14137), .A2(n15250), .ZN(n14138) );
  OAI21_X1 U25176 ( .B1(n15259), .B2(n14138), .A(n15257), .ZN(n14140) );
  INV_X1 U25177 ( .A(n14141), .ZN(n14142) );
  NAND3_X1 U25178 ( .A1(n14143), .A2(n15256), .A3(n14142), .ZN(n14144) );
  XNOR2_X1 U25179 ( .A(n15743), .B(n16431), .ZN(n18488) );
  OAI21_X1 U25180 ( .B1(n14150), .B2(n14966), .A(n14145), .ZN(n14148) );
  INV_X1 U25181 ( .A(n14146), .ZN(n14147) );
  NAND2_X1 U25182 ( .A1(n14148), .A2(n14147), .ZN(n14153) );
  NAND2_X1 U25183 ( .A1(n14150), .A2(n14149), .ZN(n14151) );
  AND3_X1 U25184 ( .A1(n14153), .A2(n14152), .A3(n14151), .ZN(n14970) );
  INV_X1 U25185 ( .A(n14154), .ZN(n14163) );
  OAI21_X1 U25186 ( .B1(n14160), .B2(n14966), .A(n14159), .ZN(n14968) );
  OAI211_X1 U25188 ( .C1(n14164), .C2(n14163), .A(n14162), .B(n51170), .ZN(
        n14165) );
  NAND2_X1 U25189 ( .A1(n14970), .A2(n14165), .ZN(n14176) );
  NAND3_X1 U25190 ( .A1(n14166), .A2(n14600), .A3(n14605), .ZN(n14168) );
  NAND2_X1 U25191 ( .A1(n14167), .A2(n14605), .ZN(n14599) );
  OAI211_X1 U25192 ( .C1(n14169), .C2(n14607), .A(n14168), .B(n14599), .ZN(
        n14174) );
  OAI211_X1 U25193 ( .C1(n14175), .C2(n14595), .A(n14174), .B(n14173), .ZN(
        n16943) );
  INV_X1 U25194 ( .A(n14177), .ZN(n14180) );
  NAND3_X1 U25195 ( .A1(n14180), .A2(n14179), .A3(n14178), .ZN(n14182) );
  NAND3_X1 U25196 ( .A1(n14188), .A2(n14187), .A3(n14186), .ZN(n14196) );
  INV_X1 U25197 ( .A(n14189), .ZN(n14195) );
  INV_X1 U25198 ( .A(n14190), .ZN(n14192) );
  OAI21_X1 U25199 ( .B1(n14193), .B2(n14192), .A(n14191), .ZN(n14194) );
  XNOR2_X1 U25200 ( .A(n17731), .B(n17730), .ZN(n18479) );
  XNOR2_X1 U25201 ( .A(n18479), .B(n566), .ZN(n15744) );
  XNOR2_X1 U25202 ( .A(n16571), .B(n17954), .ZN(n16183) );
  NAND2_X1 U25203 ( .A1(n14198), .A2(n14197), .ZN(n14201) );
  AOI21_X1 U25204 ( .B1(n14201), .B2(n14200), .A(n14199), .ZN(n14207) );
  OAI21_X1 U25205 ( .B1(n14724), .B2(n14721), .A(n14202), .ZN(n14204) );
  NAND2_X1 U25206 ( .A1(n14717), .A2(n14711), .ZN(n14203) );
  INV_X1 U25207 ( .A(n17281), .ZN(n16346) );
  XNOR2_X1 U25208 ( .A(n16346), .B(n5016), .ZN(n17948) );
  XNOR2_X1 U25209 ( .A(n17948), .B(n16183), .ZN(n14211) );
  XNOR2_X1 U25210 ( .A(n16435), .B(n48814), .ZN(n17275) );
  XNOR2_X1 U25211 ( .A(n24992), .B(n44483), .ZN(n41460) );
  INV_X1 U25212 ( .A(n28085), .ZN(n14208) );
  XNOR2_X1 U25213 ( .A(n41460), .B(n14208), .ZN(n23581) );
  XNOR2_X1 U25214 ( .A(Key[88]), .B(n4803), .ZN(n43764) );
  XNOR2_X1 U25215 ( .A(n4237), .B(n4864), .ZN(n40104) );
  XNOR2_X1 U25216 ( .A(n43764), .B(n40104), .ZN(n17181) );
  XNOR2_X1 U25217 ( .A(n4471), .B(n4845), .ZN(n28084) );
  XNOR2_X1 U25218 ( .A(n17181), .B(n28084), .ZN(n26162) );
  XNOR2_X1 U25219 ( .A(n23581), .B(n26162), .ZN(n35520) );
  XNOR2_X1 U25220 ( .A(n42889), .B(n2601), .ZN(n27299) );
  XNOR2_X1 U25221 ( .A(n27299), .B(n4026), .ZN(n35353) );
  XNOR2_X1 U25222 ( .A(n35520), .B(n35353), .ZN(n14209) );
  XNOR2_X1 U25223 ( .A(n17275), .B(n14209), .ZN(n14210) );
  XNOR2_X1 U25224 ( .A(n14211), .B(n14210), .ZN(n14212) );
  NAND2_X1 U25225 ( .A1(n18342), .A2(n18331), .ZN(n14383) );
  NAND2_X1 U25226 ( .A1(n16834), .A2(n18063), .ZN(n17436) );
  XNOR2_X1 U25227 ( .A(n19260), .B(n15883), .ZN(n14216) );
  XNOR2_X1 U25228 ( .A(n4926), .B(n4836), .ZN(n24797) );
  XNOR2_X1 U25229 ( .A(Key[85]), .B(n4691), .ZN(n23882) );
  XNOR2_X1 U25230 ( .A(n24797), .B(n23882), .ZN(n45350) );
  XNOR2_X1 U25231 ( .A(n2231), .B(n4916), .ZN(n36941) );
  XNOR2_X1 U25232 ( .A(n45350), .B(n36941), .ZN(n25374) );
  XNOR2_X1 U25233 ( .A(n25374), .B(n4838), .ZN(n19262) );
  INV_X1 U25234 ( .A(n19262), .ZN(n25281) );
  XNOR2_X1 U25235 ( .A(n4855), .B(n4247), .ZN(n45348) );
  XNOR2_X1 U25236 ( .A(n4788), .B(n4930), .ZN(n43727) );
  XNOR2_X1 U25237 ( .A(n45348), .B(n43727), .ZN(n26025) );
  XNOR2_X1 U25238 ( .A(n25281), .B(n26025), .ZN(n34818) );
  XNOR2_X1 U25239 ( .A(n42327), .B(n4869), .ZN(n14214) );
  XNOR2_X1 U25240 ( .A(n34818), .B(n14214), .ZN(n14215) );
  XNOR2_X1 U25241 ( .A(n14216), .B(n14215), .ZN(n14217) );
  XNOR2_X1 U25242 ( .A(n16064), .B(n17972), .ZN(n18460) );
  XNOR2_X1 U25243 ( .A(n14217), .B(n18460), .ZN(n14219) );
  XNOR2_X1 U25244 ( .A(n4712), .B(n4782), .ZN(n25616) );
  XNOR2_X1 U25245 ( .A(n26178), .B(n25616), .ZN(n44495) );
  INV_X1 U25246 ( .A(n44495), .ZN(n35035) );
  XNOR2_X1 U25247 ( .A(n15454), .B(n35035), .ZN(n14218) );
  XNOR2_X1 U25248 ( .A(n15876), .B(n14218), .ZN(n18706) );
  XNOR2_X1 U25249 ( .A(n18706), .B(n14219), .ZN(n14241) );
  XNOR2_X1 U25250 ( .A(n8699), .B(n45736), .ZN(n14238) );
  NAND3_X1 U25251 ( .A1(n14221), .A2(n16221), .A3(n14220), .ZN(n14222) );
  AND2_X1 U25252 ( .A1(n14234), .A2(n14224), .ZN(n14225) );
  AOI22_X1 U25253 ( .A1(n14231), .A2(n14227), .B1(n14226), .B2(n14225), .ZN(
        n14236) );
  MUX2_X1 U25254 ( .A(n14230), .B(n14229), .S(n14228), .Z(n14235) );
  XNOR2_X1 U25255 ( .A(n14238), .B(n17973), .ZN(n16384) );
  INV_X1 U25256 ( .A(n14239), .ZN(n15738) );
  XNOR2_X1 U25257 ( .A(n16384), .B(n15409), .ZN(n14240) );
  XNOR2_X1 U25258 ( .A(n14241), .B(n14240), .ZN(n14378) );
  INV_X1 U25259 ( .A(n14242), .ZN(n14246) );
  AOI21_X1 U25260 ( .B1(n15106), .B2(n14246), .A(n14245), .ZN(n14249) );
  OAI22_X1 U25261 ( .A1(n14247), .A2(n15117), .B1(n15108), .B2(n14976), .ZN(
        n14248) );
  NOR2_X1 U25262 ( .A1(n14249), .A2(n14248), .ZN(n14255) );
  NAND2_X1 U25263 ( .A1(n14250), .A2(n15103), .ZN(n14254) );
  MUX2_X1 U25264 ( .A(n14252), .B(n15113), .S(n14251), .Z(n14975) );
  NAND3_X1 U25265 ( .A1(n14975), .A2(n14974), .A3(n15118), .ZN(n14253) );
  NAND2_X1 U25266 ( .A1(n14998), .A2(n14999), .ZN(n14259) );
  NAND3_X1 U25267 ( .A1(n15133), .A2(n15126), .A3(n14257), .ZN(n14258) );
  MUX2_X1 U25268 ( .A(n14259), .B(n14258), .S(n15136), .Z(n14266) );
  INV_X1 U25269 ( .A(n15133), .ZN(n14261) );
  NOR2_X1 U25270 ( .A1(n14261), .A2(n14260), .ZN(n15127) );
  INV_X1 U25271 ( .A(n15127), .ZN(n14265) );
  NAND3_X1 U25272 ( .A1(n14262), .A2(n15138), .A3(n14270), .ZN(n14263) );
  NAND4_X1 U25273 ( .A1(n14266), .A2(n14265), .A3(n14264), .A4(n14263), .ZN(
        n14275) );
  INV_X1 U25274 ( .A(n15131), .ZN(n14269) );
  OAI211_X1 U25275 ( .C1(n14272), .C2(n15133), .A(n14271), .B(n14994), .ZN(
        n14273) );
  OAI21_X1 U25276 ( .B1(n14278), .B2(n14277), .A(n14276), .ZN(n14283) );
  INV_X1 U25277 ( .A(n14279), .ZN(n14281) );
  NAND3_X1 U25278 ( .A1(n14281), .A2(n14280), .A3(n14287), .ZN(n14282) );
  NAND2_X1 U25279 ( .A1(n14283), .A2(n14282), .ZN(n14302) );
  AOI21_X1 U25280 ( .B1(n14286), .B2(n14285), .A(n14284), .ZN(n14293) );
  OAI21_X1 U25281 ( .B1(n14289), .B2(n14288), .A(n14287), .ZN(n14292) );
  AOI22_X1 U25282 ( .A1(n14293), .A2(n14292), .B1(n14291), .B2(n14290), .ZN(
        n14301) );
  INV_X1 U25285 ( .A(n14303), .ZN(n14305) );
  INV_X1 U25286 ( .A(n14312), .ZN(n14304) );
  INV_X1 U25287 ( .A(n14306), .ZN(n14309) );
  OAI21_X1 U25288 ( .B1(n14309), .B2(n14308), .A(n14307), .ZN(n14327) );
  INV_X1 U25289 ( .A(n14319), .ZN(n14316) );
  NAND2_X1 U25290 ( .A1(n14312), .A2(n14311), .ZN(n14313) );
  OAI211_X1 U25291 ( .C1(n14316), .C2(n14315), .A(n14314), .B(n14313), .ZN(
        n14325) );
  NAND4_X1 U25292 ( .A1(n14319), .A2(n14321), .A3(n14318), .A4(n14317), .ZN(
        n14323) );
  NOR2_X1 U25293 ( .A1(n14325), .A2(n14324), .ZN(n14326) );
  XNOR2_X1 U25294 ( .A(n18592), .B(n17378), .ZN(n14377) );
  NAND2_X1 U25295 ( .A1(n14353), .A2(n14330), .ZN(n14332) );
  NAND2_X1 U25296 ( .A1(n14332), .A2(n14331), .ZN(n14335) );
  INV_X1 U25297 ( .A(n14333), .ZN(n14334) );
  NAND2_X1 U25298 ( .A1(n14335), .A2(n14334), .ZN(n14356) );
  NAND2_X1 U25299 ( .A1(n14340), .A2(n14339), .ZN(n14349) );
  NAND3_X1 U25300 ( .A1(n14343), .A2(n14342), .A3(n14341), .ZN(n14348) );
  NAND3_X1 U25301 ( .A1(n14346), .A2(n14345), .A3(n14344), .ZN(n14347) );
  NAND4_X1 U25302 ( .A1(n14350), .A2(n14349), .A3(n14348), .A4(n14347), .ZN(
        n14355) );
  OAI21_X1 U25303 ( .B1(n14353), .B2(n14352), .A(n14351), .ZN(n14354) );
  INV_X1 U25304 ( .A(n14358), .ZN(n14361) );
  NAND3_X1 U25305 ( .A1(n14359), .A2(n14552), .A3(n14369), .ZN(n14360) );
  OAI21_X1 U25306 ( .B1(n14361), .B2(n14552), .A(n14360), .ZN(n14376) );
  NAND3_X1 U25307 ( .A1(n14363), .A2(n6070), .A3(n14368), .ZN(n14364) );
  OAI21_X1 U25308 ( .B1(n14540), .B2(n14550), .A(n14366), .ZN(n14374) );
  OAI22_X1 U25309 ( .A1(n14368), .A2(n6070), .B1(n14367), .B2(n14534), .ZN(
        n14372) );
  INV_X1 U25310 ( .A(n14369), .ZN(n14371) );
  OAI21_X1 U25311 ( .B1(n14372), .B2(n14371), .A(n14370), .ZN(n14373) );
  NAND3_X1 U25312 ( .A1(n18330), .A2(n18071), .A3(n18064), .ZN(n18066) );
  NAND2_X1 U25315 ( .A1(n18059), .A2(n17545), .ZN(n14382) );
  AOI21_X1 U25316 ( .B1(n14383), .B2(n14382), .A(n17542), .ZN(n14384) );
  OR2_X1 U25317 ( .A1(n14384), .A2(n18336), .ZN(n14391) );
  INV_X1 U25319 ( .A(n18059), .ZN(n17431) );
  NAND3_X1 U25320 ( .A1(n17431), .A2(n18331), .A3(n18071), .ZN(n14388) );
  NAND4_X1 U25321 ( .A1(n18342), .A2(n18059), .A3(n403), .A4(n17553), .ZN(
        n14387) );
  INV_X1 U25322 ( .A(n17436), .ZN(n18074) );
  NAND4_X1 U25323 ( .A1(n18074), .A2(n17546), .A3(n18331), .A4(n772), .ZN(
        n18338) );
  INV_X1 U25324 ( .A(n22285), .ZN(n22697) );
  NAND2_X1 U25327 ( .A1(n14396), .A2(n14395), .ZN(n14402) );
  INV_X1 U25328 ( .A(n14397), .ZN(n14399) );
  NAND2_X1 U25329 ( .A1(n14399), .A2(n14398), .ZN(n14401) );
  MUX2_X1 U25330 ( .A(n14402), .B(n14401), .S(n14400), .Z(n14426) );
  INV_X1 U25331 ( .A(n14403), .ZN(n14404) );
  AND3_X1 U25332 ( .A1(n14406), .A2(n14405), .A3(n14404), .ZN(n14425) );
  INV_X1 U25333 ( .A(n14407), .ZN(n14409) );
  OAI21_X1 U25334 ( .B1(n14409), .B2(n14408), .A(n14410), .ZN(n14414) );
  NAND3_X1 U25335 ( .A1(n14417), .A2(n14411), .A3(n14410), .ZN(n14413) );
  MUX2_X1 U25336 ( .A(n14414), .B(n14413), .S(n14412), .Z(n14424) );
  INV_X1 U25337 ( .A(n14415), .ZN(n14416) );
  OAI22_X1 U25338 ( .A1(n14419), .A2(n14418), .B1(n14417), .B2(n14416), .ZN(
        n14422) );
  INV_X1 U25339 ( .A(n14420), .ZN(n14421) );
  NAND2_X1 U25340 ( .A1(n14422), .A2(n14421), .ZN(n14423) );
  XNOR2_X1 U25342 ( .A(n17758), .B(n19196), .ZN(n17697) );
  XNOR2_X1 U25343 ( .A(n14427), .B(n18399), .ZN(n14428) );
  XNOR2_X1 U25344 ( .A(n17697), .B(n14428), .ZN(n14466) );
  XNOR2_X1 U25345 ( .A(n4666), .B(n3367), .ZN(n41825) );
  XNOR2_X1 U25346 ( .A(n41825), .B(n4431), .ZN(n36737) );
  XNOR2_X1 U25347 ( .A(Key[75]), .B(n4637), .ZN(n42630) );
  XNOR2_X1 U25348 ( .A(n36737), .B(n2599), .ZN(n14429) );
  XNOR2_X1 U25349 ( .A(n14429), .B(n37138), .ZN(n14430) );
  XNOR2_X1 U25350 ( .A(n2117), .B(n4937), .ZN(n33930) );
  XNOR2_X1 U25351 ( .A(n33930), .B(n4739), .ZN(n25134) );
  XNOR2_X1 U25352 ( .A(n25134), .B(n4554), .ZN(n33136) );
  XNOR2_X1 U25353 ( .A(n14430), .B(n33136), .ZN(n14431) );
  XNOR2_X1 U25354 ( .A(n41183), .B(n4638), .ZN(n37013) );
  XNOR2_X1 U25355 ( .A(n14431), .B(n37013), .ZN(n14432) );
  XNOR2_X1 U25356 ( .A(n17764), .B(n14432), .ZN(n14464) );
  INV_X1 U25357 ( .A(n14433), .ZN(n14435) );
  NAND2_X1 U25358 ( .A1(n14435), .A2(n14434), .ZN(n14437) );
  NAND2_X1 U25359 ( .A1(n14455), .A2(n640), .ZN(n14440) );
  OAI21_X1 U25361 ( .B1(n14445), .B2(n14444), .A(n14443), .ZN(n14447) );
  XOR2_X1 U25362 ( .A(n640), .B(n14454), .Z(n14457) );
  AOI21_X1 U25363 ( .B1(n14455), .B2(n14454), .A(n14453), .ZN(n14456) );
  NAND3_X1 U25364 ( .A1(n14458), .A2(n14457), .A3(n14456), .ZN(n14459) );
  XNOR2_X1 U25365 ( .A(n17707), .B(n17763), .ZN(n14463) );
  XNOR2_X1 U25366 ( .A(n14464), .B(n14463), .ZN(n14465) );
  XNOR2_X1 U25367 ( .A(n14466), .B(n14465), .ZN(n14467) );
  XNOR2_X1 U25368 ( .A(n19210), .B(n14467), .ZN(n14470) );
  XNOR2_X1 U25369 ( .A(n16498), .B(n16628), .ZN(n15563) );
  XNOR2_X1 U25370 ( .A(n15563), .B(n52190), .ZN(n14468) );
  XNOR2_X1 U25371 ( .A(n15824), .B(n14468), .ZN(n14469) );
  MUX2_X1 U25372 ( .A(n14472), .B(n14471), .S(n14480), .Z(n14483) );
  NOR2_X1 U25373 ( .A1(n14474), .A2(n14473), .ZN(n14475) );
  AOI21_X1 U25374 ( .B1(n14477), .B2(n14476), .A(n14475), .ZN(n14887) );
  NAND3_X1 U25375 ( .A1(n14480), .A2(n14479), .A3(n14478), .ZN(n14481) );
  NAND2_X1 U25376 ( .A1(n15374), .A2(n15384), .ZN(n14494) );
  XNOR2_X1 U25377 ( .A(n18169), .B(n2162), .ZN(n14497) );
  XNOR2_X1 U25378 ( .A(n14497), .B(n511), .ZN(n14498) );
  XNOR2_X1 U25379 ( .A(n27483), .B(n29662), .ZN(n24229) );
  XNOR2_X1 U25380 ( .A(n24229), .B(n2605), .ZN(n34893) );
  XNOR2_X1 U25381 ( .A(n25040), .B(n41567), .ZN(n17149) );
  XNOR2_X1 U25382 ( .A(n34893), .B(n17149), .ZN(n38860) );
  INV_X1 U25383 ( .A(n42769), .ZN(n49887) );
  XNOR2_X1 U25384 ( .A(n24894), .B(n49887), .ZN(n17773) );
  INV_X1 U25385 ( .A(n17773), .ZN(n29664) );
  XNOR2_X1 U25386 ( .A(n274), .B(n1326), .ZN(n34614) );
  XNOR2_X1 U25387 ( .A(n34614), .B(n842), .ZN(n14499) );
  XNOR2_X1 U25388 ( .A(n29664), .B(n14499), .ZN(n14500) );
  XNOR2_X1 U25389 ( .A(n38860), .B(n14500), .ZN(n14501) );
  XNOR2_X1 U25390 ( .A(n18539), .B(n14501), .ZN(n14502) );
  XNOR2_X1 U25391 ( .A(n17208), .B(n14502), .ZN(n14504) );
  XNOR2_X1 U25392 ( .A(n4035), .B(Key[156]), .ZN(n25042) );
  XNOR2_X1 U25393 ( .A(n25042), .B(n4651), .ZN(n46062) );
  XNOR2_X1 U25394 ( .A(n51758), .B(n46062), .ZN(n14503) );
  XNOR2_X1 U25395 ( .A(n14503), .B(n15957), .ZN(n15582) );
  XNOR2_X1 U25396 ( .A(n14504), .B(n15582), .ZN(n14505) );
  XNOR2_X1 U25397 ( .A(n15579), .B(n16337), .ZN(n14507) );
  XNOR2_X1 U25398 ( .A(n14506), .B(n14507), .ZN(n16250) );
  XNOR2_X1 U25399 ( .A(n17364), .B(n43702), .ZN(n14509) );
  XNOR2_X1 U25400 ( .A(n14511), .B(n14510), .ZN(n14559) );
  AND2_X1 U25401 ( .A1(n51019), .A2(n14512), .ZN(n14513) );
  NAND2_X1 U25402 ( .A1(n14514), .A2(n14513), .ZN(n16034) );
  OR2_X1 U25403 ( .A1(n14516), .A2(n14515), .ZN(n16046) );
  AND2_X1 U25404 ( .A1(n16034), .A2(n16046), .ZN(n14532) );
  NAND2_X1 U25405 ( .A1(n14519), .A2(n16049), .ZN(n14517) );
  OAI21_X1 U25406 ( .B1(n16045), .B2(n14517), .A(n16043), .ZN(n14518) );
  AND2_X1 U25407 ( .A1(n16035), .A2(n14518), .ZN(n14531) );
  NAND3_X1 U25408 ( .A1(n14521), .A2(n14520), .A3(n14519), .ZN(n14524) );
  NAND3_X1 U25409 ( .A1(n16044), .A2(n14522), .A3(n51018), .ZN(n14523) );
  AND2_X1 U25410 ( .A1(n14524), .A2(n14523), .ZN(n16051) );
  NAND3_X1 U25411 ( .A1(n14525), .A2(n16049), .A3(n51019), .ZN(n14526) );
  NAND4_X1 U25412 ( .A1(n14529), .A2(n14528), .A3(n14527), .A4(n14526), .ZN(
        n14530) );
  NAND4_X1 U25413 ( .A1(n14532), .A2(n14531), .A3(n16051), .A4(n14530), .ZN(
        n14558) );
  NAND3_X1 U25414 ( .A1(n14537), .A2(n14536), .A3(n14544), .ZN(n14538) );
  AND2_X1 U25415 ( .A1(n14539), .A2(n14538), .ZN(n14557) );
  OAI211_X1 U25416 ( .C1(n14543), .C2(n14542), .A(n14541), .B(n14540), .ZN(
        n14556) );
  OAI21_X1 U25417 ( .B1(n14545), .B2(n14553), .A(n14544), .ZN(n14546) );
  NAND2_X1 U25418 ( .A1(n14549), .A2(n14548), .ZN(n14555) );
  OAI211_X1 U25419 ( .C1(n14553), .C2(n14552), .A(n14551), .B(n14550), .ZN(
        n14554) );
  XNOR2_X1 U25420 ( .A(n16464), .B(n14558), .ZN(n15680) );
  XNOR2_X1 U25421 ( .A(n15680), .B(n17804), .ZN(n15517) );
  XNOR2_X1 U25422 ( .A(n14559), .B(n15517), .ZN(n17115) );
  XNOR2_X1 U25423 ( .A(n25145), .B(n4650), .ZN(n26386) );
  XNOR2_X1 U25424 ( .A(n4641), .B(n4886), .ZN(n43662) );
  XNOR2_X1 U25425 ( .A(n26386), .B(n43662), .ZN(n34440) );
  XNOR2_X1 U25426 ( .A(n18791), .B(n34440), .ZN(n14560) );
  XNOR2_X1 U25427 ( .A(n18644), .B(n14560), .ZN(n14568) );
  INV_X1 U25428 ( .A(Key[152]), .ZN(n50431) );
  XNOR2_X1 U25429 ( .A(n50431), .B(n4746), .ZN(n42077) );
  INV_X1 U25430 ( .A(n42077), .ZN(n42995) );
  XNOR2_X1 U25431 ( .A(n42995), .B(n4558), .ZN(n28304) );
  XNOR2_X1 U25432 ( .A(n28304), .B(n48597), .ZN(n27175) );
  XNOR2_X1 U25433 ( .A(n4647), .B(n4568), .ZN(n25925) );
  XNOR2_X1 U25434 ( .A(n27175), .B(n25925), .ZN(n33519) );
  XNOR2_X1 U25435 ( .A(n17936), .B(n33519), .ZN(n14566) );
  OAI21_X1 U25436 ( .B1(n14562), .B2(n14561), .A(n2114), .ZN(n14565) );
  XNOR2_X1 U25437 ( .A(n17643), .B(n17118), .ZN(n15678) );
  XNOR2_X1 U25438 ( .A(n14566), .B(n15678), .ZN(n14567) );
  XNOR2_X1 U25439 ( .A(n14568), .B(n14567), .ZN(n14570) );
  XNOR2_X1 U25440 ( .A(n14569), .B(n14570), .ZN(n14571) );
  XNOR2_X1 U25441 ( .A(n17115), .B(n14571), .ZN(n14738) );
  NAND3_X1 U25442 ( .A1(n14575), .A2(n14574), .A3(n15161), .ZN(n14576) );
  INV_X1 U25443 ( .A(n14577), .ZN(n14578) );
  NAND2_X1 U25444 ( .A1(n14579), .A2(n15161), .ZN(n14580) );
  OAI21_X1 U25445 ( .B1(n15167), .B2(n15177), .A(n15163), .ZN(n14582) );
  NAND2_X1 U25446 ( .A1(n15159), .A2(n14582), .ZN(n14583) );
  INV_X1 U25447 ( .A(n15519), .ZN(n14584) );
  XNOR2_X1 U25448 ( .A(n16158), .B(n14584), .ZN(n14586) );
  XNOR2_X1 U25449 ( .A(n14585), .B(n14586), .ZN(n19243) );
  INV_X1 U25450 ( .A(n19243), .ZN(n14625) );
  XNOR2_X1 U25451 ( .A(n17665), .B(n18447), .ZN(n14587) );
  XNOR2_X1 U25452 ( .A(n14587), .B(n15913), .ZN(n18630) );
  XNOR2_X1 U25453 ( .A(n24861), .B(n4537), .ZN(n45403) );
  XNOR2_X1 U25454 ( .A(n45403), .B(n4618), .ZN(n26403) );
  XNOR2_X1 U25455 ( .A(n26403), .B(n27353), .ZN(n33361) );
  XNOR2_X1 U25456 ( .A(n33361), .B(n4177), .ZN(n14590) );
  BUF_X1 U25457 ( .A(Key[47]), .Z(n46552) );
  XNOR2_X1 U25458 ( .A(n2603), .B(n46552), .ZN(n14588) );
  XNOR2_X1 U25459 ( .A(n14588), .B(n32856), .ZN(n33611) );
  XNOR2_X1 U25460 ( .A(n33611), .B(n49937), .ZN(n14589) );
  XNOR2_X1 U25461 ( .A(n25897), .B(n23943), .ZN(n22776) );
  XNOR2_X1 U25462 ( .A(n14589), .B(n22776), .ZN(n34095) );
  XNOR2_X1 U25463 ( .A(n14590), .B(n34095), .ZN(n14591) );
  XNOR2_X1 U25464 ( .A(n18432), .B(n17923), .ZN(n14592) );
  XNOR2_X1 U25465 ( .A(n14593), .B(n14592), .ZN(n14594) );
  XNOR2_X1 U25466 ( .A(n18630), .B(n14594), .ZN(n14624) );
  NAND2_X1 U25467 ( .A1(n14599), .A2(n14601), .ZN(n14598) );
  NOR2_X1 U25468 ( .A1(n14601), .A2(n14600), .ZN(n14604) );
  AOI21_X1 U25469 ( .B1(n14604), .B2(n14603), .A(n14602), .ZN(n14615) );
  NOR2_X1 U25470 ( .A1(n14606), .A2(n14605), .ZN(n14608) );
  OAI21_X1 U25471 ( .B1(n14609), .B2(n14608), .A(n14607), .ZN(n14614) );
  NAND3_X1 U25472 ( .A1(n14612), .A2(n14611), .A3(n14610), .ZN(n14613) );
  XNOR2_X1 U25473 ( .A(n16450), .B(n16923), .ZN(n14616) );
  XNOR2_X1 U25474 ( .A(n16913), .B(n14616), .ZN(n14622) );
  AOI21_X1 U25475 ( .B1(n51347), .B2(n14618), .A(n14617), .ZN(n14620) );
  INV_X1 U25476 ( .A(n2200), .ZN(n16924) );
  XNOR2_X1 U25477 ( .A(n17925), .B(n16924), .ZN(n14621) );
  XNOR2_X1 U25478 ( .A(n14622), .B(n14621), .ZN(n14623) );
  XNOR2_X1 U25479 ( .A(n17947), .B(n18689), .ZN(n15972) );
  XNOR2_X1 U25480 ( .A(n17181), .B(n4676), .ZN(n45335) );
  XNOR2_X1 U25481 ( .A(n23581), .B(n45335), .ZN(n41782) );
  XNOR2_X1 U25482 ( .A(n4613), .B(n4599), .ZN(n15964) );
  XNOR2_X1 U25483 ( .A(n4733), .B(n4048), .ZN(n17182) );
  XNOR2_X1 U25484 ( .A(n15964), .B(n17182), .ZN(n37058) );
  XNOR2_X1 U25485 ( .A(n41782), .B(n37058), .ZN(n14626) );
  XNOR2_X1 U25486 ( .A(n17389), .B(n14626), .ZN(n14627) );
  XNOR2_X1 U25487 ( .A(n17954), .B(n14627), .ZN(n14628) );
  XNOR2_X1 U25488 ( .A(n15972), .B(n14628), .ZN(n14630) );
  XNOR2_X1 U25489 ( .A(n51703), .B(n4737), .ZN(n14629) );
  XNOR2_X1 U25490 ( .A(n14629), .B(n18827), .ZN(n16079) );
  XNOR2_X1 U25491 ( .A(n14630), .B(n16079), .ZN(n14678) );
  OAI21_X1 U25492 ( .B1(n14644), .B2(n14636), .A(n14635), .ZN(n14638) );
  NAND2_X1 U25493 ( .A1(n14638), .A2(n14637), .ZN(n14648) );
  OAI21_X1 U25495 ( .B1(n14642), .B2(n14641), .A(n14640), .ZN(n14645) );
  NAND3_X1 U25496 ( .A1(n14645), .A2(n14644), .A3(n2114), .ZN(n14646) );
  INV_X1 U25497 ( .A(n18475), .ZN(n14662) );
  INV_X1 U25498 ( .A(n14650), .ZN(n14661) );
  INV_X1 U25499 ( .A(n14651), .ZN(n14654) );
  INV_X1 U25500 ( .A(n14652), .ZN(n14653) );
  NAND2_X1 U25501 ( .A1(n14654), .A2(n14653), .ZN(n14659) );
  OAI21_X1 U25502 ( .B1(n14657), .B2(n14656), .A(n14655), .ZN(n14658) );
  NAND4_X1 U25503 ( .A1(n14661), .A2(n14660), .A3(n14659), .A4(n14658), .ZN(
        n17960) );
  OAI21_X1 U25504 ( .B1(n51347), .B2(n14664), .A(n14663), .ZN(n14669) );
  NAND3_X1 U25505 ( .A1(n14674), .A2(n14666), .A3(n783), .ZN(n14668) );
  NAND2_X1 U25506 ( .A1(n14671), .A2(n14670), .ZN(n14676) );
  OAI21_X1 U25507 ( .B1(n14674), .B2(n14673), .A(n14672), .ZN(n14675) );
  XNOR2_X2 U25508 ( .A(n4486), .B(n4471), .ZN(n43586) );
  XNOR2_X1 U25509 ( .A(n43586), .B(n4654), .ZN(n43878) );
  XNOR2_X1 U25510 ( .A(n18119), .B(n43878), .ZN(n15295) );
  XNOR2_X1 U25511 ( .A(n14678), .B(n14677), .ZN(n14679) );
  NAND2_X1 U25513 ( .A1(n14680), .A2(n2151), .ZN(n14684) );
  NOR2_X1 U25514 ( .A1(n14959), .A2(n14938), .ZN(n14683) );
  AOI22_X1 U25516 ( .A1(n14684), .A2(n14683), .B1(n14682), .B2(n15283), .ZN(
        n14697) );
  NAND3_X1 U25517 ( .A1(n14952), .A2(n2151), .A3(n15278), .ZN(n14685) );
  NAND2_X1 U25518 ( .A1(n14686), .A2(n14685), .ZN(n14696) );
  OAI21_X1 U25519 ( .B1(n15273), .B2(n51500), .A(n14956), .ZN(n14691) );
  NAND2_X1 U25520 ( .A1(n14946), .A2(n2151), .ZN(n14690) );
  NAND3_X1 U25521 ( .A1(n14950), .A2(n15278), .A3(n14956), .ZN(n14689) );
  NOR2_X1 U25522 ( .A1(n14962), .A2(n15278), .ZN(n14940) );
  NAND3_X1 U25523 ( .A1(n14940), .A2(n15279), .A3(n14956), .ZN(n14688) );
  NAND4_X1 U25524 ( .A1(n14691), .A2(n14690), .A3(n14689), .A4(n14688), .ZN(
        n14695) );
  OR2_X1 U25525 ( .A1(n14692), .A2(n15279), .ZN(n15288) );
  INV_X1 U25526 ( .A(n15288), .ZN(n14693) );
  NAND2_X1 U25527 ( .A1(n51724), .A2(n14693), .ZN(n14694) );
  XNOR2_X1 U25528 ( .A(n14699), .B(n15504), .ZN(n14736) );
  NAND2_X1 U25529 ( .A1(n14703), .A2(n51670), .ZN(n14705) );
  NAND4_X1 U25530 ( .A1(n14705), .A2(n14704), .A3(n14719), .A4(n14720), .ZN(
        n14706) );
  AND2_X1 U25531 ( .A1(n14707), .A2(n14706), .ZN(n14729) );
  NOR2_X1 U25532 ( .A1(n14713), .A2(n14711), .ZN(n14708) );
  AOI22_X1 U25533 ( .A1(n14710), .A2(n14709), .B1(n14721), .B2(n14708), .ZN(
        n14728) );
  OAI21_X1 U25534 ( .B1(n14713), .B2(n14712), .A(n14711), .ZN(n14714) );
  NAND2_X1 U25535 ( .A1(n14714), .A2(n14717), .ZN(n14715) );
  OAI211_X1 U25536 ( .C1(n14717), .C2(n14716), .A(n14715), .B(n14720), .ZN(
        n14727) );
  OAI21_X1 U25537 ( .B1(n14720), .B2(n14719), .A(n14718), .ZN(n14725) );
  INV_X1 U25538 ( .A(n14722), .ZN(n14723) );
  NAND4_X1 U25539 ( .A1(n14725), .A2(n14724), .A3(n13343), .A4(n14723), .ZN(
        n14726) );
  XNOR2_X1 U25540 ( .A(n18738), .B(n18134), .ZN(n14730) );
  XNOR2_X1 U25541 ( .A(n17821), .B(n14730), .ZN(n16383) );
  XNOR2_X1 U25542 ( .A(n17965), .B(n17829), .ZN(n17679) );
  XNOR2_X1 U25543 ( .A(n2203), .B(n4855), .ZN(n42258) );
  XNOR2_X1 U25544 ( .A(n42258), .B(n4655), .ZN(n24932) );
  XNOR2_X1 U25545 ( .A(n45463), .B(n49790), .ZN(n17684) );
  XNOR2_X1 U25546 ( .A(n24932), .B(n17684), .ZN(n17825) );
  XNOR2_X1 U25547 ( .A(n17825), .B(n4824), .ZN(n34125) );
  XNOR2_X1 U25548 ( .A(n4754), .B(n4782), .ZN(n26604) );
  XNOR2_X1 U25549 ( .A(n34711), .B(n26604), .ZN(n14731) );
  XNOR2_X1 U25550 ( .A(n34125), .B(n14731), .ZN(n14732) );
  XNOR2_X1 U25551 ( .A(n14732), .B(n19262), .ZN(n14733) );
  XNOR2_X1 U25552 ( .A(n17679), .B(n14733), .ZN(n14734) );
  XNOR2_X1 U25553 ( .A(n16383), .B(n14734), .ZN(n14735) );
  XNOR2_X1 U25554 ( .A(n14736), .B(n14735), .ZN(n14737) );
  NOR2_X1 U25555 ( .A1(n14744), .A2(n20468), .ZN(n14743) );
  NAND2_X1 U25556 ( .A1(n20474), .A2(n51130), .ZN(n20396) );
  INV_X1 U25557 ( .A(n20396), .ZN(n14742) );
  AND2_X1 U25558 ( .A1(n20393), .A2(n14738), .ZN(n17997) );
  INV_X1 U25559 ( .A(n17997), .ZN(n20397) );
  AOI22_X1 U25560 ( .A1(n14743), .A2(n20473), .B1(n14742), .B2(n20397), .ZN(
        n14747) );
  INV_X1 U25561 ( .A(n14744), .ZN(n14745) );
  NAND4_X1 U25562 ( .A1(n14749), .A2(n14748), .A3(n14747), .A4(n14746), .ZN(
        n14752) );
  NAND2_X1 U25563 ( .A1(n20383), .A2(n18000), .ZN(n20389) );
  MUX2_X1 U25564 ( .A(n20389), .B(n20473), .S(n20468), .Z(n20484) );
  NOR2_X1 U25565 ( .A1(n17636), .A2(n17999), .ZN(n14750) );
  INV_X1 U25566 ( .A(n20400), .ZN(n14751) );
  XNOR2_X1 U25567 ( .A(n4884), .B(n4879), .ZN(n14753) );
  XNOR2_X1 U25568 ( .A(n14753), .B(n4744), .ZN(n14754) );
  XNOR2_X1 U25569 ( .A(n14754), .B(n26525), .ZN(n17993) );
  XOR2_X1 U25570 ( .A(n4694), .B(n4627), .Z(n14755) );
  XNOR2_X1 U25571 ( .A(n17993), .B(n14755), .ZN(n33086) );
  XNOR2_X1 U25572 ( .A(n35815), .B(n4890), .ZN(n43849) );
  XNOR2_X1 U25573 ( .A(n33086), .B(n43849), .ZN(n14756) );
  XNOR2_X1 U25574 ( .A(n42721), .B(n28390), .ZN(n24625) );
  XNOR2_X1 U25575 ( .A(n4537), .B(n33221), .ZN(n16149) );
  XNOR2_X1 U25576 ( .A(n16149), .B(n7744), .ZN(n43136) );
  XNOR2_X1 U25577 ( .A(n24625), .B(n43136), .ZN(n42846) );
  XNOR2_X1 U25578 ( .A(n14756), .B(n42846), .ZN(n14757) );
  XNOR2_X1 U25579 ( .A(n18432), .B(n14757), .ZN(n14758) );
  XNOR2_X1 U25580 ( .A(n14758), .B(n17787), .ZN(n14775) );
  OAI21_X1 U25581 ( .B1(n14759), .B2(n15189), .A(n15243), .ZN(n14760) );
  NOR3_X1 U25582 ( .A1(n14766), .A2(n15244), .A3(n14765), .ZN(n14768) );
  OR2_X1 U25583 ( .A1(n15206), .A2(n15244), .ZN(n15248) );
  OAI22_X1 U25584 ( .A1(n14769), .A2(n14768), .B1(n15248), .B2(n14767), .ZN(
        n14770) );
  XNOR2_X2 U25585 ( .A(n17793), .B(n18548), .ZN(n18615) );
  XNOR2_X1 U25586 ( .A(n18615), .B(n14775), .ZN(n14776) );
  XNOR2_X1 U25587 ( .A(n14776), .B(n16454), .ZN(n14779) );
  XNOR2_X1 U25588 ( .A(n15519), .B(n51481), .ZN(n14777) );
  XNOR2_X1 U25589 ( .A(n51133), .B(n14777), .ZN(n14778) );
  XNOR2_X1 U25590 ( .A(n14778), .B(n14779), .ZN(n14804) );
  XNOR2_X1 U25591 ( .A(n18450), .B(n16158), .ZN(n16455) );
  INV_X1 U25592 ( .A(n14780), .ZN(n14781) );
  NAND2_X1 U25593 ( .A1(n14782), .A2(n14781), .ZN(n14802) );
  AND2_X1 U25594 ( .A1(n14787), .A2(n14786), .ZN(n14801) );
  INV_X1 U25595 ( .A(n14788), .ZN(n14789) );
  NOR2_X1 U25596 ( .A1(n14789), .A2(n15256), .ZN(n14793) );
  NAND2_X1 U25597 ( .A1(n14795), .A2(n15257), .ZN(n14799) );
  NAND2_X1 U25598 ( .A1(n14796), .A2(n15256), .ZN(n14798) );
  NAND4_X1 U25599 ( .A1(n14799), .A2(n14798), .A3(n51686), .A4(n14797), .ZN(
        n14800) );
  XNOR2_X1 U25600 ( .A(n16455), .B(n16527), .ZN(n16719) );
  XNOR2_X1 U25601 ( .A(n14804), .B(n16719), .ZN(n18288) );
  INV_X1 U25602 ( .A(n18288), .ZN(n15094) );
  NOR2_X1 U25603 ( .A1(n14806), .A2(n14805), .ZN(n14825) );
  NOR2_X1 U25604 ( .A1(n7906), .A2(n15384), .ZN(n14819) );
  INV_X1 U25606 ( .A(n14808), .ZN(n14811) );
  INV_X1 U25607 ( .A(n14809), .ZN(n14810) );
  NAND3_X1 U25608 ( .A1(n14811), .A2(n14810), .A3(n11853), .ZN(n14816) );
  NAND3_X1 U25609 ( .A1(n14813), .A2(n15365), .A3(n14812), .ZN(n14814) );
  NAND4_X1 U25610 ( .A1(n11853), .A2(n787), .A3(n15359), .A4(n14814), .ZN(
        n14815) );
  INV_X1 U25611 ( .A(n14818), .ZN(n15362) );
  AOI22_X1 U25612 ( .A1(n14820), .A2(n15367), .B1(n14819), .B2(n15385), .ZN(
        n14823) );
  NOR2_X1 U25613 ( .A1(n15380), .A2(n15384), .ZN(n15366) );
  NAND2_X1 U25614 ( .A1(n14821), .A2(n15366), .ZN(n14822) );
  NOR2_X1 U25615 ( .A1(n15437), .A2(n15438), .ZN(n15329) );
  AOI22_X1 U25616 ( .A1(n15329), .A2(n15342), .B1(n8697), .B2(n15437), .ZN(
        n14834) );
  INV_X1 U25617 ( .A(n14828), .ZN(n14829) );
  OAI21_X1 U25618 ( .B1(n15341), .B2(n15434), .A(n14829), .ZN(n14830) );
  INV_X1 U25619 ( .A(n15436), .ZN(n15326) );
  NOR2_X1 U25620 ( .A1(n15334), .A2(n15324), .ZN(n15444) );
  AND2_X1 U25621 ( .A1(n15437), .A2(n15325), .ZN(n14832) );
  OAI22_X1 U25622 ( .A1(n14832), .A2(n14863), .B1(n51698), .B2(n15434), .ZN(
        n14833) );
  XNOR2_X1 U25623 ( .A(n52229), .B(n14835), .ZN(n17942) );
  INV_X1 U25624 ( .A(n17942), .ZN(n14846) );
  NAND2_X1 U25625 ( .A1(n14837), .A2(n14836), .ZN(n15760) );
  INV_X1 U25626 ( .A(n15760), .ZN(n14838) );
  NAND2_X1 U25627 ( .A1(n14838), .A2(n15758), .ZN(n15763) );
  XNOR2_X1 U25628 ( .A(n4624), .B(n4558), .ZN(n25147) );
  XNOR2_X1 U25629 ( .A(n42077), .B(n25147), .ZN(n17809) );
  INV_X1 U25630 ( .A(n17809), .ZN(n35532) );
  XNOR2_X1 U25631 ( .A(n35532), .B(n37288), .ZN(n24956) );
  XNOR2_X1 U25632 ( .A(n4647), .B(n3276), .ZN(n18423) );
  XNOR2_X1 U25633 ( .A(n27174), .B(n18423), .ZN(n36698) );
  XNOR2_X1 U25634 ( .A(n24956), .B(n36698), .ZN(n16136) );
  XNOR2_X1 U25635 ( .A(n16136), .B(n49323), .ZN(n33856) );
  XNOR2_X1 U25636 ( .A(n2903), .B(n3336), .ZN(n26506) );
  XNOR2_X1 U25637 ( .A(n26506), .B(n4208), .ZN(n14839) );
  XNOR2_X1 U25638 ( .A(n46097), .B(n14839), .ZN(n34046) );
  XNOR2_X1 U25639 ( .A(n34046), .B(n47401), .ZN(n14840) );
  XNOR2_X1 U25640 ( .A(n33856), .B(n14840), .ZN(n14841) );
  XNOR2_X1 U25641 ( .A(n15763), .B(n14841), .ZN(n14842) );
  XNOR2_X1 U25642 ( .A(n14842), .B(n17802), .ZN(n14844) );
  XNOR2_X1 U25643 ( .A(n15680), .B(n17125), .ZN(n14843) );
  XNOR2_X1 U25644 ( .A(n14844), .B(n14843), .ZN(n14845) );
  XNOR2_X1 U25645 ( .A(n14846), .B(n14845), .ZN(n14852) );
  XNOR2_X1 U25646 ( .A(n14847), .B(n17127), .ZN(n18420) );
  INV_X1 U25647 ( .A(n18420), .ZN(n14850) );
  XNOR2_X1 U25648 ( .A(n14848), .B(n18791), .ZN(n15681) );
  INV_X1 U25649 ( .A(n15681), .ZN(n16703) );
  XNOR2_X1 U25650 ( .A(n16703), .B(n15511), .ZN(n14849) );
  XNOR2_X1 U25651 ( .A(n14850), .B(n14849), .ZN(n14851) );
  XNOR2_X2 U25652 ( .A(n14852), .B(n14851), .ZN(n18294) );
  INV_X1 U25653 ( .A(n18294), .ZN(n15093) );
  XNOR2_X2 U25654 ( .A(n16162), .B(n17158), .ZN(n19227) );
  XNOR2_X1 U25655 ( .A(n19227), .B(n51758), .ZN(n17912) );
  XNOR2_X1 U25656 ( .A(n24828), .B(n25042), .ZN(n25575) );
  XNOR2_X1 U25657 ( .A(n16739), .B(n4454), .ZN(n23711) );
  XNOR2_X1 U25658 ( .A(n25575), .B(n23711), .ZN(n28413) );
  XNOR2_X2 U25659 ( .A(n42769), .B(n49414), .ZN(n24430) );
  XNOR2_X1 U25660 ( .A(n28413), .B(n24430), .ZN(n33445) );
  INV_X1 U25661 ( .A(n33445), .ZN(n14854) );
  XNOR2_X1 U25662 ( .A(n4706), .B(n4536), .ZN(n27364) );
  XNOR2_X1 U25663 ( .A(n27364), .B(n4752), .ZN(n14853) );
  XNOR2_X1 U25664 ( .A(n14854), .B(n14853), .ZN(n33545) );
  XNOR2_X1 U25665 ( .A(n28270), .B(n25718), .ZN(n34479) );
  XNOR2_X1 U25666 ( .A(n34479), .B(n4847), .ZN(n14855) );
  XNOR2_X1 U25667 ( .A(n33545), .B(n14855), .ZN(n14856) );
  XNOR2_X1 U25668 ( .A(n15650), .B(n14856), .ZN(n14857) );
  XNOR2_X1 U25669 ( .A(n14857), .B(n16620), .ZN(n14858) );
  XNOR2_X1 U25670 ( .A(n17906), .B(n14859), .ZN(n16746) );
  OAI21_X1 U25671 ( .B1(n14860), .B2(n51699), .A(n15434), .ZN(n14869) );
  NAND2_X1 U25672 ( .A1(n51700), .A2(n15437), .ZN(n14862) );
  NAND4_X1 U25673 ( .A1(n14861), .A2(n15335), .A3(n15438), .A4(n15324), .ZN(
        n15445) );
  AND2_X1 U25674 ( .A1(n14862), .A2(n15445), .ZN(n14868) );
  OAI21_X1 U25675 ( .B1(n14863), .B2(n15437), .A(n15338), .ZN(n14865) );
  MUX2_X1 U25677 ( .A(n14865), .B(n14864), .S(n15435), .Z(n14867) );
  OAI21_X1 U25678 ( .B1(n15338), .B2(n15437), .A(n15326), .ZN(n14866) );
  AND4_X1 U25679 ( .A1(n1555), .A2(n14871), .A3(n1556), .A4(n14870), .ZN(
        n14874) );
  AOI22_X1 U25680 ( .A1(n14875), .A2(n14874), .B1(n14873), .B2(n14872), .ZN(
        n14881) );
  OAI21_X1 U25681 ( .B1(n14877), .B2(n7245), .A(n14876), .ZN(n14878) );
  NAND3_X1 U25682 ( .A1(n14878), .A2(n2249), .A3(n15414), .ZN(n14879) );
  INV_X1 U25684 ( .A(n18181), .ZN(n14882) );
  XNOR2_X1 U25685 ( .A(n18394), .B(n14882), .ZN(n14891) );
  OAI21_X1 U25686 ( .B1(n14885), .B2(n14884), .A(n14883), .ZN(n14888) );
  OAI211_X1 U25687 ( .C1(n14889), .C2(n14888), .A(n14887), .B(n14886), .ZN(
        n17778) );
  XNOR2_X1 U25688 ( .A(n17778), .B(n17771), .ZN(n15653) );
  INV_X1 U25689 ( .A(n15653), .ZN(n16613) );
  XNOR2_X1 U25690 ( .A(n16613), .B(n16105), .ZN(n14890) );
  XNOR2_X1 U25691 ( .A(n14890), .B(n14891), .ZN(n15962) );
  INV_X1 U25692 ( .A(n14893), .ZN(n14892) );
  INV_X1 U25693 ( .A(n4883), .ZN(n48885) );
  OR2_X1 U25694 ( .A1(n14897), .A2(n4883), .ZN(n14900) );
  NOR2_X1 U25695 ( .A1(n14894), .A2(n14893), .ZN(n14898) );
  INV_X1 U25696 ( .A(n14895), .ZN(n14896) );
  NAND4_X1 U25697 ( .A1(n14898), .A2(n4883), .A3(n14897), .A4(n14896), .ZN(
        n14899) );
  NAND3_X1 U25698 ( .A1(n14901), .A2(n14900), .A3(n14899), .ZN(n14902) );
  XNOR2_X1 U25699 ( .A(n16498), .B(n14902), .ZN(n16320) );
  XNOR2_X1 U25700 ( .A(n4605), .B(Key[159]), .ZN(n33635) );
  XNOR2_X1 U25701 ( .A(n2599), .B(n33635), .ZN(n43019) );
  XNOR2_X1 U25702 ( .A(n45105), .B(n43019), .ZN(n42592) );
  INV_X1 U25703 ( .A(Key[3]), .ZN(n47533) );
  XNOR2_X1 U25704 ( .A(n47533), .B(Key[27]), .ZN(n17880) );
  INV_X1 U25705 ( .A(n17880), .ZN(n34414) );
  XNOR2_X1 U25706 ( .A(n4565), .B(n4423), .ZN(n43863) );
  XNOR2_X1 U25707 ( .A(n34414), .B(n43863), .ZN(n35110) );
  XNOR2_X1 U25708 ( .A(n45106), .B(n4739), .ZN(n14904) );
  XNOR2_X1 U25709 ( .A(n35110), .B(n14904), .ZN(n14905) );
  XNOR2_X1 U25710 ( .A(n42592), .B(n14905), .ZN(n14906) );
  XNOR2_X1 U25711 ( .A(n14903), .B(n14906), .ZN(n14907) );
  XNOR2_X1 U25712 ( .A(n17754), .B(n14907), .ZN(n14908) );
  XNOR2_X1 U25714 ( .A(n18153), .B(n17232), .ZN(n14910) );
  XNOR2_X1 U25715 ( .A(n41155), .B(n4885), .ZN(n25683) );
  XNOR2_X1 U25716 ( .A(n18668), .B(n25683), .ZN(n14909) );
  XNOR2_X1 U25717 ( .A(n14910), .B(n14909), .ZN(n14934) );
  MUX2_X1 U25718 ( .A(n14911), .B(n7572), .S(n15770), .Z(n14913) );
  NAND3_X1 U25719 ( .A1(n14913), .A2(n14912), .A3(n15766), .ZN(n14918) );
  NOR2_X1 U25720 ( .A1(n14914), .A2(n15073), .ZN(n14916) );
  INV_X1 U25721 ( .A(n15063), .ZN(n14915) );
  NAND4_X1 U25722 ( .A1(n14916), .A2(n14929), .A3(n14915), .A4(n15068), .ZN(
        n14917) );
  AND2_X1 U25723 ( .A1(n14918), .A2(n14917), .ZN(n14933) );
  AOI21_X1 U25724 ( .B1(n14929), .B2(n2189), .A(n15063), .ZN(n14922) );
  INV_X1 U25725 ( .A(n14919), .ZN(n14920) );
  NAND2_X1 U25726 ( .A1(n15769), .A2(n15770), .ZN(n14921) );
  AND2_X1 U25727 ( .A1(n15300), .A2(n2189), .ZN(n14923) );
  NAND2_X1 U25728 ( .A1(n15067), .A2(n2189), .ZN(n15076) );
  INV_X1 U25729 ( .A(n15076), .ZN(n14927) );
  INV_X1 U25730 ( .A(n14925), .ZN(n14926) );
  NAND4_X1 U25731 ( .A1(n14929), .A2(n14927), .A3(n15307), .A4(n14926), .ZN(
        n14928) );
  INV_X1 U25732 ( .A(n15846), .ZN(n16641) );
  XNOR2_X1 U25733 ( .A(n14934), .B(n16641), .ZN(n15666) );
  AND2_X1 U25734 ( .A1(n15280), .A2(n15278), .ZN(n14937) );
  NAND4_X1 U25735 ( .A1(n14937), .A2(n14945), .A3(n14951), .A4(n14936), .ZN(
        n14943) );
  NAND2_X1 U25736 ( .A1(n14950), .A2(n14957), .ZN(n14941) );
  NAND4_X1 U25737 ( .A1(n14939), .A2(n14940), .A3(n14941), .A4(n14956), .ZN(
        n14942) );
  NAND2_X1 U25738 ( .A1(n14958), .A2(n14957), .ZN(n14944) );
  NOR2_X1 U25739 ( .A1(n14945), .A2(n14944), .ZN(n14948) );
  INV_X1 U25740 ( .A(n14946), .ZN(n14947) );
  XNOR2_X1 U25741 ( .A(n14950), .B(n51500), .ZN(n14954) );
  INV_X1 U25742 ( .A(n14951), .ZN(n14953) );
  INV_X1 U25743 ( .A(n14955), .ZN(n14963) );
  AOI21_X1 U25744 ( .B1(n15274), .B2(n14956), .A(n15279), .ZN(n14961) );
  OAI211_X1 U25745 ( .C1(n14959), .C2(n14958), .A(n14962), .B(n14957), .ZN(
        n14960) );
  XNOR2_X1 U25746 ( .A(n16412), .B(n18414), .ZN(n14965) );
  XNOR2_X1 U25747 ( .A(n15668), .B(n14965), .ZN(n16209) );
  NOR2_X1 U25749 ( .A1(n18282), .A2(n590), .ZN(n16797) );
  OAI21_X1 U25752 ( .B1(n14972), .B2(n14971), .A(n14970), .ZN(n19185) );
  XNOR2_X1 U25753 ( .A(n18827), .B(n19185), .ZN(n14973) );
  XNOR2_X1 U25754 ( .A(n14973), .B(n18832), .ZN(n14989) );
  NAND2_X1 U25755 ( .A1(n14975), .A2(n14974), .ZN(n14988) );
  OAI21_X1 U25756 ( .B1(n15108), .B2(n352), .A(n14976), .ZN(n15101) );
  INV_X1 U25757 ( .A(n15101), .ZN(n14987) );
  INV_X1 U25758 ( .A(n14977), .ZN(n14981) );
  INV_X1 U25759 ( .A(n14978), .ZN(n14979) );
  OAI21_X1 U25760 ( .B1(n14981), .B2(n14980), .A(n14979), .ZN(n14986) );
  NOR2_X1 U25761 ( .A1(n15106), .A2(n14982), .ZN(n15115) );
  OAI21_X1 U25762 ( .B1(n14984), .B2(n14983), .A(n15115), .ZN(n14985) );
  XNOR2_X1 U25763 ( .A(n16176), .B(n14989), .ZN(n17959) );
  XNOR2_X1 U25764 ( .A(n17847), .B(n4526), .ZN(n14990) );
  XNOR2_X1 U25765 ( .A(n14990), .B(n18479), .ZN(n19190) );
  NAND2_X1 U25766 ( .A1(n15133), .A2(n8514), .ZN(n14991) );
  INV_X1 U25767 ( .A(n15137), .ZN(n14997) );
  OAI21_X1 U25768 ( .B1(n14995), .B2(n14994), .A(n14993), .ZN(n14996) );
  OAI21_X1 U25769 ( .B1(n15138), .B2(n15131), .A(n14999), .ZN(n15003) );
  NAND3_X1 U25770 ( .A1(n15000), .A2(n15138), .A3(n14999), .ZN(n15002) );
  INV_X1 U25771 ( .A(n15139), .ZN(n15001) );
  XNOR2_X1 U25772 ( .A(n18483), .B(n4687), .ZN(n15004) );
  XNOR2_X1 U25773 ( .A(n19190), .B(n15889), .ZN(n15005) );
  XNOR2_X1 U25774 ( .A(n15005), .B(n17959), .ZN(n15017) );
  XNOR2_X1 U25775 ( .A(n16571), .B(n16435), .ZN(n15012) );
  XNOR2_X1 U25776 ( .A(n43586), .B(n43105), .ZN(n26244) );
  XNOR2_X1 U25777 ( .A(n2601), .B(n4048), .ZN(n15006) );
  XNOR2_X1 U25778 ( .A(n26244), .B(n15006), .ZN(n15008) );
  XNOR2_X1 U25779 ( .A(n27297), .B(n4823), .ZN(n43879) );
  INV_X1 U25780 ( .A(n33474), .ZN(n15007) );
  XNOR2_X1 U25781 ( .A(n43879), .B(n15007), .ZN(n43985) );
  XNOR2_X1 U25782 ( .A(n15008), .B(n43985), .ZN(n34462) );
  XNOR2_X1 U25783 ( .A(n40104), .B(n48814), .ZN(n25520) );
  XOR2_X1 U25784 ( .A(n4502), .B(n6031), .Z(n15009) );
  XNOR2_X1 U25785 ( .A(n25520), .B(n15009), .ZN(n33477) );
  XNOR2_X1 U25786 ( .A(n34462), .B(n33477), .ZN(n15010) );
  XNOR2_X1 U25787 ( .A(n17954), .B(n15010), .ZN(n15011) );
  XNOR2_X1 U25788 ( .A(n15012), .B(n15011), .ZN(n15013) );
  XNOR2_X1 U25789 ( .A(n15013), .B(n16431), .ZN(n15015) );
  XNOR2_X1 U25790 ( .A(n15014), .B(n18475), .ZN(n15719) );
  XNOR2_X1 U25791 ( .A(n16782), .B(n15719), .ZN(n17839) );
  XNOR2_X1 U25792 ( .A(n17839), .B(n15015), .ZN(n15016) );
  XNOR2_X1 U25795 ( .A(n18599), .B(n17821), .ZN(n15019) );
  XNOR2_X1 U25796 ( .A(n42258), .B(n41367), .ZN(n27316) );
  XNOR2_X1 U25797 ( .A(n27316), .B(n42327), .ZN(n15492) );
  INV_X1 U25798 ( .A(n15492), .ZN(n15020) );
  XNOR2_X1 U25799 ( .A(n15020), .B(n4930), .ZN(n33119) );
  XNOR2_X1 U25800 ( .A(n23882), .B(n4838), .ZN(n16476) );
  XNOR2_X1 U25801 ( .A(n4923), .B(n4712), .ZN(n15987) );
  XNOR2_X1 U25802 ( .A(n16476), .B(n15987), .ZN(n36945) );
  XNOR2_X1 U25803 ( .A(n36941), .B(n49790), .ZN(n15021) );
  XNOR2_X1 U25804 ( .A(n36945), .B(n15021), .ZN(n15022) );
  XNOR2_X1 U25805 ( .A(n33119), .B(n15022), .ZN(n15023) );
  XNOR2_X1 U25806 ( .A(n17829), .B(n15023), .ZN(n15024) );
  XNOR2_X1 U25807 ( .A(n8699), .B(n15024), .ZN(n15025) );
  XNOR2_X1 U25808 ( .A(n15026), .B(n15025), .ZN(n15027) );
  INV_X1 U25809 ( .A(n15029), .ZN(n15032) );
  AOI22_X1 U25810 ( .A1(n15035), .A2(n15032), .B1(n15031), .B2(n15030), .ZN(
        n15058) );
  NOR2_X1 U25811 ( .A1(n15033), .A2(n277), .ZN(n15037) );
  NAND2_X1 U25812 ( .A1(n15035), .A2(n15034), .ZN(n15036) );
  AOI22_X1 U25813 ( .A1(n15039), .A2(n15038), .B1(n15037), .B2(n15036), .ZN(
        n15057) );
  NOR2_X1 U25815 ( .A1(n15041), .A2(n15044), .ZN(n15042) );
  NAND2_X1 U25816 ( .A1(n15045), .A2(n15044), .ZN(n15055) );
  NAND3_X1 U25817 ( .A1(n15048), .A2(n15047), .A3(n15046), .ZN(n15053) );
  INV_X1 U25818 ( .A(n15049), .ZN(n15051) );
  NAND2_X1 U25819 ( .A1(n15051), .A2(n277), .ZN(n15052) );
  NAND4_X1 U25820 ( .A1(n15055), .A2(n15054), .A3(n15053), .A4(n15052), .ZN(
        n15056) );
  XNOR2_X1 U25821 ( .A(n4529), .B(n47268), .ZN(n42686) );
  XNOR2_X1 U25822 ( .A(n42686), .B(n28070), .ZN(n23887) );
  INV_X1 U25823 ( .A(n23887), .ZN(n33131) );
  XNOR2_X1 U25824 ( .A(n16754), .B(n33131), .ZN(n15059) );
  XNOR2_X1 U25825 ( .A(n15059), .B(n18602), .ZN(n15086) );
  OAI211_X1 U25826 ( .C1(n15062), .C2(n15766), .A(n15061), .B(n15306), .ZN(
        n15065) );
  NAND3_X1 U25827 ( .A1(n15306), .A2(n1486), .A3(n15063), .ZN(n15064) );
  NAND3_X1 U25828 ( .A1(n15065), .A2(n15303), .A3(n15064), .ZN(n15079) );
  AOI21_X1 U25829 ( .B1(n15068), .B2(n15067), .A(n15066), .ZN(n15074) );
  NAND2_X1 U25830 ( .A1(n15069), .A2(n15307), .ZN(n15072) );
  NAND4_X1 U25833 ( .A1(n15074), .A2(n15073), .A3(n15072), .A4(n15071), .ZN(
        n15075) );
  OAI21_X1 U25834 ( .B1(n15077), .B2(n15076), .A(n15075), .ZN(n15078) );
  NOR2_X1 U25835 ( .A1(n15079), .A2(n15078), .ZN(n15084) );
  INV_X1 U25836 ( .A(n15305), .ZN(n15080) );
  NAND2_X1 U25837 ( .A1(n15766), .A2(n15080), .ZN(n15082) );
  MUX2_X1 U25838 ( .A(n15304), .B(n15082), .S(n15081), .Z(n15083) );
  XNOR2_X1 U25839 ( .A(n19261), .B(n18712), .ZN(n15085) );
  XNOR2_X1 U25840 ( .A(n15086), .B(n15085), .ZN(n15088) );
  XNOR2_X1 U25841 ( .A(n17690), .B(n17297), .ZN(n15087) );
  INV_X1 U25842 ( .A(n18464), .ZN(n18603) );
  XNOR2_X1 U25843 ( .A(n15087), .B(n18603), .ZN(n15736) );
  XNOR2_X1 U25844 ( .A(n15088), .B(n15736), .ZN(n15709) );
  NAND2_X1 U25845 ( .A1(n17522), .A2(n6952), .ZN(n20014) );
  NAND2_X1 U25846 ( .A1(n590), .A2(n17522), .ZN(n15090) );
  NOR2_X1 U25847 ( .A1(n17533), .A2(n15090), .ZN(n20024) );
  NAND2_X1 U25848 ( .A1(n16798), .A2(n18287), .ZN(n17525) );
  NAND2_X1 U25850 ( .A1(n633), .A2(n20021), .ZN(n20019) );
  INV_X1 U25851 ( .A(n20015), .ZN(n17535) );
  OAI21_X1 U25852 ( .B1(n17525), .B2(n20019), .A(n17535), .ZN(n15092) );
  NAND2_X1 U25853 ( .A1(n15092), .A2(n51208), .ZN(n15098) );
  NAND3_X1 U25854 ( .A1(n18282), .A2(n590), .A3(n20021), .ZN(n17487) );
  AOI21_X1 U25855 ( .B1(n18292), .B2(n17487), .A(n6952), .ZN(n15096) );
  NAND3_X1 U25856 ( .A1(n16798), .A2(n2166), .A3(n17489), .ZN(n17516) );
  NAND3_X1 U25858 ( .A1(n18282), .A2(n51209), .A3(n20015), .ZN(n17520) );
  OAI21_X1 U25859 ( .B1(n15094), .B2(n17516), .A(n17520), .ZN(n15095) );
  NOR2_X1 U25860 ( .A1(n15096), .A2(n15095), .ZN(n15097) );
  MUX2_X1 U25861 ( .A(n15119), .B(n15107), .S(n8075), .Z(n15112) );
  AND2_X1 U25862 ( .A1(n8075), .A2(n352), .ZN(n15104) );
  INV_X1 U25863 ( .A(n15104), .ZN(n15105) );
  NAND3_X1 U25864 ( .A1(n15107), .A2(n15106), .A3(n15105), .ZN(n15111) );
  OR2_X1 U25865 ( .A1(n15109), .A2(n15108), .ZN(n15110) );
  NAND2_X1 U25866 ( .A1(n15114), .A2(n15113), .ZN(n15116) );
  NOR2_X1 U25867 ( .A1(n15116), .A2(n15115), .ZN(n15121) );
  NAND2_X1 U25868 ( .A1(n15118), .A2(n15117), .ZN(n15120) );
  MUX2_X1 U25869 ( .A(n15121), .B(n15120), .S(n15119), .Z(n15122) );
  XNOR2_X1 U25870 ( .A(n16450), .B(n51135), .ZN(n15123) );
  XNOR2_X1 U25871 ( .A(n15123), .B(n2200), .ZN(n15124) );
  XNOR2_X1 U25872 ( .A(n15125), .B(n15124), .ZN(n18186) );
  NAND3_X1 U25873 ( .A1(n15127), .A2(n15136), .A3(n15126), .ZN(n15130) );
  NAND3_X1 U25874 ( .A1(n15130), .A2(n15129), .A3(n15128), .ZN(n15141) );
  NOR3_X1 U25875 ( .A1(n15133), .A2(n15132), .A3(n15131), .ZN(n15135) );
  NAND3_X1 U25876 ( .A1(n15139), .A2(n14269), .A3(n15138), .ZN(n15140) );
  XNOR2_X1 U25877 ( .A(n51458), .B(n18550), .ZN(n15148) );
  XNOR2_X1 U25878 ( .A(n45051), .B(n33374), .ZN(n17661) );
  XNOR2_X1 U25879 ( .A(n4645), .B(n4618), .ZN(n15908) );
  XNOR2_X1 U25880 ( .A(n15908), .B(n15142), .ZN(n33845) );
  XNOR2_X1 U25881 ( .A(n17661), .B(n33845), .ZN(n24738) );
  XNOR2_X1 U25882 ( .A(n24738), .B(n17993), .ZN(n34030) );
  XNOR2_X1 U25883 ( .A(Key[23]), .B(n46552), .ZN(n25898) );
  XNOR2_X1 U25884 ( .A(n25898), .B(n4537), .ZN(n15143) );
  XNOR2_X1 U25885 ( .A(n15143), .B(n2604), .ZN(n15144) );
  XNOR2_X1 U25886 ( .A(n34030), .B(n15144), .ZN(n15145) );
  XNOR2_X1 U25887 ( .A(n16023), .B(n15145), .ZN(n15146) );
  XNOR2_X1 U25888 ( .A(n15519), .B(n15146), .ZN(n15147) );
  XNOR2_X1 U25889 ( .A(n15149), .B(n17787), .ZN(n16715) );
  AOI21_X1 U25890 ( .B1(n836), .B2(n15151), .A(n15150), .ZN(n15153) );
  XNOR2_X1 U25892 ( .A(n16715), .B(n16593), .ZN(n16521) );
  INV_X1 U25893 ( .A(n16521), .ZN(n15156) );
  NAND2_X1 U25894 ( .A1(n15160), .A2(n51452), .ZN(n15184) );
  AOI21_X1 U25895 ( .B1(n15163), .B2(n15162), .A(n15161), .ZN(n15166) );
  NAND3_X1 U25896 ( .A1(n15166), .A2(n15165), .A3(n15164), .ZN(n15170) );
  NAND3_X1 U25897 ( .A1(n15168), .A2(n15179), .A3(n15167), .ZN(n15169) );
  AND2_X1 U25898 ( .A1(n15170), .A2(n15169), .ZN(n15183) );
  NAND2_X1 U25899 ( .A1(n15172), .A2(n15171), .ZN(n15175) );
  NAND3_X1 U25900 ( .A1(n15175), .A2(n15174), .A3(n15173), .ZN(n15182) );
  OAI21_X1 U25901 ( .B1(n15178), .B2(n15177), .A(n15176), .ZN(n15180) );
  NAND2_X1 U25902 ( .A1(n15180), .A2(n15179), .ZN(n15181) );
  NAND4_X2 U25903 ( .A1(n15184), .A2(n15181), .A3(n15182), .A4(n15183), .ZN(
        n17803) );
  XNOR2_X1 U25904 ( .A(n17803), .B(n17804), .ZN(n17644) );
  XNOR2_X1 U25905 ( .A(n17938), .B(n15185), .ZN(n15186) );
  XNOR2_X1 U25908 ( .A(n18430), .B(n15680), .ZN(n15212) );
  INV_X1 U25909 ( .A(n15187), .ZN(n15191) );
  OAI21_X1 U25910 ( .B1(n15243), .B2(n15189), .A(n15188), .ZN(n15249) );
  NAND3_X1 U25911 ( .A1(n15249), .A2(n15235), .A3(n15244), .ZN(n15190) );
  AND2_X1 U25912 ( .A1(n15191), .A2(n15190), .ZN(n15211) );
  NOR2_X1 U25913 ( .A1(n15233), .A2(n15244), .ZN(n15192) );
  AOI22_X1 U25914 ( .A1(n15245), .A2(n15193), .B1(n15235), .B2(n15192), .ZN(
        n15210) );
  INV_X1 U25915 ( .A(n15194), .ZN(n15195) );
  NOR2_X1 U25916 ( .A1(n15206), .A2(n15195), .ZN(n15202) );
  INV_X1 U25917 ( .A(n15197), .ZN(n15198) );
  OAI22_X1 U25918 ( .A1(n15200), .A2(n15199), .B1(n15198), .B2(n15233), .ZN(
        n15201) );
  AOI21_X1 U25919 ( .B1(n15203), .B2(n15202), .A(n15201), .ZN(n15209) );
  NAND4_X1 U25920 ( .A1(n15207), .A2(n15206), .A3(n15205), .A4(n15204), .ZN(
        n15208) );
  XNOR2_X1 U25921 ( .A(n17125), .B(n18427), .ZN(n15606) );
  XNOR2_X1 U25922 ( .A(n15606), .B(n16372), .ZN(n17645) );
  INV_X1 U25923 ( .A(n17645), .ZN(n16247) );
  XNOR2_X1 U25924 ( .A(n15212), .B(n16247), .ZN(n18216) );
  XNOR2_X1 U25925 ( .A(n23370), .B(n49429), .ZN(n24443) );
  XNOR2_X1 U25926 ( .A(n15213), .B(n24443), .ZN(n45380) );
  XNOR2_X1 U25927 ( .A(n45380), .B(n4208), .ZN(n24723) );
  XNOR2_X1 U25928 ( .A(n24723), .B(n24057), .ZN(n34346) );
  XNOR2_X1 U25929 ( .A(n17365), .B(n34346), .ZN(n15217) );
  XNOR2_X1 U25930 ( .A(n43691), .B(n4939), .ZN(n15214) );
  XNOR2_X1 U25931 ( .A(n28304), .B(n15214), .ZN(n33625) );
  XNOR2_X1 U25932 ( .A(n33625), .B(n47737), .ZN(n15215) );
  XNOR2_X1 U25933 ( .A(n15217), .B(n15216), .ZN(n15219) );
  XNOR2_X1 U25934 ( .A(n15677), .B(n16904), .ZN(n15218) );
  XNOR2_X1 U25935 ( .A(n15218), .B(n485), .ZN(n15754) );
  XNOR2_X1 U25936 ( .A(n15754), .B(n15219), .ZN(n15223) );
  XNOR2_X1 U25937 ( .A(n18643), .B(n18791), .ZN(n15221) );
  XNOR2_X1 U25938 ( .A(n15221), .B(n15220), .ZN(n17944) );
  INV_X1 U25939 ( .A(n17944), .ZN(n15222) );
  XNOR2_X1 U25940 ( .A(n15223), .B(n15222), .ZN(n15224) );
  XNOR2_X1 U25941 ( .A(n16620), .B(n2214), .ZN(n15225) );
  XNOR2_X1 U25942 ( .A(n18169), .B(n17145), .ZN(n15478) );
  XNOR2_X1 U25943 ( .A(n15478), .B(n15225), .ZN(n16342) );
  XNOR2_X1 U25945 ( .A(n4639), .B(n3383), .ZN(n25795) );
  XNOR2_X1 U25946 ( .A(n25795), .B(n26297), .ZN(n15226) );
  XNOR2_X1 U25947 ( .A(n15226), .B(n25040), .ZN(n17716) );
  INV_X1 U25948 ( .A(n17716), .ZN(n16737) );
  XNOR2_X1 U25949 ( .A(n27483), .B(n2947), .ZN(n16608) );
  XNOR2_X1 U25950 ( .A(n16737), .B(n16608), .ZN(n42620) );
  XNOR2_X1 U25951 ( .A(n42620), .B(n25718), .ZN(n35766) );
  XNOR2_X1 U25952 ( .A(n42769), .B(n4035), .ZN(n18172) );
  XNOR2_X1 U25953 ( .A(n4482), .B(n4515), .ZN(n15227) );
  XNOR2_X1 U25954 ( .A(n18172), .B(n15227), .ZN(n15228) );
  XNOR2_X1 U25955 ( .A(n44193), .B(n15228), .ZN(n35130) );
  XNOR2_X1 U25956 ( .A(n35766), .B(n35130), .ZN(n15229) );
  XNOR2_X1 U25958 ( .A(n15231), .B(n19227), .ZN(n15232) );
  XNOR2_X1 U25959 ( .A(n16342), .B(n15232), .ZN(n15272) );
  OAI21_X1 U25960 ( .B1(n15235), .B2(n15234), .A(n15233), .ZN(n15238) );
  NAND3_X1 U25961 ( .A1(n15238), .A2(n15237), .A3(n15236), .ZN(n15239) );
  OAI21_X1 U25962 ( .B1(n15241), .B2(n15240), .A(n15239), .ZN(n15247) );
  NAND4_X1 U25963 ( .A1(n15245), .A2(n15244), .A3(n15243), .A4(n15242), .ZN(
        n15246) );
  XNOR2_X1 U25964 ( .A(n17322), .B(n16416), .ZN(n17914) );
  XNOR2_X1 U25965 ( .A(n51031), .B(n17914), .ZN(n18660) );
  INV_X1 U25966 ( .A(n15251), .ZN(n15252) );
  AOI22_X1 U25967 ( .A1(n15254), .A2(n15253), .B1(n15252), .B2(n15256), .ZN(
        n15270) );
  INV_X1 U25968 ( .A(n15255), .ZN(n15258) );
  OAI211_X1 U25969 ( .C1(n15259), .C2(n15258), .A(n15257), .B(n15256), .ZN(
        n15262) );
  AND2_X1 U25970 ( .A1(n15262), .A2(n15261), .ZN(n15269) );
  NAND2_X1 U25971 ( .A1(n15266), .A2(n15265), .ZN(n15267) );
  XNOR2_X1 U25972 ( .A(n51047), .B(n16973), .ZN(n16259) );
  XNOR2_X1 U25973 ( .A(n18660), .B(n16259), .ZN(n15271) );
  INV_X1 U25975 ( .A(n15273), .ZN(n15277) );
  NAND2_X1 U25976 ( .A1(n15274), .A2(n15279), .ZN(n15276) );
  OAI211_X1 U25977 ( .C1(n51500), .C2(n15277), .A(n15276), .B(n51724), .ZN(
        n15291) );
  AND2_X1 U25978 ( .A1(n15279), .A2(n15278), .ZN(n15282) );
  INV_X1 U25979 ( .A(n15280), .ZN(n15281) );
  OAI21_X1 U25980 ( .B1(n15283), .B2(n15282), .A(n15281), .ZN(n15290) );
  NOR2_X1 U25981 ( .A1(n15285), .A2(n51500), .ZN(n15287) );
  NAND2_X1 U25982 ( .A1(n15287), .A2(n15286), .ZN(n15289) );
  XNOR2_X1 U25984 ( .A(n16658), .B(n18696), .ZN(n15292) );
  XNOR2_X1 U25985 ( .A(n15292), .B(n16568), .ZN(n18130) );
  XNOR2_X1 U25986 ( .A(n17730), .B(n18690), .ZN(n15293) );
  XNOR2_X1 U25987 ( .A(n15295), .B(n17731), .ZN(n15296) );
  XNOR2_X1 U25988 ( .A(n15297), .B(n15296), .ZN(n15540) );
  XNOR2_X1 U25989 ( .A(n15540), .B(n18130), .ZN(n15320) );
  INV_X1 U25990 ( .A(n15298), .ZN(n15301) );
  AND2_X1 U25991 ( .A1(n15304), .A2(n15303), .ZN(n15312) );
  NAND2_X1 U25992 ( .A1(n15307), .A2(n1486), .ZN(n15308) );
  NOR2_X1 U25993 ( .A1(n15308), .A2(n15766), .ZN(n15768) );
  NAND2_X1 U25994 ( .A1(n15768), .A2(n15309), .ZN(n15310) );
  XNOR2_X1 U25995 ( .A(n16770), .B(n51014), .ZN(n17738) );
  XNOR2_X1 U25996 ( .A(n28085), .B(n40104), .ZN(n33589) );
  INV_X1 U25997 ( .A(n31432), .ZN(n42297) );
  XNOR2_X1 U25998 ( .A(n33589), .B(n42297), .ZN(n17728) );
  INV_X1 U25999 ( .A(n17728), .ZN(n24942) );
  XNOR2_X1 U26000 ( .A(n24942), .B(n4502), .ZN(n35055) );
  XNOR2_X1 U26001 ( .A(n48814), .B(n49109), .ZN(n43073) );
  XNOR2_X1 U26002 ( .A(n43073), .B(n42322), .ZN(n17180) );
  XNOR2_X1 U26003 ( .A(n17180), .B(n6031), .ZN(n35052) );
  XNOR2_X1 U26004 ( .A(n42889), .B(n4835), .ZN(n17844) );
  XNOR2_X1 U26005 ( .A(n17844), .B(n4845), .ZN(n35780) );
  XNOR2_X1 U26006 ( .A(n35052), .B(n35780), .ZN(n15314) );
  XNOR2_X1 U26007 ( .A(n35055), .B(n15314), .ZN(n15315) );
  XNOR2_X1 U26008 ( .A(n19185), .B(n15315), .ZN(n15316) );
  XNOR2_X1 U26009 ( .A(n15317), .B(n15316), .ZN(n15318) );
  XNOR2_X1 U26010 ( .A(n17738), .B(n15318), .ZN(n15319) );
  XNOR2_X1 U26011 ( .A(n17754), .B(n15321), .ZN(n15349) );
  INV_X1 U26012 ( .A(n15444), .ZN(n15322) );
  OAI21_X1 U26013 ( .B1(n15440), .B2(n15323), .A(n15322), .ZN(n15330) );
  NAND2_X1 U26014 ( .A1(n15326), .A2(n15440), .ZN(n15327) );
  NAND2_X1 U26015 ( .A1(n15438), .A2(n15440), .ZN(n15331) );
  NOR2_X1 U26016 ( .A1(n15332), .A2(n15331), .ZN(n15333) );
  OAI21_X1 U26017 ( .B1(n15333), .B2(n15443), .A(n15335), .ZN(n15347) );
  NAND2_X1 U26018 ( .A1(n15434), .A2(n15438), .ZN(n15336) );
  OAI22_X1 U26019 ( .A1(n15339), .A2(n15338), .B1(n51700), .B2(n15336), .ZN(
        n15340) );
  NAND2_X1 U26020 ( .A1(n15340), .A2(n15437), .ZN(n15346) );
  NAND3_X1 U26021 ( .A1(n15344), .A2(n15343), .A3(n15438), .ZN(n15345) );
  XNOR2_X1 U26022 ( .A(n543), .B(n15349), .ZN(n17705) );
  XNOR2_X1 U26023 ( .A(n2599), .B(n41825), .ZN(n43202) );
  XNOR2_X1 U26024 ( .A(n43202), .B(n1224), .ZN(n25555) );
  XNOR2_X1 U26025 ( .A(n33429), .B(n4565), .ZN(n26561) );
  XNOR2_X1 U26026 ( .A(n26561), .B(n4885), .ZN(n37140) );
  XNOR2_X1 U26027 ( .A(n25555), .B(n37140), .ZN(n15351) );
  XNOR2_X1 U26028 ( .A(n43368), .B(n35107), .ZN(n33050) );
  XNOR2_X1 U26029 ( .A(n33050), .B(n45106), .ZN(n27205) );
  XNOR2_X1 U26031 ( .A(n22814), .B(n42816), .ZN(n28058) );
  INV_X1 U26032 ( .A(n28058), .ZN(n15350) );
  XNOR2_X1 U26033 ( .A(n27205), .B(n15350), .ZN(n36741) );
  XNOR2_X1 U26034 ( .A(n15351), .B(n36741), .ZN(n15352) );
  XNOR2_X1 U26035 ( .A(n17891), .B(n15352), .ZN(n15353) );
  XNOR2_X1 U26036 ( .A(n15353), .B(n14903), .ZN(n15354) );
  XNOR2_X1 U26037 ( .A(n15355), .B(n15354), .ZN(n15356) );
  XNOR2_X1 U26038 ( .A(n15356), .B(n17705), .ZN(n15397) );
  XNOR2_X1 U26039 ( .A(n17879), .B(n16628), .ZN(n17343) );
  INV_X1 U26040 ( .A(n15357), .ZN(n15360) );
  NAND3_X1 U26041 ( .A1(n15360), .A2(n15359), .A3(n15358), .ZN(n15361) );
  OAI211_X1 U26042 ( .C1(n15363), .C2(n15376), .A(n15362), .B(n15361), .ZN(
        n15371) );
  INV_X1 U26043 ( .A(n15364), .ZN(n15369) );
  NAND2_X1 U26044 ( .A1(n15365), .A2(n15385), .ZN(n15379) );
  NAND3_X1 U26045 ( .A1(n15366), .A2(n15386), .A3(n15379), .ZN(n15368) );
  OAI211_X1 U26046 ( .C1(n15382), .C2(n15369), .A(n15368), .B(n15367), .ZN(
        n15370) );
  INV_X1 U26047 ( .A(n15372), .ZN(n15373) );
  NAND3_X1 U26048 ( .A1(n15374), .A2(n15380), .A3(n15373), .ZN(n15392) );
  INV_X1 U26049 ( .A(n15375), .ZN(n15377) );
  INV_X1 U26050 ( .A(n15379), .ZN(n15383) );
  NAND4_X1 U26051 ( .A1(n15383), .A2(n15382), .A3(n15381), .A4(n15380), .ZN(
        n15388) );
  NAND3_X1 U26052 ( .A1(n15386), .A2(n15385), .A3(n15384), .ZN(n15387) );
  AND2_X1 U26053 ( .A1(n15388), .A2(n15387), .ZN(n15390) );
  NAND4_X1 U26054 ( .A1(n15392), .A2(n15391), .A3(n15390), .A4(n15389), .ZN(
        n15393) );
  XNOR2_X1 U26055 ( .A(n17758), .B(n2134), .ZN(n18163) );
  XNOR2_X1 U26056 ( .A(n18163), .B(n17343), .ZN(n16732) );
  XNOR2_X1 U26057 ( .A(n18668), .B(n14427), .ZN(n15395) );
  XNOR2_X1 U26058 ( .A(n15396), .B(n15395), .ZN(n15467) );
  INV_X1 U26059 ( .A(n15399), .ZN(n19410) );
  AND2_X1 U26060 ( .A1(n18039), .A2(n19410), .ZN(n19413) );
  INV_X1 U26061 ( .A(n17869), .ZN(n19418) );
  INV_X1 U26062 ( .A(n19424), .ZN(n18037) );
  NAND2_X1 U26063 ( .A1(n18040), .A2(n15399), .ZN(n18033) );
  INV_X1 U26064 ( .A(n18033), .ZN(n17872) );
  NAND2_X1 U26065 ( .A1(n18037), .A2(n17872), .ZN(n15401) );
  XNOR2_X1 U26067 ( .A(n23882), .B(n26178), .ZN(n16385) );
  XNOR2_X1 U26068 ( .A(n36941), .B(n4667), .ZN(n35034) );
  XNOR2_X1 U26069 ( .A(n16385), .B(n35034), .ZN(n24495) );
  XNOR2_X2 U26070 ( .A(n4908), .B(n4754), .ZN(n43739) );
  XNOR2_X1 U26071 ( .A(n45736), .B(n4897), .ZN(n23495) );
  XNOR2_X1 U26072 ( .A(n43739), .B(n23495), .ZN(n24612) );
  INV_X1 U26073 ( .A(n24612), .ZN(n15404) );
  XNOR2_X1 U26074 ( .A(n24495), .B(n15404), .ZN(n22218) );
  XNOR2_X1 U26075 ( .A(n4869), .B(n4712), .ZN(n33181) );
  XNOR2_X1 U26076 ( .A(n22218), .B(n33181), .ZN(n33821) );
  XNOR2_X1 U26077 ( .A(n28070), .B(n4788), .ZN(n15405) );
  XNOR2_X1 U26078 ( .A(n24932), .B(n15405), .ZN(n34003) );
  XNOR2_X1 U26079 ( .A(n33821), .B(n34003), .ZN(n15406) );
  XNOR2_X1 U26080 ( .A(n18599), .B(n15406), .ZN(n15407) );
  XNOR2_X1 U26081 ( .A(n15407), .B(n18712), .ZN(n15408) );
  XNOR2_X1 U26082 ( .A(n15409), .B(n15408), .ZN(n15411) );
  XNOR2_X1 U26083 ( .A(n15410), .B(n18714), .ZN(n19271) );
  XNOR2_X1 U26084 ( .A(n19271), .B(n15411), .ZN(n15457) );
  XNOR2_X1 U26085 ( .A(n18749), .B(n18134), .ZN(n15491) );
  OR2_X1 U26086 ( .A1(n15417), .A2(n15424), .ZN(n15413) );
  OAI211_X1 U26087 ( .C1(n15414), .C2(n1555), .A(n15413), .B(n15412), .ZN(
        n15415) );
  INV_X1 U26088 ( .A(n15415), .ZN(n15430) );
  INV_X1 U26089 ( .A(n15416), .ZN(n15420) );
  NAND2_X1 U26090 ( .A1(n15417), .A2(n2249), .ZN(n15418) );
  AOI22_X1 U26091 ( .A1(n15421), .A2(n15420), .B1(n51023), .B2(n15418), .ZN(
        n15429) );
  NAND2_X1 U26092 ( .A1(n15427), .A2(n15426), .ZN(n15428) );
  NAND2_X1 U26093 ( .A1(n15431), .A2(n15437), .ZN(n15432) );
  AND2_X1 U26094 ( .A1(n15433), .A2(n15432), .ZN(n15453) );
  XNOR2_X1 U26095 ( .A(n15435), .B(n15434), .ZN(n15441) );
  OAI211_X1 U26096 ( .C1(n15441), .C2(n15440), .A(n15439), .B(n15438), .ZN(
        n15452) );
  OAI21_X1 U26097 ( .B1(n15444), .B2(n15443), .A(n15442), .ZN(n15451) );
  OAI21_X1 U26098 ( .B1(n15447), .B2(n15446), .A(n15445), .ZN(n15449) );
  NAND2_X1 U26099 ( .A1(n15449), .A2(n15448), .ZN(n15450) );
  XNOR2_X2 U26100 ( .A(n17288), .B(n17169), .ZN(n18457) );
  XNOR2_X1 U26101 ( .A(n15491), .B(n18591), .ZN(n15455) );
  XNOR2_X1 U26102 ( .A(n17694), .B(n15455), .ZN(n15456) );
  NOR2_X1 U26105 ( .A1(n17869), .A2(n17871), .ZN(n19422) );
  NAND2_X1 U26106 ( .A1(n17557), .A2(n18033), .ZN(n15459) );
  OAI211_X1 U26107 ( .C1(n19422), .C2(n15459), .A(n18041), .B(n18043), .ZN(
        n15463) );
  NOR2_X1 U26108 ( .A1(n18034), .A2(n18041), .ZN(n15460) );
  AOI22_X1 U26109 ( .A1(n15460), .A2(n19424), .B1(n18039), .B2(n19404), .ZN(
        n15462) );
  NAND2_X1 U26110 ( .A1(n18034), .A2(n17871), .ZN(n17558) );
  AND4_X1 U26111 ( .A1(n15463), .A2(n15462), .A3(n19408), .A4(n15461), .ZN(
        n15464) );
  XNOR2_X1 U26112 ( .A(n16412), .B(n51668), .ZN(n15466) );
  XNOR2_X1 U26113 ( .A(n15466), .B(n52194), .ZN(n16328) );
  XNOR2_X1 U26114 ( .A(n15468), .B(n15467), .ZN(n15476) );
  XNOR2_X1 U26115 ( .A(n34414), .B(n45107), .ZN(n33297) );
  INV_X1 U26116 ( .A(n33297), .ZN(n42366) );
  XNOR2_X1 U26117 ( .A(n42592), .B(n42366), .ZN(n43153) );
  XOR2_X1 U26118 ( .A(n4638), .B(n4501), .Z(n15469) );
  XNOR2_X1 U26119 ( .A(n1224), .B(n4868), .ZN(n43200) );
  XNOR2_X1 U26120 ( .A(n15469), .B(n43200), .ZN(n15470) );
  XNOR2_X1 U26121 ( .A(n43153), .B(n15470), .ZN(n15471) );
  XNOR2_X1 U26122 ( .A(n18147), .B(n15471), .ZN(n15472) );
  XNOR2_X1 U26123 ( .A(n15474), .B(n15473), .ZN(n15475) );
  XNOR2_X1 U26124 ( .A(n15476), .B(n15475), .ZN(n15477) );
  XNOR2_X1 U26125 ( .A(n461), .B(n16620), .ZN(n15479) );
  XNOR2_X1 U26126 ( .A(n15478), .B(n15479), .ZN(n15485) );
  XNOR2_X1 U26127 ( .A(n24430), .B(n38626), .ZN(n24227) );
  XNOR2_X1 U26128 ( .A(n25575), .B(n24227), .ZN(n26368) );
  INV_X1 U26129 ( .A(n16739), .ZN(n15480) );
  XNOR2_X1 U26130 ( .A(n15480), .B(n33653), .ZN(n24692) );
  XNOR2_X1 U26131 ( .A(n26368), .B(n24692), .ZN(n32807) );
  XNOR2_X1 U26132 ( .A(n4296), .B(n2947), .ZN(n16977) );
  XNOR2_X1 U26133 ( .A(n25040), .B(n16977), .ZN(n25993) );
  XNOR2_X1 U26134 ( .A(n274), .B(n4705), .ZN(n17317) );
  XNOR2_X1 U26135 ( .A(n25993), .B(n17317), .ZN(n37314) );
  XNOR2_X1 U26136 ( .A(n32807), .B(n37314), .ZN(n15481) );
  XNOR2_X1 U26137 ( .A(n16162), .B(n15481), .ZN(n15482) );
  XNOR2_X1 U26138 ( .A(n15482), .B(n2214), .ZN(n15483) );
  XNOR2_X1 U26139 ( .A(n15483), .B(n16330), .ZN(n15484) );
  XNOR2_X1 U26140 ( .A(n15484), .B(n15485), .ZN(n15490) );
  XNOR2_X1 U26141 ( .A(n15642), .B(n15486), .ZN(n15488) );
  XNOR2_X1 U26142 ( .A(n18175), .B(n4415), .ZN(n15487) );
  XNOR2_X1 U26143 ( .A(n18181), .B(n15487), .ZN(n17722) );
  XNOR2_X1 U26144 ( .A(n15488), .B(n17722), .ZN(n15489) );
  XNOR2_X1 U26145 ( .A(n15491), .B(n18714), .ZN(n15503) );
  XNOR2_X1 U26146 ( .A(n23887), .B(n4869), .ZN(n24748) );
  XNOR2_X1 U26147 ( .A(n24748), .B(n15492), .ZN(n34233) );
  XNOR2_X1 U26148 ( .A(n34233), .B(n4897), .ZN(n27470) );
  XNOR2_X1 U26149 ( .A(n4836), .B(n4916), .ZN(n15493) );
  XNOR2_X1 U26150 ( .A(n26604), .B(n15493), .ZN(n15494) );
  XNOR2_X1 U26151 ( .A(n15494), .B(n23882), .ZN(n33422) );
  XNOR2_X1 U26152 ( .A(n33422), .B(n4788), .ZN(n15495) );
  XNOR2_X1 U26153 ( .A(n27470), .B(n15495), .ZN(n15496) );
  XNOR2_X1 U26154 ( .A(n17691), .B(n15496), .ZN(n15497) );
  XNOR2_X1 U26155 ( .A(n15498), .B(n15497), .ZN(n15501) );
  XNOR2_X1 U26156 ( .A(n17690), .B(n51134), .ZN(n15499) );
  XNOR2_X1 U26157 ( .A(n560), .B(n15499), .ZN(n15500) );
  XNOR2_X1 U26158 ( .A(n15501), .B(n15500), .ZN(n15502) );
  XNOR2_X1 U26159 ( .A(n15503), .B(n15502), .ZN(n15506) );
  XNOR2_X1 U26161 ( .A(n17944), .B(n15754), .ZN(n15514) );
  XNOR2_X1 U26162 ( .A(n17364), .B(n17812), .ZN(n15510) );
  XNOR2_X1 U26163 ( .A(n4939), .B(n49323), .ZN(n35796) );
  XNOR2_X1 U26164 ( .A(n36698), .B(n35796), .ZN(n17932) );
  XNOR2_X1 U26165 ( .A(n17932), .B(n33388), .ZN(n24055) );
  XNOR2_X1 U26166 ( .A(n24055), .B(n28304), .ZN(n33720) );
  XNOR2_X1 U26167 ( .A(n34575), .B(n43968), .ZN(n15507) );
  XNOR2_X1 U26168 ( .A(n33720), .B(n15507), .ZN(n15508) );
  XNOR2_X1 U26169 ( .A(n17118), .B(n15508), .ZN(n15509) );
  XNOR2_X1 U26170 ( .A(n15509), .B(n15510), .ZN(n15512) );
  XNOR2_X1 U26171 ( .A(n15512), .B(n15511), .ZN(n15513) );
  XNOR2_X1 U26172 ( .A(n43662), .B(n3014), .ZN(n34570) );
  XNOR2_X1 U26173 ( .A(n16532), .B(n15515), .ZN(n15516) );
  XNOR2_X1 U26174 ( .A(n15518), .B(n15517), .ZN(n17372) );
  XNOR2_X1 U26175 ( .A(n15519), .B(n16920), .ZN(n15520) );
  XNOR2_X1 U26176 ( .A(n15520), .B(n16527), .ZN(n18817) );
  INV_X1 U26177 ( .A(n18817), .ZN(n15531) );
  INV_X1 U26178 ( .A(n15689), .ZN(n15529) );
  XNOR2_X1 U26179 ( .A(n18437), .B(n51642), .ZN(n15527) );
  XNOR2_X1 U26180 ( .A(n4826), .B(n4286), .ZN(n15691) );
  XNOR2_X1 U26181 ( .A(n15691), .B(n15521), .ZN(n25436) );
  XNOR2_X1 U26182 ( .A(n25436), .B(n4287), .ZN(n15522) );
  XNOR2_X1 U26183 ( .A(n15522), .B(n42721), .ZN(n15524) );
  XNOR2_X1 U26184 ( .A(n4890), .B(n4612), .ZN(n25901) );
  XNOR2_X1 U26185 ( .A(n25901), .B(n35815), .ZN(n18191) );
  XNOR2_X1 U26186 ( .A(n16149), .B(n4781), .ZN(n24626) );
  XNOR2_X1 U26187 ( .A(n18191), .B(n24626), .ZN(n15523) );
  XNOR2_X1 U26188 ( .A(n15524), .B(n15523), .ZN(n33373) );
  XNOR2_X1 U26189 ( .A(n33373), .B(n34265), .ZN(n15525) );
  XNOR2_X1 U26190 ( .A(n16450), .B(n15525), .ZN(n15526) );
  XNOR2_X1 U26191 ( .A(n15527), .B(n15526), .ZN(n15528) );
  XNOR2_X1 U26192 ( .A(n15529), .B(n15528), .ZN(n15530) );
  XNOR2_X1 U26193 ( .A(n15531), .B(n15530), .ZN(n15534) );
  XNOR2_X1 U26194 ( .A(n16023), .B(n16923), .ZN(n17678) );
  XNOR2_X1 U26195 ( .A(n17798), .B(n17678), .ZN(n15532) );
  XNOR2_X1 U26196 ( .A(n17786), .B(n4837), .ZN(n17265) );
  XNOR2_X1 U26197 ( .A(n18615), .B(n17265), .ZN(n17349) );
  XNOR2_X1 U26198 ( .A(n15532), .B(n17349), .ZN(n15533) );
  NAND2_X1 U26199 ( .A1(n15535), .A2(n20512), .ZN(n15551) );
  INV_X1 U26200 ( .A(n15551), .ZN(n15550) );
  NAND2_X1 U26201 ( .A1(n20504), .A2(n20501), .ZN(n18082) );
  XNOR2_X1 U26202 ( .A(n24992), .B(n4827), .ZN(n32520) );
  XNOR2_X1 U26203 ( .A(n16943), .B(n32520), .ZN(n17725) );
  XNOR2_X1 U26204 ( .A(n16183), .B(n17725), .ZN(n15539) );
  XNOR2_X1 U26205 ( .A(n18689), .B(n51703), .ZN(n15537) );
  XNOR2_X1 U26206 ( .A(n15537), .B(n15536), .ZN(n15538) );
  XNOR2_X1 U26207 ( .A(n15539), .B(n15538), .ZN(n15541) );
  XNOR2_X1 U26208 ( .A(n33474), .B(n27297), .ZN(n25866) );
  XNOR2_X1 U26209 ( .A(n25866), .B(n4845), .ZN(n24941) );
  XNOR2_X1 U26210 ( .A(n24941), .B(n27299), .ZN(n43592) );
  XNOR2_X1 U26211 ( .A(n40104), .B(n4737), .ZN(n15543) );
  XNOR2_X1 U26212 ( .A(n43592), .B(n15543), .ZN(n15544) );
  XNOR2_X1 U26213 ( .A(n17280), .B(n15544), .ZN(n15545) );
  XNOR2_X1 U26214 ( .A(n15545), .B(n16294), .ZN(n15546) );
  XNOR2_X1 U26215 ( .A(n16781), .B(n15546), .ZN(n15547) );
  XNOR2_X1 U26216 ( .A(n15547), .B(n16438), .ZN(n15548) );
  AND2_X1 U26217 ( .A1(n18082), .A2(n19344), .ZN(n15549) );
  INV_X1 U26218 ( .A(n20513), .ZN(n19337) );
  NAND2_X1 U26219 ( .A1(n15551), .A2(n19337), .ZN(n15552) );
  INV_X1 U26220 ( .A(n20507), .ZN(n17625) );
  NOR2_X1 U26221 ( .A1(n18085), .A2(n1517), .ZN(n15554) );
  OAI21_X1 U26222 ( .B1(n17625), .B2(n15554), .A(n18086), .ZN(n15557) );
  OAI22_X1 U26223 ( .A1(n20512), .A2(n20514), .B1(n17619), .B2(n4516), .ZN(
        n15555) );
  AND2_X1 U26224 ( .A1(n51704), .A2(n20501), .ZN(n18075) );
  NAND2_X1 U26225 ( .A1(n15555), .A2(n18075), .ZN(n15556) );
  INV_X1 U26226 ( .A(n20534), .ZN(n22288) );
  AOI21_X1 U26227 ( .B1(n22288), .B2(n20948), .A(n21114), .ZN(n15560) );
  NAND2_X1 U26228 ( .A1(n21782), .A2(n24452), .ZN(n20944) );
  NAND2_X1 U26229 ( .A1(n20942), .A2(n22701), .ZN(n21116) );
  NOR2_X1 U26230 ( .A1(n20944), .A2(n21116), .ZN(n20531) );
  INV_X1 U26231 ( .A(n20531), .ZN(n15559) );
  NAND2_X1 U26232 ( .A1(n22702), .A2(n22287), .ZN(n21777) );
  INV_X1 U26233 ( .A(n20948), .ZN(n22284) );
  OAI21_X1 U26234 ( .B1(n51695), .B2(n22287), .A(n22284), .ZN(n15561) );
  AOI21_X1 U26235 ( .B1(n21777), .B2(n15561), .A(n22703), .ZN(n15562) );
  XNOR2_X1 U26236 ( .A(n42101), .B(n4587), .ZN(n36739) );
  XNOR2_X1 U26237 ( .A(n51436), .B(n36739), .ZN(n17331) );
  INV_X1 U26238 ( .A(n15563), .ZN(n16118) );
  XNOR2_X1 U26239 ( .A(n17331), .B(n16118), .ZN(n15567) );
  XNOR2_X1 U26240 ( .A(n36737), .B(n2608), .ZN(n15564) );
  XNOR2_X1 U26241 ( .A(n17232), .B(n15564), .ZN(n15565) );
  XNOR2_X1 U26243 ( .A(n15565), .B(n18505), .ZN(n16956) );
  INV_X1 U26244 ( .A(n16956), .ZN(n15566) );
  XNOR2_X1 U26245 ( .A(n15567), .B(n15566), .ZN(n15573) );
  XNOR2_X1 U26246 ( .A(n14427), .B(n17763), .ZN(n15568) );
  XNOR2_X1 U26247 ( .A(n15568), .B(n18407), .ZN(n15847) );
  INV_X1 U26248 ( .A(n35107), .ZN(n15569) );
  XNOR2_X1 U26249 ( .A(n25470), .B(n15569), .ZN(n43654) );
  XNOR2_X1 U26250 ( .A(n43654), .B(n4451), .ZN(n35654) );
  XNOR2_X1 U26251 ( .A(n4883), .B(n4579), .ZN(n35108) );
  XNOR2_X1 U26252 ( .A(n41155), .B(n35108), .ZN(n31131) );
  XNOR2_X1 U26253 ( .A(n35654), .B(n31131), .ZN(n15570) );
  XNOR2_X1 U26254 ( .A(n2135), .B(n15570), .ZN(n15571) );
  XNOR2_X1 U26255 ( .A(n15847), .B(n15571), .ZN(n15572) );
  XNOR2_X1 U26256 ( .A(n15573), .B(n15572), .ZN(n15574) );
  XNOR2_X1 U26257 ( .A(n15649), .B(n4847), .ZN(n15576) );
  XNOR2_X1 U26258 ( .A(n15576), .B(n16416), .ZN(n16098) );
  XNOR2_X1 U26259 ( .A(n15577), .B(n18540), .ZN(n15578) );
  XNOR2_X1 U26260 ( .A(n15578), .B(n17145), .ZN(n16418) );
  XNOR2_X1 U26261 ( .A(n15579), .B(n16973), .ZN(n15808) );
  INV_X1 U26262 ( .A(n15808), .ZN(n15585) );
  XNOR2_X1 U26263 ( .A(n24229), .B(n25114), .ZN(n17148) );
  XNOR2_X1 U26264 ( .A(n25795), .B(n41567), .ZN(n26296) );
  XNOR2_X1 U26265 ( .A(n26296), .B(n4296), .ZN(n18528) );
  XNOR2_X1 U26266 ( .A(n17148), .B(n18528), .ZN(n44921) );
  XOR2_X1 U26267 ( .A(n4454), .B(n4931), .Z(n15580) );
  XNOR2_X1 U26268 ( .A(n15580), .B(n26541), .ZN(n35765) );
  XNOR2_X1 U26269 ( .A(n44921), .B(n35765), .ZN(n15581) );
  XNOR2_X1 U26270 ( .A(n461), .B(n15581), .ZN(n15583) );
  XNOR2_X1 U26271 ( .A(n15583), .B(n15582), .ZN(n15584) );
  XNOR2_X1 U26272 ( .A(n15585), .B(n15584), .ZN(n15586) );
  XNOR2_X1 U26273 ( .A(n32856), .B(n2603), .ZN(n27351) );
  XNOR2_X1 U26274 ( .A(n27351), .B(n34265), .ZN(n15587) );
  XNOR2_X1 U26275 ( .A(n15587), .B(n33374), .ZN(n24313) );
  XNOR2_X1 U26276 ( .A(n34027), .B(n49937), .ZN(n15588) );
  XNOR2_X1 U26277 ( .A(n33845), .B(n15588), .ZN(n15589) );
  XNOR2_X1 U26278 ( .A(n23943), .B(n4636), .ZN(n43850) );
  XNOR2_X1 U26279 ( .A(n15589), .B(n43850), .ZN(n15590) );
  XNOR2_X1 U26280 ( .A(n24313), .B(n15590), .ZN(n15591) );
  XNOR2_X1 U26281 ( .A(n16017), .B(n15591), .ZN(n15592) );
  XNOR2_X1 U26282 ( .A(n15592), .B(n51482), .ZN(n15595) );
  XNOR2_X1 U26283 ( .A(n17258), .B(n4826), .ZN(n18546) );
  XNOR2_X1 U26284 ( .A(n16011), .B(n18432), .ZN(n15596) );
  XNOR2_X1 U26285 ( .A(n17348), .B(n15596), .ZN(n15598) );
  XNOR2_X1 U26286 ( .A(n16913), .B(n18448), .ZN(n15597) );
  XNOR2_X1 U26287 ( .A(n15598), .B(n15597), .ZN(n16520) );
  XNOR2_X1 U26288 ( .A(n15599), .B(n16520), .ZN(n15601) );
  XNOR2_X1 U26289 ( .A(n49429), .B(Key[98]), .ZN(n16241) );
  XNOR2_X1 U26290 ( .A(n34575), .B(n16241), .ZN(n17121) );
  XNOR2_X1 U26291 ( .A(n17121), .B(n4932), .ZN(n25208) );
  XNOR2_X1 U26292 ( .A(n43293), .B(n3336), .ZN(n25078) );
  XNOR2_X1 U26293 ( .A(n25208), .B(n25078), .ZN(n33627) );
  XNOR2_X1 U26294 ( .A(n25147), .B(n26042), .ZN(n26387) );
  XNOR2_X1 U26295 ( .A(n26387), .B(n48597), .ZN(n34345) );
  XNOR2_X1 U26296 ( .A(n43968), .B(n4817), .ZN(n15602) );
  XNOR2_X1 U26297 ( .A(n34345), .B(n15602), .ZN(n15603) );
  INV_X1 U26298 ( .A(n17803), .ZN(n16028) );
  XNOR2_X1 U26299 ( .A(n15604), .B(n2225), .ZN(n15605) );
  XNOR2_X1 U26300 ( .A(n16464), .B(n17117), .ZN(n16582) );
  XNOR2_X1 U26301 ( .A(n16582), .B(n18791), .ZN(n16896) );
  XNOR2_X1 U26302 ( .A(n15606), .B(n18644), .ZN(n16907) );
  XNOR2_X1 U26303 ( .A(n15607), .B(n16907), .ZN(n15608) );
  XNOR2_X1 U26304 ( .A(n16063), .B(n18457), .ZN(n15615) );
  XNOR2_X1 U26305 ( .A(n45350), .B(n4869), .ZN(n27317) );
  XNOR2_X1 U26306 ( .A(n44493), .B(n36941), .ZN(n16280) );
  XNOR2_X1 U26307 ( .A(n25616), .B(n4897), .ZN(n25168) );
  XNOR2_X1 U26308 ( .A(n16280), .B(n25168), .ZN(n15610) );
  XNOR2_X1 U26309 ( .A(n27317), .B(n15610), .ZN(n34002) );
  XNOR2_X1 U26310 ( .A(n28071), .B(n34709), .ZN(n23888) );
  XNOR2_X1 U26311 ( .A(n23888), .B(n4655), .ZN(n33822) );
  XNOR2_X1 U26312 ( .A(n33822), .B(n4908), .ZN(n15611) );
  XNOR2_X1 U26313 ( .A(n34002), .B(n15611), .ZN(n15612) );
  XNOR2_X1 U26314 ( .A(n18466), .B(n15612), .ZN(n15613) );
  XNOR2_X1 U26315 ( .A(n15613), .B(n356), .ZN(n15614) );
  XNOR2_X1 U26316 ( .A(n15615), .B(n15614), .ZN(n15616) );
  XNOR2_X1 U26317 ( .A(n15619), .B(n16660), .ZN(n15626) );
  XNOR2_X1 U26318 ( .A(n41460), .B(n43073), .ZN(n23773) );
  XNOR2_X1 U26319 ( .A(n23773), .B(n17181), .ZN(n35781) );
  INV_X1 U26320 ( .A(n4613), .ZN(n50463) );
  XNOR2_X1 U26321 ( .A(n26586), .B(n50463), .ZN(n18117) );
  INV_X1 U26322 ( .A(n18117), .ZN(n15622) );
  XNOR2_X1 U26323 ( .A(n4585), .B(n4471), .ZN(n15620) );
  XNOR2_X1 U26324 ( .A(n43105), .B(n15620), .ZN(n15621) );
  XNOR2_X1 U26325 ( .A(n15622), .B(n15621), .ZN(n35056) );
  XNOR2_X1 U26326 ( .A(n35056), .B(n4518), .ZN(n15623) );
  XNOR2_X1 U26327 ( .A(n35781), .B(n15623), .ZN(n15624) );
  XNOR2_X1 U26328 ( .A(n18119), .B(n15624), .ZN(n15625) );
  XNOR2_X1 U26329 ( .A(n15626), .B(n15625), .ZN(n15627) );
  XNOR2_X1 U26330 ( .A(n15628), .B(n51014), .ZN(n16950) );
  AND2_X1 U26331 ( .A1(n18942), .A2(n19636), .ZN(n19887) );
  NAND2_X1 U26333 ( .A1(n51127), .A2(n19662), .ZN(n19637) );
  INV_X1 U26334 ( .A(n19637), .ZN(n19670) );
  NAND3_X1 U26335 ( .A1(n19898), .A2(n18933), .A3(n19670), .ZN(n15638) );
  AND2_X1 U26336 ( .A1(n15630), .A2(n19892), .ZN(n19657) );
  INV_X1 U26337 ( .A(n19657), .ZN(n19660) );
  NAND2_X1 U26338 ( .A1(n19893), .A2(n19892), .ZN(n19897) );
  AOI21_X1 U26339 ( .B1(n19660), .B2(n19897), .A(n18942), .ZN(n15632) );
  NAND2_X1 U26340 ( .A1(n15633), .A2(n15632), .ZN(n15637) );
  NAND2_X1 U26341 ( .A1(n18932), .A2(n19889), .ZN(n15635) );
  NAND2_X1 U26342 ( .A1(n19891), .A2(n19636), .ZN(n18941) );
  NOR2_X1 U26343 ( .A1(n18941), .A2(n19894), .ZN(n18927) );
  NAND2_X1 U26344 ( .A1(n18927), .A2(n51127), .ZN(n15634) );
  INV_X1 U26345 ( .A(n19897), .ZN(n15636) );
  XNOR2_X1 U26346 ( .A(n2126), .B(n15640), .ZN(n17770) );
  XNOR2_X1 U26347 ( .A(n511), .B(n2181), .ZN(n15641) );
  XNOR2_X1 U26348 ( .A(n17770), .B(n15641), .ZN(n15643) );
  XNOR2_X1 U26349 ( .A(n18664), .B(n15643), .ZN(n15656) );
  XNOR2_X1 U26350 ( .A(n16739), .B(n4755), .ZN(n15644) );
  XNOR2_X1 U26351 ( .A(n15644), .B(n24430), .ZN(n24585) );
  XNOR2_X1 U26352 ( .A(n33653), .B(n26541), .ZN(n28412) );
  INV_X1 U26353 ( .A(n28412), .ZN(n15645) );
  XNOR2_X1 U26354 ( .A(n24585), .B(n15645), .ZN(n46065) );
  XNOR2_X1 U26355 ( .A(n46065), .B(n25042), .ZN(n35272) );
  XNOR2_X1 U26356 ( .A(n25114), .B(n29662), .ZN(n26295) );
  XNOR2_X1 U26357 ( .A(n26295), .B(n4296), .ZN(n35674) );
  XNOR2_X1 U26358 ( .A(n4706), .B(n4665), .ZN(n21091) );
  XNOR2_X1 U26359 ( .A(n21091), .B(n4847), .ZN(n15646) );
  XNOR2_X1 U26360 ( .A(n35674), .B(n15646), .ZN(n15647) );
  XNOR2_X1 U26361 ( .A(n35272), .B(n15647), .ZN(n15648) );
  XNOR2_X1 U26362 ( .A(n15649), .B(n15648), .ZN(n15651) );
  XNOR2_X1 U26363 ( .A(n15651), .B(n15650), .ZN(n15652) );
  XNOR2_X1 U26364 ( .A(n15957), .B(n17212), .ZN(n15859) );
  XNOR2_X1 U26365 ( .A(n15652), .B(n15859), .ZN(n15654) );
  XNOR2_X1 U26366 ( .A(n18181), .B(n15653), .ZN(n18543) );
  XNOR2_X1 U26367 ( .A(n15654), .B(n17161), .ZN(n15655) );
  XNOR2_X1 U26368 ( .A(n15656), .B(n15655), .ZN(n15725) );
  INV_X1 U26369 ( .A(n15725), .ZN(n18921) );
  XNOR2_X1 U26370 ( .A(n18147), .B(n18522), .ZN(n15657) );
  XNOR2_X1 U26371 ( .A(n15658), .B(n15657), .ZN(n15665) );
  XNOR2_X1 U26372 ( .A(n33429), .B(n44934), .ZN(n44046) );
  XNOR2_X1 U26373 ( .A(n35108), .B(n45883), .ZN(n15659) );
  XNOR2_X1 U26374 ( .A(n44046), .B(n15659), .ZN(n15660) );
  XNOR2_X1 U26375 ( .A(n34414), .B(n1224), .ZN(n26358) );
  XNOR2_X1 U26376 ( .A(n15660), .B(n26358), .ZN(n15661) );
  XNOR2_X1 U26377 ( .A(n18157), .B(n15661), .ZN(n15663) );
  XNOR2_X1 U26378 ( .A(n16628), .B(n17707), .ZN(n15662) );
  XNOR2_X1 U26379 ( .A(n15663), .B(n15662), .ZN(n15664) );
  XNOR2_X1 U26380 ( .A(n43019), .B(n34411), .ZN(n35376) );
  XNOR2_X1 U26381 ( .A(n16720), .B(n35376), .ZN(n15667) );
  XNOR2_X1 U26382 ( .A(n18414), .B(n15667), .ZN(n15669) );
  INV_X1 U26383 ( .A(n20210), .ZN(n19672) );
  XNOR2_X1 U26384 ( .A(n25744), .B(n3276), .ZN(n27454) );
  XNOR2_X1 U26385 ( .A(n27454), .B(n42077), .ZN(n19246) );
  INV_X1 U26386 ( .A(n19246), .ZN(n24638) );
  XNOR2_X1 U26387 ( .A(n35796), .B(n25147), .ZN(n15671) );
  INV_X1 U26388 ( .A(n27174), .ZN(n15670) );
  XNOR2_X1 U26389 ( .A(n15671), .B(n15670), .ZN(n17360) );
  XNOR2_X1 U26390 ( .A(n24638), .B(n17360), .ZN(n42657) );
  XNOR2_X1 U26391 ( .A(n43968), .B(n2903), .ZN(n33346) );
  XNOR2_X1 U26392 ( .A(n33346), .B(n4909), .ZN(n15672) );
  XNOR2_X1 U26393 ( .A(n42657), .B(n15672), .ZN(n15673) );
  XNOR2_X1 U26394 ( .A(n18795), .B(n15673), .ZN(n15674) );
  XNOR2_X1 U26395 ( .A(n16471), .B(n15674), .ZN(n15675) );
  XNOR2_X1 U26396 ( .A(n15675), .B(n17127), .ZN(n15676) );
  XNOR2_X1 U26397 ( .A(n52229), .B(n557), .ZN(n15940) );
  XNOR2_X1 U26398 ( .A(n15940), .B(n15676), .ZN(n15685) );
  XNOR2_X1 U26399 ( .A(n15678), .B(n15867), .ZN(n15679) );
  INV_X1 U26400 ( .A(n17814), .ZN(n18212) );
  XNOR2_X1 U26401 ( .A(n15679), .B(n18212), .ZN(n15684) );
  XNOR2_X1 U26402 ( .A(n15681), .B(n15680), .ZN(n15933) );
  INV_X1 U26403 ( .A(n15933), .ZN(n15683) );
  XNOR2_X1 U26404 ( .A(n15683), .B(n15682), .ZN(n17253) );
  XNOR2_X1 U26405 ( .A(n16228), .B(n16919), .ZN(n15686) );
  XNOR2_X1 U26406 ( .A(n15686), .B(n18443), .ZN(n15687) );
  XNOR2_X1 U26407 ( .A(n15687), .B(n51481), .ZN(n17261) );
  INV_X1 U26408 ( .A(n15688), .ZN(n18194) );
  XNOR2_X1 U26409 ( .A(n15689), .B(n18820), .ZN(n15690) );
  XNOR2_X1 U26410 ( .A(n15690), .B(n17261), .ZN(n15699) );
  XNOR2_X1 U26411 ( .A(n16011), .B(n51642), .ZN(n15694) );
  XNOR2_X1 U26412 ( .A(n18191), .B(n45050), .ZN(n25651) );
  XNOR2_X1 U26413 ( .A(n25651), .B(n34027), .ZN(n43564) );
  XNOR2_X1 U26414 ( .A(n43564), .B(n4649), .ZN(n26114) );
  XNOR2_X1 U26415 ( .A(n2603), .B(n4694), .ZN(n26225) );
  XNOR2_X1 U26416 ( .A(n26225), .B(n4744), .ZN(n25655) );
  XNOR2_X1 U26417 ( .A(n25655), .B(n15691), .ZN(n34761) );
  XNOR2_X1 U26418 ( .A(n16149), .B(n4720), .ZN(n26057) );
  XNOR2_X1 U26419 ( .A(n26057), .B(n4645), .ZN(n33986) );
  XNOR2_X1 U26420 ( .A(n34761), .B(n33986), .ZN(n15692) );
  XNOR2_X1 U26421 ( .A(n26114), .B(n15692), .ZN(n15693) );
  XNOR2_X1 U26422 ( .A(n15694), .B(n15693), .ZN(n15695) );
  XNOR2_X1 U26423 ( .A(n15695), .B(n16527), .ZN(n15697) );
  XNOR2_X1 U26426 ( .A(n52209), .B(n51336), .ZN(n15696) );
  XNOR2_X1 U26427 ( .A(n15697), .B(n15696), .ZN(n15698) );
  XNOR2_X1 U26428 ( .A(n15699), .B(n15698), .ZN(n15724) );
  XNOR2_X1 U26429 ( .A(n4838), .B(n4897), .ZN(n15700) );
  XNOR2_X1 U26430 ( .A(n25013), .B(n15700), .ZN(n23796) );
  INV_X1 U26431 ( .A(n25616), .ZN(n15701) );
  XNOR2_X1 U26432 ( .A(n23796), .B(n15701), .ZN(n33896) );
  XNOR2_X1 U26433 ( .A(n34709), .B(n4926), .ZN(n43939) );
  XNOR2_X1 U26434 ( .A(n33896), .B(n43939), .ZN(n15702) );
  XNOR2_X1 U26435 ( .A(n4788), .B(n4429), .ZN(n15733) );
  XNOR2_X1 U26436 ( .A(n27316), .B(n15733), .ZN(n34713) );
  XNOR2_X1 U26437 ( .A(n15702), .B(n34713), .ZN(n15703) );
  XNOR2_X1 U26438 ( .A(n51134), .B(n15703), .ZN(n15704) );
  XNOR2_X1 U26439 ( .A(n18704), .B(n15704), .ZN(n15706) );
  XNOR2_X1 U26440 ( .A(n18739), .B(n15738), .ZN(n15877) );
  XNOR2_X1 U26441 ( .A(n16063), .B(n15877), .ZN(n15705) );
  XNOR2_X1 U26442 ( .A(n15705), .B(n15706), .ZN(n15708) );
  XNOR2_X1 U26443 ( .A(n356), .B(n18135), .ZN(n15707) );
  XNOR2_X1 U26444 ( .A(n15708), .B(n16190), .ZN(n15710) );
  INV_X1 U26445 ( .A(n15723), .ZN(n19671) );
  XNOR2_X1 U26446 ( .A(n17947), .B(n15619), .ZN(n15712) );
  XNOR2_X1 U26447 ( .A(n15712), .B(n15711), .ZN(n15718) );
  XNOR2_X1 U26448 ( .A(n16666), .B(n16943), .ZN(n18127) );
  XNOR2_X1 U26449 ( .A(n44952), .B(n43586), .ZN(n27298) );
  XNOR2_X1 U26450 ( .A(n27298), .B(n43105), .ZN(n24767) );
  INV_X1 U26451 ( .A(n24767), .ZN(n15713) );
  XNOR2_X1 U26452 ( .A(n24941), .B(n15713), .ZN(n43076) );
  XNOR2_X1 U26453 ( .A(n43764), .B(n4827), .ZN(n15714) );
  XNOR2_X1 U26454 ( .A(n24127), .B(n15714), .ZN(n35261) );
  XNOR2_X1 U26455 ( .A(n43076), .B(n35261), .ZN(n15715) );
  XNOR2_X1 U26456 ( .A(n17730), .B(n15715), .ZN(n15716) );
  XNOR2_X1 U26457 ( .A(n18127), .B(n15716), .ZN(n15717) );
  XNOR2_X1 U26458 ( .A(n15718), .B(n15717), .ZN(n15720) );
  XNOR2_X1 U26459 ( .A(n16431), .B(n15889), .ZN(n15721) );
  AOI22_X1 U26460 ( .A1(n19672), .A2(n18234), .B1(n20217), .B2(n20211), .ZN(
        n15732) );
  INV_X1 U26461 ( .A(n15724), .ZN(n19680) );
  NAND2_X1 U26463 ( .A1(n51128), .A2(n19685), .ZN(n15727) );
  INV_X1 U26464 ( .A(n19673), .ZN(n16994) );
  NAND2_X1 U26465 ( .A1(n16994), .A2(n15724), .ZN(n19689) );
  NAND2_X1 U26466 ( .A1(n19685), .A2(n51006), .ZN(n18232) );
  NAND2_X1 U26467 ( .A1(n19689), .A2(n18232), .ZN(n15726) );
  NAND3_X1 U26468 ( .A1(n15727), .A2(n15726), .A3(n19681), .ZN(n15731) );
  NAND2_X1 U26469 ( .A1(n20221), .A2(n20215), .ZN(n15730) );
  NAND2_X1 U26470 ( .A1(n20210), .A2(n19685), .ZN(n16995) );
  INV_X1 U26471 ( .A(n51521), .ZN(n19687) );
  OAI211_X1 U26472 ( .C1(n19671), .C2(n19680), .A(n19687), .B(n775), .ZN(
        n15728) );
  NAND3_X1 U26473 ( .A1(n16995), .A2(n51128), .A3(n15728), .ZN(n15729) );
  XNOR2_X1 U26474 ( .A(n18457), .B(n18460), .ZN(n16760) );
  XNOR2_X1 U26475 ( .A(n24797), .B(n43739), .ZN(n17969) );
  XNOR2_X1 U26476 ( .A(n16280), .B(n17969), .ZN(n25615) );
  XNOR2_X1 U26477 ( .A(n25615), .B(n4065), .ZN(n25169) );
  XNOR2_X1 U26478 ( .A(n25616), .B(n4923), .ZN(n45083) );
  XNOR2_X1 U26479 ( .A(n25169), .B(n45083), .ZN(n32342) );
  XNOR2_X1 U26480 ( .A(n34709), .B(n4824), .ZN(n26601) );
  XNOR2_X1 U26481 ( .A(n26601), .B(n4247), .ZN(n46146) );
  XNOR2_X1 U26482 ( .A(n46146), .B(n15733), .ZN(n36861) );
  XNOR2_X1 U26483 ( .A(n32342), .B(n36861), .ZN(n15734) );
  XNOR2_X1 U26484 ( .A(n17831), .B(n15734), .ZN(n15735) );
  XNOR2_X1 U26485 ( .A(n15736), .B(n15735), .ZN(n15737) );
  XNOR2_X1 U26486 ( .A(n16760), .B(n15737), .ZN(n15741) );
  XNOR2_X1 U26487 ( .A(n17821), .B(n18704), .ZN(n15994) );
  XNOR2_X1 U26488 ( .A(n16754), .B(n4529), .ZN(n17292) );
  XNOR2_X1 U26489 ( .A(n17292), .B(n15738), .ZN(n15739) );
  XNOR2_X1 U26490 ( .A(n15994), .B(n15739), .ZN(n15740) );
  XNOR2_X1 U26491 ( .A(n15743), .B(n18480), .ZN(n15971) );
  XNOR2_X1 U26492 ( .A(n15971), .B(n15744), .ZN(n16576) );
  XNOR2_X1 U26493 ( .A(n43764), .B(n4237), .ZN(n34215) );
  INV_X1 U26494 ( .A(n34215), .ZN(n15745) );
  INV_X1 U26495 ( .A(n4526), .ZN(n50899) );
  XNOR2_X1 U26496 ( .A(n43073), .B(n50899), .ZN(n16082) );
  INV_X1 U26497 ( .A(n16082), .ZN(n43589) );
  XNOR2_X1 U26498 ( .A(n15745), .B(n43589), .ZN(n34376) );
  XNOR2_X1 U26499 ( .A(n18126), .B(n34376), .ZN(n15968) );
  XNOR2_X1 U26500 ( .A(n16781), .B(n15968), .ZN(n15747) );
  XNOR2_X1 U26501 ( .A(n41460), .B(n31432), .ZN(n43768) );
  XNOR2_X1 U26502 ( .A(n4687), .B(n4599), .ZN(n26164) );
  XNOR2_X1 U26503 ( .A(n4275), .B(n4026), .ZN(n28090) );
  XNOR2_X1 U26504 ( .A(n26164), .B(n28090), .ZN(n33746) );
  XNOR2_X1 U26505 ( .A(n44952), .B(n4845), .ZN(n33745) );
  XNOR2_X1 U26506 ( .A(n33746), .B(n33745), .ZN(n15748) );
  XNOR2_X1 U26507 ( .A(n43768), .B(n15748), .ZN(n15749) );
  XNOR2_X1 U26508 ( .A(n16294), .B(n15749), .ZN(n15750) );
  INV_X1 U26509 ( .A(n17177), .ZN(n18476) );
  XNOR2_X1 U26510 ( .A(n18476), .B(n15750), .ZN(n15751) );
  XNOR2_X1 U26511 ( .A(n18696), .B(n17947), .ZN(n17727) );
  XNOR2_X1 U26512 ( .A(n15751), .B(n17727), .ZN(n15752) );
  AND2_X1 U26513 ( .A1(n20266), .A2(n20659), .ZN(n20652) );
  XNOR2_X1 U26514 ( .A(n17936), .B(n17117), .ZN(n15753) );
  XNOR2_X1 U26515 ( .A(n15753), .B(n18795), .ZN(n18419) );
  XNOR2_X1 U26516 ( .A(n15754), .B(n18419), .ZN(n15783) );
  XNOR2_X1 U26517 ( .A(n35796), .B(n4624), .ZN(n24725) );
  XNOR2_X1 U26518 ( .A(n17243), .B(n24725), .ZN(n33959) );
  XNOR2_X1 U26519 ( .A(n18636), .B(n4723), .ZN(n34742) );
  XNOR2_X1 U26520 ( .A(n34742), .B(n47401), .ZN(n15755) );
  XNOR2_X1 U26521 ( .A(n33959), .B(n15755), .ZN(n15757) );
  XNOR2_X1 U26522 ( .A(n23370), .B(n16241), .ZN(n15756) );
  INV_X1 U26523 ( .A(n43702), .ZN(n44015) );
  XNOR2_X1 U26524 ( .A(n15756), .B(n44015), .ZN(n19769) );
  XNOR2_X1 U26525 ( .A(n19769), .B(n25078), .ZN(n34744) );
  XNOR2_X1 U26526 ( .A(n15757), .B(n34744), .ZN(n15762) );
  INV_X1 U26527 ( .A(n15758), .ZN(n15759) );
  OAI21_X1 U26528 ( .B1(n15760), .B2(n15759), .A(n15762), .ZN(n15761) );
  OAI21_X1 U26529 ( .B1(n15763), .B2(n15762), .A(n15761), .ZN(n15765) );
  XNOR2_X1 U26530 ( .A(n17804), .B(n17643), .ZN(n15764) );
  XNOR2_X1 U26531 ( .A(n15765), .B(n15764), .ZN(n15781) );
  MUX2_X1 U26532 ( .A(n15767), .B(n15770), .S(n15766), .Z(n15779) );
  INV_X1 U26533 ( .A(n15768), .ZN(n15772) );
  INV_X1 U26534 ( .A(n15769), .ZN(n15771) );
  AOI21_X1 U26535 ( .B1(n15772), .B2(n15771), .A(n15770), .ZN(n15775) );
  INV_X1 U26536 ( .A(n15773), .ZN(n15774) );
  NOR2_X1 U26537 ( .A1(n15775), .A2(n15774), .ZN(n15776) );
  OAI211_X1 U26538 ( .C1(n15779), .C2(n15778), .A(n15777), .B(n15776), .ZN(
        n18208) );
  XNOR2_X1 U26539 ( .A(n19250), .B(n18208), .ZN(n15780) );
  XNOR2_X1 U26540 ( .A(n15780), .B(n15781), .ZN(n15782) );
  XNOR2_X1 U26541 ( .A(n15782), .B(n15783), .ZN(n15788) );
  XNOR2_X1 U26542 ( .A(n19248), .B(n18427), .ZN(n15784) );
  XNOR2_X1 U26543 ( .A(n15784), .B(n17125), .ZN(n16057) );
  XNOR2_X1 U26544 ( .A(n16532), .B(n17364), .ZN(n16704) );
  XNOR2_X1 U26545 ( .A(n17803), .B(n17365), .ZN(n15785) );
  XNOR2_X1 U26546 ( .A(n16704), .B(n15785), .ZN(n15786) );
  XNOR2_X1 U26547 ( .A(n15786), .B(n16057), .ZN(n15787) );
  XNOR2_X1 U26548 ( .A(n23943), .B(n25898), .ZN(n28391) );
  XNOR2_X1 U26549 ( .A(n28391), .B(n26525), .ZN(n15789) );
  XNOR2_X1 U26550 ( .A(n33374), .B(n4627), .ZN(n36718) );
  XNOR2_X1 U26551 ( .A(n36718), .B(n4884), .ZN(n15942) );
  XNOR2_X1 U26552 ( .A(n15789), .B(n15942), .ZN(n36802) );
  XNOR2_X1 U26553 ( .A(n34027), .B(n25901), .ZN(n32268) );
  XNOR2_X1 U26554 ( .A(n48843), .B(n4720), .ZN(n15790) );
  XNOR2_X1 U26555 ( .A(n32268), .B(n15790), .ZN(n15791) );
  XNOR2_X1 U26556 ( .A(n32856), .B(n4874), .ZN(n44887) );
  XNOR2_X1 U26557 ( .A(n15791), .B(n44887), .ZN(n15792) );
  XNOR2_X1 U26558 ( .A(n36802), .B(n15792), .ZN(n15793) );
  XNOR2_X1 U26559 ( .A(n18437), .B(n15793), .ZN(n15794) );
  XNOR2_X1 U26560 ( .A(n15794), .B(n51757), .ZN(n15795) );
  XNOR2_X1 U26562 ( .A(n15795), .B(n18446), .ZN(n15799) );
  XNOR2_X1 U26563 ( .A(n17787), .B(n15796), .ZN(n15797) );
  XNOR2_X1 U26564 ( .A(n2218), .B(n15797), .ZN(n15798) );
  INV_X1 U26566 ( .A(n18193), .ZN(n16024) );
  XNOR2_X1 U26567 ( .A(n16228), .B(n17786), .ZN(n15801) );
  XNOR2_X1 U26568 ( .A(n18194), .B(n15801), .ZN(n15802) );
  XNOR2_X1 U26569 ( .A(n16527), .B(n15802), .ZN(n15906) );
  XNOR2_X1 U26570 ( .A(n16234), .B(n15906), .ZN(n15803) );
  INV_X1 U26572 ( .A(n20650), .ZN(n16892) );
  XNOR2_X1 U26573 ( .A(n15805), .B(n2181), .ZN(n18785) );
  XNOR2_X1 U26574 ( .A(n17902), .B(n4755), .ZN(n15806) );
  XNOR2_X1 U26575 ( .A(n16980), .B(n15806), .ZN(n15807) );
  XNOR2_X1 U26576 ( .A(n15808), .B(n15807), .ZN(n18652) );
  XNOR2_X1 U26577 ( .A(n18785), .B(n18652), .ZN(n15817) );
  XNOR2_X1 U26578 ( .A(n16105), .B(n16416), .ZN(n15809) );
  XNOR2_X1 U26579 ( .A(n15809), .B(n17322), .ZN(n19216) );
  XNOR2_X1 U26580 ( .A(n26370), .B(n26296), .ZN(n25041) );
  XNOR2_X1 U26581 ( .A(n25041), .B(n28270), .ZN(n33690) );
  XNOR2_X1 U26582 ( .A(n28412), .B(n4706), .ZN(n34616) );
  XNOR2_X1 U26583 ( .A(n33690), .B(n34616), .ZN(n15810) );
  XNOR2_X1 U26584 ( .A(n17212), .B(n15810), .ZN(n15811) );
  XNOR2_X1 U26585 ( .A(n15812), .B(n15811), .ZN(n15813) );
  XNOR2_X1 U26586 ( .A(n19216), .B(n15813), .ZN(n15815) );
  XNOR2_X1 U26587 ( .A(n17208), .B(n1326), .ZN(n17908) );
  XNOR2_X1 U26588 ( .A(n17213), .B(n4880), .ZN(n18180) );
  XNOR2_X1 U26589 ( .A(n17908), .B(n18180), .ZN(n15814) );
  XNOR2_X1 U26590 ( .A(n15815), .B(n15814), .ZN(n15816) );
  XNOR2_X1 U26591 ( .A(n4554), .B(n4885), .ZN(n15818) );
  XNOR2_X1 U26592 ( .A(n41155), .B(n15818), .ZN(n25939) );
  XNOR2_X1 U26593 ( .A(n25939), .B(n4564), .ZN(n35290) );
  XNOR2_X1 U26594 ( .A(n4423), .B(Key[57]), .ZN(n24919) );
  XNOR2_X1 U26595 ( .A(n35290), .B(n24919), .ZN(n35653) );
  XNOR2_X1 U26596 ( .A(n20856), .B(n34411), .ZN(n15819) );
  XNOR2_X1 U26597 ( .A(n35653), .B(n15819), .ZN(n15820) );
  XNOR2_X1 U26598 ( .A(n43654), .B(n1224), .ZN(n31719) );
  XNOR2_X1 U26599 ( .A(n15820), .B(n31719), .ZN(n15821) );
  XNOR2_X1 U26600 ( .A(n15822), .B(n18407), .ZN(n15823) );
  XNOR2_X1 U26601 ( .A(n15824), .B(n15823), .ZN(n15826) );
  XNOR2_X1 U26602 ( .A(n18163), .B(n52194), .ZN(n15825) );
  XNOR2_X1 U26603 ( .A(n15826), .B(n15825), .ZN(n15831) );
  XNOR2_X1 U26604 ( .A(n17234), .B(n18399), .ZN(n15828) );
  XNOR2_X1 U26605 ( .A(n18756), .B(n18157), .ZN(n15827) );
  XNOR2_X1 U26606 ( .A(n15828), .B(n15827), .ZN(n15829) );
  XNOR2_X1 U26607 ( .A(n543), .B(n15829), .ZN(n15830) );
  XNOR2_X1 U26608 ( .A(n17754), .B(n51437), .ZN(n19211) );
  XNOR2_X1 U26609 ( .A(n19211), .B(n15830), .ZN(n15984) );
  OAI22_X1 U26610 ( .A1(n16892), .A2(n18846), .B1(n18847), .B2(n20656), .ZN(
        n15834) );
  NOR2_X1 U26611 ( .A1(n21664), .A2(n20266), .ZN(n15832) );
  NAND2_X1 U26613 ( .A1(n21660), .A2(n21656), .ZN(n16886) );
  OR2_X1 U26614 ( .A1(n20649), .A2(n20266), .ZN(n21655) );
  AND2_X1 U26615 ( .A1(n20657), .A2(n21661), .ZN(n21649) );
  NOR2_X1 U26616 ( .A1(n20277), .A2(n20266), .ZN(n15836) );
  NAND4_X1 U26617 ( .A1(n20650), .A2(n20649), .A3(n21660), .A4(n21664), .ZN(
        n20267) );
  INV_X1 U26618 ( .A(n20267), .ZN(n15835) );
  NAND3_X1 U26619 ( .A1(n24150), .A2(n24158), .A3(n23821), .ZN(n16004) );
  XNOR2_X1 U26620 ( .A(n17232), .B(n33050), .ZN(n15840) );
  XNOR2_X1 U26621 ( .A(n15840), .B(n18505), .ZN(n15841) );
  XNOR2_X1 U26622 ( .A(n15841), .B(n18162), .ZN(n16264) );
  XNOR2_X1 U26623 ( .A(n28058), .B(n44044), .ZN(n39719) );
  INV_X1 U26624 ( .A(n39719), .ZN(n25343) );
  XNOR2_X1 U26625 ( .A(n25343), .B(n4565), .ZN(n33053) );
  XNOR2_X1 U26626 ( .A(n4451), .B(n3367), .ZN(n22816) );
  XNOR2_X1 U26627 ( .A(n26358), .B(n22816), .ZN(n37299) );
  XNOR2_X1 U26628 ( .A(n37299), .B(n25683), .ZN(n15842) );
  XNOR2_X1 U26629 ( .A(n33053), .B(n15842), .ZN(n15843) );
  XNOR2_X1 U26630 ( .A(n19199), .B(n15843), .ZN(n15844) );
  XNOR2_X1 U26631 ( .A(n15848), .B(n15847), .ZN(n15849) );
  XNOR2_X1 U26632 ( .A(n16264), .B(n15849), .ZN(n15850) );
  INV_X1 U26633 ( .A(n15871), .ZN(n20683) );
  XNOR2_X1 U26634 ( .A(n51032), .B(n511), .ZN(n15853) );
  INV_X1 U26635 ( .A(n17914), .ZN(n15852) );
  XNOR2_X1 U26636 ( .A(n15853), .B(n15852), .ZN(n15854) );
  XNOR2_X1 U26637 ( .A(n15854), .B(n16259), .ZN(n18185) );
  XNOR2_X1 U26638 ( .A(n18169), .B(n49414), .ZN(n16422) );
  XNOR2_X1 U26639 ( .A(n16422), .B(n17771), .ZN(n16970) );
  INV_X1 U26640 ( .A(n2606), .ZN(n15855) );
  XNOR2_X1 U26641 ( .A(n15855), .B(n25040), .ZN(n18390) );
  INV_X1 U26642 ( .A(n18390), .ZN(n28271) );
  XNOR2_X1 U26643 ( .A(n26296), .B(n28271), .ZN(n15856) );
  XNOR2_X1 U26644 ( .A(n29662), .B(n4490), .ZN(n24582) );
  XNOR2_X1 U26645 ( .A(n24582), .B(n4325), .ZN(n24695) );
  XNOR2_X1 U26646 ( .A(n15856), .B(n24695), .ZN(n35480) );
  XNOR2_X1 U26647 ( .A(n25042), .B(n27364), .ZN(n43053) );
  XNOR2_X1 U26648 ( .A(n43053), .B(n33653), .ZN(n35393) );
  XNOR2_X1 U26649 ( .A(n35480), .B(n35393), .ZN(n15857) );
  XNOR2_X1 U26650 ( .A(n2121), .B(n15857), .ZN(n15858) );
  XNOR2_X1 U26651 ( .A(n17902), .B(n15858), .ZN(n15860) );
  XNOR2_X1 U26652 ( .A(n15860), .B(n15859), .ZN(n15861) );
  XNOR2_X1 U26653 ( .A(n16970), .B(n15861), .ZN(n15863) );
  INV_X1 U26654 ( .A(n18664), .ZN(n15862) );
  XNOR2_X1 U26655 ( .A(n15863), .B(n15862), .ZN(n15864) );
  XNOR2_X1 U26656 ( .A(n15864), .B(n18185), .ZN(n15872) );
  XNOR2_X1 U26659 ( .A(n19769), .B(n24057), .ZN(n18422) );
  INV_X1 U26660 ( .A(n18422), .ZN(n27173) );
  XNOR2_X1 U26661 ( .A(n27173), .B(n25426), .ZN(n22614) );
  XNOR2_X1 U26662 ( .A(n4353), .B(n4517), .ZN(n25640) );
  XNOR2_X1 U26663 ( .A(n22614), .B(n25640), .ZN(n33391) );
  XNOR2_X1 U26664 ( .A(n25147), .B(n4746), .ZN(n16900) );
  XNOR2_X1 U26665 ( .A(n4939), .B(n3276), .ZN(n28425) );
  XNOR2_X1 U26666 ( .A(n28425), .B(n49323), .ZN(n15865) );
  XNOR2_X1 U26667 ( .A(n16900), .B(n15865), .ZN(n34283) );
  XNOR2_X1 U26668 ( .A(n33391), .B(n34283), .ZN(n15866) );
  XNOR2_X1 U26669 ( .A(n16707), .B(n15869), .ZN(n15870) );
  XNOR2_X1 U26670 ( .A(n18797), .B(n19250), .ZN(n18418) );
  OAI21_X1 U26671 ( .B1(n18101), .B2(n20682), .A(n20685), .ZN(n15902) );
  INV_X1 U26672 ( .A(n17297), .ZN(n15873) );
  XNOR2_X1 U26673 ( .A(n8699), .B(n15873), .ZN(n15874) );
  XNOR2_X1 U26674 ( .A(n15874), .B(n17831), .ZN(n15875) );
  XNOR2_X1 U26675 ( .A(n576), .B(n15875), .ZN(n17175) );
  XNOR2_X1 U26676 ( .A(n18750), .B(n18457), .ZN(n16075) );
  INV_X1 U26677 ( .A(n16075), .ZN(n18705) );
  XNOR2_X1 U26678 ( .A(n44493), .B(n23495), .ZN(n15878) );
  XNOR2_X1 U26679 ( .A(n15878), .B(n43739), .ZN(n18131) );
  XNOR2_X1 U26680 ( .A(n18131), .B(n24797), .ZN(n24749) );
  XNOR2_X1 U26681 ( .A(n26178), .B(n4691), .ZN(n15879) );
  XNOR2_X1 U26682 ( .A(n26025), .B(n15879), .ZN(n15880) );
  XNOR2_X1 U26683 ( .A(n24749), .B(n15880), .ZN(n33180) );
  XNOR2_X1 U26684 ( .A(n42686), .B(n4655), .ZN(n34816) );
  XNOR2_X1 U26685 ( .A(n34816), .B(n4712), .ZN(n15881) );
  XNOR2_X1 U26686 ( .A(n33180), .B(n15881), .ZN(n15882) );
  XNOR2_X1 U26687 ( .A(n17690), .B(n15882), .ZN(n15884) );
  XNOR2_X1 U26688 ( .A(n15883), .B(n15884), .ZN(n15885) );
  XNOR2_X1 U26689 ( .A(n15885), .B(n635), .ZN(n15886) );
  XNOR2_X1 U26690 ( .A(n18705), .B(n15886), .ZN(n15887) );
  INV_X1 U26691 ( .A(n17738), .ZN(n15890) );
  XNOR2_X1 U26692 ( .A(n16294), .B(n18119), .ZN(n15891) );
  XNOR2_X1 U26693 ( .A(n18476), .B(n15891), .ZN(n15898) );
  XNOR2_X1 U26694 ( .A(n43073), .B(n43764), .ZN(n15892) );
  XNOR2_X1 U26695 ( .A(n15892), .B(n42322), .ZN(n28089) );
  XNOR2_X1 U26696 ( .A(n42297), .B(n28085), .ZN(n43265) );
  XNOR2_X1 U26697 ( .A(n28089), .B(n43265), .ZN(n18124) );
  XNOR2_X1 U26698 ( .A(n28084), .B(n4864), .ZN(n15893) );
  XNOR2_X1 U26699 ( .A(n18124), .B(n15893), .ZN(n35352) );
  XNOR2_X1 U26700 ( .A(n33474), .B(n43105), .ZN(n35518) );
  XNOR2_X1 U26701 ( .A(n35518), .B(n1341), .ZN(n15894) );
  XNOR2_X1 U26702 ( .A(n35352), .B(n15894), .ZN(n15895) );
  XNOR2_X1 U26703 ( .A(n15896), .B(n15895), .ZN(n15897) );
  XNOR2_X1 U26704 ( .A(n15899), .B(n16431), .ZN(n15901) );
  INV_X1 U26705 ( .A(n18696), .ZN(n15900) );
  XNOR2_X1 U26706 ( .A(n16568), .B(n15900), .ZN(n18489) );
  INV_X1 U26707 ( .A(n18431), .ZN(n15903) );
  XNOR2_X1 U26708 ( .A(n16919), .B(n4653), .ZN(n15904) );
  XNOR2_X1 U26709 ( .A(n16525), .B(n15904), .ZN(n15905) );
  XNOR2_X1 U26710 ( .A(n15905), .B(n2217), .ZN(n16717) );
  XNOR2_X1 U26711 ( .A(n16717), .B(n15906), .ZN(n15919) );
  XNOR2_X1 U26712 ( .A(n23943), .B(n2603), .ZN(n15907) );
  XNOR2_X1 U26713 ( .A(n15907), .B(n25898), .ZN(n24550) );
  XNOR2_X1 U26714 ( .A(n24550), .B(n17661), .ZN(n25537) );
  XNOR2_X1 U26715 ( .A(n25537), .B(n4744), .ZN(n34865) );
  XNOR2_X1 U26716 ( .A(n25901), .B(n7744), .ZN(n40847) );
  XNOR2_X1 U26717 ( .A(n40847), .B(n15908), .ZN(n33215) );
  XNOR2_X1 U26718 ( .A(n48843), .B(n33221), .ZN(n15909) );
  XNOR2_X1 U26719 ( .A(n33215), .B(n15909), .ZN(n15910) );
  XNOR2_X1 U26720 ( .A(n34865), .B(n15910), .ZN(n15911) );
  XNOR2_X1 U26721 ( .A(n52228), .B(n15911), .ZN(n15912) );
  XNOR2_X1 U26722 ( .A(n15912), .B(n51459), .ZN(n15914) );
  XNOR2_X1 U26723 ( .A(n18447), .B(n15913), .ZN(n16156) );
  XNOR2_X1 U26724 ( .A(n15914), .B(n16156), .ZN(n15917) );
  XNOR2_X1 U26725 ( .A(n51336), .B(n51482), .ZN(n15916) );
  XNOR2_X1 U26726 ( .A(n15917), .B(n15916), .ZN(n15918) );
  OR2_X1 U26727 ( .A1(n15920), .A2(n20227), .ZN(n15927) );
  NOR2_X1 U26728 ( .A1(n18102), .A2(n20683), .ZN(n15922) );
  AND3_X1 U26729 ( .A1(n1597), .A2(n20681), .A3(n20677), .ZN(n15921) );
  AOI22_X1 U26730 ( .A1(n15922), .A2(n20678), .B1(n18875), .B2(n15921), .ZN(
        n15926) );
  NAND2_X1 U26732 ( .A1(n20688), .A2(n20683), .ZN(n18867) );
  INV_X1 U26733 ( .A(n20674), .ZN(n15924) );
  OAI21_X1 U26734 ( .B1(n15924), .B2(n15923), .A(n1597), .ZN(n15925) );
  NAND2_X1 U26736 ( .A1(n18863), .A2(n20677), .ZN(n20668) );
  NOR2_X1 U26737 ( .A1(n20239), .A2(n20668), .ZN(n15929) );
  INV_X1 U26738 ( .A(n20686), .ZN(n16873) );
  MUX2_X1 U26739 ( .A(n20230), .B(n15929), .S(n16873), .Z(n15930) );
  XNOR2_X1 U26740 ( .A(n15933), .B(n15932), .ZN(n17819) );
  XNOR2_X1 U26741 ( .A(n51402), .B(n17819), .ZN(n18589) );
  XNOR2_X1 U26742 ( .A(n25744), .B(n18423), .ZN(n25325) );
  XNOR2_X1 U26743 ( .A(n35532), .B(n25325), .ZN(n24818) );
  XNOR2_X1 U26744 ( .A(n27174), .B(n49323), .ZN(n16698) );
  XNOR2_X1 U26745 ( .A(n24818), .B(n16698), .ZN(n33230) );
  XNOR2_X1 U26746 ( .A(n16241), .B(n4723), .ZN(n28309) );
  XNOR2_X1 U26747 ( .A(n4517), .B(n4208), .ZN(n24056) );
  XNOR2_X1 U26748 ( .A(n28309), .B(n24056), .ZN(n34851) );
  XNOR2_X1 U26749 ( .A(n33230), .B(n34851), .ZN(n15934) );
  XNOR2_X1 U26750 ( .A(n17643), .B(n15934), .ZN(n15935) );
  XNOR2_X1 U26751 ( .A(n18644), .B(n15935), .ZN(n15937) );
  XNOR2_X1 U26752 ( .A(n485), .B(n18208), .ZN(n15936) );
  XNOR2_X1 U26753 ( .A(n15937), .B(n15936), .ZN(n15938) );
  XNOR2_X1 U26755 ( .A(n18589), .B(n15941), .ZN(n21632) );
  XNOR2_X1 U26756 ( .A(n15942), .B(n4653), .ZN(n43563) );
  XNOR2_X1 U26757 ( .A(n43563), .B(n23943), .ZN(n15944) );
  XNOR2_X1 U26758 ( .A(n4537), .B(n4781), .ZN(n24553) );
  XNOR2_X1 U26759 ( .A(n33221), .B(n4720), .ZN(n28284) );
  XNOR2_X1 U26760 ( .A(n24553), .B(n28284), .ZN(n18555) );
  XNOR2_X1 U26761 ( .A(n34027), .B(n4890), .ZN(n24315) );
  XNOR2_X1 U26762 ( .A(n18555), .B(n24315), .ZN(n23399) );
  XNOR2_X1 U26763 ( .A(n35815), .B(n1313), .ZN(n24554) );
  XNOR2_X1 U26764 ( .A(n24554), .B(n27353), .ZN(n15943) );
  XNOR2_X1 U26765 ( .A(n23399), .B(n15943), .ZN(n32037) );
  XNOR2_X1 U26766 ( .A(n15944), .B(n32037), .ZN(n15945) );
  XNOR2_X1 U26767 ( .A(n18437), .B(n18193), .ZN(n18813) );
  INV_X1 U26768 ( .A(n18813), .ZN(n15946) );
  XNOR2_X1 U26769 ( .A(n17787), .B(n51642), .ZN(n15947) );
  XNOR2_X1 U26770 ( .A(n15947), .B(n52209), .ZN(n19239) );
  XNOR2_X1 U26771 ( .A(n17264), .B(n18615), .ZN(n15949) );
  XNOR2_X1 U26772 ( .A(n15949), .B(n18617), .ZN(n18436) );
  XNOR2_X1 U26773 ( .A(n15950), .B(n18443), .ZN(n15951) );
  XNOR2_X1 U26774 ( .A(n15951), .B(n51482), .ZN(n18553) );
  INV_X1 U26775 ( .A(n20244), .ZN(n20256) );
  INV_X1 U26776 ( .A(n21619), .ZN(n15986) );
  XNOR2_X1 U26777 ( .A(Key[180]), .B(n4752), .ZN(n41223) );
  XNOR2_X1 U26778 ( .A(n41223), .B(n26541), .ZN(n27485) );
  XNOR2_X1 U26779 ( .A(n27485), .B(n46062), .ZN(n15952) );
  XNOR2_X1 U26780 ( .A(n15952), .B(n24585), .ZN(n34365) );
  XNOR2_X1 U26781 ( .A(n4415), .B(n1336), .ZN(n18778) );
  XNOR2_X1 U26782 ( .A(n4325), .B(n4639), .ZN(n16164) );
  XNOR2_X1 U26783 ( .A(n18778), .B(n16164), .ZN(n25115) );
  XNOR2_X1 U26784 ( .A(n25115), .B(n41567), .ZN(n33655) );
  XNOR2_X1 U26785 ( .A(n33655), .B(n4490), .ZN(n15953) );
  XNOR2_X1 U26786 ( .A(n34365), .B(n15953), .ZN(n15954) );
  XNOR2_X1 U26787 ( .A(n17902), .B(n15954), .ZN(n15955) );
  XNOR2_X1 U26788 ( .A(n17208), .B(n15955), .ZN(n15959) );
  INV_X1 U26789 ( .A(n15956), .ZN(n18658) );
  XNOR2_X1 U26790 ( .A(n18658), .B(n15957), .ZN(n15958) );
  XNOR2_X1 U26791 ( .A(n15959), .B(n15958), .ZN(n15960) );
  XNOR2_X1 U26792 ( .A(n18539), .B(n16973), .ZN(n17713) );
  XNOR2_X1 U26793 ( .A(n17713), .B(n15960), .ZN(n15961) );
  XNOR2_X1 U26794 ( .A(n18785), .B(n15961), .ZN(n15963) );
  XNOR2_X1 U26795 ( .A(n24767), .B(n15964), .ZN(n33588) );
  XNOR2_X1 U26796 ( .A(n25866), .B(n1341), .ZN(n15965) );
  XNOR2_X1 U26797 ( .A(n33588), .B(n15965), .ZN(n15966) );
  XNOR2_X1 U26798 ( .A(n18483), .B(n15966), .ZN(n15967) );
  XNOR2_X1 U26799 ( .A(n15967), .B(n17731), .ZN(n15969) );
  XNOR2_X1 U26800 ( .A(n15969), .B(n15968), .ZN(n15970) );
  XNOR2_X1 U26801 ( .A(n15970), .B(n16093), .ZN(n15975) );
  INV_X1 U26802 ( .A(n15971), .ZN(n15973) );
  XNOR2_X1 U26803 ( .A(n15973), .B(n15972), .ZN(n15974) );
  XNOR2_X1 U26804 ( .A(n15975), .B(n15974), .ZN(n15977) );
  INV_X1 U26805 ( .A(n17839), .ZN(n18575) );
  XNOR2_X1 U26806 ( .A(n16438), .B(n18575), .ZN(n15976) );
  OR2_X1 U26808 ( .A1(n19981), .A2(n21613), .ZN(n21631) );
  XNOR2_X1 U26809 ( .A(n17764), .B(n4666), .ZN(n15978) );
  XNOR2_X1 U26810 ( .A(n16952), .B(n15978), .ZN(n18678) );
  XNOR2_X1 U26811 ( .A(n34414), .B(n4868), .ZN(n36823) );
  XNOR2_X1 U26812 ( .A(n36823), .B(n41155), .ZN(n18401) );
  XNOR2_X1 U26813 ( .A(n4316), .B(n4554), .ZN(n28376) );
  XNOR2_X1 U26814 ( .A(n18401), .B(n28376), .ZN(n35380) );
  XNOR2_X1 U26815 ( .A(n44044), .B(n4312), .ZN(n15979) );
  XNOR2_X1 U26816 ( .A(n15979), .B(n43863), .ZN(n35465) );
  XNOR2_X1 U26817 ( .A(n35380), .B(n35465), .ZN(n15980) );
  XNOR2_X1 U26818 ( .A(n17138), .B(n15980), .ZN(n15981) );
  XNOR2_X1 U26819 ( .A(n18678), .B(n15981), .ZN(n15982) );
  XNOR2_X1 U26820 ( .A(n15983), .B(n15982), .ZN(n15985) );
  INV_X1 U26822 ( .A(n21613), .ZN(n20696) );
  NAND3_X1 U26823 ( .A1(n21614), .A2(n20244), .A3(n8367), .ZN(n18729) );
  XNOR2_X1 U26824 ( .A(n27316), .B(n45463), .ZN(n28234) );
  XNOR2_X1 U26825 ( .A(n42686), .B(n4818), .ZN(n35838) );
  XNOR2_X1 U26826 ( .A(n35838), .B(n26601), .ZN(n37042) );
  XNOR2_X1 U26827 ( .A(n28234), .B(n37042), .ZN(n36683) );
  XNOR2_X1 U26828 ( .A(n44493), .B(n15987), .ZN(n33123) );
  XNOR2_X1 U26829 ( .A(n24797), .B(n4065), .ZN(n16556) );
  XNOR2_X1 U26830 ( .A(n33123), .B(n16556), .ZN(n31594) );
  XNOR2_X1 U26831 ( .A(n36683), .B(n31594), .ZN(n15988) );
  XNOR2_X1 U26832 ( .A(n17297), .B(n15988), .ZN(n15989) );
  XNOR2_X1 U26833 ( .A(n52142), .B(n15989), .ZN(n15991) );
  XNOR2_X1 U26834 ( .A(n15991), .B(n15990), .ZN(n15992) );
  XNOR2_X1 U26835 ( .A(n15992), .B(n18605), .ZN(n15993) );
  XNOR2_X1 U26836 ( .A(n15993), .B(n17976), .ZN(n15996) );
  XNOR2_X1 U26837 ( .A(n15995), .B(n15994), .ZN(n19272) );
  NAND2_X1 U26838 ( .A1(n21632), .A2(n20256), .ZN(n20258) );
  INV_X1 U26839 ( .A(n20258), .ZN(n15998) );
  NAND2_X1 U26840 ( .A1(n21614), .A2(n20698), .ZN(n21615) );
  NAND3_X1 U26841 ( .A1(n18731), .A2(n20240), .A3(n21619), .ZN(n20249) );
  OR2_X1 U26842 ( .A1(n16000), .A2(n21632), .ZN(n20694) );
  INV_X1 U26843 ( .A(n20694), .ZN(n16001) );
  AND2_X1 U26844 ( .A1(n21632), .A2(n20244), .ZN(n20700) );
  NAND2_X1 U26845 ( .A1(n21619), .A2(n21630), .ZN(n21624) );
  INV_X1 U26846 ( .A(n18731), .ZN(n20241) );
  NAND3_X1 U26847 ( .A1(n21624), .A2(n21617), .A3(n20241), .ZN(n16002) );
  NAND2_X1 U26848 ( .A1(n23833), .A2(n23825), .ZN(n16003) );
  NAND4_X1 U26849 ( .A1(n16004), .A2(n24159), .A3(n23832), .A4(n16003), .ZN(
        n16006) );
  NAND2_X1 U26850 ( .A1(n23826), .A2(n23833), .ZN(n16005) );
  AND2_X1 U26851 ( .A1(n16006), .A2(n16005), .ZN(n16135) );
  XNOR2_X1 U26852 ( .A(n52227), .B(n17787), .ZN(n16007) );
  XNOR2_X1 U26853 ( .A(n16007), .B(n51757), .ZN(n16015) );
  XNOR2_X1 U26854 ( .A(n17258), .B(n4636), .ZN(n16233) );
  XNOR2_X1 U26855 ( .A(n18555), .B(n25901), .ZN(n25434) );
  INV_X1 U26856 ( .A(n27186), .ZN(n28115) );
  XNOR2_X1 U26857 ( .A(n25434), .B(n28115), .ZN(n41314) );
  XNOR2_X1 U26858 ( .A(n33374), .B(n4744), .ZN(n36964) );
  XNOR2_X1 U26859 ( .A(n2603), .B(n48843), .ZN(n16008) );
  XNOR2_X1 U26860 ( .A(n36964), .B(n16008), .ZN(n16009) );
  XNOR2_X1 U26861 ( .A(n41314), .B(n16009), .ZN(n16010) );
  XNOR2_X1 U26862 ( .A(n16011), .B(n16010), .ZN(n16012) );
  XNOR2_X1 U26865 ( .A(n16015), .B(n16014), .ZN(n16022) );
  XNOR2_X1 U26866 ( .A(n16017), .B(n16016), .ZN(n16019) );
  XNOR2_X1 U26867 ( .A(n16711), .B(n18443), .ZN(n16018) );
  XNOR2_X1 U26868 ( .A(n16019), .B(n16018), .ZN(n16020) );
  XNOR2_X1 U26869 ( .A(n16020), .B(n17798), .ZN(n16021) );
  XNOR2_X1 U26870 ( .A(n16022), .B(n16021), .ZN(n16027) );
  XNOR2_X1 U26871 ( .A(n4653), .B(n4874), .ZN(n45401) );
  XNOR2_X1 U26872 ( .A(n16023), .B(n45401), .ZN(n16025) );
  XNOR2_X1 U26873 ( .A(n16025), .B(n16024), .ZN(n16026) );
  XNOR2_X1 U26874 ( .A(n17356), .B(n16026), .ZN(n16361) );
  XNOR2_X1 U26875 ( .A(n16361), .B(n16027), .ZN(n18897) );
  XNOR2_X1 U26876 ( .A(n17368), .B(n16028), .ZN(n18581) );
  XNOR2_X1 U26877 ( .A(n52229), .B(n16029), .ZN(n16030) );
  XNOR2_X1 U26878 ( .A(n16030), .B(n18581), .ZN(n16059) );
  XNOR2_X1 U26879 ( .A(n28303), .B(n24725), .ZN(n24639) );
  XNOR2_X1 U26880 ( .A(n25325), .B(n4076), .ZN(n16031) );
  XNOR2_X1 U26881 ( .A(n24639), .B(n16031), .ZN(n34047) );
  XNOR2_X1 U26882 ( .A(n4932), .B(n4517), .ZN(n16032) );
  XNOR2_X1 U26883 ( .A(n16241), .B(n16032), .ZN(n33854) );
  XNOR2_X1 U26884 ( .A(n34047), .B(n33854), .ZN(n16033) );
  XNOR2_X1 U26885 ( .A(n17117), .B(n16033), .ZN(n16055) );
  AND2_X1 U26886 ( .A1(n16035), .A2(n16034), .ZN(n16054) );
  MUX2_X1 U26887 ( .A(n16038), .B(n51019), .S(n16036), .Z(n16042) );
  NOR2_X1 U26888 ( .A1(n16040), .A2(n16039), .ZN(n16041) );
  NAND2_X1 U26889 ( .A1(n16042), .A2(n16041), .ZN(n16053) );
  OAI21_X1 U26890 ( .B1(n16045), .B2(n16044), .A(n16043), .ZN(n16047) );
  XNOR2_X1 U26893 ( .A(n16055), .B(n18790), .ZN(n16056) );
  XNOR2_X1 U26894 ( .A(n16057), .B(n16056), .ZN(n16058) );
  XNOR2_X1 U26895 ( .A(n16059), .B(n16058), .ZN(n16061) );
  XNOR2_X1 U26896 ( .A(n17127), .B(n2225), .ZN(n16060) );
  XNOR2_X1 U26897 ( .A(n17240), .B(n16060), .ZN(n16381) );
  XNOR2_X1 U26898 ( .A(n17821), .B(n18739), .ZN(n16062) );
  XNOR2_X1 U26899 ( .A(n16063), .B(n16062), .ZN(n16073) );
  XNOR2_X1 U26900 ( .A(n4691), .B(n4897), .ZN(n33121) );
  XNOR2_X1 U26901 ( .A(n4908), .B(n2203), .ZN(n16065) );
  XNOR2_X1 U26902 ( .A(n33121), .B(n16065), .ZN(n16066) );
  XNOR2_X1 U26903 ( .A(n33123), .B(n16066), .ZN(n16067) );
  XNOR2_X1 U26904 ( .A(n42686), .B(n4247), .ZN(n36943) );
  XNOR2_X1 U26905 ( .A(n16067), .B(n36943), .ZN(n16068) );
  XNOR2_X1 U26906 ( .A(n16068), .B(n33899), .ZN(n16069) );
  XNOR2_X1 U26907 ( .A(n17297), .B(n16069), .ZN(n16070) );
  XNOR2_X1 U26908 ( .A(n16071), .B(n16070), .ZN(n16072) );
  XNOR2_X1 U26909 ( .A(n16073), .B(n16072), .ZN(n16074) );
  XNOR2_X1 U26910 ( .A(n16653), .B(n16074), .ZN(n16077) );
  XNOR2_X1 U26911 ( .A(n16075), .B(n18604), .ZN(n16076) );
  XNOR2_X1 U26912 ( .A(n18476), .B(n16294), .ZN(n16078) );
  XNOR2_X1 U26913 ( .A(n16078), .B(n16781), .ZN(n16080) );
  XNOR2_X1 U26914 ( .A(n16080), .B(n16079), .ZN(n16090) );
  XNOR2_X1 U26915 ( .A(n18689), .B(n18831), .ZN(n16086) );
  XNOR2_X1 U26916 ( .A(n4823), .B(n4518), .ZN(n16297) );
  XNOR2_X1 U26917 ( .A(n16297), .B(n4486), .ZN(n16081) );
  XNOR2_X1 U26918 ( .A(n33467), .B(n16081), .ZN(n16083) );
  XNOR2_X1 U26919 ( .A(n16082), .B(n4864), .ZN(n22453) );
  XNOR2_X1 U26920 ( .A(n22453), .B(n33474), .ZN(n43769) );
  XNOR2_X1 U26921 ( .A(n16083), .B(n43769), .ZN(n16084) );
  XNOR2_X1 U26922 ( .A(n18475), .B(n16084), .ZN(n16085) );
  XNOR2_X1 U26923 ( .A(n16086), .B(n16085), .ZN(n16088) );
  XNOR2_X1 U26924 ( .A(n18690), .B(n34377), .ZN(n16087) );
  INV_X1 U26925 ( .A(n18126), .ZN(n18826) );
  XNOR2_X1 U26926 ( .A(n16087), .B(n18826), .ZN(n16352) );
  XNOR2_X1 U26927 ( .A(n16088), .B(n16352), .ZN(n16089) );
  XNOR2_X1 U26928 ( .A(n16090), .B(n16089), .ZN(n16095) );
  XNOR2_X1 U26929 ( .A(n17954), .B(n16660), .ZN(n16091) );
  XNOR2_X1 U26930 ( .A(n16091), .B(n15619), .ZN(n16092) );
  XNOR2_X1 U26931 ( .A(n16092), .B(n18701), .ZN(n17278) );
  XNOR2_X1 U26932 ( .A(n16093), .B(n17278), .ZN(n16094) );
  NAND2_X1 U26933 ( .A1(n20611), .A2(n21513), .ZN(n16111) );
  XNOR2_X1 U26934 ( .A(n17321), .B(n51758), .ZN(n16255) );
  XNOR2_X1 U26935 ( .A(n2181), .B(n16255), .ZN(n16097) );
  XNOR2_X1 U26936 ( .A(n16096), .B(n16097), .ZN(n16101) );
  XNOR2_X1 U26937 ( .A(n16099), .B(n16098), .ZN(n16100) );
  XNOR2_X1 U26938 ( .A(n16101), .B(n16100), .ZN(n16110) );
  XNOR2_X1 U26939 ( .A(n24227), .B(n24828), .ZN(n18527) );
  XNOR2_X1 U26940 ( .A(n24894), .B(n26541), .ZN(n16103) );
  INV_X1 U26941 ( .A(n33653), .ZN(n16102) );
  XNOR2_X1 U26942 ( .A(n16103), .B(n16102), .ZN(n16976) );
  XNOR2_X1 U26943 ( .A(n18527), .B(n16976), .ZN(n34480) );
  XNOR2_X1 U26944 ( .A(n24695), .B(n25795), .ZN(n33543) );
  XNOR2_X1 U26945 ( .A(n34480), .B(n33543), .ZN(n16104) );
  XNOR2_X1 U26946 ( .A(n16105), .B(n16104), .ZN(n16106) );
  XNOR2_X1 U26947 ( .A(n2162), .B(n16106), .ZN(n16107) );
  XNOR2_X1 U26948 ( .A(n16107), .B(n16973), .ZN(n16108) );
  XNOR2_X1 U26949 ( .A(n18664), .B(n16108), .ZN(n16109) );
  XNOR2_X1 U26951 ( .A(n24200), .B(n33049), .ZN(n36824) );
  XNOR2_X1 U26952 ( .A(n36824), .B(n4637), .ZN(n41831) );
  XNOR2_X1 U26953 ( .A(n16112), .B(n43863), .ZN(n24396) );
  XNOR2_X1 U26954 ( .A(n41831), .B(n24396), .ZN(n35743) );
  XNOR2_X1 U26955 ( .A(n35107), .B(n4579), .ZN(n16113) );
  XNOR2_X1 U26956 ( .A(n33297), .B(n16113), .ZN(n16114) );
  XNOR2_X1 U26957 ( .A(n35743), .B(n16114), .ZN(n16115) );
  XNOR2_X1 U26958 ( .A(n2136), .B(n16115), .ZN(n16116) );
  XNOR2_X1 U26959 ( .A(n16116), .B(n543), .ZN(n16117) );
  XNOR2_X1 U26960 ( .A(n16117), .B(n19211), .ZN(n16123) );
  XNOR2_X1 U26961 ( .A(n16118), .B(n16321), .ZN(n16121) );
  XNOR2_X1 U26962 ( .A(n19196), .B(n19199), .ZN(n16119) );
  XNOR2_X1 U26963 ( .A(n16119), .B(n18407), .ZN(n16120) );
  XNOR2_X1 U26964 ( .A(n16121), .B(n16120), .ZN(n16122) );
  XNOR2_X1 U26965 ( .A(n16123), .B(n16122), .ZN(n16124) );
  NAND2_X1 U26966 ( .A1(n20175), .A2(n21528), .ZN(n16128) );
  NAND2_X1 U26967 ( .A1(n51050), .A2(n20614), .ZN(n16863) );
  INV_X1 U26968 ( .A(n21521), .ZN(n16127) );
  NAND2_X1 U26969 ( .A1(n23827), .A2(n23821), .ZN(n24151) );
  INV_X1 U26970 ( .A(n24151), .ZN(n16130) );
  INV_X1 U26971 ( .A(n24146), .ZN(n16129) );
  OAI21_X1 U26972 ( .B1(n24148), .B2(n16130), .A(n16129), .ZN(n16134) );
  NAND2_X1 U26973 ( .A1(n23835), .A2(n23834), .ZN(n16133) );
  NAND2_X1 U26974 ( .A1(n23834), .A2(n23832), .ZN(n20587) );
  INV_X1 U26975 ( .A(n20587), .ZN(n16131) );
  NAND2_X1 U26976 ( .A1(n16131), .A2(n23271), .ZN(n16132) );
  XNOR2_X1 U26977 ( .A(n16136), .B(n4939), .ZN(n42215) );
  XNOR2_X1 U26978 ( .A(n28307), .B(n4517), .ZN(n24640) );
  XOR2_X1 U26979 ( .A(n4886), .B(n4723), .Z(n16137) );
  XNOR2_X1 U26980 ( .A(n24640), .B(n16137), .ZN(n32276) );
  XNOR2_X1 U26981 ( .A(n32276), .B(n49429), .ZN(n16138) );
  XNOR2_X1 U26982 ( .A(n42215), .B(n16138), .ZN(n16139) );
  XNOR2_X1 U26983 ( .A(n16140), .B(n16139), .ZN(n16141) );
  XNOR2_X1 U26984 ( .A(n2226), .B(n16141), .ZN(n16145) );
  INV_X1 U26985 ( .A(n18580), .ZN(n16144) );
  XNOR2_X1 U26986 ( .A(n17364), .B(n4817), .ZN(n16143) );
  XNOR2_X1 U26987 ( .A(n16144), .B(n16143), .ZN(n16467) );
  XNOR2_X1 U26988 ( .A(n16467), .B(n16145), .ZN(n16146) );
  XNOR2_X1 U26989 ( .A(n485), .B(n16471), .ZN(n18801) );
  XNOR2_X1 U26990 ( .A(n16147), .B(n18801), .ZN(n16148) );
  XNOR2_X1 U26991 ( .A(n4177), .B(n4668), .ZN(n18556) );
  XNOR2_X1 U26992 ( .A(n4649), .B(n4884), .ZN(n16596) );
  XNOR2_X1 U26993 ( .A(n18556), .B(n16596), .ZN(n26526) );
  XNOR2_X1 U26994 ( .A(n16149), .B(n1313), .ZN(n18440) );
  XNOR2_X1 U26995 ( .A(n26526), .B(n18440), .ZN(n16151) );
  XNOR2_X1 U26996 ( .A(n27186), .B(n27353), .ZN(n34266) );
  INV_X1 U26997 ( .A(n34266), .ZN(n16150) );
  XNOR2_X1 U26998 ( .A(n16151), .B(n16150), .ZN(n37275) );
  XNOR2_X1 U26999 ( .A(n35815), .B(n4612), .ZN(n42918) );
  XNOR2_X1 U27000 ( .A(n42918), .B(n4653), .ZN(n42845) );
  XNOR2_X1 U27001 ( .A(n42845), .B(n32856), .ZN(n16152) );
  XNOR2_X1 U27002 ( .A(n37275), .B(n16152), .ZN(n16153) );
  XNOR2_X1 U27003 ( .A(n16711), .B(n16153), .ZN(n16154) );
  XNOR2_X1 U27004 ( .A(n17348), .B(n16154), .ZN(n16155) );
  XNOR2_X1 U27005 ( .A(n18820), .B(n16155), .ZN(n16157) );
  XNOR2_X1 U27006 ( .A(n18196), .B(n16156), .ZN(n16231) );
  XNOR2_X1 U27007 ( .A(n16157), .B(n16231), .ZN(n16161) );
  XNOR2_X1 U27008 ( .A(n17798), .B(n16158), .ZN(n16159) );
  XNOR2_X1 U27009 ( .A(n17261), .B(n16159), .ZN(n16160) );
  INV_X1 U27010 ( .A(n20062), .ZN(n16217) );
  XNOR2_X1 U27011 ( .A(n16749), .B(n18168), .ZN(n16163) );
  XNOR2_X1 U27012 ( .A(n16163), .B(n16162), .ZN(n18774) );
  XNOR2_X1 U27013 ( .A(n18181), .B(n18774), .ZN(n16170) );
  XNOR2_X1 U27014 ( .A(n26541), .B(n4665), .ZN(n35672) );
  XNOR2_X1 U27015 ( .A(n35672), .B(n44330), .ZN(n16166) );
  XNOR2_X1 U27016 ( .A(n16164), .B(n274), .ZN(n16165) );
  XNOR2_X1 U27017 ( .A(n16165), .B(n27483), .ZN(n34298) );
  XNOR2_X1 U27018 ( .A(n16166), .B(n34298), .ZN(n16167) );
  XNOR2_X1 U27019 ( .A(n33445), .B(n16167), .ZN(n16168) );
  XNOR2_X1 U27020 ( .A(n51031), .B(n16168), .ZN(n16169) );
  XNOR2_X1 U27021 ( .A(n16613), .B(n16428), .ZN(n16171) );
  XNOR2_X1 U27022 ( .A(n16172), .B(n18540), .ZN(n16173) );
  XNOR2_X1 U27023 ( .A(n16330), .B(n16173), .ZN(n16508) );
  XNOR2_X1 U27024 ( .A(n52167), .B(n18658), .ZN(n16427) );
  XNOR2_X1 U27025 ( .A(n16427), .B(n51373), .ZN(n16261) );
  XNOR2_X1 U27026 ( .A(n16508), .B(n16261), .ZN(n16174) );
  XNOR2_X1 U27027 ( .A(n16175), .B(n16174), .ZN(n16214) );
  INV_X1 U27028 ( .A(n26586), .ZN(n16177) );
  XNOR2_X1 U27029 ( .A(n26244), .B(n16177), .ZN(n21830) );
  XNOR2_X1 U27030 ( .A(n28085), .B(n4237), .ZN(n27301) );
  XNOR2_X1 U27031 ( .A(n44483), .B(n4803), .ZN(n16178) );
  XNOR2_X1 U27032 ( .A(n27301), .B(n16178), .ZN(n33406) );
  XNOR2_X1 U27033 ( .A(n21830), .B(n33406), .ZN(n16179) );
  XNOR2_X1 U27034 ( .A(n16666), .B(n16179), .ZN(n16180) );
  XNOR2_X1 U27035 ( .A(n16180), .B(n17731), .ZN(n16181) );
  XNOR2_X1 U27036 ( .A(n27297), .B(n4204), .ZN(n24484) );
  XNOR2_X1 U27037 ( .A(n2601), .B(n4585), .ZN(n21831) );
  XNOR2_X1 U27038 ( .A(n24484), .B(n21831), .ZN(n34216) );
  XNOR2_X1 U27039 ( .A(n15619), .B(n34216), .ZN(n16182) );
  XNOR2_X1 U27040 ( .A(n566), .B(n16182), .ZN(n16184) );
  XNOR2_X1 U27041 ( .A(n16183), .B(n16184), .ZN(n16442) );
  XNOR2_X1 U27042 ( .A(n16442), .B(n16185), .ZN(n16188) );
  XNOR2_X1 U27043 ( .A(n16770), .B(n18828), .ZN(n16356) );
  XNOR2_X1 U27044 ( .A(n17284), .B(n16356), .ZN(n16187) );
  XNOR2_X1 U27045 ( .A(n16188), .B(n16187), .ZN(n19140) );
  INV_X1 U27046 ( .A(n19140), .ZN(n20067) );
  XNOR2_X1 U27047 ( .A(n17378), .B(n17381), .ZN(n16189) );
  XNOR2_X1 U27048 ( .A(n16189), .B(n16485), .ZN(n16287) );
  XNOR2_X1 U27049 ( .A(n18466), .B(n47268), .ZN(n16191) );
  XNOR2_X1 U27050 ( .A(n16191), .B(n19261), .ZN(n16192) );
  XNOR2_X1 U27051 ( .A(n51417), .B(n16192), .ZN(n16486) );
  XNOR2_X1 U27052 ( .A(n27316), .B(n25284), .ZN(n33490) );
  XNOR2_X1 U27053 ( .A(n28071), .B(n4818), .ZN(n16281) );
  XNOR2_X1 U27054 ( .A(n33490), .B(n16281), .ZN(n43252) );
  XNOR2_X1 U27055 ( .A(n4926), .B(n4065), .ZN(n18745) );
  XNOR2_X1 U27056 ( .A(n26178), .B(n18745), .ZN(n25705) );
  XNOR2_X1 U27057 ( .A(n25705), .B(n4667), .ZN(n37258) );
  XNOR2_X1 U27058 ( .A(n43252), .B(n37258), .ZN(n16193) );
  XNOR2_X1 U27059 ( .A(n52141), .B(n16193), .ZN(n16194) );
  XNOR2_X1 U27060 ( .A(n18749), .B(n16194), .ZN(n16196) );
  XNOR2_X1 U27061 ( .A(n2230), .B(n4782), .ZN(n36854) );
  XNOR2_X1 U27062 ( .A(n51378), .B(n36854), .ZN(n16195) );
  XNOR2_X1 U27063 ( .A(n16195), .B(n17821), .ZN(n16762) );
  XNOR2_X1 U27064 ( .A(n16196), .B(n16762), .ZN(n16197) );
  XNOR2_X1 U27065 ( .A(n16486), .B(n16197), .ZN(n16198) );
  INV_X1 U27066 ( .A(n20075), .ZN(n20071) );
  INV_X1 U27067 ( .A(n18148), .ZN(n16199) );
  XNOR2_X1 U27068 ( .A(n16200), .B(n16199), .ZN(n17226) );
  XNOR2_X1 U27069 ( .A(n17138), .B(n18157), .ZN(n16627) );
  XNOR2_X1 U27070 ( .A(n16201), .B(n16624), .ZN(n16202) );
  XNOR2_X1 U27071 ( .A(n16627), .B(n16202), .ZN(n16207) );
  XNOR2_X1 U27072 ( .A(n43368), .B(n4312), .ZN(n35377) );
  XNOR2_X1 U27073 ( .A(n35377), .B(n45106), .ZN(n43020) );
  XNOR2_X1 U27074 ( .A(n4638), .B(n45883), .ZN(n31129) );
  XNOR2_X1 U27075 ( .A(n43020), .B(n31129), .ZN(n34602) );
  XNOR2_X1 U27076 ( .A(n36739), .B(n4940), .ZN(n43746) );
  XNOR2_X1 U27077 ( .A(n34602), .B(n43746), .ZN(n16203) );
  XNOR2_X1 U27078 ( .A(n33049), .B(n4316), .ZN(n42241) );
  XNOR2_X1 U27079 ( .A(n43019), .B(n42241), .ZN(n43371) );
  XNOR2_X1 U27080 ( .A(n43371), .B(n4045), .ZN(n33731) );
  XNOR2_X1 U27081 ( .A(n16203), .B(n33731), .ZN(n16204) );
  XNOR2_X1 U27082 ( .A(n18404), .B(n16204), .ZN(n16205) );
  XNOR2_X1 U27083 ( .A(n17754), .B(n16205), .ZN(n16206) );
  XNOR2_X1 U27084 ( .A(n16207), .B(n16206), .ZN(n16208) );
  XNOR2_X1 U27085 ( .A(n17226), .B(n16208), .ZN(n16210) );
  NAND2_X1 U27086 ( .A1(n18303), .A2(n19141), .ZN(n20073) );
  NOR2_X1 U27087 ( .A1(n20073), .A2(n16211), .ZN(n16213) );
  NAND2_X1 U27088 ( .A1(n2101), .A2(n20067), .ZN(n20070) );
  NOR2_X1 U27089 ( .A1(n20070), .A2(n20075), .ZN(n16212) );
  NOR2_X1 U27091 ( .A1(n19487), .A2(n20067), .ZN(n16215) );
  AOI22_X1 U27093 ( .A1(n20061), .A2(n19143), .B1(n16215), .B2(n20063), .ZN(
        n19498) );
  AOI21_X1 U27094 ( .B1(n19135), .B2(n16218), .A(n20075), .ZN(n16216) );
  INV_X1 U27095 ( .A(n20061), .ZN(n18300) );
  OAI21_X1 U27096 ( .B1(n18300), .B2(n19487), .A(n19136), .ZN(n20055) );
  INV_X1 U27097 ( .A(n20070), .ZN(n17027) );
  NAND2_X1 U27098 ( .A1(n16224), .A2(n16223), .ZN(n18616) );
  XNOR2_X1 U27099 ( .A(n17661), .B(n26525), .ZN(n18190) );
  XNOR2_X1 U27100 ( .A(n18190), .B(n27351), .ZN(n46126) );
  XNOR2_X1 U27101 ( .A(n28284), .B(n3481), .ZN(n27185) );
  XNOR2_X1 U27102 ( .A(n4287), .B(n1313), .ZN(n22777) );
  XNOR2_X1 U27103 ( .A(n49937), .B(n4612), .ZN(n16225) );
  XNOR2_X1 U27104 ( .A(n22777), .B(n16225), .ZN(n16226) );
  XNOR2_X1 U27105 ( .A(n27185), .B(n16226), .ZN(n35328) );
  XNOR2_X1 U27106 ( .A(n46126), .B(n35328), .ZN(n16227) );
  XNOR2_X1 U27107 ( .A(n16228), .B(n16227), .ZN(n16229) );
  XNOR2_X1 U27108 ( .A(n16229), .B(n18616), .ZN(n16230) );
  XNOR2_X1 U27109 ( .A(n16232), .B(n16231), .ZN(n16236) );
  XNOR2_X1 U27110 ( .A(n17923), .B(n19235), .ZN(n17110) );
  XNOR2_X1 U27111 ( .A(n16233), .B(n17110), .ZN(n16604) );
  XNOR2_X1 U27112 ( .A(n16234), .B(n16604), .ZN(n16235) );
  XNOR2_X1 U27113 ( .A(n2226), .B(n556), .ZN(n16240) );
  XNOR2_X1 U27114 ( .A(n17652), .B(n16238), .ZN(n16239) );
  XNOR2_X1 U27115 ( .A(n16904), .B(n17643), .ZN(n18582) );
  XNOR2_X1 U27116 ( .A(n16241), .B(n18636), .ZN(n42342) );
  XNOR2_X1 U27117 ( .A(n42342), .B(n3014), .ZN(n25743) );
  XNOR2_X1 U27118 ( .A(n25743), .B(n4932), .ZN(n32940) );
  XNOR2_X1 U27119 ( .A(n4568), .B(n3276), .ZN(n27388) );
  XNOR2_X1 U27120 ( .A(n27174), .B(n27388), .ZN(n22616) );
  XNOR2_X1 U27121 ( .A(n22616), .B(n4939), .ZN(n37289) );
  XNOR2_X1 U27122 ( .A(n32940), .B(n37289), .ZN(n16242) );
  XNOR2_X1 U27123 ( .A(n17812), .B(n16242), .ZN(n16243) );
  XNOR2_X1 U27124 ( .A(n18582), .B(n16243), .ZN(n16245) );
  XNOR2_X1 U27125 ( .A(n18208), .B(n17365), .ZN(n16244) );
  XNOR2_X1 U27126 ( .A(n16245), .B(n16244), .ZN(n16246) );
  XNOR2_X1 U27127 ( .A(n24057), .B(n43293), .ZN(n19768) );
  XNOR2_X1 U27128 ( .A(n19768), .B(n28307), .ZN(n42339) );
  XNOR2_X1 U27129 ( .A(n16247), .B(n16248), .ZN(n16544) );
  INV_X1 U27130 ( .A(n16250), .ZN(n16258) );
  XNOR2_X1 U27131 ( .A(n16251), .B(n4705), .ZN(n24893) );
  XNOR2_X1 U27132 ( .A(n24893), .B(n25795), .ZN(n33245) );
  XNOR2_X1 U27133 ( .A(n21089), .B(n4931), .ZN(n34892) );
  XNOR2_X1 U27134 ( .A(n29662), .B(n4542), .ZN(n43054) );
  XNOR2_X1 U27135 ( .A(n34892), .B(n43054), .ZN(n16252) );
  XNOR2_X1 U27136 ( .A(n33245), .B(n16252), .ZN(n16253) );
  XNOR2_X1 U27137 ( .A(n16416), .B(n16253), .ZN(n16254) );
  XNOR2_X1 U27138 ( .A(n49414), .B(n4578), .ZN(n34891) );
  XNOR2_X1 U27139 ( .A(n18773), .B(n34891), .ZN(n18661) );
  XNOR2_X1 U27140 ( .A(n16254), .B(n18661), .ZN(n16256) );
  INV_X1 U27141 ( .A(n16743), .ZN(n17897) );
  XNOR2_X1 U27142 ( .A(n16255), .B(n17897), .ZN(n16339) );
  XNOR2_X1 U27143 ( .A(n16256), .B(n16339), .ZN(n16257) );
  XNOR2_X1 U27144 ( .A(n16258), .B(n16257), .ZN(n16263) );
  INV_X1 U27145 ( .A(n16259), .ZN(n16260) );
  XNOR2_X1 U27146 ( .A(n16261), .B(n16260), .ZN(n16262) );
  INV_X1 U27147 ( .A(n17081), .ZN(n19482) );
  INV_X1 U27148 ( .A(n16264), .ZN(n18681) );
  XNOR2_X1 U27149 ( .A(n2136), .B(n17234), .ZN(n16265) );
  INV_X1 U27150 ( .A(n4157), .ZN(n49577) );
  XNOR2_X1 U27151 ( .A(n49577), .B(n4605), .ZN(n43922) );
  INV_X1 U27152 ( .A(n43922), .ZN(n26357) );
  XNOR2_X1 U27153 ( .A(n33930), .B(n26357), .ZN(n25236) );
  XNOR2_X1 U27154 ( .A(n42101), .B(n4045), .ZN(n43369) );
  XNOR2_X1 U27155 ( .A(n25236), .B(n43369), .ZN(n33430) );
  XNOR2_X1 U27156 ( .A(n4501), .B(n4343), .ZN(n34080) );
  XNOR2_X1 U27157 ( .A(n42816), .B(n34080), .ZN(n16266) );
  XNOR2_X1 U27158 ( .A(n44046), .B(n16266), .ZN(n16267) );
  XNOR2_X1 U27159 ( .A(n33430), .B(n16267), .ZN(n16268) );
  XNOR2_X1 U27160 ( .A(n18153), .B(n16268), .ZN(n16269) );
  XNOR2_X1 U27161 ( .A(n16270), .B(n16269), .ZN(n16271) );
  XNOR2_X1 U27162 ( .A(n16272), .B(n16271), .ZN(n16273) );
  XNOR2_X1 U27163 ( .A(n18681), .B(n16273), .ZN(n16278) );
  INV_X1 U27164 ( .A(n16730), .ZN(n18671) );
  XNOR2_X1 U27165 ( .A(n18671), .B(n17343), .ZN(n16277) );
  XNOR2_X1 U27166 ( .A(n18519), .B(n16498), .ZN(n16275) );
  XNOR2_X1 U27167 ( .A(n18669), .B(n17707), .ZN(n16274) );
  XNOR2_X1 U27168 ( .A(n16275), .B(n16274), .ZN(n16276) );
  XNOR2_X1 U27169 ( .A(n16277), .B(n16276), .ZN(n17144) );
  XNOR2_X1 U27170 ( .A(n16278), .B(n17144), .ZN(n16279) );
  INV_X1 U27171 ( .A(n16279), .ZN(n21248) );
  INV_X1 U27172 ( .A(n17079), .ZN(n21256) );
  NAND2_X1 U27173 ( .A1(n21256), .A2(n18969), .ZN(n17078) );
  XNOR2_X1 U27174 ( .A(n17691), .B(n4836), .ZN(n17385) );
  XNOR2_X1 U27175 ( .A(n17965), .B(n19260), .ZN(n17168) );
  XNOR2_X1 U27176 ( .A(n17385), .B(n17168), .ZN(n16285) );
  XNOR2_X1 U27177 ( .A(n23495), .B(n25616), .ZN(n42461) );
  XNOR2_X1 U27178 ( .A(n42461), .B(n26178), .ZN(n25371) );
  XNOR2_X1 U27179 ( .A(n25371), .B(n16280), .ZN(n44090) );
  XNOR2_X1 U27180 ( .A(n44090), .B(n4908), .ZN(n35363) );
  XNOR2_X1 U27181 ( .A(n4895), .B(n4721), .ZN(n22219) );
  XNOR2_X1 U27182 ( .A(n47268), .B(n4429), .ZN(n25170) );
  XNOR2_X1 U27183 ( .A(n22219), .B(n25170), .ZN(n25372) );
  XNOR2_X1 U27184 ( .A(n25372), .B(n16281), .ZN(n35497) );
  XNOR2_X1 U27185 ( .A(n35363), .B(n35497), .ZN(n16282) );
  XNOR2_X1 U27186 ( .A(n18739), .B(n16282), .ZN(n16283) );
  XNOR2_X1 U27187 ( .A(n16283), .B(n19261), .ZN(n16284) );
  XNOR2_X1 U27188 ( .A(n16285), .B(n16284), .ZN(n16286) );
  XNOR2_X1 U27189 ( .A(n16287), .B(n16286), .ZN(n16289) );
  XNOR2_X1 U27190 ( .A(n576), .B(n18591), .ZN(n16288) );
  XNOR2_X1 U27191 ( .A(n16288), .B(n17694), .ZN(n18146) );
  XNOR2_X1 U27192 ( .A(n16290), .B(n52183), .ZN(n16291) );
  XNOR2_X1 U27193 ( .A(n16568), .B(n566), .ZN(n17189) );
  XNOR2_X1 U27194 ( .A(n16291), .B(n17189), .ZN(n17398) );
  XNOR2_X1 U27195 ( .A(n16292), .B(n16661), .ZN(n16293) );
  XNOR2_X1 U27196 ( .A(n16293), .B(n51014), .ZN(n18700) );
  XNOR2_X1 U27197 ( .A(n16294), .B(n16660), .ZN(n16301) );
  XNOR2_X1 U27198 ( .A(n17180), .B(n28085), .ZN(n16296) );
  INV_X1 U27199 ( .A(n41460), .ZN(n16295) );
  XNOR2_X1 U27200 ( .A(n16296), .B(n16295), .ZN(n16572) );
  XNOR2_X1 U27201 ( .A(n16572), .B(n16297), .ZN(n34830) );
  XNOR2_X1 U27202 ( .A(n24484), .B(n26586), .ZN(n33200) );
  XNOR2_X1 U27203 ( .A(n4733), .B(n4628), .ZN(n33192) );
  XNOR2_X1 U27204 ( .A(n33200), .B(n33192), .ZN(n16298) );
  XNOR2_X1 U27205 ( .A(n34830), .B(n16298), .ZN(n16299) );
  XNOR2_X1 U27206 ( .A(n18126), .B(n16299), .ZN(n16300) );
  XNOR2_X1 U27207 ( .A(n16301), .B(n16300), .ZN(n16302) );
  XNOR2_X1 U27208 ( .A(n16302), .B(n18701), .ZN(n16303) );
  XNOR2_X1 U27209 ( .A(n18700), .B(n16303), .ZN(n16304) );
  XNOR2_X1 U27210 ( .A(n17398), .B(n16304), .ZN(n19086) );
  OAI211_X1 U27211 ( .C1(n17083), .C2(n21248), .A(n17078), .B(n21242), .ZN(
        n16312) );
  OR2_X1 U27212 ( .A1(n21248), .A2(n19086), .ZN(n21244) );
  NOR2_X1 U27213 ( .A1(n17081), .A2(n19086), .ZN(n16305) );
  OAI21_X1 U27214 ( .B1(n18962), .B2(n21244), .A(n16306), .ZN(n16307) );
  NAND2_X1 U27215 ( .A1(n16307), .A2(n3335), .ZN(n16311) );
  INV_X1 U27216 ( .A(n19087), .ZN(n19099) );
  OAI211_X1 U27217 ( .C1(n19099), .C2(n18963), .A(n19093), .B(n16308), .ZN(
        n16309) );
  AND2_X1 U27218 ( .A1(n21251), .A2(n19086), .ZN(n21249) );
  NAND2_X1 U27219 ( .A1(n16309), .A2(n21249), .ZN(n16310) );
  XNOR2_X1 U27220 ( .A(Key[3]), .B(n2117), .ZN(n18154) );
  XNOR2_X1 U27221 ( .A(n18154), .B(n4316), .ZN(n16314) );
  XNOR2_X1 U27222 ( .A(n16314), .B(n33049), .ZN(n16316) );
  INV_X1 U27223 ( .A(n33635), .ZN(n16404) );
  XNOR2_X1 U27224 ( .A(n16404), .B(n45107), .ZN(n16315) );
  XNOR2_X1 U27225 ( .A(n16316), .B(n16315), .ZN(n16317) );
  XNOR2_X1 U27226 ( .A(n24200), .B(n4868), .ZN(n39718) );
  XNOR2_X1 U27227 ( .A(n16317), .B(n39718), .ZN(n35466) );
  XNOR2_X1 U27228 ( .A(n35466), .B(n35377), .ZN(n16318) );
  XNOR2_X1 U27229 ( .A(n17763), .B(n16318), .ZN(n16319) );
  XNOR2_X1 U27230 ( .A(n16320), .B(n16319), .ZN(n16322) );
  XNOR2_X1 U27231 ( .A(n16321), .B(n16322), .ZN(n16325) );
  XNOR2_X1 U27232 ( .A(n51438), .B(n16323), .ZN(n16324) );
  XNOR2_X1 U27233 ( .A(n17891), .B(n17138), .ZN(n16326) );
  XNOR2_X1 U27234 ( .A(n16326), .B(n18505), .ZN(n16327) );
  XNOR2_X1 U27235 ( .A(n16327), .B(n18162), .ZN(n16727) );
  XNOR2_X1 U27236 ( .A(n2180), .B(n16749), .ZN(n16331) );
  XNOR2_X1 U27237 ( .A(n16331), .B(n16330), .ZN(n18538) );
  XNOR2_X1 U27238 ( .A(n25115), .B(n26297), .ZN(n34366) );
  XNOR2_X1 U27239 ( .A(n24828), .B(n4035), .ZN(n28266) );
  XNOR2_X1 U27240 ( .A(n4847), .B(n4597), .ZN(n44329) );
  XNOR2_X1 U27241 ( .A(n33653), .B(n44329), .ZN(n16332) );
  XNOR2_X1 U27242 ( .A(n28266), .B(n16332), .ZN(n16333) );
  XNOR2_X1 U27243 ( .A(n34366), .B(n16333), .ZN(n16334) );
  XNOR2_X1 U27244 ( .A(n16334), .B(n25576), .ZN(n16335) );
  XNOR2_X1 U27245 ( .A(n17901), .B(n16335), .ZN(n16336) );
  XNOR2_X1 U27246 ( .A(n16336), .B(n17213), .ZN(n16338) );
  XNOR2_X1 U27247 ( .A(n16338), .B(n51032), .ZN(n16340) );
  XNOR2_X1 U27248 ( .A(n16340), .B(n16339), .ZN(n16341) );
  XNOR2_X1 U27249 ( .A(n18538), .B(n16341), .ZN(n16343) );
  XNOR2_X1 U27250 ( .A(n16342), .B(n16343), .ZN(n20028) );
  XNOR2_X1 U27251 ( .A(n18701), .B(n51454), .ZN(n16344) );
  XNOR2_X1 U27252 ( .A(n16345), .B(n16344), .ZN(n16355) );
  XNOR2_X1 U27253 ( .A(n16346), .B(n17731), .ZN(n16351) );
  XNOR2_X1 U27254 ( .A(n17950), .B(n4654), .ZN(n39976) );
  XNOR2_X1 U27255 ( .A(n27297), .B(n4275), .ZN(n41426) );
  XNOR2_X1 U27256 ( .A(n39976), .B(n41426), .ZN(n34379) );
  XOR2_X1 U27257 ( .A(n4823), .B(n5016), .Z(n16347) );
  XNOR2_X1 U27258 ( .A(n33589), .B(n16347), .ZN(n16348) );
  XNOR2_X1 U27259 ( .A(n34379), .B(n16348), .ZN(n16349) );
  XNOR2_X1 U27260 ( .A(n18119), .B(n16349), .ZN(n16350) );
  XNOR2_X1 U27261 ( .A(n16351), .B(n16350), .ZN(n16353) );
  XNOR2_X1 U27262 ( .A(n16353), .B(n16352), .ZN(n16354) );
  XNOR2_X1 U27263 ( .A(n16355), .B(n16354), .ZN(n16359) );
  INV_X1 U27264 ( .A(n16356), .ZN(n16357) );
  XNOR2_X1 U27265 ( .A(n16658), .B(n16781), .ZN(n17963) );
  XNOR2_X1 U27266 ( .A(n16357), .B(n17963), .ZN(n16358) );
  XNOR2_X1 U27268 ( .A(n16361), .B(n16360), .ZN(n16371) );
  XNOR2_X1 U27269 ( .A(n51757), .B(n17798), .ZN(n18559) );
  INV_X1 U27270 ( .A(n18559), .ZN(n16369) );
  XNOR2_X1 U27271 ( .A(n18437), .B(n16450), .ZN(n16365) );
  XNOR2_X1 U27272 ( .A(n25651), .B(n24861), .ZN(n16599) );
  INV_X1 U27273 ( .A(n16599), .ZN(n25095) );
  XNOR2_X1 U27274 ( .A(n28390), .B(n4535), .ZN(n42026) );
  XNOR2_X1 U27275 ( .A(n25095), .B(n42026), .ZN(n36720) );
  XNOR2_X1 U27276 ( .A(n45051), .B(n4668), .ZN(n32267) );
  XNOR2_X1 U27277 ( .A(n34265), .B(n4627), .ZN(n16362) );
  XNOR2_X1 U27278 ( .A(n32267), .B(n16362), .ZN(n16363) );
  XNOR2_X1 U27279 ( .A(n36720), .B(n16363), .ZN(n16364) );
  XNOR2_X1 U27280 ( .A(n16365), .B(n16364), .ZN(n16367) );
  XNOR2_X1 U27281 ( .A(n16711), .B(n51135), .ZN(n16366) );
  XNOR2_X1 U27282 ( .A(n16367), .B(n16366), .ZN(n16368) );
  XNOR2_X1 U27283 ( .A(n16369), .B(n16368), .ZN(n16370) );
  XNOR2_X1 U27284 ( .A(n16371), .B(n16370), .ZN(n16395) );
  XNOR2_X1 U27285 ( .A(n16470), .B(n18427), .ZN(n17116) );
  XNOR2_X1 U27286 ( .A(n16372), .B(n17116), .ZN(n16374) );
  XNOR2_X1 U27287 ( .A(n16374), .B(n557), .ZN(n16706) );
  XNOR2_X1 U27288 ( .A(n28303), .B(n17243), .ZN(n35541) );
  INV_X1 U27289 ( .A(n35796), .ZN(n16899) );
  XNOR2_X1 U27290 ( .A(n16899), .B(n27174), .ZN(n45253) );
  XNOR2_X1 U27291 ( .A(n35541), .B(n45253), .ZN(n34850) );
  XNOR2_X1 U27292 ( .A(n25640), .B(n42668), .ZN(n16375) );
  XNOR2_X1 U27293 ( .A(n17121), .B(n16375), .ZN(n33228) );
  XNOR2_X1 U27294 ( .A(n33228), .B(n4558), .ZN(n16376) );
  XNOR2_X1 U27295 ( .A(n34850), .B(n16376), .ZN(n16377) );
  XNOR2_X1 U27296 ( .A(n16464), .B(n16377), .ZN(n16378) );
  XNOR2_X1 U27297 ( .A(n16532), .B(n16378), .ZN(n16379) );
  XNOR2_X1 U27298 ( .A(n17816), .B(n16379), .ZN(n16380) );
  XNOR2_X1 U27299 ( .A(n16706), .B(n16380), .ZN(n16382) );
  NAND2_X1 U27300 ( .A1(n16821), .A2(n18380), .ZN(n16814) );
  XNOR2_X1 U27301 ( .A(n16384), .B(n16383), .ZN(n16390) );
  INV_X1 U27302 ( .A(n42539), .ZN(n26180) );
  XNOR2_X1 U27303 ( .A(n26180), .B(n41367), .ZN(n16646) );
  INV_X1 U27304 ( .A(n16646), .ZN(n26259) );
  XNOR2_X1 U27305 ( .A(n42327), .B(n4934), .ZN(n26257) );
  XNOR2_X1 U27306 ( .A(n28070), .B(n4529), .ZN(n16755) );
  XNOR2_X1 U27307 ( .A(n26257), .B(n16755), .ZN(n16557) );
  XNOR2_X1 U27308 ( .A(n26259), .B(n16557), .ZN(n31595) );
  XNOR2_X1 U27309 ( .A(n16385), .B(n44493), .ZN(n36682) );
  XNOR2_X1 U27310 ( .A(n31595), .B(n36682), .ZN(n16386) );
  XNOR2_X1 U27311 ( .A(n16754), .B(n16386), .ZN(n16387) );
  XNOR2_X1 U27312 ( .A(n52141), .B(n16387), .ZN(n16388) );
  XNOR2_X1 U27313 ( .A(n16390), .B(n16389), .ZN(n16391) );
  INV_X1 U27314 ( .A(n20028), .ZN(n20037) );
  INV_X1 U27315 ( .A(n18380), .ZN(n20029) );
  NAND3_X1 U27316 ( .A1(n18381), .A2(n20042), .A3(n7585), .ZN(n16394) );
  INV_X1 U27317 ( .A(n17047), .ZN(n16820) );
  AND2_X1 U27318 ( .A1(n18377), .A2(n16820), .ZN(n20043) );
  NAND3_X1 U27319 ( .A1(n20043), .A2(n51440), .A3(n16814), .ZN(n16393) );
  NAND2_X1 U27320 ( .A1(n20046), .A2(n20027), .ZN(n16396) );
  AND2_X1 U27321 ( .A1(n5385), .A2(n20029), .ZN(n17456) );
  NOR2_X1 U27322 ( .A1(n17046), .A2(n5385), .ZN(n16824) );
  OAI211_X1 U27323 ( .C1(n16824), .C2(n51440), .A(n20032), .B(n16814), .ZN(
        n16398) );
  INV_X1 U27325 ( .A(n20042), .ZN(n16819) );
  XNOR2_X1 U27326 ( .A(n16400), .B(n18163), .ZN(n19209) );
  XNOR2_X1 U27327 ( .A(n51435), .B(n17763), .ZN(n16402) );
  XNOR2_X1 U27328 ( .A(n17138), .B(n17232), .ZN(n16401) );
  XNOR2_X1 U27329 ( .A(n16402), .B(n16401), .ZN(n16410) );
  XNOR2_X1 U27330 ( .A(n44934), .B(n4587), .ZN(n28375) );
  XNOR2_X1 U27331 ( .A(n28375), .B(n4045), .ZN(n16403) );
  XNOR2_X1 U27332 ( .A(n45883), .B(n4213), .ZN(n33733) );
  XNOR2_X1 U27333 ( .A(n33733), .B(n2117), .ZN(n42083) );
  XNOR2_X1 U27334 ( .A(n16403), .B(n42083), .ZN(n16405) );
  XNOR2_X1 U27335 ( .A(n42241), .B(n16404), .ZN(n28251) );
  XNOR2_X1 U27336 ( .A(n16405), .B(n28251), .ZN(n16406) );
  XNOR2_X1 U27337 ( .A(n28058), .B(n45106), .ZN(n42084) );
  XNOR2_X1 U27338 ( .A(n42084), .B(n4896), .ZN(n25132) );
  XNOR2_X1 U27339 ( .A(n16406), .B(n25132), .ZN(n16407) );
  XNOR2_X1 U27340 ( .A(n18157), .B(n16407), .ZN(n16408) );
  XNOR2_X1 U27341 ( .A(n16408), .B(n18408), .ZN(n16409) );
  XNOR2_X1 U27342 ( .A(n16410), .B(n16409), .ZN(n16411) );
  XNOR2_X1 U27343 ( .A(n19209), .B(n16411), .ZN(n16415) );
  XNOR2_X1 U27344 ( .A(n2099), .B(n18414), .ZN(n17344) );
  INV_X1 U27345 ( .A(n16412), .ZN(n16955) );
  XNOR2_X1 U27346 ( .A(n16722), .B(n16955), .ZN(n16413) );
  XNOR2_X1 U27347 ( .A(n17344), .B(n16413), .ZN(n16414) );
  XNOR2_X1 U27348 ( .A(n19213), .B(n17322), .ZN(n16417) );
  XNOR2_X1 U27349 ( .A(n18777), .B(n16416), .ZN(n18533) );
  INV_X1 U27350 ( .A(n18533), .ZN(n17221) );
  XNOR2_X1 U27351 ( .A(n16417), .B(n17221), .ZN(n16419) );
  INV_X1 U27352 ( .A(n17148), .ZN(n32658) );
  XNOR2_X1 U27353 ( .A(n32658), .B(n28271), .ZN(n24429) );
  XNOR2_X1 U27354 ( .A(n24429), .B(n4665), .ZN(n34057) );
  XNOR2_X1 U27355 ( .A(n16739), .B(n4597), .ZN(n16420) );
  XNOR2_X1 U27356 ( .A(n28266), .B(n16420), .ZN(n33808) );
  XNOR2_X1 U27357 ( .A(n34057), .B(n33808), .ZN(n16421) );
  XNOR2_X1 U27358 ( .A(n17208), .B(n16421), .ZN(n16423) );
  XNOR2_X1 U27359 ( .A(n16423), .B(n16422), .ZN(n16426) );
  XNOR2_X1 U27360 ( .A(n16743), .B(n3383), .ZN(n16615) );
  XNOR2_X1 U27361 ( .A(n18773), .B(n17218), .ZN(n16424) );
  XNOR2_X1 U27362 ( .A(n16615), .B(n16424), .ZN(n16425) );
  XNOR2_X1 U27363 ( .A(n16426), .B(n16425), .ZN(n16430) );
  XNOR2_X1 U27364 ( .A(n16428), .B(n16427), .ZN(n16429) );
  XNOR2_X1 U27365 ( .A(n16431), .B(n18696), .ZN(n16432) );
  XNOR2_X1 U27366 ( .A(n16432), .B(n16568), .ZN(n16773) );
  XNOR2_X1 U27367 ( .A(n42322), .B(n31432), .ZN(n25273) );
  XNOR2_X1 U27368 ( .A(n17181), .B(n25273), .ZN(n33201) );
  XNOR2_X1 U27369 ( .A(n33201), .B(n44483), .ZN(n33837) );
  XOR2_X1 U27370 ( .A(n4654), .B(n48814), .Z(n16433) );
  XNOR2_X1 U27371 ( .A(n33837), .B(n16433), .ZN(n16434) );
  XNOR2_X1 U27372 ( .A(n18119), .B(n16434), .ZN(n16436) );
  XNOR2_X1 U27373 ( .A(n16436), .B(n16435), .ZN(n16437) );
  XNOR2_X1 U27374 ( .A(n16438), .B(n16437), .ZN(n16439) );
  XNOR2_X1 U27375 ( .A(n16773), .B(n16439), .ZN(n16444) );
  XNOR2_X1 U27376 ( .A(n16661), .B(n47679), .ZN(n18485) );
  XNOR2_X1 U27377 ( .A(n17731), .B(n16666), .ZN(n16440) );
  XNOR2_X1 U27378 ( .A(n18485), .B(n16440), .ZN(n18836) );
  INV_X1 U27379 ( .A(n18836), .ZN(n16441) );
  XNOR2_X1 U27380 ( .A(n16442), .B(n16441), .ZN(n16443) );
  NOR2_X1 U27381 ( .A1(n19055), .A2(n19534), .ZN(n19044) );
  XNOR2_X1 U27382 ( .A(n18447), .B(n51642), .ZN(n16452) );
  XNOR2_X1 U27383 ( .A(n34265), .B(n2603), .ZN(n16446) );
  XNOR2_X1 U27384 ( .A(n32856), .B(n2602), .ZN(n16445) );
  XNOR2_X1 U27385 ( .A(n16446), .B(n16445), .ZN(n32270) );
  XNOR2_X1 U27386 ( .A(n32270), .B(n17254), .ZN(n45406) );
  XNOR2_X1 U27387 ( .A(n33221), .B(n4535), .ZN(n25538) );
  XNOR2_X1 U27388 ( .A(n22777), .B(n25538), .ZN(n27349) );
  XNOR2_X1 U27389 ( .A(n45406), .B(n27349), .ZN(n35068) );
  XOR2_X1 U27390 ( .A(n4649), .B(n4874), .Z(n16447) );
  XNOR2_X1 U27391 ( .A(n16447), .B(n35815), .ZN(n16448) );
  XNOR2_X1 U27392 ( .A(n35068), .B(n16448), .ZN(n16449) );
  XNOR2_X1 U27393 ( .A(n16450), .B(n16449), .ZN(n16451) );
  XNOR2_X1 U27394 ( .A(n16452), .B(n16451), .ZN(n16453) );
  INV_X1 U27395 ( .A(n16525), .ZN(n16457) );
  XNOR2_X1 U27396 ( .A(n2217), .B(n16457), .ZN(n16458) );
  XNOR2_X1 U27397 ( .A(n28307), .B(n4121), .ZN(n18637) );
  XNOR2_X1 U27398 ( .A(n19768), .B(n18637), .ZN(n16461) );
  XNOR2_X1 U27399 ( .A(n34575), .B(n2903), .ZN(n24059) );
  INV_X1 U27400 ( .A(n23370), .ZN(n16460) );
  XNOR2_X1 U27401 ( .A(n24059), .B(n16460), .ZN(n27385) );
  XNOR2_X1 U27402 ( .A(n16461), .B(n27385), .ZN(n31928) );
  XNOR2_X1 U27403 ( .A(n36698), .B(n4558), .ZN(n16462) );
  XNOR2_X1 U27404 ( .A(n31928), .B(n16462), .ZN(n16463) );
  XNOR2_X1 U27405 ( .A(n16464), .B(n16463), .ZN(n16465) );
  XNOR2_X1 U27406 ( .A(n16465), .B(n17125), .ZN(n16466) );
  XNOR2_X1 U27407 ( .A(n16467), .B(n16468), .ZN(n16474) );
  XNOR2_X1 U27408 ( .A(n16469), .B(n18795), .ZN(n16537) );
  XNOR2_X1 U27409 ( .A(n16472), .B(n16471), .ZN(n16584) );
  XNOR2_X1 U27410 ( .A(n16584), .B(n16537), .ZN(n16473) );
  XNOR2_X1 U27411 ( .A(n16474), .B(n16473), .ZN(n16475) );
  XNOR2_X1 U27412 ( .A(n4865), .B(n2230), .ZN(n42754) );
  XNOR2_X1 U27413 ( .A(n16476), .B(n42754), .ZN(n16477) );
  XNOR2_X1 U27414 ( .A(n16477), .B(n24612), .ZN(n22518) );
  XNOR2_X1 U27415 ( .A(n25616), .B(n4926), .ZN(n16478) );
  XNOR2_X1 U27416 ( .A(n22518), .B(n16478), .ZN(n35839) );
  XNOR2_X1 U27417 ( .A(n26257), .B(n4818), .ZN(n25172) );
  XNOR2_X1 U27418 ( .A(n25172), .B(n41367), .ZN(n35038) );
  XNOR2_X1 U27419 ( .A(n35839), .B(n35038), .ZN(n16479) );
  XNOR2_X1 U27420 ( .A(n18134), .B(n16479), .ZN(n16480) );
  XNOR2_X1 U27421 ( .A(n17288), .B(n16480), .ZN(n16482) );
  XNOR2_X1 U27422 ( .A(n18135), .B(n51379), .ZN(n16481) );
  XNOR2_X1 U27423 ( .A(n16482), .B(n16481), .ZN(n16483) );
  XNOR2_X1 U27424 ( .A(n16484), .B(n17175), .ZN(n16488) );
  XNOR2_X1 U27425 ( .A(n16485), .B(n17378), .ZN(n16763) );
  XNOR2_X1 U27426 ( .A(n16763), .B(n16486), .ZN(n16487) );
  AOI21_X1 U27427 ( .B1(n20124), .B2(n20114), .A(n20158), .ZN(n16489) );
  OAI22_X1 U27429 ( .A1(n17021), .A2(n20166), .B1(n20118), .B2(n52176), .ZN(
        n16492) );
  OAI211_X1 U27430 ( .C1(n16492), .C2(n16491), .A(n16490), .B(n19538), .ZN(
        n16495) );
  NOR2_X1 U27431 ( .A1(n20124), .A2(n51815), .ZN(n19050) );
  INV_X1 U27432 ( .A(n20124), .ZN(n19545) );
  XNOR2_X1 U27433 ( .A(n52190), .B(n16641), .ZN(n16497) );
  XNOR2_X1 U27434 ( .A(n16498), .B(n51435), .ZN(n16961) );
  INV_X1 U27435 ( .A(n16961), .ZN(n16499) );
  XNOR2_X1 U27436 ( .A(n16499), .B(n18523), .ZN(n16507) );
  XNOR2_X1 U27437 ( .A(n17891), .B(n18399), .ZN(n16506) );
  XNOR2_X1 U27438 ( .A(n42816), .B(n43368), .ZN(n16501) );
  XNOR2_X1 U27439 ( .A(Key[3]), .B(n4885), .ZN(n33529) );
  XNOR2_X1 U27440 ( .A(n33529), .B(n4587), .ZN(n16500) );
  XNOR2_X1 U27441 ( .A(n16501), .B(n16500), .ZN(n16502) );
  XNOR2_X1 U27442 ( .A(n16502), .B(n45105), .ZN(n16504) );
  XNOR2_X1 U27443 ( .A(n4739), .B(n4312), .ZN(n25022) );
  XNOR2_X1 U27444 ( .A(n44934), .B(n25022), .ZN(n33931) );
  XNOR2_X1 U27445 ( .A(n25470), .B(n33931), .ZN(n16503) );
  XNOR2_X1 U27446 ( .A(n543), .B(n17343), .ZN(n18152) );
  XNOR2_X1 U27447 ( .A(n2126), .B(n17213), .ZN(n16735) );
  XNOR2_X1 U27448 ( .A(n16735), .B(n16508), .ZN(n16519) );
  XNOR2_X1 U27449 ( .A(n16509), .B(n16608), .ZN(n44539) );
  XNOR2_X1 U27450 ( .A(n4597), .B(n4515), .ZN(n26289) );
  XNOR2_X1 U27451 ( .A(n26289), .B(n4752), .ZN(n18656) );
  XNOR2_X1 U27452 ( .A(n4706), .B(n4454), .ZN(n16510) );
  XNOR2_X1 U27453 ( .A(n24828), .B(n16510), .ZN(n16511) );
  XNOR2_X1 U27454 ( .A(n18656), .B(n16511), .ZN(n33316) );
  XNOR2_X1 U27455 ( .A(n33316), .B(n4639), .ZN(n16512) );
  XNOR2_X1 U27456 ( .A(n44539), .B(n16512), .ZN(n16513) );
  XNOR2_X1 U27457 ( .A(n51758), .B(n16513), .ZN(n16514) );
  XNOR2_X1 U27458 ( .A(n16973), .B(n16514), .ZN(n16515) );
  XNOR2_X1 U27459 ( .A(n51046), .B(n16515), .ZN(n16516) );
  XNOR2_X1 U27460 ( .A(n16517), .B(n16516), .ZN(n16518) );
  XNOR2_X1 U27461 ( .A(n16521), .B(n16520), .ZN(n16531) );
  XNOR2_X1 U27462 ( .A(n23943), .B(n4884), .ZN(n36717) );
  XNOR2_X1 U27463 ( .A(n44887), .B(n36717), .ZN(n16522) );
  XNOR2_X1 U27464 ( .A(n18190), .B(n16522), .ZN(n30526) );
  XNOR2_X1 U27465 ( .A(n42026), .B(n2604), .ZN(n37104) );
  XNOR2_X1 U27466 ( .A(n37104), .B(n4890), .ZN(n16523) );
  XNOR2_X1 U27467 ( .A(n30526), .B(n16523), .ZN(n16524) );
  XNOR2_X1 U27468 ( .A(n16525), .B(n16524), .ZN(n16526) );
  XNOR2_X1 U27469 ( .A(n18617), .B(n16526), .ZN(n16529) );
  XNOR2_X1 U27470 ( .A(n16527), .B(n17798), .ZN(n16528) );
  XNOR2_X1 U27471 ( .A(n16529), .B(n16528), .ZN(n16530) );
  NAND2_X1 U27472 ( .A1(n18352), .A2(n574), .ZN(n16566) );
  XNOR2_X1 U27473 ( .A(n16533), .B(n16534), .ZN(n16536) );
  XNOR2_X1 U27474 ( .A(n16535), .B(n16536), .ZN(n16538) );
  XNOR2_X1 U27475 ( .A(n4817), .B(n49323), .ZN(n25209) );
  XNOR2_X1 U27476 ( .A(n25209), .B(n47737), .ZN(n25148) );
  XNOR2_X1 U27477 ( .A(n4647), .B(n47401), .ZN(n42349) );
  XNOR2_X1 U27478 ( .A(n25148), .B(n42349), .ZN(n36977) );
  XNOR2_X1 U27479 ( .A(n34742), .B(n49429), .ZN(n16539) );
  XNOR2_X1 U27480 ( .A(n36977), .B(n16539), .ZN(n16540) );
  XNOR2_X1 U27481 ( .A(n17364), .B(n16540), .ZN(n16541) );
  XNOR2_X1 U27482 ( .A(n16541), .B(n17365), .ZN(n16542) );
  NAND2_X1 U27483 ( .A1(n16807), .A2(n574), .ZN(n19077) );
  NAND2_X1 U27484 ( .A1(n19077), .A2(n20147), .ZN(n20139) );
  NAND2_X1 U27485 ( .A1(n20135), .A2(n18362), .ZN(n16547) );
  NAND2_X1 U27486 ( .A1(n20139), .A2(n16547), .ZN(n16565) );
  INV_X1 U27487 ( .A(n35034), .ZN(n16548) );
  XNOR2_X1 U27488 ( .A(n18599), .B(n16548), .ZN(n16549) );
  XNOR2_X1 U27489 ( .A(n16549), .B(n51134), .ZN(n16550) );
  XNOR2_X1 U27490 ( .A(n16550), .B(n635), .ZN(n18709) );
  XNOR2_X1 U27491 ( .A(n17973), .B(n18712), .ZN(n16551) );
  XNOR2_X1 U27492 ( .A(n16551), .B(n560), .ZN(n16554) );
  XNOR2_X1 U27493 ( .A(n17690), .B(n18466), .ZN(n16552) );
  XNOR2_X1 U27494 ( .A(n18749), .B(n16552), .ZN(n16553) );
  XNOR2_X1 U27495 ( .A(n16554), .B(n16553), .ZN(n16555) );
  XNOR2_X1 U27496 ( .A(n18709), .B(n16555), .ZN(n16564) );
  XNOR2_X1 U27497 ( .A(n16754), .B(n52142), .ZN(n16933) );
  XNOR2_X1 U27498 ( .A(n25371), .B(n16556), .ZN(n37043) );
  XNOR2_X1 U27499 ( .A(n16557), .B(n49790), .ZN(n25988) );
  XNOR2_X1 U27500 ( .A(n37043), .B(n25988), .ZN(n16558) );
  XNOR2_X1 U27501 ( .A(n17829), .B(n16558), .ZN(n16560) );
  XNOR2_X1 U27502 ( .A(n16559), .B(n16560), .ZN(n16561) );
  XNOR2_X1 U27503 ( .A(n16933), .B(n16561), .ZN(n16562) );
  XNOR2_X1 U27504 ( .A(n17694), .B(n16562), .ZN(n16563) );
  MUX2_X1 U27505 ( .A(n16566), .B(n16565), .S(n52037), .Z(n16581) );
  NAND2_X1 U27506 ( .A1(n16546), .A2(n18346), .ZN(n19071) );
  NOR2_X1 U27507 ( .A1(n51756), .A2(n20134), .ZN(n16567) );
  XOR2_X1 U27508 ( .A(n4835), .B(n4275), .Z(n16569) );
  XNOR2_X1 U27509 ( .A(n21831), .B(n16569), .ZN(n43314) );
  XNOR2_X1 U27510 ( .A(n43314), .B(n4803), .ZN(n16570) );
  XNOR2_X1 U27511 ( .A(n16571), .B(n16570), .ZN(n16574) );
  INV_X1 U27512 ( .A(n16572), .ZN(n16573) );
  XNOR2_X1 U27513 ( .A(n16573), .B(n4237), .ZN(n33287) );
  XNOR2_X1 U27514 ( .A(n33287), .B(n4048), .ZN(n43881) );
  XNOR2_X1 U27515 ( .A(n16574), .B(n43881), .ZN(n16575) );
  NAND2_X1 U27516 ( .A1(n20132), .A2(n20134), .ZN(n20145) );
  NOR2_X1 U27517 ( .A1(n20145), .A2(n52037), .ZN(n16579) );
  NAND2_X1 U27518 ( .A1(n17071), .A2(n16579), .ZN(n16580) );
  XNOR2_X1 U27519 ( .A(n16582), .B(n17938), .ZN(n16583) );
  XNOR2_X1 U27520 ( .A(n16583), .B(n19244), .ZN(n16585) );
  XNOR2_X1 U27521 ( .A(n16585), .B(n16584), .ZN(n16591) );
  INV_X1 U27522 ( .A(n17360), .ZN(n16586) );
  XNOR2_X1 U27523 ( .A(n16586), .B(n28303), .ZN(n43552) );
  XNOR2_X1 U27524 ( .A(n43552), .B(n27388), .ZN(n37084) );
  XNOR2_X1 U27525 ( .A(n28307), .B(n4932), .ZN(n37082) );
  XNOR2_X1 U27526 ( .A(n24057), .B(n4723), .ZN(n16587) );
  XNOR2_X1 U27527 ( .A(n37082), .B(n16587), .ZN(n30953) );
  XNOR2_X1 U27528 ( .A(n37084), .B(n30953), .ZN(n16588) );
  XNOR2_X1 U27529 ( .A(n17118), .B(n16588), .ZN(n16589) );
  XNOR2_X1 U27530 ( .A(n16589), .B(n2225), .ZN(n16590) );
  XNOR2_X1 U27531 ( .A(n17356), .B(n18820), .ZN(n16595) );
  XNOR2_X1 U27532 ( .A(n51133), .B(n16593), .ZN(n16594) );
  XNOR2_X1 U27533 ( .A(n16595), .B(n16594), .ZN(n16606) );
  XNOR2_X1 U27534 ( .A(n18447), .B(n2200), .ZN(n16602) );
  XNOR2_X1 U27535 ( .A(n45051), .B(n4879), .ZN(n24972) );
  XNOR2_X1 U27536 ( .A(n24972), .B(n16596), .ZN(n35622) );
  XNOR2_X1 U27537 ( .A(n28390), .B(n7744), .ZN(n25094) );
  XNOR2_X1 U27538 ( .A(n25094), .B(n33221), .ZN(n16597) );
  XNOR2_X1 U27539 ( .A(n35622), .B(n16597), .ZN(n16598) );
  XNOR2_X1 U27540 ( .A(n16599), .B(n16598), .ZN(n16600) );
  XNOR2_X1 U27541 ( .A(n51135), .B(n16600), .ZN(n16601) );
  XNOR2_X1 U27542 ( .A(n16602), .B(n16601), .ZN(n16603) );
  XNOR2_X1 U27543 ( .A(n16603), .B(n51482), .ZN(n16605) );
  NAND2_X1 U27544 ( .A1(n21233), .A2(n16678), .ZN(n17412) );
  INV_X1 U27545 ( .A(n17412), .ZN(n21230) );
  XNOR2_X1 U27546 ( .A(n17158), .B(n18540), .ZN(n16612) );
  XNOR2_X1 U27547 ( .A(n33653), .B(n4536), .ZN(n25792) );
  XNOR2_X1 U27548 ( .A(n25792), .B(n4035), .ZN(n16607) );
  XNOR2_X1 U27549 ( .A(n25791), .B(n16607), .ZN(n34790) );
  XNOR2_X1 U27550 ( .A(n16608), .B(n26297), .ZN(n33949) );
  XNOR2_X1 U27551 ( .A(n33949), .B(n4665), .ZN(n16609) );
  XNOR2_X1 U27552 ( .A(n34790), .B(n16609), .ZN(n16610) );
  XNOR2_X1 U27553 ( .A(n16612), .B(n16611), .ZN(n16614) );
  XNOR2_X1 U27554 ( .A(n16613), .B(n16614), .ZN(n16619) );
  XNOR2_X1 U27555 ( .A(n18533), .B(n16615), .ZN(n16617) );
  XNOR2_X1 U27556 ( .A(n17146), .B(n18661), .ZN(n16616) );
  XNOR2_X1 U27557 ( .A(n16616), .B(n16617), .ZN(n16618) );
  XNOR2_X1 U27558 ( .A(n16618), .B(n16619), .ZN(n16623) );
  INV_X1 U27559 ( .A(n16620), .ZN(n16621) );
  XNOR2_X1 U27560 ( .A(n18394), .B(n16621), .ZN(n17916) );
  XNOR2_X1 U27561 ( .A(n51046), .B(n2214), .ZN(n16622) );
  XNOR2_X1 U27562 ( .A(n17916), .B(n16622), .ZN(n17327) );
  XNOR2_X1 U27563 ( .A(n17891), .B(n16624), .ZN(n16626) );
  XNOR2_X1 U27564 ( .A(n4316), .B(n4157), .ZN(n34424) );
  XNOR2_X1 U27565 ( .A(n19199), .B(n34424), .ZN(n16625) );
  INV_X1 U27566 ( .A(n18770), .ZN(n16637) );
  XNOR2_X1 U27567 ( .A(n16628), .B(n17763), .ZN(n16629) );
  XNOR2_X1 U27568 ( .A(n17879), .B(n16629), .ZN(n16957) );
  XNOR2_X1 U27569 ( .A(n18755), .B(n19203), .ZN(n16634) );
  XNOR2_X1 U27570 ( .A(n42101), .B(n4937), .ZN(n28252) );
  XNOR2_X1 U27571 ( .A(n28252), .B(n33635), .ZN(n45111) );
  XNOR2_X1 U27572 ( .A(n45111), .B(n4940), .ZN(n33299) );
  XNOR2_X1 U27573 ( .A(n45106), .B(n33733), .ZN(n41827) );
  XNOR2_X1 U27574 ( .A(n42816), .B(n4896), .ZN(n16630) );
  XNOR2_X1 U27575 ( .A(n41827), .B(n16630), .ZN(n34166) );
  XNOR2_X1 U27576 ( .A(n34166), .B(n33297), .ZN(n16631) );
  XNOR2_X1 U27577 ( .A(n33299), .B(n16631), .ZN(n16632) );
  XNOR2_X1 U27578 ( .A(n17707), .B(n16632), .ZN(n16633) );
  XNOR2_X1 U27579 ( .A(n16634), .B(n16633), .ZN(n16635) );
  XNOR2_X1 U27580 ( .A(n16635), .B(n16957), .ZN(n16636) );
  XNOR2_X1 U27581 ( .A(n16636), .B(n16637), .ZN(n16644) );
  XNOR2_X1 U27582 ( .A(n16720), .B(n14903), .ZN(n16639) );
  XNOR2_X1 U27583 ( .A(n2135), .B(n18407), .ZN(n16638) );
  XNOR2_X1 U27584 ( .A(n16639), .B(n16638), .ZN(n16642) );
  INV_X1 U27585 ( .A(n51668), .ZN(n16640) );
  XNOR2_X1 U27586 ( .A(n16641), .B(n16640), .ZN(n17334) );
  XNOR2_X1 U27587 ( .A(n16642), .B(n17334), .ZN(n16643) );
  XNOR2_X1 U27588 ( .A(n576), .B(n17168), .ZN(n16645) );
  XNOR2_X1 U27589 ( .A(n51379), .B(n18749), .ZN(n16652) );
  XNOR2_X1 U27590 ( .A(n4895), .B(n4930), .ZN(n17164) );
  XNOR2_X1 U27591 ( .A(n16646), .B(n17164), .ZN(n35592) );
  XNOR2_X1 U27592 ( .A(n42754), .B(n4908), .ZN(n28232) );
  XNOR2_X1 U27593 ( .A(n23495), .B(n18745), .ZN(n16647) );
  XNOR2_X1 U27594 ( .A(n28232), .B(n16647), .ZN(n35252) );
  XNOR2_X1 U27595 ( .A(n35252), .B(n23887), .ZN(n16648) );
  XNOR2_X1 U27596 ( .A(n35592), .B(n16648), .ZN(n16649) );
  XNOR2_X1 U27597 ( .A(n18747), .B(n16649), .ZN(n16650) );
  XNOR2_X1 U27598 ( .A(n17288), .B(n18599), .ZN(n19267) );
  XNOR2_X1 U27599 ( .A(n16653), .B(n19267), .ZN(n17968) );
  INV_X1 U27600 ( .A(n17968), .ZN(n16654) );
  NAND2_X1 U27601 ( .A1(n19512), .A2(n16655), .ZN(n16676) );
  XNOR2_X1 U27602 ( .A(n17950), .B(n43105), .ZN(n25271) );
  INV_X1 U27603 ( .A(n25866), .ZN(n16656) );
  XNOR2_X1 U27604 ( .A(n25271), .B(n16656), .ZN(n33914) );
  XNOR2_X1 U27605 ( .A(n17177), .B(n33914), .ZN(n16657) );
  XNOR2_X1 U27606 ( .A(n16658), .B(n16657), .ZN(n16659) );
  XNOR2_X1 U27607 ( .A(n16659), .B(n16781), .ZN(n17397) );
  XNOR2_X1 U27608 ( .A(n17959), .B(n17397), .ZN(n16672) );
  XNOR2_X1 U27609 ( .A(n16661), .B(n16660), .ZN(n18573) );
  XNOR2_X1 U27610 ( .A(n51703), .B(n18119), .ZN(n16663) );
  XNOR2_X1 U27611 ( .A(n16663), .B(n17281), .ZN(n16946) );
  XNOR2_X1 U27612 ( .A(n18573), .B(n16946), .ZN(n16670) );
  XNOR2_X1 U27613 ( .A(n47679), .B(n4502), .ZN(n44161) );
  XNOR2_X1 U27614 ( .A(n4803), .B(n4518), .ZN(n27247) );
  XNOR2_X1 U27615 ( .A(n44161), .B(n27247), .ZN(n43074) );
  XNOR2_X1 U27616 ( .A(n43074), .B(n42322), .ZN(n34729) );
  XNOR2_X1 U27617 ( .A(n33192), .B(n4237), .ZN(n16664) );
  XNOR2_X1 U27618 ( .A(n34729), .B(n16664), .ZN(n16665) );
  XNOR2_X1 U27619 ( .A(n16666), .B(n16665), .ZN(n16667) );
  XNOR2_X1 U27620 ( .A(n16667), .B(n17731), .ZN(n16668) );
  XNOR2_X1 U27621 ( .A(n18701), .B(n16668), .ZN(n16669) );
  XNOR2_X1 U27622 ( .A(n16670), .B(n16669), .ZN(n16671) );
  NAND3_X1 U27624 ( .A1(n19518), .A2(n770), .A3(n19503), .ZN(n16674) );
  AOI21_X1 U27625 ( .B1(n16676), .B2(n19503), .A(n16675), .ZN(n16686) );
  OAI22_X1 U27626 ( .A1(n21233), .A2(n19521), .B1(n21223), .B2(n21227), .ZN(
        n16680) );
  OAI22_X1 U27627 ( .A1(n21222), .A2(n19520), .B1(n21232), .B2(n21234), .ZN(
        n16679) );
  OAI21_X1 U27628 ( .B1(n16680), .B2(n16679), .A(n19504), .ZN(n16683) );
  MUX2_X1 U27629 ( .A(n21224), .B(n16681), .S(n17412), .Z(n16682) );
  AOI22_X1 U27632 ( .A1(n19110), .A2(n6226), .B1(n16684), .B2(n21235), .ZN(
        n16685) );
  OAI211_X1 U27634 ( .C1(n23160), .C2(n21948), .A(n21953), .B(n6010), .ZN(
        n16693) );
  AND2_X1 U27635 ( .A1(n21957), .A2(n51123), .ZN(n19590) );
  INV_X1 U27636 ( .A(n19590), .ZN(n16690) );
  NAND2_X1 U27637 ( .A1(n23467), .A2(n23157), .ZN(n16689) );
  NAND2_X1 U27638 ( .A1(n16690), .A2(n16689), .ZN(n16691) );
  NAND2_X1 U27639 ( .A1(n16691), .A2(n23465), .ZN(n16692) );
  XNOR2_X1 U27640 ( .A(n24057), .B(n4886), .ZN(n42740) );
  XNOR2_X1 U27641 ( .A(n17121), .B(n42740), .ZN(n16697) );
  XNOR2_X1 U27642 ( .A(n24640), .B(n23370), .ZN(n16696) );
  XNOR2_X1 U27643 ( .A(n16697), .B(n16696), .ZN(n33960) );
  XNOR2_X1 U27644 ( .A(n42349), .B(n4624), .ZN(n25210) );
  XNOR2_X1 U27645 ( .A(n25210), .B(n4746), .ZN(n16699) );
  XNOR2_X1 U27646 ( .A(n16699), .B(n16698), .ZN(n34743) );
  XNOR2_X1 U27647 ( .A(n33960), .B(n34743), .ZN(n16700) );
  XNOR2_X1 U27648 ( .A(n17936), .B(n16700), .ZN(n16702) );
  XNOR2_X1 U27649 ( .A(n16704), .B(n17365), .ZN(n17239) );
  XNOR2_X1 U27650 ( .A(n32270), .B(n32267), .ZN(n16709) );
  XNOR2_X1 U27651 ( .A(n7744), .B(n4890), .ZN(n16708) );
  XNOR2_X1 U27652 ( .A(n28116), .B(n16708), .ZN(n36803) );
  XNOR2_X1 U27653 ( .A(n16709), .B(n36803), .ZN(n16710) );
  XNOR2_X1 U27654 ( .A(n16711), .B(n51642), .ZN(n16712) );
  XNOR2_X1 U27655 ( .A(n16713), .B(n16712), .ZN(n16714) );
  XNOR2_X1 U27656 ( .A(n18446), .B(n16714), .ZN(n16716) );
  XNOR2_X1 U27657 ( .A(n16715), .B(n16716), .ZN(n16718) );
  XNOR2_X1 U27658 ( .A(n36741), .B(n4638), .ZN(n26356) );
  XNOR2_X1 U27659 ( .A(n26356), .B(n4451), .ZN(n42781) );
  XNOR2_X1 U27660 ( .A(n18399), .B(n42781), .ZN(n16725) );
  XNOR2_X1 U27661 ( .A(n35290), .B(n4316), .ZN(n44935) );
  XNOR2_X1 U27662 ( .A(n44935), .B(n4605), .ZN(n16723) );
  XNOR2_X1 U27663 ( .A(n14427), .B(n16723), .ZN(n16724) );
  XNOR2_X1 U27664 ( .A(n16725), .B(n16724), .ZN(n16726) );
  XNOR2_X1 U27665 ( .A(n16728), .B(n16727), .ZN(n16734) );
  XNOR2_X1 U27666 ( .A(n2099), .B(n16729), .ZN(n16731) );
  XNOR2_X1 U27667 ( .A(n16732), .B(n16731), .ZN(n16733) );
  XNOR2_X1 U27668 ( .A(n51046), .B(n19227), .ZN(n16736) );
  XNOR2_X1 U27669 ( .A(n16736), .B(n16735), .ZN(n16748) );
  XNOR2_X1 U27670 ( .A(n24229), .B(n4325), .ZN(n16738) );
  XNOR2_X1 U27671 ( .A(n16738), .B(n16737), .ZN(n34613) );
  XNOR2_X1 U27672 ( .A(n16739), .B(n4482), .ZN(n16740) );
  XNOR2_X1 U27673 ( .A(n16740), .B(n27364), .ZN(n33689) );
  XNOR2_X1 U27674 ( .A(n33689), .B(n274), .ZN(n16741) );
  XNOR2_X1 U27675 ( .A(n34613), .B(n16741), .ZN(n16742) );
  XNOR2_X1 U27676 ( .A(n18175), .B(n16742), .ZN(n16744) );
  XNOR2_X1 U27677 ( .A(n16743), .B(n16744), .ZN(n16745) );
  XNOR2_X1 U27678 ( .A(n16746), .B(n16745), .ZN(n16747) );
  XNOR2_X1 U27679 ( .A(n16748), .B(n16747), .ZN(n16753) );
  INV_X1 U27680 ( .A(n16749), .ZN(n16750) );
  XNOR2_X1 U27681 ( .A(n17208), .B(n16750), .ZN(n16752) );
  XNOR2_X1 U27682 ( .A(n17771), .B(n41223), .ZN(n16751) );
  XNOR2_X1 U27683 ( .A(n16752), .B(n16751), .ZN(n18397) );
  XNOR2_X1 U27684 ( .A(n16754), .B(n17690), .ZN(n16757) );
  XNOR2_X1 U27685 ( .A(n16755), .B(n4930), .ZN(n24610) );
  XNOR2_X1 U27686 ( .A(n24610), .B(n4824), .ZN(n24496) );
  XNOR2_X1 U27687 ( .A(n24496), .B(n4721), .ZN(n32341) );
  XNOR2_X1 U27688 ( .A(n36682), .B(n24612), .ZN(n36859) );
  XNOR2_X1 U27689 ( .A(n32341), .B(n36859), .ZN(n16756) );
  XNOR2_X1 U27690 ( .A(n16757), .B(n16756), .ZN(n16759) );
  XNOR2_X1 U27692 ( .A(n16762), .B(n16763), .ZN(n16764) );
  XNOR2_X1 U27693 ( .A(n576), .B(n16765), .ZN(n16766) );
  AND2_X1 U27694 ( .A1(n17498), .A2(n16767), .ZN(n16796) );
  INV_X1 U27695 ( .A(n19186), .ZN(n16768) );
  XNOR2_X1 U27696 ( .A(n16768), .B(n17731), .ZN(n16769) );
  XNOR2_X1 U27697 ( .A(n16769), .B(n566), .ZN(n16771) );
  XNOR2_X1 U27698 ( .A(n16770), .B(n16771), .ZN(n16772) );
  XNOR2_X1 U27699 ( .A(n16773), .B(n16772), .ZN(n16786) );
  XNOR2_X1 U27700 ( .A(n42322), .B(n4823), .ZN(n25521) );
  XNOR2_X1 U27701 ( .A(n44483), .B(n31432), .ZN(n16774) );
  XNOR2_X1 U27702 ( .A(n25521), .B(n16774), .ZN(n16776) );
  INV_X1 U27703 ( .A(n33589), .ZN(n16775) );
  XNOR2_X1 U27704 ( .A(n16776), .B(n16775), .ZN(n33749) );
  XNOR2_X1 U27705 ( .A(n33746), .B(n16777), .ZN(n34558) );
  XNOR2_X1 U27706 ( .A(n33749), .B(n34558), .ZN(n16778) );
  XNOR2_X1 U27707 ( .A(n17954), .B(n16778), .ZN(n16779) );
  XNOR2_X1 U27708 ( .A(n16779), .B(n18832), .ZN(n16780) );
  XNOR2_X1 U27709 ( .A(n16781), .B(n16780), .ZN(n16784) );
  XNOR2_X1 U27710 ( .A(n16782), .B(n18828), .ZN(n16783) );
  XNOR2_X1 U27711 ( .A(n16784), .B(n16783), .ZN(n16785) );
  XNOR2_X1 U27712 ( .A(n16786), .B(n16785), .ZN(n17499) );
  INV_X1 U27713 ( .A(n17499), .ZN(n20094) );
  INV_X1 U27714 ( .A(n20093), .ZN(n17505) );
  AND2_X1 U27715 ( .A1(n20094), .A2(n20095), .ZN(n20105) );
  INV_X1 U27716 ( .A(n18315), .ZN(n16787) );
  OAI211_X1 U27718 ( .C1(n17505), .C2(n20101), .A(n16790), .B(n16789), .ZN(
        n16791) );
  AND2_X1 U27719 ( .A1(n20100), .A2(n16792), .ZN(n17504) );
  INV_X1 U27720 ( .A(n17504), .ZN(n17600) );
  NAND2_X1 U27721 ( .A1(n16791), .A2(n17600), .ZN(n16795) );
  NAND2_X1 U27722 ( .A1(n20086), .A2(n18315), .ZN(n18312) );
  NAND3_X1 U27723 ( .A1(n18312), .A2(n16788), .A3(n20097), .ZN(n16793) );
  NAND2_X1 U27724 ( .A1(n16793), .A2(n18313), .ZN(n16794) );
  NAND4_X1 U27725 ( .A1(n590), .A2(n17489), .A3(n18287), .A4(n20021), .ZN(
        n20020) );
  INV_X1 U27726 ( .A(n18282), .ZN(n16799) );
  OAI21_X1 U27727 ( .B1(n16799), .B2(n16798), .A(n20013), .ZN(n16800) );
  INV_X1 U27728 ( .A(n18291), .ZN(n17529) );
  OR2_X1 U27729 ( .A1(n20014), .A2(n18294), .ZN(n20010) );
  NOR2_X1 U27730 ( .A1(n16807), .A2(n18344), .ZN(n16802) );
  NOR2_X1 U27731 ( .A1(n16802), .A2(n18360), .ZN(n16803) );
  NAND2_X1 U27732 ( .A1(n19076), .A2(n19077), .ZN(n17067) );
  NAND2_X1 U27733 ( .A1(n17067), .A2(n17065), .ZN(n16805) );
  NAND3_X1 U27734 ( .A1(n19076), .A2(n19061), .A3(n18352), .ZN(n19074) );
  NAND3_X1 U27735 ( .A1(n51403), .A2(n52037), .A3(n20132), .ZN(n20138) );
  NAND2_X1 U27736 ( .A1(n19071), .A2(n20138), .ZN(n16810) );
  AOI21_X1 U27737 ( .B1(n1416), .B2(n16808), .A(n52037), .ZN(n16809) );
  INV_X1 U27738 ( .A(n16811), .ZN(n16812) );
  NOR2_X1 U27739 ( .A1(n18383), .A2(n20028), .ZN(n16818) );
  NOR2_X1 U27740 ( .A1(n16814), .A2(n5881), .ZN(n16816) );
  INV_X1 U27741 ( .A(n16814), .ZN(n16823) );
  NOR2_X1 U27742 ( .A1(n16818), .A2(n16817), .ZN(n16832) );
  AND2_X1 U27743 ( .A1(n16820), .A2(n20029), .ZN(n17050) );
  NAND2_X1 U27744 ( .A1(n18376), .A2(n16821), .ZN(n17458) );
  INV_X1 U27745 ( .A(n16824), .ZN(n16825) );
  INV_X1 U27746 ( .A(n20027), .ZN(n20040) );
  AOI22_X1 U27747 ( .A1(n17049), .A2(n20045), .B1(n20040), .B2(n51440), .ZN(
        n16828) );
  NAND2_X1 U27748 ( .A1(n16823), .A2(n20042), .ZN(n16827) );
  NAND2_X1 U27749 ( .A1(n5881), .A2(n16820), .ZN(n17448) );
  NAND2_X1 U27750 ( .A1(n18064), .A2(n18070), .ZN(n16833) );
  OAI211_X1 U27751 ( .C1(n18326), .C2(n403), .A(n16833), .B(n18332), .ZN(
        n16839) );
  AOI22_X1 U27752 ( .A1(n18330), .A2(n17440), .B1(n18071), .B2(n17544), .ZN(
        n16838) );
  NAND2_X1 U27753 ( .A1(n17431), .A2(n18074), .ZN(n16837) );
  OAI211_X1 U27754 ( .C1(n772), .C2(n17542), .A(n18062), .B(n17545), .ZN(
        n16835) );
  OAI211_X1 U27755 ( .C1(n18074), .C2(n17542), .A(n18060), .B(n16835), .ZN(
        n16836) );
  INV_X1 U27756 ( .A(n19399), .ZN(n18025) );
  NAND2_X1 U27757 ( .A1(n18025), .A2(n19396), .ZN(n16840) );
  INV_X1 U27759 ( .A(n17484), .ZN(n17577) );
  INV_X1 U27760 ( .A(n18015), .ZN(n16844) );
  AOI22_X1 U27761 ( .A1(n16844), .A2(n16843), .B1(n19398), .B2(n764), .ZN(
        n16847) );
  NAND3_X1 U27762 ( .A1(n18025), .A2(n18024), .A3(n16844), .ZN(n19386) );
  OAI21_X1 U27763 ( .B1(n17568), .B2(n19388), .A(n19395), .ZN(n16846) );
  NAND2_X1 U27764 ( .A1(n18024), .A2(n17484), .ZN(n18011) );
  NOR2_X1 U27765 ( .A1(n18022), .A2(n18023), .ZN(n18017) );
  INV_X1 U27766 ( .A(n18017), .ZN(n17582) );
  NAND3_X1 U27767 ( .A1(n18012), .A2(n18013), .A3(n18024), .ZN(n16845) );
  NOR2_X1 U27768 ( .A1(n23480), .A2(n2130), .ZN(n21969) );
  AND3_X1 U27769 ( .A1(n23480), .A2(n23477), .A3(n23481), .ZN(n16848) );
  NAND2_X1 U27770 ( .A1(n23485), .A2(n16848), .ZN(n16852) );
  NOR2_X1 U27771 ( .A1(n23483), .A2(n21981), .ZN(n21339) );
  NAND3_X1 U27772 ( .A1(n23489), .A2(n23488), .A3(n23480), .ZN(n16851) );
  NAND2_X1 U27773 ( .A1(n21970), .A2(n23480), .ZN(n16850) );
  XNOR2_X1 U27774 ( .A(n28126), .B(n22762), .ZN(n26125) );
  INV_X1 U27775 ( .A(n26125), .ZN(n16855) );
  XNOR2_X1 U27776 ( .A(n16855), .B(n16856), .ZN(n17426) );
  NAND3_X1 U27777 ( .A1(n20175), .A2(n6903), .A3(n21528), .ZN(n16857) );
  AOI21_X1 U27778 ( .B1(n16859), .B2(n21520), .A(n20609), .ZN(n16862) );
  NAND3_X1 U27779 ( .A1(n52210), .A2(n51049), .A3(n18898), .ZN(n16858) );
  MUX2_X1 U27780 ( .A(n16859), .B(n20612), .S(n6903), .Z(n16860) );
  AND2_X1 U27781 ( .A1(n51050), .A2(n20188), .ZN(n21515) );
  AOI22_X1 U27782 ( .A1(n16862), .A2(n16861), .B1(n16860), .B2(n21515), .ZN(
        n16871) );
  NAND2_X1 U27783 ( .A1(n21525), .A2(n20188), .ZN(n16864) );
  OAI22_X1 U27784 ( .A1(n16865), .A2(n16864), .B1(n18898), .B2(n16863), .ZN(
        n16869) );
  INV_X1 U27785 ( .A(n20608), .ZN(n18894) );
  INV_X1 U27786 ( .A(n21520), .ZN(n20178) );
  NAND2_X1 U27787 ( .A1(n18903), .A2(n21530), .ZN(n16866) );
  NAND2_X1 U27788 ( .A1(n16125), .A2(n6903), .ZN(n18896) );
  AOI21_X1 U27789 ( .B1(n16867), .B2(n16866), .A(n18896), .ZN(n16868) );
  NOR2_X1 U27790 ( .A1(n16869), .A2(n16868), .ZN(n16870) );
  AND2_X1 U27791 ( .A1(n20232), .A2(n498), .ZN(n20671) );
  OAI21_X1 U27792 ( .B1(n20678), .B2(n20232), .A(n18102), .ZN(n16874) );
  OAI21_X1 U27794 ( .B1(n20678), .B2(n18873), .A(n20683), .ZN(n16875) );
  NAND2_X1 U27795 ( .A1(n16875), .A2(n20232), .ZN(n16878) );
  NAND2_X1 U27796 ( .A1(n20675), .A2(n18863), .ZN(n16877) );
  OAI21_X1 U27797 ( .B1(n20682), .B2(n20677), .A(n51090), .ZN(n18100) );
  AND2_X1 U27799 ( .A1(n19894), .A2(n19636), .ZN(n19890) );
  NAND4_X1 U27800 ( .A1(n18936), .A2(n19890), .A3(n19663), .A4(n51127), .ZN(
        n16879) );
  XNOR2_X1 U27801 ( .A(n6043), .B(n19662), .ZN(n16880) );
  AND2_X1 U27802 ( .A1(n19658), .A2(n19892), .ZN(n19664) );
  OAI211_X1 U27803 ( .C1(n19664), .C2(n18942), .A(n19893), .B(n16881), .ZN(
        n16883) );
  OAI21_X1 U27804 ( .B1(n52186), .B2(n20270), .A(n20266), .ZN(n16884) );
  AOI21_X1 U27805 ( .B1(n16885), .B2(n3344), .A(n16884), .ZN(n16888) );
  OAI21_X1 U27806 ( .B1(n52186), .B2(n16886), .A(n20272), .ZN(n16887) );
  OAI21_X1 U27807 ( .B1(n16888), .B2(n16887), .A(n20659), .ZN(n16895) );
  NOR2_X1 U27808 ( .A1(n18846), .A2(n3370), .ZN(n16889) );
  NOR2_X1 U27809 ( .A1(n18846), .A2(n21663), .ZN(n16890) );
  OAI211_X1 U27810 ( .C1(n21653), .C2(n16892), .A(n21654), .B(n20660), .ZN(
        n16893) );
  INV_X1 U27811 ( .A(n24287), .ZN(n24295) );
  XNOR2_X1 U27812 ( .A(n16897), .B(n16896), .ZN(n16898) );
  XNOR2_X1 U27813 ( .A(n25325), .B(n16899), .ZN(n26204) );
  XNOR2_X1 U27814 ( .A(n26204), .B(n16900), .ZN(n37476) );
  XNOR2_X1 U27815 ( .A(n4641), .B(n4295), .ZN(n16901) );
  XNOR2_X1 U27816 ( .A(n16901), .B(n49429), .ZN(n16902) );
  XNOR2_X1 U27817 ( .A(n19768), .B(n16902), .ZN(n33719) );
  XNOR2_X1 U27818 ( .A(n37476), .B(n33719), .ZN(n16903) );
  XNOR2_X1 U27819 ( .A(n17364), .B(n16903), .ZN(n16905) );
  XNOR2_X1 U27820 ( .A(n16905), .B(n16904), .ZN(n16906) );
  XNOR2_X1 U27821 ( .A(n16906), .B(n18797), .ZN(n16908) );
  XNOR2_X1 U27822 ( .A(n16908), .B(n16907), .ZN(n16909) );
  XNOR2_X1 U27823 ( .A(n16911), .B(n16910), .ZN(n18633) );
  XNOR2_X1 U27824 ( .A(n52228), .B(n1354), .ZN(n19237) );
  XNOR2_X1 U27825 ( .A(n17798), .B(n19237), .ZN(n16912) );
  XNOR2_X1 U27826 ( .A(n18633), .B(n16912), .ZN(n16929) );
  XNOR2_X1 U27827 ( .A(n16913), .B(n51757), .ZN(n18815) );
  XNOR2_X1 U27828 ( .A(n33221), .B(n4618), .ZN(n16914) );
  XNOR2_X1 U27829 ( .A(n24861), .B(n16914), .ZN(n16915) );
  XNOR2_X1 U27830 ( .A(n16915), .B(n25901), .ZN(n16916) );
  XNOR2_X1 U27831 ( .A(n16916), .B(n25436), .ZN(n34268) );
  XNOR2_X1 U27832 ( .A(n34266), .B(n33374), .ZN(n16917) );
  XNOR2_X1 U27833 ( .A(n34268), .B(n16917), .ZN(n16918) );
  XNOR2_X1 U27834 ( .A(n16919), .B(n16918), .ZN(n16921) );
  XNOR2_X1 U27835 ( .A(n16921), .B(n16920), .ZN(n16922) );
  XNOR2_X1 U27836 ( .A(n18815), .B(n16922), .ZN(n16927) );
  XNOR2_X1 U27837 ( .A(n18431), .B(n16923), .ZN(n16925) );
  XNOR2_X1 U27838 ( .A(n23495), .B(n26604), .ZN(n24384) );
  XNOR2_X1 U27839 ( .A(n24384), .B(n4712), .ZN(n34234) );
  XNOR2_X1 U27840 ( .A(n4667), .B(n4916), .ZN(n34232) );
  XNOR2_X1 U27841 ( .A(n34816), .B(n34232), .ZN(n16930) );
  XNOR2_X1 U27842 ( .A(n34234), .B(n16930), .ZN(n16931) );
  XNOR2_X1 U27843 ( .A(n16931), .B(n33899), .ZN(n16932) );
  XNOR2_X1 U27844 ( .A(n19261), .B(n16932), .ZN(n16934) );
  XNOR2_X1 U27845 ( .A(n16934), .B(n16933), .ZN(n16935) );
  XNOR2_X1 U27846 ( .A(n17831), .B(n51134), .ZN(n18138) );
  XNOR2_X1 U27847 ( .A(n16935), .B(n18138), .ZN(n16936) );
  XNOR2_X1 U27848 ( .A(n16937), .B(n16936), .ZN(n16940) );
  XNOR2_X1 U27849 ( .A(n576), .B(n355), .ZN(n17380) );
  XNOR2_X1 U27850 ( .A(n17380), .B(n18604), .ZN(n16939) );
  XNOR2_X1 U27852 ( .A(n34377), .B(n4471), .ZN(n42712) );
  XNOR2_X1 U27853 ( .A(n35518), .B(n18117), .ZN(n27244) );
  XNOR2_X1 U27854 ( .A(n42712), .B(n27244), .ZN(n32752) );
  XNOR2_X1 U27855 ( .A(n35052), .B(n4827), .ZN(n16941) );
  XNOR2_X1 U27856 ( .A(n16942), .B(n18827), .ZN(n16945) );
  XNOR2_X1 U27857 ( .A(n16943), .B(n18831), .ZN(n16944) );
  XNOR2_X1 U27858 ( .A(n16945), .B(n16944), .ZN(n16947) );
  XNOR2_X1 U27859 ( .A(n16947), .B(n16946), .ZN(n16949) );
  XNOR2_X1 U27860 ( .A(n16949), .B(n16948), .ZN(n16951) );
  XNOR2_X1 U27861 ( .A(n16951), .B(n16950), .ZN(n19648) );
  NAND2_X1 U27862 ( .A1(n19868), .A2(n19648), .ZN(n19873) );
  NOR2_X1 U27863 ( .A1(n19873), .A2(n19649), .ZN(n18253) );
  XNOR2_X1 U27864 ( .A(n16954), .B(n16955), .ZN(n17225) );
  XNOR2_X1 U27865 ( .A(n16957), .B(n16956), .ZN(n16958) );
  XNOR2_X1 U27866 ( .A(n637), .B(n17707), .ZN(n16959) );
  XNOR2_X1 U27867 ( .A(n16960), .B(n16959), .ZN(n16962) );
  XNOR2_X1 U27868 ( .A(n16961), .B(n16962), .ZN(n17761) );
  XNOR2_X1 U27869 ( .A(n42816), .B(n2112), .ZN(n42240) );
  XNOR2_X1 U27870 ( .A(n17764), .B(n42240), .ZN(n16963) );
  XNOR2_X1 U27871 ( .A(n34414), .B(n4312), .ZN(n41828) );
  XNOR2_X1 U27872 ( .A(n36824), .B(n41828), .ZN(n24397) );
  XNOR2_X1 U27873 ( .A(n4940), .B(n4451), .ZN(n16964) );
  XNOR2_X1 U27874 ( .A(n24397), .B(n16964), .ZN(n16965) );
  XNOR2_X1 U27875 ( .A(n19199), .B(n16965), .ZN(n16966) );
  XNOR2_X1 U27876 ( .A(n17758), .B(n16966), .ZN(n16967) );
  XNOR2_X1 U27877 ( .A(n18161), .B(n16967), .ZN(n16968) );
  XNOR2_X1 U27878 ( .A(n17761), .B(n16968), .ZN(n16969) );
  MUX2_X1 U27879 ( .A(n19640), .B(n18253), .S(n374), .Z(n16985) );
  XNOR2_X1 U27880 ( .A(n18394), .B(n16970), .ZN(n16971) );
  XNOR2_X1 U27881 ( .A(n16972), .B(n16971), .ZN(n16984) );
  XNOR2_X1 U27882 ( .A(n17322), .B(n4639), .ZN(n16974) );
  XNOR2_X1 U27883 ( .A(n16974), .B(n16973), .ZN(n16975) );
  XNOR2_X1 U27884 ( .A(n51047), .B(n16975), .ZN(n17156) );
  XNOR2_X1 U27885 ( .A(n18539), .B(n18175), .ZN(n16979) );
  INV_X1 U27886 ( .A(n16976), .ZN(n25957) );
  XNOR2_X1 U27887 ( .A(n25957), .B(n4651), .ZN(n25309) );
  XNOR2_X1 U27888 ( .A(n25309), .B(n25575), .ZN(n37316) );
  XNOR2_X1 U27889 ( .A(n25114), .B(n16977), .ZN(n41562) );
  XNOR2_X1 U27890 ( .A(n4880), .B(n75), .ZN(n17318) );
  XNOR2_X1 U27891 ( .A(n41562), .B(n17318), .ZN(n32806) );
  XNOR2_X1 U27892 ( .A(n37316), .B(n32806), .ZN(n16978) );
  XNOR2_X1 U27893 ( .A(n16979), .B(n16978), .ZN(n16981) );
  XNOR2_X1 U27894 ( .A(n16980), .B(n17212), .ZN(n18176) );
  XNOR2_X1 U27895 ( .A(n16981), .B(n18176), .ZN(n16982) );
  XNOR2_X1 U27896 ( .A(n17156), .B(n16982), .ZN(n16983) );
  XNOR2_X1 U27897 ( .A(n16984), .B(n16983), .ZN(n19869) );
  NAND2_X1 U27898 ( .A1(n16985), .A2(n19865), .ZN(n16992) );
  INV_X1 U27900 ( .A(n19648), .ZN(n19866) );
  NAND2_X1 U27901 ( .A1(n51039), .A2(n19866), .ZN(n19864) );
  NOR2_X1 U27902 ( .A1(n19867), .A2(n19864), .ZN(n18910) );
  NAND2_X1 U27903 ( .A1(n19866), .A2(n374), .ZN(n19642) );
  AOI21_X1 U27904 ( .B1(n18910), .B2(n19650), .A(n18254), .ZN(n16991) );
  INV_X1 U27905 ( .A(n19873), .ZN(n19030) );
  NAND3_X1 U27906 ( .A1(n19031), .A2(n19030), .A3(n19846), .ZN(n16990) );
  OAI21_X1 U27907 ( .B1(n19847), .B2(n19846), .A(n19865), .ZN(n16988) );
  AND2_X1 U27908 ( .A1(n19866), .A2(n19647), .ZN(n19858) );
  NAND2_X1 U27909 ( .A1(n19858), .A2(n19870), .ZN(n16987) );
  NAND4_X1 U27910 ( .A1(n16988), .A2(n19873), .A3(n19871), .A4(n16987), .ZN(
        n16989) );
  NOR2_X1 U27912 ( .A1(n24295), .A2(n52206), .ZN(n20985) );
  NOR2_X1 U27913 ( .A1(n21905), .A2(n23504), .ZN(n24293) );
  INV_X1 U27914 ( .A(n24293), .ZN(n16993) );
  NAND2_X1 U27915 ( .A1(n19679), .A2(n20211), .ZN(n20207) );
  AOI21_X1 U27916 ( .B1(n20207), .B2(n19671), .A(n51006), .ZN(n16996) );
  OAI211_X1 U27917 ( .C1(n16996), .C2(n20217), .A(n4681), .B(n16995), .ZN(
        n16997) );
  NAND3_X1 U27918 ( .A1(n16998), .A2(n19676), .A3(n16997), .ZN(n17004) );
  AOI21_X1 U27919 ( .B1(n19673), .B2(n19679), .A(n20211), .ZN(n16999) );
  AND2_X1 U27920 ( .A1(n19689), .A2(n16999), .ZN(n17002) );
  OAI22_X1 U27921 ( .A1(n51128), .A2(n20216), .B1(n19689), .B2(n20207), .ZN(
        n17001) );
  MUX2_X1 U27922 ( .A(n17002), .B(n17001), .S(n19685), .Z(n17003) );
  NAND2_X1 U27923 ( .A1(n52207), .A2(n23510), .ZN(n17006) );
  INV_X1 U27925 ( .A(n21082), .ZN(n21911) );
  OAI21_X1 U27926 ( .B1(n24291), .B2(n17006), .A(n21911), .ZN(n17008) );
  AOI21_X1 U27927 ( .B1(n24280), .B2(n21902), .A(n24289), .ZN(n17007) );
  NOR2_X1 U27928 ( .A1(n17008), .A2(n17007), .ZN(n17010) );
  INV_X1 U27930 ( .A(n24282), .ZN(n21086) );
  INV_X1 U27931 ( .A(n24291), .ZN(n20981) );
  NAND2_X1 U27932 ( .A1(n20981), .A2(n7519), .ZN(n17009) );
  INV_X1 U27933 ( .A(n24866), .ZN(n23725) );
  INV_X1 U27934 ( .A(n17093), .ZN(n17016) );
  INV_X1 U27935 ( .A(n17094), .ZN(n17015) );
  OAI21_X1 U27936 ( .B1(n19048), .B2(n19056), .A(n20114), .ZN(n17012) );
  NAND2_X1 U27937 ( .A1(n17012), .A2(n19543), .ZN(n17014) );
  NAND3_X1 U27938 ( .A1(n20123), .A2(n51126), .A3(n19544), .ZN(n17013) );
  OAI211_X1 U27939 ( .C1(n17016), .C2(n17015), .A(n17014), .B(n17013), .ZN(
        n17017) );
  NAND2_X1 U27940 ( .A1(n20158), .A2(n20155), .ZN(n17099) );
  OAI21_X1 U27941 ( .B1(n17099), .B2(n5058), .A(n20116), .ZN(n17019) );
  AOI22_X1 U27942 ( .A1(n17019), .A2(n52401), .B1(n19540), .B2(n17018), .ZN(
        n17020) );
  OR2_X1 U27943 ( .A1(n17020), .A2(n20166), .ZN(n17023) );
  AND2_X1 U27944 ( .A1(n20114), .A2(n19056), .ZN(n20110) );
  INV_X1 U27945 ( .A(n19143), .ZN(n20056) );
  NAND2_X1 U27946 ( .A1(n18303), .A2(n20075), .ZN(n17024) );
  NAND2_X1 U27947 ( .A1(n20073), .A2(n17024), .ZN(n17025) );
  AOI22_X1 U27948 ( .A1(n17026), .A2(n19135), .B1(n20056), .B2(n17025), .ZN(
        n17030) );
  AOI22_X1 U27949 ( .A1(n20056), .A2(n17027), .B1(n20075), .B2(n2101), .ZN(
        n17029) );
  NAND2_X1 U27950 ( .A1(n19143), .A2(n4459), .ZN(n17033) );
  NOR2_X1 U27951 ( .A1(n20072), .A2(n20075), .ZN(n20057) );
  NAND3_X1 U27952 ( .A1(n17033), .A2(n20057), .A3(n20060), .ZN(n17028) );
  INV_X1 U27953 ( .A(n19135), .ZN(n18304) );
  NAND2_X1 U27954 ( .A1(n20082), .A2(n20075), .ZN(n17031) );
  AOI21_X1 U27955 ( .B1(n20067), .B2(n20052), .A(n17031), .ZN(n17032) );
  OAI21_X1 U27956 ( .B1(n17033), .B2(n18304), .A(n17032), .ZN(n17034) );
  OAI21_X1 U27957 ( .B1(n17035), .B2(n21237), .A(n21235), .ZN(n17043) );
  OAI21_X1 U27958 ( .B1(n17036), .B2(n19113), .A(n21231), .ZN(n17037) );
  NOR2_X1 U27959 ( .A1(n770), .A2(n19503), .ZN(n17038) );
  AOI22_X1 U27960 ( .A1(n17313), .A2(n17038), .B1(n761), .B2(n19113), .ZN(
        n17042) );
  AND2_X1 U27961 ( .A1(n19510), .A2(n19503), .ZN(n19505) );
  NAND2_X1 U27962 ( .A1(n19505), .A2(n21233), .ZN(n17040) );
  NAND2_X1 U27963 ( .A1(n6226), .A2(n19504), .ZN(n19509) );
  NAND4_X1 U27964 ( .A1(n17040), .A2(n17039), .A3(n19520), .A4(n19509), .ZN(
        n17041) );
  NAND2_X1 U27965 ( .A1(n17046), .A2(n5881), .ZN(n20030) );
  OAI211_X1 U27966 ( .C1(n17047), .C2(n7920), .A(n20030), .B(n20027), .ZN(
        n17048) );
  OAI211_X1 U27967 ( .C1(n17050), .C2(n5881), .A(n17049), .B(n5385), .ZN(
        n17051) );
  AND2_X1 U27968 ( .A1(n23546), .A2(n23360), .ZN(n23364) );
  INV_X1 U27969 ( .A(n23364), .ZN(n23352) );
  OR2_X1 U27970 ( .A1(n17057), .A2(n20094), .ZN(n17503) );
  AND2_X1 U27972 ( .A1(n18316), .A2(n20097), .ZN(n17053) );
  NOR2_X1 U27973 ( .A1(n20085), .A2(n17053), .ZN(n17064) );
  INV_X1 U27974 ( .A(n17056), .ZN(n20096) );
  NAND2_X1 U27975 ( .A1(n20096), .A2(n20088), .ZN(n17506) );
  INV_X1 U27976 ( .A(n17506), .ZN(n17055) );
  OAI21_X1 U27977 ( .B1(n18318), .B2(n17505), .A(n17600), .ZN(n17054) );
  OAI21_X1 U27978 ( .B1(n17055), .B2(n17603), .A(n17054), .ZN(n17063) );
  NOR2_X1 U27979 ( .A1(n17056), .A2(n20088), .ZN(n20103) );
  NOR2_X1 U27980 ( .A1(n17057), .A2(n20104), .ZN(n17058) );
  OAI21_X1 U27981 ( .B1(n20103), .B2(n17058), .A(n20105), .ZN(n17062) );
  INV_X1 U27982 ( .A(n20092), .ZN(n20087) );
  OAI21_X1 U27983 ( .B1(n17504), .B2(n20087), .A(n20101), .ZN(n17060) );
  AND2_X1 U27984 ( .A1(n8624), .A2(n20095), .ZN(n20090) );
  INV_X1 U27985 ( .A(n18318), .ZN(n17599) );
  NAND3_X1 U27986 ( .A1(n17060), .A2(n20090), .A3(n17599), .ZN(n17061) );
  INV_X1 U27987 ( .A(n19061), .ZN(n17066) );
  INV_X1 U27988 ( .A(n19071), .ZN(n20148) );
  OAI22_X1 U27989 ( .A1(n17067), .A2(n20147), .B1(n20148), .B2(n18344), .ZN(
        n17068) );
  NAND2_X1 U27990 ( .A1(n17068), .A2(n18345), .ZN(n17073) );
  INV_X1 U27991 ( .A(n18354), .ZN(n17070) );
  INV_X1 U27993 ( .A(n51675), .ZN(n20721) );
  NOR2_X1 U27994 ( .A1(n21155), .A2(n23563), .ZN(n20726) );
  NAND2_X1 U27995 ( .A1(n22275), .A2(n20726), .ZN(n17075) );
  NAND2_X1 U27996 ( .A1(n51677), .A2(n23360), .ZN(n21154) );
  NAND2_X1 U27997 ( .A1(n23568), .A2(n23546), .ZN(n23350) );
  AND2_X1 U27999 ( .A1(n17081), .A2(n19477), .ZN(n21243) );
  AOI21_X1 U28000 ( .B1(n17076), .B2(n21243), .A(n51132), .ZN(n17077) );
  AOI22_X1 U28002 ( .A1(n19099), .A2(n21243), .B1(n17079), .B2(n21254), .ZN(
        n17080) );
  NAND2_X1 U28003 ( .A1(n18969), .A2(n17083), .ZN(n19102) );
  NAND3_X1 U28004 ( .A1(n19475), .A2(n19087), .A3(n17081), .ZN(n19094) );
  NAND2_X1 U28005 ( .A1(n21245), .A2(n19477), .ZN(n17082) );
  AOI21_X1 U28008 ( .B1(n3335), .B2(n18963), .A(n17084), .ZN(n17085) );
  MUX2_X1 U28010 ( .A(n17086), .B(n17085), .S(n18966), .Z(n17087) );
  INV_X1 U28011 ( .A(n17087), .ZN(n17088) );
  MUX2_X1 U28012 ( .A(n19055), .B(n20116), .S(n20124), .Z(n17097) );
  NOR2_X1 U28013 ( .A1(n17090), .A2(n5058), .ZN(n17092) );
  NOR2_X1 U28014 ( .A1(n4081), .A2(n19534), .ZN(n17091) );
  AOI22_X1 U28015 ( .A1(n17092), .A2(n20125), .B1(n19540), .B2(n17091), .ZN(
        n17096) );
  NAND3_X1 U28016 ( .A1(n19540), .A2(n20125), .A3(n19048), .ZN(n20112) );
  INV_X1 U28017 ( .A(n20166), .ZN(n19045) );
  NAND2_X1 U28018 ( .A1(n16490), .A2(n20157), .ZN(n17098) );
  OR2_X1 U28019 ( .A1(n17099), .A2(n17098), .ZN(n19052) );
  INV_X1 U28021 ( .A(n24313), .ZN(n17103) );
  XNOR2_X1 U28022 ( .A(n17103), .B(n23943), .ZN(n33696) );
  XNOR2_X1 U28023 ( .A(n25094), .B(n35815), .ZN(n34590) );
  XOR2_X1 U28024 ( .A(n4720), .B(n4537), .Z(n17104) );
  XNOR2_X1 U28025 ( .A(n1354), .B(n46552), .ZN(n44885) );
  XNOR2_X1 U28026 ( .A(n17104), .B(n44885), .ZN(n17105) );
  XNOR2_X1 U28027 ( .A(n34590), .B(n17105), .ZN(n17106) );
  XNOR2_X1 U28028 ( .A(n33696), .B(n17106), .ZN(n17107) );
  XNOR2_X1 U28029 ( .A(n17108), .B(n17107), .ZN(n17109) );
  XNOR2_X1 U28030 ( .A(n18196), .B(n17109), .ZN(n17112) );
  XNOR2_X1 U28031 ( .A(n51459), .B(n17110), .ZN(n17111) );
  INV_X1 U28032 ( .A(n17115), .ZN(n17132) );
  XNOR2_X1 U28033 ( .A(n17116), .B(n19244), .ZN(n17120) );
  XNOR2_X1 U28034 ( .A(n17118), .B(n17117), .ZN(n17119) );
  XNOR2_X1 U28035 ( .A(n17938), .B(n17119), .ZN(n17369) );
  XNOR2_X1 U28036 ( .A(n17120), .B(n17369), .ZN(n17130) );
  XNOR2_X1 U28037 ( .A(n17121), .B(n4641), .ZN(n41597) );
  XNOR2_X1 U28038 ( .A(n25078), .B(n24057), .ZN(n25207) );
  XNOR2_X1 U28039 ( .A(n41597), .B(n25207), .ZN(n35640) );
  XNOR2_X1 U28040 ( .A(n37288), .B(n4076), .ZN(n17122) );
  XNOR2_X1 U28041 ( .A(n17122), .B(n25147), .ZN(n26205) );
  XNOR2_X1 U28042 ( .A(n4589), .B(n4568), .ZN(n17123) );
  XNOR2_X1 U28043 ( .A(n26205), .B(n17123), .ZN(n35220) );
  XNOR2_X1 U28044 ( .A(n35640), .B(n35220), .ZN(n17124) );
  XNOR2_X1 U28045 ( .A(n17646), .B(n17124), .ZN(n17126) );
  XNOR2_X1 U28046 ( .A(n17126), .B(n17125), .ZN(n17128) );
  XNOR2_X1 U28047 ( .A(n17128), .B(n17127), .ZN(n17129) );
  XNOR2_X1 U28048 ( .A(n17130), .B(n17129), .ZN(n17131) );
  XNOR2_X1 U28049 ( .A(n33635), .B(n4637), .ZN(n37008) );
  XNOR2_X1 U28050 ( .A(n17763), .B(n37008), .ZN(n17133) );
  XNOR2_X1 U28051 ( .A(n17758), .B(n18407), .ZN(n17140) );
  XNOR2_X1 U28052 ( .A(n28058), .B(n25470), .ZN(n33934) );
  XNOR2_X1 U28053 ( .A(n4937), .B(n4157), .ZN(n34773) );
  XNOR2_X1 U28054 ( .A(n41155), .B(n34773), .ZN(n17135) );
  XNOR2_X1 U28055 ( .A(n33931), .B(n17135), .ZN(n17136) );
  XNOR2_X1 U28056 ( .A(n33934), .B(n17136), .ZN(n17137) );
  XNOR2_X1 U28057 ( .A(n17138), .B(n17137), .ZN(n17139) );
  XNOR2_X1 U28058 ( .A(n17140), .B(n17139), .ZN(n17141) );
  XNOR2_X1 U28059 ( .A(n17142), .B(n17141), .ZN(n17143) );
  XNOR2_X1 U28060 ( .A(n17146), .B(n17145), .ZN(n17714) );
  XNOR2_X1 U28061 ( .A(n18540), .B(n18773), .ZN(n17154) );
  XNOR2_X1 U28062 ( .A(n24894), .B(n4659), .ZN(n24830) );
  XNOR2_X1 U28063 ( .A(n18172), .B(n4536), .ZN(n17147) );
  XNOR2_X1 U28064 ( .A(n24830), .B(n17147), .ZN(n36876) );
  XNOR2_X1 U28065 ( .A(n17148), .B(n36876), .ZN(n17151) );
  XNOR2_X1 U28066 ( .A(n17149), .B(n75), .ZN(n32627) );
  XNOR2_X1 U28067 ( .A(n32627), .B(n4578), .ZN(n17150) );
  XNOR2_X1 U28068 ( .A(n17151), .B(n17150), .ZN(n17152) );
  XNOR2_X1 U28069 ( .A(n17321), .B(n17152), .ZN(n17153) );
  XNOR2_X1 U28070 ( .A(n17154), .B(n17153), .ZN(n17155) );
  XNOR2_X1 U28071 ( .A(n17714), .B(n17155), .ZN(n17157) );
  INV_X1 U28072 ( .A(n17158), .ZN(n17160) );
  XNOR2_X1 U28073 ( .A(n17902), .B(n18175), .ZN(n17159) );
  AOI21_X1 U28074 ( .B1(n19702), .B2(n21178), .A(n19703), .ZN(n17197) );
  XNOR2_X1 U28075 ( .A(n42461), .B(n2231), .ZN(n17162) );
  INV_X1 U28076 ( .A(n45350), .ZN(n18461) );
  XNOR2_X1 U28077 ( .A(n17162), .B(n18461), .ZN(n26443) );
  XNOR2_X1 U28078 ( .A(n44493), .B(n4754), .ZN(n23884) );
  XNOR2_X1 U28079 ( .A(n26443), .B(n23884), .ZN(n34536) );
  XNOR2_X1 U28080 ( .A(n2203), .B(n4429), .ZN(n17163) );
  XNOR2_X1 U28081 ( .A(n41367), .B(n17163), .ZN(n23886) );
  XNOR2_X1 U28082 ( .A(n23886), .B(n49790), .ZN(n45085) );
  XNOR2_X1 U28083 ( .A(n45085), .B(n17164), .ZN(n33769) );
  XNOR2_X1 U28084 ( .A(n34536), .B(n33769), .ZN(n17165) );
  XNOR2_X1 U28085 ( .A(n17829), .B(n17165), .ZN(n17166) );
  XNOR2_X1 U28086 ( .A(n18602), .B(n17166), .ZN(n17167) );
  XNOR2_X1 U28087 ( .A(n17168), .B(n17167), .ZN(n17173) );
  XNOR2_X1 U28088 ( .A(n17171), .B(n356), .ZN(n17172) );
  XNOR2_X1 U28089 ( .A(n17173), .B(n17172), .ZN(n17174) );
  XNOR2_X1 U28090 ( .A(n17175), .B(n17174), .ZN(n17176) );
  INV_X1 U28091 ( .A(n21185), .ZN(n19832) );
  XNOR2_X1 U28092 ( .A(n17177), .B(n17731), .ZN(n17179) );
  XNOR2_X1 U28093 ( .A(n17181), .B(n17180), .ZN(n26243) );
  XNOR2_X1 U28094 ( .A(n44483), .B(n4676), .ZN(n26242) );
  XNOR2_X1 U28095 ( .A(n26242), .B(n1341), .ZN(n17390) );
  XNOR2_X1 U28096 ( .A(n26243), .B(n17390), .ZN(n36836) );
  XNOR2_X1 U28097 ( .A(n4486), .B(n4317), .ZN(n18118) );
  XNOR2_X1 U28098 ( .A(n18118), .B(n17182), .ZN(n43766) );
  XNOR2_X1 U28099 ( .A(n43105), .B(n4628), .ZN(n17183) );
  XNOR2_X1 U28100 ( .A(n43766), .B(n17183), .ZN(n32495) );
  XNOR2_X1 U28101 ( .A(n36836), .B(n32495), .ZN(n17184) );
  XNOR2_X1 U28102 ( .A(n17389), .B(n17184), .ZN(n17185) );
  XNOR2_X1 U28103 ( .A(n17186), .B(n17185), .ZN(n17187) );
  XNOR2_X1 U28104 ( .A(n18701), .B(n18123), .ZN(n17191) );
  XNOR2_X1 U28105 ( .A(n18488), .B(n17191), .ZN(n17192) );
  INV_X1 U28106 ( .A(n19839), .ZN(n21188) );
  AND2_X1 U28107 ( .A1(n21186), .A2(n17201), .ZN(n19840) );
  OAI21_X1 U28108 ( .B1(n19702), .B2(n17194), .A(n19840), .ZN(n17196) );
  INV_X1 U28109 ( .A(n19834), .ZN(n19828) );
  MUX2_X1 U28110 ( .A(n17197), .B(n17196), .S(n18973), .Z(n17207) );
  NAND2_X1 U28111 ( .A1(n21186), .A2(n21173), .ZN(n19699) );
  AND2_X1 U28112 ( .A1(n21173), .A2(n21188), .ZN(n18975) );
  AND3_X1 U28113 ( .A1(n19699), .A2(n18975), .A3(n19832), .ZN(n17200) );
  AND2_X1 U28114 ( .A1(n21188), .A2(n19826), .ZN(n21175) );
  MUX2_X1 U28115 ( .A(n21175), .B(n51434), .S(n19828), .Z(n17199) );
  INV_X1 U28116 ( .A(n19837), .ZN(n19705) );
  NOR2_X1 U28117 ( .A1(n19705), .A2(n21185), .ZN(n17198) );
  INV_X1 U28118 ( .A(n21174), .ZN(n17202) );
  NAND3_X1 U28119 ( .A1(n17202), .A2(n21171), .A3(n17201), .ZN(n17206) );
  NAND3_X1 U28120 ( .A1(n21178), .A2(n21181), .A3(n19826), .ZN(n19829) );
  INV_X1 U28121 ( .A(n19829), .ZN(n17203) );
  NAND2_X1 U28122 ( .A1(n17204), .A2(n21185), .ZN(n17205) );
  XNOR2_X1 U28123 ( .A(n18773), .B(n17901), .ZN(n17209) );
  XNOR2_X1 U28124 ( .A(n17209), .B(n17208), .ZN(n17210) );
  XNOR2_X1 U28125 ( .A(n17211), .B(n17210), .ZN(n17784) );
  XNOR2_X1 U28126 ( .A(n51373), .B(n17213), .ZN(n17220) );
  XNOR2_X1 U28127 ( .A(n3383), .B(n4542), .ZN(n36994) );
  XNOR2_X1 U28128 ( .A(n36994), .B(n4705), .ZN(n17214) );
  XNOR2_X1 U28129 ( .A(n17214), .B(n26297), .ZN(n25959) );
  XNOR2_X1 U28130 ( .A(n25959), .B(n25114), .ZN(n33164) );
  XNOR2_X1 U28131 ( .A(n25575), .B(n42769), .ZN(n17215) );
  XNOR2_X1 U28132 ( .A(n33164), .B(n17215), .ZN(n17216) );
  XNOR2_X1 U28133 ( .A(n25957), .B(n4659), .ZN(n25255) );
  XNOR2_X1 U28134 ( .A(n17216), .B(n25255), .ZN(n17217) );
  XNOR2_X1 U28135 ( .A(n17218), .B(n17217), .ZN(n17219) );
  XNOR2_X1 U28136 ( .A(n17220), .B(n17219), .ZN(n17222) );
  XNOR2_X1 U28137 ( .A(n17222), .B(n17221), .ZN(n17223) );
  XNOR2_X1 U28138 ( .A(n17784), .B(n17223), .ZN(n17224) );
  INV_X1 U28139 ( .A(n36824), .ZN(n17228) );
  XNOR2_X1 U28140 ( .A(n43019), .B(n4564), .ZN(n17227) );
  XNOR2_X1 U28141 ( .A(n17228), .B(n17227), .ZN(n33795) );
  XNOR2_X1 U28142 ( .A(n4793), .B(n4896), .ZN(n41496) );
  XNOR2_X1 U28143 ( .A(n41496), .B(n4343), .ZN(n17229) );
  XNOR2_X1 U28144 ( .A(n4940), .B(n4501), .ZN(n27203) );
  XNOR2_X1 U28145 ( .A(n17229), .B(n27203), .ZN(n43370) );
  XNOR2_X1 U28146 ( .A(n44934), .B(n4213), .ZN(n34072) );
  XNOR2_X1 U28147 ( .A(n43370), .B(n34072), .ZN(n17230) );
  XNOR2_X1 U28148 ( .A(n33795), .B(n17230), .ZN(n17231) );
  XNOR2_X1 U28149 ( .A(n17232), .B(n17231), .ZN(n17233) );
  XNOR2_X1 U28150 ( .A(n51437), .B(n17233), .ZN(n17235) );
  XNOR2_X1 U28151 ( .A(n17879), .B(n17234), .ZN(n17756) );
  XNOR2_X1 U28152 ( .A(n17756), .B(n17235), .ZN(n17237) );
  XNOR2_X1 U28153 ( .A(n18408), .B(n2135), .ZN(n18507) );
  XNOR2_X1 U28154 ( .A(n17237), .B(n17236), .ZN(n17238) );
  XNOR2_X1 U28155 ( .A(n17240), .B(n17239), .ZN(n17252) );
  XNOR2_X1 U28156 ( .A(n17646), .B(n17812), .ZN(n17248) );
  BUF_X1 U28157 ( .A(Key[50]), .Z(n42668) );
  XNOR2_X1 U28158 ( .A(n42668), .B(n3014), .ZN(n24820) );
  XNOR2_X1 U28159 ( .A(n35796), .B(n24820), .ZN(n17241) );
  XNOR2_X1 U28160 ( .A(n35532), .B(n17241), .ZN(n17242) );
  XNOR2_X1 U28161 ( .A(n17242), .B(n37082), .ZN(n17244) );
  INV_X1 U28162 ( .A(n4589), .ZN(n48122) );
  XNOR2_X1 U28163 ( .A(n37288), .B(n48122), .ZN(n37473) );
  XNOR2_X1 U28164 ( .A(n17243), .B(n37473), .ZN(n35795) );
  XNOR2_X1 U28165 ( .A(n17244), .B(n35795), .ZN(n17245) );
  XNOR2_X1 U28166 ( .A(n17246), .B(n17245), .ZN(n17247) );
  XNOR2_X1 U28167 ( .A(n17248), .B(n17247), .ZN(n17251) );
  XNOR2_X1 U28168 ( .A(n17938), .B(n17803), .ZN(n17249) );
  XNOR2_X1 U28170 ( .A(n34266), .B(n18191), .ZN(n28283) );
  XNOR2_X1 U28171 ( .A(n28283), .B(n4537), .ZN(n34451) );
  XNOR2_X1 U28172 ( .A(n17254), .B(n32856), .ZN(n33508) );
  XNOR2_X1 U28173 ( .A(n4636), .B(n4720), .ZN(n17255) );
  XNOR2_X1 U28174 ( .A(n33508), .B(n17255), .ZN(n17256) );
  XNOR2_X1 U28175 ( .A(n34451), .B(n17256), .ZN(n17257) );
  INV_X1 U28176 ( .A(n17258), .ZN(n17677) );
  XNOR2_X1 U28177 ( .A(n17259), .B(n17677), .ZN(n17260) );
  XNOR2_X1 U28178 ( .A(n51133), .B(n17260), .ZN(n17263) );
  INV_X1 U28179 ( .A(n17261), .ZN(n17262) );
  XNOR2_X1 U28180 ( .A(n17263), .B(n17262), .ZN(n17271) );
  XNOR2_X1 U28181 ( .A(n18616), .B(n51135), .ZN(n17918) );
  XNOR2_X1 U28182 ( .A(n17264), .B(n18447), .ZN(n17266) );
  XNOR2_X1 U28183 ( .A(n17266), .B(n17265), .ZN(n17267) );
  XNOR2_X1 U28184 ( .A(n17918), .B(n17267), .ZN(n17269) );
  XNOR2_X1 U28185 ( .A(n17269), .B(n17268), .ZN(n17270) );
  NAND3_X1 U28186 ( .A1(n2182), .A2(n21276), .A3(n19776), .ZN(n19020) );
  XNOR2_X1 U28187 ( .A(n18123), .B(n566), .ZN(n17277) );
  XNOR2_X1 U28188 ( .A(n34377), .B(n26244), .ZN(n18570) );
  XNOR2_X1 U28189 ( .A(n26586), .B(n4317), .ZN(n22454) );
  XNOR2_X1 U28190 ( .A(n18570), .B(n22454), .ZN(n33072) );
  XNOR2_X1 U28191 ( .A(n44483), .B(n4518), .ZN(n28087) );
  XNOR2_X1 U28192 ( .A(n28087), .B(n1341), .ZN(n41949) );
  XNOR2_X1 U28193 ( .A(n41949), .B(n4275), .ZN(n17272) );
  XNOR2_X1 U28194 ( .A(n33072), .B(n17272), .ZN(n17273) );
  XNOR2_X1 U28195 ( .A(n18483), .B(n17273), .ZN(n17274) );
  XNOR2_X1 U28196 ( .A(n17275), .B(n17274), .ZN(n17276) );
  XNOR2_X1 U28197 ( .A(n17277), .B(n17276), .ZN(n17279) );
  XNOR2_X1 U28198 ( .A(n17279), .B(n17278), .ZN(n17286) );
  XNOR2_X1 U28199 ( .A(n17280), .B(n5016), .ZN(n17282) );
  XNOR2_X1 U28200 ( .A(n17282), .B(n17281), .ZN(n17726) );
  XNOR2_X1 U28201 ( .A(n17726), .B(n18485), .ZN(n17283) );
  XNOR2_X1 U28202 ( .A(n17284), .B(n17283), .ZN(n17285) );
  INV_X1 U28203 ( .A(n19452), .ZN(n19118) );
  XNOR2_X1 U28204 ( .A(n17288), .B(n51417), .ZN(n17290) );
  XNOR2_X1 U28205 ( .A(n17290), .B(n18704), .ZN(n17291) );
  XNOR2_X1 U28206 ( .A(n17291), .B(n18605), .ZN(n17837) );
  XNOR2_X1 U28207 ( .A(n18602), .B(n17292), .ZN(n18142) );
  XNOR2_X1 U28208 ( .A(n18738), .B(n33490), .ZN(n18600) );
  INV_X1 U28209 ( .A(n18600), .ZN(n17293) );
  XNOR2_X1 U28210 ( .A(n17381), .B(n17293), .ZN(n17294) );
  XNOR2_X1 U28211 ( .A(n18142), .B(n17294), .ZN(n17302) );
  XNOR2_X1 U28212 ( .A(n17691), .B(n17973), .ZN(n17299) );
  XNOR2_X1 U28213 ( .A(n4836), .B(n45736), .ZN(n26603) );
  XNOR2_X1 U28214 ( .A(n25616), .B(n26603), .ZN(n17295) );
  XNOR2_X1 U28215 ( .A(n28232), .B(n17295), .ZN(n34494) );
  XNOR2_X1 U28216 ( .A(n28071), .B(n4429), .ZN(n33495) );
  XNOR2_X1 U28217 ( .A(n34494), .B(n33495), .ZN(n17296) );
  XNOR2_X1 U28218 ( .A(n17297), .B(n17296), .ZN(n17298) );
  XNOR2_X1 U28219 ( .A(n17299), .B(n17298), .ZN(n17300) );
  XNOR2_X1 U28220 ( .A(n17300), .B(n17378), .ZN(n17301) );
  XNOR2_X1 U28221 ( .A(n17302), .B(n17301), .ZN(n17303) );
  XNOR2_X1 U28222 ( .A(n17837), .B(n17303), .ZN(n19019) );
  NOR2_X1 U28223 ( .A1(n19122), .A2(n51013), .ZN(n17304) );
  INV_X1 U28224 ( .A(n19459), .ZN(n19779) );
  AOI22_X1 U28225 ( .A1(n17304), .A2(n19779), .B1(n19775), .B2(n19023), .ZN(
        n17307) );
  INV_X1 U28226 ( .A(n19466), .ZN(n19782) );
  OAI21_X1 U28227 ( .B1(n19122), .B2(n2182), .A(n19776), .ZN(n17305) );
  NAND2_X1 U28228 ( .A1(n17305), .A2(n51013), .ZN(n17306) );
  AND2_X1 U28229 ( .A1(n24207), .A2(n22639), .ZN(n23598) );
  NOR2_X1 U28230 ( .A1(n17309), .A2(n21234), .ZN(n17413) );
  INV_X1 U28231 ( .A(n19508), .ZN(n17310) );
  NOR2_X1 U28232 ( .A1(n17311), .A2(n5177), .ZN(n19114) );
  OAI211_X1 U28233 ( .C1(n21239), .C2(n19518), .A(n17416), .B(n17415), .ZN(
        n17312) );
  INV_X1 U28234 ( .A(n17312), .ZN(n17411) );
  INV_X1 U28235 ( .A(n21235), .ZN(n19108) );
  AOI21_X1 U28236 ( .B1(n17314), .B2(n19108), .A(n19510), .ZN(n17315) );
  INV_X1 U28237 ( .A(n17417), .ZN(n17410) );
  XNOR2_X1 U28238 ( .A(n28412), .B(n4035), .ZN(n21090) );
  XNOR2_X1 U28239 ( .A(n21090), .B(n23711), .ZN(n24521) );
  XNOR2_X1 U28240 ( .A(n17318), .B(n17317), .ZN(n25793) );
  XNOR2_X1 U28241 ( .A(n24227), .B(n25793), .ZN(n27230) );
  XNOR2_X1 U28242 ( .A(n24521), .B(n27230), .ZN(n36756) );
  XNOR2_X1 U28243 ( .A(n36756), .B(n43054), .ZN(n17319) );
  XNOR2_X1 U28244 ( .A(n17320), .B(n17319), .ZN(n17324) );
  XNOR2_X1 U28245 ( .A(n17322), .B(n17321), .ZN(n17323) );
  XNOR2_X1 U28246 ( .A(n17324), .B(n17323), .ZN(n17325) );
  XNOR2_X1 U28247 ( .A(n17326), .B(n17325), .ZN(n17329) );
  INV_X1 U28248 ( .A(n17327), .ZN(n17328) );
  XNOR2_X1 U28249 ( .A(n17329), .B(n17328), .ZN(n17401) );
  INV_X1 U28250 ( .A(n17401), .ZN(n19820) );
  XNOR2_X1 U28251 ( .A(n17234), .B(n17758), .ZN(n17330) );
  XNOR2_X1 U28252 ( .A(n17331), .B(n17330), .ZN(n17333) );
  XNOR2_X1 U28253 ( .A(n17333), .B(n17332), .ZN(n17336) );
  INV_X1 U28254 ( .A(n17334), .ZN(n17335) );
  XNOR2_X1 U28255 ( .A(n34080), .B(n4316), .ZN(n17337) );
  XNOR2_X1 U28256 ( .A(n37008), .B(n17337), .ZN(n17338) );
  XNOR2_X1 U28257 ( .A(n41155), .B(n4638), .ZN(n41497) );
  XNOR2_X1 U28258 ( .A(n17338), .B(n41497), .ZN(n17339) );
  XNOR2_X1 U28259 ( .A(n33297), .B(n42240), .ZN(n32553) );
  XNOR2_X1 U28260 ( .A(n17339), .B(n32553), .ZN(n17340) );
  XNOR2_X1 U28261 ( .A(n18153), .B(n17340), .ZN(n17341) );
  XNOR2_X1 U28262 ( .A(n18407), .B(n17341), .ZN(n17342) );
  XNOR2_X1 U28263 ( .A(n17343), .B(n17342), .ZN(n17345) );
  XNOR2_X1 U28264 ( .A(n17344), .B(n17345), .ZN(n17346) );
  XNOR2_X1 U28265 ( .A(n18443), .B(n18193), .ZN(n17347) );
  XNOR2_X1 U28266 ( .A(n17348), .B(n17347), .ZN(n17350) );
  XNOR2_X1 U28267 ( .A(n17350), .B(n17349), .ZN(n17352) );
  XNOR2_X1 U28268 ( .A(n17351), .B(n17352), .ZN(n17359) );
  XNOR2_X1 U28269 ( .A(n43564), .B(n24626), .ZN(n34333) );
  XNOR2_X1 U28270 ( .A(n49937), .B(n1354), .ZN(n41660) );
  XNOR2_X1 U28271 ( .A(n33611), .B(n41660), .ZN(n17353) );
  XNOR2_X1 U28272 ( .A(n34333), .B(n17353), .ZN(n17354) );
  XNOR2_X1 U28273 ( .A(n18616), .B(n17354), .ZN(n17355) );
  XNOR2_X1 U28274 ( .A(n51133), .B(n17355), .ZN(n17357) );
  XNOR2_X1 U28275 ( .A(n17356), .B(n17357), .ZN(n17358) );
  XNOR2_X1 U28276 ( .A(n17358), .B(n17359), .ZN(n17406) );
  INV_X1 U28277 ( .A(n17406), .ZN(n19725) );
  XNOR2_X1 U28278 ( .A(n48597), .B(n4076), .ZN(n18206) );
  XNOR2_X1 U28279 ( .A(n17360), .B(n18206), .ZN(n27453) );
  XNOR2_X1 U28280 ( .A(n4817), .B(n3276), .ZN(n43560) );
  XNOR2_X1 U28281 ( .A(n27453), .B(n43560), .ZN(n35342) );
  XNOR2_X1 U28282 ( .A(n24057), .B(n26506), .ZN(n35539) );
  XNOR2_X1 U28283 ( .A(n35539), .B(n43691), .ZN(n17361) );
  XNOR2_X1 U28284 ( .A(n35342), .B(n17361), .ZN(n17362) );
  XNOR2_X1 U28285 ( .A(n17812), .B(n17362), .ZN(n17363) );
  XNOR2_X1 U28286 ( .A(n17364), .B(n18795), .ZN(n17366) );
  XNOR2_X1 U28287 ( .A(n17366), .B(n17365), .ZN(n18646) );
  XNOR2_X1 U28288 ( .A(n17367), .B(n18646), .ZN(n17371) );
  XNOR2_X1 U28289 ( .A(n17368), .B(n18208), .ZN(n18802) );
  XNOR2_X1 U28290 ( .A(n18802), .B(n17369), .ZN(n17370) );
  XNOR2_X1 U28291 ( .A(n17371), .B(n17370), .ZN(n17373) );
  INV_X1 U28292 ( .A(n23888), .ZN(n17374) );
  XNOR2_X1 U28293 ( .A(n24748), .B(n17374), .ZN(n41403) );
  XNOR2_X1 U28294 ( .A(n24384), .B(n4838), .ZN(n34397) );
  XNOR2_X1 U28295 ( .A(n34397), .B(n2231), .ZN(n17375) );
  XNOR2_X1 U28296 ( .A(n41403), .B(n17375), .ZN(n17376) );
  XNOR2_X1 U28297 ( .A(n18466), .B(n17376), .ZN(n17377) );
  XNOR2_X1 U28298 ( .A(n17378), .B(n17377), .ZN(n17379) );
  XNOR2_X1 U28299 ( .A(n17380), .B(n17379), .ZN(n17383) );
  XNOR2_X1 U28300 ( .A(n17382), .B(n17381), .ZN(n18743) );
  XNOR2_X1 U28301 ( .A(n17383), .B(n18743), .ZN(n17388) );
  XNOR2_X1 U28302 ( .A(n41367), .B(n2203), .ZN(n33567) );
  XNOR2_X1 U28303 ( .A(n17384), .B(n18739), .ZN(n18141) );
  XNOR2_X1 U28304 ( .A(n18141), .B(n17385), .ZN(n17386) );
  XNOR2_X1 U28305 ( .A(n17976), .B(n17386), .ZN(n17387) );
  XNOR2_X1 U28307 ( .A(n18475), .B(n17389), .ZN(n17393) );
  XNOR2_X1 U28308 ( .A(n17390), .B(n25521), .ZN(n36665) );
  XNOR2_X1 U28309 ( .A(n4585), .B(n4486), .ZN(n31431) );
  XNOR2_X1 U28310 ( .A(n36665), .B(n31431), .ZN(n17391) );
  XNOR2_X1 U28311 ( .A(n18119), .B(n17391), .ZN(n17392) );
  XNOR2_X1 U28312 ( .A(n17393), .B(n17392), .ZN(n17395) );
  XNOR2_X1 U28313 ( .A(n18126), .B(n15619), .ZN(n17394) );
  XNOR2_X1 U28314 ( .A(n17395), .B(n17394), .ZN(n17396) );
  XNOR2_X1 U28315 ( .A(n17397), .B(n17396), .ZN(n17399) );
  XNOR2_X1 U28316 ( .A(n17398), .B(n17399), .ZN(n21198) );
  NAND2_X1 U28317 ( .A1(n2229), .A2(n21213), .ZN(n17400) );
  NAND3_X1 U28318 ( .A1(n19808), .A2(n21208), .A3(n17400), .ZN(n17409) );
  INV_X1 U28319 ( .A(n17405), .ZN(n19007) );
  NAND2_X1 U28320 ( .A1(n17406), .A2(n19007), .ZN(n19813) );
  NAND2_X1 U28321 ( .A1(n21214), .A2(n19823), .ZN(n17402) );
  NAND2_X1 U28322 ( .A1(n17406), .A2(n2229), .ZN(n19733) );
  NAND2_X1 U28323 ( .A1(n19809), .A2(n6078), .ZN(n21211) );
  AOI21_X1 U28324 ( .B1(n17402), .B2(n19733), .A(n21211), .ZN(n17403) );
  NOR2_X1 U28325 ( .A1(n18108), .A2(n17403), .ZN(n17408) );
  NAND2_X1 U28326 ( .A1(n19823), .A2(n19822), .ZN(n21199) );
  INV_X1 U28327 ( .A(n21214), .ZN(n17404) );
  AND2_X1 U28329 ( .A1(n17405), .A2(n17406), .ZN(n19009) );
  NOR2_X1 U28330 ( .A1(n21215), .A2(n19009), .ZN(n18112) );
  AOI21_X1 U28331 ( .B1(n17411), .B2(n17410), .A(n23068), .ZN(n23591) );
  OAI21_X1 U28332 ( .B1(n24206), .B2(n23598), .A(n23591), .ZN(n17424) );
  NAND3_X1 U28333 ( .A1(n17413), .A2(n21233), .A3(n17412), .ZN(n17414) );
  OAI211_X1 U28334 ( .C1(n17418), .C2(n23068), .A(n22638), .B(n23613), .ZN(
        n17422) );
  NOR2_X1 U28335 ( .A1(n17420), .A2(n52155), .ZN(n22643) );
  INV_X1 U28336 ( .A(n22643), .ZN(n17421) );
  NAND4_X1 U28337 ( .A1(n17424), .A2(n17423), .A3(n17422), .A4(n17421), .ZN(
        n25909) );
  XNOR2_X1 U28338 ( .A(n23725), .B(n26053), .ZN(n17425) );
  XNOR2_X1 U28339 ( .A(n17426), .B(n17425), .ZN(n18281) );
  INV_X1 U28340 ( .A(n403), .ZN(n17541) );
  NAND2_X1 U28341 ( .A1(n17546), .A2(n17440), .ZN(n17427) );
  AND2_X1 U28342 ( .A1(n18060), .A2(n18062), .ZN(n17439) );
  AOI21_X1 U28343 ( .B1(n17553), .B2(n17428), .A(n17439), .ZN(n17429) );
  NAND2_X1 U28344 ( .A1(n17431), .A2(n18071), .ZN(n18340) );
  INV_X1 U28345 ( .A(n18342), .ZN(n17433) );
  AND2_X1 U28346 ( .A1(n18340), .A2(n17434), .ZN(n17445) );
  AOI21_X1 U28347 ( .B1(n17436), .B2(n17435), .A(n17546), .ZN(n17438) );
  OAI21_X1 U28348 ( .B1(n17438), .B2(n17437), .A(n18064), .ZN(n17444) );
  INV_X1 U28349 ( .A(n17439), .ZN(n17442) );
  NAND4_X1 U28350 ( .A1(n17442), .A2(n17441), .A3(n17553), .A4(n17546), .ZN(
        n17443) );
  INV_X1 U28351 ( .A(n17446), .ZN(n17450) );
  INV_X1 U28352 ( .A(n17447), .ZN(n17449) );
  INV_X1 U28353 ( .A(n17448), .ZN(n17460) );
  AOI22_X1 U28354 ( .A1(n17450), .A2(n51440), .B1(n17449), .B2(n17460), .ZN(
        n17455) );
  OAI21_X1 U28355 ( .B1(n18376), .B2(n5385), .A(n6711), .ZN(n17452) );
  OAI21_X1 U28356 ( .B1(n17452), .B2(n51440), .A(n20032), .ZN(n17453) );
  NAND3_X1 U28357 ( .A1(n17455), .A2(n17454), .A3(n17453), .ZN(n17465) );
  INV_X1 U28358 ( .A(n17456), .ZN(n18373) );
  NAND3_X1 U28359 ( .A1(n17457), .A2(n20037), .A3(n18373), .ZN(n17463) );
  INV_X1 U28360 ( .A(n17458), .ZN(n17459) );
  AOI22_X1 U28361 ( .A1(n17460), .A2(n17459), .B1(n20040), .B2(n20046), .ZN(
        n17462) );
  NAND3_X1 U28362 ( .A1(n17463), .A2(n17462), .A3(n17461), .ZN(n17464) );
  OR2_X2 U28363 ( .A1(n17465), .A2(n17464), .ZN(n23341) );
  OAI21_X1 U28364 ( .B1(n17871), .B2(n18034), .A(n19408), .ZN(n17468) );
  INV_X1 U28365 ( .A(n18034), .ZN(n19426) );
  AND2_X1 U28366 ( .A1(n2222), .A2(n19426), .ZN(n17467) );
  INV_X1 U28367 ( .A(n18032), .ZN(n17469) );
  INV_X1 U28369 ( .A(n19408), .ZN(n17476) );
  AOI21_X1 U28370 ( .B1(n17474), .B2(n18032), .A(n18041), .ZN(n17475) );
  OAI211_X1 U28371 ( .C1(n17476), .C2(n19425), .A(n17475), .B(n2222), .ZN(
        n21746) );
  OAI22_X1 U28372 ( .A1(n18023), .A2(n19396), .B1(n18015), .B2(n19388), .ZN(
        n17477) );
  NAND2_X1 U28373 ( .A1(n17477), .A2(n3714), .ZN(n17483) );
  OAI211_X1 U28376 ( .C1(n17479), .C2(n17568), .A(n17478), .B(n19398), .ZN(
        n17482) );
  AND3_X1 U28377 ( .A1(n17569), .A2(n17568), .A3(n17479), .ZN(n18021) );
  INV_X1 U28378 ( .A(n18021), .ZN(n17481) );
  INV_X1 U28379 ( .A(n19398), .ZN(n18007) );
  NAND3_X1 U28380 ( .A1(n19395), .A2(n18007), .A3(n19389), .ZN(n17480) );
  MUX2_X1 U28381 ( .A(n19389), .B(n17484), .S(n19396), .Z(n17574) );
  INV_X1 U28382 ( .A(n17574), .ZN(n17486) );
  NAND2_X1 U28383 ( .A1(n18012), .A2(n3865), .ZN(n17485) );
  NAND2_X1 U28384 ( .A1(n23341), .A2(n21744), .ZN(n23338) );
  INV_X1 U28385 ( .A(n23338), .ZN(n21148) );
  NAND2_X1 U28386 ( .A1(n17487), .A2(n633), .ZN(n17488) );
  NAND2_X1 U28387 ( .A1(n17488), .A2(n18287), .ZN(n17495) );
  NOR2_X1 U28388 ( .A1(n20014), .A2(n17489), .ZN(n17490) );
  INV_X1 U28389 ( .A(n18285), .ZN(n17492) );
  OAI21_X1 U28390 ( .B1(n17491), .B2(n17490), .A(n17492), .ZN(n17494) );
  INV_X1 U28392 ( .A(n20086), .ZN(n18317) );
  NAND3_X1 U28393 ( .A1(n18317), .A2(n20096), .A3(n16788), .ZN(n17497) );
  OAI211_X1 U28394 ( .C1(n17600), .C2(n20087), .A(n17498), .B(n17497), .ZN(
        n17500) );
  NAND2_X1 U28395 ( .A1(n17596), .A2(n20095), .ZN(n17502) );
  NAND2_X1 U28396 ( .A1(n20092), .A2(n20094), .ZN(n17501) );
  INV_X1 U28397 ( .A(n18316), .ZN(n17604) );
  NAND3_X1 U28398 ( .A1(n18322), .A2(n17604), .A3(n17506), .ZN(n17508) );
  AOI21_X1 U28399 ( .B1(n17506), .B2(n18318), .A(n17505), .ZN(n17507) );
  NAND3_X1 U28400 ( .A1(n1024), .A2(n22256), .A3(n21744), .ZN(n17511) );
  NOR2_X1 U28401 ( .A1(n17511), .A2(n21756), .ZN(n17512) );
  NAND2_X1 U28402 ( .A1(n22263), .A2(n17513), .ZN(n17514) );
  NAND2_X1 U28403 ( .A1(n21756), .A2(n21755), .ZN(n22261) );
  NAND2_X1 U28404 ( .A1(n18287), .A2(n590), .ZN(n18286) );
  OAI21_X1 U28405 ( .B1(n18282), .B2(n18286), .A(n17516), .ZN(n17518) );
  INV_X1 U28406 ( .A(n20019), .ZN(n17517) );
  NAND3_X1 U28407 ( .A1(n51208), .A2(n6952), .A3(n20015), .ZN(n17519) );
  OAI21_X1 U28408 ( .B1(n17523), .B2(n17522), .A(n17521), .ZN(n17524) );
  NAND2_X1 U28409 ( .A1(n17524), .A2(n633), .ZN(n17531) );
  INV_X1 U28410 ( .A(n17525), .ZN(n20011) );
  NAND3_X1 U28412 ( .A1(n20013), .A2(n16798), .A3(n2166), .ZN(n17527) );
  NAND2_X1 U28413 ( .A1(n17528), .A2(n17527), .ZN(n17530) );
  AOI22_X1 U28414 ( .A1(n17531), .A2(n20011), .B1(n17530), .B2(n17529), .ZN(
        n17539) );
  INV_X1 U28415 ( .A(n17533), .ZN(n20022) );
  AOI22_X1 U28416 ( .A1(n20022), .A2(n20023), .B1(n17534), .B2(n6952), .ZN(
        n17536) );
  MUX2_X1 U28417 ( .A(n17537), .B(n17536), .S(n17535), .Z(n17538) );
  NOR2_X1 U28418 ( .A1(n17542), .A2(n17553), .ZN(n17543) );
  AOI22_X1 U28419 ( .A1(n18326), .A2(n17543), .B1(n18062), .B2(n17542), .ZN(
        n17551) );
  NAND3_X1 U28420 ( .A1(n18071), .A2(n18331), .A3(n17544), .ZN(n17550) );
  NAND3_X1 U28421 ( .A1(n18074), .A2(n18064), .A3(n17545), .ZN(n17549) );
  NOR2_X1 U28422 ( .A1(n17546), .A2(n18063), .ZN(n17547) );
  OAI21_X1 U28423 ( .B1(n18332), .B2(n17547), .A(n18326), .ZN(n17548) );
  AND4_X1 U28424 ( .A1(n17551), .A2(n17550), .A3(n17549), .A4(n17548), .ZN(
        n17552) );
  NOR2_X1 U28425 ( .A1(n18032), .A2(n18039), .ZN(n18031) );
  AOI22_X1 U28426 ( .A1(n17557), .A2(n6332), .B1(n19410), .B2(n18040), .ZN(
        n17554) );
  OAI21_X1 U28427 ( .B1(n18031), .B2(n17554), .A(n18037), .ZN(n17563) );
  INV_X1 U28428 ( .A(n17870), .ZN(n17556) );
  NAND3_X1 U28429 ( .A1(n19411), .A2(n17873), .A3(n6332), .ZN(n17555) );
  NAND3_X1 U28430 ( .A1(n19424), .A2(n19426), .A3(n19417), .ZN(n17562) );
  OAI21_X1 U28431 ( .B1(n8378), .B2(n17557), .A(n18043), .ZN(n17560) );
  NOR2_X1 U28432 ( .A1(n22155), .A2(n22140), .ZN(n19565) );
  NAND3_X1 U28433 ( .A1(n19396), .A2(n17577), .A3(n19388), .ZN(n17564) );
  INV_X1 U28434 ( .A(n19395), .ZN(n17565) );
  NOR2_X1 U28435 ( .A1(n18009), .A2(n17568), .ZN(n17570) );
  OAI211_X1 U28436 ( .C1(n18008), .C2(n17570), .A(n17569), .B(n17575), .ZN(
        n17571) );
  INV_X1 U28440 ( .A(n17575), .ZN(n17578) );
  INV_X1 U28441 ( .A(n19397), .ZN(n17581) );
  INV_X1 U28442 ( .A(n19348), .ZN(n17585) );
  INV_X1 U28443 ( .A(n18081), .ZN(n17621) );
  OAI22_X1 U28444 ( .A1(n17585), .A2(n17621), .B1(n18080), .B2(n20512), .ZN(
        n17586) );
  NAND2_X1 U28445 ( .A1(n17586), .A2(n19344), .ZN(n17593) );
  NAND3_X1 U28446 ( .A1(n18086), .A2(n20513), .A3(n18081), .ZN(n20519) );
  NAND3_X1 U28447 ( .A1(n18086), .A2(n20503), .A3(n489), .ZN(n17587) );
  INV_X1 U28448 ( .A(n17627), .ZN(n17626) );
  NAND3_X1 U28449 ( .A1(n17626), .A2(n17589), .A3(n18081), .ZN(n17588) );
  AND2_X1 U28450 ( .A1(n18077), .A2(n17588), .ZN(n17592) );
  NAND3_X1 U28451 ( .A1(n17589), .A2(n20507), .A3(n18081), .ZN(n19335) );
  NAND2_X1 U28452 ( .A1(n20513), .A2(n489), .ZN(n18076) );
  NAND2_X1 U28453 ( .A1(n19335), .A2(n18076), .ZN(n17590) );
  NAND2_X1 U28454 ( .A1(n17590), .A2(n18075), .ZN(n17591) );
  NOR2_X1 U28455 ( .A1(n51661), .A2(n22140), .ZN(n22146) );
  AOI21_X1 U28456 ( .B1(n20092), .B2(n20088), .A(n20094), .ZN(n17594) );
  NAND2_X1 U28457 ( .A1(n18312), .A2(n17594), .ZN(n17598) );
  OAI21_X1 U28458 ( .B1(n20100), .B2(n20104), .A(n20086), .ZN(n17595) );
  NAND2_X1 U28459 ( .A1(n17596), .A2(n17595), .ZN(n17597) );
  AND2_X1 U28460 ( .A1(n17599), .A2(n20096), .ZN(n17602) );
  AND2_X1 U28461 ( .A1(n18316), .A2(n17600), .ZN(n17601) );
  NAND2_X1 U28463 ( .A1(n17607), .A2(n20097), .ZN(n17606) );
  INV_X1 U28465 ( .A(n21934), .ZN(n17610) );
  NAND2_X1 U28466 ( .A1(n22154), .A2(n22155), .ZN(n22156) );
  INV_X1 U28467 ( .A(n21935), .ZN(n17609) );
  OAI21_X1 U28468 ( .B1(n20952), .B2(n19560), .A(n22154), .ZN(n17614) );
  NOR2_X1 U28469 ( .A1(n17612), .A2(n2488), .ZN(n17613) );
  INV_X1 U28470 ( .A(n22152), .ZN(n21025) );
  XNOR2_X1 U28472 ( .A(n24736), .B(n24344), .ZN(n17996) );
  NAND2_X1 U28473 ( .A1(n18075), .A2(n17625), .ZN(n17617) );
  INV_X1 U28474 ( .A(n20511), .ZN(n17624) );
  NAND2_X1 U28475 ( .A1(n20515), .A2(n18085), .ZN(n17620) );
  AND2_X1 U28476 ( .A1(n19337), .A2(n17620), .ZN(n17623) );
  NAND3_X1 U28477 ( .A1(n20508), .A2(n19344), .A3(n18081), .ZN(n17630) );
  NAND3_X1 U28478 ( .A1(n17627), .A2(n20513), .A3(n18081), .ZN(n17628) );
  NAND2_X1 U28480 ( .A1(n51704), .A2(n18085), .ZN(n19345) );
  NAND2_X1 U28481 ( .A1(n19335), .A2(n19345), .ZN(n17633) );
  NAND2_X1 U28482 ( .A1(n17633), .A2(n20501), .ZN(n22355) );
  NAND2_X1 U28483 ( .A1(n20472), .A2(n20383), .ZN(n20388) );
  AND2_X1 U28484 ( .A1(n17639), .A2(n20478), .ZN(n20476) );
  NAND3_X1 U28485 ( .A1(n20462), .A2(n20466), .A3(n20389), .ZN(n17634) );
  OAI211_X1 U28486 ( .C1(n20388), .C2(n17636), .A(n17635), .B(n17634), .ZN(
        n17637) );
  INV_X1 U28487 ( .A(n17637), .ZN(n17642) );
  OAI21_X1 U28488 ( .B1(n20399), .B2(n19371), .A(n20474), .ZN(n17638) );
  NAND2_X1 U28489 ( .A1(n17638), .A2(n20477), .ZN(n17641) );
  AND2_X1 U28490 ( .A1(n17639), .A2(n20474), .ZN(n20460) );
  INV_X1 U28491 ( .A(n20460), .ZN(n17640) );
  NAND3_X1 U28492 ( .A1(n17640), .A2(n17997), .A3(n20468), .ZN(n18006) );
  NAND4_X1 U28494 ( .A1(n17642), .A2(n17641), .A3(n18006), .A4(n20465), .ZN(
        n22367) );
  XNOR2_X1 U28495 ( .A(n17644), .B(n17643), .ZN(n17943) );
  XNOR2_X1 U28496 ( .A(n17645), .B(n17943), .ZN(n17650) );
  XNOR2_X1 U28497 ( .A(n17646), .B(n4589), .ZN(n18579) );
  XNOR2_X1 U28498 ( .A(n17647), .B(n17648), .ZN(n17649) );
  XNOR2_X1 U28499 ( .A(n17652), .B(n17651), .ZN(n17659) );
  XNOR2_X1 U28500 ( .A(n43293), .B(n24820), .ZN(n35093) );
  XNOR2_X1 U28501 ( .A(n35093), .B(n43691), .ZN(n17653) );
  XNOR2_X1 U28502 ( .A(n27388), .B(n18206), .ZN(n35641) );
  XNOR2_X1 U28503 ( .A(n17653), .B(n35641), .ZN(n17655) );
  XNOR2_X1 U28504 ( .A(n4353), .B(n49429), .ZN(n26207) );
  XNOR2_X1 U28505 ( .A(n23370), .B(n26207), .ZN(n17654) );
  XNOR2_X1 U28506 ( .A(n46097), .B(n17654), .ZN(n35221) );
  XNOR2_X1 U28507 ( .A(n17655), .B(n35221), .ZN(n17656) );
  XNOR2_X1 U28508 ( .A(n17812), .B(n17656), .ZN(n17657) );
  XNOR2_X1 U28509 ( .A(n17657), .B(n18790), .ZN(n17658) );
  XNOR2_X1 U28510 ( .A(n17659), .B(n17658), .ZN(n17660) );
  XNOR2_X1 U28511 ( .A(n17661), .B(n25897), .ZN(n25382) );
  XNOR2_X1 U28512 ( .A(n2602), .B(n4837), .ZN(n25380) );
  XNOR2_X1 U28513 ( .A(n25380), .B(n4286), .ZN(n25097) );
  XNOR2_X1 U28514 ( .A(n25382), .B(n25097), .ZN(n34589) );
  XNOR2_X1 U28515 ( .A(n27185), .B(n24553), .ZN(n33698) );
  XNOR2_X1 U28516 ( .A(n49937), .B(n48843), .ZN(n17662) );
  XNOR2_X1 U28517 ( .A(n33698), .B(n17662), .ZN(n17663) );
  XNOR2_X1 U28518 ( .A(n34589), .B(n17663), .ZN(n17664) );
  XNOR2_X1 U28519 ( .A(n17665), .B(n17664), .ZN(n17666) );
  XNOR2_X1 U28520 ( .A(n52227), .B(n17786), .ZN(n17668) );
  XNOR2_X1 U28521 ( .A(n18437), .B(n17923), .ZN(n17667) );
  XNOR2_X1 U28522 ( .A(n17668), .B(n17667), .ZN(n17669) );
  XNOR2_X1 U28523 ( .A(n17669), .B(n17670), .ZN(n17675) );
  XNOR2_X1 U28524 ( .A(n51458), .B(n17788), .ZN(n17673) );
  INV_X1 U28525 ( .A(n18196), .ZN(n17672) );
  XNOR2_X1 U28526 ( .A(n17673), .B(n17672), .ZN(n17674) );
  XNOR2_X1 U28527 ( .A(n18447), .B(n18443), .ZN(n17676) );
  XNOR2_X1 U28528 ( .A(n17787), .B(n17676), .ZN(n18198) );
  XNOR2_X1 U28529 ( .A(n17678), .B(n17677), .ZN(n18619) );
  XNOR2_X1 U28530 ( .A(n47268), .B(n4247), .ZN(n35251) );
  XNOR2_X1 U28531 ( .A(n19261), .B(n35251), .ZN(n18593) );
  XNOR2_X1 U28532 ( .A(n18457), .B(n18593), .ZN(n17682) );
  XNOR2_X1 U28533 ( .A(n18602), .B(n51134), .ZN(n17680) );
  XNOR2_X1 U28534 ( .A(n17680), .B(n17679), .ZN(n17681) );
  XNOR2_X1 U28535 ( .A(n17682), .B(n17681), .ZN(n17689) );
  XNOR2_X1 U28536 ( .A(n44495), .B(n34232), .ZN(n25779) );
  XNOR2_X1 U28537 ( .A(n43739), .B(n26603), .ZN(n46144) );
  XNOR2_X1 U28538 ( .A(n46144), .B(n23882), .ZN(n17683) );
  XNOR2_X1 U28539 ( .A(n25779), .B(n17683), .ZN(n33768) );
  XNOR2_X1 U28540 ( .A(n17684), .B(n4721), .ZN(n42329) );
  XNOR2_X1 U28541 ( .A(n42329), .B(n2203), .ZN(n17685) );
  XNOR2_X1 U28542 ( .A(n18749), .B(n17686), .ZN(n17687) );
  XNOR2_X1 U28543 ( .A(n17687), .B(n18714), .ZN(n17688) );
  XNOR2_X1 U28544 ( .A(n17689), .B(n17688), .ZN(n17696) );
  XNOR2_X1 U28545 ( .A(n17690), .B(n17973), .ZN(n17693) );
  XNOR2_X1 U28546 ( .A(n17693), .B(n17692), .ZN(n17834) );
  XNOR2_X1 U28547 ( .A(n17834), .B(n17694), .ZN(n17695) );
  XNOR2_X2 U28548 ( .A(n17696), .B(n17695), .ZN(n21468) );
  INV_X1 U28549 ( .A(n21468), .ZN(n20487) );
  XNOR2_X1 U28550 ( .A(n17697), .B(n2135), .ZN(n18768) );
  XNOR2_X1 U28551 ( .A(n18147), .B(n19199), .ZN(n17703) );
  XNOR2_X1 U28552 ( .A(n33050), .B(n20856), .ZN(n34255) );
  XNOR2_X1 U28553 ( .A(n4739), .B(n4868), .ZN(n43150) );
  XNOR2_X1 U28554 ( .A(n34255), .B(n43150), .ZN(n34776) );
  XNOR2_X1 U28555 ( .A(n45107), .B(n4045), .ZN(n18513) );
  XNOR2_X1 U28556 ( .A(n4637), .B(n4605), .ZN(n20857) );
  XNOR2_X1 U28557 ( .A(n18513), .B(n20857), .ZN(n33933) );
  XNOR2_X1 U28558 ( .A(n22814), .B(n4793), .ZN(n27204) );
  XNOR2_X1 U28559 ( .A(n4937), .B(n4501), .ZN(n17698) );
  XNOR2_X1 U28560 ( .A(n27204), .B(n17698), .ZN(n17699) );
  XNOR2_X1 U28561 ( .A(n33933), .B(n17699), .ZN(n17700) );
  XNOR2_X1 U28562 ( .A(n34776), .B(n17700), .ZN(n17701) );
  XNOR2_X1 U28563 ( .A(n17764), .B(n17701), .ZN(n17702) );
  XNOR2_X1 U28564 ( .A(n17703), .B(n17702), .ZN(n17704) );
  XNOR2_X1 U28565 ( .A(n18768), .B(n17704), .ZN(n17706) );
  XNOR2_X1 U28566 ( .A(n17706), .B(n17705), .ZN(n17711) );
  XNOR2_X1 U28567 ( .A(n19198), .B(n17756), .ZN(n17709) );
  XNOR2_X1 U28568 ( .A(n17707), .B(n18668), .ZN(n17708) );
  XNOR2_X1 U28569 ( .A(n18148), .B(n17708), .ZN(n17894) );
  XNOR2_X1 U28570 ( .A(n17709), .B(n17894), .ZN(n17710) );
  NAND2_X1 U28571 ( .A1(n20487), .A2(n20314), .ZN(n17712) );
  INV_X1 U28572 ( .A(n20314), .ZN(n17740) );
  XNOR2_X1 U28573 ( .A(n17714), .B(n17713), .ZN(n17721) );
  XNOR2_X1 U28574 ( .A(n17901), .B(n2121), .ZN(n17715) );
  XNOR2_X1 U28575 ( .A(n461), .B(n17715), .ZN(n17719) );
  XNOR2_X1 U28576 ( .A(n17716), .B(n4705), .ZN(n25720) );
  XNOR2_X1 U28577 ( .A(n25720), .B(n26370), .ZN(n36878) );
  XNOR2_X1 U28578 ( .A(n24227), .B(n24830), .ZN(n32657) );
  XNOR2_X1 U28579 ( .A(n36878), .B(n32657), .ZN(n17717) );
  XNOR2_X1 U28580 ( .A(n52167), .B(n17717), .ZN(n17718) );
  XNOR2_X1 U28581 ( .A(n17719), .B(n17718), .ZN(n17720) );
  XNOR2_X1 U28582 ( .A(n17721), .B(n17720), .ZN(n17724) );
  XNOR2_X1 U28583 ( .A(n18660), .B(n17722), .ZN(n17723) );
  XNOR2_X1 U28584 ( .A(n17728), .B(n43073), .ZN(n32497) );
  XNOR2_X1 U28585 ( .A(n43766), .B(n4204), .ZN(n36837) );
  XNOR2_X1 U28586 ( .A(n32497), .B(n36837), .ZN(n17729) );
  XNOR2_X1 U28587 ( .A(n17730), .B(n17729), .ZN(n17732) );
  XNOR2_X1 U28588 ( .A(n17732), .B(n17731), .ZN(n17733) );
  XNOR2_X1 U28589 ( .A(n18831), .B(n42889), .ZN(n18565) );
  INV_X1 U28590 ( .A(n18565), .ZN(n17735) );
  XNOR2_X1 U28591 ( .A(n18475), .B(n18690), .ZN(n17734) );
  XNOR2_X1 U28592 ( .A(n17735), .B(n17734), .ZN(n17736) );
  XNOR2_X1 U28593 ( .A(n17736), .B(n18564), .ZN(n17737) );
  XNOR2_X1 U28594 ( .A(n17738), .B(n17737), .ZN(n17739) );
  AND2_X1 U28595 ( .A1(n21463), .A2(n21450), .ZN(n19352) );
  NAND2_X1 U28596 ( .A1(n21468), .A2(n20493), .ZN(n21452) );
  INV_X1 U28597 ( .A(n21452), .ZN(n19364) );
  NAND2_X1 U28598 ( .A1(n19364), .A2(n20314), .ZN(n17742) );
  NAND2_X1 U28599 ( .A1(n21460), .A2(n21469), .ZN(n17741) );
  AND3_X1 U28600 ( .A1(n17743), .A2(n17742), .A3(n17741), .ZN(n17749) );
  NAND2_X1 U28601 ( .A1(n21463), .A2(n21465), .ZN(n17744) );
  AND2_X1 U28602 ( .A1(n52146), .A2(n17744), .ZN(n17746) );
  OAI21_X1 U28603 ( .B1(n21464), .B2(n21468), .A(n21451), .ZN(n17745) );
  AOI22_X1 U28604 ( .A1(n17747), .A2(n17746), .B1(n17745), .B2(n20316), .ZN(
        n17748) );
  XNOR2_X1 U28605 ( .A(n45105), .B(n4739), .ZN(n17751) );
  XNOR2_X1 U28606 ( .A(n41496), .B(n4638), .ZN(n25685) );
  XNOR2_X1 U28607 ( .A(n27203), .B(n24919), .ZN(n17750) );
  XNOR2_X1 U28608 ( .A(n25685), .B(n17750), .ZN(n34878) );
  XNOR2_X1 U28609 ( .A(n17751), .B(n34878), .ZN(n17752) );
  XNOR2_X1 U28610 ( .A(n43202), .B(n4885), .ZN(n42419) );
  XNOR2_X1 U28611 ( .A(n17752), .B(n42419), .ZN(n17753) );
  XNOR2_X1 U28612 ( .A(n17891), .B(n17753), .ZN(n17755) );
  XNOR2_X1 U28613 ( .A(n17758), .B(n17757), .ZN(n17759) );
  XNOR2_X1 U28614 ( .A(n17759), .B(n2136), .ZN(n18673) );
  XNOR2_X1 U28615 ( .A(n17760), .B(n18673), .ZN(n17762) );
  XNOR2_X1 U28616 ( .A(n17762), .B(n17761), .ZN(n17769) );
  XNOR2_X1 U28617 ( .A(n17764), .B(n17763), .ZN(n17765) );
  XNOR2_X1 U28618 ( .A(n17766), .B(n17765), .ZN(n17767) );
  XNOR2_X1 U28619 ( .A(n17768), .B(n17767), .ZN(n18526) );
  XNOR2_X1 U28620 ( .A(n17770), .B(n19216), .ZN(n17783) );
  XNOR2_X1 U28621 ( .A(n2162), .B(n17771), .ZN(n17772) );
  XNOR2_X1 U28622 ( .A(n461), .B(n17772), .ZN(n17781) );
  XNOR2_X1 U28623 ( .A(n26541), .B(n4515), .ZN(n28267) );
  XNOR2_X1 U28624 ( .A(n25575), .B(n28267), .ZN(n17775) );
  XNOR2_X1 U28625 ( .A(n25793), .B(n17773), .ZN(n17774) );
  XNOR2_X1 U28626 ( .A(n17775), .B(n17774), .ZN(n31807) );
  XNOR2_X1 U28627 ( .A(n38626), .B(n3383), .ZN(n24523) );
  XNOR2_X1 U28628 ( .A(n24523), .B(n2605), .ZN(n17776) );
  XNOR2_X1 U28629 ( .A(n31807), .B(n17776), .ZN(n17777) );
  XNOR2_X1 U28630 ( .A(n18539), .B(n17777), .ZN(n17779) );
  XNOR2_X1 U28631 ( .A(n17779), .B(n17778), .ZN(n17780) );
  XNOR2_X1 U28632 ( .A(n17781), .B(n17780), .ZN(n17782) );
  XNOR2_X1 U28634 ( .A(n17787), .B(n17786), .ZN(n17789) );
  XNOR2_X1 U28635 ( .A(n17789), .B(n17788), .ZN(n17796) );
  XNOR2_X1 U28636 ( .A(n25097), .B(n26525), .ZN(n34332) );
  XNOR2_X1 U28637 ( .A(n34332), .B(n1354), .ZN(n17791) );
  XNOR2_X1 U28638 ( .A(n27186), .B(n42721), .ZN(n17790) );
  XNOR2_X1 U28639 ( .A(n17790), .B(n26403), .ZN(n33612) );
  XNOR2_X1 U28640 ( .A(n17791), .B(n33612), .ZN(n17792) );
  XNOR2_X1 U28641 ( .A(n17793), .B(n17792), .ZN(n17794) );
  XNOR2_X1 U28642 ( .A(n17795), .B(n17796), .ZN(n17797) );
  XNOR2_X1 U28643 ( .A(n17797), .B(n18553), .ZN(n17801) );
  XNOR2_X1 U28644 ( .A(n17798), .B(n2218), .ZN(n17799) );
  XNOR2_X1 U28645 ( .A(n51414), .B(n17799), .ZN(n17800) );
  XNOR2_X1 U28646 ( .A(n17804), .B(n47737), .ZN(n17805) );
  XNOR2_X1 U28647 ( .A(n17806), .B(n17805), .ZN(n18806) );
  XNOR2_X1 U28648 ( .A(n17807), .B(n18806), .ZN(n17818) );
  XNOR2_X1 U28649 ( .A(n23370), .B(n24820), .ZN(n24641) );
  XNOR2_X1 U28650 ( .A(n18636), .B(n4886), .ZN(n17808) );
  XNOR2_X1 U28651 ( .A(n24641), .B(n17808), .ZN(n35340) );
  XNOR2_X1 U28652 ( .A(n35340), .B(n17809), .ZN(n17810) );
  XNOR2_X1 U28653 ( .A(n17810), .B(n35541), .ZN(n17811) );
  XNOR2_X1 U28654 ( .A(n17812), .B(n17811), .ZN(n17813) );
  XNOR2_X1 U28655 ( .A(n17814), .B(n17813), .ZN(n17815) );
  XNOR2_X1 U28656 ( .A(n17816), .B(n17815), .ZN(n17817) );
  XNOR2_X1 U28657 ( .A(n18464), .B(n17821), .ZN(n17824) );
  XNOR2_X1 U28658 ( .A(n18712), .B(n51134), .ZN(n17823) );
  XNOR2_X1 U28659 ( .A(n17824), .B(n17823), .ZN(n17833) );
  XNOR2_X1 U28660 ( .A(n25284), .B(n41740), .ZN(n24925) );
  XNOR2_X1 U28661 ( .A(n24925), .B(n17825), .ZN(n34398) );
  XNOR2_X1 U28662 ( .A(n4916), .B(n4782), .ZN(n17826) );
  XNOR2_X1 U28663 ( .A(n17826), .B(n4923), .ZN(n17827) );
  XNOR2_X1 U28664 ( .A(n46144), .B(n17827), .ZN(n33568) );
  XNOR2_X1 U28665 ( .A(n34398), .B(n33568), .ZN(n17828) );
  XNOR2_X1 U28666 ( .A(n17829), .B(n17828), .ZN(n17830) );
  XNOR2_X1 U28667 ( .A(n17831), .B(n17830), .ZN(n17832) );
  XNOR2_X1 U28668 ( .A(n17833), .B(n17832), .ZN(n17835) );
  XNOR2_X1 U28669 ( .A(n17835), .B(n17834), .ZN(n17836) );
  INV_X1 U28670 ( .A(n17856), .ZN(n20427) );
  NAND2_X1 U28671 ( .A1(n20434), .A2(n20427), .ZN(n20358) );
  OAI21_X1 U28673 ( .B1(n18053), .B2(n20358), .A(n20362), .ZN(n17855) );
  XNOR2_X1 U28674 ( .A(n17840), .B(n17839), .ZN(n17842) );
  XNOR2_X1 U28675 ( .A(n17841), .B(n51454), .ZN(n18568) );
  XNOR2_X1 U28676 ( .A(n52183), .B(n18564), .ZN(n17850) );
  XNOR2_X1 U28677 ( .A(n18570), .B(n17844), .ZN(n42293) );
  XNOR2_X1 U28678 ( .A(n42293), .B(n4048), .ZN(n36667) );
  XNOR2_X1 U28679 ( .A(n31432), .B(n4526), .ZN(n17845) );
  XNOR2_X1 U28680 ( .A(n36667), .B(n17845), .ZN(n17846) );
  XNOR2_X1 U28681 ( .A(n17847), .B(n17846), .ZN(n17848) );
  XNOR2_X1 U28682 ( .A(n17848), .B(n18696), .ZN(n17849) );
  INV_X1 U28684 ( .A(n20349), .ZN(n17853) );
  NAND3_X1 U28685 ( .A1(n20434), .A2(n19173), .A3(n20428), .ZN(n17852) );
  INV_X1 U28686 ( .A(n19326), .ZN(n17858) );
  NAND2_X1 U28687 ( .A1(n18053), .A2(n20426), .ZN(n19331) );
  NAND2_X1 U28688 ( .A1(n19170), .A2(n20422), .ZN(n18052) );
  INV_X1 U28689 ( .A(n18052), .ZN(n17857) );
  OAI211_X1 U28690 ( .C1(n50), .C2(n17858), .A(n19331), .B(n17857), .ZN(n17863) );
  NOR2_X1 U28691 ( .A1(n20343), .A2(n20427), .ZN(n17860) );
  OAI22_X1 U28692 ( .A1(n17860), .A2(n19322), .B1(n19324), .B2(n20428), .ZN(
        n17861) );
  NAND2_X1 U28693 ( .A1(n19424), .A2(n19418), .ZN(n17866) );
  NAND3_X1 U28694 ( .A1(n19404), .A2(n19418), .A3(n17871), .ZN(n17865) );
  AND3_X1 U28695 ( .A1(n17867), .A2(n17866), .A3(n17865), .ZN(n17878) );
  NAND2_X1 U28696 ( .A1(n17868), .A2(n17469), .ZN(n17877) );
  NAND3_X1 U28697 ( .A1(n17870), .A2(n17869), .A3(n18043), .ZN(n19434) );
  AOI21_X1 U28698 ( .B1(n17872), .B2(n6605), .A(n18041), .ZN(n17875) );
  NAND2_X1 U28699 ( .A1(n22918), .A2(n22359), .ZN(n22362) );
  NAND3_X1 U28700 ( .A1(n19576), .A2(n2175), .A3(n22362), .ZN(n17990) );
  NAND2_X1 U28701 ( .A1(n22913), .A2(n5542), .ZN(n17989) );
  XNOR2_X1 U28702 ( .A(n17879), .B(n14903), .ZN(n17885) );
  XNOR2_X1 U28703 ( .A(n45107), .B(n42630), .ZN(n17881) );
  XNOR2_X1 U28704 ( .A(n17881), .B(n17880), .ZN(n18759) );
  XNOR2_X1 U28705 ( .A(n18759), .B(n4605), .ZN(n24843) );
  XNOR2_X1 U28706 ( .A(n41496), .B(n28376), .ZN(n17882) );
  XNOR2_X1 U28707 ( .A(n28252), .B(n17882), .ZN(n17883) );
  XNOR2_X1 U28708 ( .A(n24843), .B(n17883), .ZN(n34071) );
  XNOR2_X1 U28709 ( .A(n18399), .B(n34071), .ZN(n17884) );
  XNOR2_X1 U28710 ( .A(n17885), .B(n17884), .ZN(n17886) );
  XNOR2_X1 U28711 ( .A(n14427), .B(n18409), .ZN(n17888) );
  XNOR2_X1 U28712 ( .A(n51668), .B(n17890), .ZN(n18769) );
  XNOR2_X1 U28713 ( .A(n44044), .B(n4343), .ZN(n33295) );
  XNOR2_X1 U28714 ( .A(n33295), .B(n22814), .ZN(n33793) );
  XNOR2_X1 U28715 ( .A(n19199), .B(n33793), .ZN(n17893) );
  INV_X1 U28716 ( .A(n17891), .ZN(n17892) );
  XNOR2_X1 U28717 ( .A(n17893), .B(n17892), .ZN(n18677) );
  XNOR2_X1 U28718 ( .A(n2113), .B(n18677), .ZN(n17895) );
  XNOR2_X1 U28719 ( .A(n17895), .B(n17894), .ZN(n17896) );
  XNOR2_X1 U28720 ( .A(n18780), .B(n32627), .ZN(n17898) );
  XNOR2_X1 U28721 ( .A(n17898), .B(n17897), .ZN(n19223) );
  XNOR2_X1 U28722 ( .A(n38626), .B(n4482), .ZN(n17899) );
  INV_X1 U28723 ( .A(n24430), .ZN(n43640) );
  XNOR2_X1 U28724 ( .A(n17899), .B(n43640), .ZN(n25956) );
  XNOR2_X1 U28725 ( .A(n25956), .B(n33653), .ZN(n18776) );
  XNOR2_X1 U28726 ( .A(n18776), .B(n21089), .ZN(n33166) );
  XNOR2_X1 U28727 ( .A(n33166), .B(n36994), .ZN(n17900) );
  XNOR2_X1 U28729 ( .A(n17902), .B(n17901), .ZN(n17903) );
  XNOR2_X1 U28730 ( .A(n17904), .B(n17903), .ZN(n17905) );
  XNOR2_X1 U28731 ( .A(n19223), .B(n17905), .ZN(n17910) );
  XNOR2_X1 U28732 ( .A(n17908), .B(n17907), .ZN(n17909) );
  XNOR2_X1 U28733 ( .A(n17911), .B(n17912), .ZN(n17917) );
  XNOR2_X1 U28734 ( .A(n17914), .B(n2215), .ZN(n17915) );
  XNOR2_X1 U28735 ( .A(n17916), .B(n17915), .ZN(n18787) );
  XNOR2_X1 U28736 ( .A(n17918), .B(n18619), .ZN(n17919) );
  XNOR2_X1 U28737 ( .A(n18817), .B(n17919), .ZN(n17930) );
  XNOR2_X1 U28738 ( .A(n51133), .B(n18617), .ZN(n17928) );
  XNOR2_X1 U28739 ( .A(n28116), .B(n25434), .ZN(n26223) );
  XNOR2_X1 U28740 ( .A(n4744), .B(n4879), .ZN(n17920) );
  XNOR2_X1 U28741 ( .A(n28391), .B(n17920), .ZN(n34450) );
  XNOR2_X1 U28742 ( .A(n34450), .B(n41660), .ZN(n17921) );
  XNOR2_X1 U28743 ( .A(n26223), .B(n17921), .ZN(n17922) );
  XNOR2_X1 U28744 ( .A(n17923), .B(n17922), .ZN(n17924) );
  XNOR2_X1 U28745 ( .A(n17925), .B(n17924), .ZN(n17926) );
  XNOR2_X1 U28746 ( .A(n18615), .B(n17926), .ZN(n17927) );
  XNOR2_X1 U28747 ( .A(n17928), .B(n17927), .ZN(n17929) );
  XNOR2_X1 U28748 ( .A(n43691), .B(n4568), .ZN(n24537) );
  XNOR2_X1 U28749 ( .A(n42995), .B(n48597), .ZN(n23845) );
  XNOR2_X1 U28750 ( .A(n24537), .B(n23845), .ZN(n17931) );
  XNOR2_X1 U28751 ( .A(n17932), .B(n17931), .ZN(n35081) );
  XNOR2_X1 U28752 ( .A(n23370), .B(n43702), .ZN(n26385) );
  XOR2_X1 U28753 ( .A(n3336), .B(n42668), .Z(n17933) );
  XNOR2_X1 U28754 ( .A(n26385), .B(n17933), .ZN(n35798) );
  XNOR2_X1 U28755 ( .A(n35798), .B(n4909), .ZN(n17934) );
  XNOR2_X1 U28756 ( .A(n35081), .B(n17934), .ZN(n17935) );
  XNOR2_X1 U28757 ( .A(n17936), .B(n17935), .ZN(n17937) );
  XNOR2_X1 U28758 ( .A(n19250), .B(n17937), .ZN(n17941) );
  XNOR2_X1 U28759 ( .A(n17938), .B(n18790), .ZN(n17939) );
  XNOR2_X1 U28760 ( .A(n17939), .B(n2225), .ZN(n17940) );
  XNOR2_X1 U28761 ( .A(n17944), .B(n17943), .ZN(n17945) );
  INV_X1 U28762 ( .A(n21373), .ZN(n20802) );
  XNOR2_X1 U28763 ( .A(n17947), .B(n18690), .ZN(n17949) );
  XNOR2_X1 U28764 ( .A(n17948), .B(n17949), .ZN(n17957) );
  XNOR2_X1 U28765 ( .A(n17950), .B(n43586), .ZN(n41924) );
  XOR2_X1 U28766 ( .A(n4599), .B(n4733), .Z(n17951) );
  XNOR2_X1 U28767 ( .A(n25866), .B(n17951), .ZN(n17952) );
  XNOR2_X1 U28768 ( .A(n41924), .B(n17952), .ZN(n36928) );
  XNOR2_X1 U28769 ( .A(n1341), .B(n4502), .ZN(n43262) );
  XNOR2_X1 U28770 ( .A(n4803), .B(n4864), .ZN(n18686) );
  XNOR2_X1 U28771 ( .A(n43262), .B(n18686), .ZN(n33071) );
  XNOR2_X1 U28772 ( .A(n36928), .B(n33071), .ZN(n17953) );
  XNOR2_X1 U28773 ( .A(n17954), .B(n17953), .ZN(n17955) );
  XNOR2_X1 U28774 ( .A(n18697), .B(n17955), .ZN(n17956) );
  XNOR2_X1 U28775 ( .A(n17957), .B(n17956), .ZN(n17958) );
  XNOR2_X1 U28776 ( .A(n17959), .B(n17958), .ZN(n17964) );
  XNOR2_X1 U28777 ( .A(n17961), .B(n18696), .ZN(n17962) );
  NAND3_X1 U28778 ( .A1(n21388), .A2(n20375), .A3(n20795), .ZN(n21372) );
  INV_X1 U28779 ( .A(n20416), .ZN(n21396) );
  XNOR2_X1 U28780 ( .A(n23887), .B(n42258), .ZN(n23494) );
  XNOR2_X1 U28781 ( .A(n23494), .B(n42539), .ZN(n37257) );
  XNOR2_X1 U28782 ( .A(n37257), .B(n4824), .ZN(n41961) );
  XNOR2_X1 U28783 ( .A(n41961), .B(n4721), .ZN(n34495) );
  XNOR2_X1 U28784 ( .A(n17966), .B(n18714), .ZN(n17967) );
  XNOR2_X1 U28785 ( .A(n17969), .B(n4691), .ZN(n35036) );
  XOR2_X1 U28786 ( .A(n2230), .B(n45736), .Z(n17970) );
  XNOR2_X1 U28787 ( .A(n35036), .B(n17970), .ZN(n17971) );
  XNOR2_X1 U28788 ( .A(n17972), .B(n17971), .ZN(n17974) );
  XNOR2_X1 U28789 ( .A(n17974), .B(n17973), .ZN(n17975) );
  XNOR2_X1 U28790 ( .A(n17975), .B(n635), .ZN(n17977) );
  XNOR2_X1 U28791 ( .A(n17977), .B(n17976), .ZN(n17978) );
  AOI21_X1 U28792 ( .B1(n21372), .B2(n21396), .A(n21397), .ZN(n17980) );
  OR2_X1 U28794 ( .A1(n581), .A2(n21389), .ZN(n20371) );
  INV_X1 U28795 ( .A(n20371), .ZN(n17981) );
  NAND4_X1 U28796 ( .A1(n20416), .A2(n5923), .A3(n21397), .A4(n21369), .ZN(
        n17982) );
  NAND2_X1 U28797 ( .A1(n1860), .A2(n581), .ZN(n20792) );
  NAND2_X1 U28798 ( .A1(n21370), .A2(n20791), .ZN(n17983) );
  AND2_X1 U28799 ( .A1(n17983), .A2(n20373), .ZN(n17985) );
  OAI211_X1 U28800 ( .C1(n581), .C2(n20415), .A(n21377), .B(n20805), .ZN(
        n17984) );
  NAND2_X1 U28801 ( .A1(n22901), .A2(n22919), .ZN(n22349) );
  NOR2_X1 U28802 ( .A1(n22349), .A2(n22367), .ZN(n17987) );
  INV_X1 U28803 ( .A(n2174), .ZN(n22363) );
  AND2_X1 U28804 ( .A1(n2175), .A2(n22918), .ZN(n22170) );
  INV_X1 U28805 ( .A(n22908), .ZN(n22902) );
  NOR2_X1 U28806 ( .A1(n22918), .A2(n2175), .ZN(n22354) );
  INV_X1 U28807 ( .A(n22349), .ZN(n17991) );
  NAND2_X1 U28808 ( .A1(n22354), .A2(n17991), .ZN(n17992) );
  XNOR2_X1 U28809 ( .A(n24550), .B(n17993), .ZN(n40849) );
  XNOR2_X1 U28810 ( .A(n42920), .B(n4177), .ZN(n17994) );
  XNOR2_X1 U28811 ( .A(n17996), .B(n17995), .ZN(n18279) );
  INV_X1 U28812 ( .A(n20388), .ZN(n17998) );
  INV_X1 U28813 ( .A(n20387), .ZN(n20459) );
  OAI21_X1 U28814 ( .B1(n20459), .B2(n17998), .A(n20477), .ZN(n18001) );
  NAND2_X1 U28815 ( .A1(n17999), .A2(n17639), .ZN(n18003) );
  INV_X1 U28816 ( .A(n18002), .ZN(n19372) );
  NAND3_X1 U28817 ( .A1(n18003), .A2(n20397), .A3(n19372), .ZN(n18004) );
  AOI22_X1 U28818 ( .A1(n19392), .A2(n18008), .B1(n18007), .B2(n18013), .ZN(
        n18020) );
  NAND2_X1 U28819 ( .A1(n3714), .A2(n18009), .ZN(n19390) );
  OAI211_X1 U28820 ( .C1(n19387), .C2(n18013), .A(n18012), .B(n18011), .ZN(
        n18019) );
  NOR2_X1 U28821 ( .A1(n18015), .A2(n3865), .ZN(n18016) );
  OAI21_X1 U28822 ( .B1(n18017), .B2(n18016), .A(n19395), .ZN(n18018) );
  OAI211_X1 U28823 ( .C1(n18020), .C2(n19390), .A(n18019), .B(n18018), .ZN(
        n18030) );
  INV_X1 U28824 ( .A(n18022), .ZN(n19400) );
  NAND3_X1 U28825 ( .A1(n18025), .A2(n18023), .A3(n18024), .ZN(n18026) );
  NAND4_X1 U28826 ( .A1(n19402), .A2(n18028), .A3(n18027), .A4(n18026), .ZN(
        n18029) );
  NAND2_X1 U28827 ( .A1(n18031), .A2(n19425), .ZN(n18038) );
  AND2_X1 U28828 ( .A1(n18034), .A2(n18033), .ZN(n18035) );
  AOI22_X1 U28829 ( .A1(n18038), .A2(n18037), .B1(n18036), .B2(n18035), .ZN(
        n18049) );
  NOR2_X1 U28830 ( .A1(n51374), .A2(n18039), .ZN(n18042) );
  AOI22_X1 U28831 ( .A1(n19404), .A2(n18042), .B1(n18041), .B2(n18040), .ZN(
        n18045) );
  OAI211_X1 U28832 ( .C1(n18047), .C2(n18046), .A(n18045), .B(n18044), .ZN(
        n18048) );
  NAND3_X1 U28833 ( .A1(n20436), .A2(n40), .A3(n20363), .ZN(n20356) );
  INV_X1 U28834 ( .A(n20357), .ZN(n19332) );
  AOI21_X1 U28835 ( .B1(n20356), .B2(n18050), .A(n20360), .ZN(n18056) );
  NAND2_X1 U28836 ( .A1(n20349), .A2(n20359), .ZN(n18054) );
  AOI21_X1 U28837 ( .B1(n18054), .B2(n18053), .A(n18052), .ZN(n18055) );
  NOR2_X1 U28838 ( .A1(n20348), .A2(n20359), .ZN(n20425) );
  NAND2_X1 U28839 ( .A1(n20347), .A2(n20428), .ZN(n20345) );
  AOI22_X1 U28840 ( .A1(n18064), .A2(n18063), .B1(n18062), .B2(n772), .ZN(
        n18068) );
  INV_X1 U28841 ( .A(n18065), .ZN(n18067) );
  OAI21_X1 U28842 ( .B1(n18068), .B2(n18067), .A(n18066), .ZN(n18069) );
  OAI21_X1 U28843 ( .B1(n18072), .B2(n18342), .A(n18341), .ZN(n18073) );
  OAI21_X1 U28844 ( .B1(n22186), .B2(n22190), .A(n20564), .ZN(n18095) );
  AOI21_X1 U28845 ( .B1(n20561), .B2(n21712), .A(n21106), .ZN(n18094) );
  MUX2_X1 U28846 ( .A(n20512), .B(n18081), .S(n18085), .Z(n18078) );
  INV_X1 U28847 ( .A(n18075), .ZN(n19341) );
  OAI211_X1 U28848 ( .C1(n18078), .C2(n19341), .A(n18077), .B(n18076), .ZN(
        n18079) );
  INV_X1 U28849 ( .A(n18079), .ZN(n18093) );
  NOR2_X1 U28850 ( .A1(n18080), .A2(n19344), .ZN(n19343) );
  AND2_X1 U28851 ( .A1(n20507), .A2(n18081), .ZN(n18084) );
  NOR2_X1 U28852 ( .A1(n18082), .A2(n20503), .ZN(n18083) );
  AOI22_X1 U28853 ( .A1(n19343), .A2(n489), .B1(n18084), .B2(n18083), .ZN(
        n18092) );
  OAI211_X1 U28854 ( .C1(n18087), .C2(n18086), .A(n18085), .B(n17619), .ZN(
        n18091) );
  NAND2_X1 U28855 ( .A1(n20508), .A2(n18088), .ZN(n20517) );
  INV_X1 U28856 ( .A(n20517), .ZN(n18089) );
  AND2_X1 U28857 ( .A1(n51705), .A2(n19344), .ZN(n19339) );
  OAI211_X1 U28858 ( .C1(n18089), .C2(n19339), .A(n20504), .B(n20512), .ZN(
        n18090) );
  NAND4_X2 U28859 ( .A1(n18092), .A2(n18093), .A3(n18090), .A4(n18091), .ZN(
        n21714) );
  OAI21_X1 U28860 ( .B1(n18095), .B2(n18094), .A(n21713), .ZN(n18099) );
  NAND2_X1 U28861 ( .A1(n21713), .A2(n22176), .ZN(n21104) );
  NAND2_X1 U28862 ( .A1(n463), .A2(n21105), .ZN(n21716) );
  OAI21_X1 U28863 ( .B1(n19916), .B2(n21104), .A(n21716), .ZN(n18096) );
  INV_X1 U28864 ( .A(n18096), .ZN(n18098) );
  OAI21_X1 U28866 ( .B1(n22191), .B2(n22189), .A(n21717), .ZN(n18097) );
  AND2_X1 U28867 ( .A1(n1597), .A2(n498), .ZN(n18872) );
  INV_X1 U28868 ( .A(n18101), .ZN(n18862) );
  NAND2_X1 U28869 ( .A1(n18863), .A2(n20682), .ZN(n18103) );
  INV_X1 U28870 ( .A(n20231), .ZN(n18105) );
  NAND2_X1 U28871 ( .A1(n21200), .A2(n6078), .ZN(n19008) );
  INV_X1 U28872 ( .A(n19008), .ZN(n18106) );
  NAND4_X1 U28873 ( .A1(n18106), .A2(n19820), .A3(n19819), .A4(n21197), .ZN(
        n21205) );
  NAND3_X1 U28874 ( .A1(n18106), .A2(n19822), .A3(n21197), .ZN(n18107) );
  NAND3_X1 U28875 ( .A1(n21205), .A2(n21196), .A3(n18107), .ZN(n18110) );
  INV_X1 U28876 ( .A(n18108), .ZN(n18109) );
  NAND2_X1 U28877 ( .A1(n18110), .A2(n18109), .ZN(n18116) );
  NAND2_X1 U28878 ( .A1(n19820), .A2(n2229), .ZN(n21194) );
  OR2_X1 U28879 ( .A1(n21194), .A2(n21213), .ZN(n19726) );
  INV_X1 U28880 ( .A(n19726), .ZN(n18111) );
  OAI21_X1 U28881 ( .B1(n18112), .B2(n18111), .A(n19734), .ZN(n18115) );
  NAND2_X1 U28882 ( .A1(n6078), .A2(n19007), .ZN(n21201) );
  OR2_X1 U28883 ( .A1(n21215), .A2(n21201), .ZN(n19807) );
  NOR2_X1 U28884 ( .A1(n21215), .A2(n19725), .ZN(n21209) );
  INV_X1 U28885 ( .A(n21199), .ZN(n19012) );
  OAI21_X1 U28886 ( .B1(n21209), .B2(n19012), .A(n2456), .ZN(n18113) );
  XNOR2_X1 U28887 ( .A(n18483), .B(n18475), .ZN(n18121) );
  XNOR2_X1 U28888 ( .A(n18117), .B(n4654), .ZN(n27433) );
  XNOR2_X1 U28889 ( .A(n27433), .B(n18118), .ZN(n28729) );
  XNOR2_X1 U28890 ( .A(n18121), .B(n18120), .ZN(n18122) );
  INV_X1 U28891 ( .A(n18124), .ZN(n18125) );
  XNOR2_X1 U28892 ( .A(n18125), .B(n4827), .ZN(n43316) );
  XNOR2_X1 U28893 ( .A(n43316), .B(n6031), .ZN(n37060) );
  XNOR2_X1 U28894 ( .A(n18126), .B(n37060), .ZN(n18128) );
  XNOR2_X1 U28895 ( .A(n18128), .B(n18127), .ZN(n18129) );
  INV_X1 U28896 ( .A(n19796), .ZN(n18997) );
  XNOR2_X1 U28897 ( .A(n18131), .B(n4916), .ZN(n27318) );
  XNOR2_X1 U28898 ( .A(n27318), .B(n44495), .ZN(n34124) );
  XNOR2_X1 U28899 ( .A(n28071), .B(n4869), .ZN(n42460) );
  XNOR2_X1 U28900 ( .A(n42460), .B(n4926), .ZN(n18132) );
  XNOR2_X1 U28901 ( .A(n34124), .B(n18132), .ZN(n18133) );
  XNOR2_X1 U28902 ( .A(n18134), .B(n18133), .ZN(n18136) );
  XNOR2_X1 U28903 ( .A(n18135), .B(n18136), .ZN(n18137) );
  XNOR2_X1 U28904 ( .A(n18138), .B(n18137), .ZN(n18140) );
  XNOR2_X1 U28905 ( .A(n18139), .B(n18140), .ZN(n18144) );
  XNOR2_X1 U28906 ( .A(n18142), .B(n18141), .ZN(n18143) );
  XNOR2_X1 U28907 ( .A(n18144), .B(n18143), .ZN(n18145) );
  XNOR2_X1 U28908 ( .A(n18147), .B(n18409), .ZN(n18149) );
  XNOR2_X1 U28909 ( .A(n637), .B(n18153), .ZN(n18159) );
  XNOR2_X1 U28910 ( .A(n34255), .B(n45883), .ZN(n42824) );
  XNOR2_X1 U28911 ( .A(n42101), .B(n18154), .ZN(n37009) );
  XNOR2_X1 U28912 ( .A(n37009), .B(n4666), .ZN(n18155) );
  XNOR2_X1 U28913 ( .A(n42824), .B(n18155), .ZN(n18156) );
  XNOR2_X1 U28914 ( .A(n18157), .B(n18156), .ZN(n18158) );
  XNOR2_X1 U28915 ( .A(n18159), .B(n18158), .ZN(n18160) );
  XNOR2_X1 U28916 ( .A(n18160), .B(n18161), .ZN(n18165) );
  XNOR2_X1 U28917 ( .A(n18163), .B(n52190), .ZN(n18164) );
  XNOR2_X1 U28918 ( .A(n18165), .B(n18164), .ZN(n18166) );
  XNOR2_X1 U28919 ( .A(n18539), .B(n51758), .ZN(n18170) );
  XNOR2_X1 U28920 ( .A(n18169), .B(n18170), .ZN(n18179) );
  XNOR2_X1 U28921 ( .A(n25795), .B(n4665), .ZN(n25578) );
  XNOR2_X1 U28922 ( .A(n18171), .B(n25578), .ZN(n29661) );
  XNOR2_X1 U28923 ( .A(n29661), .B(n4659), .ZN(n43057) );
  XNOR2_X1 U28924 ( .A(n33653), .B(n4454), .ZN(n25722) );
  XNOR2_X1 U28925 ( .A(n18172), .B(n4651), .ZN(n24896) );
  XNOR2_X1 U28926 ( .A(n25722), .B(n24896), .ZN(n37122) );
  XNOR2_X1 U28927 ( .A(n37122), .B(n29662), .ZN(n18173) );
  XNOR2_X1 U28928 ( .A(n43057), .B(n18173), .ZN(n18174) );
  XNOR2_X1 U28929 ( .A(n18175), .B(n18174), .ZN(n18177) );
  XNOR2_X1 U28930 ( .A(n18177), .B(n18176), .ZN(n18178) );
  XNOR2_X1 U28931 ( .A(n18179), .B(n18178), .ZN(n18183) );
  XNOR2_X1 U28932 ( .A(n18181), .B(n18180), .ZN(n18182) );
  XNOR2_X1 U28933 ( .A(n18183), .B(n18182), .ZN(n18184) );
  INV_X1 U28934 ( .A(n21304), .ZN(n19806) );
  XNOR2_X1 U28935 ( .A(n18633), .B(n18186), .ZN(n18201) );
  XNOR2_X1 U28936 ( .A(n2602), .B(n49937), .ZN(n34028) );
  XNOR2_X1 U28937 ( .A(n4649), .B(n4286), .ZN(n18187) );
  XNOR2_X1 U28938 ( .A(n2603), .B(n18187), .ZN(n18188) );
  XNOR2_X1 U28939 ( .A(n34028), .B(n18188), .ZN(n18189) );
  XNOR2_X1 U28940 ( .A(n18190), .B(n18189), .ZN(n33362) );
  XNOR2_X1 U28941 ( .A(n18191), .B(n24553), .ZN(n34096) );
  XNOR2_X1 U28942 ( .A(n33362), .B(n34096), .ZN(n18192) );
  XNOR2_X1 U28943 ( .A(n18193), .B(n18192), .ZN(n18195) );
  XNOR2_X1 U28944 ( .A(n18194), .B(n18195), .ZN(n18197) );
  XNOR2_X1 U28945 ( .A(n51133), .B(n18197), .ZN(n18199) );
  XNOR2_X1 U28946 ( .A(n18199), .B(n18198), .ZN(n18200) );
  XNOR2_X1 U28947 ( .A(n16532), .B(n18202), .ZN(n18203) );
  XNOR2_X1 U28948 ( .A(n18579), .B(n18203), .ZN(n18211) );
  XNOR2_X1 U28949 ( .A(n19768), .B(n42342), .ZN(n18205) );
  XNOR2_X1 U28950 ( .A(n23370), .B(n4353), .ZN(n18793) );
  XNOR2_X1 U28951 ( .A(n2183), .B(n4800), .ZN(n41272) );
  XNOR2_X1 U28952 ( .A(n18793), .B(n41272), .ZN(n18204) );
  XNOR2_X1 U28953 ( .A(n18205), .B(n18204), .ZN(n33520) );
  XNOR2_X1 U28954 ( .A(n18206), .B(n4558), .ZN(n27390) );
  XNOR2_X1 U28955 ( .A(n27390), .B(n35796), .ZN(n34439) );
  XNOR2_X1 U28956 ( .A(n33520), .B(n34439), .ZN(n18207) );
  XNOR2_X1 U28957 ( .A(n18209), .B(n18208), .ZN(n18210) );
  XNOR2_X1 U28958 ( .A(n18211), .B(n18210), .ZN(n18214) );
  XNOR2_X1 U28959 ( .A(n2226), .B(n18212), .ZN(n18213) );
  XNOR2_X1 U28960 ( .A(n18214), .B(n18213), .ZN(n18215) );
  NAND2_X1 U28961 ( .A1(n18888), .A2(n3683), .ZN(n18985) );
  OAI22_X1 U28962 ( .A1(n18996), .A2(n21305), .B1(n18985), .B2(n18999), .ZN(
        n18221) );
  INV_X1 U28963 ( .A(n18999), .ZN(n18882) );
  NAND3_X1 U28964 ( .A1(n18882), .A2(n18888), .A3(n509), .ZN(n18218) );
  OAI211_X1 U28965 ( .C1(n18995), .C2(n19792), .A(n18219), .B(n18218), .ZN(
        n18220) );
  AOI21_X1 U28966 ( .B1(n19794), .B2(n18221), .A(n18220), .ZN(n18226) );
  NOR2_X1 U28967 ( .A1(n18222), .A2(n18996), .ZN(n18224) );
  NAND2_X1 U28968 ( .A1(n18217), .A2(n19711), .ZN(n18223) );
  NAND2_X1 U28969 ( .A1(n20221), .A2(n20209), .ZN(n18918) );
  NAND2_X1 U28970 ( .A1(n19685), .A2(n19680), .ZN(n18227) );
  NOR2_X1 U28971 ( .A1(n18227), .A2(n20210), .ZN(n20222) );
  INV_X1 U28972 ( .A(n20222), .ZN(n18228) );
  NOR2_X1 U28973 ( .A1(n20210), .A2(n51006), .ZN(n18916) );
  OAI21_X1 U28974 ( .B1(n19687), .B2(n19680), .A(n20215), .ZN(n18229) );
  INV_X1 U28975 ( .A(n20207), .ZN(n19691) );
  NAND2_X1 U28976 ( .A1(n18229), .A2(n19691), .ZN(n18230) );
  OAI21_X1 U28977 ( .B1(n2118), .B2(n19689), .A(n18230), .ZN(n18231) );
  NAND2_X1 U28978 ( .A1(n18231), .A2(n19685), .ZN(n18241) );
  NOR2_X1 U28979 ( .A1(n18232), .A2(n775), .ZN(n18233) );
  AOI22_X1 U28980 ( .A1(n18233), .A2(n18234), .B1(n20217), .B2(n19688), .ZN(
        n18237) );
  INV_X1 U28981 ( .A(n20220), .ZN(n18236) );
  NAND2_X1 U28982 ( .A1(n18236), .A2(n8707), .ZN(n18235) );
  NAND3_X1 U28983 ( .A1(n20220), .A2(n19687), .A3(n19671), .ZN(n20208) );
  NAND3_X1 U28984 ( .A1(n20217), .A2(n19689), .A3(n19675), .ZN(n18238) );
  NAND3_X1 U28985 ( .A1(n19898), .A2(n18933), .A3(n19892), .ZN(n18250) );
  INV_X1 U28986 ( .A(n18932), .ZN(n19885) );
  AND2_X1 U28987 ( .A1(n18942), .A2(n19662), .ZN(n19632) );
  INV_X1 U28988 ( .A(n19887), .ZN(n18244) );
  INV_X1 U28989 ( .A(n19664), .ZN(n18243) );
  OAI22_X1 U28990 ( .A1(n18244), .A2(n18243), .B1(n19894), .B2(n19893), .ZN(
        n18245) );
  AOI22_X1 U28991 ( .A1(n51127), .A2(n19885), .B1(n19896), .B2(n18246), .ZN(
        n18249) );
  NOR2_X1 U28992 ( .A1(n18942), .A2(n19662), .ZN(n18247) );
  NAND4_X1 U28993 ( .A1(n19884), .A2(n18247), .A3(n18944), .A4(n19893), .ZN(
        n18248) );
  OR2_X1 U28994 ( .A1(n22837), .A2(n22492), .ZN(n20289) );
  OAI211_X1 U28995 ( .C1(n22834), .C2(n22822), .A(n21066), .B(n20289), .ZN(
        n18271) );
  NOR2_X1 U28996 ( .A1(n19870), .A2(n19865), .ZN(n19849) );
  INV_X1 U28997 ( .A(n19849), .ZN(n18252) );
  NAND3_X1 U28998 ( .A1(n19848), .A2(n19640), .A3(n374), .ZN(n18251) );
  AND2_X1 U28999 ( .A1(n18251), .A2(n18252), .ZN(n18260) );
  INV_X1 U29000 ( .A(n18253), .ZN(n18256) );
  INV_X1 U29001 ( .A(n18254), .ZN(n18255) );
  AND2_X1 U29002 ( .A1(n18256), .A2(n18255), .ZN(n18259) );
  NAND2_X1 U29003 ( .A1(n18910), .A2(n19863), .ZN(n18258) );
  NAND3_X1 U29004 ( .A1(n19650), .A2(n19869), .A3(n19848), .ZN(n18257) );
  NAND4_X1 U29005 ( .A1(n18260), .A2(n18259), .A3(n18258), .A4(n18257), .ZN(
        n18270) );
  NOR2_X1 U29006 ( .A1(n19866), .A2(n19851), .ZN(n18263) );
  INV_X1 U29007 ( .A(n585), .ZN(n19645) );
  OAI211_X1 U29008 ( .C1(n19853), .C2(n18263), .A(n51039), .B(n19645), .ZN(
        n18267) );
  NAND2_X1 U29009 ( .A1(n19639), .A2(n19033), .ZN(n19857) );
  INV_X1 U29010 ( .A(n19857), .ZN(n18264) );
  NAND2_X1 U29011 ( .A1(n18264), .A2(n51039), .ZN(n18266) );
  INV_X1 U29012 ( .A(n19867), .ZN(n19861) );
  INV_X1 U29013 ( .A(n19640), .ZN(n19852) );
  NAND3_X1 U29014 ( .A1(n19861), .A2(n19852), .A3(n19647), .ZN(n18265) );
  NAND4_X1 U29015 ( .A1(n18268), .A2(n18267), .A3(n18266), .A4(n18265), .ZN(
        n18269) );
  NAND2_X1 U29016 ( .A1(n18271), .A2(n22831), .ZN(n18278) );
  NAND2_X1 U29017 ( .A1(n22494), .A2(n22832), .ZN(n18272) );
  NOR2_X1 U29018 ( .A1(n22832), .A2(n22492), .ZN(n21068) );
  AOI21_X1 U29019 ( .B1(n21073), .B2(n18272), .A(n21068), .ZN(n18277) );
  NAND4_X1 U29021 ( .A1(n22832), .A2(n22834), .A3(n22830), .A4(n22826), .ZN(
        n18273) );
  OAI21_X1 U29022 ( .B1(n22504), .B2(n20297), .A(n18273), .ZN(n18274) );
  INV_X1 U29023 ( .A(n18274), .ZN(n18276) );
  INV_X1 U29024 ( .A(n21066), .ZN(n18275) );
  NAND2_X1 U29025 ( .A1(n18275), .A2(n22491), .ZN(n20293) );
  XNOR2_X1 U29026 ( .A(n25161), .B(n26119), .ZN(n25387) );
  XNOR2_X1 U29027 ( .A(n18279), .B(n25387), .ZN(n18280) );
  XNOR2_X1 U29028 ( .A(n18281), .B(n18280), .ZN(n19441) );
  NAND2_X1 U29029 ( .A1(n18282), .A2(n16798), .ZN(n18284) );
  AOI21_X1 U29030 ( .B1(n18285), .B2(n18284), .A(n18283), .ZN(n18298) );
  INV_X1 U29031 ( .A(n18286), .ZN(n18290) );
  NAND3_X1 U29032 ( .A1(n18288), .A2(n18287), .A3(n20021), .ZN(n18289) );
  OAI211_X1 U29033 ( .C1(n18290), .C2(n6952), .A(n20025), .B(n18289), .ZN(
        n18297) );
  OR2_X1 U29034 ( .A1(n18292), .A2(n18291), .ZN(n18296) );
  AOI22_X1 U29035 ( .A1(n20015), .A2(n18294), .B1(n51209), .B2(n2166), .ZN(
        n18295) );
  INV_X1 U29036 ( .A(n22121), .ZN(n21725) );
  AOI21_X1 U29037 ( .B1(n18304), .B2(n19491), .A(n19132), .ZN(n20079) );
  INV_X1 U29038 ( .A(n19500), .ZN(n18299) );
  AND2_X1 U29039 ( .A1(n19487), .A2(n20067), .ZN(n18306) );
  NOR2_X1 U29040 ( .A1(n18300), .A2(n20071), .ZN(n18301) );
  AOI22_X1 U29041 ( .A1(n18306), .A2(n18301), .B1(n20056), .B2(n20061), .ZN(
        n18309) );
  AOI21_X1 U29042 ( .B1(n20062), .B2(n2101), .A(n20067), .ZN(n18302) );
  OAI21_X1 U29043 ( .B1(n18304), .B2(n18303), .A(n18302), .ZN(n18308) );
  OAI21_X1 U29044 ( .B1(n20082), .B2(n20062), .A(n16218), .ZN(n18305) );
  AOI21_X1 U29045 ( .B1(n18306), .B2(n18305), .A(n20075), .ZN(n18307) );
  INV_X1 U29047 ( .A(n23213), .ZN(n23211) );
  NAND2_X1 U29048 ( .A1(n20105), .A2(n20086), .ZN(n18311) );
  NAND2_X1 U29049 ( .A1(n20093), .A2(n20097), .ZN(n18310) );
  OAI211_X1 U29050 ( .C1(n18312), .C2(n16788), .A(n18311), .B(n18310), .ZN(
        n18314) );
  NAND4_X1 U29051 ( .A1(n16787), .A2(n20100), .A3(n7131), .A4(n20104), .ZN(
        n18321) );
  NAND3_X1 U29052 ( .A1(n18318), .A2(n20092), .A3(n20090), .ZN(n18319) );
  NOR2_X1 U29053 ( .A1(n20097), .A2(n20087), .ZN(n18324) );
  AND2_X1 U29054 ( .A1(n18328), .A2(n18329), .ZN(n18335) );
  NAND4_X1 U29056 ( .A1(n18341), .A2(n18340), .A3(n18339), .A4(n18338), .ZN(
        n18343) );
  AND2_X1 U29057 ( .A1(n18343), .A2(n18342), .ZN(n20966) );
  NOR2_X1 U29059 ( .A1(n20137), .A2(n19064), .ZN(n18351) );
  OR2_X1 U29060 ( .A1(n20144), .A2(n51756), .ZN(n18347) );
  NAND3_X1 U29061 ( .A1(n18349), .A2(n18348), .A3(n18347), .ZN(n18350) );
  AOI21_X1 U29062 ( .B1(n18351), .B2(n20139), .A(n18350), .ZN(n18368) );
  NAND3_X1 U29063 ( .A1(n18352), .A2(n574), .A3(n51403), .ZN(n18353) );
  OAI211_X1 U29064 ( .C1(n19078), .C2(n19071), .A(n18354), .B(n18353), .ZN(
        n18355) );
  NAND3_X1 U29068 ( .A1(n19076), .A2(n19077), .A3(n18362), .ZN(n18363) );
  OAI21_X1 U29069 ( .B1(n19078), .B2(n19076), .A(n18363), .ZN(n18364) );
  NAND2_X1 U29070 ( .A1(n18364), .A2(n19075), .ZN(n18365) );
  NOR2_X1 U29071 ( .A1(n51355), .A2(n23219), .ZN(n18370) );
  OAI21_X1 U29072 ( .B1(n18371), .B2(n18370), .A(n20304), .ZN(n18372) );
  MUX2_X1 U29073 ( .A(n20046), .B(n51440), .S(n18377), .Z(n18379) );
  NAND2_X1 U29074 ( .A1(n18375), .A2(n20044), .ZN(n18378) );
  NAND2_X1 U29075 ( .A1(n18377), .A2(n18376), .ZN(n20035) );
  NAND2_X1 U29076 ( .A1(n18381), .A2(n6711), .ZN(n18382) );
  INV_X1 U29077 ( .A(n18387), .ZN(n18385) );
  NAND2_X1 U29078 ( .A1(n18387), .A2(n23219), .ZN(n23217) );
  NAND2_X1 U29079 ( .A1(n23207), .A2(n417), .ZN(n22115) );
  OAI21_X1 U29080 ( .B1(n18369), .B2(n22116), .A(n22115), .ZN(n18388) );
  INV_X1 U29081 ( .A(n23229), .ZN(n23218) );
  NAND2_X1 U29082 ( .A1(n23218), .A2(n22121), .ZN(n22119) );
  INV_X1 U29083 ( .A(n22119), .ZN(n21726) );
  XNOR2_X1 U29084 ( .A(n18528), .B(n18390), .ZN(n24581) );
  XNOR2_X1 U29085 ( .A(n24581), .B(n29662), .ZN(n33315) );
  XNOR2_X1 U29086 ( .A(n28267), .B(n24430), .ZN(n34154) );
  XNOR2_X1 U29087 ( .A(n34154), .B(n4415), .ZN(n18391) );
  XNOR2_X1 U29088 ( .A(n33315), .B(n18391), .ZN(n18392) );
  XNOR2_X1 U29089 ( .A(n461), .B(n18392), .ZN(n18396) );
  XNOR2_X1 U29090 ( .A(n2162), .B(n18658), .ZN(n18393) );
  XNOR2_X1 U29091 ( .A(n16201), .B(n18399), .ZN(n18406) );
  XNOR2_X1 U29092 ( .A(n35107), .B(n4213), .ZN(n33296) );
  XNOR2_X1 U29093 ( .A(n39719), .B(n33296), .ZN(n45310) );
  XNOR2_X1 U29094 ( .A(n33429), .B(n4587), .ZN(n26359) );
  XNOR2_X1 U29095 ( .A(n4554), .B(n4637), .ZN(n34508) );
  XNOR2_X1 U29096 ( .A(n26359), .B(n34508), .ZN(n18400) );
  XNOR2_X1 U29097 ( .A(n18401), .B(n18400), .ZN(n18402) );
  XNOR2_X1 U29098 ( .A(n45310), .B(n18402), .ZN(n18403) );
  XNOR2_X1 U29099 ( .A(n51436), .B(n18403), .ZN(n18405) );
  XNOR2_X1 U29100 ( .A(n18406), .B(n18405), .ZN(n18413) );
  XNOR2_X1 U29101 ( .A(n18408), .B(n18407), .ZN(n18411) );
  XNOR2_X1 U29102 ( .A(n19196), .B(n18409), .ZN(n18410) );
  XNOR2_X1 U29103 ( .A(n18411), .B(n18410), .ZN(n18412) );
  XNOR2_X1 U29104 ( .A(n18412), .B(n18413), .ZN(n18416) );
  XNOR2_X1 U29105 ( .A(n19198), .B(n18414), .ZN(n18415) );
  XNOR2_X1 U29106 ( .A(n18416), .B(n18415), .ZN(n18417) );
  XNOR2_X1 U29107 ( .A(n18418), .B(n18419), .ZN(n18421) );
  XNOR2_X1 U29108 ( .A(n4353), .B(n4295), .ZN(n23846) );
  XNOR2_X1 U29109 ( .A(n18422), .B(n23846), .ZN(n36979) );
  XNOR2_X1 U29110 ( .A(n25148), .B(n18423), .ZN(n43692) );
  XNOR2_X1 U29111 ( .A(n4624), .B(n4076), .ZN(n25641) );
  XNOR2_X1 U29112 ( .A(n43692), .B(n25641), .ZN(n33105) );
  XNOR2_X1 U29113 ( .A(n33105), .B(n34575), .ZN(n18424) );
  XNOR2_X1 U29114 ( .A(n36979), .B(n18424), .ZN(n18425) );
  XNOR2_X1 U29115 ( .A(n18426), .B(n18790), .ZN(n18428) );
  XNOR2_X1 U29116 ( .A(n18428), .B(n18798), .ZN(n18429) );
  XNOR2_X1 U29117 ( .A(n51135), .B(n18432), .ZN(n18433) );
  XNOR2_X1 U29118 ( .A(n18433), .B(n2200), .ZN(n18434) );
  XNOR2_X1 U29119 ( .A(n2217), .B(n18434), .ZN(n19240) );
  INV_X1 U29120 ( .A(n19240), .ZN(n18435) );
  XNOR2_X1 U29121 ( .A(n18435), .B(n18436), .ZN(n18454) );
  XNOR2_X1 U29122 ( .A(n18437), .B(n18438), .ZN(n18445) );
  XNOR2_X1 U29123 ( .A(n32267), .B(n4874), .ZN(n18439) );
  XNOR2_X1 U29124 ( .A(n24550), .B(n18439), .ZN(n37102) );
  XNOR2_X1 U29125 ( .A(n24315), .B(n18440), .ZN(n30525) );
  XNOR2_X1 U29126 ( .A(n34265), .B(n4826), .ZN(n37103) );
  XNOR2_X1 U29127 ( .A(n30525), .B(n37103), .ZN(n18441) );
  XNOR2_X1 U29128 ( .A(n37102), .B(n18441), .ZN(n18442) );
  XNOR2_X1 U29129 ( .A(n18443), .B(n18442), .ZN(n18444) );
  XNOR2_X1 U29130 ( .A(n18448), .B(n18447), .ZN(n18818) );
  INV_X1 U29131 ( .A(n18818), .ZN(n18449) );
  XNOR2_X1 U29132 ( .A(n18450), .B(n18449), .ZN(n18451) );
  XNOR2_X1 U29133 ( .A(n18452), .B(n18451), .ZN(n18453) );
  INV_X1 U29134 ( .A(n20624), .ZN(n20742) );
  XNOR2_X1 U29135 ( .A(n18712), .B(n4865), .ZN(n18456) );
  XNOR2_X1 U29136 ( .A(n18457), .B(n18456), .ZN(n18742) );
  XNOR2_X1 U29137 ( .A(n18750), .B(n635), .ZN(n18470) );
  XNOR2_X1 U29138 ( .A(n18460), .B(n18459), .ZN(n18468) );
  XNOR2_X1 U29139 ( .A(n27318), .B(n18461), .ZN(n42541) );
  XNOR2_X1 U29140 ( .A(n37042), .B(n2203), .ZN(n18462) );
  XNOR2_X1 U29141 ( .A(n42541), .B(n18462), .ZN(n18463) );
  XNOR2_X1 U29142 ( .A(n18464), .B(n18463), .ZN(n18465) );
  XNOR2_X1 U29143 ( .A(n18466), .B(n18465), .ZN(n18467) );
  XNOR2_X1 U29144 ( .A(n18468), .B(n18467), .ZN(n18469) );
  XNOR2_X1 U29145 ( .A(n33201), .B(n24992), .ZN(n45478) );
  XNOR2_X1 U29146 ( .A(n33474), .B(n4835), .ZN(n18702) );
  XNOR2_X1 U29147 ( .A(n18702), .B(n4599), .ZN(n44954) );
  XNOR2_X1 U29148 ( .A(n31431), .B(n4026), .ZN(n18473) );
  XNOR2_X1 U29149 ( .A(n44954), .B(n18473), .ZN(n33285) );
  XNOR2_X1 U29150 ( .A(n45478), .B(n33285), .ZN(n18474) );
  XNOR2_X1 U29151 ( .A(n18475), .B(n18474), .ZN(n18477) );
  XNOR2_X1 U29152 ( .A(n18477), .B(n18476), .ZN(n18478) );
  XNOR2_X1 U29153 ( .A(n18478), .B(n18828), .ZN(n18482) );
  XNOR2_X1 U29154 ( .A(n18479), .B(n51454), .ZN(n18481) );
  XNOR2_X1 U29155 ( .A(n18481), .B(n18482), .ZN(n18487) );
  XNOR2_X1 U29156 ( .A(n18831), .B(n18483), .ZN(n18484) );
  XNOR2_X1 U29157 ( .A(n18484), .B(n18832), .ZN(n18694) );
  XNOR2_X1 U29158 ( .A(n18694), .B(n18485), .ZN(n18486) );
  XNOR2_X1 U29159 ( .A(n18487), .B(n18486), .ZN(n18493) );
  INV_X1 U29160 ( .A(n18488), .ZN(n18491) );
  INV_X1 U29161 ( .A(n18489), .ZN(n18490) );
  XNOR2_X1 U29162 ( .A(n18491), .B(n18490), .ZN(n18492) );
  INV_X1 U29164 ( .A(n20642), .ZN(n20627) );
  INV_X1 U29165 ( .A(n21538), .ZN(n20751) );
  OAI21_X1 U29166 ( .B1(n20751), .B2(n18495), .A(n18494), .ZN(n18498) );
  INV_X1 U29168 ( .A(n21533), .ZN(n20749) );
  NAND2_X1 U29169 ( .A1(n18496), .A2(n20197), .ZN(n18497) );
  AND2_X1 U29170 ( .A1(n20745), .A2(n51485), .ZN(n20195) );
  NOR2_X1 U29171 ( .A1(n20745), .A2(n21543), .ZN(n18499) );
  OAI21_X1 U29173 ( .B1(n20195), .B2(n18499), .A(n21541), .ZN(n18502) );
  NOR2_X1 U29174 ( .A1(n20737), .A2(n21540), .ZN(n20625) );
  INV_X1 U29175 ( .A(n20625), .ZN(n18501) );
  NAND3_X1 U29176 ( .A1(n20752), .A2(n20736), .A3(n21544), .ZN(n18500) );
  XNOR2_X1 U29178 ( .A(n14903), .B(n18505), .ZN(n18506) );
  XNOR2_X1 U29180 ( .A(n4605), .B(n4451), .ZN(n18508) );
  XNOR2_X1 U29181 ( .A(n34411), .B(n18508), .ZN(n18511) );
  XNOR2_X1 U29182 ( .A(n4637), .B(n3367), .ZN(n18509) );
  XNOR2_X1 U29183 ( .A(n18509), .B(n4940), .ZN(n18510) );
  XNOR2_X1 U29184 ( .A(n18511), .B(n18510), .ZN(n25468) );
  INV_X1 U29185 ( .A(n33049), .ZN(n18512) );
  XNOR2_X1 U29186 ( .A(n18513), .B(n18512), .ZN(n18514) );
  XNOR2_X1 U29187 ( .A(n25468), .B(n18514), .ZN(n34165) );
  XNOR2_X1 U29188 ( .A(n33296), .B(n4431), .ZN(n18515) );
  XNOR2_X1 U29189 ( .A(n18515), .B(n33295), .ZN(n18516) );
  XNOR2_X1 U29190 ( .A(n34165), .B(n18516), .ZN(n18517) );
  XNOR2_X1 U29191 ( .A(n19199), .B(n18517), .ZN(n18518) );
  XNOR2_X1 U29192 ( .A(n18519), .B(n18518), .ZN(n18520) );
  XNOR2_X1 U29194 ( .A(n18524), .B(n2113), .ZN(n18675) );
  XNOR2_X1 U29195 ( .A(n4755), .B(n4659), .ZN(n19218) );
  XNOR2_X1 U29196 ( .A(n25042), .B(n19218), .ZN(n27228) );
  XNOR2_X1 U29197 ( .A(n18527), .B(n27228), .ZN(n33951) );
  XNOR2_X1 U29198 ( .A(n33951), .B(n26541), .ZN(n18529) );
  XNOR2_X1 U29199 ( .A(n18528), .B(n4542), .ZN(n34789) );
  XNOR2_X1 U29200 ( .A(n18529), .B(n34789), .ZN(n18530) );
  XNOR2_X1 U29201 ( .A(n2121), .B(n18530), .ZN(n18532) );
  XNOR2_X1 U29202 ( .A(n18533), .B(n18532), .ZN(n18536) );
  XNOR2_X1 U29203 ( .A(n462), .B(n52168), .ZN(n19228) );
  XNOR2_X1 U29204 ( .A(n19228), .B(n18536), .ZN(n18537) );
  XNOR2_X1 U29205 ( .A(n18537), .B(n18538), .ZN(n18545) );
  XNOR2_X1 U29206 ( .A(n18539), .B(n842), .ZN(n18541) );
  XNOR2_X1 U29207 ( .A(n18540), .B(n18541), .ZN(n18662) );
  XNOR2_X1 U29208 ( .A(n18662), .B(n19227), .ZN(n18542) );
  XNOR2_X1 U29209 ( .A(n18543), .B(n18542), .ZN(n18544) );
  INV_X1 U29211 ( .A(n19943), .ZN(n18563) );
  XNOR2_X1 U29212 ( .A(n18546), .B(n18818), .ZN(n18552) );
  XNOR2_X1 U29213 ( .A(n52227), .B(n51642), .ZN(n18549) );
  XNOR2_X1 U29214 ( .A(n18550), .B(n18549), .ZN(n18551) );
  XNOR2_X1 U29215 ( .A(n18552), .B(n18551), .ZN(n18554) );
  XNOR2_X1 U29216 ( .A(n18554), .B(n18553), .ZN(n18562) );
  XNOR2_X1 U29217 ( .A(n18555), .B(n34027), .ZN(n24458) );
  XNOR2_X1 U29218 ( .A(n24458), .B(n4287), .ZN(n42723) );
  XNOR2_X1 U29219 ( .A(n24314), .B(n35815), .ZN(n23397) );
  XNOR2_X1 U29220 ( .A(n42723), .B(n23397), .ZN(n35623) );
  XNOR2_X1 U29221 ( .A(n43850), .B(n4879), .ZN(n24459) );
  XNOR2_X1 U29222 ( .A(n24459), .B(n18556), .ZN(n35233) );
  XNOR2_X1 U29223 ( .A(n35623), .B(n35233), .ZN(n18557) );
  XNOR2_X1 U29224 ( .A(n18616), .B(n18557), .ZN(n18558) );
  XNOR2_X1 U29225 ( .A(n18617), .B(n18558), .ZN(n18560) );
  XNOR2_X1 U29226 ( .A(n18560), .B(n18559), .ZN(n18561) );
  XNOR2_X1 U29227 ( .A(n18564), .B(n18828), .ZN(n18567) );
  XNOR2_X1 U29228 ( .A(n18697), .B(n18565), .ZN(n18566) );
  XNOR2_X1 U29229 ( .A(n18567), .B(n18566), .ZN(n18569) );
  XNOR2_X1 U29230 ( .A(n18569), .B(n18568), .ZN(n18578) );
  XNOR2_X1 U29231 ( .A(n4204), .B(n4317), .ZN(n19182) );
  XNOR2_X1 U29232 ( .A(n18570), .B(n19182), .ZN(n34731) );
  XNOR2_X1 U29233 ( .A(n43074), .B(n24992), .ZN(n33915) );
  XNOR2_X1 U29234 ( .A(n34731), .B(n33915), .ZN(n18571) );
  XNOR2_X1 U29235 ( .A(n19185), .B(n18571), .ZN(n18572) );
  XNOR2_X1 U29236 ( .A(n18572), .B(n19186), .ZN(n18574) );
  XNOR2_X1 U29237 ( .A(n18574), .B(n18573), .ZN(n18576) );
  XNOR2_X1 U29238 ( .A(n18576), .B(n18575), .ZN(n18577) );
  XNOR2_X1 U29239 ( .A(n18580), .B(n18579), .ZN(n19253) );
  XNOR2_X1 U29240 ( .A(n19253), .B(n18581), .ZN(n18587) );
  XNOR2_X1 U29241 ( .A(n24818), .B(n33388), .ZN(n44220) );
  XNOR2_X1 U29242 ( .A(n37082), .B(n49429), .ZN(n26101) );
  XNOR2_X1 U29243 ( .A(n26101), .B(n4295), .ZN(n18583) );
  XNOR2_X1 U29244 ( .A(n44220), .B(n18583), .ZN(n18584) );
  XNOR2_X1 U29245 ( .A(n18798), .B(n18584), .ZN(n18585) );
  XNOR2_X1 U29246 ( .A(n18648), .B(n18585), .ZN(n18586) );
  XNOR2_X1 U29247 ( .A(n18587), .B(n18586), .ZN(n18588) );
  INV_X1 U29248 ( .A(n18610), .ZN(n20325) );
  NAND2_X1 U29249 ( .A1(n21420), .A2(n3493), .ZN(n18590) );
  AND2_X1 U29250 ( .A1(n20325), .A2(n52139), .ZN(n19162) );
  NAND3_X1 U29251 ( .A1(n21427), .A2(n3493), .A3(n52139), .ZN(n18607) );
  XNOR2_X1 U29252 ( .A(n18591), .B(n635), .ZN(n18595) );
  XNOR2_X1 U29253 ( .A(n24797), .B(n4908), .ZN(n35590) );
  XNOR2_X1 U29254 ( .A(n45463), .B(n4865), .ZN(n18596) );
  XNOR2_X1 U29255 ( .A(n35590), .B(n18596), .ZN(n18597) );
  XNOR2_X1 U29256 ( .A(n18597), .B(n35034), .ZN(n18598) );
  XNOR2_X1 U29257 ( .A(n18599), .B(n18598), .ZN(n18601) );
  XNOR2_X1 U29258 ( .A(n18602), .B(n18603), .ZN(n19266) );
  AOI22_X1 U29259 ( .A1(n19162), .A2(n21442), .B1(n18607), .B2(n21421), .ZN(
        n18609) );
  INV_X1 U29260 ( .A(n21420), .ZN(n21440) );
  NAND2_X1 U29261 ( .A1(n21440), .A2(n19947), .ZN(n18608) );
  NAND2_X1 U29262 ( .A1(n20840), .A2(n20322), .ZN(n21436) );
  NAND2_X1 U29263 ( .A1(n21436), .A2(n20329), .ZN(n18613) );
  NAND2_X1 U29264 ( .A1(n21427), .A2(n20326), .ZN(n21443) );
  INV_X1 U29265 ( .A(n21443), .ZN(n20839) );
  AND2_X1 U29266 ( .A1(n19947), .A2(n21425), .ZN(n21439) );
  OAI21_X1 U29267 ( .B1(n20836), .B2(n20839), .A(n21439), .ZN(n18612) );
  INV_X1 U29269 ( .A(n20327), .ZN(n21422) );
  NAND3_X1 U29270 ( .A1(n21422), .A2(n21426), .A3(n20322), .ZN(n18611) );
  NOR2_X1 U29272 ( .A1(n24186), .A2(n24187), .ZN(n23194) );
  XNOR2_X1 U29273 ( .A(n18615), .B(n18616), .ZN(n18618) );
  XNOR2_X1 U29274 ( .A(n18618), .B(n18617), .ZN(n18620) );
  XNOR2_X1 U29275 ( .A(n18620), .B(n18619), .ZN(n18632) );
  XNOR2_X1 U29276 ( .A(n27349), .B(n42025), .ZN(n18623) );
  XNOR2_X1 U29277 ( .A(n32856), .B(n4890), .ZN(n18621) );
  XNOR2_X1 U29278 ( .A(n18621), .B(n33374), .ZN(n18622) );
  XNOR2_X1 U29279 ( .A(n18623), .B(n18622), .ZN(n18625) );
  XNOR2_X1 U29280 ( .A(n28391), .B(n35816), .ZN(n18624) );
  XNOR2_X1 U29281 ( .A(n18625), .B(n18624), .ZN(n18626) );
  XNOR2_X1 U29282 ( .A(n19235), .B(n18626), .ZN(n18627) );
  XNOR2_X1 U29283 ( .A(n52209), .B(n18627), .ZN(n18629) );
  XNOR2_X1 U29284 ( .A(n18630), .B(n18629), .ZN(n18631) );
  INV_X1 U29285 ( .A(n18633), .ZN(n18634) );
  XNOR2_X1 U29286 ( .A(n18636), .B(n4909), .ZN(n25924) );
  XNOR2_X1 U29287 ( .A(n25924), .B(n18637), .ZN(n18639) );
  INV_X1 U29288 ( .A(n26385), .ZN(n18638) );
  XNOR2_X1 U29289 ( .A(n18639), .B(n18638), .ZN(n36697) );
  XNOR2_X1 U29290 ( .A(n27454), .B(n49323), .ZN(n31926) );
  XNOR2_X1 U29291 ( .A(n43293), .B(n49429), .ZN(n18640) );
  XNOR2_X1 U29292 ( .A(n31926), .B(n18640), .ZN(n18641) );
  XNOR2_X1 U29293 ( .A(n36697), .B(n18641), .ZN(n18642) );
  XNOR2_X1 U29294 ( .A(n18643), .B(n18642), .ZN(n18645) );
  XNOR2_X1 U29295 ( .A(n18644), .B(n18645), .ZN(n18647) );
  XNOR2_X1 U29296 ( .A(n18646), .B(n18647), .ZN(n18650) );
  XNOR2_X1 U29297 ( .A(n18648), .B(n18806), .ZN(n18649) );
  XOR2_X1 U29298 ( .A(n18650), .B(n18649), .Z(n18651) );
  INV_X1 U29299 ( .A(n20768), .ZN(n21600) );
  XNOR2_X1 U29300 ( .A(n25040), .B(n4542), .ZN(n18653) );
  XNOR2_X1 U29301 ( .A(n26370), .B(n18653), .ZN(n18655) );
  INV_X1 U29302 ( .A(n26296), .ZN(n18654) );
  XNOR2_X1 U29303 ( .A(n18655), .B(n18654), .ZN(n24827) );
  XNOR2_X1 U29304 ( .A(n18656), .B(n4651), .ZN(n34059) );
  XNOR2_X1 U29305 ( .A(n24827), .B(n34059), .ZN(n18657) );
  XNOR2_X1 U29306 ( .A(n18658), .B(n18657), .ZN(n18659) );
  XNOR2_X1 U29307 ( .A(n18661), .B(n18662), .ZN(n18663) );
  XNOR2_X1 U29308 ( .A(n18664), .B(n18663), .ZN(n18665) );
  XNOR2_X1 U29309 ( .A(n34414), .B(n4157), .ZN(n18666) );
  XNOR2_X1 U29310 ( .A(n44046), .B(n18666), .ZN(n18667) );
  XNOR2_X1 U29311 ( .A(n18668), .B(n18667), .ZN(n18670) );
  XNOR2_X1 U29312 ( .A(n18670), .B(n18669), .ZN(n18672) );
  XNOR2_X1 U29313 ( .A(n18671), .B(n18672), .ZN(n18674) );
  XNOR2_X1 U29314 ( .A(n18674), .B(n18673), .ZN(n18676) );
  XNOR2_X1 U29315 ( .A(n18676), .B(n18675), .ZN(n18683) );
  INV_X1 U29316 ( .A(n18677), .ZN(n18679) );
  XNOR2_X1 U29317 ( .A(n18679), .B(n18678), .ZN(n18680) );
  XNOR2_X1 U29318 ( .A(n18681), .B(n18680), .ZN(n18682) );
  NAND2_X1 U29319 ( .A1(n18685), .A2(n18684), .ZN(n18721) );
  NAND2_X1 U29320 ( .A1(n5150), .A2(n21355), .ZN(n19293) );
  OR2_X1 U29321 ( .A1(n19293), .A2(n21364), .ZN(n20765) );
  INV_X1 U29322 ( .A(n43265), .ZN(n26418) );
  XNOR2_X1 U29323 ( .A(n26418), .B(n18686), .ZN(n18687) );
  XNOR2_X1 U29324 ( .A(n23773), .B(n18687), .ZN(n34015) );
  XNOR2_X1 U29325 ( .A(n34015), .B(n4613), .ZN(n18688) );
  XNOR2_X1 U29326 ( .A(n18689), .B(n18688), .ZN(n18691) );
  XNOR2_X1 U29327 ( .A(n18690), .B(n18691), .ZN(n18693) );
  XNOR2_X1 U29328 ( .A(n18693), .B(n566), .ZN(n18695) );
  XNOR2_X1 U29329 ( .A(n18695), .B(n18694), .ZN(n18699) );
  XNOR2_X1 U29330 ( .A(n18697), .B(n18696), .ZN(n18698) );
  XNOR2_X1 U29331 ( .A(n15619), .B(n18701), .ZN(n19192) );
  XNOR2_X1 U29332 ( .A(n44952), .B(n4628), .ZN(n26419) );
  XNOR2_X1 U29333 ( .A(n26419), .B(n18702), .ZN(n33404) );
  XNOR2_X1 U29334 ( .A(n19192), .B(n33404), .ZN(n18824) );
  INV_X1 U29335 ( .A(n21351), .ZN(n21599) );
  XNOR2_X1 U29336 ( .A(n4895), .B(n4934), .ZN(n35831) );
  XNOR2_X1 U29337 ( .A(n19260), .B(n35831), .ZN(n18703) );
  XNOR2_X1 U29338 ( .A(n18704), .B(n18703), .ZN(n18752) );
  XNOR2_X1 U29339 ( .A(n18705), .B(n18752), .ZN(n18708) );
  INV_X1 U29340 ( .A(n18706), .ZN(n18707) );
  XNOR2_X1 U29341 ( .A(n18708), .B(n18707), .ZN(n18719) );
  INV_X1 U29342 ( .A(n18709), .ZN(n18717) );
  XNOR2_X1 U29343 ( .A(n35838), .B(n24928), .ZN(n18710) );
  XNOR2_X1 U29344 ( .A(n35036), .B(n18710), .ZN(n18711) );
  XNOR2_X1 U29345 ( .A(n18712), .B(n18711), .ZN(n18713) );
  XNOR2_X1 U29346 ( .A(n18715), .B(n18714), .ZN(n18716) );
  XNOR2_X1 U29347 ( .A(n18717), .B(n18716), .ZN(n18718) );
  INV_X1 U29348 ( .A(n18726), .ZN(n21601) );
  AND2_X1 U29349 ( .A1(n21601), .A2(n21599), .ZN(n19290) );
  NAND3_X1 U29350 ( .A1(n762), .A2(n21356), .A3(n20768), .ZN(n21609) );
  INV_X1 U29351 ( .A(n18724), .ZN(n19285) );
  NAND2_X1 U29352 ( .A1(n19284), .A2(n21354), .ZN(n21598) );
  OAI22_X1 U29353 ( .A1(n19293), .A2(n19285), .B1(n21598), .B2(n21604), .ZN(
        n18722) );
  OAI21_X1 U29354 ( .B1(n19286), .B2(n18722), .A(n21349), .ZN(n18723) );
  OR2_X1 U29355 ( .A1(n18724), .A2(n21601), .ZN(n20767) );
  NAND2_X1 U29356 ( .A1(n21356), .A2(n18724), .ZN(n18725) );
  MUX2_X1 U29357 ( .A(n20767), .B(n18725), .S(n19289), .Z(n18727) );
  BUF_X2 U29358 ( .A(n18726), .Z(n21362) );
  NAND2_X1 U29359 ( .A1(n21362), .A2(n19284), .ZN(n19927) );
  AND2_X1 U29360 ( .A1(n19284), .A2(n21351), .ZN(n20758) );
  NAND2_X1 U29361 ( .A1(n20696), .A2(n21620), .ZN(n21633) );
  OR2_X1 U29362 ( .A1(n21633), .A2(n21630), .ZN(n19977) );
  NAND2_X1 U29363 ( .A1(n21615), .A2(n21629), .ZN(n18730) );
  INV_X1 U29364 ( .A(n20700), .ZN(n20259) );
  NAND4_X1 U29365 ( .A1(n19977), .A2(n18730), .A3(n20259), .A4(n18729), .ZN(
        n18737) );
  AOI22_X1 U29366 ( .A1(n18731), .A2(n21617), .B1(n20240), .B2(n21630), .ZN(
        n18736) );
  AND2_X1 U29367 ( .A1(n20258), .A2(n20698), .ZN(n20695) );
  INV_X1 U29368 ( .A(n20695), .ZN(n18733) );
  NAND2_X1 U29369 ( .A1(n21615), .A2(n21619), .ZN(n18732) );
  NAND2_X1 U29370 ( .A1(n20259), .A2(n21614), .ZN(n21638) );
  AND2_X1 U29371 ( .A1(n21614), .A2(n19981), .ZN(n20247) );
  NAND3_X1 U29372 ( .A1(n21638), .A2(n21639), .A3(n20247), .ZN(n18734) );
  XNOR2_X1 U29373 ( .A(n51378), .B(n18739), .ZN(n18740) );
  XNOR2_X1 U29374 ( .A(n18742), .B(n18741), .ZN(n18744) );
  XNOR2_X1 U29375 ( .A(n44493), .B(n18745), .ZN(n42755) );
  XNOR2_X1 U29376 ( .A(n42755), .B(n43739), .ZN(n32738) );
  XNOR2_X1 U29377 ( .A(n37257), .B(n32738), .ZN(n18746) );
  XNOR2_X1 U29378 ( .A(n18747), .B(n18746), .ZN(n18748) );
  XNOR2_X1 U29379 ( .A(n18748), .B(n18749), .ZN(n18751) );
  XNOR2_X1 U29380 ( .A(n18750), .B(n18751), .ZN(n18753) );
  XNOR2_X1 U29381 ( .A(n18752), .B(n18753), .ZN(n18754) );
  INV_X1 U29382 ( .A(n21578), .ZN(n21560) );
  XNOR2_X1 U29383 ( .A(n18755), .B(n18756), .ZN(n18757) );
  XNOR2_X1 U29384 ( .A(n51437), .B(n18757), .ZN(n18767) );
  INV_X1 U29385 ( .A(n18759), .ZN(n18761) );
  INV_X1 U29386 ( .A(n24200), .ZN(n18760) );
  XNOR2_X1 U29387 ( .A(n18761), .B(n18760), .ZN(n34601) );
  XNOR2_X1 U29388 ( .A(n2112), .B(n4868), .ZN(n18762) );
  XNOR2_X1 U29389 ( .A(n35107), .B(n18762), .ZN(n33734) );
  XNOR2_X1 U29390 ( .A(n42083), .B(n33734), .ZN(n18763) );
  XNOR2_X1 U29391 ( .A(n34601), .B(n18763), .ZN(n18764) );
  XNOR2_X1 U29392 ( .A(n19203), .B(n18764), .ZN(n18765) );
  XNOR2_X1 U29393 ( .A(n18765), .B(n18505), .ZN(n18766) );
  XNOR2_X1 U29394 ( .A(n18769), .B(n18770), .ZN(n18771) );
  NAND2_X1 U29395 ( .A1(n21584), .A2(n21560), .ZN(n18789) );
  XNOR2_X1 U29396 ( .A(n18773), .B(n4578), .ZN(n19222) );
  XNOR2_X1 U29397 ( .A(n18774), .B(n19222), .ZN(n18784) );
  XNOR2_X1 U29398 ( .A(n24894), .B(n26289), .ZN(n18775) );
  XNOR2_X1 U29399 ( .A(n18776), .B(n18775), .ZN(n25992) );
  XNOR2_X1 U29400 ( .A(n25992), .B(n4880), .ZN(n41563) );
  XNOR2_X1 U29401 ( .A(n18777), .B(n41563), .ZN(n18782) );
  XNOR2_X1 U29402 ( .A(n25578), .B(n18778), .ZN(n33443) );
  XNOR2_X1 U29403 ( .A(n33443), .B(n842), .ZN(n18779) );
  XNOR2_X1 U29404 ( .A(n2162), .B(n18779), .ZN(n18781) );
  XNOR2_X1 U29405 ( .A(n18782), .B(n18781), .ZN(n18783) );
  XNOR2_X1 U29406 ( .A(n18784), .B(n18783), .ZN(n18786) );
  XNOR2_X1 U29407 ( .A(n18785), .B(n18786), .ZN(n18788) );
  MUX2_X1 U29408 ( .A(n21560), .B(n18789), .S(n21569), .Z(n20777) );
  XNOR2_X1 U29409 ( .A(n18791), .B(n18790), .ZN(n19245) );
  XNOR2_X1 U29410 ( .A(n28303), .B(n35796), .ZN(n18792) );
  XNOR2_X1 U29411 ( .A(n24638), .B(n18792), .ZN(n32277) );
  XNOR2_X1 U29412 ( .A(n28309), .B(n18793), .ZN(n36789) );
  XNOR2_X1 U29413 ( .A(n32277), .B(n36789), .ZN(n18794) );
  XNOR2_X1 U29414 ( .A(n18795), .B(n18794), .ZN(n18796) );
  XNOR2_X1 U29415 ( .A(n19245), .B(n18796), .ZN(n18800) );
  XNOR2_X1 U29416 ( .A(n52229), .B(n18798), .ZN(n18799) );
  XNOR2_X1 U29417 ( .A(n18802), .B(n18801), .ZN(n18803) );
  XNOR2_X1 U29418 ( .A(n2226), .B(n19244), .ZN(n18805) );
  XNOR2_X1 U29419 ( .A(n18806), .B(n18805), .ZN(n18807) );
  XNOR2_X1 U29420 ( .A(n18808), .B(n18807), .ZN(n19989) );
  XNOR2_X1 U29421 ( .A(n26526), .B(n4645), .ZN(n18809) );
  XNOR2_X1 U29422 ( .A(n25434), .B(n18809), .ZN(n18810) );
  XNOR2_X1 U29423 ( .A(n18810), .B(n37104), .ZN(n32930) );
  XNOR2_X1 U29424 ( .A(n25898), .B(n4627), .ZN(n37273) );
  XNOR2_X1 U29425 ( .A(n32930), .B(n37273), .ZN(n18811) );
  XNOR2_X1 U29426 ( .A(n19235), .B(n18811), .ZN(n18812) );
  XNOR2_X1 U29427 ( .A(n18813), .B(n18812), .ZN(n18814) );
  XNOR2_X1 U29428 ( .A(n18814), .B(n18815), .ZN(n18816) );
  XNOR2_X1 U29429 ( .A(n18817), .B(n18816), .ZN(n18822) );
  XNOR2_X1 U29430 ( .A(n18818), .B(n2217), .ZN(n18821) );
  NAND2_X1 U29431 ( .A1(n20777), .A2(n20601), .ZN(n18845) );
  NAND2_X1 U29432 ( .A1(n777), .A2(n18823), .ZN(n21568) );
  INV_X1 U29433 ( .A(n21568), .ZN(n21580) );
  XNOR2_X1 U29434 ( .A(n18824), .B(n18825), .ZN(n18839) );
  XNOR2_X1 U29435 ( .A(n18827), .B(n18826), .ZN(n18829) );
  XNOR2_X1 U29436 ( .A(n18829), .B(n18828), .ZN(n18835) );
  XNOR2_X1 U29437 ( .A(n41924), .B(n34215), .ZN(n18830) );
  XNOR2_X1 U29438 ( .A(n18831), .B(n18830), .ZN(n18833) );
  XNOR2_X1 U29439 ( .A(n18832), .B(n18833), .ZN(n18834) );
  XNOR2_X1 U29440 ( .A(n18835), .B(n18834), .ZN(n18837) );
  XNOR2_X1 U29441 ( .A(n18837), .B(n18836), .ZN(n18838) );
  AND2_X1 U29442 ( .A1(n21556), .A2(n21559), .ZN(n18840) );
  AOI22_X1 U29443 ( .A1(n18841), .A2(n20781), .B1(n21567), .B2(n18840), .ZN(
        n18844) );
  NAND2_X1 U29444 ( .A1(n20781), .A2(n21566), .ZN(n18842) );
  MUX2_X1 U29445 ( .A(n18842), .B(n21560), .S(n21412), .Z(n18843) );
  INV_X1 U29447 ( .A(n21663), .ZN(n20276) );
  OAI22_X1 U29448 ( .A1(n18847), .A2(n21648), .B1(n18846), .B2(n20276), .ZN(
        n18849) );
  NAND3_X1 U29449 ( .A1(n21664), .A2(n20270), .A3(n20266), .ZN(n20647) );
  NAND2_X1 U29450 ( .A1(n20267), .A2(n20647), .ZN(n18850) );
  NAND2_X1 U29451 ( .A1(n18850), .A2(n21649), .ZN(n18854) );
  XNOR2_X1 U29452 ( .A(n21660), .B(n21664), .ZN(n18851) );
  OAI211_X1 U29453 ( .C1(n18851), .C2(n3370), .A(n21654), .B(n20650), .ZN(
        n18852) );
  AND2_X1 U29454 ( .A1(n22605), .A2(n2210), .ZN(n22603) );
  INV_X1 U29455 ( .A(n22603), .ZN(n18856) );
  OAI21_X1 U29456 ( .B1(n24190), .B2(n4328), .A(n18856), .ZN(n18858) );
  NAND2_X1 U29457 ( .A1(n24190), .A2(n2210), .ZN(n23762) );
  INV_X1 U29458 ( .A(n23762), .ZN(n18857) );
  AOI21_X1 U29459 ( .B1(n4462), .B2(n18858), .A(n18857), .ZN(n18861) );
  AND2_X1 U29460 ( .A1(n24188), .A2(n2210), .ZN(n23872) );
  INV_X1 U29461 ( .A(n24190), .ZN(n24183) );
  OAI211_X1 U29462 ( .C1(n23872), .C2(n24180), .A(n24183), .B(n24189), .ZN(
        n18859) );
  NAND2_X1 U29463 ( .A1(n24186), .A2(n24187), .ZN(n23203) );
  INV_X1 U29464 ( .A(n23203), .ZN(n23764) );
  NAND2_X1 U29465 ( .A1(n18859), .A2(n23764), .ZN(n18860) );
  NOR2_X1 U29467 ( .A1(n20239), .A2(n760), .ZN(n18866) );
  NAND3_X1 U29468 ( .A1(n18862), .A2(n1597), .A3(n20230), .ZN(n18864) );
  INV_X1 U29469 ( .A(n18867), .ZN(n18871) );
  OAI22_X1 U29470 ( .A1(n20679), .A2(n18101), .B1(n20685), .B2(n51090), .ZN(
        n18870) );
  OAI21_X1 U29471 ( .B1(n18871), .B2(n18870), .A(n18869), .ZN(n18880) );
  NOR2_X1 U29472 ( .A1(n18872), .A2(n20668), .ZN(n18876) );
  NOR2_X1 U29473 ( .A1(n1597), .A2(n18873), .ZN(n18874) );
  AOI22_X1 U29474 ( .A1(n20679), .A2(n18876), .B1(n18875), .B2(n18874), .ZN(
        n18879) );
  NAND2_X1 U29475 ( .A1(n20679), .A2(n760), .ZN(n18877) );
  INV_X1 U29476 ( .A(n23317), .ZN(n23312) );
  OR2_X1 U29477 ( .A1(n18985), .A2(n21300), .ZN(n19715) );
  NAND2_X1 U29478 ( .A1(n18992), .A2(n18882), .ZN(n21290) );
  INV_X1 U29479 ( .A(n18996), .ZN(n19713) );
  NAND2_X1 U29480 ( .A1(n19713), .A2(n19792), .ZN(n18883) );
  INV_X1 U29481 ( .A(n19793), .ZN(n21296) );
  NAND2_X1 U29483 ( .A1(n18992), .A2(n766), .ZN(n18885) );
  NAND2_X1 U29484 ( .A1(n18886), .A2(n18885), .ZN(n18887) );
  AOI22_X1 U29487 ( .A1(n19721), .A2(n19792), .B1(n19797), .B2(n21293), .ZN(
        n18891) );
  NAND2_X1 U29488 ( .A1(n18992), .A2(n19796), .ZN(n18990) );
  NAND2_X1 U29490 ( .A1(n23312), .A2(n23314), .ZN(n21004) );
  INV_X1 U29491 ( .A(n18896), .ZN(n21524) );
  OAI211_X1 U29492 ( .C1(n18898), .C2(n52210), .A(n20608), .B(n21524), .ZN(
        n18900) );
  NAND2_X1 U29493 ( .A1(n18900), .A2(n18899), .ZN(n18901) );
  NAND3_X1 U29494 ( .A1(n18903), .A2(n21525), .A3(n20611), .ZN(n18904) );
  NAND2_X1 U29495 ( .A1(n19861), .A2(n19848), .ZN(n18906) );
  AND2_X1 U29496 ( .A1(n19643), .A2(n19649), .ZN(n18907) );
  OAI21_X1 U29497 ( .B1(n19030), .B2(n18907), .A(n19851), .ZN(n18913) );
  INV_X1 U29498 ( .A(n19870), .ZN(n19850) );
  NAND2_X1 U29499 ( .A1(n19643), .A2(n51039), .ZN(n19744) );
  INV_X1 U29500 ( .A(n19744), .ZN(n18909) );
  AND2_X1 U29501 ( .A1(n19846), .A2(n19647), .ZN(n18908) );
  AOI22_X1 U29502 ( .A1(n19850), .A2(n18909), .B1(n19853), .B2(n18908), .ZN(
        n18912) );
  NAND2_X1 U29503 ( .A1(n18910), .A2(n585), .ZN(n18911) );
  NAND2_X1 U29504 ( .A1(n19685), .A2(n20211), .ZN(n18914) );
  AND2_X1 U29505 ( .A1(n19688), .A2(n18914), .ZN(n18915) );
  AOI22_X1 U29506 ( .A1(n18915), .A2(n20209), .B1(n775), .B2(n19671), .ZN(
        n18919) );
  NAND2_X1 U29507 ( .A1(n18916), .A2(n19689), .ZN(n18917) );
  NAND4_X1 U29508 ( .A1(n18920), .A2(n18919), .A3(n18918), .A4(n18917), .ZN(
        n18925) );
  NAND2_X1 U29509 ( .A1(n20217), .A2(n20215), .ZN(n18923) );
  NAND2_X1 U29510 ( .A1(n20212), .A2(n18921), .ZN(n18922) );
  AOI21_X1 U29511 ( .B1(n20208), .B2(n18923), .A(n18922), .ZN(n18924) );
  NAND3_X1 U29512 ( .A1(n21864), .A2(n23317), .A3(n23316), .ZN(n18926) );
  NAND4_X1 U29514 ( .A1(n19884), .A2(n19636), .A3(n19894), .A4(n19662), .ZN(
        n18930) );
  NAND3_X1 U29515 ( .A1(n19896), .A2(n19887), .A3(n51127), .ZN(n18929) );
  INV_X1 U29516 ( .A(n18927), .ZN(n18928) );
  INV_X1 U29517 ( .A(n18931), .ZN(n18952) );
  AND2_X1 U29518 ( .A1(n18935), .A2(n18934), .ZN(n18951) );
  INV_X1 U29519 ( .A(n19896), .ZN(n18939) );
  OAI22_X1 U29521 ( .A1(n18939), .A2(n18938), .B1(n51127), .B2(n18937), .ZN(
        n18940) );
  NAND2_X1 U29522 ( .A1(n18940), .A2(n18942), .ZN(n18950) );
  OAI21_X1 U29523 ( .B1(n19659), .B2(n19891), .A(n19893), .ZN(n18948) );
  INV_X1 U29524 ( .A(n18941), .ZN(n18943) );
  AOI21_X1 U29525 ( .B1(n18943), .B2(n19663), .A(n18942), .ZN(n18947) );
  NAND2_X1 U29527 ( .A1(n18945), .A2(n51127), .ZN(n18946) );
  NAND3_X1 U29528 ( .A1(n18948), .A2(n18947), .A3(n18946), .ZN(n18949) );
  NAND4_X2 U29529 ( .A1(n18952), .A2(n18949), .A3(n18950), .A4(n18951), .ZN(
        n23306) );
  NAND2_X1 U29530 ( .A1(n22255), .A2(n23314), .ZN(n18959) );
  AND2_X1 U29531 ( .A1(n8303), .A2(n23306), .ZN(n18953) );
  OAI22_X1 U29532 ( .A1(n23320), .A2(n18953), .B1(n22251), .B2(n441), .ZN(
        n18954) );
  NAND2_X1 U29533 ( .A1(n18954), .A2(n23303), .ZN(n18958) );
  OAI21_X1 U29534 ( .B1(n23310), .B2(n23316), .A(n23317), .ZN(n18956) );
  NOR2_X1 U29535 ( .A1(n23314), .A2(n21873), .ZN(n22958) );
  INV_X1 U29536 ( .A(n23306), .ZN(n22964) );
  NAND2_X1 U29537 ( .A1(n22964), .A2(n441), .ZN(n23311) );
  INV_X1 U29538 ( .A(n23311), .ZN(n18955) );
  OAI21_X1 U29539 ( .B1(n18956), .B2(n22958), .A(n18955), .ZN(n18957) );
  AND2_X1 U29541 ( .A1(n19087), .A2(n3335), .ZN(n18965) );
  INV_X1 U29542 ( .A(n21253), .ZN(n19478) );
  NAND2_X1 U29543 ( .A1(n19097), .A2(n19478), .ZN(n18964) );
  AND2_X1 U29546 ( .A1(n19475), .A2(n19087), .ZN(n19473) );
  INV_X1 U29547 ( .A(n21243), .ZN(n19085) );
  AOI21_X1 U29548 ( .B1(n19473), .B2(n21257), .A(n18968), .ZN(n18971) );
  AOI22_X1 U29549 ( .A1(n21250), .A2(n21249), .B1(n21245), .B2(n18969), .ZN(
        n18970) );
  INV_X1 U29550 ( .A(n19840), .ZN(n19701) );
  NAND2_X1 U29551 ( .A1(n21186), .A2(n51434), .ZN(n21182) );
  NAND2_X1 U29552 ( .A1(n19828), .A2(n21173), .ZN(n21180) );
  MUX2_X1 U29553 ( .A(n19701), .B(n21182), .S(n21180), .Z(n18978) );
  INV_X1 U29554 ( .A(n18973), .ZN(n18974) );
  INV_X1 U29556 ( .A(n19524), .ZN(n19841) );
  INV_X1 U29557 ( .A(n18975), .ZN(n18976) );
  NAND4_X1 U29558 ( .A1(n18978), .A2(n18977), .A3(n19526), .A4(n2299), .ZN(
        n18984) );
  NAND2_X1 U29559 ( .A1(n19524), .A2(n19837), .ZN(n21187) );
  AOI21_X1 U29560 ( .B1(n19703), .B2(n21173), .A(n19832), .ZN(n18981) );
  NAND2_X1 U29561 ( .A1(n19834), .A2(n17201), .ZN(n19523) );
  NAND2_X1 U29562 ( .A1(n21186), .A2(n19826), .ZN(n19525) );
  INV_X1 U29563 ( .A(n19525), .ZN(n18979) );
  NAND3_X1 U29564 ( .A1(n19523), .A2(n18979), .A3(n17201), .ZN(n18980) );
  NAND3_X1 U29565 ( .A1(n21187), .A2(n18981), .A3(n18980), .ZN(n18983) );
  INV_X1 U29566 ( .A(n19529), .ZN(n21172) );
  OAI21_X1 U29567 ( .B1(n19826), .B2(n21172), .A(n19700), .ZN(n18982) );
  OR2_X1 U29568 ( .A1(n22979), .A2(n22978), .ZN(n19754) );
  INV_X1 U29569 ( .A(n18985), .ZN(n21295) );
  NAND2_X1 U29570 ( .A1(n18992), .A2(n21293), .ZN(n18987) );
  AOI21_X1 U29571 ( .B1(n18999), .B2(n18987), .A(n18986), .ZN(n18988) );
  NOR2_X1 U29572 ( .A1(n18992), .A2(n18996), .ZN(n19720) );
  OAI21_X1 U29573 ( .B1(n18992), .B2(n21300), .A(n18991), .ZN(n18993) );
  OAI211_X1 U29574 ( .C1(n19794), .C2(n21300), .A(n18994), .B(n18993), .ZN(
        n19004) );
  NAND3_X1 U29575 ( .A1(n19716), .A2(n21295), .A3(n18996), .ZN(n19001) );
  NAND2_X1 U29576 ( .A1(n18997), .A2(n509), .ZN(n18998) );
  OAI22_X1 U29577 ( .A1(n18999), .A2(n18998), .B1(n19796), .B2(n19795), .ZN(
        n19000) );
  NAND3_X1 U29578 ( .A1(n19002), .A2(n19001), .A3(n19000), .ZN(n19003) );
  AND2_X1 U29579 ( .A1(n21214), .A2(n6078), .ZN(n19006) );
  INV_X1 U29580 ( .A(n21215), .ZN(n19732) );
  NAND2_X1 U29581 ( .A1(n19820), .A2(n21200), .ZN(n19727) );
  INV_X1 U29582 ( .A(n19727), .ZN(n19005) );
  INV_X1 U29583 ( .A(n19813), .ZN(n19011) );
  OAI22_X1 U29585 ( .A1(n19009), .A2(n19008), .B1(n19814), .B2(n19007), .ZN(
        n19010) );
  NAND3_X1 U29586 ( .A1(n19010), .A2(n19819), .A3(n19823), .ZN(n19015) );
  OAI21_X1 U29587 ( .B1(n19011), .B2(n21200), .A(n2229), .ZN(n19014) );
  NOR2_X1 U29588 ( .A1(n21200), .A2(n21213), .ZN(n19013) );
  NAND2_X1 U29589 ( .A1(n22989), .A2(n22977), .ZN(n19757) );
  NAND2_X1 U29590 ( .A1(n19754), .A2(n19757), .ZN(n19036) );
  NOR2_X1 U29591 ( .A1(n21283), .A2(n19122), .ZN(n21286) );
  AOI21_X1 U29592 ( .B1(n19023), .B2(n51013), .A(n21269), .ZN(n19017) );
  NAND2_X1 U29593 ( .A1(n21270), .A2(n19452), .ZN(n19461) );
  OAI22_X1 U29594 ( .A1(n19455), .A2(n21283), .B1(n19785), .B2(n19461), .ZN(
        n19018) );
  INV_X1 U29595 ( .A(n19019), .ZN(n21287) );
  AND2_X1 U29596 ( .A1(n19452), .A2(n21287), .ZN(n19784) );
  INV_X1 U29597 ( .A(n19784), .ZN(n19021) );
  OAI21_X1 U29598 ( .B1(n19785), .B2(n19021), .A(n19020), .ZN(n19022) );
  INV_X1 U29599 ( .A(n19022), .ZN(n19026) );
  NAND2_X1 U29600 ( .A1(n19023), .A2(n21269), .ZN(n19024) );
  OAI211_X1 U29601 ( .C1(n21271), .C2(n51013), .A(n19122), .B(n19024), .ZN(
        n19025) );
  NAND2_X1 U29602 ( .A1(n19643), .A2(n19866), .ZN(n19027) );
  OAI22_X1 U29603 ( .A1(n585), .A2(n19027), .B1(n19846), .B2(n19642), .ZN(
        n19029) );
  OAI21_X1 U29604 ( .B1(n19873), .B2(n19033), .A(n19640), .ZN(n19028) );
  AOI22_X1 U29605 ( .A1(n19029), .A2(n19647), .B1(n19028), .B2(n19639), .ZN(
        n19035) );
  INV_X1 U29606 ( .A(n19865), .ZN(n19874) );
  OAI211_X1 U29607 ( .C1(n19851), .C2(n19033), .A(n19032), .B(n19848), .ZN(
        n19034) );
  NAND2_X1 U29608 ( .A1(n19036), .A2(n19758), .ZN(n19043) );
  INV_X1 U29609 ( .A(n22999), .ZN(n19042) );
  NAND2_X1 U29610 ( .A1(n22558), .A2(n22989), .ZN(n22992) );
  AND2_X1 U29611 ( .A1(n22978), .A2(n22983), .ZN(n19762) );
  NAND2_X1 U29612 ( .A1(n22982), .A2(n22977), .ZN(n19761) );
  NAND3_X1 U29613 ( .A1(n22992), .A2(n19762), .A3(n19038), .ZN(n19041) );
  OR2_X1 U29614 ( .A1(n22978), .A2(n22983), .ZN(n22993) );
  NAND3_X1 U29615 ( .A1(n22985), .A2(n22557), .A3(n22982), .ZN(n19755) );
  INV_X1 U29616 ( .A(n19755), .ZN(n19039) );
  NAND2_X1 U29617 ( .A1(n22993), .A2(n19039), .ZN(n19040) );
  XNOR2_X1 U29618 ( .A(n26530), .B(n25548), .ZN(n25831) );
  OAI211_X1 U29619 ( .C1(n19044), .C2(n51815), .A(n52176), .B(n19047), .ZN(
        n19053) );
  MUX2_X1 U29620 ( .A(n20156), .B(n19535), .S(n20124), .Z(n19046) );
  OAI21_X1 U29621 ( .B1(n19050), .B2(n19049), .A(n19543), .ZN(n19051) );
  NAND3_X1 U29622 ( .A1(n20158), .A2(n20157), .A3(n20156), .ZN(n19054) );
  OAI211_X1 U29623 ( .C1(n20158), .C2(n19056), .A(n19055), .B(n19054), .ZN(
        n19058) );
  NAND2_X1 U29624 ( .A1(n19058), .A2(n51815), .ZN(n19060) );
  INV_X1 U29625 ( .A(n19067), .ZN(n19063) );
  OAI21_X1 U29626 ( .B1(n19063), .B2(n19062), .A(n19061), .ZN(n19084) );
  AOI21_X1 U29627 ( .B1(n19065), .B2(n20143), .A(n19064), .ZN(n19069) );
  NAND2_X1 U29628 ( .A1(n19067), .A2(n19066), .ZN(n19068) );
  NAND2_X1 U29629 ( .A1(n19069), .A2(n19068), .ZN(n19083) );
  NAND2_X1 U29630 ( .A1(n19071), .A2(n19070), .ZN(n19072) );
  AND3_X1 U29631 ( .A1(n19073), .A2(n19074), .A3(n19072), .ZN(n19082) );
  INV_X1 U29632 ( .A(n19077), .ZN(n19079) );
  OAI21_X1 U29633 ( .B1(n19079), .B2(n20144), .A(n19078), .ZN(n19080) );
  NAND2_X1 U29634 ( .A1(n20130), .A2(n19080), .ZN(n19081) );
  AOI21_X1 U29635 ( .B1(n19087), .B2(n19086), .A(n19085), .ZN(n19092) );
  AND2_X1 U29636 ( .A1(n3335), .A2(n51222), .ZN(n19103) );
  NAND2_X1 U29637 ( .A1(n19475), .A2(n19103), .ZN(n19091) );
  INV_X1 U29638 ( .A(n19089), .ZN(n19090) );
  OAI21_X1 U29639 ( .B1(n21253), .B2(n19099), .A(n19093), .ZN(n19096) );
  INV_X1 U29640 ( .A(n19094), .ZN(n19095) );
  AOI22_X1 U29641 ( .A1(n21249), .A2(n19096), .B1(n19095), .B2(n19472), .ZN(
        n19107) );
  OAI21_X1 U29642 ( .B1(n19099), .B2(n19098), .A(n19097), .ZN(n19100) );
  OAI21_X1 U29643 ( .B1(n19101), .B2(n19100), .A(n21242), .ZN(n19106) );
  NAND2_X1 U29644 ( .A1(n19104), .A2(n19103), .ZN(n19105) );
  NOR2_X1 U29645 ( .A1(n19108), .A2(n19518), .ZN(n19109) );
  INV_X1 U29646 ( .A(n19505), .ZN(n19111) );
  AOI22_X1 U29647 ( .A1(n19114), .A2(n19520), .B1(n19514), .B2(n19510), .ZN(
        n19115) );
  NAND2_X1 U29648 ( .A1(n23237), .A2(n22654), .ZN(n22132) );
  AND2_X1 U29649 ( .A1(n21276), .A2(n19777), .ZN(n19120) );
  NAND2_X1 U29650 ( .A1(n21281), .A2(n19120), .ZN(n19130) );
  INV_X1 U29651 ( .A(n19455), .ZN(n21272) );
  OAI21_X1 U29652 ( .B1(n21272), .B2(n19459), .A(n51013), .ZN(n19117) );
  OAI21_X1 U29653 ( .B1(n21283), .B2(n19452), .A(n21269), .ZN(n19116) );
  AND2_X1 U29654 ( .A1(n19117), .A2(n19116), .ZN(n19129) );
  AND2_X1 U29655 ( .A1(n19778), .A2(n19777), .ZN(n19786) );
  NAND3_X1 U29656 ( .A1(n19786), .A2(n21271), .A3(n51013), .ZN(n19126) );
  NAND4_X1 U29657 ( .A1(n19455), .A2(n21287), .A3(n2182), .A4(n21269), .ZN(
        n19125) );
  INV_X1 U29658 ( .A(n19120), .ZN(n19121) );
  NAND2_X1 U29659 ( .A1(n19122), .A2(n19121), .ZN(n19123) );
  OAI211_X1 U29660 ( .C1(n19775), .C2(n51013), .A(n19123), .B(n5229), .ZN(
        n19124) );
  NAND4_X1 U29661 ( .A1(n19127), .A2(n19126), .A3(n19125), .A4(n19124), .ZN(
        n19128) );
  NOR2_X1 U29663 ( .A1(n19131), .A2(n20075), .ZN(n19134) );
  OAI22_X1 U29664 ( .A1(n20052), .A2(n20072), .B1(n19132), .B2(n2101), .ZN(
        n19133) );
  NOR2_X1 U29665 ( .A1(n19134), .A2(n19133), .ZN(n19147) );
  OAI22_X1 U29666 ( .A1(n20060), .A2(n19136), .B1(n19135), .B2(n20073), .ZN(
        n19137) );
  NAND2_X1 U29667 ( .A1(n19137), .A2(n19499), .ZN(n19146) );
  INV_X1 U29668 ( .A(n19138), .ZN(n19139) );
  NAND2_X1 U29669 ( .A1(n19139), .A2(n19493), .ZN(n19145) );
  NAND2_X1 U29670 ( .A1(n2101), .A2(n4459), .ZN(n19142) );
  OAI211_X1 U29671 ( .C1(n20063), .C2(n20075), .A(n19143), .B(n19142), .ZN(
        n19144) );
  NAND4_X2 U29672 ( .A1(n19146), .A2(n19147), .A3(n19145), .A4(n19144), .ZN(
        n23257) );
  NAND2_X1 U29673 ( .A1(n23238), .A2(n23257), .ZN(n21851) );
  INV_X1 U29674 ( .A(n21851), .ZN(n19148) );
  NAND2_X1 U29675 ( .A1(n22132), .A2(n19148), .ZN(n19155) );
  INV_X1 U29676 ( .A(n19149), .ZN(n23245) );
  AND2_X1 U29677 ( .A1(n22658), .A2(n23245), .ZN(n19151) );
  INV_X1 U29678 ( .A(n23257), .ZN(n23246) );
  NAND2_X1 U29679 ( .A1(n23246), .A2(n23244), .ZN(n22123) );
  INV_X1 U29680 ( .A(n22123), .ZN(n19150) );
  NOR2_X1 U29681 ( .A1(n23247), .A2(n23246), .ZN(n22650) );
  NAND3_X1 U29682 ( .A1(n22650), .A2(n22124), .A3(n628), .ZN(n19153) );
  INV_X1 U29683 ( .A(n28287), .ZN(n19320) );
  INV_X1 U29684 ( .A(n21430), .ZN(n19157) );
  NOR2_X1 U29685 ( .A1(n19157), .A2(n21420), .ZN(n19159) );
  NOR2_X1 U29686 ( .A1(n19159), .A2(n19158), .ZN(n19169) );
  INV_X1 U29687 ( .A(n20837), .ZN(n19160) );
  OAI21_X1 U29688 ( .B1(n19160), .B2(n21442), .A(n19957), .ZN(n19161) );
  NAND2_X1 U29689 ( .A1(n19161), .A2(n21443), .ZN(n19168) );
  OAI21_X1 U29690 ( .B1(n21427), .B2(n5500), .A(n21424), .ZN(n19164) );
  INV_X1 U29691 ( .A(n19162), .ZN(n19163) );
  NAND2_X1 U29692 ( .A1(n19164), .A2(n19163), .ZN(n19165) );
  NAND2_X1 U29693 ( .A1(n19165), .A2(n21422), .ZN(n19167) );
  AND2_X1 U29694 ( .A1(n5499), .A2(n52139), .ZN(n19956) );
  INV_X1 U29695 ( .A(n20321), .ZN(n19945) );
  NAND4_X2 U29696 ( .A1(n19169), .A2(n19168), .A3(n19167), .A4(n19166), .ZN(
        n22426) );
  INV_X1 U29697 ( .A(n20420), .ZN(n19172) );
  NAND2_X1 U29698 ( .A1(n20359), .A2(n20422), .ZN(n19175) );
  NAND3_X1 U29699 ( .A1(n20354), .A2(n19170), .A3(n19175), .ZN(n19171) );
  NAND2_X1 U29700 ( .A1(n40), .A2(n20435), .ZN(n19327) );
  NAND2_X1 U29701 ( .A1(n20432), .A2(n20422), .ZN(n19176) );
  NAND2_X1 U29702 ( .A1(n19178), .A2(n20426), .ZN(n19179) );
  XNOR2_X1 U29703 ( .A(n26419), .B(n19182), .ZN(n42549) );
  XNOR2_X1 U29704 ( .A(n24992), .B(n4502), .ZN(n33199) );
  XNOR2_X1 U29705 ( .A(n33199), .B(n43586), .ZN(n42973) );
  XNOR2_X1 U29706 ( .A(n42549), .B(n42973), .ZN(n19183) );
  XNOR2_X1 U29707 ( .A(n19183), .B(n33201), .ZN(n19184) );
  XNOR2_X1 U29708 ( .A(n19185), .B(n19184), .ZN(n19187) );
  XNOR2_X1 U29709 ( .A(n19186), .B(n19187), .ZN(n19189) );
  XNOR2_X1 U29710 ( .A(n19188), .B(n19189), .ZN(n19191) );
  XNOR2_X1 U29711 ( .A(n19191), .B(n19190), .ZN(n19193) );
  XNOR2_X1 U29712 ( .A(n19193), .B(n19192), .ZN(n19195) );
  XNOR2_X1 U29713 ( .A(n19195), .B(n19194), .ZN(n19965) );
  XNOR2_X1 U29714 ( .A(n14903), .B(n19196), .ZN(n19197) );
  XNOR2_X1 U29715 ( .A(n19198), .B(n19197), .ZN(n19207) );
  XNOR2_X1 U29716 ( .A(n14427), .B(n19199), .ZN(n19205) );
  XNOR2_X1 U29717 ( .A(n34411), .B(n4045), .ZN(n24505) );
  XNOR2_X1 U29718 ( .A(n24505), .B(n43922), .ZN(n24708) );
  XNOR2_X1 U29719 ( .A(n24708), .B(n4431), .ZN(n45307) );
  XNOR2_X1 U29720 ( .A(n42630), .B(Key[189]), .ZN(n34252) );
  XNOR2_X1 U29721 ( .A(n45307), .B(n34252), .ZN(n19201) );
  XNOR2_X1 U29722 ( .A(n4423), .B(n4896), .ZN(n19200) );
  XNOR2_X1 U29723 ( .A(n33934), .B(n19200), .ZN(n33432) );
  XNOR2_X1 U29724 ( .A(n19201), .B(n33432), .ZN(n19202) );
  XNOR2_X1 U29725 ( .A(n19203), .B(n19202), .ZN(n19204) );
  XNOR2_X1 U29726 ( .A(n19205), .B(n19204), .ZN(n19206) );
  XNOR2_X1 U29727 ( .A(n19207), .B(n19206), .ZN(n19208) );
  XNOR2_X1 U29728 ( .A(n19210), .B(n19211), .ZN(n19212) );
  XNOR2_X1 U29729 ( .A(n51047), .B(n2181), .ZN(n19215) );
  XNOR2_X1 U29730 ( .A(n19216), .B(n19215), .ZN(n19226) );
  XNOR2_X1 U29731 ( .A(n4482), .B(n4597), .ZN(n19217) );
  XNOR2_X1 U29732 ( .A(n19218), .B(n19217), .ZN(n19219) );
  XNOR2_X1 U29733 ( .A(n19219), .B(n24430), .ZN(n33242) );
  XNOR2_X1 U29734 ( .A(n33242), .B(n3383), .ZN(n19220) );
  XNOR2_X1 U29735 ( .A(n19220), .B(n34893), .ZN(n19221) );
  XNOR2_X1 U29736 ( .A(n19222), .B(n19221), .ZN(n19224) );
  XNOR2_X1 U29737 ( .A(n19223), .B(n19224), .ZN(n19225) );
  XNOR2_X1 U29738 ( .A(n19226), .B(n19225), .ZN(n19232) );
  XNOR2_X1 U29739 ( .A(n19228), .B(n19227), .ZN(n19230) );
  XNOR2_X1 U29740 ( .A(n19229), .B(n19230), .ZN(n19231) );
  XNOR2_X1 U29741 ( .A(n2220), .B(n21495), .ZN(n19276) );
  XNOR2_X1 U29742 ( .A(n4287), .B(n3481), .ZN(n25822) );
  XNOR2_X1 U29743 ( .A(n25822), .B(n4535), .ZN(n35553) );
  XNOR2_X1 U29744 ( .A(n33986), .B(n35553), .ZN(n19233) );
  XNOR2_X1 U29745 ( .A(n40849), .B(n19233), .ZN(n19234) );
  XNOR2_X1 U29746 ( .A(n19235), .B(n19234), .ZN(n19236) );
  XNOR2_X1 U29747 ( .A(n19237), .B(n19236), .ZN(n19238) );
  XNOR2_X1 U29748 ( .A(n19239), .B(n19238), .ZN(n19241) );
  XNOR2_X1 U29749 ( .A(n19241), .B(n19240), .ZN(n19242) );
  XNOR2_X1 U29750 ( .A(n19242), .B(n19243), .ZN(n19280) );
  INV_X1 U29751 ( .A(n19280), .ZN(n20821) );
  XNOR2_X1 U29752 ( .A(n19245), .B(n19244), .ZN(n19252) );
  XNOR2_X1 U29753 ( .A(n46097), .B(n26385), .ZN(n26041) );
  XNOR2_X1 U29754 ( .A(n26041), .B(n35539), .ZN(n37291) );
  XNOR2_X1 U29755 ( .A(n19246), .B(n4121), .ZN(n32941) );
  XNOR2_X1 U29756 ( .A(n37291), .B(n32941), .ZN(n19247) );
  XNOR2_X1 U29757 ( .A(n19248), .B(n19247), .ZN(n19249) );
  XNOR2_X1 U29758 ( .A(n19250), .B(n19249), .ZN(n19251) );
  XNOR2_X1 U29759 ( .A(n19252), .B(n19251), .ZN(n19257) );
  NAND2_X1 U29762 ( .A1(n20821), .A2(n20825), .ZN(n21485) );
  XNOR2_X1 U29763 ( .A(n19260), .B(n19261), .ZN(n19265) );
  XNOR2_X1 U29764 ( .A(n19262), .B(n24612), .ZN(n35499) );
  XNOR2_X1 U29765 ( .A(n25372), .B(n42258), .ZN(n35361) );
  XNOR2_X1 U29766 ( .A(n4923), .B(n4934), .ZN(n42537) );
  XNOR2_X1 U29767 ( .A(n35361), .B(n42537), .ZN(n19263) );
  XNOR2_X1 U29768 ( .A(n35499), .B(n19263), .ZN(n19264) );
  XNOR2_X1 U29769 ( .A(n19265), .B(n19264), .ZN(n19269) );
  XNOR2_X1 U29770 ( .A(n19267), .B(n19266), .ZN(n19268) );
  XNOR2_X1 U29771 ( .A(n19269), .B(n19268), .ZN(n19270) );
  XNOR2_X1 U29772 ( .A(n19271), .B(n19270), .ZN(n19273) );
  OAI21_X1 U29773 ( .B1(n21485), .B2(n21495), .A(n20334), .ZN(n19275) );
  INV_X1 U29774 ( .A(n20334), .ZN(n19966) );
  NAND2_X1 U29775 ( .A1(n20815), .A2(n21492), .ZN(n19967) );
  NAND3_X1 U29777 ( .A1(n21494), .A2(n20826), .A3(n2221), .ZN(n19279) );
  INV_X1 U29778 ( .A(n19965), .ZN(n21486) );
  AND2_X1 U29779 ( .A1(n21486), .A2(n20334), .ZN(n20827) );
  AND2_X1 U29781 ( .A1(n2221), .A2(n19969), .ZN(n20813) );
  INV_X1 U29782 ( .A(n20813), .ZN(n20449) );
  NAND2_X1 U29783 ( .A1(n20334), .A2(n20441), .ZN(n21490) );
  INV_X1 U29785 ( .A(n20815), .ZN(n21491) );
  INV_X1 U29787 ( .A(n21356), .ZN(n21596) );
  AOI21_X1 U29788 ( .B1(n21350), .B2(n52208), .A(n21596), .ZN(n19287) );
  OR2_X1 U29789 ( .A1(n21360), .A2(n19285), .ZN(n21597) );
  INV_X1 U29790 ( .A(n19286), .ZN(n20771) );
  OAI211_X1 U29791 ( .C1(n19289), .C2(n21354), .A(n19288), .B(n21596), .ZN(
        n19292) );
  NAND2_X1 U29792 ( .A1(n19290), .A2(n21359), .ZN(n19291) );
  INV_X1 U29793 ( .A(n19293), .ZN(n21592) );
  NOR2_X1 U29794 ( .A1(n21351), .A2(n21601), .ZN(n19295) );
  NAND2_X1 U29795 ( .A1(n19296), .A2(n19295), .ZN(n19930) );
  INV_X1 U29796 ( .A(n19930), .ZN(n19297) );
  NAND2_X1 U29797 ( .A1(n19297), .A2(n21350), .ZN(n19298) );
  NAND2_X1 U29799 ( .A1(n20375), .A2(n5923), .ZN(n21374) );
  NAND2_X1 U29800 ( .A1(n21389), .A2(n20415), .ZN(n20794) );
  NAND2_X1 U29801 ( .A1(n20408), .A2(n20375), .ZN(n21383) );
  OAI21_X1 U29802 ( .B1(n21383), .B2(n21389), .A(n358), .ZN(n19301) );
  NAND2_X1 U29803 ( .A1(n19301), .A2(n21388), .ZN(n19304) );
  NAND4_X1 U29804 ( .A1(n20416), .A2(n769), .A3(n20805), .A4(n21375), .ZN(
        n19303) );
  INV_X1 U29805 ( .A(n20791), .ZN(n20380) );
  OAI211_X1 U29806 ( .C1(n21397), .C2(n21388), .A(n21396), .B(n20380), .ZN(
        n19302) );
  MUX2_X1 U29807 ( .A(n22426), .B(n23992), .S(n23982), .Z(n19305) );
  AOI22_X1 U29808 ( .A1(n23036), .A2(n23982), .B1(n22427), .B2(n19305), .ZN(
        n19319) );
  NAND2_X1 U29809 ( .A1(n21449), .A2(n20493), .ZN(n19310) );
  INV_X1 U29810 ( .A(n21449), .ZN(n21459) );
  NAND3_X1 U29811 ( .A1(n19364), .A2(n21460), .A3(n21474), .ZN(n21475) );
  NAND3_X1 U29813 ( .A1(n19351), .A2(n19357), .A3(n21450), .ZN(n19306) );
  INV_X1 U29814 ( .A(n20316), .ZN(n19363) );
  OAI222_X1 U29815 ( .A1(n19363), .A2(n21474), .B1(n21458), .B2(n21469), .C1(
        n767), .C2(n52146), .ZN(n19307) );
  NAND3_X1 U29817 ( .A1(n20316), .A2(n20493), .A3(n21464), .ZN(n19309) );
  NAND3_X1 U29818 ( .A1(n21460), .A2(n20493), .A3(n19362), .ZN(n19308) );
  OAI211_X1 U29819 ( .C1(n19310), .C2(n21458), .A(n19309), .B(n19308), .ZN(
        n19311) );
  NAND2_X1 U29820 ( .A1(n19311), .A2(n20487), .ZN(n19312) );
  NAND2_X1 U29821 ( .A1(n6967), .A2(n23982), .ZN(n23037) );
  OAI21_X1 U29822 ( .B1(n23998), .B2(n23981), .A(n23037), .ZN(n19315) );
  INV_X1 U29823 ( .A(n22426), .ZN(n23984) );
  NOR2_X1 U29824 ( .A1(n23995), .A2(n23984), .ZN(n19314) );
  NOR2_X1 U29825 ( .A1(n19315), .A2(n19314), .ZN(n19318) );
  OAI21_X1 U29827 ( .B1(n23992), .B2(n23987), .A(n22428), .ZN(n19316) );
  NAND2_X1 U29828 ( .A1(n22534), .A2(n19316), .ZN(n19317) );
  NAND2_X1 U29829 ( .A1(n22426), .A2(n24000), .ZN(n23996) );
  XNOR2_X1 U29830 ( .A(n26529), .B(n19320), .ZN(n25442) );
  INV_X1 U29831 ( .A(n25442), .ZN(n27506) );
  AOI21_X1 U29832 ( .B1(n5875), .B2(n20426), .A(n20435), .ZN(n19321) );
  INV_X1 U29833 ( .A(n20423), .ZN(n19323) );
  NAND2_X1 U29834 ( .A1(n19326), .A2(n20428), .ZN(n19329) );
  INV_X1 U29835 ( .A(n19327), .ZN(n19328) );
  NAND2_X1 U29836 ( .A1(n19332), .A2(n6452), .ZN(n19333) );
  OAI21_X1 U29837 ( .B1(n19337), .B2(n489), .A(n19335), .ZN(n19338) );
  INV_X1 U29838 ( .A(n19339), .ZN(n19340) );
  OAI211_X1 U29839 ( .C1(n20504), .C2(n8687), .A(n19341), .B(n19340), .ZN(
        n19342) );
  AND2_X1 U29840 ( .A1(n20507), .A2(n19344), .ZN(n19347) );
  INV_X1 U29841 ( .A(n19345), .ZN(n19346) );
  AOI21_X1 U29842 ( .B1(n19348), .B2(n19347), .A(n19346), .ZN(n19350) );
  INV_X1 U29843 ( .A(n19352), .ZN(n21455) );
  OR2_X1 U29844 ( .A1(n19353), .A2(n21455), .ZN(n19369) );
  NAND3_X1 U29845 ( .A1(n20316), .A2(n20488), .A3(n21465), .ZN(n20495) );
  INV_X1 U29846 ( .A(n20495), .ZN(n19355) );
  NOR2_X1 U29847 ( .A1(n21458), .A2(n21462), .ZN(n19354) );
  NOR2_X1 U29848 ( .A1(n19355), .A2(n19354), .ZN(n19368) );
  INV_X1 U29849 ( .A(n19356), .ZN(n19358) );
  OAI21_X1 U29850 ( .B1(n19363), .B2(n19359), .A(n767), .ZN(n19360) );
  NAND3_X1 U29851 ( .A1(n19361), .A2(n21449), .A3(n19360), .ZN(n19367) );
  NAND2_X1 U29852 ( .A1(n19362), .A2(n21460), .ZN(n20490) );
  INV_X1 U29853 ( .A(n20490), .ZN(n21457) );
  OAI22_X1 U29854 ( .A1(n19363), .A2(n21464), .B1(n21469), .B2(n20314), .ZN(
        n19365) );
  OAI21_X1 U29855 ( .B1(n21457), .B2(n19365), .A(n19364), .ZN(n19366) );
  AND2_X1 U29856 ( .A1(n21887), .A2(n22857), .ZN(n22866) );
  OAI21_X1 U29857 ( .B1(n22849), .B2(n22866), .A(n22844), .ZN(n19403) );
  NAND3_X1 U29858 ( .A1(n20462), .A2(n20477), .A3(n20389), .ZN(n19374) );
  NAND4_X1 U29859 ( .A1(n19372), .A2(n19371), .A3(n19370), .A4(n20477), .ZN(
        n19373) );
  AND2_X1 U29860 ( .A1(n19374), .A2(n19373), .ZN(n19379) );
  INV_X1 U29861 ( .A(n20389), .ZN(n20461) );
  INV_X1 U29863 ( .A(n19380), .ZN(n19383) );
  INV_X1 U29864 ( .A(n20473), .ZN(n20479) );
  AOI21_X1 U29866 ( .B1(n19383), .B2(n19382), .A(n19381), .ZN(n19384) );
  OAI21_X1 U29867 ( .B1(n19387), .B2(n18023), .A(n19386), .ZN(n19394) );
  NAND2_X1 U29868 ( .A1(n19389), .A2(n19388), .ZN(n19391) );
  OAI21_X1 U29869 ( .B1(n19400), .B2(n19399), .A(n19398), .ZN(n19401) );
  NOR2_X1 U29870 ( .A1(n17469), .A2(n19405), .ZN(n19406) );
  NAND2_X1 U29871 ( .A1(n19411), .A2(n8378), .ZN(n19407) );
  NAND3_X1 U29873 ( .A1(n19412), .A2(n19411), .A3(n19423), .ZN(n19421) );
  INV_X1 U29874 ( .A(n19413), .ZN(n19415) );
  OAI21_X1 U29875 ( .B1(n19415), .B2(n8378), .A(n6332), .ZN(n19416) );
  NAND2_X1 U29876 ( .A1(n19416), .A2(n19426), .ZN(n19420) );
  NAND3_X1 U29877 ( .A1(n2222), .A2(n19418), .A3(n19417), .ZN(n19419) );
  INV_X1 U29878 ( .A(n19422), .ZN(n19431) );
  INV_X1 U29879 ( .A(n19423), .ZN(n19430) );
  OAI211_X1 U29881 ( .C1(n19431), .C2(n19430), .A(n19429), .B(n19428), .ZN(
        n19432) );
  INV_X1 U29882 ( .A(n19432), .ZN(n19435) );
  AND2_X1 U29883 ( .A1(n22856), .A2(n4413), .ZN(n21015) );
  AOI21_X1 U29884 ( .B1(n19436), .B2(n22328), .A(n21015), .ZN(n19440) );
  OAI21_X1 U29885 ( .B1(n19603), .B2(n22857), .A(n22859), .ZN(n19438) );
  NAND2_X1 U29886 ( .A1(n22856), .A2(n22857), .ZN(n19604) );
  OAI21_X1 U29887 ( .B1(n21885), .B2(n22859), .A(n19604), .ZN(n19437) );
  NOR2_X1 U29888 ( .A1(n23982), .A2(n23992), .ZN(n22416) );
  NAND2_X1 U29889 ( .A1(n22416), .A2(n22426), .ZN(n19442) );
  AND2_X1 U29890 ( .A1(n19442), .A2(n23037), .ZN(n19444) );
  NAND2_X1 U29891 ( .A1(n23989), .A2(n23981), .ZN(n19443) );
  MUX2_X1 U29892 ( .A(n19444), .B(n19443), .S(n23998), .Z(n19451) );
  NOR2_X1 U29893 ( .A1(n23992), .A2(n24000), .ZN(n19445) );
  NOR2_X1 U29894 ( .A1(n22428), .A2(n19445), .ZN(n19446) );
  NOR2_X1 U29895 ( .A1(n22426), .A2(n24000), .ZN(n22430) );
  NAND2_X1 U29896 ( .A1(n23987), .A2(n23992), .ZN(n23027) );
  OAI22_X1 U29897 ( .A1(n23991), .A2(n19446), .B1(n22430), .B2(n23027), .ZN(
        n19450) );
  NAND2_X1 U29898 ( .A1(n19447), .A2(n23028), .ZN(n19449) );
  INV_X1 U29899 ( .A(n23028), .ZN(n23990) );
  NAND4_X1 U29900 ( .A1(n19451), .A2(n19450), .A3(n19449), .A4(n19448), .ZN(
        n23840) );
  INV_X1 U29901 ( .A(n23840), .ZN(n28424) );
  NOR2_X1 U29902 ( .A1(n19774), .A2(n21276), .ZN(n21263) );
  AOI21_X1 U29903 ( .B1(n19452), .B2(n19777), .A(n51013), .ZN(n19454) );
  OAI211_X1 U29904 ( .C1(n21263), .C2(n21271), .A(n19454), .B(n19453), .ZN(
        n19458) );
  NOR2_X1 U29905 ( .A1(n19459), .A2(n51013), .ZN(n19788) );
  NAND3_X1 U29906 ( .A1(n19788), .A2(n19775), .A3(n21269), .ZN(n19457) );
  AND2_X1 U29907 ( .A1(n19455), .A2(n51013), .ZN(n21264) );
  NAND3_X1 U29908 ( .A1(n21264), .A2(n19777), .A3(n19779), .ZN(n19456) );
  NAND2_X1 U29909 ( .A1(n19462), .A2(n51013), .ZN(n21284) );
  AND2_X1 U29910 ( .A1(n19019), .A2(n19777), .ZN(n21268) );
  NAND2_X1 U29911 ( .A1(n21268), .A2(n19778), .ZN(n19460) );
  MUX2_X1 U29912 ( .A(n21284), .B(n19460), .S(n19459), .Z(n19470) );
  INV_X1 U29913 ( .A(n19461), .ZN(n19463) );
  NAND3_X1 U29915 ( .A1(n19473), .A2(n19472), .A3(n19482), .ZN(n19485) );
  NAND3_X1 U29916 ( .A1(n19475), .A2(n3335), .A3(n19474), .ZN(n19476) );
  NAND2_X1 U29917 ( .A1(n19476), .A2(n21253), .ZN(n19481) );
  NOR2_X1 U29918 ( .A1(n19477), .A2(n51132), .ZN(n19479) );
  OAI21_X1 U29919 ( .B1(n21245), .B2(n19479), .A(n19478), .ZN(n19480) );
  NAND2_X1 U29920 ( .A1(n19481), .A2(n19480), .ZN(n19484) );
  NOR2_X1 U29921 ( .A1(n19487), .A2(n16218), .ZN(n19489) );
  OAI21_X1 U29922 ( .B1(n19490), .B2(n19489), .A(n19488), .ZN(n19497) );
  NAND2_X1 U29924 ( .A1(n20082), .A2(n20062), .ZN(n20054) );
  NAND2_X1 U29925 ( .A1(n20072), .A2(n20054), .ZN(n19492) );
  OAI211_X1 U29926 ( .C1(n19494), .C2(n19493), .A(n19492), .B(n20078), .ZN(
        n19495) );
  NAND4_X1 U29927 ( .A1(n19498), .A2(n19497), .A3(n19496), .A4(n19495), .ZN(
        n19502) );
  NAND2_X1 U29928 ( .A1(n19500), .A2(n19499), .ZN(n20083) );
  NOR2_X1 U29929 ( .A1(n20083), .A2(n20073), .ZN(n19501) );
  NAND2_X1 U29930 ( .A1(n6226), .A2(n19503), .ZN(n19507) );
  NAND2_X1 U29931 ( .A1(n19505), .A2(n21227), .ZN(n19506) );
  OAI211_X1 U29932 ( .C1(n19508), .C2(n19507), .A(n21229), .B(n19506), .ZN(
        n19516) );
  NAND3_X1 U29933 ( .A1(n19520), .A2(n19510), .A3(n19509), .ZN(n19511) );
  INV_X1 U29935 ( .A(n19549), .ZN(n19550) );
  MUX2_X1 U29936 ( .A(n8311), .B(n19528), .S(n21180), .Z(n19533) );
  NAND4_X1 U29937 ( .A1(n19524), .A2(n19523), .A3(n19522), .A4(n8311), .ZN(
        n19532) );
  NAND3_X1 U29938 ( .A1(n19526), .A2(n51434), .A3(n19525), .ZN(n19531) );
  OAI211_X1 U29939 ( .C1(n19702), .C2(n8311), .A(n19528), .B(n19527), .ZN(
        n19530) );
  OAI21_X1 U29940 ( .B1(n20158), .B2(n19534), .A(n20124), .ZN(n19539) );
  NOR2_X1 U29941 ( .A1(n19535), .A2(n20157), .ZN(n19536) );
  AOI22_X1 U29944 ( .A1(n19541), .A2(n19540), .B1(n20158), .B2(n20125), .ZN(
        n19547) );
  OAI211_X1 U29945 ( .C1(n19545), .C2(n19544), .A(n19543), .B(n19542), .ZN(
        n19546) );
  OAI21_X1 U29946 ( .B1(n22018), .B2(n19550), .A(n22003), .ZN(n22583) );
  OAI21_X1 U29947 ( .B1(n22587), .B2(n20903), .A(n22593), .ZN(n19551) );
  NAND2_X1 U29948 ( .A1(n22583), .A2(n19551), .ZN(n19558) );
  INV_X1 U29949 ( .A(n19554), .ZN(n23438) );
  INV_X1 U29950 ( .A(n22593), .ZN(n22023) );
  AOI22_X1 U29951 ( .A1(n22012), .A2(n23438), .B1(n22021), .B2(n22584), .ZN(
        n19557) );
  INV_X1 U29952 ( .A(n23446), .ZN(n22011) );
  AND2_X1 U29953 ( .A1(n23445), .A2(n22586), .ZN(n22004) );
  OAI211_X1 U29954 ( .C1(n22023), .C2(n22011), .A(n21318), .B(n22004), .ZN(
        n19553) );
  NAND3_X1 U29956 ( .A1(n22589), .A2(n23436), .A3(n19554), .ZN(n19552) );
  NAND2_X1 U29957 ( .A1(n19555), .A2(n23434), .ZN(n19556) );
  XNOR2_X1 U29958 ( .A(n28424), .B(n26044), .ZN(n19586) );
  NOR2_X1 U29959 ( .A1(n50991), .A2(n22140), .ZN(n22151) );
  MUX2_X1 U29960 ( .A(n19559), .B(n19562), .S(n21025), .Z(n19572) );
  INV_X1 U29962 ( .A(n22155), .ZN(n21027) );
  XNOR2_X1 U29963 ( .A(n51660), .B(n21027), .ZN(n19567) );
  OR2_X1 U29964 ( .A1(n50992), .A2(n22155), .ZN(n20956) );
  INV_X1 U29965 ( .A(n20956), .ZN(n19564) );
  NAND3_X1 U29966 ( .A1(n19565), .A2(n50991), .A3(n22157), .ZN(n19566) );
  AND2_X1 U29967 ( .A1(n50991), .A2(n22155), .ZN(n22141) );
  OAI21_X1 U29968 ( .B1(n52381), .B2(n19568), .A(n22141), .ZN(n19569) );
  NAND2_X1 U29969 ( .A1(n22916), .A2(n22918), .ZN(n22350) );
  INV_X1 U29970 ( .A(n22367), .ZN(n19578) );
  NAND2_X1 U29971 ( .A1(n19578), .A2(n2175), .ZN(n19573) );
  AOI21_X1 U29972 ( .B1(n22360), .B2(n19573), .A(n22349), .ZN(n19574) );
  NOR2_X1 U29973 ( .A1(n19575), .A2(n19574), .ZN(n19585) );
  NOR2_X1 U29974 ( .A1(n22165), .A2(n19577), .ZN(n21036) );
  INV_X1 U29975 ( .A(n21036), .ZN(n19584) );
  NOR2_X1 U29976 ( .A1(n19578), .A2(n22919), .ZN(n21038) );
  AND2_X1 U29977 ( .A1(n22901), .A2(n22918), .ZN(n22168) );
  INV_X1 U29978 ( .A(n22168), .ZN(n19579) );
  AOI21_X1 U29979 ( .B1(n22363), .B2(n21038), .A(n19579), .ZN(n19580) );
  OAI211_X1 U29980 ( .C1(n22167), .C2(n22165), .A(n19580), .B(n22914), .ZN(
        n19583) );
  AOI21_X1 U29981 ( .B1(n22362), .B2(n22918), .A(n22167), .ZN(n19581) );
  OR2_X1 U29982 ( .A1(n19581), .A2(n22902), .ZN(n19582) );
  XNOR2_X1 U29983 ( .A(n751), .B(n19586), .ZN(n19628) );
  INV_X1 U29984 ( .A(n23469), .ZN(n19587) );
  NAND2_X1 U29985 ( .A1(n19587), .A2(n21947), .ZN(n19601) );
  NAND2_X1 U29987 ( .A1(n21962), .A2(n23154), .ZN(n19588) );
  AOI22_X1 U29988 ( .A1(n19589), .A2(n19588), .B1(n23156), .B2(n23154), .ZN(
        n19600) );
  NAND3_X1 U29989 ( .A1(n19591), .A2(n23464), .A3(n19590), .ZN(n19594) );
  NOR2_X1 U29990 ( .A1(n21957), .A2(n21947), .ZN(n21950) );
  NAND3_X1 U29991 ( .A1(n19592), .A2(n21950), .A3(n6010), .ZN(n19593) );
  NOR2_X1 U29993 ( .A1(n23153), .A2(n23157), .ZN(n19595) );
  NAND2_X1 U29994 ( .A1(n51250), .A2(n19595), .ZN(n19597) );
  AND2_X1 U29995 ( .A1(n21167), .A2(n19597), .ZN(n19598) );
  NAND2_X1 U29996 ( .A1(n22861), .A2(n21887), .ZN(n19602) );
  INV_X1 U29997 ( .A(n19610), .ZN(n19606) );
  INV_X1 U29998 ( .A(n19604), .ZN(n22327) );
  OAI211_X1 U29999 ( .C1(n22849), .C2(n22864), .A(n4413), .B(n21887), .ZN(
        n19605) );
  OAI211_X1 U30000 ( .C1(n22334), .C2(n19606), .A(n22327), .B(n19605), .ZN(
        n19607) );
  OAI21_X1 U30001 ( .B1(n19608), .B2(n22851), .A(n19607), .ZN(n19619) );
  NAND3_X1 U30002 ( .A1(n19611), .A2(n23020), .A3(n22857), .ZN(n19617) );
  NAND3_X1 U30003 ( .A1(n19611), .A2(n22859), .A3(n23020), .ZN(n19615) );
  OAI21_X1 U30004 ( .B1(n21885), .B2(n22857), .A(n4413), .ZN(n19613) );
  NAND2_X1 U30005 ( .A1(n19613), .A2(n19612), .ZN(n19614) );
  NAND4_X1 U30006 ( .A1(n19617), .A2(n19616), .A3(n19615), .A4(n19614), .ZN(
        n19618) );
  XNOR2_X1 U30007 ( .A(n25213), .B(n25747), .ZN(n19627) );
  AND2_X1 U30008 ( .A1(n23483), .A2(n23479), .ZN(n19620) );
  NAND2_X1 U30009 ( .A1(n8076), .A2(n2130), .ZN(n20995) );
  INV_X1 U30010 ( .A(n20995), .ZN(n19624) );
  NAND3_X1 U30011 ( .A1(n23485), .A2(n21970), .A3(n21975), .ZN(n19623) );
  XNOR2_X1 U30012 ( .A(n23480), .B(n21975), .ZN(n19621) );
  AOI21_X1 U30013 ( .B1(n23489), .B2(n23477), .A(n19621), .ZN(n19622) );
  NAND4_X1 U30015 ( .A1(n23485), .A2(n21970), .A3(n21987), .A4(n23481), .ZN(
        n20999) );
  NAND2_X1 U30016 ( .A1(n21983), .A2(n21970), .ZN(n19625) );
  OR2_X1 U30018 ( .A1(n19886), .A2(n19894), .ZN(n19631) );
  NAND2_X1 U30019 ( .A1(n19886), .A2(n19887), .ZN(n19630) );
  MUX2_X1 U30020 ( .A(n19631), .B(n19630), .S(n19897), .Z(n19634) );
  NAND2_X1 U30021 ( .A1(n19898), .A2(n19632), .ZN(n19633) );
  MUX2_X1 U30022 ( .A(n19884), .B(n19886), .S(n19636), .Z(n19638) );
  NOR2_X1 U30023 ( .A1(n19707), .A2(n19708), .ZN(n19656) );
  MUX2_X1 U30024 ( .A(n19643), .B(n19639), .S(n19647), .Z(n19641) );
  NOR2_X1 U30025 ( .A1(n19641), .A2(n19640), .ZN(n19651) );
  INV_X1 U30026 ( .A(n19642), .ZN(n19644) );
  NAND3_X1 U30027 ( .A1(n19645), .A2(n19644), .A3(n19643), .ZN(n19646) );
  MUX2_X1 U30028 ( .A(n19650), .B(n19649), .S(n19648), .Z(n19742) );
  INV_X1 U30029 ( .A(n19651), .ZN(n19654) );
  INV_X1 U30030 ( .A(n19652), .ZN(n19653) );
  NAND3_X1 U30031 ( .A1(n19654), .A2(n19653), .A3(n19744), .ZN(n19655) );
  OAI21_X1 U30032 ( .B1(n19743), .B2(n19742), .A(n19655), .ZN(n19698) );
  NOR2_X1 U30033 ( .A1(n19656), .A2(n19698), .ZN(n22728) );
  OAI211_X1 U30034 ( .C1(n19663), .C2(n19662), .A(n19891), .B(n19893), .ZN(
        n19667) );
  AOI22_X1 U30036 ( .A1(n19675), .A2(n18236), .B1(n19674), .B2(n4681), .ZN(
        n19677) );
  INV_X1 U30037 ( .A(n19689), .ZN(n19684) );
  MUX2_X1 U30038 ( .A(n19679), .B(n775), .S(n51006), .Z(n19683) );
  OAI21_X1 U30039 ( .B1(n19684), .B2(n19683), .A(n19682), .ZN(n19686) );
  NAND2_X1 U30040 ( .A1(n19686), .A2(n19685), .ZN(n19695) );
  AOI22_X1 U30042 ( .A1(n19690), .A2(n19689), .B1(n20209), .B2(n19691), .ZN(
        n19694) );
  NAND3_X1 U30043 ( .A1(n20217), .A2(n20212), .A3(n19691), .ZN(n19692) );
  OAI21_X1 U30044 ( .B1(n19698), .B2(n19709), .A(n5370), .ZN(n22735) );
  OR2_X1 U30045 ( .A1(n22728), .A2(n22735), .ZN(n20574) );
  NAND2_X1 U30046 ( .A1(n20574), .A2(n23814), .ZN(n20581) );
  NAND2_X1 U30047 ( .A1(n5371), .A2(n23814), .ZN(n22374) );
  INV_X1 U30048 ( .A(n19797), .ZN(n21291) );
  OAI22_X1 U30049 ( .A1(n19712), .A2(n7874), .B1(n19711), .B2(n21291), .ZN(
        n21308) );
  NAND3_X1 U30050 ( .A1(n21291), .A2(n19713), .A3(n509), .ZN(n19714) );
  AND2_X1 U30051 ( .A1(n19714), .A2(n19715), .ZN(n19724) );
  NAND2_X1 U30052 ( .A1(n19716), .A2(n19800), .ZN(n19719) );
  OAI211_X1 U30053 ( .C1(n19796), .C2(n21304), .A(n18217), .B(n19801), .ZN(
        n19717) );
  NAND2_X1 U30054 ( .A1(n21305), .A2(n19717), .ZN(n19718) );
  MUX2_X1 U30055 ( .A(n21293), .B(n19721), .S(n509), .Z(n19722) );
  OAI21_X1 U30056 ( .B1(n19722), .B2(n21296), .A(n19792), .ZN(n19723) );
  NAND2_X1 U30057 ( .A1(n22374), .A2(n22375), .ZN(n22384) );
  NOR2_X1 U30058 ( .A1(n19726), .A2(n19725), .ZN(n19810) );
  INV_X1 U30059 ( .A(n19810), .ZN(n19728) );
  NAND2_X1 U30060 ( .A1(n21212), .A2(n6078), .ZN(n19729) );
  OR2_X1 U30061 ( .A1(n19727), .A2(n19729), .ZN(n19812) );
  NAND2_X1 U30062 ( .A1(n19728), .A2(n19812), .ZN(n19741) );
  INV_X1 U30063 ( .A(n21208), .ZN(n19815) );
  NAND2_X1 U30064 ( .A1(n19815), .A2(n21214), .ZN(n19740) );
  INV_X1 U30065 ( .A(n19729), .ZN(n19821) );
  NAND2_X1 U30066 ( .A1(n21200), .A2(n19822), .ZN(n19730) );
  OAI211_X1 U30067 ( .C1(n21215), .C2(n19821), .A(n19814), .B(n19730), .ZN(
        n19731) );
  NAND2_X1 U30068 ( .A1(n19731), .A2(n19813), .ZN(n19738) );
  NAND4_X1 U30069 ( .A1(n19733), .A2(n19809), .A3(n21213), .A4(n19823), .ZN(
        n19736) );
  NAND2_X1 U30070 ( .A1(n19734), .A2(n19822), .ZN(n19735) );
  NAND4_X1 U30071 ( .A1(n19738), .A2(n19737), .A3(n19736), .A4(n19735), .ZN(
        n19739) );
  NAND2_X1 U30073 ( .A1(n353), .A2(n50977), .ZN(n22377) );
  NOR2_X1 U30074 ( .A1(n22377), .A2(n22740), .ZN(n22395) );
  OAI21_X1 U30075 ( .B1(n20581), .B2(n22384), .A(n19745), .ZN(n23820) );
  NAND2_X1 U30076 ( .A1(n5095), .A2(n22390), .ZN(n19749) );
  NAND2_X1 U30077 ( .A1(n753), .A2(n50976), .ZN(n19746) );
  NAND2_X1 U30078 ( .A1(n22386), .A2(n19746), .ZN(n19747) );
  AOI22_X1 U30079 ( .A1(n22739), .A2(n51753), .B1(n19748), .B2(n19747), .ZN(
        n23818) );
  INV_X1 U30080 ( .A(n19749), .ZN(n23812) );
  NAND2_X1 U30081 ( .A1(n23812), .A2(n51753), .ZN(n19751) );
  NAND3_X1 U30082 ( .A1(n23813), .A2(n23814), .A3(n22741), .ZN(n19750) );
  MUX2_X1 U30083 ( .A(n19751), .B(n19750), .S(n22736), .Z(n19752) );
  NAND2_X1 U30084 ( .A1(n23818), .A2(n19752), .ZN(n19753) );
  OR2_X1 U30085 ( .A1(n23820), .A2(n19753), .ZN(n25929) );
  NAND2_X1 U30086 ( .A1(n22995), .A2(n22557), .ZN(n20918) );
  OAI21_X1 U30087 ( .B1(n22434), .B2(n20918), .A(n19755), .ZN(n19756) );
  OAI21_X1 U30088 ( .B1(n22555), .B2(n19756), .A(n22983), .ZN(n19767) );
  OAI21_X1 U30089 ( .B1(n22990), .B2(n22978), .A(n19758), .ZN(n19760) );
  INV_X1 U30090 ( .A(n19762), .ZN(n19759) );
  NAND3_X1 U30091 ( .A1(n19760), .A2(n22989), .A3(n19759), .ZN(n19765) );
  NOR2_X1 U30092 ( .A1(n19761), .A2(n22995), .ZN(n19763) );
  OAI21_X1 U30093 ( .B1(n22999), .B2(n19763), .A(n19762), .ZN(n19764) );
  XNOR2_X1 U30094 ( .A(n19768), .B(n25640), .ZN(n19771) );
  INV_X1 U30095 ( .A(n19769), .ZN(n19770) );
  XNOR2_X1 U30096 ( .A(n19771), .B(n19770), .ZN(n42433) );
  XNOR2_X1 U30097 ( .A(n42433), .B(n43692), .ZN(n19772) );
  XNOR2_X1 U30098 ( .A(n25320), .B(n19772), .ZN(n19773) );
  XNOR2_X1 U30099 ( .A(n19773), .B(n25929), .ZN(n19922) );
  OAI21_X1 U30100 ( .B1(n19776), .B2(n21269), .A(n19785), .ZN(n21262) );
  NAND2_X1 U30101 ( .A1(n21287), .A2(n19777), .ZN(n21279) );
  NAND3_X1 U30102 ( .A1(n21262), .A2(n21270), .A3(n21279), .ZN(n19781) );
  NAND3_X1 U30103 ( .A1(n19779), .A2(n19782), .A3(n19778), .ZN(n19780) );
  NOR2_X1 U30104 ( .A1(n19785), .A2(n19784), .ZN(n19787) );
  OAI21_X1 U30105 ( .B1(n19788), .B2(n19787), .A(n19786), .ZN(n19789) );
  INV_X1 U30106 ( .A(n19901), .ZN(n22876) );
  NAND2_X1 U30107 ( .A1(n19796), .A2(n19795), .ZN(n21301) );
  OAI21_X1 U30108 ( .B1(n21301), .B2(n21300), .A(n19797), .ZN(n19802) );
  XNOR2_X1 U30109 ( .A(n509), .B(n7874), .ZN(n19798) );
  OAI21_X1 U30111 ( .B1(n19800), .B2(n19799), .A(n509), .ZN(n19803) );
  OAI21_X1 U30112 ( .B1(n19803), .B2(n19802), .A(n19801), .ZN(n19804) );
  AND2_X1 U30113 ( .A1(n22876), .A2(n23101), .ZN(n22890) );
  NAND2_X1 U30114 ( .A1(n19808), .A2(n19807), .ZN(n19811) );
  OAI21_X1 U30115 ( .B1(n19812), .B2(n21197), .A(n21218), .ZN(n19818) );
  NAND2_X1 U30116 ( .A1(n19813), .A2(n2229), .ZN(n19816) );
  OAI22_X1 U30117 ( .A1(n19816), .A2(n19815), .B1(n19814), .B2(n21213), .ZN(
        n19817) );
  OAI21_X1 U30118 ( .B1(n19823), .B2(n21213), .A(n19822), .ZN(n19824) );
  NOR2_X1 U30119 ( .A1(n19826), .A2(n21188), .ZN(n19827) );
  NAND4_X1 U30120 ( .A1(n19828), .A2(n21186), .A3(n19827), .A4(n17201), .ZN(
        n19830) );
  NAND2_X1 U30122 ( .A1(n19833), .A2(n19832), .ZN(n19845) );
  NAND4_X1 U30123 ( .A1(n19834), .A2(n21173), .A3(n21181), .A4(n21185), .ZN(
        n19835) );
  OAI21_X1 U30124 ( .B1(n21172), .B2(n21186), .A(n19835), .ZN(n19836) );
  INV_X1 U30125 ( .A(n19836), .ZN(n19844) );
  OAI211_X1 U30126 ( .C1(n51434), .C2(n21178), .A(n21180), .B(n19838), .ZN(
        n19843) );
  NAND3_X1 U30127 ( .A1(n19841), .A2(n21185), .A3(n19840), .ZN(n19842) );
  NAND4_X1 U30128 ( .A1(n19845), .A2(n19844), .A3(n19843), .A4(n19842), .ZN(
        n22875) );
  NOR2_X1 U30129 ( .A1(n25056), .A2(n51654), .ZN(n23099) );
  NAND2_X1 U30130 ( .A1(n19861), .A2(n19850), .ZN(n19856) );
  NAND2_X1 U30131 ( .A1(n19852), .A2(n19851), .ZN(n19855) );
  NAND2_X1 U30132 ( .A1(n19853), .A2(n585), .ZN(n19854) );
  NAND4_X1 U30133 ( .A1(n19857), .A2(n19856), .A3(n19855), .A4(n19854), .ZN(
        n19859) );
  NAND2_X1 U30134 ( .A1(n19859), .A2(n19858), .ZN(n19880) );
  NOR2_X1 U30135 ( .A1(n585), .A2(n19873), .ZN(n19862) );
  AOI22_X1 U30136 ( .A1(n19862), .A2(n19874), .B1(n51039), .B2(n19861), .ZN(
        n19879) );
  OAI21_X1 U30137 ( .B1(n19865), .B2(n19864), .A(n19863), .ZN(n19877) );
  NOR2_X1 U30138 ( .A1(n19867), .A2(n19866), .ZN(n19876) );
  NAND3_X1 U30139 ( .A1(n19870), .A2(n19869), .A3(n51039), .ZN(n19872) );
  OAI211_X1 U30140 ( .C1(n19874), .C2(n19873), .A(n19872), .B(n19871), .ZN(
        n19875) );
  OAI21_X1 U30141 ( .B1(n19877), .B2(n19876), .A(n19875), .ZN(n19878) );
  INV_X1 U30142 ( .A(n25056), .ZN(n23100) );
  NAND2_X1 U30143 ( .A1(n22876), .A2(n52174), .ZN(n22772) );
  INV_X1 U30144 ( .A(n23101), .ZN(n22884) );
  NAND3_X1 U30145 ( .A1(n22772), .A2(n22884), .A3(n7806), .ZN(n19881) );
  NAND2_X1 U30146 ( .A1(n25056), .A2(n52175), .ZN(n19904) );
  NAND4_X1 U30147 ( .A1(n19883), .A2(n19882), .A3(n19881), .A4(n19904), .ZN(
        n19900) );
  OAI211_X1 U30148 ( .C1(n19885), .C2(n19887), .A(n19889), .B(n19884), .ZN(
        n19888) );
  NAND3_X1 U30149 ( .A1(n19896), .A2(n19895), .A3(n19894), .ZN(n19899) );
  NAND2_X1 U30150 ( .A1(n25057), .A2(n51654), .ZN(n19906) );
  NOR2_X1 U30151 ( .A1(n23101), .A2(n52174), .ZN(n23098) );
  NAND2_X1 U30152 ( .A1(n19906), .A2(n23098), .ZN(n19903) );
  NAND3_X1 U30153 ( .A1(n22763), .A2(n25057), .A3(n23101), .ZN(n19902) );
  INV_X1 U30154 ( .A(n19904), .ZN(n19905) );
  NAND2_X1 U30155 ( .A1(n22890), .A2(n19905), .ZN(n19909) );
  INV_X1 U30156 ( .A(n19906), .ZN(n19907) );
  NAND2_X1 U30157 ( .A1(n19907), .A2(n52174), .ZN(n19908) );
  XNOR2_X1 U30158 ( .A(n25927), .B(n43691), .ZN(n19921) );
  NAND2_X1 U30159 ( .A1(n7119), .A2(n21714), .ZN(n21699) );
  NAND4_X1 U30160 ( .A1(n7119), .A2(n21713), .A3(n22184), .A4(n52048), .ZN(
        n19911) );
  OAI22_X1 U30161 ( .A1(n21699), .A2(n20568), .B1(n19911), .B2(n22186), .ZN(
        n19912) );
  INV_X1 U30162 ( .A(n19912), .ZN(n19920) );
  INV_X1 U30163 ( .A(n21104), .ZN(n22185) );
  NOR2_X1 U30164 ( .A1(n21700), .A2(n52048), .ZN(n21710) );
  INV_X1 U30165 ( .A(n19914), .ZN(n19913) );
  OAI211_X1 U30166 ( .C1(n21710), .C2(n21712), .A(n19913), .B(n463), .ZN(
        n19919) );
  INV_X1 U30167 ( .A(n21716), .ZN(n19915) );
  OAI211_X1 U30168 ( .C1(n22178), .C2(n52048), .A(n19915), .B(n19914), .ZN(
        n19918) );
  XNOR2_X1 U30169 ( .A(n19921), .B(n27177), .ZN(n23850) );
  XNOR2_X1 U30170 ( .A(n23850), .B(n19922), .ZN(n19923) );
  NAND2_X1 U30171 ( .A1(n21355), .A2(n21601), .ZN(n19924) );
  OAI211_X1 U30172 ( .C1(n20758), .C2(n21604), .A(n20760), .B(n19924), .ZN(
        n19929) );
  NOR2_X1 U30173 ( .A1(n21362), .A2(n21364), .ZN(n19925) );
  OAI211_X1 U30174 ( .C1(n21349), .C2(n19925), .A(n762), .B(n21359), .ZN(
        n19928) );
  NAND4_X1 U30175 ( .A1(n19929), .A2(n19928), .A3(n19927), .A4(n19926), .ZN(
        n19932) );
  AOI21_X1 U30176 ( .B1(n19930), .B2(n21591), .A(n21604), .ZN(n19931) );
  OR2_X2 U30177 ( .A1(n19932), .A2(n19931), .ZN(n24034) );
  NAND2_X1 U30178 ( .A1(n19933), .A2(n20745), .ZN(n19934) );
  NAND2_X1 U30179 ( .A1(n19934), .A2(n18495), .ZN(n19938) );
  NAND3_X1 U30180 ( .A1(n20746), .A2(n21547), .A3(n20745), .ZN(n19937) );
  NAND3_X1 U30181 ( .A1(n51485), .A2(n20627), .A3(n20201), .ZN(n19935) );
  INV_X1 U30182 ( .A(n20746), .ZN(n20193) );
  NAND3_X1 U30183 ( .A1(n20752), .A2(n21537), .A3(n21544), .ZN(n19940) );
  INV_X1 U30184 ( .A(n24030), .ZN(n22107) );
  NOR2_X1 U30185 ( .A1(n24034), .A2(n5204), .ZN(n20005) );
  NOR2_X1 U30186 ( .A1(n21421), .A2(n52139), .ZN(n19944) );
  AOI21_X1 U30187 ( .B1(n19944), .B2(n20840), .A(n19943), .ZN(n19946) );
  NAND3_X1 U30189 ( .A1(n20841), .A2(n21435), .A3(n20839), .ZN(n19949) );
  NAND3_X1 U30190 ( .A1(n20329), .A2(n21426), .A3(n21420), .ZN(n19948) );
  AND2_X1 U30191 ( .A1(n19949), .A2(n19948), .ZN(n19963) );
  OAI211_X1 U30192 ( .C1(n21420), .C2(n20327), .A(n19950), .B(n21435), .ZN(
        n19954) );
  OAI21_X1 U30193 ( .B1(n21442), .B2(n21424), .A(n3493), .ZN(n19951) );
  AOI21_X1 U30194 ( .B1(n19951), .B2(n52139), .A(n21421), .ZN(n19953) );
  OAI211_X1 U30195 ( .C1(n20325), .C2(n21442), .A(n21424), .B(n52139), .ZN(
        n19952) );
  NAND3_X1 U30196 ( .A1(n19954), .A2(n19953), .A3(n19952), .ZN(n19962) );
  NOR2_X1 U30197 ( .A1(n20322), .A2(n19955), .ZN(n20330) );
  INV_X1 U30198 ( .A(n20322), .ZN(n21429) );
  NAND2_X1 U30199 ( .A1(n21429), .A2(n20838), .ZN(n19960) );
  INV_X1 U30200 ( .A(n19956), .ZN(n19958) );
  OAI211_X1 U30201 ( .C1(n19958), .C2(n21442), .A(n20838), .B(n19957), .ZN(
        n19959) );
  OAI211_X1 U30202 ( .C1(n20330), .C2(n20838), .A(n19960), .B(n19959), .ZN(
        n19961) );
  INV_X1 U30203 ( .A(n22101), .ZN(n23392) );
  INV_X1 U30204 ( .A(n24043), .ZN(n19976) );
  NAND3_X1 U30205 ( .A1(n21492), .A2(n20451), .A3(n21485), .ZN(n20833) );
  OAI211_X1 U30206 ( .C1(n51754), .C2(n21480), .A(n19967), .B(n20833), .ZN(
        n19968) );
  INV_X1 U30207 ( .A(n19968), .ZN(n19975) );
  INV_X1 U30208 ( .A(n21485), .ZN(n19970) );
  AND2_X1 U30209 ( .A1(n2220), .A2(n20825), .ZN(n20820) );
  NOR2_X1 U30210 ( .A1(n20820), .A2(n20812), .ZN(n19972) );
  NAND2_X1 U30211 ( .A1(n20451), .A2(n21480), .ZN(n20818) );
  OR2_X1 U30212 ( .A1(n20818), .A2(n20811), .ZN(n20454) );
  NOR2_X1 U30213 ( .A1(n20336), .A2(n20441), .ZN(n21496) );
  INV_X1 U30214 ( .A(n20826), .ZN(n21482) );
  OAI21_X1 U30215 ( .B1(n21496), .B2(n21482), .A(n20829), .ZN(n19974) );
  INV_X1 U30216 ( .A(n24041), .ZN(n22575) );
  MUX2_X1 U30217 ( .A(n19976), .B(n23393), .S(n22575), .Z(n20009) );
  NAND2_X1 U30218 ( .A1(n24041), .A2(n24030), .ZN(n23664) );
  NAND2_X1 U30219 ( .A1(n20258), .A2(n19981), .ZN(n20251) );
  NOR2_X1 U30220 ( .A1(n20251), .A2(n21637), .ZN(n21628) );
  INV_X1 U30221 ( .A(n19977), .ZN(n21636) );
  NAND2_X1 U30222 ( .A1(n21628), .A2(n21636), .ZN(n19986) );
  NAND2_X1 U30223 ( .A1(n19978), .A2(n21633), .ZN(n19980) );
  NAND2_X1 U30224 ( .A1(n20698), .A2(n20244), .ZN(n20254) );
  AOI21_X1 U30225 ( .B1(n20241), .B2(n20254), .A(n21637), .ZN(n19979) );
  AND3_X1 U30226 ( .A1(n21622), .A2(n21632), .A3(n21614), .ZN(n19983) );
  XNOR2_X1 U30227 ( .A(n19981), .B(n21613), .ZN(n19982) );
  AOI22_X1 U30228 ( .A1(n19983), .A2(n19982), .B1(n20253), .B2(n20259), .ZN(
        n19985) );
  INV_X1 U30229 ( .A(n23670), .ZN(n20001) );
  NAND2_X1 U30230 ( .A1(n21555), .A2(n21412), .ZN(n19988) );
  AOI21_X1 U30231 ( .B1(n21556), .B2(n21412), .A(n21560), .ZN(n19987) );
  INV_X1 U30233 ( .A(n21576), .ZN(n19992) );
  OAI21_X1 U30234 ( .B1(n19987), .B2(n19992), .A(n21558), .ZN(n19991) );
  NAND2_X1 U30235 ( .A1(n21556), .A2(n21584), .ZN(n20605) );
  NAND3_X1 U30236 ( .A1(n19992), .A2(n21580), .A3(n21412), .ZN(n19995) );
  NOR2_X1 U30237 ( .A1(n21569), .A2(n20600), .ZN(n21402) );
  NOR2_X1 U30238 ( .A1(n21402), .A2(n19993), .ZN(n19994) );
  NOR2_X1 U30239 ( .A1(n24025), .A2(n354), .ZN(n20000) );
  OAI211_X1 U30240 ( .C1(n24041), .C2(n24034), .A(n7494), .B(n354), .ZN(n19998) );
  INV_X1 U30241 ( .A(n19998), .ZN(n19999) );
  NOR2_X1 U30243 ( .A1(n22101), .A2(n24034), .ZN(n23671) );
  INV_X1 U30244 ( .A(n23671), .ZN(n22577) );
  NAND2_X1 U30245 ( .A1(n22577), .A2(n23674), .ZN(n20002) );
  NOR2_X1 U30246 ( .A1(n24041), .A2(n24030), .ZN(n23667) );
  NAND2_X1 U30247 ( .A1(n20002), .A2(n22098), .ZN(n22574) );
  INV_X1 U30248 ( .A(n23666), .ZN(n22573) );
  OAI21_X1 U30249 ( .B1(n24025), .B2(n24030), .A(n22573), .ZN(n20003) );
  NAND2_X1 U30250 ( .A1(n20003), .A2(n22575), .ZN(n20004) );
  NAND2_X1 U30251 ( .A1(n22574), .A2(n20004), .ZN(n20007) );
  NOR2_X1 U30252 ( .A1(n24033), .A2(n354), .ZN(n22103) );
  OAI21_X1 U30253 ( .B1(n22103), .B2(n20005), .A(n22097), .ZN(n20006) );
  INV_X1 U30254 ( .A(n20012), .ZN(n20016) );
  MUX2_X1 U30256 ( .A(n20028), .B(n7920), .S(n20027), .Z(n20034) );
  INV_X1 U30257 ( .A(n20043), .ZN(n20031) );
  OAI211_X1 U30258 ( .C1(n20046), .C2(n20031), .A(n20030), .B(n7585), .ZN(
        n20033) );
  MUX2_X1 U30259 ( .A(n20034), .B(n20033), .S(n6515), .Z(n20051) );
  INV_X1 U30260 ( .A(n20035), .ZN(n20036) );
  NAND2_X1 U30261 ( .A1(n20036), .A2(n20044), .ZN(n20038) );
  AOI22_X1 U30262 ( .A1(n20039), .A2(n20038), .B1(n16820), .B2(n20037), .ZN(
        n20049) );
  NAND3_X1 U30263 ( .A1(n20041), .A2(n20040), .A3(n20042), .ZN(n20047) );
  NOR2_X1 U30264 ( .A1(n20049), .A2(n20048), .ZN(n20050) );
  NAND2_X1 U30265 ( .A1(n20052), .A2(n20082), .ZN(n20053) );
  NAND4_X1 U30266 ( .A1(n20055), .A2(n20071), .A3(n20054), .A4(n20053), .ZN(
        n20059) );
  NAND2_X1 U30267 ( .A1(n20057), .A2(n20056), .ZN(n20058) );
  OAI211_X1 U30268 ( .C1(n20073), .C2(n20060), .A(n20059), .B(n20058), .ZN(
        n20069) );
  AOI21_X1 U30269 ( .B1(n20063), .B2(n20062), .A(n20061), .ZN(n20066) );
  OAI21_X1 U30270 ( .B1(n20078), .B2(n20082), .A(n20071), .ZN(n20064) );
  AOI21_X1 U30271 ( .B1(n20066), .B2(n20065), .A(n20064), .ZN(n20068) );
  OAI22_X1 U30272 ( .A1(n20072), .A2(n20071), .B1(n20070), .B2(n20082), .ZN(
        n20077) );
  INV_X1 U30273 ( .A(n20073), .ZN(n20074) );
  AOI22_X1 U30274 ( .A1(n20077), .A2(n20076), .B1(n20075), .B2(n20074), .ZN(
        n20081) );
  NAND2_X1 U30275 ( .A1(n20079), .A2(n20078), .ZN(n20080) );
  NOR2_X1 U30276 ( .A1(n20084), .A2(n23414), .ZN(n24268) );
  OAI22_X1 U30277 ( .A1(n20089), .A2(n20088), .B1(n20087), .B2(n20086), .ZN(
        n20091) );
  NAND2_X1 U30278 ( .A1(n20093), .A2(n20092), .ZN(n20099) );
  OAI22_X1 U30279 ( .A1(n20096), .A2(n20095), .B1(n20094), .B2(n20104), .ZN(
        n20098) );
  MUX2_X1 U30280 ( .A(n20099), .B(n20098), .S(n20097), .Z(n20108) );
  NOR2_X1 U30281 ( .A1(n20101), .A2(n20100), .ZN(n20102) );
  OAI21_X1 U30282 ( .B1(n20103), .B2(n20102), .A(n16788), .ZN(n20107) );
  NAND2_X1 U30283 ( .A1(n20105), .A2(n20104), .ZN(n20106) );
  INV_X1 U30284 ( .A(n23411), .ZN(n23410) );
  NAND2_X1 U30285 ( .A1(n20111), .A2(n20110), .ZN(n20113) );
  INV_X1 U30287 ( .A(n20165), .ZN(n20129) );
  NAND2_X1 U30288 ( .A1(n20155), .A2(n20114), .ZN(n20115) );
  OAI21_X1 U30289 ( .B1(n20116), .B2(n20115), .A(n20158), .ZN(n20117) );
  NAND2_X1 U30290 ( .A1(n20117), .A2(n5058), .ZN(n20163) );
  OAI21_X1 U30291 ( .B1(n20119), .B2(n20118), .A(n20124), .ZN(n20121) );
  OAI211_X1 U30293 ( .C1(n20125), .C2(n20124), .A(n20123), .B(n20122), .ZN(
        n20126) );
  NAND3_X1 U30295 ( .A1(n20165), .A2(n20164), .A3(n20166), .ZN(n20128) );
  OAI21_X1 U30296 ( .B1(n20129), .B2(n20163), .A(n20128), .ZN(n20890) );
  OR2_X1 U30297 ( .A1(n20131), .A2(n20139), .ZN(n20154) );
  AOI22_X1 U30298 ( .A1(n20136), .A2(n20135), .B1(n20134), .B2(n52037), .ZN(
        n20153) );
  INV_X1 U30301 ( .A(n20139), .ZN(n20140) );
  INV_X1 U30303 ( .A(n20143), .ZN(n20150) );
  OAI211_X1 U30304 ( .C1(n20147), .C2(n51756), .A(n20145), .B(n20144), .ZN(
        n20149) );
  OAI21_X1 U30305 ( .B1(n20150), .B2(n20149), .A(n20148), .ZN(n20151) );
  OAI21_X1 U30306 ( .B1(n23417), .B2(n23408), .A(n23412), .ZN(n24267) );
  NOR2_X1 U30307 ( .A1(n24268), .A2(n24267), .ZN(n20173) );
  NAND2_X1 U30308 ( .A1(n20156), .A2(n20155), .ZN(n20159) );
  AOI21_X1 U30309 ( .B1(n20159), .B2(n20158), .A(n52176), .ZN(n20160) );
  NAND2_X1 U30310 ( .A1(n20162), .A2(n22037), .ZN(n20168) );
  NAND2_X1 U30311 ( .A1(n23414), .A2(n23411), .ZN(n22048) );
  INV_X1 U30312 ( .A(n20163), .ZN(n20167) );
  OAI211_X1 U30313 ( .C1(n20167), .C2(n20166), .A(n20165), .B(n20164), .ZN(
        n22036) );
  INV_X1 U30314 ( .A(n22036), .ZN(n22320) );
  NAND3_X1 U30315 ( .A1(n22048), .A2(n22320), .A3(n22037), .ZN(n20171) );
  OAI21_X1 U30316 ( .B1(n23423), .B2(n20168), .A(n20171), .ZN(n24272) );
  NAND3_X1 U30317 ( .A1(n23410), .A2(n22320), .A3(n2676), .ZN(n20169) );
  NOR2_X1 U30318 ( .A1(n23417), .A2(n20169), .ZN(n24266) );
  NAND3_X1 U30319 ( .A1(n23425), .A2(n22317), .A3(n23426), .ZN(n20170) );
  INV_X1 U30322 ( .A(n23417), .ZN(n20895) );
  NOR2_X1 U30323 ( .A1(n22034), .A2(n20895), .ZN(n20889) );
  AND2_X1 U30324 ( .A1(n23414), .A2(n23412), .ZN(n22314) );
  INV_X1 U30325 ( .A(n22314), .ZN(n22318) );
  NOR2_X1 U30326 ( .A1(n22318), .A2(n23408), .ZN(n23428) );
  AOI21_X1 U30327 ( .B1(n20889), .B2(n23407), .A(n23428), .ZN(n24271) );
  OAI211_X1 U30328 ( .C1(n20173), .C2(n24272), .A(n20172), .B(n24271), .ZN(
        n20174) );
  NAND2_X1 U30329 ( .A1(n20175), .A2(n21515), .ZN(n20182) );
  NAND2_X1 U30331 ( .A1(n51625), .A2(n21515), .ZN(n20181) );
  NAND3_X1 U30332 ( .A1(n20178), .A2(n21530), .A3(n20609), .ZN(n20180) );
  NAND3_X1 U30333 ( .A1(n20178), .A2(n20608), .A3(n20614), .ZN(n20179) );
  NAND3_X1 U30334 ( .A1(n20608), .A2(n20611), .A3(n51049), .ZN(n20183) );
  NAND2_X1 U30335 ( .A1(n21521), .A2(n51049), .ZN(n20186) );
  NAND2_X1 U30336 ( .A1(n20187), .A2(n20186), .ZN(n20191) );
  NAND3_X1 U30337 ( .A1(n20615), .A2(n20614), .A3(n20188), .ZN(n20189) );
  AOI21_X1 U30338 ( .B1(n21514), .B2(n20189), .A(n21513), .ZN(n20190) );
  MUX2_X1 U30339 ( .A(n20191), .B(n20190), .S(n20609), .Z(n20192) );
  NAND3_X1 U30340 ( .A1(n21548), .A2(n21533), .A3(n20197), .ZN(n20634) );
  AND2_X1 U30342 ( .A1(n20744), .A2(n20634), .ZN(n20206) );
  NAND2_X1 U30343 ( .A1(n20196), .A2(n21541), .ZN(n20205) );
  OAI211_X1 U30344 ( .C1(n21533), .C2(n51129), .A(n20742), .B(n21540), .ZN(
        n20200) );
  NAND4_X1 U30345 ( .A1(n20198), .A2(n20627), .A3(n21547), .A4(n20197), .ZN(
        n20199) );
  AND2_X1 U30346 ( .A1(n20200), .A2(n20199), .ZN(n20204) );
  XNOR2_X1 U30347 ( .A(n20641), .B(n20201), .ZN(n21542) );
  INV_X1 U30348 ( .A(n21542), .ZN(n20202) );
  NAND2_X1 U30349 ( .A1(n20202), .A2(n21548), .ZN(n20203) );
  OAI21_X1 U30350 ( .B1(n20212), .B2(n20211), .A(n20210), .ZN(n20213) );
  OAI21_X1 U30351 ( .B1(n51954), .B2(n20218), .A(n20217), .ZN(n20226) );
  AND2_X1 U30352 ( .A1(n20220), .A2(n51006), .ZN(n20223) );
  OAI22_X1 U30353 ( .A1(n51954), .A2(n20223), .B1(n20222), .B2(n20221), .ZN(
        n20225) );
  INV_X1 U30354 ( .A(n20668), .ZN(n20228) );
  NAND2_X1 U30355 ( .A1(n20228), .A2(n20681), .ZN(n20238) );
  OAI211_X1 U30356 ( .C1(n20678), .C2(n20681), .A(n20683), .B(n20232), .ZN(
        n20229) );
  AND2_X1 U30357 ( .A1(n20678), .A2(n20681), .ZN(n20235) );
  NAND2_X1 U30358 ( .A1(n20685), .A2(n1597), .ZN(n20234) );
  OAI211_X2 U30359 ( .C1(n20239), .C2(n20238), .A(n20237), .B(n20236), .ZN(
        n24247) );
  INV_X1 U30360 ( .A(n20875), .ZN(n21813) );
  AND2_X1 U30361 ( .A1(n24245), .A2(n24237), .ZN(n23456) );
  NAND2_X1 U30362 ( .A1(n21637), .A2(n21620), .ZN(n20243) );
  MUX2_X1 U30363 ( .A(n20243), .B(n20242), .S(n20241), .Z(n20265) );
  NAND3_X1 U30364 ( .A1(n21617), .A2(n20244), .A3(n21613), .ZN(n20245) );
  OAI211_X1 U30365 ( .C1(n20251), .C2(n20250), .A(n20249), .B(n20248), .ZN(
        n20252) );
  INV_X1 U30366 ( .A(n20252), .ZN(n20264) );
  NAND4_X1 U30367 ( .A1(n21614), .A2(n21617), .A3(n20698), .A4(n20256), .ZN(
        n20257) );
  OAI21_X1 U30368 ( .B1(n20258), .B2(n20698), .A(n20257), .ZN(n20261) );
  NOR2_X1 U30369 ( .A1(n20259), .A2(n21614), .ZN(n20260) );
  OAI211_X1 U30370 ( .C1(n20261), .C2(n20260), .A(n8367), .B(n21629), .ZN(
        n20262) );
  INV_X1 U30371 ( .A(n21653), .ZN(n20269) );
  AND2_X1 U30372 ( .A1(n52186), .A2(n20659), .ZN(n20274) );
  OAI211_X1 U30373 ( .C1(n20270), .C2(n20269), .A(n20268), .B(n20267), .ZN(
        n20271) );
  NAND2_X1 U30374 ( .A1(n20271), .A2(n20658), .ZN(n20280) );
  INV_X1 U30375 ( .A(n20272), .ZN(n20273) );
  OAI21_X1 U30376 ( .B1(n20273), .B2(n21664), .A(n21661), .ZN(n20279) );
  INV_X1 U30377 ( .A(n20274), .ZN(n20275) );
  NAND3_X1 U30378 ( .A1(n20277), .A2(n20276), .A3(n20275), .ZN(n20278) );
  AND2_X1 U30379 ( .A1(n23785), .A2(n21810), .ZN(n23455) );
  OAI21_X1 U30380 ( .B1(n23455), .B2(n23784), .A(n24250), .ZN(n20281) );
  NOR2_X1 U30381 ( .A1(n24237), .A2(n1497), .ZN(n20881) );
  INV_X1 U30382 ( .A(n20881), .ZN(n21819) );
  NAND2_X1 U30383 ( .A1(n24247), .A2(n21820), .ZN(n21818) );
  NOR3_X1 U30384 ( .A1(n21811), .A2(n21818), .A3(n21810), .ZN(n20283) );
  AND2_X1 U30385 ( .A1(n24250), .A2(n24247), .ZN(n23454) );
  NAND2_X1 U30386 ( .A1(n21811), .A2(n24245), .ZN(n20872) );
  INV_X1 U30389 ( .A(n21818), .ZN(n20285) );
  AOI21_X1 U30390 ( .B1(n20289), .B2(n320), .A(n22823), .ZN(n20292) );
  NAND2_X1 U30392 ( .A1(n22490), .A2(n22830), .ZN(n20290) );
  NOR2_X1 U30393 ( .A1(n22503), .A2(n20290), .ZN(n20291) );
  INV_X1 U30394 ( .A(n21070), .ZN(n22502) );
  OAI22_X1 U30395 ( .A1(n20292), .A2(n20291), .B1(n22502), .B2(n320), .ZN(
        n20303) );
  INV_X1 U30396 ( .A(n20293), .ZN(n20295) );
  NOR2_X1 U30397 ( .A1(n22830), .A2(n22491), .ZN(n20296) );
  NAND2_X1 U30398 ( .A1(n20296), .A2(n22832), .ZN(n21071) );
  NAND3_X1 U30399 ( .A1(n22832), .A2(n22491), .A3(n22509), .ZN(n22820) );
  NAND2_X1 U30400 ( .A1(n21071), .A2(n22820), .ZN(n20294) );
  OAI21_X1 U30402 ( .B1(n22492), .B2(n22491), .A(n22509), .ZN(n22828) );
  INV_X1 U30403 ( .A(n22828), .ZN(n22225) );
  NOR2_X1 U30404 ( .A1(n22826), .A2(n22491), .ZN(n22824) );
  OAI21_X1 U30405 ( .B1(n22503), .B2(n20297), .A(n22496), .ZN(n22229) );
  OAI21_X1 U30406 ( .B1(n22225), .B2(n22824), .A(n22229), .ZN(n20301) );
  NOR2_X1 U30407 ( .A1(n22822), .A2(n20298), .ZN(n20299) );
  OAI21_X1 U30408 ( .B1(n20299), .B2(n21068), .A(n21073), .ZN(n20300) );
  XNOR2_X1 U30410 ( .A(n22695), .B(n25915), .ZN(n25333) );
  OAI21_X1 U30411 ( .B1(n23225), .B2(n51355), .A(n20304), .ZN(n20308) );
  NOR2_X1 U30412 ( .A1(n22121), .A2(n23229), .ZN(n23223) );
  INV_X1 U30414 ( .A(n20306), .ZN(n20307) );
  INV_X1 U30415 ( .A(n23225), .ZN(n21722) );
  AOI22_X1 U30416 ( .A1(n21722), .A2(n2102), .B1(n23223), .B2(n23207), .ZN(
        n20313) );
  NAND2_X1 U30417 ( .A1(n51355), .A2(n2102), .ZN(n21723) );
  AOI21_X1 U30418 ( .B1(n413), .B2(n23230), .A(n23207), .ZN(n20310) );
  NAND2_X1 U30419 ( .A1(n20311), .A2(n20310), .ZN(n20312) );
  OAI211_X1 U30420 ( .C1(n21462), .C2(n20493), .A(n21460), .B(n21451), .ZN(
        n20315) );
  MUX2_X1 U30421 ( .A(n20315), .B(n20314), .S(n21468), .Z(n20319) );
  NAND3_X1 U30422 ( .A1(n20316), .A2(n21465), .A3(n21474), .ZN(n20318) );
  NOR2_X1 U30423 ( .A1(n20327), .A2(n52139), .ZN(n20843) );
  NAND2_X1 U30424 ( .A1(n20843), .A2(n21427), .ZN(n21444) );
  OAI21_X1 U30425 ( .B1(n20327), .B2(n21424), .A(n20838), .ZN(n20320) );
  NAND2_X1 U30427 ( .A1(n21439), .A2(n21443), .ZN(n20323) );
  OAI22_X1 U30428 ( .A1(n20327), .A2(n20326), .B1(n20325), .B2(n21425), .ZN(
        n20328) );
  OAI22_X1 U30429 ( .A1(n20826), .A2(n20812), .B1(n21485), .B2(n20448), .ZN(
        n20333) );
  NAND2_X1 U30430 ( .A1(n20333), .A2(n20813), .ZN(n20342) );
  NAND3_X1 U30431 ( .A1(n20334), .A2(n21495), .A3(n20825), .ZN(n20335) );
  NAND2_X1 U30432 ( .A1(n20336), .A2(n20335), .ZN(n20337) );
  NAND2_X1 U30433 ( .A1(n20815), .A2(n763), .ZN(n20340) );
  NAND2_X1 U30434 ( .A1(n2220), .A2(n21486), .ZN(n20338) );
  OAI211_X1 U30435 ( .C1(n763), .C2(n21483), .A(n20826), .B(n20338), .ZN(
        n20339) );
  NAND2_X1 U30436 ( .A1(n23045), .A2(n22748), .ZN(n22080) );
  AND2_X1 U30437 ( .A1(n20434), .A2(n20432), .ZN(n20344) );
  OAI22_X1 U30438 ( .A1(n20345), .A2(n20344), .B1(n6452), .B2(n20343), .ZN(
        n20346) );
  NAND3_X1 U30439 ( .A1(n20346), .A2(n20426), .A3(n20435), .ZN(n20370) );
  INV_X1 U30440 ( .A(n20347), .ZN(n20352) );
  OAI21_X1 U30441 ( .B1(n20354), .B2(n20435), .A(n20426), .ZN(n20350) );
  AOI22_X1 U30442 ( .A1(n20352), .A2(n20351), .B1(n20350), .B2(n20349), .ZN(
        n20369) );
  NAND2_X1 U30443 ( .A1(n20428), .A2(n20426), .ZN(n20353) );
  NAND4_X1 U30444 ( .A1(n20357), .A2(n20359), .A3(n20354), .A4(n20353), .ZN(
        n20355) );
  AND2_X1 U30445 ( .A1(n20356), .A2(n20355), .ZN(n20368) );
  AOI21_X1 U30446 ( .B1(n20358), .B2(n20359), .A(n20357), .ZN(n20366) );
  NAND2_X1 U30447 ( .A1(n20430), .A2(n20426), .ZN(n20431) );
  OAI21_X1 U30448 ( .B1(n20360), .B2(n20359), .A(n20427), .ZN(n20361) );
  NAND2_X1 U30449 ( .A1(n20431), .A2(n20361), .ZN(n20365) );
  INV_X1 U30450 ( .A(n20362), .ZN(n20364) );
  AOI22_X1 U30451 ( .A1(n20366), .A2(n20365), .B1(n20364), .B2(n20363), .ZN(
        n20367) );
  NAND4_X2 U30452 ( .A1(n20367), .A2(n20369), .A3(n20370), .A4(n20368), .ZN(
        n23052) );
  AND2_X1 U30453 ( .A1(n20371), .A2(n20791), .ZN(n20411) );
  OAI21_X1 U30454 ( .B1(n20408), .B2(n20375), .A(n581), .ZN(n20372) );
  NAND2_X1 U30455 ( .A1(n20411), .A2(n20372), .ZN(n20374) );
  INV_X1 U30456 ( .A(n20377), .ZN(n20379) );
  INV_X1 U30457 ( .A(n21369), .ZN(n21386) );
  NAND2_X1 U30458 ( .A1(n21386), .A2(n21388), .ZN(n20378) );
  NAND3_X1 U30459 ( .A1(n20380), .A2(n1860), .A3(n358), .ZN(n20413) );
  OAI21_X1 U30460 ( .B1(n581), .B2(n20413), .A(n21373), .ZN(n20381) );
  NAND2_X1 U30461 ( .A1(n20385), .A2(n20476), .ZN(n20403) );
  NOR2_X1 U30462 ( .A1(n20394), .A2(n20466), .ZN(n20386) );
  NAND4_X1 U30466 ( .A1(n17639), .A2(n3745), .A3(n20394), .A4(n20393), .ZN(
        n20395) );
  OAI21_X1 U30467 ( .B1(n20397), .B2(n20396), .A(n20395), .ZN(n20398) );
  AOI21_X1 U30468 ( .B1(n4098), .B2(n20399), .A(n20398), .ZN(n20401) );
  NAND2_X1 U30469 ( .A1(n424), .A2(n23054), .ZN(n22090) );
  INV_X1 U30470 ( .A(n23052), .ZN(n22201) );
  NOR2_X1 U30471 ( .A1(n23054), .A2(n23044), .ZN(n22072) );
  OAI211_X1 U30472 ( .C1(n23052), .C2(n23054), .A(n23049), .B(n23044), .ZN(
        n20404) );
  AND2_X1 U30473 ( .A1(n20404), .A2(n22753), .ZN(n20406) );
  NOR2_X1 U30474 ( .A1(n23052), .A2(n23044), .ZN(n22197) );
  OAI21_X1 U30475 ( .B1(n424), .B2(n22748), .A(n22197), .ZN(n22199) );
  NOR2_X1 U30476 ( .A1(n22201), .A2(n22087), .ZN(n22947) );
  AOI22_X1 U30477 ( .A1(n20406), .A2(n22199), .B1(n22947), .B2(n23048), .ZN(
        n20407) );
  XNOR2_X1 U30478 ( .A(n26100), .B(n26395), .ZN(n20538) );
  INV_X1 U30479 ( .A(n20408), .ZN(n20788) );
  OAI21_X1 U30480 ( .B1(n21397), .B2(n20412), .A(n20411), .ZN(n20419) );
  INV_X1 U30481 ( .A(n20413), .ZN(n20414) );
  AND2_X1 U30482 ( .A1(n21388), .A2(n21389), .ZN(n20797) );
  NAND2_X1 U30483 ( .A1(n20414), .A2(n20797), .ZN(n20418) );
  NAND2_X1 U30484 ( .A1(n20416), .A2(n20415), .ZN(n20417) );
  OAI21_X1 U30485 ( .B1(n20422), .B2(n20421), .A(n20420), .ZN(n20424) );
  AOI22_X1 U30486 ( .A1(n20430), .A2(n20429), .B1(n20428), .B2(n20427), .ZN(
        n20439) );
  INV_X1 U30487 ( .A(n20431), .ZN(n20433) );
  NAND2_X1 U30488 ( .A1(n20433), .A2(n20432), .ZN(n20438) );
  NAND3_X1 U30489 ( .A1(n20436), .A2(n20435), .A3(n20434), .ZN(n20437) );
  NAND4_X2 U30490 ( .A1(n20440), .A2(n20439), .A3(n20438), .A4(n20437), .ZN(
        n22306) );
  NAND2_X1 U30491 ( .A1(n22714), .A2(n22306), .ZN(n20542) );
  OAI21_X1 U30492 ( .B1(n20811), .B2(n20826), .A(n20447), .ZN(n20445) );
  NAND2_X1 U30493 ( .A1(n21491), .A2(n20812), .ZN(n20444) );
  NAND2_X1 U30494 ( .A1(n21486), .A2(n20441), .ZN(n20442) );
  OAI22_X1 U30495 ( .A1(n21482), .A2(n20824), .B1(n20811), .B2(n20442), .ZN(
        n20443) );
  AOI21_X1 U30496 ( .B1(n20445), .B2(n20444), .A(n20443), .ZN(n20457) );
  INV_X1 U30497 ( .A(n21480), .ZN(n20446) );
  NAND2_X1 U30498 ( .A1(n20810), .A2(n20813), .ZN(n20456) );
  INV_X1 U30499 ( .A(n20448), .ZN(n20452) );
  NOR2_X1 U30500 ( .A1(n20449), .A2(n20825), .ZN(n20450) );
  AOI22_X1 U30501 ( .A1(n20453), .A2(n20452), .B1(n20451), .B2(n20450), .ZN(
        n20455) );
  NAND4_X2 U30502 ( .A1(n20457), .A2(n20455), .A3(n20456), .A4(n20454), .ZN(
        n22464) );
  AOI22_X1 U30503 ( .A1(n20460), .A2(n20459), .B1(n20480), .B2(n20458), .ZN(
        n20464) );
  NAND3_X1 U30504 ( .A1(n20462), .A2(n20461), .A3(n17639), .ZN(n20463) );
  INV_X1 U30505 ( .A(n20467), .ZN(n20470) );
  NOR2_X1 U30506 ( .A1(n20468), .A2(n20473), .ZN(n20469) );
  OAI21_X1 U30507 ( .B1(n20470), .B2(n20469), .A(n20477), .ZN(n20486) );
  NAND2_X1 U30508 ( .A1(n20480), .A2(n20477), .ZN(n20482) );
  NAND2_X1 U30509 ( .A1(n20484), .A2(n20483), .ZN(n20485) );
  OAI21_X1 U30510 ( .B1(n20542), .B2(n22464), .A(n22709), .ZN(n20522) );
  NAND2_X1 U30511 ( .A1(n20489), .A2(n20488), .ZN(n20491) );
  NAND4_X1 U30512 ( .A1(n21451), .A2(n21449), .A3(n20493), .A4(n21450), .ZN(
        n20494) );
  AND2_X2 U30514 ( .A1(n20500), .A2(n20499), .ZN(n22488) );
  NAND2_X1 U30515 ( .A1(n632), .A2(n20501), .ZN(n20502) );
  NAND4_X1 U30516 ( .A1(n17619), .A2(n20504), .A3(n20503), .A4(n20502), .ZN(
        n20510) );
  AOI21_X1 U30517 ( .B1(n20513), .B2(n20507), .A(n20506), .ZN(n20509) );
  MUX2_X1 U30518 ( .A(n20510), .B(n20509), .S(n20508), .Z(n20521) );
  OAI21_X1 U30519 ( .B1(n20513), .B2(n20512), .A(n20511), .ZN(n20520) );
  AOI21_X1 U30520 ( .B1(n20515), .B2(n51705), .A(n20514), .ZN(n20516) );
  NAND2_X1 U30521 ( .A1(n20517), .A2(n20516), .ZN(n20518) );
  NAND2_X1 U30522 ( .A1(n22488), .A2(n22470), .ZN(n22711) );
  INV_X1 U30523 ( .A(n22711), .ZN(n22717) );
  INV_X1 U30524 ( .A(n22306), .ZN(n22471) );
  OAI211_X1 U30525 ( .C1(n22476), .C2(n22470), .A(n22462), .B(n22479), .ZN(
        n20526) );
  INV_X1 U30526 ( .A(n21130), .ZN(n22715) );
  OAI21_X1 U30527 ( .B1(n22715), .B2(n20523), .A(n22308), .ZN(n20525) );
  NAND2_X1 U30529 ( .A1(n20548), .A2(n51124), .ZN(n20524) );
  NAND2_X1 U30530 ( .A1(n22306), .A2(n22464), .ZN(n22461) );
  NOR2_X1 U30531 ( .A1(n22481), .A2(n22470), .ZN(n22720) );
  OAI211_X1 U30532 ( .C1(n22720), .C2(n22464), .A(n22711), .B(n21130), .ZN(
        n20527) );
  OAI211_X1 U30533 ( .C1(n22481), .C2(n22479), .A(n51124), .B(n22306), .ZN(
        n20528) );
  NAND2_X1 U30534 ( .A1(n20531), .A2(n21780), .ZN(n20537) );
  NAND2_X1 U30535 ( .A1(n21117), .A2(n21767), .ZN(n20532) );
  AND2_X1 U30536 ( .A1(n22701), .A2(n21767), .ZN(n21125) );
  NAND2_X1 U30537 ( .A1(n20948), .A2(n21125), .ZN(n20533) );
  NAND3_X1 U30538 ( .A1(n20534), .A2(n51081), .A3(n22703), .ZN(n20536) );
  INV_X1 U30539 ( .A(n21782), .ZN(n20943) );
  NOR2_X1 U30540 ( .A1(n21767), .A2(n24452), .ZN(n20939) );
  AOI21_X1 U30541 ( .B1(n20943), .B2(n20942), .A(n20939), .ZN(n20535) );
  NOR2_X1 U30542 ( .A1(n21780), .A2(n22701), .ZN(n22699) );
  XNOR2_X2 U30543 ( .A(n28104), .B(n26390), .ZN(n27452) );
  XNOR2_X1 U30544 ( .A(n20538), .B(n27452), .ZN(n20539) );
  XNOR2_X1 U30545 ( .A(n25333), .B(n20539), .ZN(n20540) );
  OR2_X1 U30546 ( .A1(n27618), .A2(n27729), .ZN(n22341) );
  INV_X1 U30547 ( .A(n20542), .ZN(n20543) );
  NAND3_X1 U30548 ( .A1(n20543), .A2(n22721), .A3(n2083), .ZN(n20545) );
  AND2_X1 U30549 ( .A1(n22714), .A2(n22479), .ZN(n20547) );
  NAND2_X1 U30550 ( .A1(n51124), .A2(n22462), .ZN(n22713) );
  NAND3_X1 U30551 ( .A1(n20547), .A2(n22711), .A3(n22713), .ZN(n20544) );
  AND2_X1 U30552 ( .A1(n20545), .A2(n20544), .ZN(n20554) );
  NAND2_X1 U30553 ( .A1(n22464), .A2(n51124), .ZN(n22482) );
  NOR2_X1 U30554 ( .A1(n22482), .A2(n22714), .ZN(n20546) );
  AND2_X1 U30555 ( .A1(n22306), .A2(n22479), .ZN(n22722) );
  OAI21_X1 U30556 ( .B1(n21130), .B2(n22464), .A(n22716), .ZN(n20551) );
  NAND2_X1 U30557 ( .A1(n22306), .A2(n22488), .ZN(n20549) );
  OAI211_X1 U30558 ( .C1(n22462), .C2(n22479), .A(n22711), .B(n20549), .ZN(
        n20550) );
  NOR2_X1 U30559 ( .A1(n24207), .A2(n23613), .ZN(n24205) );
  NAND2_X1 U30560 ( .A1(n24206), .A2(n24205), .ZN(n23601) );
  NAND2_X1 U30561 ( .A1(n24208), .A2(n52155), .ZN(n20556) );
  NAND3_X1 U30562 ( .A1(n23601), .A2(n24211), .A3(n20556), .ZN(n20560) );
  NOR2_X1 U30563 ( .A1(n24207), .A2(n22639), .ZN(n23081) );
  INV_X1 U30564 ( .A(n23081), .ZN(n23077) );
  NAND2_X1 U30565 ( .A1(n24211), .A2(n23068), .ZN(n23078) );
  OAI21_X1 U30566 ( .B1(n23077), .B2(n23080), .A(n23078), .ZN(n20557) );
  NAND3_X1 U30567 ( .A1(n23604), .A2(n23068), .A3(n22639), .ZN(n20559) );
  NAND2_X1 U30568 ( .A1(n17418), .A2(n52155), .ZN(n23072) );
  INV_X1 U30569 ( .A(n23591), .ZN(n23597) );
  OR2_X1 U30570 ( .A1(n23072), .A2(n23597), .ZN(n20558) );
  NAND2_X1 U30571 ( .A1(n20561), .A2(n22184), .ZN(n20562) );
  MUX2_X1 U30572 ( .A(n20563), .B(n20562), .S(n52048), .Z(n20565) );
  NAND3_X1 U30573 ( .A1(n22178), .A2(n21712), .A3(n52048), .ZN(n20566) );
  NAND2_X1 U30574 ( .A1(n21105), .A2(n21714), .ZN(n21702) );
  NOR2_X1 U30575 ( .A1(n21702), .A2(n22186), .ZN(n20567) );
  XNOR2_X1 U30576 ( .A(n35107), .B(n4423), .ZN(n43537) );
  XNOR2_X1 U30577 ( .A(n43537), .B(n4666), .ZN(n20571) );
  XNOR2_X1 U30578 ( .A(n51666), .B(n20571), .ZN(n20572) );
  INV_X1 U30579 ( .A(n22377), .ZN(n20573) );
  NAND3_X1 U30580 ( .A1(n20574), .A2(n20573), .A3(n21062), .ZN(n20578) );
  NAND2_X1 U30581 ( .A1(n22377), .A2(n22390), .ZN(n20575) );
  AOI21_X1 U30583 ( .B1(n23811), .B2(n753), .A(n22741), .ZN(n20576) );
  NAND3_X1 U30584 ( .A1(n20576), .A2(n22386), .A3(n8310), .ZN(n20577) );
  XNOR2_X1 U30585 ( .A(n22375), .B(n753), .ZN(n20579) );
  AOI21_X1 U30586 ( .B1(n20581), .B2(n20580), .A(n50976), .ZN(n20582) );
  AND2_X1 U30587 ( .A1(n23827), .A2(n23825), .ZN(n23822) );
  INV_X1 U30588 ( .A(n23822), .ZN(n20584) );
  AOI22_X1 U30589 ( .A1(n24158), .A2(n24157), .B1(n20584), .B2(n23826), .ZN(
        n20586) );
  OR2_X1 U30590 ( .A1(n23827), .A2(n23825), .ZN(n20592) );
  OAI211_X1 U30591 ( .C1(n20587), .C2(n24157), .A(n20586), .B(n20585), .ZN(
        n20599) );
  AND2_X1 U30593 ( .A1(n23827), .A2(n24158), .ZN(n23267) );
  NAND3_X1 U30594 ( .A1(n23267), .A2(n23828), .A3(n23821), .ZN(n20589) );
  NAND2_X1 U30595 ( .A1(n20590), .A2(n20589), .ZN(n20591) );
  NAND2_X1 U30596 ( .A1(n20591), .A2(n23833), .ZN(n20598) );
  NAND2_X1 U30597 ( .A1(n23824), .A2(n1941), .ZN(n20595) );
  NAND2_X1 U30598 ( .A1(n23822), .A2(n23821), .ZN(n20594) );
  NAND2_X1 U30599 ( .A1(n20592), .A2(n23832), .ZN(n20593) );
  NAND3_X1 U30600 ( .A1(n20595), .A2(n20594), .A3(n20593), .ZN(n20596) );
  NAND2_X1 U30601 ( .A1(n20596), .A2(n24150), .ZN(n20597) );
  INV_X1 U30602 ( .A(n21569), .ZN(n21565) );
  NAND3_X1 U30603 ( .A1(n21565), .A2(n21407), .A3(n21556), .ZN(n21574) );
  NAND2_X1 U30604 ( .A1(n21403), .A2(n20601), .ZN(n20602) );
  OAI211_X1 U30605 ( .C1(n21413), .C2(n21569), .A(n20603), .B(n20602), .ZN(
        n20604) );
  NAND4_X1 U30606 ( .A1(n20605), .A2(n51711), .A3(n21569), .A4(n21583), .ZN(
        n20606) );
  OAI22_X1 U30607 ( .A1(n21521), .A2(n20609), .B1(n20608), .B2(n20607), .ZN(
        n20610) );
  NAND2_X1 U30608 ( .A1(n20610), .A2(n21515), .ZN(n20622) );
  AOI22_X1 U30609 ( .A1(n21513), .A2(n21528), .B1(n20611), .B2(n20615), .ZN(
        n20621) );
  NAND2_X1 U30610 ( .A1(n21531), .A2(n20612), .ZN(n20620) );
  AOI21_X1 U30611 ( .B1(n7431), .B2(n16125), .A(n52213), .ZN(n20617) );
  OAI211_X1 U30613 ( .C1(n20617), .C2(n21520), .A(n21514), .B(n20616), .ZN(
        n20618) );
  NAND2_X1 U30614 ( .A1(n20618), .A2(n21521), .ZN(n20619) );
  NAND2_X1 U30615 ( .A1(n23706), .A2(n23535), .ZN(n20711) );
  OAI22_X1 U30616 ( .A1(n20736), .A2(n20624), .B1(n20746), .B2(n20623), .ZN(
        n20626) );
  OAI21_X1 U30617 ( .B1(n20626), .B2(n20625), .A(n21541), .ZN(n20637) );
  OAI21_X1 U30618 ( .B1(n20629), .B2(n18495), .A(n20752), .ZN(n20636) );
  NAND2_X1 U30621 ( .A1(n21542), .A2(n20638), .ZN(n20640) );
  NAND2_X1 U30622 ( .A1(n21548), .A2(n20736), .ZN(n20639) );
  AOI21_X1 U30623 ( .B1(n20640), .B2(n20639), .A(n20738), .ZN(n20645) );
  NAND3_X1 U30624 ( .A1(n20742), .A2(n20641), .A3(n21547), .ZN(n20643) );
  NAND2_X1 U30625 ( .A1(n21663), .A2(n21661), .ZN(n20651) );
  NAND2_X1 U30626 ( .A1(n21647), .A2(n20651), .ZN(n20654) );
  NAND2_X1 U30627 ( .A1(n20651), .A2(n20658), .ZN(n20653) );
  NAND3_X1 U30628 ( .A1(n20654), .A2(n20653), .A3(n20652), .ZN(n20666) );
  NAND2_X1 U30629 ( .A1(n20655), .A2(n21649), .ZN(n20665) );
  NOR2_X1 U30630 ( .A1(n20657), .A2(n20656), .ZN(n20663) );
  XNOR2_X1 U30631 ( .A(n20658), .B(n21661), .ZN(n20662) );
  OAI21_X1 U30632 ( .B1(n20660), .B2(n21661), .A(n20659), .ZN(n20661) );
  OAI211_X1 U30633 ( .C1(n20663), .C2(n21646), .A(n20662), .B(n20661), .ZN(
        n20664) );
  NAND3_X1 U30634 ( .A1(n20672), .A2(n20671), .A3(n20670), .ZN(n20673) );
  OAI211_X1 U30635 ( .C1(n20675), .C2(n18101), .A(n20674), .B(n20673), .ZN(
        n20676) );
  INV_X1 U30636 ( .A(n20676), .ZN(n20691) );
  OAI211_X1 U30637 ( .C1(n20688), .C2(n20681), .A(n1597), .B(n20680), .ZN(
        n20690) );
  OAI22_X1 U30638 ( .A1(n20685), .A2(n20684), .B1(n20683), .B2(n20682), .ZN(
        n20687) );
  OAI21_X1 U30639 ( .B1(n20688), .B2(n20687), .A(n20686), .ZN(n20689) );
  NAND3_X1 U30640 ( .A1(n20697), .A2(n8367), .A3(n21619), .ZN(n20703) );
  NAND3_X1 U30641 ( .A1(n20700), .A2(n20698), .A3(n21629), .ZN(n20702) );
  OAI21_X1 U30642 ( .B1(n20698), .B2(n21629), .A(n21630), .ZN(n20699) );
  AOI22_X1 U30643 ( .A1(n20700), .A2(n20699), .B1(n21620), .B2(n21614), .ZN(
        n20701) );
  NOR2_X1 U30644 ( .A1(n24332), .A2(n457), .ZN(n23708) );
  INV_X1 U30645 ( .A(n23708), .ZN(n20706) );
  OAI211_X1 U30646 ( .C1(n23703), .C2(n23694), .A(n20707), .B(n20706), .ZN(
        n20710) );
  NAND2_X1 U30647 ( .A1(n24332), .A2(n5415), .ZN(n22236) );
  INV_X1 U30648 ( .A(n22236), .ZN(n24331) );
  INV_X1 U30649 ( .A(n23694), .ZN(n20708) );
  NAND3_X1 U30650 ( .A1(n24331), .A2(n23702), .A3(n20708), .ZN(n20709) );
  NOR2_X1 U30651 ( .A1(n24332), .A2(n23531), .ZN(n24326) );
  INV_X1 U30652 ( .A(n24326), .ZN(n23540) );
  INV_X1 U30653 ( .A(n23693), .ZN(n24329) );
  NAND2_X1 U30654 ( .A1(n23531), .A2(n23535), .ZN(n23704) );
  NAND3_X1 U30655 ( .A1(n23540), .A2(n24329), .A3(n23704), .ZN(n20717) );
  NOR2_X1 U30656 ( .A1(n20711), .A2(n457), .ZN(n24338) );
  INV_X1 U30657 ( .A(n24338), .ZN(n20716) );
  OAI21_X1 U30658 ( .B1(n50990), .B2(n5415), .A(n3822), .ZN(n20712) );
  AOI21_X1 U30659 ( .B1(n20712), .B2(n24332), .A(n23531), .ZN(n20713) );
  OAI21_X1 U30660 ( .B1(n23538), .B2(n24332), .A(n20713), .ZN(n20715) );
  NOR2_X1 U30661 ( .A1(n23374), .A2(n457), .ZN(n23375) );
  NAND2_X1 U30662 ( .A1(n23375), .A2(n50990), .ZN(n20714) );
  NAND4_X1 U30663 ( .A1(n20717), .A2(n20716), .A3(n20715), .A4(n20714), .ZN(
        n20718) );
  AND2_X1 U30664 ( .A1(n23547), .A2(n21155), .ZN(n23362) );
  OAI21_X1 U30665 ( .B1(n23362), .B2(n20720), .A(n23364), .ZN(n20725) );
  AND2_X1 U30666 ( .A1(n20721), .A2(n23547), .ZN(n21157) );
  INV_X1 U30667 ( .A(n23350), .ZN(n23553) );
  NAND2_X1 U30668 ( .A1(n21157), .A2(n23553), .ZN(n20724) );
  NOR2_X1 U30669 ( .A1(n23562), .A2(n51676), .ZN(n23361) );
  NAND2_X1 U30670 ( .A1(n23361), .A2(n23360), .ZN(n20722) );
  NOR2_X1 U30671 ( .A1(n8205), .A2(n21155), .ZN(n20729) );
  INV_X1 U30672 ( .A(n20727), .ZN(n20728) );
  OAI21_X1 U30673 ( .B1(n23549), .B2(n20729), .A(n20728), .ZN(n20734) );
  NOR2_X1 U30674 ( .A1(n23547), .A2(n23563), .ZN(n23356) );
  INV_X1 U30675 ( .A(n23356), .ZN(n20731) );
  NOR2_X1 U30676 ( .A1(n23360), .A2(n23546), .ZN(n21156) );
  AND2_X1 U30677 ( .A1(n21156), .A2(n23547), .ZN(n23357) );
  INV_X1 U30678 ( .A(n23357), .ZN(n20730) );
  OAI21_X1 U30679 ( .B1(n20731), .B2(n23570), .A(n20730), .ZN(n20732) );
  NAND2_X1 U30680 ( .A1(n51677), .A2(n23568), .ZN(n23554) );
  NAND2_X1 U30681 ( .A1(n20732), .A2(n752), .ZN(n20733) );
  NOR2_X1 U30682 ( .A1(n20737), .A2(n20736), .ZN(n20748) );
  NOR2_X1 U30684 ( .A1(n20739), .A2(n20738), .ZN(n20740) );
  NAND2_X1 U30685 ( .A1(n20742), .A2(n20745), .ZN(n20743) );
  AND2_X1 U30686 ( .A1(n20744), .A2(n20743), .ZN(n20755) );
  NOR2_X1 U30687 ( .A1(n20746), .A2(n20745), .ZN(n20747) );
  OAI21_X1 U30688 ( .B1(n20748), .B2(n20747), .A(n21541), .ZN(n20754) );
  OAI21_X1 U30689 ( .B1(n20752), .B2(n20751), .A(n20750), .ZN(n20753) );
  NAND2_X1 U30690 ( .A1(n21599), .A2(n52208), .ZN(n20757) );
  OAI21_X1 U30691 ( .B1(n21360), .B2(n20757), .A(n21601), .ZN(n20764) );
  OAI21_X1 U30692 ( .B1(n21599), .B2(n21364), .A(n21362), .ZN(n20763) );
  INV_X1 U30693 ( .A(n20758), .ZN(n21607) );
  NAND2_X1 U30694 ( .A1(n21604), .A2(n21351), .ZN(n20759) );
  AOI22_X1 U30695 ( .A1(n20764), .A2(n20763), .B1(n20762), .B2(n20761), .ZN(
        n20774) );
  INV_X1 U30696 ( .A(n20765), .ZN(n20766) );
  OAI211_X1 U30697 ( .C1(n20766), .C2(n21358), .A(n21362), .B(n20768), .ZN(
        n20773) );
  INV_X1 U30698 ( .A(n20767), .ZN(n20770) );
  NOR2_X1 U30699 ( .A1(n20768), .A2(n21362), .ZN(n20769) );
  AOI22_X1 U30700 ( .A1(n20770), .A2(n21350), .B1(n20769), .B2(n21592), .ZN(
        n20772) );
  NAND2_X1 U30701 ( .A1(n23641), .A2(n23637), .ZN(n22625) );
  INV_X1 U30702 ( .A(n21566), .ZN(n20775) );
  NOR3_X1 U30703 ( .A1(n20775), .A2(n21555), .A3(n51755), .ZN(n20776) );
  NAND2_X1 U30704 ( .A1(n20777), .A2(n20776), .ZN(n20786) );
  AOI22_X1 U30705 ( .A1(n951), .A2(n21565), .B1(n21407), .B2(n21584), .ZN(
        n20785) );
  AND2_X1 U30706 ( .A1(n21559), .A2(n20778), .ZN(n20780) );
  NAND2_X1 U30707 ( .A1(n20788), .A2(n581), .ZN(n20790) );
  NOR2_X1 U30708 ( .A1(n1860), .A2(n5923), .ZN(n20789) );
  OAI22_X1 U30709 ( .A1(n21369), .A2(n21396), .B1(n20792), .B2(n20791), .ZN(
        n20793) );
  OAI21_X1 U30710 ( .B1(n20798), .B2(n20797), .A(n20796), .ZN(n20799) );
  NAND2_X1 U30711 ( .A1(n20799), .A2(n769), .ZN(n20803) );
  NAND2_X1 U30712 ( .A1(n358), .A2(n21389), .ZN(n20800) );
  NOR2_X1 U30713 ( .A1(n21396), .A2(n20800), .ZN(n20801) );
  NAND2_X1 U30714 ( .A1(n20805), .A2(n1860), .ZN(n20806) );
  NOR2_X1 U30715 ( .A1(n21382), .A2(n20806), .ZN(n20807) );
  OR2_X2 U30716 ( .A1(n20808), .A2(n20807), .ZN(n23961) );
  AOI21_X1 U30717 ( .B1(n23950), .B2(n23090), .A(n23961), .ZN(n20809) );
  OAI21_X1 U30718 ( .B1(n22625), .B2(n23950), .A(n20809), .ZN(n20851) );
  INV_X1 U30719 ( .A(n20827), .ZN(n20814) );
  OAI211_X1 U30720 ( .C1(n20815), .C2(n20814), .A(n20828), .B(n20813), .ZN(
        n20816) );
  INV_X1 U30721 ( .A(n20817), .ZN(n20819) );
  INV_X1 U30722 ( .A(n20820), .ZN(n20823) );
  NAND2_X1 U30723 ( .A1(n20821), .A2(n21495), .ZN(n20822) );
  NAND2_X1 U30724 ( .A1(n20830), .A2(n20829), .ZN(n20831) );
  NAND3_X1 U30725 ( .A1(n20839), .A2(n20838), .A3(n20837), .ZN(n20845) );
  NOR2_X1 U30726 ( .A1(n21425), .A2(n5500), .ZN(n20842) );
  AOI21_X1 U30727 ( .B1(n20843), .B2(n21420), .A(n20842), .ZN(n20844) );
  AND2_X1 U30728 ( .A1(n23955), .A2(n559), .ZN(n23965) );
  INV_X1 U30729 ( .A(n23965), .ZN(n20850) );
  AND2_X1 U30730 ( .A1(n23090), .A2(n559), .ZN(n20849) );
  INV_X1 U30731 ( .A(n23950), .ZN(n23958) );
  AND2_X1 U30732 ( .A1(n23958), .A2(n23955), .ZN(n20853) );
  AND2_X1 U30733 ( .A1(n22623), .A2(n23961), .ZN(n23959) );
  AOI22_X1 U30734 ( .A1(n20853), .A2(n23959), .B1(n20852), .B2(n23950), .ZN(
        n20855) );
  AND2_X1 U30735 ( .A1(n23961), .A2(n559), .ZN(n23635) );
  AOI22_X1 U30736 ( .A1(n23953), .A2(n23622), .B1(n23635), .B2(n23956), .ZN(
        n20854) );
  NAND3_X1 U30737 ( .A1(n23963), .A2(n22623), .A3(n23955), .ZN(n23633) );
  INV_X1 U30738 ( .A(n33793), .ZN(n33638) );
  XNOR2_X1 U30739 ( .A(n33638), .B(n20856), .ZN(n43539) );
  XNOR2_X1 U30740 ( .A(n33049), .B(n20857), .ZN(n20858) );
  XNOR2_X1 U30741 ( .A(n25134), .B(n20858), .ZN(n44136) );
  XNOR2_X1 U30742 ( .A(n43539), .B(n44136), .ZN(n20859) );
  XNOR2_X1 U30743 ( .A(n51424), .B(n20859), .ZN(n20860) );
  NOR2_X1 U30744 ( .A1(n21756), .A2(n21755), .ZN(n22260) );
  OAI21_X1 U30745 ( .B1(n21758), .B2(n629), .A(n23338), .ZN(n20861) );
  NAND3_X1 U30746 ( .A1(n20861), .A2(n21756), .A3(n23334), .ZN(n20862) );
  AND2_X1 U30747 ( .A1(n20862), .A2(n20863), .ZN(n20871) );
  NAND2_X1 U30748 ( .A1(n21737), .A2(n1024), .ZN(n20867) );
  AOI21_X1 U30749 ( .B1(n21756), .B2(n23336), .A(n629), .ZN(n20864) );
  OAI21_X1 U30750 ( .B1(n21756), .B2(n23341), .A(n20868), .ZN(n23343) );
  NAND2_X1 U30752 ( .A1(n24237), .A2(n21810), .ZN(n24246) );
  INV_X1 U30753 ( .A(n24246), .ZN(n21806) );
  NAND4_X1 U30754 ( .A1(n21806), .A2(n24238), .A3(n24247), .A4(n24245), .ZN(
        n20874) );
  NAND4_X1 U30755 ( .A1(n20872), .A2(n24250), .A3(n23784), .A4(n23785), .ZN(
        n20873) );
  AND2_X1 U30756 ( .A1(n20873), .A2(n20874), .ZN(n20885) );
  NAND3_X1 U30757 ( .A1(n20875), .A2(n21810), .A3(n21820), .ZN(n20878) );
  NAND4_X1 U30758 ( .A1(n24239), .A2(n21811), .A3(n24238), .A4(n21823), .ZN(
        n20877) );
  AND2_X1 U30759 ( .A1(n20877), .A2(n20878), .ZN(n20884) );
  XNOR2_X1 U30760 ( .A(n24245), .B(n21820), .ZN(n20880) );
  OAI211_X1 U30761 ( .C1(n20880), .C2(n6744), .A(n20879), .B(n23785), .ZN(
        n20883) );
  OAI21_X1 U30762 ( .B1(n23455), .B2(n21820), .A(n20881), .ZN(n20882) );
  NAND2_X1 U30763 ( .A1(n23414), .A2(n2676), .ZN(n20888) );
  OAI21_X1 U30764 ( .B1(n22045), .B2(n20889), .A(n23411), .ZN(n20900) );
  AND2_X1 U30765 ( .A1(n23417), .A2(n23412), .ZN(n22050) );
  XNOR2_X1 U30766 ( .A(n23410), .B(n20890), .ZN(n20891) );
  OAI211_X1 U30767 ( .C1(n22050), .C2(n23426), .A(n452), .B(n20892), .ZN(
        n20899) );
  NAND2_X1 U30768 ( .A1(n24266), .A2(n23422), .ZN(n20898) );
  OAI21_X1 U30769 ( .B1(n23407), .B2(n22037), .A(n23411), .ZN(n20894) );
  OAI21_X1 U30770 ( .B1(n23411), .B2(n22037), .A(n22036), .ZN(n20893) );
  AOI21_X1 U30771 ( .B1(n20895), .B2(n20894), .A(n20893), .ZN(n20896) );
  OAI21_X1 U30772 ( .B1(n22037), .B2(n23424), .A(n20896), .ZN(n20897) );
  NAND2_X1 U30773 ( .A1(n20903), .A2(n23445), .ZN(n22020) );
  NOR2_X1 U30774 ( .A1(n22020), .A2(n22011), .ZN(n21328) );
  NAND2_X1 U30775 ( .A1(n22586), .A2(n22593), .ZN(n20901) );
  AOI21_X1 U30776 ( .B1(n20903), .B2(n20901), .A(n23445), .ZN(n20902) );
  NOR2_X1 U30777 ( .A1(n7689), .A2(n23442), .ZN(n22010) );
  AND2_X1 U30778 ( .A1(n23446), .A2(n23436), .ZN(n20910) );
  OAI22_X1 U30779 ( .A1(n21328), .A2(n20902), .B1(n22010), .B2(n20910), .ZN(
        n20914) );
  AND2_X1 U30780 ( .A1(n23446), .A2(n3513), .ZN(n21326) );
  NOR2_X1 U30781 ( .A1(n22586), .A2(n22593), .ZN(n20905) );
  NAND2_X1 U30782 ( .A1(n20903), .A2(n22586), .ZN(n20904) );
  AND2_X1 U30783 ( .A1(n23445), .A2(n22593), .ZN(n21325) );
  AOI22_X1 U30784 ( .A1(n21326), .A2(n20905), .B1(n20904), .B2(n21325), .ZN(
        n20913) );
  NOR2_X1 U30785 ( .A1(n23445), .A2(n22586), .ZN(n21329) );
  NOR2_X1 U30786 ( .A1(n5609), .A2(n22593), .ZN(n20906) );
  OAI21_X1 U30787 ( .B1(n21329), .B2(n20906), .A(n3513), .ZN(n20909) );
  OAI21_X1 U30788 ( .B1(n23445), .B2(n22593), .A(n23442), .ZN(n20907) );
  AOI21_X1 U30789 ( .B1(n23446), .B2(n22586), .A(n20907), .ZN(n20908) );
  OAI211_X1 U30790 ( .C1(n3513), .C2(n23441), .A(n20909), .B(n20908), .ZN(
        n20912) );
  NAND2_X1 U30791 ( .A1(n20910), .A2(n22593), .ZN(n20911) );
  NOR2_X1 U30792 ( .A1(n22445), .A2(n22434), .ZN(n20916) );
  NAND2_X1 U30793 ( .A1(n22978), .A2(n22995), .ZN(n20915) );
  OAI211_X1 U30794 ( .C1(n22562), .C2(n22985), .A(n20916), .B(n20915), .ZN(
        n20927) );
  OR2_X1 U30795 ( .A1(n22995), .A2(n22983), .ZN(n20917) );
  AOI21_X1 U30796 ( .B1(n20918), .B2(n20917), .A(n22989), .ZN(n20926) );
  NAND4_X1 U30797 ( .A1(n22979), .A2(n22978), .A3(n22557), .A4(n3691), .ZN(
        n20921) );
  NAND2_X1 U30798 ( .A1(n22995), .A2(n22434), .ZN(n20919) );
  AND2_X1 U30799 ( .A1(n22983), .A2(n22977), .ZN(n22980) );
  NAND2_X1 U30800 ( .A1(n20919), .A2(n22980), .ZN(n20920) );
  AND2_X1 U30801 ( .A1(n20920), .A2(n20921), .ZN(n20925) );
  NAND3_X1 U30802 ( .A1(n22436), .A2(n22557), .A3(n23001), .ZN(n20923) );
  INV_X1 U30803 ( .A(n22978), .ZN(n22986) );
  NAND2_X1 U30804 ( .A1(n22986), .A2(n22982), .ZN(n20922) );
  NAND2_X1 U30805 ( .A1(n22658), .A2(n23247), .ZN(n21836) );
  NAND2_X1 U30806 ( .A1(n23238), .A2(n23246), .ZN(n22653) );
  INV_X1 U30807 ( .A(n22653), .ZN(n20929) );
  INV_X1 U30809 ( .A(n23241), .ZN(n20928) );
  OAI21_X1 U30810 ( .B1(n23237), .B2(n5292), .A(n23238), .ZN(n20931) );
  NAND3_X1 U30811 ( .A1(n20931), .A2(n22123), .A3(n23254), .ZN(n20936) );
  OAI211_X1 U30812 ( .C1(n22653), .C2(n757), .A(n20932), .B(n21847), .ZN(
        n20933) );
  OAI21_X1 U30813 ( .B1(n21852), .B2(n23241), .A(n20933), .ZN(n20935) );
  NOR2_X1 U30814 ( .A1(n23254), .A2(n52133), .ZN(n23239) );
  NAND3_X1 U30815 ( .A1(n23239), .A2(n5294), .A3(n22658), .ZN(n20934) );
  NAND4_X2 U30816 ( .A1(n20937), .A2(n20935), .A3(n20936), .A4(n20934), .ZN(
        n28381) );
  XNOR2_X1 U30817 ( .A(n27424), .B(n28381), .ZN(n24716) );
  INV_X1 U30818 ( .A(n24716), .ZN(n26272) );
  XNOR2_X1 U30819 ( .A(n26272), .B(n24855), .ZN(n26013) );
  INV_X1 U30820 ( .A(n20941), .ZN(n20938) );
  OAI21_X1 U30821 ( .B1(n20938), .B2(n21780), .A(n22290), .ZN(n20951) );
  INV_X1 U30822 ( .A(n20939), .ZN(n20940) );
  OR2_X1 U30823 ( .A1(n20941), .A2(n20940), .ZN(n21786) );
  AND2_X1 U30824 ( .A1(n21782), .A2(n22701), .ZN(n21121) );
  NAND2_X1 U30825 ( .A1(n21121), .A2(n21780), .ZN(n20945) );
  OAI21_X1 U30826 ( .B1(n21779), .B2(n20948), .A(n20942), .ZN(n20949) );
  OAI211_X2 U30827 ( .C1(n21765), .C2(n20951), .A(n20950), .B(n20949), .ZN(
        n25346) );
  NAND3_X1 U30828 ( .A1(n22154), .A2(n22142), .A3(n22151), .ZN(n21938) );
  NOR2_X1 U30829 ( .A1(n20954), .A2(n20953), .ZN(n20963) );
  INV_X1 U30830 ( .A(n20958), .ZN(n20961) );
  NAND2_X1 U30831 ( .A1(n21027), .A2(n22157), .ZN(n20955) );
  NAND3_X1 U30832 ( .A1(n22145), .A2(n21026), .A3(n20952), .ZN(n20959) );
  OAI211_X1 U30833 ( .C1(n20961), .C2(n975), .A(n20960), .B(n20959), .ZN(
        n20962) );
  OAI21_X1 U30834 ( .B1(n51355), .B2(n21725), .A(n413), .ZN(n20971) );
  INV_X1 U30835 ( .A(n20965), .ZN(n20968) );
  INV_X1 U30836 ( .A(n20966), .ZN(n20967) );
  NAND3_X1 U30837 ( .A1(n20968), .A2(n20967), .A3(n2102), .ZN(n20969) );
  NAND2_X1 U30838 ( .A1(n22115), .A2(n20969), .ZN(n20970) );
  OAI21_X1 U30839 ( .B1(n20972), .B2(n20971), .A(n20970), .ZN(n20979) );
  NAND2_X1 U30840 ( .A1(n23225), .A2(n23230), .ZN(n20973) );
  NOR2_X1 U30841 ( .A1(n51355), .A2(n413), .ZN(n22406) );
  XNOR2_X1 U30842 ( .A(n23218), .B(n22121), .ZN(n20975) );
  XNOR2_X1 U30846 ( .A(n27419), .B(n24849), .ZN(n20980) );
  XNOR2_X1 U30847 ( .A(n25346), .B(n20980), .ZN(n21001) );
  AND2_X1 U30848 ( .A1(n24295), .A2(n52207), .ZN(n23511) );
  OAI21_X1 U30849 ( .B1(n21900), .B2(n52206), .A(n24295), .ZN(n20982) );
  INV_X1 U30850 ( .A(n20985), .ZN(n20986) );
  NOR2_X1 U30852 ( .A1(n23513), .A2(n21904), .ZN(n24278) );
  INV_X1 U30853 ( .A(n24278), .ZN(n20989) );
  NAND2_X1 U30854 ( .A1(n23483), .A2(n21975), .ZN(n23478) );
  NOR2_X1 U30855 ( .A1(n23480), .A2(n21975), .ZN(n21986) );
  NAND2_X1 U30856 ( .A1(n21986), .A2(n21970), .ZN(n20990) );
  NOR2_X1 U30857 ( .A1(n23489), .A2(n21970), .ZN(n21968) );
  AND2_X1 U30858 ( .A1(n23483), .A2(n23489), .ZN(n20993) );
  NAND2_X1 U30859 ( .A1(n21970), .A2(n21981), .ZN(n20997) );
  NAND4_X1 U30860 ( .A1(n20997), .A2(n20996), .A3(n21975), .A4(n20995), .ZN(
        n20998) );
  INV_X1 U30861 ( .A(n51119), .ZN(n21000) );
  XNOR2_X1 U30862 ( .A(n21001), .B(n21000), .ZN(n23688) );
  XNOR2_X1 U30863 ( .A(n26013), .B(n23688), .ZN(n21002) );
  NOR2_X1 U30864 ( .A1(n22341), .A2(n597), .ZN(n26806) );
  NAND3_X1 U30865 ( .A1(n23306), .A2(n23317), .A3(n21873), .ZN(n21003) );
  NAND2_X1 U30866 ( .A1(n21004), .A2(n21003), .ZN(n21006) );
  AOI21_X1 U30867 ( .B1(n21006), .B2(n22251), .A(n21005), .ZN(n24018) );
  NOR2_X1 U30868 ( .A1(n23317), .A2(n21873), .ZN(n22252) );
  NAND2_X1 U30869 ( .A1(n22252), .A2(n756), .ZN(n21008) );
  AOI21_X1 U30870 ( .B1(n23303), .B2(n23306), .A(n8303), .ZN(n21007) );
  NAND2_X1 U30871 ( .A1(n23316), .A2(n21873), .ZN(n22961) );
  NAND4_X1 U30872 ( .A1(n21008), .A2(n21007), .A3(n22961), .A4(n21010), .ZN(
        n21009) );
  AND2_X1 U30874 ( .A1(n23316), .A2(n441), .ZN(n22960) );
  OAI21_X1 U30875 ( .B1(n942), .B2(n23314), .A(n756), .ZN(n21011) );
  INV_X1 U30876 ( .A(n22866), .ZN(n21014) );
  OAI211_X1 U30877 ( .C1(n22859), .C2(n22857), .A(n22334), .B(n22849), .ZN(
        n21013) );
  NAND2_X1 U30878 ( .A1(n22851), .A2(n21877), .ZN(n21012) );
  NAND4_X1 U30879 ( .A1(n22328), .A2(n21014), .A3(n21013), .A4(n21012), .ZN(
        n23025) );
  NOR2_X1 U30880 ( .A1(n22851), .A2(n22861), .ZN(n22333) );
  NOR2_X1 U30881 ( .A1(n22864), .A2(n22857), .ZN(n21886) );
  OR2_X1 U30882 ( .A1(n21886), .A2(n21887), .ZN(n22855) );
  NAND2_X1 U30883 ( .A1(n22333), .A2(n22855), .ZN(n23019) );
  NAND2_X1 U30884 ( .A1(n21017), .A2(n23019), .ZN(n25039) );
  XNOR2_X1 U30885 ( .A(n26377), .B(n25039), .ZN(n24700) );
  MUX2_X1 U30886 ( .A(n21020), .B(n21019), .S(n51660), .Z(n21034) );
  NAND3_X1 U30887 ( .A1(n52381), .A2(n22142), .A3(n21026), .ZN(n21033) );
  AOI21_X1 U30888 ( .B1(n21921), .B2(n22140), .A(n51661), .ZN(n21022) );
  INV_X1 U30889 ( .A(n22141), .ZN(n21937) );
  OR2_X1 U30890 ( .A1(n21022), .A2(n21937), .ZN(n21032) );
  OAI21_X1 U30891 ( .B1(n22149), .B2(n21027), .A(n21026), .ZN(n21028) );
  OAI21_X1 U30892 ( .B1(n21030), .B2(n21029), .A(n21028), .ZN(n21031) );
  NOR2_X1 U30893 ( .A1(n21041), .A2(n22362), .ZN(n21035) );
  NOR2_X1 U30894 ( .A1(n21036), .A2(n21035), .ZN(n21046) );
  NOR2_X1 U30895 ( .A1(n22908), .A2(n22901), .ZN(n21039) );
  NAND4_X1 U30897 ( .A1(n21041), .A2(n22165), .A3(n21040), .A4(n22919), .ZN(
        n21044) );
  NAND2_X1 U30898 ( .A1(n5737), .A2(n22919), .ZN(n22348) );
  OAI21_X1 U30899 ( .B1(n22348), .B2(n22901), .A(n22169), .ZN(n21042) );
  NAND2_X1 U30900 ( .A1(n22913), .A2(n21042), .ZN(n21043) );
  NAND4_X2 U30901 ( .A1(n21046), .A2(n21045), .A3(n21044), .A4(n21043), .ZN(
        n28274) );
  XNOR2_X1 U30902 ( .A(n27235), .B(n24700), .ZN(n23719) );
  INV_X1 U30903 ( .A(n23719), .ZN(n21080) );
  INV_X1 U30904 ( .A(n23409), .ZN(n22035) );
  NAND2_X1 U30905 ( .A1(n22035), .A2(n452), .ZN(n21048) );
  INV_X1 U30906 ( .A(n22046), .ZN(n21051) );
  NAND2_X1 U30907 ( .A1(n21051), .A2(n23407), .ZN(n21047) );
  NAND2_X1 U30908 ( .A1(n21049), .A2(n23414), .ZN(n21059) );
  INV_X1 U30909 ( .A(n23408), .ZN(n21050) );
  OAI21_X1 U30910 ( .B1(n2676), .B2(n23411), .A(n23417), .ZN(n21052) );
  NAND2_X1 U30911 ( .A1(n21052), .A2(n21051), .ZN(n21057) );
  NAND2_X1 U30912 ( .A1(n21053), .A2(n22320), .ZN(n21055) );
  NAND2_X1 U30913 ( .A1(n23417), .A2(n23409), .ZN(n21054) );
  NAND4_X1 U30914 ( .A1(n21055), .A2(n23410), .A3(n23426), .A4(n21054), .ZN(
        n21056) );
  OR2_X1 U30915 ( .A1(n22375), .A2(n50976), .ZN(n22732) );
  OAI21_X1 U30916 ( .B1(n22298), .B2(n22736), .A(n5371), .ZN(n21061) );
  NAND2_X1 U30917 ( .A1(n22386), .A2(n51753), .ZN(n21060) );
  NAND2_X1 U30918 ( .A1(n50977), .A2(n22390), .ZN(n22373) );
  XNOR2_X1 U30919 ( .A(n26147), .B(n26152), .ZN(n21079) );
  NAND2_X1 U30920 ( .A1(n22835), .A2(n22832), .ZN(n21064) );
  NAND4_X1 U30921 ( .A1(n21066), .A2(n22508), .A3(n21065), .A4(n21064), .ZN(
        n24258) );
  NAND2_X1 U30922 ( .A1(n24258), .A2(n22223), .ZN(n21078) );
  AOI21_X1 U30923 ( .B1(n21068), .B2(n22831), .A(n22491), .ZN(n24255) );
  INV_X1 U30924 ( .A(n24255), .ZN(n21069) );
  NAND2_X1 U30925 ( .A1(n24258), .A2(n21069), .ZN(n21077) );
  OR2_X1 U30927 ( .A1(n22832), .A2(n22506), .ZN(n22827) );
  INV_X1 U30928 ( .A(n22827), .ZN(n21072) );
  OR2_X1 U30929 ( .A1(n21072), .A2(n22826), .ZN(n21075) );
  NOR2_X1 U30930 ( .A1(n21074), .A2(n22830), .ZN(n22224) );
  AND2_X1 U30931 ( .A1(n22224), .A2(n21075), .ZN(n24259) );
  INV_X1 U30932 ( .A(n24259), .ZN(n21076) );
  NAND4_X1 U30933 ( .A1(n21078), .A2(n21077), .A3(n24256), .A4(n21076), .ZN(
        n25996) );
  XNOR2_X1 U30934 ( .A(n21079), .B(n25996), .ZN(n23718) );
  AND2_X1 U30935 ( .A1(n24290), .A2(n52207), .ZN(n21081) );
  NAND2_X1 U30936 ( .A1(n23504), .A2(n23513), .ZN(n24279) );
  INV_X1 U30937 ( .A(n21083), .ZN(n21084) );
  NAND3_X1 U30938 ( .A1(n7247), .A2(n24287), .A3(n52207), .ZN(n21909) );
  AND2_X1 U30939 ( .A1(n21084), .A2(n21909), .ZN(n21087) );
  NOR2_X1 U30940 ( .A1(n24290), .A2(n52206), .ZN(n21908) );
  NOR2_X1 U30941 ( .A1(n24283), .A2(n24287), .ZN(n21907) );
  XNOR2_X1 U30942 ( .A(n21090), .B(n21089), .ZN(n43786) );
  XNOR2_X1 U30943 ( .A(n25115), .B(n25040), .ZN(n42477) );
  XNOR2_X1 U30944 ( .A(n42477), .B(n21091), .ZN(n21092) );
  XNOR2_X1 U30945 ( .A(n43786), .B(n21092), .ZN(n21093) );
  XNOR2_X1 U30946 ( .A(n24905), .B(n21093), .ZN(n21112) );
  NOR2_X1 U30947 ( .A1(n21095), .A2(n21106), .ZN(n21709) );
  NAND2_X1 U30948 ( .A1(n52048), .A2(n21714), .ZN(n21096) );
  NOR2_X1 U30949 ( .A1(n22186), .A2(n21096), .ZN(n21097) );
  NOR2_X1 U30950 ( .A1(n21709), .A2(n21097), .ZN(n21103) );
  INV_X1 U30951 ( .A(n22191), .ZN(n21099) );
  OAI21_X1 U30952 ( .B1(n21700), .B2(n21713), .A(n21712), .ZN(n21098) );
  NAND4_X1 U30953 ( .A1(n21100), .A2(n21099), .A3(n21106), .A4(n21098), .ZN(
        n21102) );
  NOR2_X1 U30954 ( .A1(n21104), .A2(n21700), .ZN(n21109) );
  NOR2_X1 U30955 ( .A1(n21715), .A2(n21700), .ZN(n21108) );
  NAND2_X1 U30956 ( .A1(n21105), .A2(n52048), .ZN(n22180) );
  OAI21_X1 U30957 ( .B1(n7119), .B2(n21106), .A(n22180), .ZN(n21107) );
  AOI22_X1 U30958 ( .A1(n21110), .A2(n21109), .B1(n21108), .B2(n21107), .ZN(
        n21111) );
  XNOR2_X1 U30959 ( .A(n24891), .B(n24430), .ZN(n25306) );
  XNOR2_X1 U30960 ( .A(n25306), .B(n21112), .ZN(n21138) );
  NAND2_X1 U30961 ( .A1(n21782), .A2(n22702), .ZN(n21113) );
  INV_X1 U30962 ( .A(n21115), .ZN(n21775) );
  NAND2_X1 U30963 ( .A1(n21116), .A2(n21117), .ZN(n21119) );
  OAI21_X1 U30964 ( .B1(n21117), .B2(n21767), .A(n51080), .ZN(n21118) );
  NAND4_X1 U30965 ( .A1(n21120), .A2(n21782), .A3(n21119), .A4(n21118), .ZN(
        n21128) );
  INV_X1 U30966 ( .A(n22290), .ZN(n21771) );
  INV_X1 U30967 ( .A(n21121), .ZN(n21124) );
  AND2_X1 U30968 ( .A1(n21122), .A2(n22702), .ZN(n21123) );
  OAI211_X1 U30969 ( .C1(n21125), .C2(n21782), .A(n21124), .B(n21123), .ZN(
        n21126) );
  NAND4_X2 U30970 ( .A1(n21127), .A2(n21129), .A3(n21128), .A4(n21126), .ZN(
        n25249) );
  NAND3_X1 U30971 ( .A1(n22306), .A2(n22470), .A3(n22464), .ZN(n22466) );
  OAI211_X1 U30972 ( .C1(n2083), .C2(n22464), .A(n22478), .B(n21130), .ZN(
        n21133) );
  NAND3_X1 U30973 ( .A1(n22476), .A2(n51124), .A3(n2083), .ZN(n21132) );
  OAI21_X1 U30974 ( .B1(n22715), .B2(n22462), .A(n22308), .ZN(n21135) );
  NOR2_X1 U30975 ( .A1(n22464), .A2(n22479), .ZN(n22458) );
  OAI211_X1 U30976 ( .C1(n22458), .C2(n22306), .A(n22717), .B(n22481), .ZN(
        n21134) );
  NAND2_X1 U30977 ( .A1(n21135), .A2(n21134), .ZN(n21136) );
  XNOR2_X2 U30978 ( .A(n25249), .B(n25050), .ZN(n28276) );
  XNOR2_X1 U30979 ( .A(n21138), .B(n28276), .ZN(n21139) );
  AOI21_X1 U30981 ( .B1(n21144), .B2(n21758), .A(n51200), .ZN(n21142) );
  NAND2_X1 U30982 ( .A1(n21756), .A2(n21144), .ZN(n21141) );
  OAI21_X1 U30983 ( .B1(n21737), .B2(n1024), .A(n22256), .ZN(n21146) );
  NAND2_X1 U30984 ( .A1(n21147), .A2(n21146), .ZN(n23008) );
  NAND2_X1 U30985 ( .A1(n22260), .A2(n21148), .ZN(n23332) );
  OAI21_X1 U30987 ( .B1(n23334), .B2(n23336), .A(n1024), .ZN(n21149) );
  NAND2_X1 U30989 ( .A1(n23007), .A2(n23013), .ZN(n23290) );
  NOR3_X1 U30990 ( .A1(n23547), .A2(n21155), .A3(n23360), .ZN(n23552) );
  NAND2_X1 U30991 ( .A1(n23552), .A2(n51677), .ZN(n21152) );
  OAI21_X1 U30992 ( .B1(n22275), .B2(n21155), .A(n23364), .ZN(n21151) );
  AND2_X1 U30993 ( .A1(n21152), .A2(n21151), .ZN(n21161) );
  NAND2_X1 U30994 ( .A1(n23563), .A2(n23568), .ZN(n23566) );
  MUX2_X1 U30995 ( .A(n23566), .B(n23574), .S(n23351), .Z(n21160) );
  NOR2_X1 U30996 ( .A1(n23563), .A2(n23568), .ZN(n21153) );
  NOR2_X1 U30997 ( .A1(n21154), .A2(n21153), .ZN(n21158) );
  AND2_X1 U30998 ( .A1(n21156), .A2(n21155), .ZN(n23559) );
  NOR2_X1 U30999 ( .A1(n51675), .A2(n23546), .ZN(n23569) );
  NOR2_X1 U31000 ( .A1(n23472), .A2(n21953), .ZN(n21162) );
  NAND3_X1 U31001 ( .A1(n21163), .A2(n21162), .A3(n23150), .ZN(n21170) );
  OAI21_X1 U31002 ( .B1(n23154), .B2(n23466), .A(n21164), .ZN(n21165) );
  AOI21_X1 U31003 ( .B1(n23472), .B2(n21166), .A(n21165), .ZN(n21169) );
  INV_X1 U31004 ( .A(n21946), .ZN(n23471) );
  OAI21_X1 U31005 ( .B1(n23467), .B2(n51123), .A(n21947), .ZN(n23158) );
  NAND2_X1 U31006 ( .A1(n23471), .A2(n23158), .ZN(n21168) );
  NAND4_X2 U31007 ( .A1(n21169), .A2(n21170), .A3(n21168), .A4(n21167), .ZN(
        n27224) );
  INV_X1 U31008 ( .A(n21175), .ZN(n21176) );
  NAND3_X1 U31009 ( .A1(n5271), .A2(n21177), .A3(n21176), .ZN(n21179) );
  MUX2_X1 U31010 ( .A(n21179), .B(n21178), .S(n21185), .Z(n21192) );
  INV_X1 U31011 ( .A(n21180), .ZN(n21184) );
  NAND2_X1 U31012 ( .A1(n21182), .A2(n21181), .ZN(n21183) );
  OAI211_X1 U31013 ( .C1(n21186), .C2(n21185), .A(n21184), .B(n21183), .ZN(
        n21191) );
  INV_X1 U31014 ( .A(n21187), .ZN(n21189) );
  NAND2_X1 U31015 ( .A1(n21189), .A2(n21188), .ZN(n21190) );
  INV_X1 U31016 ( .A(n21194), .ZN(n21195) );
  NAND3_X1 U31017 ( .A1(n21199), .A2(n21198), .A3(n21197), .ZN(n21203) );
  NAND2_X1 U31018 ( .A1(n21201), .A2(n21200), .ZN(n21202) );
  AOI21_X1 U31019 ( .B1(n21204), .B2(n21203), .A(n21202), .ZN(n21207) );
  INV_X1 U31020 ( .A(n21205), .ZN(n21206) );
  NOR2_X1 U31021 ( .A1(n21207), .A2(n21206), .ZN(n21221) );
  INV_X1 U31022 ( .A(n21218), .ZN(n21210) );
  OAI21_X1 U31023 ( .B1(n21210), .B2(n21209), .A(n21208), .ZN(n21220) );
  INV_X1 U31024 ( .A(n21211), .ZN(n21217) );
  OAI22_X1 U31025 ( .A1(n21215), .A2(n21214), .B1(n21213), .B2(n2229), .ZN(
        n21216) );
  NAND3_X1 U31026 ( .A1(n21218), .A2(n21217), .A3(n21216), .ZN(n21219) );
  OAI22_X1 U31027 ( .A1(n21232), .A2(n21223), .B1(n21222), .B2(n21227), .ZN(
        n21226) );
  NOR2_X1 U31028 ( .A1(n21224), .A2(n21230), .ZN(n21225) );
  NOR2_X1 U31029 ( .A1(n21226), .A2(n21225), .ZN(n21241) );
  NAND2_X1 U31030 ( .A1(n761), .A2(n21227), .ZN(n21228) );
  OAI21_X1 U31031 ( .B1(n21234), .B2(n21233), .A(n21232), .ZN(n21236) );
  OAI21_X1 U31032 ( .B1(n21237), .B2(n21236), .A(n21235), .ZN(n21238) );
  INV_X1 U31033 ( .A(n22061), .ZN(n23166) );
  NAND2_X1 U31034 ( .A1(n21243), .A2(n21242), .ZN(n21247) );
  OAI21_X1 U31035 ( .B1(n21254), .B2(n51132), .A(n21244), .ZN(n21246) );
  MUX2_X1 U31036 ( .A(n21247), .B(n21246), .S(n21245), .Z(n21261) );
  AOI22_X1 U31037 ( .A1(n21250), .A2(n21254), .B1(n21249), .B2(n21248), .ZN(
        n21260) );
  NOR2_X1 U31038 ( .A1(n21252), .A2(n51132), .ZN(n21255) );
  NAND2_X1 U31039 ( .A1(n21257), .A2(n21256), .ZN(n21258) );
  NAND4_X2 U31040 ( .A1(n21261), .A2(n21260), .A3(n21259), .A4(n21258), .ZN(
        n23167) );
  INV_X1 U31041 ( .A(n23167), .ZN(n22674) );
  INV_X1 U31042 ( .A(n21262), .ZN(n21267) );
  INV_X1 U31043 ( .A(n21263), .ZN(n21266) );
  INV_X1 U31044 ( .A(n21264), .ZN(n21265) );
  AOI21_X1 U31045 ( .B1(n21267), .B2(n21266), .A(n21265), .ZN(n21278) );
  INV_X1 U31046 ( .A(n21268), .ZN(n21275) );
  NAND3_X1 U31047 ( .A1(n21271), .A2(n21270), .A3(n21269), .ZN(n21274) );
  NAND3_X1 U31048 ( .A1(n5229), .A2(n21272), .A3(n21287), .ZN(n21273) );
  OAI211_X1 U31049 ( .C1(n21276), .C2(n21275), .A(n21274), .B(n21273), .ZN(
        n21277) );
  NOR2_X1 U31050 ( .A1(n21278), .A2(n21277), .ZN(n21289) );
  INV_X1 U31051 ( .A(n21279), .ZN(n21280) );
  NAND2_X1 U31052 ( .A1(n21281), .A2(n21280), .ZN(n21288) );
  OAI21_X1 U31053 ( .B1(n21284), .B2(n21283), .A(n21282), .ZN(n21285) );
  INV_X1 U31054 ( .A(n21290), .ZN(n21292) );
  AOI22_X1 U31055 ( .A1(n21292), .A2(n21296), .B1(n21291), .B2(n21293), .ZN(
        n21299) );
  OAI21_X1 U31056 ( .B1(n21295), .B2(n21302), .A(n21294), .ZN(n21297) );
  INV_X1 U31057 ( .A(n21301), .ZN(n21307) );
  AOI21_X1 U31058 ( .B1(n21308), .B2(n21307), .A(n21306), .ZN(n22543) );
  NOR2_X1 U31059 ( .A1(n23182), .A2(n23167), .ZN(n22785) );
  INV_X1 U31060 ( .A(n22785), .ZN(n21309) );
  OAI21_X1 U31061 ( .B1(n21309), .B2(n5269), .A(n23183), .ZN(n21310) );
  OR2_X1 U31062 ( .A1(n23175), .A2(n23166), .ZN(n22058) );
  NAND2_X1 U31063 ( .A1(n21311), .A2(n23184), .ZN(n21312) );
  AND2_X1 U31064 ( .A1(n51021), .A2(n23182), .ZN(n23170) );
  NAND2_X1 U31065 ( .A1(n23170), .A2(n23178), .ZN(n22068) );
  OAI21_X1 U31066 ( .B1(n21314), .B2(n23175), .A(n22055), .ZN(n21315) );
  AND2_X1 U31067 ( .A1(n23178), .A2(n7811), .ZN(n22536) );
  NAND2_X1 U31068 ( .A1(n21315), .A2(n22536), .ZN(n21316) );
  AOI21_X1 U31069 ( .B1(n22019), .B2(n3513), .A(n21319), .ZN(n21324) );
  AOI22_X1 U31070 ( .A1(n23433), .A2(n23436), .B1(n23446), .B2(n23442), .ZN(
        n21323) );
  NAND2_X1 U31072 ( .A1(n3513), .A2(n23445), .ZN(n21321) );
  NAND4_X1 U31073 ( .A1(n21319), .A2(n23434), .A3(n3513), .A4(n22593), .ZN(
        n21320) );
  OAI21_X1 U31074 ( .B1(n22009), .B2(n21321), .A(n21320), .ZN(n21322) );
  AOI21_X1 U31075 ( .B1(n21324), .B2(n21323), .A(n21322), .ZN(n21333) );
  INV_X1 U31076 ( .A(n23441), .ZN(n22591) );
  AOI22_X1 U31077 ( .A1(n22591), .A2(n21326), .B1(n21325), .B2(n22586), .ZN(
        n21332) );
  OAI21_X1 U31078 ( .B1(n23436), .B2(n22586), .A(n22023), .ZN(n21327) );
  NAND2_X1 U31079 ( .A1(n21328), .A2(n21327), .ZN(n21331) );
  NAND2_X1 U31080 ( .A1(n22008), .A2(n22010), .ZN(n21330) );
  NAND2_X1 U31081 ( .A1(n21977), .A2(n21981), .ZN(n21334) );
  OAI22_X1 U31082 ( .A1(n23489), .A2(n21334), .B1(n21977), .B2(n21981), .ZN(
        n21338) );
  AND2_X1 U31083 ( .A1(n23483), .A2(n2130), .ZN(n21337) );
  NAND2_X1 U31084 ( .A1(n23480), .A2(n8076), .ZN(n23482) );
  NAND3_X1 U31085 ( .A1(n21975), .A2(n2130), .A3(n23479), .ZN(n21335) );
  OAI21_X1 U31086 ( .B1(n23482), .B2(n23483), .A(n21335), .ZN(n21336) );
  AOI22_X1 U31087 ( .A1(n21338), .A2(n21337), .B1(n21336), .B2(n23489), .ZN(
        n21348) );
  NAND3_X1 U31088 ( .A1(n21339), .A2(n23489), .A3(n21986), .ZN(n21340) );
  AND2_X1 U31089 ( .A1(n21341), .A2(n21340), .ZN(n21347) );
  NOR2_X1 U31090 ( .A1(n23489), .A2(n23477), .ZN(n21342) );
  NOR2_X1 U31091 ( .A1(n21342), .A2(n21983), .ZN(n21346) );
  INV_X1 U31092 ( .A(n21343), .ZN(n21344) );
  NAND3_X1 U31093 ( .A1(n21344), .A2(n21975), .A3(n23482), .ZN(n21345) );
  NOR2_X1 U31094 ( .A1(n21362), .A2(n21354), .ZN(n21357) );
  AOI22_X1 U31095 ( .A1(n21358), .A2(n21357), .B1(n21356), .B2(n21355), .ZN(
        n21367) );
  OAI22_X1 U31096 ( .A1(n21361), .A2(n20768), .B1(n21360), .B2(n21359), .ZN(
        n21363) );
  NAND2_X1 U31097 ( .A1(n21363), .A2(n21362), .ZN(n21366) );
  NAND2_X1 U31098 ( .A1(n762), .A2(n21364), .ZN(n21365) );
  NAND4_X2 U31099 ( .A1(n21368), .A2(n21367), .A3(n21366), .A4(n21365), .ZN(
        n23142) );
  NAND2_X1 U31100 ( .A1(n21370), .A2(n21369), .ZN(n21371) );
  INV_X1 U31101 ( .A(n21374), .ZN(n21378) );
  INV_X1 U31102 ( .A(n21375), .ZN(n21376) );
  NAND2_X1 U31103 ( .A1(n2257), .A2(n21388), .ZN(n21379) );
  NOR2_X1 U31104 ( .A1(n21396), .A2(n358), .ZN(n21387) );
  INV_X1 U31105 ( .A(n21383), .ZN(n21384) );
  AOI22_X1 U31106 ( .A1(n21387), .A2(n21386), .B1(n21385), .B2(n21384), .ZN(
        n21401) );
  NOR2_X1 U31107 ( .A1(n21398), .A2(n21390), .ZN(n21395) );
  AOI21_X1 U31108 ( .B1(n21393), .B2(n581), .A(n358), .ZN(n21394) );
  OAI21_X1 U31109 ( .B1(n21395), .B2(n21394), .A(n1860), .ZN(n21400) );
  NAND3_X1 U31110 ( .A1(n21398), .A2(n21397), .A3(n21396), .ZN(n21399) );
  INV_X1 U31111 ( .A(n21402), .ZN(n21411) );
  NAND2_X1 U31112 ( .A1(n21403), .A2(n21555), .ZN(n21405) );
  NAND2_X1 U31113 ( .A1(n21407), .A2(n21406), .ZN(n21408) );
  NAND4_X1 U31114 ( .A1(n21411), .A2(n21410), .A3(n21409), .A4(n21408), .ZN(
        n21419) );
  NAND2_X1 U31115 ( .A1(n21413), .A2(n21412), .ZN(n21417) );
  XNOR2_X1 U31116 ( .A(n51710), .B(n21578), .ZN(n21416) );
  OAI211_X1 U31117 ( .C1(n18823), .C2(n21584), .A(n21568), .B(n51755), .ZN(
        n21415) );
  OAI22_X1 U31118 ( .A1(n21417), .A2(n21576), .B1(n21416), .B2(n21415), .ZN(
        n21418) );
  OR2_X2 U31119 ( .A1(n21419), .A2(n21418), .ZN(n23895) );
  OR2_X1 U31120 ( .A1(n23141), .A2(n23895), .ZN(n21503) );
  OAI211_X1 U31121 ( .C1(n21423), .C2(n21422), .A(n21421), .B(n21420), .ZN(
        n21434) );
  NOR2_X1 U31122 ( .A1(n21425), .A2(n21424), .ZN(n21428) );
  OAI21_X1 U31123 ( .B1(n21428), .B2(n21427), .A(n21426), .ZN(n21433) );
  NAND2_X1 U31124 ( .A1(n21430), .A2(n21429), .ZN(n21431) );
  NOR2_X1 U31125 ( .A1(n21435), .A2(n3493), .ZN(n21437) );
  OAI21_X1 U31126 ( .B1(n21438), .B2(n21437), .A(n4433), .ZN(n21447) );
  NAND2_X1 U31127 ( .A1(n21440), .A2(n21439), .ZN(n21446) );
  NAND3_X1 U31128 ( .A1(n21443), .A2(n21442), .A3(n52139), .ZN(n21445) );
  NAND4_X1 U31129 ( .A1(n21447), .A2(n21446), .A3(n21445), .A4(n21444), .ZN(
        n21448) );
  NAND2_X1 U31130 ( .A1(n21449), .A2(n21463), .ZN(n21454) );
  NAND2_X1 U31131 ( .A1(n21451), .A2(n21450), .ZN(n21453) );
  AOI21_X1 U31132 ( .B1(n21454), .B2(n21453), .A(n21452), .ZN(n21456) );
  INV_X1 U31133 ( .A(n21458), .ZN(n21461) );
  AOI21_X1 U31135 ( .B1(n21464), .B2(n21463), .A(n1618), .ZN(n21467) );
  OAI21_X1 U31136 ( .B1(n21467), .B2(n21466), .A(n21465), .ZN(n21472) );
  AOI21_X1 U31137 ( .B1(n21470), .B2(n21469), .A(n21468), .ZN(n21471) );
  OAI211_X1 U31138 ( .C1(n21474), .C2(n21473), .A(n21472), .B(n21471), .ZN(
        n21476) );
  NAND2_X1 U31139 ( .A1(n23924), .A2(n22521), .ZN(n23898) );
  OAI21_X1 U31141 ( .B1(n23902), .B2(n23143), .A(n23913), .ZN(n21501) );
  OAI211_X1 U31142 ( .C1(n21483), .C2(n2221), .A(n21482), .B(n51754), .ZN(
        n21489) );
  NAND2_X1 U31143 ( .A1(n2220), .A2(n21483), .ZN(n21488) );
  NAND3_X1 U31144 ( .A1(n763), .A2(n21486), .A3(n21485), .ZN(n21487) );
  AND3_X1 U31145 ( .A1(n21489), .A2(n21488), .A3(n21487), .ZN(n21499) );
  INV_X1 U31146 ( .A(n21490), .ZN(n21493) );
  OAI211_X1 U31147 ( .C1(n21494), .C2(n21493), .A(n21492), .B(n21491), .ZN(
        n21498) );
  NAND2_X1 U31148 ( .A1(n21496), .A2(n21495), .ZN(n21497) );
  NAND3_X1 U31149 ( .A1(n22524), .A2(n21501), .A3(n23906), .ZN(n23901) );
  OAI211_X1 U31150 ( .C1(n21503), .C2(n23898), .A(n21502), .B(n23901), .ZN(
        n21504) );
  NAND2_X1 U31151 ( .A1(n23135), .A2(n23142), .ZN(n22801) );
  OR2_X1 U31152 ( .A1(n51033), .A2(n22521), .ZN(n21505) );
  NOR2_X1 U31153 ( .A1(n22801), .A2(n21505), .ZN(n22685) );
  NAND2_X1 U31155 ( .A1(n51034), .A2(n23143), .ZN(n22682) );
  NOR2_X1 U31156 ( .A1(n23923), .A2(n22682), .ZN(n21506) );
  NOR2_X1 U31157 ( .A1(n22685), .A2(n21506), .ZN(n21511) );
  INV_X1 U31158 ( .A(n23136), .ZN(n22523) );
  OR2_X1 U31159 ( .A1(n23141), .A2(n23906), .ZN(n21508) );
  XNOR2_X1 U31160 ( .A(n23924), .B(n23142), .ZN(n21507) );
  NAND4_X1 U31161 ( .A1(n21508), .A2(n23143), .A3(n21507), .A4(n23923), .ZN(
        n21509) );
  NOR2_X1 U31163 ( .A1(n21514), .A2(n21513), .ZN(n21516) );
  OAI21_X1 U31164 ( .B1(n21517), .B2(n21516), .A(n21515), .ZN(n21532) );
  INV_X1 U31165 ( .A(n21518), .ZN(n21522) );
  NAND2_X1 U31166 ( .A1(n21523), .A2(n20611), .ZN(n21529) );
  NAND2_X1 U31167 ( .A1(n21525), .A2(n21524), .ZN(n21526) );
  NAND2_X1 U31168 ( .A1(n18495), .A2(n51485), .ZN(n21535) );
  OAI211_X1 U31169 ( .C1(n21538), .C2(n21537), .A(n21536), .B(n21535), .ZN(
        n21539) );
  INV_X1 U31170 ( .A(n21539), .ZN(n21554) );
  NAND3_X1 U31171 ( .A1(n21544), .A2(n21543), .A3(n21542), .ZN(n21545) );
  AND2_X1 U31172 ( .A1(n21546), .A2(n21545), .ZN(n21553) );
  NAND2_X1 U31173 ( .A1(n21550), .A2(n51129), .ZN(n21551) );
  OAI22_X1 U31174 ( .A1(n21557), .A2(n21556), .B1(n21569), .B2(n21555), .ZN(
        n21562) );
  INV_X1 U31175 ( .A(n21558), .ZN(n21561) );
  OAI211_X1 U31176 ( .C1(n21562), .C2(n21561), .A(n21560), .B(n21559), .ZN(
        n21590) );
  NAND4_X1 U31177 ( .A1(n21563), .A2(n21566), .A3(n21568), .A4(n21584), .ZN(
        n21573) );
  NAND3_X1 U31178 ( .A1(n21565), .A2(n21564), .A3(n21580), .ZN(n21572) );
  NAND3_X1 U31179 ( .A1(n21567), .A2(n21566), .A3(n18823), .ZN(n21571) );
  NAND4_X1 U31180 ( .A1(n21569), .A2(n51711), .A3(n21578), .A4(n21568), .ZN(
        n21570) );
  OAI21_X1 U31181 ( .B1(n21576), .B2(n21575), .A(n21574), .ZN(n21577) );
  INV_X1 U31182 ( .A(n21577), .ZN(n21588) );
  AOI21_X1 U31183 ( .B1(n21580), .B2(n51710), .A(n21578), .ZN(n21585) );
  INV_X1 U31184 ( .A(n21581), .ZN(n21582) );
  NAND2_X1 U31185 ( .A1(n21586), .A2(n5167), .ZN(n21587) );
  OAI211_X1 U31188 ( .C1(n21600), .C2(n21604), .A(n21599), .B(n21598), .ZN(
        n21602) );
  NAND2_X1 U31189 ( .A1(n21602), .A2(n21601), .ZN(n21610) );
  NAND2_X1 U31190 ( .A1(n21604), .A2(n21603), .ZN(n21606) );
  AOI21_X1 U31191 ( .B1(n21607), .B2(n21606), .A(n52208), .ZN(n21608) );
  AOI21_X1 U31192 ( .B1(n21610), .B2(n21609), .A(n21608), .ZN(n21611) );
  NAND2_X1 U31194 ( .A1(n21613), .A2(n21614), .ZN(n21616) );
  OAI211_X1 U31195 ( .C1(n21618), .C2(n21617), .A(n21616), .B(n21615), .ZN(
        n21621) );
  NAND3_X1 U31196 ( .A1(n21621), .A2(n21620), .A3(n21619), .ZN(n21627) );
  INV_X1 U31197 ( .A(n21622), .ZN(n21623) );
  NAND3_X1 U31198 ( .A1(n21638), .A2(n21624), .A3(n21623), .ZN(n21625) );
  NAND2_X1 U31199 ( .A1(n21628), .A2(n21639), .ZN(n21643) );
  OAI21_X1 U31200 ( .B1(n21631), .B2(n21630), .A(n21629), .ZN(n21635) );
  AND2_X1 U31201 ( .A1(n21633), .A2(n21632), .ZN(n21634) );
  INV_X1 U31202 ( .A(n21638), .ZN(n21640) );
  NAND2_X1 U31203 ( .A1(n21640), .A2(n21639), .ZN(n21641) );
  AND2_X1 U31204 ( .A1(n24105), .A2(n24413), .ZN(n23736) );
  INV_X1 U31205 ( .A(n23736), .ZN(n21645) );
  NOR2_X1 U31206 ( .A1(n21647), .A2(n21646), .ZN(n21651) );
  NOR2_X1 U31207 ( .A1(n21648), .A2(n21660), .ZN(n21650) );
  OAI21_X1 U31208 ( .B1(n21651), .B2(n21650), .A(n21649), .ZN(n21668) );
  INV_X1 U31209 ( .A(n21655), .ZN(n21659) );
  NOR2_X1 U31210 ( .A1(n21664), .A2(n21656), .ZN(n21658) );
  OAI21_X1 U31211 ( .B1(n21659), .B2(n21658), .A(n21657), .ZN(n21666) );
  NAND2_X1 U31212 ( .A1(n21661), .A2(n21660), .ZN(n21662) );
  OAI211_X1 U31213 ( .C1(n21657), .C2(n21664), .A(n21663), .B(n21662), .ZN(
        n21665) );
  NAND2_X1 U31214 ( .A1(n24117), .A2(n51001), .ZN(n21669) );
  NOR2_X1 U31215 ( .A1(n23521), .A2(n21669), .ZN(n21670) );
  INV_X1 U31216 ( .A(n24074), .ZN(n23124) );
  OAI21_X1 U31217 ( .B1(n21670), .B2(n23124), .A(n24413), .ZN(n21678) );
  INV_X1 U31218 ( .A(n23129), .ZN(n24098) );
  NAND2_X1 U31219 ( .A1(n24105), .A2(n24098), .ZN(n24071) );
  NAND2_X1 U31220 ( .A1(n51001), .A2(n24098), .ZN(n21672) );
  NAND3_X1 U31221 ( .A1(n23730), .A2(n24071), .A3(n21672), .ZN(n21673) );
  AND2_X1 U31222 ( .A1(n21673), .A2(n21674), .ZN(n21677) );
  AOI21_X1 U31223 ( .B1(n4726), .B2(n24414), .A(n24117), .ZN(n21675) );
  OAI211_X1 U31224 ( .C1(n23731), .C2(n24409), .A(n21675), .B(n24119), .ZN(
        n21676) );
  XNOR2_X1 U31225 ( .A(n21680), .B(n25962), .ZN(n24531) );
  MUX2_X1 U31226 ( .A(n52175), .B(n51654), .S(n25056), .Z(n21682) );
  NAND2_X1 U31227 ( .A1(n21682), .A2(n22884), .ZN(n21685) );
  AND2_X1 U31228 ( .A1(n23101), .A2(n51654), .ZN(n22212) );
  NOR2_X1 U31229 ( .A1(n25056), .A2(n52175), .ZN(n21683) );
  AOI22_X1 U31230 ( .A1(n22874), .A2(n51654), .B1(n22212), .B2(n21683), .ZN(
        n21684) );
  NAND2_X1 U31231 ( .A1(n25064), .A2(n22876), .ZN(n25055) );
  MUX2_X1 U31232 ( .A(n21685), .B(n21684), .S(n25055), .Z(n21697) );
  INV_X1 U31234 ( .A(n22215), .ZN(n21691) );
  NAND2_X1 U31235 ( .A1(n25057), .A2(n25056), .ZN(n23095) );
  NOR2_X1 U31236 ( .A1(n23095), .A2(n22890), .ZN(n21690) );
  NAND2_X1 U31237 ( .A1(n51654), .A2(n52174), .ZN(n23093) );
  NAND3_X1 U31238 ( .A1(n25064), .A2(n23092), .A3(n23101), .ZN(n21687) );
  OAI211_X1 U31239 ( .C1(n23093), .C2(n22768), .A(n21688), .B(n21687), .ZN(
        n21689) );
  NAND3_X1 U31240 ( .A1(n23102), .A2(n7806), .A3(n23101), .ZN(n21693) );
  NAND2_X1 U31241 ( .A1(n23101), .A2(n52174), .ZN(n22765) );
  INV_X1 U31242 ( .A(n22765), .ZN(n22209) );
  NAND2_X1 U31243 ( .A1(n22207), .A2(n22209), .ZN(n21692) );
  MUX2_X1 U31244 ( .A(n21693), .B(n21692), .S(n25056), .Z(n21696) );
  INV_X1 U31245 ( .A(n23099), .ZN(n21694) );
  INV_X1 U31246 ( .A(n52175), .ZN(n22885) );
  NAND2_X1 U31247 ( .A1(n25056), .A2(n51654), .ZN(n22208) );
  OAI21_X1 U31248 ( .B1(n21694), .B2(n22885), .A(n22208), .ZN(n21695) );
  OAI21_X1 U31249 ( .B1(n21699), .B2(n21711), .A(n21716), .ZN(n21706) );
  NOR2_X1 U31250 ( .A1(n52048), .A2(n22184), .ZN(n21701) );
  AOI21_X1 U31251 ( .B1(n7119), .B2(n21701), .A(n21700), .ZN(n21705) );
  OAI21_X1 U31252 ( .B1(n463), .B2(n52048), .A(n21713), .ZN(n21704) );
  NOR2_X1 U31253 ( .A1(n21709), .A2(n21708), .ZN(n21720) );
  MUX2_X1 U31254 ( .A(n463), .B(n21715), .S(n21714), .Z(n21718) );
  NAND3_X1 U31255 ( .A1(n21718), .A2(n21717), .A3(n21716), .ZN(n21719) );
  NAND4_X2 U31256 ( .A1(n21721), .A2(n21720), .A3(n2270), .A4(n21719), .ZN(
        n28213) );
  INV_X1 U31257 ( .A(n24945), .ZN(n21764) );
  NAND3_X1 U31258 ( .A1(n23231), .A2(n22116), .A3(n23213), .ZN(n22401) );
  NAND2_X1 U31259 ( .A1(n21722), .A2(n22119), .ZN(n22402) );
  NAND2_X1 U31260 ( .A1(n22401), .A2(n22402), .ZN(n21724) );
  NAND2_X1 U31261 ( .A1(n6313), .A2(n413), .ZN(n23220) );
  NOR2_X1 U31262 ( .A1(n23213), .A2(n22116), .ZN(n22405) );
  NOR2_X1 U31263 ( .A1(n51355), .A2(n418), .ZN(n21728) );
  AND3_X1 U31264 ( .A1(n23230), .A2(n2102), .A3(n23207), .ZN(n21727) );
  AOI21_X1 U31265 ( .B1(n21734), .B2(n21737), .A(n21758), .ZN(n21735) );
  OAI21_X1 U31266 ( .B1(n21736), .B2(n21735), .A(n21756), .ZN(n21763) );
  NAND4_X1 U31267 ( .A1(n22262), .A2(n22256), .A3(n21755), .A4(n21737), .ZN(
        n21740) );
  NAND3_X1 U31269 ( .A1(n21755), .A2(n23341), .A3(n23336), .ZN(n21738) );
  OAI211_X1 U31270 ( .C1(n21740), .C2(n22257), .A(n21739), .B(n21738), .ZN(
        n21741) );
  INV_X1 U31271 ( .A(n21741), .ZN(n21762) );
  NAND2_X1 U31272 ( .A1(n21742), .A2(n629), .ZN(n21743) );
  AND2_X1 U31274 ( .A1(n21743), .A2(n23328), .ZN(n21761) );
  NAND2_X1 U31275 ( .A1(n21756), .A2(n21744), .ZN(n21754) );
  XNOR2_X1 U31276 ( .A(n23341), .B(n629), .ZN(n21753) );
  INV_X1 U31278 ( .A(n21748), .ZN(n21749) );
  NOR3_X1 U31279 ( .A1(n21751), .A2(n21750), .A3(n21749), .ZN(n21752) );
  AND3_X1 U31280 ( .A1(n21754), .A2(n21753), .A3(n21752), .ZN(n21759) );
  NOR2_X1 U31281 ( .A1(n21757), .A2(n21756), .ZN(n23345) );
  OAI21_X1 U31282 ( .B1(n21759), .B2(n23345), .A(n21758), .ZN(n21760) );
  NAND4_X2 U31283 ( .A1(n21762), .A2(n21760), .A3(n21763), .A4(n21761), .ZN(
        n27295) );
  XNOR2_X1 U31284 ( .A(n25003), .B(n27295), .ZN(n23745) );
  NAND2_X1 U31285 ( .A1(n22288), .A2(n22701), .ZN(n21766) );
  INV_X1 U31286 ( .A(n21769), .ZN(n21772) );
  NAND3_X1 U31287 ( .A1(n21772), .A2(n21771), .A3(n21770), .ZN(n21773) );
  OAI21_X1 U31288 ( .B1(n22291), .B2(n51695), .A(n22289), .ZN(n21776) );
  NAND2_X1 U31289 ( .A1(n21776), .A2(n21775), .ZN(n21788) );
  INV_X1 U31290 ( .A(n21777), .ZN(n21781) );
  NAND2_X1 U31291 ( .A1(n21778), .A2(n21781), .ZN(n22292) );
  AND2_X1 U31292 ( .A1(n22287), .A2(n21780), .ZN(n21783) );
  NAND2_X1 U31293 ( .A1(n23831), .A2(n24146), .ZN(n21791) );
  INV_X1 U31294 ( .A(n23834), .ZN(n23273) );
  OAI22_X1 U31295 ( .A1(n24161), .A2(n23832), .B1(n23273), .B2(n24159), .ZN(
        n21804) );
  INV_X1 U31296 ( .A(n24161), .ZN(n21792) );
  AND2_X1 U31297 ( .A1(n23832), .A2(n24158), .ZN(n23277) );
  NOR2_X1 U31298 ( .A1(n21792), .A2(n23277), .ZN(n21793) );
  AOI22_X1 U31299 ( .A1(n23835), .A2(n21793), .B1(n24148), .B2(n23268), .ZN(
        n21803) );
  MUX2_X1 U31300 ( .A(n24159), .B(n23824), .S(n24150), .Z(n21800) );
  NAND2_X1 U31301 ( .A1(n23833), .A2(n3520), .ZN(n21794) );
  NOR2_X1 U31302 ( .A1(n21794), .A2(n23832), .ZN(n21795) );
  NAND3_X1 U31304 ( .A1(n23826), .A2(n24158), .A3(n23833), .ZN(n21797) );
  NAND3_X1 U31305 ( .A1(n23827), .A2(n23833), .A3(n23832), .ZN(n21796) );
  NAND4_X1 U31306 ( .A1(n24149), .A2(n21798), .A3(n21797), .A4(n21796), .ZN(
        n21799) );
  AOI21_X1 U31307 ( .B1(n21801), .B2(n21800), .A(n21799), .ZN(n21802) );
  OAI211_X2 U31308 ( .C1(n21805), .C2(n21804), .A(n21803), .B(n21802), .ZN(
        n25508) );
  NOR2_X1 U31309 ( .A1(n24237), .A2(n24247), .ZN(n23451) );
  INV_X1 U31310 ( .A(n23451), .ZN(n23786) );
  NAND2_X1 U31311 ( .A1(n23786), .A2(n24250), .ZN(n23787) );
  NAND4_X1 U31312 ( .A1(n23787), .A2(n21810), .A3(n24245), .A4(n23785), .ZN(
        n21809) );
  NAND3_X1 U31313 ( .A1(n21806), .A2(n24238), .A3(n24245), .ZN(n21808) );
  NAND4_X1 U31314 ( .A1(n24242), .A2(n21823), .A3(n21811), .A4(n23785), .ZN(
        n21807) );
  AND3_X1 U31315 ( .A1(n21809), .A2(n21808), .A3(n21807), .ZN(n21827) );
  NAND2_X1 U31316 ( .A1(n21812), .A2(n21820), .ZN(n21816) );
  NAND2_X1 U31317 ( .A1(n21813), .A2(n24238), .ZN(n21814) );
  NAND2_X1 U31319 ( .A1(n21819), .A2(n21818), .ZN(n23782) );
  OAI211_X1 U31320 ( .C1(n24247), .C2(n21820), .A(n24239), .B(n23785), .ZN(
        n21821) );
  OR2_X1 U31321 ( .A1(n23782), .A2(n21821), .ZN(n21825) );
  NAND4_X1 U31322 ( .A1(n23782), .A2(n21823), .A3(n24238), .A4(n21822), .ZN(
        n21824) );
  XNOR2_X1 U31323 ( .A(n32520), .B(n4803), .ZN(n28211) );
  XNOR2_X1 U31324 ( .A(n28211), .B(n21828), .ZN(n44956) );
  XNOR2_X1 U31325 ( .A(n41426), .B(n4676), .ZN(n21829) );
  XNOR2_X1 U31326 ( .A(n44956), .B(n21829), .ZN(n21832) );
  INV_X1 U31327 ( .A(n21830), .ZN(n43267) );
  XNOR2_X1 U31328 ( .A(n43267), .B(n21831), .ZN(n42676) );
  XNOR2_X1 U31329 ( .A(n21832), .B(n42676), .ZN(n21833) );
  XNOR2_X1 U31330 ( .A(n25353), .B(n21833), .ZN(n21859) );
  NAND2_X1 U31331 ( .A1(n23257), .A2(n52133), .ZN(n21835) );
  INV_X1 U31332 ( .A(n21835), .ZN(n21834) );
  NAND2_X1 U31333 ( .A1(n23245), .A2(n757), .ZN(n21842) );
  OAI21_X1 U31334 ( .B1(n23245), .B2(n21835), .A(n21842), .ZN(n21839) );
  NAND3_X1 U31335 ( .A1(n21839), .A2(n21838), .A3(n21837), .ZN(n21840) );
  AND2_X1 U31336 ( .A1(n21841), .A2(n21840), .ZN(n21858) );
  NOR3_X1 U31337 ( .A1(n22658), .A2(n23257), .A3(n23254), .ZN(n21846) );
  INV_X1 U31338 ( .A(n21842), .ZN(n21845) );
  NAND2_X1 U31339 ( .A1(n23254), .A2(n52133), .ZN(n21843) );
  NOR2_X1 U31340 ( .A1(n23238), .A2(n21843), .ZN(n21844) );
  AOI21_X1 U31341 ( .B1(n21846), .B2(n21845), .A(n21844), .ZN(n21857) );
  OR2_X1 U31342 ( .A1(n23238), .A2(n23257), .ZN(n22134) );
  NOR2_X1 U31343 ( .A1(n22134), .A2(n22129), .ZN(n23253) );
  NAND2_X1 U31344 ( .A1(n22658), .A2(n23254), .ZN(n22133) );
  NAND2_X1 U31345 ( .A1(n22658), .A2(n757), .ZN(n22655) );
  INV_X1 U31346 ( .A(n22655), .ZN(n21850) );
  NAND2_X1 U31347 ( .A1(n23238), .A2(n23254), .ZN(n22649) );
  INV_X1 U31348 ( .A(n22649), .ZN(n21849) );
  NAND3_X1 U31349 ( .A1(n21850), .A2(n5294), .A3(n21849), .ZN(n21854) );
  NAND3_X1 U31350 ( .A1(n21852), .A2(n22129), .A3(n21851), .ZN(n21853) );
  AND2_X1 U31351 ( .A1(n21854), .A2(n21853), .ZN(n21855) );
  XNOR2_X1 U31352 ( .A(n21859), .B(n28214), .ZN(n21894) );
  OR2_X1 U31353 ( .A1(n22964), .A2(n23317), .ZN(n21866) );
  NAND2_X1 U31354 ( .A1(n23314), .A2(n23316), .ZN(n21860) );
  NOR2_X1 U31355 ( .A1(n756), .A2(n23306), .ZN(n21862) );
  INV_X1 U31356 ( .A(n21864), .ZN(n22962) );
  NAND3_X1 U31357 ( .A1(n21864), .A2(n23317), .A3(n23314), .ZN(n21865) );
  OAI21_X1 U31358 ( .B1(n22962), .B2(n21866), .A(n21865), .ZN(n21868) );
  OAI21_X1 U31360 ( .B1(n22254), .B2(n23316), .A(n22249), .ZN(n21869) );
  AND2_X1 U31361 ( .A1(n441), .A2(n23306), .ZN(n22955) );
  NAND2_X1 U31362 ( .A1(n21869), .A2(n22955), .ZN(n21870) );
  NAND2_X1 U31363 ( .A1(n23314), .A2(n21873), .ZN(n22959) );
  INV_X1 U31364 ( .A(n22959), .ZN(n21874) );
  NOR2_X1 U31365 ( .A1(n22849), .A2(n22856), .ZN(n21875) );
  NOR2_X1 U31366 ( .A1(n23021), .A2(n22864), .ZN(n22332) );
  INV_X1 U31367 ( .A(n22862), .ZN(n21876) );
  NAND4_X1 U31368 ( .A1(n22332), .A2(n22329), .A3(n21876), .A4(n22861), .ZN(
        n21878) );
  NOR2_X1 U31369 ( .A1(n21887), .A2(n22857), .ZN(n21888) );
  INV_X1 U31370 ( .A(n22865), .ZN(n21879) );
  NAND2_X1 U31371 ( .A1(n21880), .A2(n22849), .ZN(n21883) );
  NAND2_X1 U31372 ( .A1(n21880), .A2(n22859), .ZN(n21882) );
  AOI21_X1 U31373 ( .B1(n21885), .B2(n23020), .A(n22329), .ZN(n21881) );
  OAI211_X1 U31374 ( .C1(n21885), .C2(n23021), .A(n22851), .B(n22864), .ZN(
        n21892) );
  INV_X1 U31375 ( .A(n21886), .ZN(n21891) );
  NAND2_X1 U31376 ( .A1(n23020), .A2(n21887), .ZN(n22847) );
  INV_X1 U31377 ( .A(n21888), .ZN(n21889) );
  OAI211_X1 U31378 ( .C1(n22847), .C2(n23021), .A(n21889), .B(n22861), .ZN(
        n21890) );
  XNOR2_X1 U31379 ( .A(n26584), .B(n26160), .ZN(n25352) );
  XNOR2_X1 U31380 ( .A(n25352), .B(n21894), .ZN(n21997) );
  NAND2_X1 U31381 ( .A1(n23509), .A2(n23513), .ZN(n21896) );
  NOR2_X1 U31383 ( .A1(n24287), .A2(n24292), .ZN(n21899) );
  NAND3_X1 U31384 ( .A1(n24278), .A2(n7519), .A3(n24277), .ZN(n21901) );
  OAI211_X1 U31385 ( .C1(n21902), .C2(n23502), .A(n23508), .B(n21901), .ZN(
        n21903) );
  INV_X1 U31386 ( .A(n21903), .ZN(n21916) );
  NOR2_X1 U31387 ( .A1(n21905), .A2(n52206), .ZN(n21906) );
  NAND3_X1 U31388 ( .A1(n21908), .A2(n755), .A3(n21907), .ZN(n21910) );
  OAI211_X1 U31389 ( .C1(n24292), .C2(n21911), .A(n21910), .B(n21909), .ZN(
        n21912) );
  INV_X1 U31390 ( .A(n21912), .ZN(n21914) );
  OAI21_X1 U31391 ( .B1(n21921), .B2(n21937), .A(n21920), .ZN(n21924) );
  NAND2_X1 U31392 ( .A1(n22154), .A2(n22140), .ZN(n21922) );
  OAI22_X1 U31393 ( .A1(n21922), .A2(n22152), .B1(n22154), .B2(n2476), .ZN(
        n21923) );
  NOR2_X1 U31394 ( .A1(n21924), .A2(n21923), .ZN(n21943) );
  NAND4_X1 U31395 ( .A1(n22149), .A2(n22144), .A3(n21928), .A4(n22155), .ZN(
        n21930) );
  XNOR2_X1 U31396 ( .A(n50992), .B(n22140), .ZN(n21927) );
  NOR2_X1 U31397 ( .A1(n51661), .A2(n22155), .ZN(n21926) );
  NAND4_X1 U31398 ( .A1(n21928), .A2(n21927), .A3(n21926), .A4(n22144), .ZN(
        n21929) );
  AND2_X1 U31399 ( .A1(n21930), .A2(n21929), .ZN(n21942) );
  INV_X1 U31400 ( .A(n22149), .ZN(n21933) );
  INV_X1 U31401 ( .A(n21931), .ZN(n21932) );
  NAND4_X1 U31402 ( .A1(n21933), .A2(n22142), .A3(n22155), .A4(n21932), .ZN(
        n21936) );
  NAND2_X1 U31403 ( .A1(n21935), .A2(n21934), .ZN(n22161) );
  AND2_X1 U31404 ( .A1(n21936), .A2(n22161), .ZN(n21941) );
  NAND2_X1 U31405 ( .A1(n21938), .A2(n21937), .ZN(n21939) );
  NAND2_X1 U31406 ( .A1(n21939), .A2(n51661), .ZN(n21940) );
  INV_X1 U31407 ( .A(n24655), .ZN(n21944) );
  NAND2_X1 U31408 ( .A1(n21945), .A2(n51123), .ZN(n23152) );
  MUX2_X1 U31409 ( .A(n21946), .B(n23152), .S(n23473), .Z(n21967) );
  AND2_X1 U31410 ( .A1(n21947), .A2(n21957), .ZN(n21949) );
  OAI22_X1 U31411 ( .A1(n21949), .A2(n23467), .B1(n21948), .B2(n23157), .ZN(
        n21956) );
  NAND4_X1 U31413 ( .A1(n23465), .A2(n21953), .A3(n23153), .A4(n21957), .ZN(
        n21954) );
  NAND4_X1 U31414 ( .A1(n23473), .A2(n21957), .A3(n51123), .A4(n23157), .ZN(
        n21958) );
  NOR2_X1 U31415 ( .A1(n21960), .A2(n21959), .ZN(n21961) );
  NAND2_X1 U31416 ( .A1(n23147), .A2(n23467), .ZN(n21964) );
  MUX2_X1 U31417 ( .A(n21964), .B(n21963), .S(n23160), .Z(n21965) );
  INV_X1 U31418 ( .A(n21969), .ZN(n23484) );
  NAND2_X1 U31419 ( .A1(n23480), .A2(n2130), .ZN(n21979) );
  NAND2_X1 U31420 ( .A1(n21990), .A2(n23483), .ZN(n21972) );
  NAND3_X1 U31421 ( .A1(n21973), .A2(n21978), .A3(n21972), .ZN(n21995) );
  NAND2_X1 U31422 ( .A1(n21977), .A2(n21975), .ZN(n21976) );
  INV_X1 U31423 ( .A(n21979), .ZN(n21980) );
  NAND3_X1 U31424 ( .A1(n23485), .A2(n21981), .A3(n21980), .ZN(n21985) );
  INV_X1 U31425 ( .A(n23478), .ZN(n21982) );
  INV_X1 U31426 ( .A(n21983), .ZN(n21984) );
  INV_X1 U31427 ( .A(n21986), .ZN(n21989) );
  INV_X1 U31428 ( .A(n21987), .ZN(n21988) );
  NAND3_X1 U31429 ( .A1(n21992), .A2(n23485), .A3(n21991), .ZN(n21993) );
  XNOR2_X1 U31430 ( .A(n27289), .B(n24373), .ZN(n21996) );
  XNOR2_X1 U31431 ( .A(n21997), .B(n21996), .ZN(n21998) );
  NAND3_X1 U31432 ( .A1(n23446), .A2(n23436), .A3(n23442), .ZN(n22002) );
  INV_X1 U31433 ( .A(n21999), .ZN(n22000) );
  NAND2_X1 U31434 ( .A1(n22000), .A2(n22589), .ZN(n22001) );
  MUX2_X1 U31435 ( .A(n22002), .B(n22001), .S(n23441), .Z(n22030) );
  INV_X1 U31436 ( .A(n22003), .ZN(n22007) );
  INV_X1 U31437 ( .A(n22004), .ZN(n22005) );
  NOR2_X1 U31438 ( .A1(n22007), .A2(n22006), .ZN(n22029) );
  NOR2_X1 U31439 ( .A1(n22009), .A2(n23436), .ZN(n23444) );
  INV_X1 U31440 ( .A(n23444), .ZN(n22015) );
  NAND2_X1 U31441 ( .A1(n23438), .A2(n22010), .ZN(n22014) );
  OAI211_X1 U31442 ( .C1(n22016), .C2(n22015), .A(n22014), .B(n22013), .ZN(
        n22017) );
  INV_X1 U31443 ( .A(n22017), .ZN(n22028) );
  MUX2_X1 U31444 ( .A(n22019), .B(n22590), .S(n23446), .Z(n22026) );
  INV_X1 U31445 ( .A(n22020), .ZN(n22024) );
  OAI21_X1 U31446 ( .B1(n22024), .B2(n22023), .A(n22022), .ZN(n22025) );
  NAND4_X1 U31447 ( .A1(n22026), .A2(n23434), .A3(n22025), .A4(n23440), .ZN(
        n22027) );
  AND2_X1 U31448 ( .A1(n22035), .A2(n23411), .ZN(n22032) );
  AND2_X1 U31449 ( .A1(n23409), .A2(n23412), .ZN(n22031) );
  MUX2_X1 U31450 ( .A(n22032), .B(n22031), .S(n23417), .Z(n22043) );
  NAND3_X1 U31453 ( .A1(n22033), .A2(n452), .A3(n23426), .ZN(n22042) );
  OAI21_X1 U31454 ( .B1(n22034), .B2(n23421), .A(n23407), .ZN(n22041) );
  NAND3_X1 U31455 ( .A1(n23417), .A2(n22035), .A3(n22037), .ZN(n22039) );
  NAND3_X1 U31456 ( .A1(n23411), .A2(n22037), .A3(n22036), .ZN(n22038) );
  NAND3_X1 U31457 ( .A1(n22039), .A2(n23414), .A3(n22038), .ZN(n22040) );
  OAI211_X1 U31458 ( .C1(n22043), .C2(n22042), .A(n22041), .B(n22040), .ZN(
        n22054) );
  NOR2_X1 U31459 ( .A1(n23424), .A2(n23411), .ZN(n22044) );
  NOR2_X1 U31460 ( .A1(n22045), .A2(n22044), .ZN(n22053) );
  NOR2_X1 U31461 ( .A1(n23417), .A2(n22046), .ZN(n22047) );
  NOR2_X1 U31462 ( .A1(n24266), .A2(n22047), .ZN(n22052) );
  NAND2_X1 U31463 ( .A1(n22048), .A2(n22320), .ZN(n22049) );
  NAND4_X1 U31464 ( .A1(n22050), .A2(n22049), .A3(n23407), .A4(n23408), .ZN(
        n22051) );
  NAND2_X1 U31465 ( .A1(n7811), .A2(n23182), .ZN(n23179) );
  AND2_X1 U31466 ( .A1(n23179), .A2(n23171), .ZN(n22056) );
  NAND2_X1 U31467 ( .A1(n23175), .A2(n23182), .ZN(n22783) );
  OR2_X1 U31468 ( .A1(n22783), .A2(n3876), .ZN(n22677) );
  OAI211_X1 U31469 ( .C1(n22535), .C2(n22536), .A(n22056), .B(n22677), .ZN(
        n22060) );
  NOR2_X1 U31470 ( .A1(n23175), .A2(n23167), .ZN(n22057) );
  AOI21_X1 U31471 ( .B1(n23178), .B2(n22057), .A(n23171), .ZN(n23169) );
  OAI21_X1 U31472 ( .B1(n22793), .B2(n22058), .A(n23169), .ZN(n22059) );
  AND2_X1 U31473 ( .A1(n22061), .A2(n23167), .ZN(n22788) );
  INV_X1 U31474 ( .A(n22788), .ZN(n22062) );
  NAND2_X1 U31475 ( .A1(n22062), .A2(n23175), .ZN(n22063) );
  NOR2_X1 U31476 ( .A1(n22063), .A2(n23178), .ZN(n22065) );
  NOR2_X1 U31477 ( .A1(n22784), .A2(n5269), .ZN(n22064) );
  AOI22_X1 U31478 ( .A1(n22066), .A2(n22065), .B1(n22793), .B2(n22064), .ZN(
        n22069) );
  NOR2_X1 U31479 ( .A1(n51021), .A2(n23182), .ZN(n22668) );
  INV_X1 U31481 ( .A(n22090), .ZN(n22070) );
  INV_X1 U31482 ( .A(n23044), .ZN(n23053) );
  NAND2_X1 U31483 ( .A1(n23049), .A2(n23048), .ZN(n22751) );
  INV_X1 U31484 ( .A(n22751), .ZN(n22071) );
  AND2_X1 U31485 ( .A1(n23054), .A2(n23045), .ZN(n22934) );
  NAND2_X1 U31486 ( .A1(n22071), .A2(n22934), .ZN(n22078) );
  INV_X1 U31487 ( .A(n22072), .ZN(n22074) );
  NOR2_X1 U31488 ( .A1(n23048), .A2(n23054), .ZN(n23050) );
  INV_X1 U31489 ( .A(n23050), .ZN(n22073) );
  INV_X1 U31490 ( .A(n22944), .ZN(n22075) );
  NOR2_X1 U31491 ( .A1(n23045), .A2(n23044), .ZN(n22082) );
  INV_X1 U31492 ( .A(n22080), .ZN(n22081) );
  MUX2_X1 U31493 ( .A(n22082), .B(n22081), .S(n23049), .Z(n22084) );
  NAND2_X1 U31494 ( .A1(n23052), .A2(n22085), .ZN(n22936) );
  INV_X1 U31495 ( .A(n22936), .ZN(n22083) );
  NAND2_X1 U31496 ( .A1(n22084), .A2(n22083), .ZN(n22094) );
  AND2_X1 U31497 ( .A1(n22085), .A2(n424), .ZN(n22749) );
  NAND2_X1 U31498 ( .A1(n22943), .A2(n22749), .ZN(n22949) );
  NAND2_X1 U31499 ( .A1(n22086), .A2(n23045), .ZN(n23063) );
  NOR3_X1 U31500 ( .A1(n22087), .A2(n23052), .A3(n23048), .ZN(n22091) );
  INV_X1 U31501 ( .A(n22088), .ZN(n22752) );
  INV_X1 U31502 ( .A(n23060), .ZN(n22089) );
  INV_X1 U31503 ( .A(n24028), .ZN(n22096) );
  NAND2_X1 U31504 ( .A1(n24026), .A2(n22107), .ZN(n23668) );
  MUX2_X1 U31505 ( .A(n22096), .B(n23668), .S(n23392), .Z(n22113) );
  NAND2_X1 U31506 ( .A1(n22099), .A2(n22098), .ZN(n22106) );
  NAND4_X1 U31507 ( .A1(n22100), .A2(n24025), .A3(n24036), .A4(n24041), .ZN(
        n22104) );
  INV_X1 U31508 ( .A(n23674), .ZN(n22102) );
  NAND2_X1 U31509 ( .A1(n22575), .A2(n354), .ZN(n23394) );
  NOR2_X1 U31510 ( .A1(n23394), .A2(n24026), .ZN(n22109) );
  NOR2_X1 U31511 ( .A1(n24041), .A2(n22107), .ZN(n23395) );
  AOI22_X1 U31512 ( .A1(n24043), .A2(n22109), .B1(n22108), .B2(n23666), .ZN(
        n22111) );
  NOR2_X1 U31513 ( .A1(n24041), .A2(n354), .ZN(n24032) );
  NAND3_X1 U31514 ( .A1(n24032), .A2(n24033), .A3(n24030), .ZN(n23673) );
  XNOR2_X1 U31515 ( .A(n27258), .B(n22114), .ZN(n25864) );
  INV_X1 U31516 ( .A(n25864), .ZN(n24489) );
  NAND2_X1 U31517 ( .A1(n413), .A2(n22121), .ZN(n22122) );
  NOR2_X1 U31518 ( .A1(n22124), .A2(n22123), .ZN(n22652) );
  NOR2_X1 U31520 ( .A1(n22652), .A2(n22127), .ZN(n22139) );
  NAND2_X1 U31521 ( .A1(n22129), .A2(n757), .ZN(n23259) );
  NAND2_X1 U31522 ( .A1(n22129), .A2(n23245), .ZN(n23256) );
  NAND2_X1 U31523 ( .A1(n23259), .A2(n23256), .ZN(n22130) );
  NAND2_X1 U31524 ( .A1(n22130), .A2(n22650), .ZN(n22138) );
  MUX2_X1 U31525 ( .A(n23254), .B(n52134), .S(n23247), .Z(n22131) );
  NAND2_X1 U31526 ( .A1(n22132), .A2(n22131), .ZN(n22137) );
  INV_X1 U31527 ( .A(n22133), .ZN(n22135) );
  INV_X1 U31528 ( .A(n22134), .ZN(n23242) );
  NAND3_X1 U31529 ( .A1(n22142), .A2(n22141), .A3(n22140), .ZN(n22148) );
  OAI211_X1 U31530 ( .C1(n22146), .C2(n22143), .A(n22145), .B(n22144), .ZN(
        n22147) );
  OAI21_X1 U31531 ( .B1(n22149), .B2(n22148), .A(n22147), .ZN(n22150) );
  INV_X1 U31532 ( .A(n22150), .ZN(n22162) );
  OR2_X1 U31533 ( .A1(n22151), .A2(n51661), .ZN(n22153) );
  OAI211_X1 U31534 ( .C1(n22155), .C2(n22154), .A(n22153), .B(n22152), .ZN(
        n22160) );
  INV_X1 U31535 ( .A(n22156), .ZN(n22158) );
  NAND2_X1 U31536 ( .A1(n22158), .A2(n22157), .ZN(n22159) );
  OAI211_X1 U31538 ( .C1(n22914), .C2(n22916), .A(n22909), .B(n22169), .ZN(
        n22163) );
  NAND2_X1 U31539 ( .A1(n22163), .A2(n22165), .ZN(n22174) );
  NOR2_X1 U31540 ( .A1(n22164), .A2(n22348), .ZN(n22166) );
  AOI22_X1 U31541 ( .A1(n22913), .A2(n22166), .B1(n22165), .B2(n22168), .ZN(
        n22173) );
  NAND2_X1 U31542 ( .A1(n22168), .A2(n22167), .ZN(n22172) );
  NAND3_X1 U31543 ( .A1(n22170), .A2(n22902), .A3(n22169), .ZN(n22171) );
  XNOR2_X1 U31544 ( .A(n750), .B(n23879), .ZN(n25702) );
  INV_X1 U31545 ( .A(n25702), .ZN(n22234) );
  NAND2_X1 U31547 ( .A1(n22177), .A2(n22190), .ZN(n22195) );
  INV_X1 U31548 ( .A(n22183), .ZN(n22187) );
  NAND4_X1 U31549 ( .A1(n22187), .A2(n22186), .A3(n22185), .A4(n22184), .ZN(
        n22193) );
  AOI22_X1 U31550 ( .A1(n22191), .A2(n22190), .B1(n22189), .B2(n463), .ZN(
        n22192) );
  NOR2_X1 U31551 ( .A1(n23052), .A2(n23045), .ZN(n22941) );
  NAND3_X1 U31552 ( .A1(n22749), .A2(n22941), .A3(n23054), .ZN(n22196) );
  NAND2_X1 U31553 ( .A1(n23049), .A2(n23045), .ZN(n22200) );
  NAND3_X1 U31554 ( .A1(n22196), .A2(n22937), .A3(n22200), .ZN(n22198) );
  INV_X1 U31555 ( .A(n22197), .ZN(n23051) );
  NAND2_X1 U31556 ( .A1(n22198), .A2(n23051), .ZN(n22206) );
  NAND2_X1 U31557 ( .A1(n22199), .A2(n22753), .ZN(n22205) );
  AND2_X1 U31558 ( .A1(n23045), .A2(n23044), .ZN(n22930) );
  INV_X1 U31559 ( .A(n22930), .ZN(n22203) );
  AND2_X1 U31560 ( .A1(n23048), .A2(n22748), .ZN(n22931) );
  NAND2_X1 U31561 ( .A1(n22200), .A2(n22931), .ZN(n22202) );
  MUX2_X1 U31562 ( .A(n22203), .B(n22202), .S(n22201), .Z(n22204) );
  INV_X1 U31563 ( .A(n23098), .ZN(n22880) );
  INV_X1 U31564 ( .A(n22208), .ZN(n22210) );
  NAND2_X1 U31565 ( .A1(n23102), .A2(n22212), .ZN(n22213) );
  XNOR2_X1 U31566 ( .A(n22218), .B(n4782), .ZN(n42959) );
  XNOR2_X1 U31567 ( .A(n35838), .B(n4788), .ZN(n28233) );
  XNOR2_X1 U31568 ( .A(n28233), .B(n22219), .ZN(n40304) );
  XNOR2_X1 U31569 ( .A(n42959), .B(n40304), .ZN(n22220) );
  XNOR2_X1 U31570 ( .A(n25778), .B(n22220), .ZN(n22231) );
  NAND2_X1 U31571 ( .A1(n22492), .A2(n22823), .ZN(n22222) );
  NAND2_X1 U31572 ( .A1(n22826), .A2(n22506), .ZN(n22497) );
  INV_X1 U31573 ( .A(n22497), .ZN(n22221) );
  AOI22_X1 U31574 ( .A1(n22834), .A2(n22222), .B1(n22221), .B2(n22832), .ZN(
        n22228) );
  NAND2_X1 U31575 ( .A1(n22224), .A2(n22223), .ZN(n22227) );
  NAND3_X1 U31576 ( .A1(n22225), .A2(n8586), .A3(n22830), .ZN(n22226) );
  XNOR2_X1 U31577 ( .A(n24792), .B(n22231), .ZN(n22232) );
  XNOR2_X1 U31578 ( .A(n24171), .B(n22232), .ZN(n22233) );
  XNOR2_X1 U31579 ( .A(n22234), .B(n22233), .ZN(n22283) );
  NOR2_X1 U31580 ( .A1(n23706), .A2(n23535), .ZN(n23530) );
  NAND2_X1 U31581 ( .A1(n23530), .A2(n23531), .ZN(n22235) );
  INV_X1 U31582 ( .A(n23704), .ZN(n23528) );
  AND3_X1 U31583 ( .A1(n23528), .A2(n23703), .A3(n23694), .ZN(n22240) );
  NAND2_X1 U31584 ( .A1(n23637), .A2(n23090), .ZN(n23631) );
  INV_X1 U31585 ( .A(n23631), .ZN(n23964) );
  INV_X1 U31586 ( .A(n23953), .ZN(n22243) );
  NOR2_X1 U31587 ( .A1(n23641), .A2(n23961), .ZN(n22244) );
  NOR2_X1 U31588 ( .A1(n22244), .A2(n22623), .ZN(n22242) );
  NOR2_X1 U31589 ( .A1(n23955), .A2(n23958), .ZN(n22630) );
  NOR2_X1 U31590 ( .A1(n22623), .A2(n23961), .ZN(n23634) );
  AOI22_X1 U31591 ( .A1(n22242), .A2(n22630), .B1(n22241), .B2(n23634), .ZN(
        n22247) );
  OAI21_X1 U31592 ( .B1(n22244), .B2(n23963), .A(n22243), .ZN(n22246) );
  NAND4_X1 U31593 ( .A1(n23623), .A2(n23958), .A3(n23622), .A4(n23959), .ZN(
        n22245) );
  AOI21_X1 U31594 ( .B1(n8303), .B2(n23314), .A(n22964), .ZN(n22253) );
  NOR2_X1 U31596 ( .A1(n22256), .A2(n629), .ZN(n23330) );
  INV_X1 U31597 ( .A(n22257), .ZN(n22258) );
  NAND3_X1 U31598 ( .A1(n23330), .A2(n22262), .A3(n22258), .ZN(n22259) );
  NAND4_X1 U31599 ( .A1(n22264), .A2(n629), .A3(n22263), .A4(n22262), .ZN(
        n22265) );
  INV_X1 U31601 ( .A(n22635), .ZN(n22266) );
  NAND2_X1 U31602 ( .A1(n24206), .A2(n22266), .ZN(n23602) );
  INV_X1 U31603 ( .A(n24207), .ZN(n23606) );
  AND3_X1 U31604 ( .A1(n22641), .A2(n23606), .A3(n23066), .ZN(n22267) );
  NAND2_X1 U31605 ( .A1(n23597), .A2(n22268), .ZN(n22269) );
  OAI21_X1 U31606 ( .B1(n24206), .B2(n22269), .A(n23077), .ZN(n22270) );
  OAI21_X1 U31608 ( .B1(n22275), .B2(n23360), .A(n23570), .ZN(n22279) );
  XNOR2_X1 U31609 ( .A(n23360), .B(n23563), .ZN(n22277) );
  OAI211_X1 U31610 ( .C1(n23356), .C2(n51677), .A(n22279), .B(n22278), .ZN(
        n22280) );
  XNOR2_X1 U31611 ( .A(n22283), .B(n25289), .ZN(n22339) );
  OAI211_X1 U31612 ( .C1(n22288), .C2(n22287), .A(n22286), .B(n22285), .ZN(
        n22295) );
  NAND3_X1 U31613 ( .A1(n2084), .A2(n22698), .A3(n22702), .ZN(n22294) );
  NAND3_X1 U31614 ( .A1(n22291), .A2(n51694), .A3(n22290), .ZN(n22293) );
  NAND2_X1 U31615 ( .A1(n753), .A2(n51753), .ZN(n22301) );
  NAND3_X1 U31616 ( .A1(n22729), .A2(n22733), .A3(n22301), .ZN(n22296) );
  NAND2_X1 U31617 ( .A1(n22297), .A2(n22296), .ZN(n22305) );
  INV_X1 U31618 ( .A(n22298), .ZN(n22299) );
  OAI21_X1 U31619 ( .B1(n22373), .B2(n22299), .A(n5371), .ZN(n22300) );
  OAI211_X1 U31620 ( .C1(n5371), .C2(n51753), .A(n22300), .B(n22736), .ZN(
        n22304) );
  INV_X1 U31621 ( .A(n22395), .ZN(n22303) );
  NAND4_X1 U31622 ( .A1(n5371), .A2(n22741), .A3(n22375), .A4(n22301), .ZN(
        n22302) );
  XNOR2_X1 U31624 ( .A(n24757), .B(n25703), .ZN(n24793) );
  AND2_X1 U31625 ( .A1(n22306), .A2(n22481), .ZN(n22307) );
  AOI22_X1 U31626 ( .A1(n22717), .A2(n22307), .B1(n22462), .B2(n22714), .ZN(
        n22311) );
  INV_X1 U31627 ( .A(n22464), .ZN(n22718) );
  NOR2_X1 U31628 ( .A1(n23411), .A2(n23412), .ZN(n22312) );
  AOI22_X1 U31629 ( .A1(n22313), .A2(n22312), .B1(n23407), .B2(n23411), .ZN(
        n22324) );
  NAND2_X1 U31630 ( .A1(n23417), .A2(n23414), .ZN(n22323) );
  OAI21_X1 U31631 ( .B1(n23421), .B2(n22315), .A(n22314), .ZN(n22316) );
  NAND2_X1 U31632 ( .A1(n22316), .A2(n23423), .ZN(n22322) );
  NAND2_X1 U31633 ( .A1(n23417), .A2(n22317), .ZN(n22319) );
  OAI211_X1 U31634 ( .C1(n23422), .C2(n22320), .A(n22319), .B(n22318), .ZN(
        n22321) );
  XNOR2_X1 U31635 ( .A(n51720), .B(n4934), .ZN(n25881) );
  NAND2_X1 U31636 ( .A1(n22325), .A2(n23020), .ZN(n22326) );
  NAND3_X1 U31637 ( .A1(n22328), .A2(n22327), .A3(n22326), .ZN(n22337) );
  OAI21_X1 U31638 ( .B1(n22329), .B2(n23020), .A(n22861), .ZN(n22330) );
  INV_X1 U31639 ( .A(n22330), .ZN(n22331) );
  AOI22_X1 U31640 ( .A1(n22332), .A2(n22331), .B1(n22866), .B2(n22864), .ZN(
        n22336) );
  XNOR2_X1 U31641 ( .A(n25881), .B(n27473), .ZN(n22338) );
  XNOR2_X1 U31642 ( .A(n23793), .B(n22338), .ZN(n24392) );
  AND2_X1 U31643 ( .A1(n27632), .A2(n27732), .ZN(n27721) );
  OAI21_X1 U31644 ( .B1(n26806), .B2(n26888), .A(n27721), .ZN(n22343) );
  INV_X1 U31645 ( .A(n27633), .ZN(n22344) );
  INV_X1 U31646 ( .A(n27638), .ZN(n27635) );
  OAI22_X1 U31647 ( .A1(n22344), .A2(n24569), .B1(n27629), .B2(n27635), .ZN(
        n22340) );
  INV_X1 U31648 ( .A(n27632), .ZN(n24570) );
  INV_X1 U31649 ( .A(n22341), .ZN(n27621) );
  INV_X1 U31650 ( .A(n26888), .ZN(n27720) );
  OAI211_X1 U31651 ( .C1(n27621), .C2(n27720), .A(n27730), .B(n27627), .ZN(
        n22342) );
  NAND2_X1 U31652 ( .A1(n27627), .A2(n2144), .ZN(n22345) );
  OAI21_X1 U31653 ( .B1(n22346), .B2(n22345), .A(n27723), .ZN(n22347) );
  NAND2_X1 U31654 ( .A1(n22369), .A2(n22907), .ZN(n22353) );
  AND2_X1 U31655 ( .A1(n22348), .A2(n22367), .ZN(n22352) );
  NAND2_X1 U31656 ( .A1(n22908), .A2(n22349), .ZN(n22351) );
  NAND3_X1 U31657 ( .A1(n22354), .A2(n22908), .A3(n5542), .ZN(n22897) );
  NAND4_X1 U31658 ( .A1(n22357), .A2(n22356), .A3(n22355), .A4(n2175), .ZN(
        n22358) );
  NOR2_X1 U31659 ( .A1(n22901), .A2(n22367), .ZN(n22912) );
  INV_X1 U31660 ( .A(n22362), .ZN(n22364) );
  NAND2_X1 U31661 ( .A1(n5737), .A2(n22901), .ZN(n22920) );
  OAI21_X1 U31662 ( .B1(n22364), .B2(n22902), .A(n22899), .ZN(n22365) );
  AND2_X1 U31663 ( .A1(n22918), .A2(n22367), .ZN(n22903) );
  NAND3_X1 U31664 ( .A1(n22903), .A2(n22908), .A3(n22909), .ZN(n22371) );
  NAND2_X1 U31665 ( .A1(n22368), .A2(n22908), .ZN(n22370) );
  MUX2_X1 U31666 ( .A(n22371), .B(n22370), .S(n22369), .Z(n22372) );
  INV_X1 U31667 ( .A(n22373), .ZN(n22389) );
  NOR2_X1 U31668 ( .A1(n22374), .A2(n22389), .ZN(n22382) );
  NAND2_X1 U31669 ( .A1(n23811), .A2(n22375), .ZN(n22392) );
  OAI22_X1 U31670 ( .A1(n22392), .A2(n22733), .B1(n23811), .B2(n22375), .ZN(
        n22381) );
  INV_X1 U31671 ( .A(n22376), .ZN(n22378) );
  NAND2_X1 U31672 ( .A1(n22378), .A2(n22377), .ZN(n22380) );
  NAND2_X1 U31673 ( .A1(n22386), .A2(n22379), .ZN(n22737) );
  AOI22_X1 U31674 ( .A1(n22382), .A2(n22381), .B1(n22380), .B2(n22737), .ZN(
        n22399) );
  NAND2_X1 U31675 ( .A1(n22388), .A2(n22736), .ZN(n22383) );
  OR2_X1 U31676 ( .A1(n22384), .A2(n22383), .ZN(n22398) );
  INV_X1 U31677 ( .A(n22385), .ZN(n22387) );
  NAND2_X1 U31678 ( .A1(n22389), .A2(n23814), .ZN(n22393) );
  NAND3_X1 U31679 ( .A1(n22736), .A2(n22390), .A3(n51753), .ZN(n22391) );
  OAI21_X1 U31680 ( .B1(n22393), .B2(n22392), .A(n22391), .ZN(n22394) );
  NAND3_X2 U31681 ( .A1(n22397), .A2(n22398), .A3(n22399), .ZN(n23621) );
  INV_X1 U31682 ( .A(n23621), .ZN(n24660) );
  XNOR2_X1 U31683 ( .A(n27289), .B(n24660), .ZN(n25188) );
  XNOR2_X1 U31684 ( .A(n22400), .B(n25188), .ZN(n22415) );
  INV_X1 U31685 ( .A(n22405), .ZN(n22408) );
  NAND3_X1 U31686 ( .A1(n22406), .A2(n2102), .A3(n23207), .ZN(n22407) );
  OAI211_X1 U31687 ( .C1(n22408), .C2(n51355), .A(n23230), .B(n22407), .ZN(
        n22409) );
  XNOR2_X1 U31688 ( .A(n27250), .B(n24810), .ZN(n27440) );
  XNOR2_X1 U31689 ( .A(n24945), .B(n27440), .ZN(n23652) );
  XNOR2_X1 U31690 ( .A(n22415), .B(n23652), .ZN(n22517) );
  NOR2_X1 U31691 ( .A1(n23029), .A2(n23986), .ZN(n22417) );
  NAND2_X1 U31693 ( .A1(n23981), .A2(n23982), .ZN(n22533) );
  NOR3_X1 U31694 ( .A1(n23989), .A2(n23986), .A3(n22533), .ZN(n22419) );
  NAND2_X1 U31695 ( .A1(n24003), .A2(n23982), .ZN(n23031) );
  OAI21_X1 U31696 ( .B1(n23037), .B2(n22426), .A(n23031), .ZN(n22418) );
  NOR2_X1 U31697 ( .A1(n22419), .A2(n22418), .ZN(n22432) );
  AND2_X1 U31698 ( .A1(n22426), .A2(n23981), .ZN(n23999) );
  INV_X1 U31699 ( .A(n22420), .ZN(n22422) );
  NAND2_X1 U31700 ( .A1(n23982), .A2(n23992), .ZN(n22421) );
  NAND3_X1 U31701 ( .A1(n22422), .A2(n23986), .A3(n22421), .ZN(n22423) );
  AOI21_X1 U31702 ( .B1(n23983), .B2(n23999), .A(n22423), .ZN(n22425) );
  INV_X1 U31703 ( .A(n23032), .ZN(n22424) );
  INV_X1 U31704 ( .A(n22428), .ZN(n22429) );
  AND2_X1 U31705 ( .A1(n22532), .A2(n24006), .ZN(n22431) );
  AND2_X1 U31706 ( .A1(n22995), .A2(n22977), .ZN(n22556) );
  AOI22_X1 U31707 ( .A1(n22999), .A2(n22434), .B1(n22556), .B2(n22983), .ZN(
        n22439) );
  NAND3_X1 U31708 ( .A1(n22979), .A2(n22557), .A3(n22983), .ZN(n22435) );
  OAI211_X1 U31709 ( .C1(n22979), .C2(n22436), .A(n22435), .B(n23001), .ZN(
        n22437) );
  AND2_X1 U31710 ( .A1(n22439), .A2(n22438), .ZN(n22451) );
  NAND2_X1 U31711 ( .A1(n3691), .A2(n22978), .ZN(n22994) );
  NOR2_X1 U31712 ( .A1(n22994), .A2(n22990), .ZN(n22564) );
  NAND2_X1 U31713 ( .A1(n22564), .A2(n23001), .ZN(n22450) );
  INV_X1 U31714 ( .A(n22980), .ZN(n22440) );
  AOI21_X1 U31715 ( .B1(n22982), .B2(n22440), .A(n22978), .ZN(n22444) );
  OAI211_X1 U31716 ( .C1(n22557), .C2(n22989), .A(n22441), .B(n22979), .ZN(
        n22442) );
  INV_X1 U31717 ( .A(n22442), .ZN(n22443) );
  OR2_X1 U31718 ( .A1(n22978), .A2(n22989), .ZN(n23000) );
  INV_X1 U31719 ( .A(n23000), .ZN(n22563) );
  AOI22_X1 U31720 ( .A1(n22444), .A2(n22443), .B1(n22563), .B2(n22556), .ZN(
        n22449) );
  NAND4_X1 U31721 ( .A1(n22979), .A2(n22985), .A3(n22445), .A4(n22982), .ZN(
        n22446) );
  NAND2_X1 U31722 ( .A1(n22447), .A2(n22986), .ZN(n22448) );
  XNOR2_X1 U31723 ( .A(n25755), .B(n22452), .ZN(n27310) );
  XNOR2_X1 U31724 ( .A(n26436), .B(n27310), .ZN(n22515) );
  INV_X1 U31725 ( .A(n22453), .ZN(n34463) );
  XNOR2_X1 U31726 ( .A(n42712), .B(n34463), .ZN(n22456) );
  XNOR2_X1 U31727 ( .A(n35518), .B(n22454), .ZN(n42711) );
  XNOR2_X1 U31728 ( .A(n42711), .B(n24992), .ZN(n22455) );
  XNOR2_X1 U31729 ( .A(n22456), .B(n22455), .ZN(n22457) );
  XNOR2_X1 U31730 ( .A(n27303), .B(n22457), .ZN(n22489) );
  NAND2_X1 U31731 ( .A1(n22458), .A2(n22471), .ZN(n22460) );
  INV_X1 U31732 ( .A(n22722), .ZN(n22719) );
  INV_X1 U31733 ( .A(n22720), .ZN(n22459) );
  MUX2_X1 U31734 ( .A(n22460), .B(n22719), .S(n22459), .Z(n22487) );
  INV_X1 U31735 ( .A(n22461), .ZN(n22463) );
  NAND3_X1 U31736 ( .A1(n22463), .A2(n2083), .A3(n22462), .ZN(n22468) );
  NAND2_X1 U31737 ( .A1(n22464), .A2(n22481), .ZN(n22710) );
  INV_X1 U31738 ( .A(n22710), .ZN(n22465) );
  NAND2_X1 U31739 ( .A1(n22465), .A2(n2083), .ZN(n22467) );
  NAND4_X1 U31740 ( .A1(n22469), .A2(n22468), .A3(n22467), .A4(n22466), .ZN(
        n22475) );
  MUX2_X1 U31741 ( .A(n22714), .B(n2083), .S(n22488), .Z(n22473) );
  NAND3_X1 U31742 ( .A1(n22718), .A2(n22471), .A3(n22470), .ZN(n22472) );
  NOR2_X1 U31743 ( .A1(n22473), .A2(n22472), .ZN(n22474) );
  NOR2_X1 U31744 ( .A1(n22475), .A2(n22474), .ZN(n22486) );
  INV_X1 U31745 ( .A(n22478), .ZN(n22480) );
  OAI211_X1 U31746 ( .C1(n22482), .C2(n22481), .A(n22480), .B(n22479), .ZN(
        n22483) );
  NAND3_X1 U31747 ( .A1(n22484), .A2(n22488), .A3(n22483), .ZN(n22485) );
  OAI211_X1 U31748 ( .C1(n22488), .C2(n22487), .A(n22486), .B(n22485), .ZN(
        n23651) );
  XNOR2_X1 U31749 ( .A(n22489), .B(n25669), .ZN(n22513) );
  NAND2_X1 U31750 ( .A1(n22823), .A2(n22491), .ZN(n22493) );
  NAND4_X1 U31751 ( .A1(n22493), .A2(n22492), .A3(n22831), .A4(n22826), .ZN(
        n22495) );
  NAND2_X1 U31752 ( .A1(n22495), .A2(n22494), .ZN(n22501) );
  NAND2_X1 U31753 ( .A1(n22496), .A2(n22832), .ZN(n22500) );
  NAND3_X1 U31754 ( .A1(n22832), .A2(n22831), .A3(n22506), .ZN(n22498) );
  AOI21_X1 U31755 ( .B1(n22501), .B2(n22500), .A(n22499), .ZN(n22512) );
  NAND3_X1 U31756 ( .A1(n22832), .A2(n22509), .A3(n22826), .ZN(n22505) );
  OAI22_X1 U31757 ( .A1(n22830), .A2(n22509), .B1(n22826), .B2(n22506), .ZN(
        n22507) );
  OAI211_X1 U31758 ( .C1(n22832), .C2(n22509), .A(n22508), .B(n22507), .ZN(
        n22510) );
  XNOR2_X2 U31759 ( .A(n25353), .B(n25506), .ZN(n25762) );
  XNOR2_X1 U31761 ( .A(n22513), .B(n27256), .ZN(n22514) );
  XNOR2_X1 U31762 ( .A(n22515), .B(n22514), .ZN(n22516) );
  XNOR2_X1 U31763 ( .A(n22518), .B(n45083), .ZN(n42331) );
  XNOR2_X1 U31764 ( .A(n42331), .B(n45085), .ZN(n22519) );
  XNOR2_X1 U31765 ( .A(n26176), .B(n22519), .ZN(n22529) );
  NOR2_X1 U31766 ( .A1(n51034), .A2(n23906), .ZN(n22520) );
  AND2_X1 U31767 ( .A1(n22521), .A2(n23142), .ZN(n22803) );
  INV_X1 U31768 ( .A(n22803), .ZN(n23905) );
  NAND3_X1 U31769 ( .A1(n23921), .A2(n22524), .A3(n23905), .ZN(n22522) );
  NAND3_X1 U31771 ( .A1(n22523), .A2(n23913), .A3(n23904), .ZN(n22527) );
  AND2_X1 U31772 ( .A1(n51033), .A2(n23906), .ZN(n22804) );
  NAND2_X1 U31773 ( .A1(n22804), .A2(n23895), .ZN(n22526) );
  NOR2_X1 U31774 ( .A1(n6207), .A2(n51033), .ZN(n23897) );
  NAND3_X1 U31775 ( .A1(n23897), .A2(n23924), .A3(n22524), .ZN(n22525) );
  NAND4_X2 U31776 ( .A1(n22528), .A2(n22527), .A3(n22526), .A4(n22525), .ZN(
        n24795) );
  XNOR2_X1 U31777 ( .A(n22529), .B(n24795), .ZN(n22530) );
  XNOR2_X1 U31778 ( .A(n25609), .B(n22530), .ZN(n22570) );
  NOR2_X1 U31779 ( .A1(n23982), .A2(n23981), .ZN(n23033) );
  INV_X1 U31780 ( .A(n23172), .ZN(n22540) );
  NOR2_X1 U31781 ( .A1(n23178), .A2(n23166), .ZN(n22542) );
  NOR2_X1 U31782 ( .A1(n22542), .A2(n23183), .ZN(n22539) );
  INV_X1 U31783 ( .A(n22536), .ZN(n22537) );
  NAND2_X1 U31784 ( .A1(n22537), .A2(n23172), .ZN(n22538) );
  OAI211_X1 U31785 ( .C1(n22541), .C2(n22540), .A(n22539), .B(n22538), .ZN(
        n22553) );
  INV_X1 U31786 ( .A(n22543), .ZN(n22546) );
  INV_X1 U31787 ( .A(n22544), .ZN(n22545) );
  NAND3_X1 U31788 ( .A1(n22674), .A2(n22546), .A3(n22545), .ZN(n22547) );
  NAND2_X1 U31789 ( .A1(n22548), .A2(n22547), .ZN(n22672) );
  INV_X1 U31790 ( .A(n22783), .ZN(n22549) );
  NAND2_X1 U31791 ( .A1(n22672), .A2(n22549), .ZN(n22551) );
  NAND2_X1 U31792 ( .A1(n22789), .A2(n23182), .ZN(n22550) );
  NAND2_X1 U31793 ( .A1(n22556), .A2(n22989), .ZN(n22561) );
  INV_X1 U31794 ( .A(n22558), .ZN(n22559) );
  AND2_X1 U31795 ( .A1(n22560), .A2(n22561), .ZN(n22566) );
  NAND3_X1 U31796 ( .A1(n22563), .A2(n22982), .A3(n22562), .ZN(n22565) );
  XNOR2_X2 U31797 ( .A(n26264), .B(n25889), .ZN(n25608) );
  INV_X1 U31798 ( .A(n25608), .ZN(n22568) );
  XNOR2_X1 U31799 ( .A(n22569), .B(n22568), .ZN(n26032) );
  INV_X1 U31800 ( .A(n42686), .ZN(n45082) );
  XNOR2_X1 U31801 ( .A(n26610), .B(n45082), .ZN(n22571) );
  XNOR2_X1 U31802 ( .A(n23879), .B(n22571), .ZN(n22598) );
  MUX2_X1 U31803 ( .A(n22573), .B(n22572), .S(n24036), .Z(n22582) );
  NAND3_X1 U31806 ( .A1(n22576), .A2(n24042), .A3(n23392), .ZN(n22580) );
  OAI21_X1 U31807 ( .B1(n22578), .B2(n23395), .A(n22577), .ZN(n22579) );
  INV_X1 U31808 ( .A(n22583), .ZN(n22597) );
  NOR2_X1 U31809 ( .A1(n22585), .A2(n23446), .ZN(n22588) );
  AOI22_X1 U31810 ( .A1(n22588), .A2(n23441), .B1(n22587), .B2(n22586), .ZN(
        n22596) );
  INV_X1 U31811 ( .A(n22589), .ZN(n22592) );
  OAI21_X1 U31812 ( .B1(n22592), .B2(n22591), .A(n22590), .ZN(n22595) );
  NAND4_X1 U31813 ( .A1(n23438), .A2(n3513), .A3(n23433), .A4(n22593), .ZN(
        n22594) );
  XNOR2_X1 U31814 ( .A(n26600), .B(n25775), .ZN(n25700) );
  XNOR2_X1 U31815 ( .A(n22598), .B(n25700), .ZN(n25012) );
  XNOR2_X1 U31816 ( .A(n25738), .B(n25590), .ZN(n24545) );
  INV_X1 U31817 ( .A(n24189), .ZN(n23751) );
  NAND2_X1 U31818 ( .A1(n24187), .A2(n2210), .ZN(n23201) );
  NAND3_X1 U31819 ( .A1(n22601), .A2(n24188), .A3(n23201), .ZN(n22602) );
  NAND2_X1 U31820 ( .A1(n24190), .A2(n24186), .ZN(n23747) );
  NAND2_X1 U31821 ( .A1(n4328), .A2(n23756), .ZN(n22604) );
  AOI21_X1 U31822 ( .B1(n23747), .B2(n22604), .A(n23201), .ZN(n22608) );
  OR2_X1 U31823 ( .A1(n24190), .A2(n23756), .ZN(n23763) );
  NAND2_X1 U31824 ( .A1(n24177), .A2(n22606), .ZN(n22607) );
  NOR2_X1 U31825 ( .A1(n22608), .A2(n22607), .ZN(n22612) );
  AOI22_X1 U31826 ( .A1(n23750), .A2(n23871), .B1(n24179), .B2(n23764), .ZN(
        n22611) );
  NAND2_X1 U31827 ( .A1(n22609), .A2(n24187), .ZN(n22610) );
  XNOR2_X1 U31828 ( .A(n27382), .B(n47401), .ZN(n27446) );
  INV_X1 U31829 ( .A(n22614), .ZN(n22615) );
  XNOR2_X1 U31830 ( .A(n22615), .B(n23846), .ZN(n44292) );
  XNOR2_X1 U31831 ( .A(n22616), .B(n4076), .ZN(n46098) );
  XNOR2_X1 U31832 ( .A(n46098), .B(n4121), .ZN(n22617) );
  XNOR2_X1 U31833 ( .A(n44292), .B(n22617), .ZN(n22618) );
  XNOR2_X1 U31834 ( .A(n28311), .B(n22618), .ZN(n22619) );
  XNOR2_X1 U31835 ( .A(n27446), .B(n22619), .ZN(n22620) );
  XNOR2_X1 U31836 ( .A(n24545), .B(n22620), .ZN(n22665) );
  OR2_X1 U31837 ( .A1(n23963), .A2(n23959), .ZN(n22622) );
  NAND2_X1 U31838 ( .A1(n23959), .A2(n23090), .ZN(n22621) );
  MUX2_X1 U31839 ( .A(n22622), .B(n22621), .S(n23638), .Z(n22634) );
  OR2_X1 U31840 ( .A1(n22624), .A2(n23090), .ZN(n23645) );
  INV_X1 U31841 ( .A(n23645), .ZN(n23962) );
  NOR2_X1 U31842 ( .A1(n23638), .A2(n22625), .ZN(n22626) );
  AOI22_X1 U31843 ( .A1(n23962), .A2(n23635), .B1(n22626), .B2(n559), .ZN(
        n22633) );
  NOR2_X1 U31844 ( .A1(n23641), .A2(n559), .ZN(n22627) );
  OAI211_X1 U31845 ( .C1(n23953), .C2(n22627), .A(n23950), .B(n23961), .ZN(
        n22632) );
  OR2_X1 U31846 ( .A1(n5069), .A2(n23961), .ZN(n22629) );
  OAI211_X1 U31847 ( .C1(n22630), .C2(n22629), .A(n23964), .B(n22628), .ZN(
        n22631) );
  NAND2_X1 U31848 ( .A1(n23075), .A2(n22639), .ZN(n22637) );
  NAND2_X1 U31849 ( .A1(n22635), .A2(n23081), .ZN(n22636) );
  OAI211_X1 U31850 ( .C1(n22638), .C2(n22637), .A(n24206), .B(n22636), .ZN(
        n22648) );
  NOR2_X1 U31851 ( .A1(n23078), .A2(n22639), .ZN(n22640) );
  NAND2_X1 U31852 ( .A1(n52155), .A2(n17420), .ZN(n23076) );
  NAND2_X1 U31853 ( .A1(n22641), .A2(n24211), .ZN(n23611) );
  OAI21_X1 U31854 ( .B1(n22644), .B2(n22643), .A(n22642), .ZN(n22646) );
  NAND3_X1 U31855 ( .A1(n24208), .A2(n23080), .A3(n52155), .ZN(n22645) );
  NAND4_X2 U31856 ( .A1(n22648), .A2(n22647), .A3(n22646), .A4(n22645), .ZN(
        n26210) );
  XNOR2_X1 U31857 ( .A(n28424), .B(n27177), .ZN(n22663) );
  NOR2_X1 U31858 ( .A1(n23243), .A2(n23237), .ZN(n22651) );
  OAI22_X1 U31859 ( .A1(n22652), .A2(n22651), .B1(n22650), .B2(n22649), .ZN(
        n22662) );
  NAND2_X1 U31860 ( .A1(n22655), .A2(n23254), .ZN(n22657) );
  NAND2_X1 U31861 ( .A1(n23239), .A2(n23247), .ZN(n22656) );
  NAND3_X1 U31862 ( .A1(n22657), .A2(n23241), .A3(n22656), .ZN(n22661) );
  NAND3_X1 U31863 ( .A1(n22658), .A2(n52134), .A3(n23245), .ZN(n22659) );
  MUX2_X1 U31864 ( .A(n22659), .B(n23256), .S(n23247), .Z(n22660) );
  NAND4_X2 U31865 ( .A1(n22662), .A2(n8706), .A3(n22661), .A4(n22660), .ZN(
        n25920) );
  XNOR2_X1 U31866 ( .A(n22663), .B(n25920), .ZN(n22664) );
  XNOR2_X1 U31867 ( .A(n25638), .B(n22664), .ZN(n24087) );
  XNOR2_X1 U31868 ( .A(n24087), .B(n22665), .ZN(n22696) );
  NAND2_X1 U31869 ( .A1(n51021), .A2(n23167), .ZN(n22666) );
  MUX2_X1 U31870 ( .A(n22666), .B(n23183), .S(n23182), .Z(n22667) );
  NAND2_X1 U31871 ( .A1(n23178), .A2(n5269), .ZN(n22787) );
  OR2_X1 U31872 ( .A1(n22667), .A2(n22787), .ZN(n22680) );
  NOR2_X1 U31873 ( .A1(n22668), .A2(n5269), .ZN(n22671) );
  AND2_X1 U31874 ( .A1(n51021), .A2(n7811), .ZN(n23185) );
  NAND2_X1 U31875 ( .A1(n23170), .A2(n23183), .ZN(n22669) );
  NAND4_X1 U31876 ( .A1(n22672), .A2(n22671), .A3(n22670), .A4(n22669), .ZN(
        n22679) );
  AND2_X1 U31877 ( .A1(n23178), .A2(n23167), .ZN(n23164) );
  NAND3_X1 U31878 ( .A1(n23164), .A2(n3876), .A3(n22673), .ZN(n22678) );
  NAND3_X1 U31879 ( .A1(n23178), .A2(n23175), .A3(n23183), .ZN(n22676) );
  NAND3_X1 U31880 ( .A1(n23184), .A2(n22674), .A3(n23183), .ZN(n22675) );
  AOI21_X1 U31882 ( .B1(n23134), .B2(n23904), .A(n22683), .ZN(n22694) );
  NAND2_X1 U31883 ( .A1(n23142), .A2(n23895), .ZN(n22684) );
  OAI22_X1 U31884 ( .A1(n23141), .A2(n23143), .B1(n22796), .B2(n22684), .ZN(
        n22686) );
  NOR2_X1 U31885 ( .A1(n22686), .A2(n22685), .ZN(n22693) );
  OAI21_X1 U31886 ( .B1(n22688), .B2(n22804), .A(n22521), .ZN(n22689) );
  NAND3_X1 U31887 ( .A1(n22690), .A2(n22805), .A3(n22689), .ZN(n22692) );
  NOR2_X1 U31888 ( .A1(n23913), .A2(n23902), .ZN(n22795) );
  NAND2_X1 U31889 ( .A1(n23904), .A2(n22795), .ZN(n22691) );
  NAND2_X1 U31890 ( .A1(n22704), .A2(n22697), .ZN(n22707) );
  OAI21_X1 U31891 ( .B1(n51695), .B2(n22699), .A(n22698), .ZN(n22706) );
  AOI21_X1 U31892 ( .B1(n22703), .B2(n22702), .A(n22701), .ZN(n22705) );
  OAI21_X1 U31893 ( .B1(n22711), .B2(n22710), .A(n22709), .ZN(n22712) );
  INV_X1 U31894 ( .A(n22712), .ZN(n22726) );
  NAND3_X1 U31895 ( .A1(n22715), .A2(n22714), .A3(n22713), .ZN(n22725) );
  OAI211_X1 U31896 ( .C1(n22719), .C2(n22718), .A(n22717), .B(n22716), .ZN(
        n22724) );
  INV_X1 U31898 ( .A(n22728), .ZN(n22730) );
  AOI21_X1 U31899 ( .B1(n22733), .B2(n22732), .A(n22731), .ZN(n22734) );
  OAI211_X1 U31900 ( .C1(n5371), .C2(n22738), .A(n22737), .B(n51753), .ZN(
        n22745) );
  INV_X1 U31901 ( .A(n22739), .ZN(n22744) );
  NAND3_X1 U31902 ( .A1(n22742), .A2(n22741), .A3(n22740), .ZN(n22743) );
  XNOR2_X1 U31903 ( .A(n25821), .B(n28398), .ZN(n26055) );
  XNOR2_X1 U31904 ( .A(n26055), .B(n27346), .ZN(n26414) );
  INV_X1 U31905 ( .A(n22943), .ZN(n23061) );
  NAND2_X1 U31906 ( .A1(n22930), .A2(n22748), .ZN(n22750) );
  OAI211_X1 U31907 ( .C1(n23061), .C2(n22934), .A(n22750), .B(n22749), .ZN(
        n22760) );
  INV_X1 U31908 ( .A(n22932), .ZN(n22759) );
  NAND2_X1 U31909 ( .A1(n22752), .A2(n22751), .ZN(n22758) );
  NAND2_X1 U31910 ( .A1(n23052), .A2(n23044), .ZN(n22754) );
  INV_X1 U31911 ( .A(n22937), .ZN(n22755) );
  NAND2_X1 U31912 ( .A1(n22756), .A2(n22755), .ZN(n22757) );
  XNOR2_X2 U31913 ( .A(n25161), .B(n26402), .ZN(n28121) );
  XNOR2_X1 U31914 ( .A(n28121), .B(n24344), .ZN(n22761) );
  XNOR2_X1 U31915 ( .A(n26414), .B(n22761), .ZN(n27195) );
  XNOR2_X1 U31916 ( .A(n27502), .B(n4618), .ZN(n26518) );
  AOI22_X1 U31917 ( .A1(n23097), .A2(n23095), .B1(n22767), .B2(n22766), .ZN(
        n22773) );
  AND2_X1 U31918 ( .A1(n52175), .A2(n7806), .ZN(n22889) );
  NAND3_X1 U31919 ( .A1(n22889), .A2(n23092), .A3(n23101), .ZN(n22770) );
  XNOR2_X1 U31920 ( .A(n26518), .B(n25542), .ZN(n22782) );
  XNOR2_X1 U31921 ( .A(n32856), .B(n46552), .ZN(n43848) );
  XOR2_X1 U31922 ( .A(n4627), .B(n4874), .Z(n22774) );
  XNOR2_X1 U31923 ( .A(n43848), .B(n22774), .ZN(n22775) );
  XNOR2_X1 U31924 ( .A(n22776), .B(n22775), .ZN(n45055) );
  XNOR2_X1 U31925 ( .A(n24315), .B(n22777), .ZN(n42355) );
  XNOR2_X1 U31926 ( .A(n42355), .B(n45051), .ZN(n22778) );
  XNOR2_X1 U31927 ( .A(n45055), .B(n22778), .ZN(n22779) );
  XNOR2_X1 U31928 ( .A(n28396), .B(n22779), .ZN(n22780) );
  XNOR2_X1 U31929 ( .A(n28287), .B(n25548), .ZN(n26116) );
  XNOR2_X1 U31930 ( .A(n22780), .B(n26116), .ZN(n22781) );
  XNOR2_X1 U31931 ( .A(n22782), .B(n22781), .ZN(n22812) );
  AND2_X1 U31932 ( .A1(n22784), .A2(n22783), .ZN(n22794) );
  AND2_X1 U31933 ( .A1(n22785), .A2(n23183), .ZN(n22786) );
  OAI22_X1 U31934 ( .A1(n22787), .A2(n22786), .B1(n23166), .B2(n23183), .ZN(
        n22791) );
  NAND2_X1 U31935 ( .A1(n22789), .A2(n22788), .ZN(n22790) );
  INV_X1 U31936 ( .A(n22795), .ZN(n22798) );
  INV_X1 U31937 ( .A(n22796), .ZN(n23914) );
  INV_X1 U31940 ( .A(n23923), .ZN(n23896) );
  OAI21_X1 U31941 ( .B1(n23926), .B2(n23896), .A(n23904), .ZN(n22808) );
  INV_X1 U31942 ( .A(n22801), .ZN(n22802) );
  NAND3_X1 U31943 ( .A1(n23898), .A2(n23926), .A3(n22802), .ZN(n22807) );
  OAI21_X1 U31944 ( .B1(n22805), .B2(n22804), .A(n22803), .ZN(n22806) );
  XNOR2_X1 U31945 ( .A(n22810), .B(n25829), .ZN(n22811) );
  XNOR2_X1 U31946 ( .A(n22812), .B(n22811), .ZN(n22813) );
  INV_X1 U31947 ( .A(n34255), .ZN(n22815) );
  XNOR2_X1 U31948 ( .A(n22815), .B(n22814), .ZN(n43204) );
  XNOR2_X1 U31949 ( .A(n45107), .B(n22816), .ZN(n42082) );
  XNOR2_X1 U31950 ( .A(n42101), .B(n4868), .ZN(n22817) );
  XNOR2_X1 U31951 ( .A(n42082), .B(n22817), .ZN(n22818) );
  XNOR2_X1 U31952 ( .A(n43204), .B(n22818), .ZN(n22819) );
  XNOR2_X1 U31953 ( .A(n27419), .B(n22819), .ZN(n22842) );
  NAND2_X1 U31954 ( .A1(n22821), .A2(n22830), .ZN(n22841) );
  NAND2_X1 U31955 ( .A1(n22832), .A2(n22823), .ZN(n22825) );
  NAND3_X1 U31956 ( .A1(n22832), .A2(n22831), .A3(n22830), .ZN(n22833) );
  OAI21_X1 U31957 ( .B1(n22835), .B2(n22834), .A(n22833), .ZN(n22836) );
  XNOR2_X1 U31958 ( .A(n22842), .B(n25947), .ZN(n22843) );
  XNOR2_X1 U31959 ( .A(n52184), .B(n22843), .ZN(n22873) );
  INV_X1 U31960 ( .A(n22844), .ZN(n22848) );
  NAND2_X1 U31961 ( .A1(n23021), .A2(n22864), .ZN(n22845) );
  OAI22_X1 U31962 ( .A1(n22848), .A2(n22847), .B1(n22846), .B2(n22845), .ZN(
        n22853) );
  NAND2_X1 U31963 ( .A1(n22849), .A2(n22864), .ZN(n22850) );
  NOR2_X1 U31964 ( .A1(n22851), .A2(n22850), .ZN(n22852) );
  NOR2_X1 U31965 ( .A1(n22853), .A2(n22852), .ZN(n22872) );
  NAND2_X1 U31967 ( .A1(n22858), .A2(n22857), .ZN(n22863) );
  NAND2_X1 U31968 ( .A1(n22859), .A2(n4413), .ZN(n22860) );
  NAND4_X1 U31969 ( .A1(n22863), .A2(n22862), .A3(n22861), .A4(n22860), .ZN(
        n22870) );
  NOR2_X1 U31970 ( .A1(n22865), .A2(n22864), .ZN(n22867) );
  OAI21_X1 U31971 ( .B1(n22868), .B2(n22867), .A(n22866), .ZN(n22869) );
  XNOR2_X1 U31972 ( .A(n27218), .B(n22873), .ZN(n22929) );
  NAND3_X1 U31974 ( .A1(n25064), .A2(n22876), .A3(n7806), .ZN(n22877) );
  AND2_X1 U31975 ( .A1(n22878), .A2(n22877), .ZN(n22895) );
  NOR2_X1 U31976 ( .A1(n25064), .A2(n23101), .ZN(n22879) );
  NAND2_X1 U31977 ( .A1(n22880), .A2(n23093), .ZN(n22881) );
  NAND4_X1 U31978 ( .A1(n22882), .A2(n22881), .A3(n23100), .A4(n23105), .ZN(
        n22894) );
  NAND2_X1 U31979 ( .A1(n51654), .A2(n23092), .ZN(n22883) );
  XNOR2_X1 U31980 ( .A(n22883), .B(n25064), .ZN(n22888) );
  INV_X1 U31981 ( .A(n22883), .ZN(n22886) );
  AOI21_X1 U31982 ( .B1(n22886), .B2(n22885), .A(n22884), .ZN(n22887) );
  NAND2_X1 U31983 ( .A1(n22888), .A2(n22887), .ZN(n22893) );
  XNOR2_X1 U31984 ( .A(n25064), .B(n25056), .ZN(n22891) );
  OAI21_X1 U31985 ( .B1(n22891), .B2(n22890), .A(n22889), .ZN(n22892) );
  INV_X1 U31987 ( .A(n22900), .ZN(n22925) );
  NAND4_X1 U31988 ( .A1(n22903), .A2(n22902), .A3(n2175), .A4(n22901), .ZN(
        n22906) );
  AND2_X1 U31990 ( .A1(n22906), .A2(n22905), .ZN(n22924) );
  AND2_X1 U31991 ( .A1(n22908), .A2(n22907), .ZN(n22911) );
  INV_X1 U31992 ( .A(n22909), .ZN(n22910) );
  INV_X1 U31993 ( .A(n22914), .ZN(n22922) );
  NAND2_X1 U31994 ( .A1(n22916), .A2(n2175), .ZN(n22917) );
  OAI211_X1 U31995 ( .C1(n22920), .C2(n5542), .A(n22918), .B(n22917), .ZN(
        n22921) );
  NAND2_X1 U31996 ( .A1(n22922), .A2(n22921), .ZN(n22923) );
  XNOR2_X1 U31997 ( .A(n28381), .B(n44044), .ZN(n22926) );
  XNOR2_X1 U31998 ( .A(n27420), .B(n22927), .ZN(n26137) );
  INV_X1 U31999 ( .A(n26137), .ZN(n22928) );
  XNOR2_X1 U32000 ( .A(n22929), .B(n22928), .ZN(n22975) );
  XNOR2_X1 U32001 ( .A(n25240), .B(n51665), .ZN(n22953) );
  OAI22_X1 U32002 ( .A1(n22937), .A2(n22936), .B1(n22935), .B2(n22934), .ZN(
        n22938) );
  NOR2_X1 U32003 ( .A1(n22939), .A2(n22938), .ZN(n22951) );
  NOR2_X1 U32004 ( .A1(n23048), .A2(n23053), .ZN(n22942) );
  NOR2_X1 U32005 ( .A1(n23048), .A2(n23044), .ZN(n22940) );
  AOI22_X1 U32006 ( .A1(n22943), .A2(n22942), .B1(n22941), .B2(n22940), .ZN(
        n22950) );
  AOI21_X1 U32007 ( .B1(n22944), .B2(n23045), .A(n23054), .ZN(n22945) );
  OAI21_X1 U32008 ( .B1(n22947), .B2(n424), .A(n22945), .ZN(n22948) );
  NAND4_X2 U32009 ( .A1(n22951), .A2(n22949), .A3(n22948), .A4(n22950), .ZN(
        n28049) );
  XNOR2_X1 U32010 ( .A(n28049), .B(n4157), .ZN(n22952) );
  XNOR2_X1 U32011 ( .A(n22953), .B(n22952), .ZN(n27418) );
  OAI21_X1 U32013 ( .B1(n22957), .B2(n22956), .A(n23303), .ZN(n22972) );
  AOI22_X1 U32014 ( .A1(n22960), .A2(n22959), .B1(n22958), .B2(n441), .ZN(
        n22971) );
  NAND3_X1 U32015 ( .A1(n22962), .A2(n22961), .A3(n942), .ZN(n22965) );
  OAI21_X1 U32016 ( .B1(n23316), .B2(n23314), .A(n23312), .ZN(n22963) );
  NAND3_X1 U32017 ( .A1(n23314), .A2(n23316), .A3(n8303), .ZN(n22967) );
  NAND2_X1 U32018 ( .A1(n23311), .A2(n22967), .ZN(n22968) );
  XNOR2_X1 U32019 ( .A(n27418), .B(n27217), .ZN(n22974) );
  XNOR2_X1 U32020 ( .A(n22975), .B(n22974), .ZN(n23109) );
  XNOR2_X1 U32021 ( .A(n28274), .B(n3383), .ZN(n22976) );
  XNOR2_X1 U32022 ( .A(n22976), .B(n26540), .ZN(n24438) );
  AOI21_X1 U32023 ( .B1(n22981), .B2(n22989), .A(n22980), .ZN(n22988) );
  AND2_X1 U32024 ( .A1(n22982), .A2(n22983), .ZN(n22984) );
  OAI21_X1 U32025 ( .B1(n22986), .B2(n22985), .A(n22984), .ZN(n22987) );
  OAI211_X1 U32026 ( .C1(n22990), .C2(n22989), .A(n22988), .B(n22987), .ZN(
        n22991) );
  NOR2_X1 U32027 ( .A1(n23001), .A2(n22995), .ZN(n22996) );
  NAND3_X1 U32028 ( .A1(n23000), .A2(n22999), .A3(n22998), .ZN(n23004) );
  OR2_X1 U32029 ( .A1(n23002), .A2(n23001), .ZN(n23003) );
  XNOR2_X1 U32030 ( .A(n2082), .B(n25124), .ZN(n25574) );
  INV_X1 U32031 ( .A(n25574), .ZN(n23005) );
  XNOR2_X1 U32032 ( .A(n24438), .B(n23005), .ZN(n23018) );
  XNOR2_X1 U32033 ( .A(n27483), .B(n41567), .ZN(n44332) );
  XNOR2_X1 U32034 ( .A(n46065), .B(n44332), .ZN(n23006) );
  XNOR2_X1 U32035 ( .A(n26147), .B(n23006), .ZN(n23014) );
  INV_X1 U32036 ( .A(n4847), .ZN(n50586) );
  AND2_X1 U32037 ( .A1(n23332), .A2(n4847), .ZN(n23009) );
  NAND4_X1 U32038 ( .A1(n23010), .A2(n23009), .A3(n23013), .A4(n23008), .ZN(
        n23011) );
  XNOR2_X1 U32039 ( .A(n23014), .B(n26548), .ZN(n23016) );
  INV_X1 U32040 ( .A(n25457), .ZN(n23206) );
  XNOR2_X1 U32041 ( .A(n23016), .B(n23015), .ZN(n23017) );
  INV_X1 U32042 ( .A(n23019), .ZN(n23026) );
  AOI21_X1 U32043 ( .B1(n2352), .B2(n23021), .A(n23020), .ZN(n23022) );
  OAI21_X1 U32044 ( .B1(n23026), .B2(n23025), .A(n23024), .ZN(n23042) );
  INV_X1 U32045 ( .A(n23033), .ZN(n23034) );
  NAND2_X1 U32046 ( .A1(n23034), .A2(n23992), .ZN(n23035) );
  OAI21_X1 U32047 ( .B1(n23037), .B2(n24000), .A(n24001), .ZN(n23040) );
  NAND4_X1 U32048 ( .A1(n23984), .A2(n23983), .A3(n24002), .A4(n23981), .ZN(
        n23038) );
  NAND3_X1 U32049 ( .A1(n23038), .A2(n23986), .A3(n23996), .ZN(n23039) );
  XNOR2_X1 U32050 ( .A(n25308), .B(n46062), .ZN(n23043) );
  NAND2_X1 U32051 ( .A1(n22201), .A2(n23044), .ZN(n23047) );
  NOR2_X1 U32052 ( .A1(n23047), .A2(n23045), .ZN(n23046) );
  OAI21_X1 U32053 ( .B1(n2381), .B2(n23046), .A(n23049), .ZN(n23065) );
  INV_X1 U32054 ( .A(n23047), .ZN(n23059) );
  AOI21_X1 U32055 ( .B1(n23051), .B2(n23050), .A(n23049), .ZN(n23057) );
  NAND3_X1 U32056 ( .A1(n23055), .A2(n23054), .A3(n23053), .ZN(n23056) );
  OAI211_X1 U32057 ( .C1(n23059), .C2(n23058), .A(n23057), .B(n23056), .ZN(
        n23064) );
  OR2_X1 U32058 ( .A1(n23061), .A2(n23060), .ZN(n23062) );
  NAND2_X1 U32059 ( .A1(n52155), .A2(n23613), .ZN(n23067) );
  NAND3_X1 U32060 ( .A1(n23067), .A2(n23066), .A3(n17420), .ZN(n23070) );
  NOR2_X1 U32061 ( .A1(n23590), .A2(n23068), .ZN(n23610) );
  NAND2_X1 U32062 ( .A1(n24205), .A2(n23610), .ZN(n23069) );
  OAI211_X1 U32063 ( .C1(n23595), .C2(n23070), .A(n23592), .B(n23069), .ZN(
        n23071) );
  INV_X1 U32064 ( .A(n23071), .ZN(n23085) );
  INV_X1 U32065 ( .A(n24206), .ZN(n23074) );
  NAND4_X1 U32066 ( .A1(n23074), .A2(n23073), .A3(n23075), .A4(n23072), .ZN(
        n23084) );
  NOR2_X1 U32067 ( .A1(n24211), .A2(n23075), .ZN(n23607) );
  NAND3_X1 U32068 ( .A1(n23077), .A2(n23607), .A3(n23076), .ZN(n23083) );
  INV_X1 U32069 ( .A(n23078), .ZN(n23079) );
  OAI21_X1 U32070 ( .B1(n23081), .B2(n23080), .A(n23079), .ZN(n23082) );
  NAND4_X2 U32071 ( .A1(n23085), .A2(n23084), .A3(n23083), .A4(n23082), .ZN(
        n27374) );
  AOI21_X1 U32072 ( .B1(n23955), .B2(n23090), .A(n23950), .ZN(n23086) );
  NAND2_X1 U32073 ( .A1(n23087), .A2(n23955), .ZN(n23088) );
  OR2_X1 U32074 ( .A1(n23090), .A2(n23957), .ZN(n23625) );
  INV_X1 U32075 ( .A(n25726), .ZN(n25790) );
  OR2_X1 U32076 ( .A1(n23093), .A2(n23092), .ZN(n23294) );
  NAND3_X1 U32079 ( .A1(n23295), .A2(n25064), .A3(n23294), .ZN(n25053) );
  OAI21_X1 U32080 ( .B1(n23102), .B2(n25064), .A(n23101), .ZN(n23103) );
  INV_X1 U32081 ( .A(n24904), .ZN(n23107) );
  XNOR2_X1 U32082 ( .A(n28410), .B(n24691), .ZN(n25999) );
  XNOR2_X1 U32083 ( .A(n25999), .B(n25790), .ZN(n25965) );
  NAND2_X1 U32084 ( .A1(n2109), .A2(n28809), .ZN(n30722) );
  INV_X1 U32085 ( .A(n28809), .ZN(n27162) );
  OAI22_X1 U32086 ( .A1(n4020), .A2(n30722), .B1(n30709), .B2(n28810), .ZN(
        n23111) );
  NAND2_X1 U32087 ( .A1(n2169), .A2(n2205), .ZN(n28808) );
  NAND3_X1 U32088 ( .A1(n27588), .A2(n28810), .A3(n27162), .ZN(n23110) );
  OAI21_X1 U32089 ( .B1(n30716), .B2(n30711), .A(n28810), .ZN(n23113) );
  NAND2_X1 U32090 ( .A1(n30724), .A2(n23113), .ZN(n23114) );
  NAND3_X1 U32091 ( .A1(n30716), .A2(n27162), .A3(n29853), .ZN(n27592) );
  MUX2_X1 U32092 ( .A(n23114), .B(n27592), .S(n2205), .Z(n23115) );
  NAND2_X1 U32093 ( .A1(n32254), .A2(n31778), .ZN(n32236) );
  INV_X1 U32094 ( .A(n51751), .ZN(n25553) );
  XNOR2_X1 U32095 ( .A(n25346), .B(n25553), .ZN(n26362) );
  XNOR2_X1 U32096 ( .A(n26362), .B(n51120), .ZN(n23121) );
  XNOR2_X1 U32097 ( .A(n33050), .B(n45883), .ZN(n43151) );
  XNOR2_X1 U32098 ( .A(n36823), .B(n36737), .ZN(n23116) );
  XNOR2_X1 U32099 ( .A(n43151), .B(n23116), .ZN(n23117) );
  XNOR2_X1 U32100 ( .A(n41831), .B(n23117), .ZN(n23118) );
  XNOR2_X1 U32101 ( .A(n26573), .B(n23118), .ZN(n23119) );
  XNOR2_X1 U32102 ( .A(n51119), .B(n23119), .ZN(n23120) );
  INV_X1 U32103 ( .A(n24855), .ZN(n24405) );
  XNOR2_X1 U32104 ( .A(n24405), .B(n24705), .ZN(n23123) );
  XNOR2_X1 U32105 ( .A(n2106), .B(n51667), .ZN(n24218) );
  XNOR2_X1 U32106 ( .A(n25935), .B(n24218), .ZN(n23188) );
  NOR2_X1 U32107 ( .A1(n24413), .A2(n24117), .ZN(n24100) );
  NOR2_X1 U32108 ( .A1(n24100), .A2(n23124), .ZN(n23125) );
  MUX2_X1 U32109 ( .A(n23125), .B(n24412), .S(n24106), .Z(n23131) );
  OAI211_X1 U32110 ( .C1(n24113), .C2(n24411), .A(n24412), .B(n24071), .ZN(
        n24408) );
  OAI21_X1 U32111 ( .B1(n24105), .B2(n24409), .A(n24413), .ZN(n23126) );
  AND2_X1 U32112 ( .A1(n51001), .A2(n23129), .ZN(n24065) );
  NAND2_X1 U32113 ( .A1(n23126), .A2(n24065), .ZN(n24419) );
  OR2_X1 U32114 ( .A1(n24070), .A2(n24116), .ZN(n24407) );
  INV_X1 U32115 ( .A(n23127), .ZN(n24101) );
  INV_X1 U32116 ( .A(n24413), .ZN(n24112) );
  NAND3_X1 U32117 ( .A1(n24101), .A2(n24112), .A3(n24111), .ZN(n23128) );
  AND4_X1 U32118 ( .A1(n24408), .A2(n24419), .A3(n24407), .A4(n23128), .ZN(
        n23130) );
  OAI211_X1 U32119 ( .C1(n24111), .C2(n23131), .A(n23130), .B(n24420), .ZN(
        n23146) );
  AOI21_X1 U32120 ( .B1(n23911), .B2(n6207), .A(n23926), .ZN(n23133) );
  AOI21_X1 U32121 ( .B1(n23926), .B2(n23913), .A(n23906), .ZN(n23132) );
  OAI22_X1 U32122 ( .A1(n23133), .A2(n23135), .B1(n23132), .B2(n23924), .ZN(
        n23140) );
  NAND2_X1 U32123 ( .A1(n51034), .A2(n23142), .ZN(n23909) );
  OAI21_X1 U32124 ( .B1(n23908), .B2(n23909), .A(n23925), .ZN(n23139) );
  NOR2_X1 U32125 ( .A1(n23135), .A2(n51034), .ZN(n23919) );
  NAND2_X1 U32126 ( .A1(n23921), .A2(n23919), .ZN(n23137) );
  AND2_X1 U32127 ( .A1(n23137), .A2(n23136), .ZN(n23138) );
  AND2_X1 U32128 ( .A1(n23902), .A2(n23924), .ZN(n23907) );
  OAI211_X1 U32129 ( .C1(n23907), .C2(n23913), .A(n23143), .B(n23142), .ZN(
        n23145) );
  NAND3_X1 U32130 ( .A1(n23923), .A2(n23143), .A3(n23906), .ZN(n23144) );
  XNOR2_X1 U32131 ( .A(n23146), .B(n27211), .ZN(n23187) );
  INV_X1 U32132 ( .A(n23147), .ZN(n23148) );
  OAI21_X1 U32133 ( .B1(n23150), .B2(n51123), .A(n23148), .ZN(n23151) );
  AOI21_X1 U32134 ( .B1(n23154), .B2(n23467), .A(n23153), .ZN(n23155) );
  OAI211_X1 U32135 ( .C1(n23472), .C2(n23160), .A(n23159), .B(n23158), .ZN(
        n23162) );
  NAND2_X1 U32136 ( .A1(n23471), .A2(n23467), .ZN(n23161) );
  INV_X1 U32137 ( .A(n23164), .ZN(n23165) );
  INV_X1 U32139 ( .A(n23170), .ZN(n23173) );
  OAI21_X1 U32140 ( .B1(n23173), .B2(n23172), .A(n23171), .ZN(n23174) );
  NAND3_X1 U32141 ( .A1(n23176), .A2(n23178), .A3(n23175), .ZN(n23181) );
  NAND3_X1 U32142 ( .A1(n23179), .A2(n23178), .A3(n51021), .ZN(n23180) );
  NAND4_X1 U32143 ( .A1(n23185), .A2(n23184), .A3(n23183), .A4(n23182), .ZN(
        n23186) );
  INV_X1 U32144 ( .A(n26287), .ZN(n26569) );
  XNOR2_X1 U32145 ( .A(n23188), .B(n26569), .ZN(n23189) );
  OAI21_X1 U32146 ( .B1(n23191), .B2(n23756), .A(n24187), .ZN(n23192) );
  NAND2_X1 U32147 ( .A1(n23193), .A2(n23192), .ZN(n23199) );
  INV_X1 U32148 ( .A(n24182), .ZN(n23195) );
  NAND2_X1 U32149 ( .A1(n23196), .A2(n23195), .ZN(n23197) );
  NOR2_X1 U32150 ( .A1(n23200), .A2(n24187), .ZN(n23767) );
  INV_X1 U32151 ( .A(n23747), .ZN(n23766) );
  OAI21_X1 U32152 ( .B1(n23203), .B2(n23756), .A(n23201), .ZN(n23202) );
  NAND2_X1 U32153 ( .A1(n23202), .A2(n24188), .ZN(n23205) );
  NOR2_X1 U32154 ( .A1(n23203), .A2(n2210), .ZN(n23864) );
  AND2_X1 U32155 ( .A1(n24190), .A2(n24180), .ZN(n23865) );
  NAND2_X1 U32156 ( .A1(n23864), .A2(n23865), .ZN(n23204) );
  XNOR2_X1 U32157 ( .A(n26304), .B(n23206), .ZN(n27363) );
  NOR2_X1 U32158 ( .A1(n23230), .A2(n23207), .ZN(n23210) );
  AOI22_X1 U32159 ( .A1(n23211), .A2(n23210), .B1(n23209), .B2(n413), .ZN(
        n23216) );
  OAI21_X1 U32160 ( .B1(n23213), .B2(n23219), .A(n23212), .ZN(n23214) );
  NAND2_X1 U32161 ( .A1(n23214), .A2(n51355), .ZN(n23215) );
  AND3_X1 U32162 ( .A1(n23216), .A2(n23217), .A3(n23215), .ZN(n23236) );
  NAND3_X1 U32163 ( .A1(n23220), .A2(n23219), .A3(n23218), .ZN(n23222) );
  NAND2_X1 U32164 ( .A1(n23222), .A2(n51355), .ZN(n23228) );
  INV_X1 U32165 ( .A(n23223), .ZN(n23226) );
  OAI21_X1 U32166 ( .B1(n23226), .B2(n23225), .A(n18369), .ZN(n23227) );
  NAND2_X1 U32167 ( .A1(n23228), .A2(n23227), .ZN(n23234) );
  NOR2_X1 U32168 ( .A1(n23230), .A2(n2102), .ZN(n23232) );
  INV_X1 U32169 ( .A(n23237), .ZN(n23240) );
  OAI21_X1 U32170 ( .B1(n23240), .B2(n23239), .A(n23238), .ZN(n23252) );
  NAND2_X1 U32171 ( .A1(n23243), .A2(n23242), .ZN(n23250) );
  OAI211_X1 U32172 ( .C1(n23246), .C2(n23254), .A(n23245), .B(n52134), .ZN(
        n23248) );
  NAND2_X1 U32173 ( .A1(n23248), .A2(n5292), .ZN(n23249) );
  NAND4_X1 U32174 ( .A1(n23252), .A2(n23251), .A3(n23250), .A4(n23249), .ZN(
        n23265) );
  OAI21_X1 U32175 ( .B1(n23255), .B2(n23254), .A(n23253), .ZN(n23264) );
  INV_X1 U32176 ( .A(n23256), .ZN(n23258) );
  NAND2_X1 U32177 ( .A1(n23258), .A2(n23257), .ZN(n23263) );
  INV_X1 U32178 ( .A(n23259), .ZN(n23260) );
  NAND2_X1 U32179 ( .A1(n23261), .A2(n23260), .ZN(n23262) );
  XNOR2_X1 U32180 ( .A(n27363), .B(n26556), .ZN(n23285) );
  INV_X1 U32181 ( .A(n4639), .ZN(n23266) );
  XNOR2_X1 U32182 ( .A(n26152), .B(n23266), .ZN(n23283) );
  NAND3_X1 U32183 ( .A1(n24150), .A2(n24158), .A3(n23828), .ZN(n23270) );
  NAND3_X1 U32184 ( .A1(n23268), .A2(n24150), .A3(n23828), .ZN(n23269) );
  INV_X1 U32185 ( .A(n23272), .ZN(n23282) );
  OAI211_X1 U32186 ( .C1(n23824), .C2(n24157), .A(n23832), .B(n23825), .ZN(
        n23275) );
  INV_X1 U32187 ( .A(n23824), .ZN(n24147) );
  NAND4_X1 U32188 ( .A1(n24147), .A2(n23833), .A3(n23832), .A4(n23273), .ZN(
        n23274) );
  NAND2_X1 U32189 ( .A1(n23278), .A2(n23277), .ZN(n23280) );
  NAND2_X1 U32190 ( .A1(n23835), .A2(n24145), .ZN(n23279) );
  XNOR2_X1 U32191 ( .A(n51647), .B(n23283), .ZN(n25252) );
  INV_X1 U32192 ( .A(n25252), .ZN(n23284) );
  XNOR2_X1 U32193 ( .A(n23285), .B(n23284), .ZN(n23287) );
  XNOR2_X1 U32194 ( .A(n23287), .B(n23286), .ZN(n23300) );
  XNOR2_X1 U32195 ( .A(n24047), .B(n4931), .ZN(n27368) );
  XNOR2_X1 U32196 ( .A(n24430), .B(n4536), .ZN(n43528) );
  XNOR2_X1 U32197 ( .A(n34057), .B(n43528), .ZN(n23288) );
  XNOR2_X1 U32198 ( .A(n28274), .B(n23288), .ZN(n23289) );
  XNOR2_X1 U32199 ( .A(n27368), .B(n23289), .ZN(n23293) );
  INV_X1 U32200 ( .A(n23290), .ZN(n23292) );
  XNOR2_X1 U32201 ( .A(n25124), .B(n27232), .ZN(n23291) );
  XNOR2_X1 U32202 ( .A(n24578), .B(n23293), .ZN(n23298) );
  INV_X1 U32203 ( .A(n23294), .ZN(n25058) );
  NAND2_X1 U32204 ( .A1(n25058), .A2(n25056), .ZN(n25054) );
  AND2_X1 U32205 ( .A1(n23295), .A2(n23294), .ZN(n25065) );
  INV_X1 U32206 ( .A(n25065), .ZN(n23296) );
  MUX2_X1 U32207 ( .A(n25054), .B(n23296), .S(n25064), .Z(n23297) );
  NAND3_X1 U32208 ( .A1(n23297), .A2(n25052), .A3(n25061), .ZN(n24526) );
  XNOR2_X1 U32209 ( .A(n28276), .B(n24526), .ZN(n24235) );
  XNOR2_X1 U32210 ( .A(n23298), .B(n24235), .ZN(n23299) );
  XNOR2_X1 U32211 ( .A(n23300), .B(n23299), .ZN(n27566) );
  NAND2_X1 U32212 ( .A1(n23301), .A2(n27566), .ZN(n29907) );
  XNOR2_X1 U32213 ( .A(n751), .B(n43560), .ZN(n23302) );
  XNOR2_X1 U32214 ( .A(n25088), .B(n23302), .ZN(n24306) );
  AND2_X1 U32215 ( .A1(n441), .A2(n23303), .ZN(n23305) );
  NAND2_X1 U32216 ( .A1(n23305), .A2(n756), .ZN(n23309) );
  MUX2_X1 U32217 ( .A(n23309), .B(n23319), .S(n23317), .Z(n23327) );
  NAND3_X1 U32218 ( .A1(n23305), .A2(n23310), .A3(n23316), .ZN(n23308) );
  MUX2_X1 U32219 ( .A(n23308), .B(n23307), .S(n23306), .Z(n23326) );
  INV_X1 U32220 ( .A(n23309), .ZN(n23315) );
  NOR2_X1 U32221 ( .A1(n23311), .A2(n23310), .ZN(n23313) );
  AOI22_X1 U32222 ( .A1(n23315), .A2(n23314), .B1(n23313), .B2(n23312), .ZN(
        n23325) );
  OAI21_X1 U32223 ( .B1(n23318), .B2(n942), .A(n23316), .ZN(n23323) );
  NAND3_X1 U32224 ( .A1(n23323), .A2(n23322), .A3(n23321), .ZN(n23324) );
  NAND2_X1 U32226 ( .A1(n23345), .A2(n23330), .ZN(n23331) );
  AND2_X1 U32227 ( .A1(n23332), .A2(n23331), .ZN(n23348) );
  OAI22_X1 U32228 ( .A1(n23335), .A2(n23334), .B1(n23342), .B2(n23333), .ZN(
        n23340) );
  NAND2_X1 U32229 ( .A1(n1024), .A2(n23336), .ZN(n23337) );
  AOI21_X1 U32230 ( .B1(n23342), .B2(n23338), .A(n23337), .ZN(n23339) );
  NOR2_X1 U32231 ( .A1(n23340), .A2(n23339), .ZN(n23347) );
  INV_X1 U32232 ( .A(n23343), .ZN(n23344) );
  NOR2_X1 U32233 ( .A1(n23350), .A2(n51676), .ZN(n23354) );
  OAI21_X1 U32234 ( .B1(n22274), .B2(n23352), .A(n23351), .ZN(n23353) );
  OAI21_X1 U32235 ( .B1(n23355), .B2(n23354), .A(n23353), .ZN(n23368) );
  OR2_X1 U32236 ( .A1(n23356), .A2(n23360), .ZN(n23359) );
  NOR2_X1 U32237 ( .A1(n23554), .A2(n23570), .ZN(n23358) );
  AOI21_X1 U32238 ( .B1(n23359), .B2(n23358), .A(n23357), .ZN(n23367) );
  OR2_X1 U32239 ( .A1(n23361), .A2(n23360), .ZN(n23557) );
  OAI21_X1 U32240 ( .B1(n23557), .B2(n23363), .A(n23362), .ZN(n23366) );
  OAI21_X1 U32241 ( .B1(n23559), .B2(n23364), .A(n23363), .ZN(n23365) );
  NAND4_X1 U32242 ( .A1(n23368), .A2(n23367), .A3(n23366), .A4(n23365), .ZN(
        n25589) );
  XNOR2_X1 U32243 ( .A(n24306), .B(n23369), .ZN(n23391) );
  XNOR2_X1 U32244 ( .A(n23370), .B(n25426), .ZN(n23371) );
  XNOR2_X1 U32245 ( .A(n33346), .B(n23371), .ZN(n44221) );
  XNOR2_X1 U32246 ( .A(n43552), .B(n44221), .ZN(n23372) );
  XNOR2_X1 U32247 ( .A(n26100), .B(n23372), .ZN(n23385) );
  OAI211_X1 U32249 ( .C1(n24332), .C2(n23702), .A(n24336), .B(n5415), .ZN(
        n23373) );
  AND2_X1 U32250 ( .A1(n50990), .A2(n457), .ZN(n23692) );
  OAI21_X1 U32251 ( .B1(n24326), .B2(n24324), .A(n23692), .ZN(n23377) );
  OAI21_X1 U32252 ( .B1(n23375), .B2(n50990), .A(n23695), .ZN(n23376) );
  NAND2_X1 U32253 ( .A1(n23377), .A2(n23376), .ZN(n23382) );
  NAND2_X1 U32254 ( .A1(n23530), .A2(n24332), .ZN(n23380) );
  NOR2_X1 U32255 ( .A1(n23382), .A2(n23381), .ZN(n23383) );
  XNOR2_X1 U32257 ( .A(n23385), .B(n369), .ZN(n23387) );
  XNOR2_X1 U32258 ( .A(n26044), .B(n26509), .ZN(n23386) );
  XNOR2_X1 U32259 ( .A(n23386), .B(n26395), .ZN(n24083) );
  XNOR2_X1 U32260 ( .A(n23387), .B(n24083), .ZN(n23389) );
  XNOR2_X1 U32261 ( .A(n23388), .B(n27452), .ZN(n28318) );
  XNOR2_X1 U32262 ( .A(n28318), .B(n23389), .ZN(n23390) );
  XNOR2_X1 U32263 ( .A(n26125), .B(n25548), .ZN(n23971) );
  XNOR2_X1 U32264 ( .A(n28295), .B(n23971), .ZN(n23406) );
  XNOR2_X1 U32265 ( .A(n24556), .B(n1354), .ZN(n26229) );
  OAI21_X1 U32266 ( .B1(n23666), .B2(n23674), .A(n23395), .ZN(n23396) );
  XNOR2_X1 U32267 ( .A(n25825), .B(n4826), .ZN(n27355) );
  XNOR2_X1 U32268 ( .A(n26229), .B(n27355), .ZN(n23404) );
  INV_X1 U32269 ( .A(n23397), .ZN(n23398) );
  XNOR2_X1 U32270 ( .A(n23399), .B(n23398), .ZN(n42647) );
  XNOR2_X1 U32271 ( .A(n4884), .B(n4837), .ZN(n46122) );
  XNOR2_X1 U32272 ( .A(n43848), .B(n46122), .ZN(n23400) );
  XNOR2_X1 U32273 ( .A(n42647), .B(n23400), .ZN(n23401) );
  XNOR2_X1 U32274 ( .A(n23404), .B(n23403), .ZN(n23405) );
  XNOR2_X1 U32275 ( .A(n23406), .B(n23405), .ZN(n23462) );
  XNOR2_X1 U32276 ( .A(n28398), .B(n28121), .ZN(n27509) );
  NOR2_X1 U32277 ( .A1(n23408), .A2(n23407), .ZN(n23419) );
  NAND3_X1 U32278 ( .A1(n23410), .A2(n452), .A3(n23409), .ZN(n23416) );
  NAND4_X1 U32279 ( .A1(n23414), .A2(n452), .A3(n23412), .A4(n23411), .ZN(
        n23415) );
  OAI21_X1 U32280 ( .B1(n23417), .B2(n23416), .A(n23415), .ZN(n23418) );
  AOI21_X1 U32281 ( .B1(n23420), .B2(n23419), .A(n23418), .ZN(n23432) );
  NOR2_X1 U32282 ( .A1(n23426), .A2(n23425), .ZN(n23427) );
  INV_X1 U32283 ( .A(n23428), .ZN(n23429) );
  NAND2_X1 U32284 ( .A1(n23437), .A2(n23436), .ZN(n23439) );
  NAND2_X1 U32285 ( .A1(n23439), .A2(n23438), .ZN(n23450) );
  OAI22_X1 U32286 ( .A1(n23441), .A2(n23446), .B1(n23440), .B2(n23445), .ZN(
        n23443) );
  NAND2_X1 U32287 ( .A1(n23443), .A2(n23442), .ZN(n23449) );
  OAI21_X1 U32288 ( .B1(n23446), .B2(n23445), .A(n23444), .ZN(n23448) );
  AND2_X1 U32289 ( .A1(n23451), .A2(n23785), .ZN(n24249) );
  OAI21_X1 U32290 ( .B1(n6744), .B2(n24246), .A(n24242), .ZN(n23459) );
  NAND3_X1 U32291 ( .A1(n24244), .A2(n24248), .A3(n24247), .ZN(n23453) );
  AND2_X1 U32292 ( .A1(n23452), .A2(n23453), .ZN(n23458) );
  OAI21_X1 U32293 ( .B1(n23456), .B2(n23455), .A(n23454), .ZN(n23457) );
  INV_X1 U32294 ( .A(n26531), .ZN(n23460) );
  XNOR2_X1 U32295 ( .A(n23460), .B(n26119), .ZN(n24873) );
  XNOR2_X1 U32296 ( .A(n24873), .B(n52201), .ZN(n25450) );
  INV_X1 U32297 ( .A(n25450), .ZN(n24980) );
  XNOR2_X1 U32298 ( .A(n27509), .B(n24980), .ZN(n23461) );
  XNOR2_X1 U32299 ( .A(n24171), .B(n24936), .ZN(n28231) );
  INV_X1 U32300 ( .A(n23472), .ZN(n23474) );
  NAND3_X1 U32301 ( .A1(n23474), .A2(n2076), .A3(n23473), .ZN(n23475) );
  NAND3_X1 U32302 ( .A1(n23490), .A2(n23489), .A3(n23488), .ZN(n23491) );
  XNOR2_X1 U32303 ( .A(n51750), .B(n23879), .ZN(n27469) );
  XNOR2_X1 U32304 ( .A(n28231), .B(n27469), .ZN(n23501) );
  XNOR2_X1 U32305 ( .A(n27322), .B(n51720), .ZN(n23498) );
  XNOR2_X1 U32306 ( .A(n4788), .B(n4721), .ZN(n23492) );
  XNOR2_X1 U32307 ( .A(n45463), .B(n23492), .ZN(n23493) );
  XNOR2_X1 U32308 ( .A(n23494), .B(n23493), .ZN(n44977) );
  XNOR2_X1 U32309 ( .A(n36945), .B(n23495), .ZN(n42689) );
  XNOR2_X1 U32310 ( .A(n44977), .B(n42689), .ZN(n23496) );
  XNOR2_X1 U32311 ( .A(n51648), .B(n23496), .ZN(n23497) );
  XNOR2_X1 U32312 ( .A(n23498), .B(n23497), .ZN(n23499) );
  XNOR2_X1 U32313 ( .A(n26264), .B(n51749), .ZN(n23801) );
  XNOR2_X1 U32314 ( .A(n23801), .B(n27473), .ZN(n24170) );
  XNOR2_X1 U32315 ( .A(n23499), .B(n24170), .ZN(n23500) );
  NOR2_X1 U32316 ( .A1(n23503), .A2(n23502), .ZN(n23505) );
  MUX2_X1 U32317 ( .A(n23506), .B(n23505), .S(n23504), .Z(n23517) );
  NAND2_X1 U32318 ( .A1(n24285), .A2(n23508), .ZN(n24284) );
  NOR2_X1 U32319 ( .A1(n24290), .A2(n23510), .ZN(n24288) );
  INV_X1 U32320 ( .A(n23511), .ZN(n23512) );
  NAND3_X1 U32321 ( .A1(n24288), .A2(n23513), .A3(n23512), .ZN(n23514) );
  XNOR2_X1 U32322 ( .A(n27479), .B(n25613), .ZN(n23523) );
  AND2_X1 U32323 ( .A1(n24105), .A2(n24117), .ZN(n24102) );
  INV_X1 U32324 ( .A(n24102), .ZN(n23520) );
  NAND2_X1 U32325 ( .A1(n24065), .A2(n24105), .ZN(n24068) );
  NAND3_X1 U32326 ( .A1(n24113), .A2(n23730), .A3(n24111), .ZN(n23522) );
  XNOR2_X1 U32327 ( .A(n24616), .B(n28352), .ZN(n24390) );
  XNOR2_X1 U32328 ( .A(n24390), .B(n24795), .ZN(n27325) );
  XNOR2_X1 U32329 ( .A(n26584), .B(n23525), .ZN(n23527) );
  INV_X1 U32330 ( .A(n26160), .ZN(n23526) );
  XNOR2_X1 U32331 ( .A(n23527), .B(n23526), .ZN(n23580) );
  MUX2_X1 U32332 ( .A(n23528), .B(n3816), .S(n5415), .Z(n23529) );
  NOR2_X1 U32333 ( .A1(n457), .A2(n50990), .ZN(n23539) );
  INV_X1 U32335 ( .A(n24330), .ZN(n23700) );
  INV_X1 U32336 ( .A(n23530), .ZN(n23533) );
  OR2_X1 U32340 ( .A1(n23538), .A2(n24329), .ZN(n23542) );
  INV_X1 U32341 ( .A(n23539), .ZN(n23541) );
  NAND4_X1 U32342 ( .A1(n23542), .A2(n23704), .A3(n23541), .A4(n23540), .ZN(
        n23543) );
  OAI21_X1 U32343 ( .B1(n51677), .B2(n23568), .A(n23546), .ZN(n23548) );
  AND2_X1 U32344 ( .A1(n23548), .A2(n23547), .ZN(n23550) );
  INV_X1 U32345 ( .A(n23552), .ZN(n23556) );
  NAND2_X1 U32347 ( .A1(n23558), .A2(n23557), .ZN(n23577) );
  INV_X1 U32348 ( .A(n23559), .ZN(n23560) );
  NAND2_X1 U32349 ( .A1(n23561), .A2(n51676), .ZN(n23576) );
  OAI21_X1 U32350 ( .B1(n51676), .B2(n23563), .A(n8205), .ZN(n23565) );
  NOR2_X1 U32351 ( .A1(n17074), .A2(n23568), .ZN(n23572) );
  INV_X1 U32352 ( .A(n23569), .ZN(n23571) );
  AOI21_X1 U32353 ( .B1(n23572), .B2(n23571), .A(n23570), .ZN(n23573) );
  XNOR2_X1 U32354 ( .A(n26435), .B(n26589), .ZN(n23579) );
  XNOR2_X1 U32355 ( .A(n26239), .B(n23580), .ZN(n24654) );
  XNOR2_X1 U32356 ( .A(n4048), .B(n4026), .ZN(n45333) );
  XNOR2_X1 U32357 ( .A(n25493), .B(n45333), .ZN(n27306) );
  XNOR2_X1 U32358 ( .A(n25860), .B(n27306), .ZN(n23588) );
  INV_X1 U32359 ( .A(n23581), .ZN(n23583) );
  XNOR2_X1 U32360 ( .A(n25520), .B(n4803), .ZN(n23582) );
  XNOR2_X1 U32361 ( .A(n23583), .B(n23582), .ZN(n44072) );
  XNOR2_X1 U32362 ( .A(n42549), .B(n42322), .ZN(n23584) );
  XNOR2_X1 U32363 ( .A(n44072), .B(n23584), .ZN(n23585) );
  XNOR2_X1 U32364 ( .A(n28214), .B(n23585), .ZN(n23586) );
  XNOR2_X1 U32365 ( .A(n23586), .B(n25506), .ZN(n23587) );
  XNOR2_X1 U32366 ( .A(n23588), .B(n23587), .ZN(n23589) );
  XNOR2_X1 U32367 ( .A(n24654), .B(n23589), .ZN(n23654) );
  NAND3_X1 U32368 ( .A1(n23614), .A2(n23613), .A3(n17420), .ZN(n23603) );
  NAND3_X1 U32371 ( .A1(n23599), .A2(n23598), .A3(n23597), .ZN(n23600) );
  AND3_X1 U32372 ( .A1(n23602), .A2(n23601), .A3(n23600), .ZN(n23619) );
  INV_X1 U32373 ( .A(n23603), .ZN(n23608) );
  INV_X1 U32374 ( .A(n23604), .ZN(n23605) );
  AOI22_X1 U32375 ( .A1(n23608), .A2(n23607), .B1(n23606), .B2(n23605), .ZN(
        n23618) );
  INV_X1 U32376 ( .A(n24208), .ZN(n23617) );
  INV_X1 U32377 ( .A(n23610), .ZN(n23612) );
  OAI21_X1 U32378 ( .B1(n23613), .B2(n23612), .A(n23611), .ZN(n23616) );
  INV_X1 U32379 ( .A(n23614), .ZN(n23615) );
  XNOR2_X2 U32380 ( .A(n27309), .B(n23621), .ZN(n26235) );
  NAND2_X1 U32381 ( .A1(n23637), .A2(n23961), .ZN(n23624) );
  NAND2_X1 U32382 ( .A1(n5068), .A2(n23624), .ZN(n23629) );
  INV_X1 U32383 ( .A(n23625), .ZN(n23626) );
  OAI211_X1 U32384 ( .C1(n23626), .C2(n23958), .A(n23955), .B(n23961), .ZN(
        n23627) );
  INV_X1 U32385 ( .A(n23627), .ZN(n23628) );
  AOI21_X1 U32386 ( .B1(n23630), .B2(n23629), .A(n23628), .ZN(n23650) );
  NAND4_X1 U32387 ( .A1(n23963), .A2(n23638), .A3(n5069), .A4(n23637), .ZN(
        n23632) );
  MUX2_X1 U32388 ( .A(n23633), .B(n23632), .S(n23641), .Z(n23648) );
  INV_X1 U32389 ( .A(n23634), .ZN(n23951) );
  INV_X1 U32390 ( .A(n23635), .ZN(n23636) );
  OAI21_X1 U32391 ( .B1(n23951), .B2(n23950), .A(n23636), .ZN(n23640) );
  NAND2_X1 U32392 ( .A1(n23637), .A2(n559), .ZN(n23642) );
  OAI21_X1 U32393 ( .B1(n23638), .B2(n23642), .A(n23641), .ZN(n23639) );
  NOR2_X1 U32394 ( .A1(n23955), .A2(n23641), .ZN(n23952) );
  NAND2_X1 U32395 ( .A1(n23642), .A2(n23950), .ZN(n23643) );
  NAND2_X1 U32396 ( .A1(n23952), .A2(n23643), .ZN(n23644) );
  XNOR2_X2 U32398 ( .A(n26235), .B(n27439), .ZN(n28218) );
  XNOR2_X1 U32399 ( .A(n28218), .B(n23652), .ZN(n23653) );
  OR2_X1 U32400 ( .A1(n29907), .A2(n30785), .ZN(n29895) );
  NAND3_X1 U32401 ( .A1(n26828), .A2(n30783), .A3(n23658), .ZN(n23656) );
  NAND3_X1 U32402 ( .A1(n29909), .A2(n29908), .A3(n30789), .ZN(n23655) );
  NAND2_X1 U32404 ( .A1(n30790), .A2(n1042), .ZN(n23659) );
  OR2_X1 U32405 ( .A1(n29899), .A2(n23659), .ZN(n26833) );
  NAND2_X1 U32406 ( .A1(n29900), .A2(n27566), .ZN(n30794) );
  OAI21_X1 U32407 ( .B1(n27570), .B2(n23660), .A(n30794), .ZN(n23662) );
  OR2_X1 U32408 ( .A1(n30794), .A2(n29901), .ZN(n27411) );
  NOR2_X1 U32409 ( .A1(n32236), .A2(n32252), .ZN(n30839) );
  XNOR2_X1 U32410 ( .A(n23977), .B(n2106), .ZN(n24511) );
  OAI21_X1 U32411 ( .B1(n24028), .B2(n23665), .A(n24033), .ZN(n23678) );
  NAND3_X1 U32412 ( .A1(n23668), .A2(n24041), .A3(n24034), .ZN(n23669) );
  AND2_X1 U32413 ( .A1(n23673), .A2(n23672), .ZN(n23677) );
  NAND3_X1 U32414 ( .A1(n23675), .A2(n23674), .A3(n24030), .ZN(n23676) );
  XNOR2_X1 U32415 ( .A(n28048), .B(n25946), .ZN(n24842) );
  BUF_X2 U32416 ( .A(n24842), .Z(n28249) );
  XNOR2_X1 U32417 ( .A(n28249), .B(n24511), .ZN(n23686) );
  XNOR2_X1 U32418 ( .A(n26565), .B(n28381), .ZN(n23684) );
  XNOR2_X1 U32419 ( .A(n45107), .B(n4605), .ZN(n23679) );
  XNOR2_X1 U32420 ( .A(n23679), .B(n41155), .ZN(n23680) );
  XNOR2_X1 U32421 ( .A(n42630), .B(n43150), .ZN(n25341) );
  XNOR2_X1 U32422 ( .A(n23680), .B(n25341), .ZN(n23681) );
  XNOR2_X1 U32423 ( .A(n42241), .B(n34411), .ZN(n33254) );
  XNOR2_X1 U32424 ( .A(n23681), .B(n33254), .ZN(n44350) );
  XNOR2_X1 U32425 ( .A(n2608), .B(n4312), .ZN(n42102) );
  XNOR2_X1 U32426 ( .A(n44350), .B(n42102), .ZN(n23682) );
  XNOR2_X1 U32427 ( .A(n23684), .B(n23683), .ZN(n23685) );
  XNOR2_X1 U32428 ( .A(n23686), .B(n23685), .ZN(n23687) );
  XNOR2_X1 U32429 ( .A(n23687), .B(n23688), .ZN(n23691) );
  XNOR2_X1 U32430 ( .A(n51667), .B(n28049), .ZN(n24856) );
  XNOR2_X1 U32431 ( .A(n24856), .B(n24855), .ZN(n25035) );
  XNOR2_X1 U32432 ( .A(n25816), .B(n25127), .ZN(n23689) );
  XNOR2_X1 U32433 ( .A(n25035), .B(n23689), .ZN(n23690) );
  XNOR2_X1 U32434 ( .A(n23691), .B(n23690), .ZN(n23809) );
  INV_X1 U32435 ( .A(n23809), .ZN(n27600) );
  AOI21_X1 U32436 ( .B1(n24332), .B2(n23702), .A(n5415), .ZN(n23698) );
  INV_X1 U32437 ( .A(n23692), .ZN(n23697) );
  NAND4_X1 U32438 ( .A1(n23695), .A2(n24336), .A3(n23694), .A4(n23693), .ZN(
        n23696) );
  NAND4_X1 U32439 ( .A1(n23701), .A2(n23703), .A3(n24336), .A4(n23700), .ZN(
        n23710) );
  XNOR2_X1 U32440 ( .A(n23711), .B(n42769), .ZN(n43906) );
  XNOR2_X1 U32441 ( .A(n43906), .B(n46062), .ZN(n23715) );
  XNOR2_X1 U32442 ( .A(n25040), .B(n29662), .ZN(n23713) );
  XNOR2_X1 U32443 ( .A(n4415), .B(n75), .ZN(n24694) );
  XNOR2_X1 U32444 ( .A(n2605), .B(n24694), .ZN(n23712) );
  XNOR2_X1 U32445 ( .A(n23713), .B(n23712), .ZN(n23714) );
  XNOR2_X1 U32446 ( .A(n23714), .B(n26296), .ZN(n45289) );
  XNOR2_X1 U32447 ( .A(n23715), .B(n45289), .ZN(n23716) );
  XNOR2_X1 U32448 ( .A(n25724), .B(n23716), .ZN(n23717) );
  XNOR2_X1 U32449 ( .A(n26556), .B(n488), .ZN(n26155) );
  XNOR2_X1 U32450 ( .A(n25726), .B(n28276), .ZN(n24577) );
  INV_X1 U32451 ( .A(n24577), .ZN(n24052) );
  XNOR2_X1 U32452 ( .A(n23719), .B(n24052), .ZN(n23720) );
  XNOR2_X1 U32453 ( .A(n23721), .B(n23720), .ZN(n23858) );
  INV_X1 U32454 ( .A(n23858), .ZN(n30667) );
  INV_X1 U32455 ( .A(n42846), .ZN(n36968) );
  XNOR2_X1 U32456 ( .A(n43850), .B(n23722), .ZN(n41313) );
  XNOR2_X1 U32457 ( .A(n36968), .B(n41313), .ZN(n23723) );
  XNOR2_X1 U32458 ( .A(n28396), .B(n23723), .ZN(n23724) );
  XNOR2_X1 U32459 ( .A(n23725), .B(n23724), .ZN(n23726) );
  XNOR2_X1 U32460 ( .A(n23726), .B(n25387), .ZN(n23729) );
  INV_X1 U32461 ( .A(n26530), .ZN(n23727) );
  XNOR2_X1 U32462 ( .A(n24344), .B(n23727), .ZN(n24464) );
  XNOR2_X1 U32463 ( .A(n51752), .B(n24464), .ZN(n23728) );
  XNOR2_X1 U32464 ( .A(n23729), .B(n23728), .ZN(n23743) );
  NAND2_X1 U32465 ( .A1(n24097), .A2(n24105), .ZN(n23740) );
  OAI21_X1 U32466 ( .B1(n23732), .B2(n23731), .A(n24414), .ZN(n23733) );
  NAND2_X1 U32467 ( .A1(n23733), .A2(n24100), .ZN(n23739) );
  NOR2_X1 U32468 ( .A1(n23734), .A2(n24119), .ZN(n23735) );
  NOR2_X1 U32469 ( .A1(n24072), .A2(n23735), .ZN(n23738) );
  NOR2_X1 U32470 ( .A1(n24409), .A2(n24412), .ZN(n24120) );
  OAI21_X1 U32471 ( .B1(n23736), .B2(n24065), .A(n24120), .ZN(n23737) );
  XNOR2_X1 U32472 ( .A(n28126), .B(n25444), .ZN(n23741) );
  XNOR2_X1 U32473 ( .A(n23741), .B(n27502), .ZN(n24631) );
  INV_X1 U32474 ( .A(n1354), .ZN(n49867) );
  XNOR2_X1 U32475 ( .A(n25540), .B(n49867), .ZN(n23742) );
  XNOR2_X1 U32476 ( .A(n24556), .B(n23742), .ZN(n24310) );
  XNOR2_X1 U32477 ( .A(n24631), .B(n24310), .ZN(n25103) );
  XNOR2_X1 U32478 ( .A(n24319), .B(n25829), .ZN(n24872) );
  NOR2_X1 U32479 ( .A1(n24687), .A2(n27609), .ZN(n23808) );
  NAND2_X1 U32480 ( .A1(n23858), .A2(n23809), .ZN(n26909) );
  NOR2_X1 U32481 ( .A1(n26909), .A2(n30665), .ZN(n23807) );
  MUX2_X1 U32482 ( .A(n23746), .B(n24186), .S(n2210), .Z(n23749) );
  AND2_X1 U32483 ( .A1(n4462), .A2(n23747), .ZN(n23748) );
  NAND2_X1 U32484 ( .A1(n23749), .A2(n23748), .ZN(n23771) );
  NAND2_X1 U32485 ( .A1(n24190), .A2(n23751), .ZN(n23753) );
  OAI211_X1 U32486 ( .C1(n23754), .C2(n4462), .A(n23753), .B(n23752), .ZN(
        n23760) );
  XNOR2_X1 U32487 ( .A(n2210), .B(n24188), .ZN(n23758) );
  NOR2_X1 U32488 ( .A1(n24188), .A2(n22605), .ZN(n24192) );
  NAND2_X1 U32489 ( .A1(n24192), .A2(n24190), .ZN(n23757) );
  AND4_X1 U32491 ( .A1(n23757), .A2(n23758), .A3(n24187), .A4(n23869), .ZN(
        n23759) );
  NOR2_X1 U32492 ( .A1(n23760), .A2(n23759), .ZN(n23770) );
  INV_X1 U32493 ( .A(n23763), .ZN(n23765) );
  OAI21_X1 U32494 ( .B1(n24179), .B2(n23767), .A(n23766), .ZN(n23768) );
  XNOR2_X1 U32495 ( .A(n25755), .B(n23772), .ZN(n24651) );
  XNOR2_X1 U32496 ( .A(n27242), .B(n24651), .ZN(n24814) );
  INV_X1 U32497 ( .A(n24814), .ZN(n23937) );
  XNOR2_X1 U32498 ( .A(n23773), .B(n31432), .ZN(n45071) );
  XNOR2_X1 U32499 ( .A(n42712), .B(n4835), .ZN(n23774) );
  XNOR2_X1 U32500 ( .A(n26589), .B(n28213), .ZN(n24132) );
  XNOR2_X1 U32501 ( .A(n23775), .B(n24132), .ZN(n23776) );
  XNOR2_X1 U32502 ( .A(n23776), .B(n51512), .ZN(n23779) );
  XNOR2_X1 U32503 ( .A(n25860), .B(n27289), .ZN(n23778) );
  XNOR2_X1 U32504 ( .A(n34215), .B(n4737), .ZN(n44155) );
  XNOR2_X1 U32505 ( .A(n27309), .B(n44155), .ZN(n25763) );
  XNOR2_X1 U32506 ( .A(n25506), .B(n4204), .ZN(n24128) );
  XNOR2_X1 U32507 ( .A(n25763), .B(n24128), .ZN(n23777) );
  XNOR2_X1 U32508 ( .A(n51719), .B(n41367), .ZN(n23791) );
  NAND2_X1 U32509 ( .A1(n23782), .A2(n24245), .ZN(n23783) );
  MUX2_X1 U32510 ( .A(n24246), .B(n23783), .S(n24238), .Z(n23790) );
  OR2_X1 U32511 ( .A1(n23787), .A2(n24248), .ZN(n23788) );
  XNOR2_X1 U32512 ( .A(n23791), .B(n25483), .ZN(n25010) );
  INV_X1 U32513 ( .A(n25010), .ZN(n23792) );
  XNOR2_X1 U32514 ( .A(n23793), .B(n23792), .ZN(n23795) );
  XNOR2_X1 U32516 ( .A(n23794), .B(n51750), .ZN(n24756) );
  XNOR2_X1 U32517 ( .A(n24756), .B(n23795), .ZN(n23805) );
  XNOR2_X1 U32518 ( .A(n23796), .B(n4712), .ZN(n42876) );
  XNOR2_X1 U32519 ( .A(n43739), .B(n4895), .ZN(n23797) );
  XNOR2_X1 U32520 ( .A(n42876), .B(n23797), .ZN(n23798) );
  XNOR2_X1 U32521 ( .A(n41403), .B(n23798), .ZN(n23799) );
  XNOR2_X1 U32522 ( .A(n25778), .B(n23799), .ZN(n23800) );
  XNOR2_X1 U32523 ( .A(n23801), .B(n23800), .ZN(n23802) );
  XNOR2_X1 U32524 ( .A(n23802), .B(n28357), .ZN(n23803) );
  XNOR2_X1 U32525 ( .A(n24171), .B(n25700), .ZN(n27480) );
  INV_X1 U32526 ( .A(n27480), .ZN(n24608) );
  XNOR2_X1 U32527 ( .A(n24608), .B(n23803), .ZN(n23804) );
  INV_X1 U32528 ( .A(n27602), .ZN(n30670) );
  OAI21_X1 U32529 ( .B1(n23808), .B2(n23807), .A(n23806), .ZN(n23856) );
  NAND2_X1 U32530 ( .A1(n30663), .A2(n27602), .ZN(n30664) );
  OAI21_X1 U32532 ( .B1(n30664), .B2(n51492), .A(n26856), .ZN(n23854) );
  AND2_X1 U32533 ( .A1(n30662), .A2(n27609), .ZN(n24679) );
  XNOR2_X1 U32534 ( .A(n27382), .B(n26100), .ZN(n28438) );
  NAND3_X1 U32535 ( .A1(n23812), .A2(n23811), .A3(n51753), .ZN(n23817) );
  NAND3_X1 U32536 ( .A1(n23815), .A2(n23814), .A3(n23813), .ZN(n23816) );
  NAND3_X1 U32537 ( .A1(n23818), .A2(n23817), .A3(n23816), .ZN(n23819) );
  NAND4_X1 U32538 ( .A1(n23822), .A2(n24150), .A3(n24159), .A4(n23832), .ZN(
        n23823) );
  NAND2_X1 U32539 ( .A1(n23826), .A2(n23825), .ZN(n24154) );
  NAND3_X1 U32540 ( .A1(n24148), .A2(n23830), .A3(n23829), .ZN(n23838) );
  NAND2_X1 U32541 ( .A1(n23831), .A2(n24161), .ZN(n23837) );
  OAI211_X1 U32542 ( .C1(n23835), .C2(n23834), .A(n23833), .B(n23832), .ZN(
        n23836) );
  XNOR2_X1 U32544 ( .A(n23840), .B(n25920), .ZN(n27384) );
  INV_X1 U32545 ( .A(n27384), .ZN(n27447) );
  XNOR2_X1 U32546 ( .A(n28427), .B(n43662), .ZN(n24825) );
  INV_X1 U32547 ( .A(n24825), .ZN(n23842) );
  XNOR2_X1 U32548 ( .A(n23843), .B(n25143), .ZN(n23844) );
  XNOR2_X1 U32549 ( .A(n23844), .B(n28317), .ZN(n23853) );
  XNOR2_X1 U32550 ( .A(n28311), .B(n25320), .ZN(n26106) );
  XNOR2_X1 U32551 ( .A(n26204), .B(n23845), .ZN(n43970) );
  XNOR2_X1 U32552 ( .A(n23846), .B(n4909), .ZN(n23847) );
  XNOR2_X1 U32553 ( .A(n23847), .B(n24057), .ZN(n45254) );
  XNOR2_X1 U32554 ( .A(n43970), .B(n45254), .ZN(n23848) );
  XNOR2_X1 U32555 ( .A(n25213), .B(n23848), .ZN(n23849) );
  XNOR2_X1 U32556 ( .A(n26106), .B(n23849), .ZN(n23851) );
  XNOR2_X1 U32557 ( .A(n23850), .B(n23851), .ZN(n23852) );
  XNOR2_X1 U32558 ( .A(n27452), .B(n47737), .ZN(n25084) );
  NAND3_X1 U32559 ( .A1(n23854), .A2(n24679), .A3(n3819), .ZN(n23855) );
  OR2_X1 U32560 ( .A1(n30664), .A2(n26909), .ZN(n26860) );
  NAND2_X1 U32561 ( .A1(n23859), .A2(n27602), .ZN(n26914) );
  OR2_X1 U32562 ( .A1(n26914), .A2(n51492), .ZN(n24683) );
  NOR2_X1 U32563 ( .A1(n26914), .A2(n30665), .ZN(n27607) );
  NAND2_X1 U32564 ( .A1(n51492), .A2(n27600), .ZN(n30661) );
  NOR2_X1 U32565 ( .A1(n30661), .A2(n27604), .ZN(n23860) );
  AND2_X1 U32566 ( .A1(n23859), .A2(n23861), .ZN(n27605) );
  AOI22_X1 U32567 ( .A1(n27607), .A2(n23860), .B1(n27605), .B2(n30670), .ZN(
        n23863) );
  INV_X1 U32568 ( .A(n23864), .ZN(n23877) );
  INV_X1 U32569 ( .A(n23865), .ZN(n23867) );
  OR2_X1 U32570 ( .A1(n23867), .A2(n4328), .ZN(n23876) );
  INV_X1 U32573 ( .A(n23872), .ZN(n23873) );
  MUX2_X1 U32574 ( .A(n23874), .B(n23873), .S(n24183), .Z(n23875) );
  XNOR2_X1 U32575 ( .A(n26448), .B(n51720), .ZN(n23878) );
  XNOR2_X1 U32576 ( .A(n25291), .B(n23878), .ZN(n28067) );
  XNOR2_X1 U32577 ( .A(n27272), .B(n51749), .ZN(n25485) );
  XNOR2_X1 U32578 ( .A(n51648), .B(n4923), .ZN(n25604) );
  INV_X1 U32579 ( .A(n25883), .ZN(n23880) );
  INV_X1 U32580 ( .A(n28242), .ZN(n23881) );
  XNOR2_X1 U32581 ( .A(n23882), .B(n4926), .ZN(n23883) );
  XNOR2_X1 U32582 ( .A(n23884), .B(n23883), .ZN(n42261) );
  XNOR2_X1 U32583 ( .A(n24936), .B(n42261), .ZN(n23885) );
  XNOR2_X1 U32584 ( .A(n23885), .B(n24757), .ZN(n27265) );
  XNOR2_X1 U32585 ( .A(n23887), .B(n23886), .ZN(n23889) );
  XNOR2_X1 U32586 ( .A(n23889), .B(n23888), .ZN(n44497) );
  XNOR2_X1 U32587 ( .A(n27322), .B(n44497), .ZN(n23890) );
  XNOR2_X1 U32588 ( .A(n23890), .B(n24795), .ZN(n23891) );
  XNOR2_X1 U32589 ( .A(n27265), .B(n23891), .ZN(n23892) );
  XNOR2_X1 U32590 ( .A(n23892), .B(n27330), .ZN(n23893) );
  XNOR2_X1 U32591 ( .A(n27241), .B(n25669), .ZN(n23894) );
  NOR2_X1 U32592 ( .A1(n23895), .A2(n23906), .ZN(n23903) );
  AOI21_X1 U32593 ( .B1(n23897), .B2(n23903), .A(n23896), .ZN(n23900) );
  INV_X1 U32594 ( .A(n23898), .ZN(n23899) );
  MUX2_X1 U32595 ( .A(n23901), .B(n23900), .S(n23899), .Z(n23929) );
  NAND3_X1 U32597 ( .A1(n23907), .A2(n23906), .A3(n23905), .ZN(n23917) );
  INV_X1 U32598 ( .A(n23909), .ZN(n23910) );
  NAND3_X1 U32599 ( .A1(n23912), .A2(n23911), .A3(n23910), .ZN(n23916) );
  INV_X1 U32600 ( .A(n23919), .ZN(n23920) );
  NOR2_X1 U32601 ( .A1(n23921), .A2(n23920), .ZN(n23922) );
  NAND2_X1 U32602 ( .A1(n23927), .A2(n23926), .ZN(n23928) );
  XNOR2_X1 U32603 ( .A(n23621), .B(n28220), .ZN(n23930) );
  XNOR2_X1 U32604 ( .A(n43768), .B(n34463), .ZN(n23933) );
  XNOR2_X1 U32605 ( .A(n43766), .B(n4613), .ZN(n23931) );
  XNOR2_X1 U32606 ( .A(n43764), .B(n43263), .ZN(n24479) );
  XNOR2_X1 U32607 ( .A(n23931), .B(n24479), .ZN(n23932) );
  XNOR2_X1 U32608 ( .A(n23933), .B(n23932), .ZN(n23934) );
  XNOR2_X1 U32609 ( .A(n25501), .B(n23934), .ZN(n23936) );
  XNOR2_X1 U32610 ( .A(n26589), .B(n27303), .ZN(n23935) );
  INV_X1 U32611 ( .A(n24091), .ZN(n30683) );
  XNOR2_X1 U32612 ( .A(n24319), .B(n24548), .ZN(n23940) );
  XNOR2_X1 U32613 ( .A(n23940), .B(n25829), .ZN(n28131) );
  XNOR2_X1 U32614 ( .A(n23941), .B(n471), .ZN(n23948) );
  INV_X1 U32615 ( .A(n34451), .ZN(n23942) );
  XNOR2_X1 U32616 ( .A(n23942), .B(n1313), .ZN(n42227) );
  XNOR2_X1 U32617 ( .A(n23943), .B(n4694), .ZN(n23944) );
  XNOR2_X1 U32618 ( .A(n25436), .B(n23944), .ZN(n44522) );
  XNOR2_X1 U32619 ( .A(n42227), .B(n44522), .ZN(n23945) );
  XNOR2_X1 U32620 ( .A(n24344), .B(n23945), .ZN(n23946) );
  XNOR2_X1 U32621 ( .A(n25229), .B(n25909), .ZN(n25446) );
  XNOR2_X1 U32622 ( .A(n23946), .B(n25446), .ZN(n23947) );
  XNOR2_X1 U32623 ( .A(n23948), .B(n23947), .ZN(n23949) );
  XNOR2_X1 U32624 ( .A(n23949), .B(n28131), .ZN(n23973) );
  AND2_X1 U32625 ( .A1(n23951), .A2(n23950), .ZN(n23954) );
  AOI21_X1 U32626 ( .B1(n23954), .B2(n23953), .A(n23952), .ZN(n23969) );
  OAI211_X1 U32627 ( .C1(n23958), .C2(n559), .A(n23956), .B(n23955), .ZN(
        n23960) );
  NAND2_X1 U32628 ( .A1(n23960), .A2(n23959), .ZN(n23968) );
  NAND2_X1 U32629 ( .A1(n23962), .A2(n23961), .ZN(n23967) );
  XNOR2_X1 U32630 ( .A(n28121), .B(n51121), .ZN(n23970) );
  XNOR2_X1 U32631 ( .A(n23971), .B(n23970), .ZN(n23972) );
  XNOR2_X1 U32632 ( .A(n23973), .B(n23972), .ZN(n29933) );
  XNOR2_X1 U32634 ( .A(n28257), .B(n4343), .ZN(n23975) );
  XNOR2_X1 U32635 ( .A(n23975), .B(n27197), .ZN(n23976) );
  XNOR2_X1 U32636 ( .A(n25805), .B(n23976), .ZN(n27341) );
  INV_X1 U32637 ( .A(n27424), .ZN(n27200) );
  XNOR2_X1 U32638 ( .A(n27200), .B(n51751), .ZN(n23978) );
  XNOR2_X1 U32639 ( .A(n23978), .B(n23977), .ZN(n25475) );
  XNOR2_X1 U32640 ( .A(n26571), .B(n51380), .ZN(n24915) );
  INV_X1 U32641 ( .A(n24915), .ZN(n23979) );
  XNOR2_X1 U32642 ( .A(n23980), .B(n23979), .ZN(n24015) );
  NAND3_X1 U32643 ( .A1(n23983), .A2(n23982), .A3(n23981), .ZN(n23985) );
  OAI211_X1 U32644 ( .C1(n23987), .C2(n23986), .A(n23985), .B(n23984), .ZN(
        n23988) );
  OAI21_X1 U32645 ( .B1(n23990), .B2(n23989), .A(n23988), .ZN(n23994) );
  AOI21_X1 U32646 ( .B1(n23994), .B2(n23993), .A(n23992), .ZN(n24008) );
  OAI211_X1 U32647 ( .C1(n24001), .C2(n24000), .A(n23999), .B(n23998), .ZN(
        n24005) );
  NAND2_X1 U32648 ( .A1(n24003), .A2(n24002), .ZN(n24004) );
  XNOR2_X1 U32649 ( .A(n27196), .B(n4793), .ZN(n26279) );
  INV_X1 U32650 ( .A(n28251), .ZN(n24009) );
  XNOR2_X1 U32651 ( .A(n24010), .B(n24009), .ZN(n40222) );
  XNOR2_X1 U32652 ( .A(n33733), .B(n35107), .ZN(n42934) );
  XNOR2_X1 U32653 ( .A(n42934), .B(n4565), .ZN(n24011) );
  XNOR2_X1 U32654 ( .A(n26279), .B(n24012), .ZN(n24013) );
  XNOR2_X1 U32655 ( .A(n25035), .B(n24013), .ZN(n24014) );
  AND2_X1 U32656 ( .A1(n24091), .A2(n29940), .ZN(n30399) );
  INV_X1 U32657 ( .A(n24016), .ZN(n24021) );
  INV_X1 U32658 ( .A(n24017), .ZN(n24020) );
  INV_X1 U32659 ( .A(n24018), .ZN(n24019) );
  OAI21_X1 U32660 ( .B1(n24021), .B2(n24020), .A(n24019), .ZN(n24022) );
  XNOR2_X1 U32661 ( .A(n28038), .B(n25724), .ZN(n24046) );
  OAI21_X1 U32662 ( .B1(n24033), .B2(n24026), .A(n24025), .ZN(n24027) );
  NAND2_X1 U32663 ( .A1(n24028), .A2(n24027), .ZN(n24045) );
  AOI21_X1 U32664 ( .B1(n24036), .B2(n354), .A(n24041), .ZN(n24031) );
  OAI21_X1 U32665 ( .B1(n24031), .B2(n24030), .A(n24033), .ZN(n24040) );
  NAND2_X1 U32666 ( .A1(n24036), .A2(n24041), .ZN(n24039) );
  INV_X1 U32667 ( .A(n24032), .ZN(n24037) );
  AOI21_X1 U32668 ( .B1(n7494), .B2(n24034), .A(n22101), .ZN(n24035) );
  OAI21_X1 U32669 ( .B1(n24037), .B2(n24036), .A(n24035), .ZN(n24038) );
  OAI21_X1 U32670 ( .B1(n24043), .B2(n24042), .A(n24041), .ZN(n24044) );
  XNOR2_X1 U32671 ( .A(n24046), .B(n51416), .ZN(n25259) );
  XNOR2_X1 U32672 ( .A(n24047), .B(n44330), .ZN(n25071) );
  XNOR2_X1 U32673 ( .A(n25457), .B(n1326), .ZN(n25727) );
  INV_X1 U32674 ( .A(n38860), .ZN(n24048) );
  XNOR2_X1 U32675 ( .A(n24048), .B(n4659), .ZN(n37121) );
  XNOR2_X1 U32676 ( .A(n37121), .B(n43053), .ZN(n24049) );
  XNOR2_X1 U32677 ( .A(n26375), .B(n24049), .ZN(n24050) );
  XNOR2_X1 U32678 ( .A(n25047), .B(n24050), .ZN(n24051) );
  XNOR2_X1 U32679 ( .A(n24051), .B(n488), .ZN(n24053) );
  XNOR2_X1 U32680 ( .A(n24053), .B(n24052), .ZN(n24054) );
  NOR2_X1 U32681 ( .A1(n24091), .A2(n402), .ZN(n24088) );
  XNOR2_X1 U32682 ( .A(n28430), .B(n27450), .ZN(n24063) );
  XNOR2_X1 U32683 ( .A(n24055), .B(n4568), .ZN(n42998) );
  XNOR2_X1 U32684 ( .A(n24057), .B(n24056), .ZN(n24058) );
  XNOR2_X1 U32685 ( .A(n24059), .B(n24058), .ZN(n37474) );
  XNOR2_X1 U32686 ( .A(n37474), .B(n42995), .ZN(n24060) );
  XNOR2_X1 U32687 ( .A(n42998), .B(n24060), .ZN(n24061) );
  XNOR2_X1 U32688 ( .A(n25213), .B(n24061), .ZN(n24062) );
  XNOR2_X1 U32689 ( .A(n24063), .B(n24062), .ZN(n24082) );
  OAI21_X1 U32690 ( .B1(n24098), .B2(n24411), .A(n24105), .ZN(n24064) );
  INV_X1 U32691 ( .A(n24064), .ZN(n24066) );
  AOI21_X1 U32692 ( .B1(n24067), .B2(n24066), .A(n24065), .ZN(n24081) );
  NAND2_X1 U32693 ( .A1(n24068), .A2(n24413), .ZN(n24080) );
  NAND4_X1 U32694 ( .A1(n24112), .A2(n24111), .A3(n24412), .A4(n24105), .ZN(
        n24069) );
  OAI211_X1 U32695 ( .C1(n24071), .C2(n24074), .A(n24070), .B(n24069), .ZN(
        n24073) );
  NOR2_X1 U32696 ( .A1(n24073), .A2(n24072), .ZN(n24079) );
  AOI21_X1 U32697 ( .B1(n4726), .B2(n24413), .A(n24098), .ZN(n24077) );
  INV_X1 U32698 ( .A(n24113), .ZN(n24075) );
  NAND2_X1 U32699 ( .A1(n24413), .A2(n24412), .ZN(n24410) );
  OAI21_X1 U32700 ( .B1(n24075), .B2(n24074), .A(n24410), .ZN(n24076) );
  OAI21_X1 U32701 ( .B1(n24077), .B2(n24414), .A(n24076), .ZN(n24078) );
  OAI211_X1 U32702 ( .C1(n24081), .C2(n24080), .A(n24079), .B(n24078), .ZN(
        n24302) );
  XNOR2_X1 U32703 ( .A(n24082), .B(n370), .ZN(n24085) );
  INV_X1 U32704 ( .A(n24083), .ZN(n24084) );
  XNOR2_X1 U32705 ( .A(n24085), .B(n24084), .ZN(n24086) );
  AOI22_X1 U32706 ( .A1(n30399), .A2(n30696), .B1(n24088), .B2(n734), .ZN(
        n24089) );
  OAI211_X1 U32707 ( .C1(n27528), .C2(n402), .A(n24089), .B(n30396), .ZN(
        n24090) );
  INV_X1 U32708 ( .A(n24090), .ZN(n24362) );
  NAND2_X1 U32709 ( .A1(n30683), .A2(n29940), .ZN(n29931) );
  AND2_X1 U32710 ( .A1(n30692), .A2(n51113), .ZN(n30690) );
  NAND2_X1 U32711 ( .A1(n24093), .A2(n30690), .ZN(n24095) );
  OAI21_X1 U32712 ( .B1(n1906), .B2(n30688), .A(n30392), .ZN(n24094) );
  NAND2_X1 U32713 ( .A1(n24096), .A2(n29938), .ZN(n24361) );
  OR2_X1 U32714 ( .A1(n32251), .A2(n31781), .ZN(n31241) );
  XNOR2_X1 U32715 ( .A(n24105), .B(n24117), .ZN(n24099) );
  NAND4_X1 U32716 ( .A1(n24099), .A2(n24409), .A3(n24098), .A4(n24413), .ZN(
        n24109) );
  NAND2_X1 U32717 ( .A1(n24101), .A2(n24100), .ZN(n24104) );
  NAND2_X1 U32718 ( .A1(n24102), .A2(n24106), .ZN(n24103) );
  AOI21_X1 U32719 ( .B1(n24105), .B2(n24409), .A(n24414), .ZN(n24108) );
  NAND3_X1 U32720 ( .A1(n24109), .A2(n24108), .A3(n24107), .ZN(n24110) );
  NAND4_X1 U32721 ( .A1(n24113), .A2(n24117), .A3(n24112), .A4(n24111), .ZN(
        n24114) );
  OAI211_X1 U32722 ( .C1(n24117), .C2(n24116), .A(n24115), .B(n24114), .ZN(
        n24126) );
  INV_X1 U32723 ( .A(n24120), .ZN(n24118) );
  NAND2_X1 U32724 ( .A1(n24118), .A2(n24414), .ZN(n24124) );
  INV_X1 U32725 ( .A(n24119), .ZN(n24121) );
  INV_X1 U32726 ( .A(n24127), .ZN(n42291) );
  XNOR2_X1 U32728 ( .A(n27290), .B(n25360), .ZN(n24129) );
  XNOR2_X1 U32729 ( .A(n51483), .B(n24128), .ZN(n26237) );
  XNOR2_X1 U32730 ( .A(n24129), .B(n26237), .ZN(n24135) );
  XNOR2_X1 U32731 ( .A(n42293), .B(n44483), .ZN(n24130) );
  XNOR2_X1 U32732 ( .A(n27295), .B(n24130), .ZN(n24131) );
  XNOR2_X1 U32733 ( .A(n24132), .B(n24131), .ZN(n24133) );
  XNOR2_X1 U32734 ( .A(n25188), .B(n24133), .ZN(n24134) );
  XNOR2_X1 U32735 ( .A(n24134), .B(n24135), .ZN(n24139) );
  INV_X1 U32736 ( .A(n25352), .ZN(n26248) );
  XNOR2_X1 U32737 ( .A(n25669), .B(n4526), .ZN(n25859) );
  XNOR2_X1 U32738 ( .A(n26248), .B(n25859), .ZN(n25529) );
  INV_X1 U32739 ( .A(n25529), .ZN(n24137) );
  XNOR2_X1 U32740 ( .A(n25860), .B(n25664), .ZN(n27311) );
  INV_X1 U32741 ( .A(n27311), .ZN(n24136) );
  XNOR2_X1 U32742 ( .A(n24137), .B(n24136), .ZN(n24138) );
  XNOR2_X1 U32743 ( .A(n24138), .B(n24139), .ZN(n24265) );
  XNOR2_X1 U32744 ( .A(n750), .B(n24140), .ZN(n24143) );
  XNOR2_X1 U32745 ( .A(n24616), .B(n41740), .ZN(n24141) );
  XNOR2_X1 U32746 ( .A(n24141), .B(n28353), .ZN(n26268) );
  INV_X1 U32747 ( .A(n26268), .ZN(n24142) );
  XNOR2_X1 U32748 ( .A(n24143), .B(n24142), .ZN(n24165) );
  XNOR2_X1 U32749 ( .A(n24144), .B(n24757), .ZN(n24164) );
  NOR2_X1 U32751 ( .A1(n24151), .A2(n24150), .ZN(n24152) );
  NOR2_X1 U32752 ( .A1(n24153), .A2(n24152), .ZN(n24163) );
  INV_X1 U32753 ( .A(n24154), .ZN(n24156) );
  NAND4_X1 U32754 ( .A1(n24161), .A2(n24160), .A3(n24159), .A4(n24158), .ZN(
        n24162) );
  XNOR2_X1 U32755 ( .A(n24164), .B(n25610), .ZN(n28364) );
  XNOR2_X1 U32756 ( .A(n24165), .B(n28364), .ZN(n24175) );
  XNOR2_X1 U32757 ( .A(n25013), .B(n4865), .ZN(n24383) );
  XNOR2_X1 U32758 ( .A(n24383), .B(n4712), .ZN(n24166) );
  XNOR2_X1 U32759 ( .A(n24166), .B(n25372), .ZN(n24167) );
  XNOR2_X1 U32760 ( .A(n24749), .B(n24167), .ZN(n43355) );
  XNOR2_X1 U32761 ( .A(n25778), .B(n43355), .ZN(n24168) );
  XNOR2_X1 U32762 ( .A(n24168), .B(n25708), .ZN(n24169) );
  XNOR2_X1 U32763 ( .A(n24170), .B(n24169), .ZN(n24173) );
  XNOR2_X1 U32764 ( .A(n24171), .B(n25882), .ZN(n24172) );
  XNOR2_X1 U32765 ( .A(n24173), .B(n24172), .ZN(n24174) );
  XNOR2_X1 U32766 ( .A(n24175), .B(n24174), .ZN(n29923) );
  AND2_X1 U32767 ( .A1(n24265), .A2(n738), .ZN(n29917) );
  NAND2_X1 U32768 ( .A1(n24191), .A2(n24187), .ZN(n24176) );
  AND2_X1 U32769 ( .A1(n24177), .A2(n24176), .ZN(n24178) );
  NAND2_X1 U32770 ( .A1(n24179), .A2(n24183), .ZN(n24197) );
  OAI21_X1 U32771 ( .B1(n24188), .B2(n24187), .A(n24180), .ZN(n24181) );
  OAI21_X1 U32772 ( .B1(n24182), .B2(n24187), .A(n24181), .ZN(n24184) );
  NAND3_X1 U32773 ( .A1(n24189), .A2(n24188), .A3(n24187), .ZN(n24194) );
  NAND3_X1 U32774 ( .A1(n24192), .A2(n24191), .A3(n24190), .ZN(n24193) );
  NAND3_X1 U32775 ( .A1(n24197), .A2(n24196), .A3(n24195), .ZN(n24198) );
  XNOR2_X2 U32776 ( .A(n25937), .B(n25682), .ZN(n25806) );
  XNOR2_X1 U32777 ( .A(n24716), .B(n25806), .ZN(n25141) );
  INV_X1 U32778 ( .A(n25141), .ZN(n27335) );
  XNOR2_X1 U32779 ( .A(n24200), .B(n2608), .ZN(n24201) );
  XNOR2_X1 U32780 ( .A(n36737), .B(n4637), .ZN(n39720) );
  XNOR2_X1 U32781 ( .A(n24201), .B(n39720), .ZN(n24203) );
  INV_X1 U32782 ( .A(n43020), .ZN(n24202) );
  XNOR2_X1 U32783 ( .A(n24203), .B(n24202), .ZN(n24204) );
  XNOR2_X1 U32784 ( .A(n51751), .B(n24204), .ZN(n24215) );
  NAND3_X1 U32785 ( .A1(n24206), .A2(n24205), .A3(n24211), .ZN(n24210) );
  NAND3_X1 U32786 ( .A1(n24208), .A2(n24211), .A3(n24207), .ZN(n24209) );
  OAI211_X1 U32787 ( .C1(n24212), .C2(n24211), .A(n24210), .B(n24209), .ZN(
        n24214) );
  XNOR2_X1 U32788 ( .A(n25805), .B(n24216), .ZN(n24217) );
  XNOR2_X1 U32789 ( .A(n27335), .B(n24217), .ZN(n24221) );
  XNOR2_X1 U32792 ( .A(n24221), .B(n24220), .ZN(n24226) );
  XNOR2_X1 U32793 ( .A(n26565), .B(n4501), .ZN(n24222) );
  XNOR2_X1 U32794 ( .A(n51380), .B(n24222), .ZN(n24421) );
  INV_X1 U32795 ( .A(n42816), .ZN(n24223) );
  XNOR2_X1 U32796 ( .A(n25935), .B(n24224), .ZN(n27339) );
  XNOR2_X1 U32797 ( .A(n24421), .B(n27339), .ZN(n24225) );
  XNOR2_X1 U32798 ( .A(n25124), .B(n26152), .ZN(n24233) );
  XNOR2_X1 U32799 ( .A(n24227), .B(n4752), .ZN(n24228) );
  XNOR2_X1 U32800 ( .A(n28413), .B(n24228), .ZN(n43805) );
  XNOR2_X1 U32801 ( .A(n24229), .B(n4639), .ZN(n24892) );
  XNOR2_X1 U32802 ( .A(n842), .B(n4665), .ZN(n24230) );
  XNOR2_X1 U32803 ( .A(n24892), .B(n24230), .ZN(n45422) );
  XNOR2_X1 U32804 ( .A(n43805), .B(n45422), .ZN(n24231) );
  XNOR2_X1 U32805 ( .A(n27224), .B(n24231), .ZN(n24232) );
  XNOR2_X1 U32806 ( .A(n24233), .B(n24232), .ZN(n24234) );
  XNOR2_X1 U32807 ( .A(n51056), .B(n24234), .ZN(n24236) );
  XNOR2_X1 U32808 ( .A(n24236), .B(n24235), .ZN(n24262) );
  NAND2_X1 U32809 ( .A1(n24249), .A2(n24244), .ZN(n24252) );
  XNOR2_X1 U32810 ( .A(n26375), .B(n26544), .ZN(n24260) );
  NAND3_X1 U32811 ( .A1(n24256), .A2(n24255), .A3(n24254), .ZN(n24257) );
  XNOR2_X1 U32813 ( .A(n26547), .B(n24260), .ZN(n24261) );
  XNOR2_X1 U32814 ( .A(n24261), .B(n27235), .ZN(n28409) );
  XNOR2_X1 U32815 ( .A(n24262), .B(n28409), .ZN(n24264) );
  INV_X1 U32816 ( .A(n27372), .ZN(n26384) );
  XNOR2_X1 U32817 ( .A(n24264), .B(n26384), .ZN(n24351) );
  INV_X1 U32818 ( .A(n24351), .ZN(n29924) );
  AND2_X1 U32819 ( .A1(n24265), .A2(n29923), .ZN(n24348) );
  AND2_X1 U32820 ( .A1(n27558), .A2(n24351), .ZN(n29916) );
  INV_X1 U32821 ( .A(n24269), .ZN(n24270) );
  XNOR2_X1 U32822 ( .A(n45380), .B(n45253), .ZN(n24273) );
  XNOR2_X1 U32823 ( .A(n25320), .B(n24273), .ZN(n24274) );
  XNOR2_X1 U32824 ( .A(n26093), .B(n24274), .ZN(n24275) );
  XNOR2_X1 U32825 ( .A(n28104), .B(n4121), .ZN(n25319) );
  XNOR2_X1 U32826 ( .A(n25319), .B(n25215), .ZN(n25153) );
  XNOR2_X1 U32827 ( .A(n26395), .B(n42740), .ZN(n24442) );
  NAND2_X1 U32828 ( .A1(n24284), .A2(n24283), .ZN(n24300) );
  INV_X1 U32829 ( .A(n24285), .ZN(n24286) );
  OAI21_X1 U32830 ( .B1(n24288), .B2(n24287), .A(n24286), .ZN(n24299) );
  NAND2_X1 U32831 ( .A1(n24293), .A2(n24292), .ZN(n24294) );
  INV_X1 U32832 ( .A(n24297), .ZN(n24298) );
  NAND4_X2 U32833 ( .A1(n24298), .A2(n24301), .A3(n24300), .A4(n24299), .ZN(
        n26508) );
  XNOR2_X1 U32834 ( .A(n24442), .B(n749), .ZN(n24305) );
  XNOR2_X1 U32835 ( .A(n28424), .B(n28430), .ZN(n24303) );
  XNOR2_X1 U32836 ( .A(n24305), .B(n24304), .ZN(n24307) );
  XNOR2_X1 U32837 ( .A(n24307), .B(n24306), .ZN(n24308) );
  XNOR2_X1 U32838 ( .A(n24548), .B(n26530), .ZN(n24309) );
  XNOR2_X1 U32839 ( .A(n26221), .B(n24309), .ZN(n24312) );
  INV_X1 U32840 ( .A(n24310), .ZN(n24311) );
  XNOR2_X1 U32841 ( .A(n24312), .B(n24311), .ZN(n24322) );
  XNOR2_X1 U32842 ( .A(n24313), .B(n43850), .ZN(n41663) );
  XNOR2_X1 U32843 ( .A(n24314), .B(n4537), .ZN(n24316) );
  XNOR2_X1 U32844 ( .A(n24316), .B(n24315), .ZN(n43304) );
  XNOR2_X1 U32845 ( .A(n41663), .B(n43304), .ZN(n24317) );
  XNOR2_X1 U32846 ( .A(n24318), .B(n26119), .ZN(n24320) );
  XNOR2_X1 U32847 ( .A(n24319), .B(n24320), .ZN(n24321) );
  XNOR2_X1 U32848 ( .A(n24322), .B(n24321), .ZN(n24347) );
  INV_X1 U32849 ( .A(n27501), .ZN(n24323) );
  XNOR2_X1 U32850 ( .A(n26053), .B(n24323), .ZN(n24345) );
  INV_X1 U32851 ( .A(n24324), .ZN(n24337) );
  NAND2_X1 U32852 ( .A1(n24337), .A2(n24336), .ZN(n24325) );
  NAND2_X1 U32853 ( .A1(n24326), .A2(n24325), .ZN(n24327) );
  AND2_X1 U32854 ( .A1(n24328), .A2(n24327), .ZN(n24343) );
  OAI21_X1 U32855 ( .B1(n24331), .B2(n24330), .A(n24329), .ZN(n24342) );
  NOR2_X1 U32856 ( .A1(n24337), .A2(n24336), .ZN(n24339) );
  OAI21_X1 U32857 ( .B1(n24339), .B2(n24338), .A(n3816), .ZN(n24340) );
  XNOR2_X1 U32858 ( .A(n2212), .B(n24345), .ZN(n25833) );
  XNOR2_X1 U32859 ( .A(n25833), .B(n27509), .ZN(n24346) );
  XNOR2_X1 U32860 ( .A(n24347), .B(n24346), .ZN(n30769) );
  INV_X1 U32861 ( .A(n24348), .ZN(n30751) );
  NAND2_X1 U32862 ( .A1(n24349), .A2(n30751), .ZN(n26928) );
  AOI22_X1 U32864 ( .A1(n24352), .A2(n26842), .B1(n51696), .B2(n730), .ZN(
        n24353) );
  NAND2_X1 U32865 ( .A1(n31241), .A2(n31244), .ZN(n24359) );
  NAND2_X1 U32866 ( .A1(n32243), .A2(n31781), .ZN(n24357) );
  OAI22_X1 U32868 ( .A1(n24357), .A2(n32247), .B1(n29364), .B2(n622), .ZN(
        n24358) );
  AOI21_X1 U32869 ( .B1(n30839), .B2(n24359), .A(n24358), .ZN(n24368) );
  INV_X1 U32870 ( .A(n24360), .ZN(n24364) );
  OAI211_X1 U32871 ( .C1(n24364), .C2(n24363), .A(n24362), .B(n24361), .ZN(
        n32230) );
  INV_X1 U32872 ( .A(n32236), .ZN(n24366) );
  XNOR2_X1 U32873 ( .A(n27250), .B(n25003), .ZN(n26592) );
  XNOR2_X1 U32875 ( .A(n26592), .B(n26581), .ZN(n24371) );
  XNOR2_X1 U32876 ( .A(n25755), .B(n43105), .ZN(n24369) );
  XNOR2_X1 U32877 ( .A(n24369), .B(n28214), .ZN(n25865) );
  INV_X1 U32878 ( .A(n25865), .ZN(n24370) );
  XNOR2_X1 U32879 ( .A(n24371), .B(n24370), .ZN(n24372) );
  XNOR2_X1 U32880 ( .A(n28218), .B(n24372), .ZN(n26174) );
  INV_X1 U32881 ( .A(n26174), .ZN(n24382) );
  XNOR2_X1 U32882 ( .A(n51483), .B(n24373), .ZN(n24378) );
  XNOR2_X1 U32883 ( .A(n25353), .B(n27241), .ZN(n26591) );
  INV_X1 U32884 ( .A(n41782), .ZN(n28731) );
  INV_X1 U32885 ( .A(n43314), .ZN(n24374) );
  XNOR2_X1 U32886 ( .A(n28731), .B(n24374), .ZN(n24375) );
  XNOR2_X1 U32887 ( .A(n28213), .B(n24375), .ZN(n24376) );
  XNOR2_X1 U32888 ( .A(n26591), .B(n24376), .ZN(n24377) );
  XNOR2_X1 U32889 ( .A(n24378), .B(n24377), .ZN(n24380) );
  XNOR2_X1 U32890 ( .A(n26435), .B(n27295), .ZN(n25268) );
  XNOR2_X1 U32891 ( .A(n26589), .B(n5016), .ZN(n24379) );
  XNOR2_X1 U32892 ( .A(n25268), .B(n24379), .ZN(n24762) );
  XNOR2_X1 U32893 ( .A(n24762), .B(n24380), .ZN(n24381) );
  INV_X1 U32894 ( .A(n24451), .ZN(n27576) );
  INV_X1 U32895 ( .A(n41961), .ZN(n24385) );
  XNOR2_X1 U32896 ( .A(n24384), .B(n24383), .ZN(n43251) );
  XNOR2_X1 U32897 ( .A(n24385), .B(n43251), .ZN(n24386) );
  XNOR2_X1 U32898 ( .A(n25775), .B(n24386), .ZN(n24387) );
  XNOR2_X1 U32899 ( .A(n24387), .B(n28353), .ZN(n24388) );
  XNOR2_X1 U32900 ( .A(n26611), .B(n25481), .ZN(n24747) );
  XNOR2_X1 U32901 ( .A(n24388), .B(n24747), .ZN(n24391) );
  XNOR2_X1 U32902 ( .A(n25889), .B(n24795), .ZN(n24389) );
  XNOR2_X1 U32903 ( .A(n24390), .B(n24389), .ZN(n28080) );
  XNOR2_X1 U32904 ( .A(n24391), .B(n28080), .ZN(n24393) );
  XNOR2_X1 U32905 ( .A(n24393), .B(n24392), .ZN(n24395) );
  XNOR2_X1 U32906 ( .A(n28242), .B(n51750), .ZN(n26192) );
  INV_X1 U32907 ( .A(n26192), .ZN(n24394) );
  XNOR2_X1 U32908 ( .A(n24394), .B(n24395), .ZN(n26823) );
  XNOR2_X1 U32910 ( .A(n33635), .B(n4451), .ZN(n25938) );
  XNOR2_X1 U32911 ( .A(n24396), .B(n25938), .ZN(n45442) );
  XNOR2_X1 U32912 ( .A(n45442), .B(n4431), .ZN(n24398) );
  XNOR2_X1 U32913 ( .A(n24398), .B(n24397), .ZN(n24399) );
  XNOR2_X1 U32914 ( .A(n28257), .B(n24849), .ZN(n24401) );
  INV_X1 U32915 ( .A(n25346), .ZN(n24400) );
  XNOR2_X1 U32916 ( .A(n24401), .B(n24400), .ZN(n24516) );
  INV_X1 U32917 ( .A(n24516), .ZN(n24402) );
  XNOR2_X1 U32918 ( .A(n26008), .B(n24405), .ZN(n26130) );
  XNOR2_X1 U32919 ( .A(n24406), .B(n26130), .ZN(n24425) );
  NOR2_X1 U32920 ( .A1(n24410), .A2(n24409), .ZN(n24418) );
  XNOR2_X1 U32921 ( .A(n24411), .B(n24412), .ZN(n24415) );
  AOI21_X1 U32922 ( .B1(n24415), .B2(n24414), .A(n24413), .ZN(n24417) );
  XNOR2_X1 U32923 ( .A(n28371), .B(n24593), .ZN(n24423) );
  INV_X1 U32924 ( .A(n24421), .ZN(n24422) );
  XNOR2_X1 U32925 ( .A(n24422), .B(n24423), .ZN(n24424) );
  XNOR2_X1 U32926 ( .A(n25249), .B(n27374), .ZN(n24519) );
  XNOR2_X1 U32927 ( .A(n51647), .B(n27224), .ZN(n24426) );
  XNOR2_X1 U32928 ( .A(n24519), .B(n24426), .ZN(n24427) );
  XNOR2_X1 U32929 ( .A(n28040), .B(n25996), .ZN(n24912) );
  XNOR2_X1 U32930 ( .A(n24912), .B(n24427), .ZN(n24428) );
  XNOR2_X1 U32931 ( .A(n26155), .B(n24428), .ZN(n24441) );
  INV_X1 U32932 ( .A(n24429), .ZN(n42773) );
  XNOR2_X1 U32933 ( .A(n4325), .B(n4752), .ZN(n42831) );
  XNOR2_X1 U32934 ( .A(n42831), .B(n4035), .ZN(n24431) );
  XNOR2_X1 U32935 ( .A(n24431), .B(n24430), .ZN(n24432) );
  XNOR2_X1 U32936 ( .A(n42773), .B(n24432), .ZN(n24433) );
  XNOR2_X1 U32937 ( .A(n24891), .B(n24433), .ZN(n24434) );
  XNOR2_X1 U32938 ( .A(n24434), .B(n26304), .ZN(n24435) );
  INV_X1 U32939 ( .A(n24830), .ZN(n42283) );
  XNOR2_X1 U32940 ( .A(n25308), .B(n42283), .ZN(n24436) );
  XNOR2_X1 U32941 ( .A(n24905), .B(n24436), .ZN(n26555) );
  INV_X1 U32942 ( .A(n26555), .ZN(n24437) );
  XNOR2_X1 U32943 ( .A(n24438), .B(n24437), .ZN(n24439) );
  NAND2_X1 U32944 ( .A1(n1484), .A2(n26772), .ZN(n27680) );
  OR2_X1 U32945 ( .A1(n27580), .A2(n27680), .ZN(n26825) );
  XNOR2_X1 U32946 ( .A(n368), .B(n24442), .ZN(n24447) );
  XNOR2_X1 U32947 ( .A(n43552), .B(n25925), .ZN(n43675) );
  XNOR2_X1 U32948 ( .A(n24443), .B(n3014), .ZN(n42741) );
  XNOR2_X1 U32949 ( .A(n43675), .B(n42741), .ZN(n24444) );
  XNOR2_X1 U32950 ( .A(n26100), .B(n24444), .ZN(n24445) );
  XNOR2_X1 U32951 ( .A(n24445), .B(n25215), .ZN(n24446) );
  XNOR2_X1 U32952 ( .A(n24447), .B(n24446), .ZN(n24450) );
  XNOR2_X1 U32953 ( .A(n26093), .B(n25929), .ZN(n26214) );
  XNOR2_X1 U32954 ( .A(n28431), .B(n2164), .ZN(n24448) );
  XNOR2_X1 U32955 ( .A(n24448), .B(n26214), .ZN(n24449) );
  XNOR2_X1 U32956 ( .A(n25920), .B(n25429), .ZN(n25737) );
  NOR2_X1 U32957 ( .A1(n27685), .A2(n27690), .ZN(n26962) );
  BUF_X2 U32958 ( .A(n24451), .Z(n26955) );
  INV_X1 U32959 ( .A(n26823), .ZN(n26960) );
  AND2_X1 U32960 ( .A1(n26955), .A2(n26960), .ZN(n27679) );
  NAND2_X1 U32961 ( .A1(n26962), .A2(n27679), .ZN(n24470) );
  INV_X1 U32962 ( .A(n4177), .ZN(n49387) );
  OAI211_X1 U32963 ( .C1(n4177), .C2(n24455), .A(n24454), .B(n24453), .ZN(
        n24456) );
  XNOR2_X1 U32964 ( .A(n24554), .B(n25901), .ZN(n24457) );
  XNOR2_X1 U32965 ( .A(n24458), .B(n24457), .ZN(n43234) );
  XNOR2_X1 U32966 ( .A(n24459), .B(n34265), .ZN(n42029) );
  XNOR2_X1 U32967 ( .A(n43234), .B(n42029), .ZN(n24460) );
  XNOR2_X1 U32968 ( .A(n25540), .B(n24460), .ZN(n24461) );
  XNOR2_X1 U32969 ( .A(n24463), .B(n24462), .ZN(n24465) );
  XNOR2_X1 U32970 ( .A(n24736), .B(n4645), .ZN(n25154) );
  XNOR2_X1 U32971 ( .A(n26125), .B(n471), .ZN(n24466) );
  NAND3_X1 U32972 ( .A1(n27679), .A2(n24467), .A3(n26771), .ZN(n24469) );
  AND4_X1 U32973 ( .A1(n26825), .A2(n24470), .A3(n24469), .A4(n24468), .ZN(
        n24478) );
  AND3_X1 U32974 ( .A1(n27680), .A2(n6290), .A3(n26960), .ZN(n24473) );
  INV_X1 U32975 ( .A(n27677), .ZN(n24471) );
  OAI21_X1 U32976 ( .B1(n24471), .B2(n27576), .A(n8481), .ZN(n24472) );
  AOI22_X1 U32977 ( .A1(n26810), .A2(n24473), .B1(n24472), .B2(n27686), .ZN(
        n24477) );
  NAND2_X1 U32978 ( .A1(n26955), .A2(n26823), .ZN(n26774) );
  NAND2_X1 U32979 ( .A1(n27681), .A2(n1484), .ZN(n24474) );
  NOR2_X1 U32980 ( .A1(n26774), .A2(n24474), .ZN(n26776) );
  NAND2_X1 U32981 ( .A1(n27677), .A2(n27576), .ZN(n27581) );
  OAI211_X1 U32982 ( .C1(n26776), .C2(n27578), .A(n6290), .B(n27581), .ZN(
        n24476) );
  NAND2_X1 U32983 ( .A1(n26819), .A2(n26814), .ZN(n24475) );
  XNOR2_X1 U32984 ( .A(n24945), .B(n27290), .ZN(n25002) );
  INV_X1 U32985 ( .A(n25002), .ZN(n25267) );
  XNOR2_X1 U32986 ( .A(n27289), .B(n25267), .ZN(n25768) );
  INV_X1 U32987 ( .A(n25768), .ZN(n24491) );
  XNOR2_X1 U32988 ( .A(n41949), .B(n24479), .ZN(n24480) );
  XNOR2_X1 U32989 ( .A(n24480), .B(n43267), .ZN(n24481) );
  XNOR2_X1 U32990 ( .A(n24810), .B(n24481), .ZN(n24483) );
  INV_X1 U32991 ( .A(n26159), .ZN(n24482) );
  XNOR2_X1 U32992 ( .A(n24483), .B(n24482), .ZN(n24487) );
  XNOR2_X1 U32993 ( .A(n24484), .B(n4687), .ZN(n44070) );
  XNOR2_X1 U32994 ( .A(n25506), .B(n44070), .ZN(n24991) );
  INV_X1 U32995 ( .A(n24991), .ZN(n24485) );
  XNOR2_X1 U32996 ( .A(n24485), .B(n24651), .ZN(n24486) );
  INV_X1 U32998 ( .A(n24563), .ZN(n26779) );
  INV_X1 U32999 ( .A(n24791), .ZN(n24492) );
  XNOR2_X1 U33000 ( .A(n750), .B(n24492), .ZN(n24493) );
  XNOR2_X1 U33001 ( .A(n25483), .B(n51720), .ZN(n26187) );
  XNOR2_X1 U33002 ( .A(n24493), .B(n26187), .ZN(n24623) );
  XNOR2_X1 U33003 ( .A(n24494), .B(n24623), .ZN(n24504) );
  XNOR2_X1 U33004 ( .A(n24495), .B(n4712), .ZN(n46148) );
  XNOR2_X1 U33005 ( .A(n46148), .B(n46144), .ZN(n24497) );
  XNOR2_X1 U33006 ( .A(n24496), .B(n28071), .ZN(n44367) );
  XNOR2_X1 U33007 ( .A(n24497), .B(n44367), .ZN(n24498) );
  XNOR2_X1 U33008 ( .A(n26264), .B(n24498), .ZN(n24499) );
  XNOR2_X1 U33009 ( .A(n26611), .B(n24499), .ZN(n24501) );
  XNOR2_X1 U33010 ( .A(n25481), .B(n25775), .ZN(n24500) );
  XNOR2_X1 U33011 ( .A(n24501), .B(n24500), .ZN(n24502) );
  XNOR2_X1 U33012 ( .A(n28364), .B(n24502), .ZN(n24503) );
  XNOR2_X1 U33013 ( .A(n26013), .B(n25554), .ZN(n25699) );
  INV_X1 U33014 ( .A(n25681), .ZN(n24916) );
  INV_X1 U33015 ( .A(n35654), .ZN(n24507) );
  XNOR2_X1 U33016 ( .A(n45105), .B(n24505), .ZN(n42780) );
  XNOR2_X1 U33017 ( .A(n4579), .B(n2112), .ZN(n44043) );
  XNOR2_X1 U33018 ( .A(n2608), .B(n44043), .ZN(n26131) );
  XNOR2_X1 U33019 ( .A(n42780), .B(n26131), .ZN(n24506) );
  XNOR2_X1 U33020 ( .A(n24507), .B(n24506), .ZN(n24508) );
  XNOR2_X1 U33021 ( .A(n51423), .B(n24508), .ZN(n24509) );
  XNOR2_X1 U33022 ( .A(n24509), .B(n28048), .ZN(n24510) );
  XNOR2_X1 U33023 ( .A(n24916), .B(n24510), .ZN(n24513) );
  XNOR2_X1 U33025 ( .A(n24513), .B(n24512), .ZN(n24517) );
  XNOR2_X1 U33026 ( .A(n24514), .B(n28383), .ZN(n24515) );
  INV_X1 U33027 ( .A(n25724), .ZN(n24518) );
  XNOR2_X1 U33028 ( .A(n26147), .B(n24518), .ZN(n24579) );
  XNOR2_X1 U33029 ( .A(n24519), .B(n24579), .ZN(n24529) );
  INV_X1 U33030 ( .A(n34891), .ZN(n24520) );
  XNOR2_X1 U33031 ( .A(n24521), .B(n24520), .ZN(n45125) );
  XNOR2_X1 U33032 ( .A(n25040), .B(n4296), .ZN(n24522) );
  XNOR2_X1 U33033 ( .A(n24582), .B(n24522), .ZN(n42384) );
  XNOR2_X1 U33034 ( .A(n42384), .B(n24523), .ZN(n24524) );
  XNOR2_X1 U33035 ( .A(n45125), .B(n24524), .ZN(n24525) );
  XNOR2_X1 U33036 ( .A(n51647), .B(n24525), .ZN(n24527) );
  XNOR2_X1 U33037 ( .A(n24527), .B(n24526), .ZN(n24528) );
  XNOR2_X1 U33038 ( .A(n24529), .B(n24528), .ZN(n24530) );
  XNOR2_X1 U33039 ( .A(n26100), .B(n28430), .ZN(n24532) );
  XNOR2_X1 U33040 ( .A(n26508), .B(n25920), .ZN(n26094) );
  XNOR2_X1 U33041 ( .A(n24532), .B(n26094), .ZN(n24533) );
  XNOR2_X1 U33042 ( .A(n28103), .B(n4932), .ZN(n24534) );
  XNOR2_X1 U33043 ( .A(n24534), .B(n28431), .ZN(n24535) );
  XNOR2_X1 U33044 ( .A(n24535), .B(n51502), .ZN(n26516) );
  XNOR2_X1 U33045 ( .A(n24536), .B(n26516), .ZN(n24547) );
  XNOR2_X1 U33046 ( .A(n28106), .B(n26390), .ZN(n24542) );
  XNOR2_X1 U33047 ( .A(n42339), .B(n42342), .ZN(n24539) );
  XNOR2_X1 U33048 ( .A(n24537), .B(n4746), .ZN(n24538) );
  XNOR2_X1 U33049 ( .A(n24538), .B(n24725), .ZN(n45039) );
  XNOR2_X1 U33050 ( .A(n24539), .B(n45039), .ZN(n24540) );
  XNOR2_X1 U33051 ( .A(n25740), .B(n24540), .ZN(n24541) );
  XNOR2_X1 U33052 ( .A(n24542), .B(n24541), .ZN(n24543) );
  XNOR2_X1 U33053 ( .A(n28302), .B(n24543), .ZN(n24544) );
  XNOR2_X1 U33054 ( .A(n24545), .B(n24544), .ZN(n24546) );
  XNOR2_X1 U33055 ( .A(n24548), .B(n26531), .ZN(n28400) );
  XNOR2_X1 U33056 ( .A(n28400), .B(n25154), .ZN(n24549) );
  XNOR2_X1 U33057 ( .A(n26536), .B(n26053), .ZN(n24634) );
  XNOR2_X1 U33058 ( .A(n24634), .B(n24549), .ZN(n24560) );
  XNOR2_X1 U33059 ( .A(n25445), .B(n4668), .ZN(n26120) );
  XNOR2_X1 U33060 ( .A(n25897), .B(n41660), .ZN(n24552) );
  INV_X1 U33061 ( .A(n24550), .ZN(n24551) );
  XNOR2_X1 U33062 ( .A(n24552), .B(n24551), .ZN(n44310) );
  XNOR2_X1 U33063 ( .A(n24554), .B(n24553), .ZN(n46124) );
  XNOR2_X1 U33064 ( .A(n44310), .B(n46124), .ZN(n24555) );
  XNOR2_X1 U33065 ( .A(n24556), .B(n24555), .ZN(n24557) );
  XNOR2_X1 U33066 ( .A(n26120), .B(n24557), .ZN(n24558) );
  XNOR2_X1 U33067 ( .A(n24631), .B(n24558), .ZN(n24559) );
  AND2_X1 U33068 ( .A1(n27764), .A2(n27765), .ZN(n29469) );
  NAND2_X1 U33069 ( .A1(n27015), .A2(n29469), .ZN(n24561) );
  INV_X1 U33070 ( .A(n26690), .ZN(n24568) );
  INV_X1 U33071 ( .A(n29467), .ZN(n26788) );
  OR2_X1 U33072 ( .A1(n24563), .A2(n26788), .ZN(n27012) );
  INV_X1 U33073 ( .A(n27012), .ZN(n24562) );
  INV_X1 U33074 ( .A(n27764), .ZN(n26781) );
  AND2_X1 U33075 ( .A1(n26781), .A2(n29467), .ZN(n27007) );
  INV_X1 U33076 ( .A(n27765), .ZN(n29463) );
  NAND3_X1 U33077 ( .A1(n29471), .A2(n27764), .A3(n27758), .ZN(n24566) );
  NAND2_X1 U33078 ( .A1(n26788), .A2(n27764), .ZN(n24564) );
  OAI211_X1 U33079 ( .C1(n27007), .C2(n27758), .A(n7973), .B(n24564), .ZN(
        n24565) );
  OR2_X1 U33080 ( .A1(n737), .A2(n2144), .ZN(n26803) );
  AOI22_X1 U33082 ( .A1(n27621), .A2(n27632), .B1(n27730), .B2(n22344), .ZN(
        n24575) );
  OAI211_X1 U33083 ( .C1(n26890), .C2(n27623), .A(n24571), .B(n27720), .ZN(
        n24574) );
  NAND2_X1 U33084 ( .A1(n27635), .A2(n597), .ZN(n26887) );
  NOR2_X1 U33087 ( .A1(n29650), .A2(n30824), .ZN(n24782) );
  XNOR2_X1 U33088 ( .A(n51646), .B(n26152), .ZN(n24900) );
  XNOR2_X1 U33089 ( .A(n24577), .B(n24900), .ZN(n26294) );
  XNOR2_X1 U33090 ( .A(n24905), .B(n25308), .ZN(n28035) );
  XNOR2_X1 U33091 ( .A(n24579), .B(n28035), .ZN(n24590) );
  INV_X1 U33092 ( .A(n24891), .ZN(n24580) );
  XNOR2_X1 U33093 ( .A(n26540), .B(n24580), .ZN(n24837) );
  INV_X1 U33094 ( .A(n24581), .ZN(n24583) );
  XNOR2_X1 U33095 ( .A(n24583), .B(n24582), .ZN(n42275) );
  XNOR2_X1 U33096 ( .A(n4706), .B(n4578), .ZN(n24584) );
  XNOR2_X1 U33097 ( .A(n24585), .B(n24584), .ZN(n44537) );
  XNOR2_X1 U33098 ( .A(n42275), .B(n44537), .ZN(n24586) );
  XNOR2_X1 U33099 ( .A(n25047), .B(n24586), .ZN(n24587) );
  XNOR2_X1 U33100 ( .A(n24587), .B(n26544), .ZN(n24588) );
  XNOR2_X1 U33101 ( .A(n24588), .B(n24837), .ZN(n24589) );
  XNOR2_X1 U33102 ( .A(n24590), .B(n24589), .ZN(n24591) );
  XNOR2_X1 U33103 ( .A(n25554), .B(n28048), .ZN(n24592) );
  XNOR2_X1 U33104 ( .A(n25816), .B(n24592), .ZN(n24594) );
  XNOR2_X1 U33105 ( .A(n24594), .B(n24593), .ZN(n24596) );
  INV_X1 U33106 ( .A(n25035), .ZN(n24595) );
  XNOR2_X1 U33107 ( .A(n24595), .B(n24596), .ZN(n24607) );
  XNOR2_X1 U33108 ( .A(n51119), .B(n26272), .ZN(n24605) );
  XNOR2_X1 U33109 ( .A(n4423), .B(n4343), .ZN(n24597) );
  XNOR2_X1 U33110 ( .A(n35108), .B(n24597), .ZN(n43744) );
  XNOR2_X1 U33111 ( .A(n2608), .B(n4940), .ZN(n24598) );
  XNOR2_X1 U33112 ( .A(n43744), .B(n24598), .ZN(n24599) );
  XNOR2_X1 U33113 ( .A(n42419), .B(n24599), .ZN(n24600) );
  XNOR2_X1 U33114 ( .A(n24600), .B(n42780), .ZN(n24601) );
  XNOR2_X1 U33115 ( .A(n25813), .B(n24601), .ZN(n24602) );
  XNOR2_X1 U33116 ( .A(n24602), .B(n25947), .ZN(n24603) );
  XNOR2_X1 U33117 ( .A(n25937), .B(n24849), .ZN(n26572) );
  XNOR2_X1 U33118 ( .A(n24603), .B(n26572), .ZN(n24604) );
  XNOR2_X1 U33119 ( .A(n24605), .B(n24604), .ZN(n24606) );
  XNOR2_X1 U33120 ( .A(n27479), .B(n27473), .ZN(n24609) );
  XNOR2_X1 U33121 ( .A(n24608), .B(n24609), .ZN(n24803) );
  XNOR2_X1 U33122 ( .A(n25889), .B(n24757), .ZN(n24618) );
  XNOR2_X1 U33123 ( .A(n26259), .B(n24610), .ZN(n39538) );
  XNOR2_X1 U33124 ( .A(n4667), .B(n4782), .ZN(n24611) );
  XNOR2_X1 U33125 ( .A(n24612), .B(n24611), .ZN(n43040) );
  XNOR2_X1 U33126 ( .A(n42327), .B(n4836), .ZN(n24613) );
  XNOR2_X1 U33127 ( .A(n43040), .B(n24613), .ZN(n24614) );
  XNOR2_X1 U33128 ( .A(n39538), .B(n24614), .ZN(n24615) );
  XNOR2_X1 U33129 ( .A(n24616), .B(n24615), .ZN(n24617) );
  XNOR2_X1 U33130 ( .A(n24618), .B(n24617), .ZN(n24621) );
  XNOR2_X1 U33131 ( .A(n51750), .B(n24619), .ZN(n24620) );
  XNOR2_X1 U33132 ( .A(n24621), .B(n24620), .ZN(n24622) );
  XNOR2_X1 U33133 ( .A(n24623), .B(n24622), .ZN(n24624) );
  NAND2_X1 U33135 ( .A1(n26731), .A2(n51679), .ZN(n26733) );
  INV_X1 U33136 ( .A(n24625), .ZN(n24627) );
  XNOR2_X1 U33137 ( .A(n24627), .B(n24626), .ZN(n43032) );
  XNOR2_X1 U33138 ( .A(n26526), .B(n4879), .ZN(n36291) );
  XNOR2_X1 U33139 ( .A(n43849), .B(n2603), .ZN(n36966) );
  XNOR2_X1 U33140 ( .A(n36291), .B(n36966), .ZN(n24628) );
  XNOR2_X1 U33141 ( .A(n43032), .B(n24628), .ZN(n24629) );
  XNOR2_X1 U33142 ( .A(n24631), .B(n24632), .ZN(n24633) );
  XNOR2_X1 U33143 ( .A(n24634), .B(n24633), .ZN(n24635) );
  XNOR2_X1 U33144 ( .A(n24872), .B(n25450), .ZN(n27511) );
  XNOR2_X1 U33145 ( .A(n27511), .B(n24635), .ZN(n26998) );
  XNOR2_X1 U33146 ( .A(n25429), .B(n27177), .ZN(n24732) );
  XNOR2_X1 U33147 ( .A(n26210), .B(n26390), .ZN(n24636) );
  XNOR2_X1 U33148 ( .A(n28106), .B(n24636), .ZN(n26047) );
  XNOR2_X1 U33149 ( .A(n24637), .B(n26047), .ZN(n24646) );
  XNOR2_X1 U33150 ( .A(n24639), .B(n24638), .ZN(n44508) );
  XNOR2_X1 U33151 ( .A(n24641), .B(n24640), .ZN(n42214) );
  XNOR2_X1 U33152 ( .A(n44508), .B(n42214), .ZN(n24642) );
  XNOR2_X1 U33153 ( .A(n26508), .B(n24642), .ZN(n24643) );
  XNOR2_X1 U33154 ( .A(n751), .B(n24643), .ZN(n24644) );
  XNOR2_X1 U33155 ( .A(n24646), .B(n24645), .ZN(n24648) );
  XNOR2_X1 U33156 ( .A(n27384), .B(n27445), .ZN(n25087) );
  XNOR2_X1 U33157 ( .A(n25087), .B(n28438), .ZN(n26218) );
  INV_X1 U33158 ( .A(n26218), .ZN(n24647) );
  AND2_X1 U33159 ( .A1(n26998), .A2(n27711), .ZN(n26991) );
  AND2_X1 U33160 ( .A1(n24649), .A2(n24675), .ZN(n24673) );
  INV_X1 U33161 ( .A(n24673), .ZN(n29419) );
  NAND2_X1 U33162 ( .A1(n26991), .A2(n29419), .ZN(n29407) );
  NOR2_X1 U33163 ( .A1(n27709), .A2(n24673), .ZN(n26734) );
  INV_X1 U33164 ( .A(n25353), .ZN(n24650) );
  XNOR2_X1 U33165 ( .A(n24651), .B(n24650), .ZN(n24653) );
  INV_X1 U33166 ( .A(n27242), .ZN(n24652) );
  XNOR2_X1 U33167 ( .A(n24653), .B(n24652), .ZN(n28096) );
  XNOR2_X1 U33168 ( .A(n28096), .B(n24654), .ZN(n24667) );
  XNOR2_X1 U33169 ( .A(n27309), .B(n24810), .ZN(n24656) );
  XNOR2_X1 U33170 ( .A(n24655), .B(n4585), .ZN(n25351) );
  XNOR2_X1 U33171 ( .A(n24656), .B(n25351), .ZN(n24663) );
  XNOR2_X1 U33172 ( .A(n41949), .B(n33746), .ZN(n24658) );
  INV_X1 U33173 ( .A(n26243), .ZN(n24657) );
  XNOR2_X1 U33174 ( .A(n24658), .B(n24657), .ZN(n40996) );
  XNOR2_X1 U33175 ( .A(n40996), .B(n43586), .ZN(n24659) );
  XNOR2_X1 U33176 ( .A(n25495), .B(n24659), .ZN(n24661) );
  XNOR2_X1 U33177 ( .A(n24661), .B(n24660), .ZN(n24662) );
  XNOR2_X1 U33178 ( .A(n24663), .B(n24662), .ZN(n24665) );
  XNOR2_X1 U33179 ( .A(n2080), .B(n26432), .ZN(n28216) );
  XNOR2_X1 U33180 ( .A(n28216), .B(n27241), .ZN(n26170) );
  INV_X1 U33181 ( .A(n26170), .ZN(n24664) );
  XNOR2_X1 U33182 ( .A(n24665), .B(n24664), .ZN(n24666) );
  NAND2_X1 U33184 ( .A1(n29413), .A2(n51678), .ZN(n29408) );
  OAI21_X1 U33185 ( .B1(n26731), .B2(n26989), .A(n29408), .ZN(n24668) );
  INV_X1 U33186 ( .A(n27709), .ZN(n27707) );
  NAND3_X1 U33187 ( .A1(n27707), .A2(n26985), .A3(n51351), .ZN(n24669) );
  OAI211_X1 U33188 ( .C1(n26733), .C2(n29407), .A(n24670), .B(n24669), .ZN(
        n24671) );
  INV_X1 U33189 ( .A(n24671), .ZN(n24677) );
  INV_X1 U33190 ( .A(n26998), .ZN(n29418) );
  AND2_X1 U33191 ( .A1(n29418), .A2(n7362), .ZN(n26901) );
  AND2_X1 U33192 ( .A1(n26989), .A2(n51679), .ZN(n29426) );
  AND2_X1 U33195 ( .A1(n24649), .A2(n29422), .ZN(n24674) );
  INV_X1 U33196 ( .A(n24674), .ZN(n27710) );
  NAND3_X1 U33197 ( .A1(n29428), .A2(n27706), .A3(n27710), .ZN(n26900) );
  AND2_X1 U33198 ( .A1(n26900), .A2(n24672), .ZN(n24676) );
  OAI211_X1 U33199 ( .C1(n29422), .C2(n26905), .A(n29418), .B(n27711), .ZN(
        n26904) );
  NAND2_X1 U33200 ( .A1(n26991), .A2(n24673), .ZN(n26737) );
  INV_X1 U33201 ( .A(n29408), .ZN(n29411) );
  OAI21_X1 U33202 ( .B1(n26859), .B2(n27600), .A(n26909), .ZN(n24678) );
  NAND2_X1 U33203 ( .A1(n24678), .A2(n27601), .ZN(n24682) );
  INV_X1 U33204 ( .A(n24679), .ZN(n24680) );
  OR2_X1 U33205 ( .A1(n26914), .A2(n24680), .ZN(n26853) );
  INV_X1 U33206 ( .A(n26856), .ZN(n30658) );
  NAND2_X1 U33207 ( .A1(n30658), .A2(n27608), .ZN(n24681) );
  INV_X1 U33209 ( .A(n26914), .ZN(n26911) );
  INV_X1 U33210 ( .A(n24683), .ZN(n24686) );
  INV_X1 U33211 ( .A(n30664), .ZN(n30676) );
  AOI21_X1 U33212 ( .B1(n26909), .B2(n27609), .A(n27604), .ZN(n24684) );
  OR2_X1 U33213 ( .A1(n24684), .A2(n26855), .ZN(n24685) );
  OAI211_X1 U33214 ( .C1(n24686), .C2(n30676), .A(n24685), .B(n24687), .ZN(
        n24689) );
  NOR2_X1 U33215 ( .A1(n26859), .A2(n30673), .ZN(n26920) );
  NAND2_X1 U33216 ( .A1(n26920), .A2(n27599), .ZN(n24688) );
  NAND4_X2 U33217 ( .A1(n24689), .A2(n24690), .A3(n30678), .A4(n24688), .ZN(
        n31306) );
  XNOR2_X1 U33218 ( .A(n26540), .B(n26544), .ZN(n24699) );
  INV_X1 U33219 ( .A(n24692), .ZN(n26144) );
  XNOR2_X1 U33220 ( .A(n26144), .B(n24828), .ZN(n24693) );
  XNOR2_X1 U33221 ( .A(n24693), .B(n25956), .ZN(n44059) );
  XNOR2_X1 U33222 ( .A(n44059), .B(n4755), .ZN(n24696) );
  XNOR2_X1 U33223 ( .A(n24695), .B(n24694), .ZN(n42520) );
  XNOR2_X1 U33224 ( .A(n24696), .B(n42520), .ZN(n24697) );
  XNOR2_X1 U33225 ( .A(n25249), .B(n24697), .ZN(n24698) );
  XNOR2_X1 U33226 ( .A(n24699), .B(n24698), .ZN(n24701) );
  XNOR2_X1 U33227 ( .A(n24701), .B(n24700), .ZN(n24702) );
  XNOR2_X1 U33228 ( .A(n26548), .B(n51647), .ZN(n26374) );
  XNOR2_X1 U33229 ( .A(n24702), .B(n26374), .ZN(n24703) );
  XNOR2_X1 U33230 ( .A(n25946), .B(n24849), .ZN(n25130) );
  XNOR2_X1 U33231 ( .A(n24705), .B(n25130), .ZN(n24706) );
  XNOR2_X1 U33232 ( .A(n27217), .B(n24706), .ZN(n24720) );
  INV_X1 U33233 ( .A(n24707), .ZN(n24711) );
  INV_X1 U33234 ( .A(n24708), .ZN(n34254) );
  XNOR2_X1 U33235 ( .A(n42816), .B(n4739), .ZN(n43018) );
  XNOR2_X1 U33236 ( .A(n43018), .B(n4883), .ZN(n24709) );
  XNOR2_X1 U33237 ( .A(n34254), .B(n24709), .ZN(n24710) );
  XNOR2_X1 U33238 ( .A(n24711), .B(n24710), .ZN(n24712) );
  XNOR2_X1 U33239 ( .A(n27419), .B(n24712), .ZN(n24714) );
  XNOR2_X1 U33240 ( .A(n28257), .B(n25554), .ZN(n24713) );
  XNOR2_X1 U33241 ( .A(n24714), .B(n24713), .ZN(n24715) );
  XNOR2_X1 U33242 ( .A(n26008), .B(n24715), .ZN(n24718) );
  XNOR2_X1 U33243 ( .A(n24716), .B(n25240), .ZN(n24717) );
  XNOR2_X1 U33244 ( .A(n24717), .B(n25806), .ZN(n26354) );
  XNOR2_X1 U33245 ( .A(n24718), .B(n26354), .ZN(n24719) );
  XNOR2_X1 U33246 ( .A(n24721), .B(n24722), .ZN(n24731) );
  INV_X1 U33247 ( .A(n24723), .ZN(n24724) );
  XNOR2_X1 U33248 ( .A(n24724), .B(n24820), .ZN(n42563) );
  XNOR2_X1 U33249 ( .A(n24725), .B(n48597), .ZN(n44010) );
  XNOR2_X1 U33250 ( .A(n44010), .B(n42349), .ZN(n24726) );
  XNOR2_X1 U33251 ( .A(n42563), .B(n24726), .ZN(n24727) );
  XNOR2_X1 U33252 ( .A(n26044), .B(n24727), .ZN(n24728) );
  XNOR2_X1 U33253 ( .A(n24728), .B(n28431), .ZN(n24729) );
  XNOR2_X1 U33254 ( .A(n26214), .B(n24732), .ZN(n24733) );
  XNOR2_X1 U33255 ( .A(n25084), .B(n24733), .ZN(n24734) );
  XNOR2_X1 U33256 ( .A(n25833), .B(n24735), .ZN(n24746) );
  XNOR2_X1 U33257 ( .A(n24737), .B(n27502), .ZN(n25226) );
  XNOR2_X1 U33258 ( .A(n33611), .B(n34265), .ZN(n24739) );
  XNOR2_X1 U33259 ( .A(n24739), .B(n24738), .ZN(n41865) );
  XNOR2_X1 U33260 ( .A(n43136), .B(n4649), .ZN(n24740) );
  XNOR2_X1 U33261 ( .A(n41865), .B(n24740), .ZN(n24741) );
  XNOR2_X1 U33262 ( .A(n25548), .B(n24741), .ZN(n24742) );
  XNOR2_X1 U33263 ( .A(n25161), .B(n24742), .ZN(n24743) );
  XNOR2_X1 U33264 ( .A(n25226), .B(n24743), .ZN(n24744) );
  INV_X1 U33265 ( .A(n26055), .ZN(n25164) );
  XNOR2_X1 U33266 ( .A(n24744), .B(n25164), .ZN(n24745) );
  NAND2_X1 U33267 ( .A1(n27668), .A2(n26937), .ZN(n27670) );
  XNOR2_X1 U33268 ( .A(n24747), .B(n25608), .ZN(n24753) );
  XNOR2_X1 U33269 ( .A(n24748), .B(n4824), .ZN(n41872) );
  XNOR2_X1 U33270 ( .A(n41872), .B(n4934), .ZN(n24750) );
  XNOR2_X1 U33271 ( .A(n24749), .B(n44495), .ZN(n43109) );
  XNOR2_X1 U33272 ( .A(n24750), .B(n43109), .ZN(n24751) );
  XNOR2_X1 U33273 ( .A(n25176), .B(n24751), .ZN(n24752) );
  XNOR2_X1 U33274 ( .A(n24753), .B(n24752), .ZN(n24755) );
  XNOR2_X1 U33275 ( .A(n26175), .B(n25708), .ZN(n24754) );
  XNOR2_X1 U33276 ( .A(n750), .B(n24754), .ZN(n26452) );
  XNOR2_X1 U33277 ( .A(n24755), .B(n26452), .ZN(n24760) );
  INV_X1 U33278 ( .A(n24756), .ZN(n24758) );
  XNOR2_X1 U33279 ( .A(n24758), .B(n26190), .ZN(n24759) );
  XNOR2_X2 U33280 ( .A(n24759), .B(n24760), .ZN(n26944) );
  NAND2_X1 U33281 ( .A1(n24761), .A2(n26944), .ZN(n24780) );
  XNOR2_X1 U33282 ( .A(n26170), .B(n24762), .ZN(n24764) );
  XNOR2_X1 U33283 ( .A(n24763), .B(n25664), .ZN(n27240) );
  XNOR2_X1 U33284 ( .A(n27257), .B(n27291), .ZN(n26171) );
  XOR2_X1 U33285 ( .A(n4317), .B(n4599), .Z(n24765) );
  XNOR2_X1 U33286 ( .A(n24765), .B(n33474), .ZN(n24766) );
  XNOR2_X1 U33287 ( .A(n24767), .B(n24766), .ZN(n42893) );
  XNOR2_X1 U33288 ( .A(n42889), .B(n4237), .ZN(n34728) );
  XNOR2_X1 U33289 ( .A(n34728), .B(n24992), .ZN(n24768) );
  XNOR2_X1 U33290 ( .A(n24768), .B(n26242), .ZN(n24769) );
  XNOR2_X1 U33291 ( .A(n42893), .B(n24769), .ZN(n24770) );
  XNOR2_X1 U33292 ( .A(n25003), .B(n24770), .ZN(n24771) );
  XNOR2_X1 U33293 ( .A(n25762), .B(n24771), .ZN(n24772) );
  XNOR2_X1 U33294 ( .A(n25005), .B(n24772), .ZN(n24773) );
  NAND2_X1 U33295 ( .A1(n26944), .A2(n447), .ZN(n26949) );
  NOR2_X1 U33296 ( .A1(n26949), .A2(n3765), .ZN(n27066) );
  NOR2_X1 U33297 ( .A1(n27070), .A2(n2642), .ZN(n24775) );
  AOI21_X1 U33298 ( .B1(n27066), .B2(n27665), .A(n24775), .ZN(n24779) );
  OAI21_X1 U33299 ( .B1(n27653), .B2(n27669), .A(n27067), .ZN(n24778) );
  OAI21_X1 U33300 ( .B1(n26743), .B2(n26937), .A(n27669), .ZN(n24777) );
  OAI21_X1 U33301 ( .B1(n31302), .B2(n31306), .A(n30644), .ZN(n29403) );
  NAND2_X1 U33302 ( .A1(n30833), .A2(n30825), .ZN(n24781) );
  AOI22_X1 U33303 ( .A1(n24782), .A2(n29403), .B1(n51085), .B2(n24781), .ZN(
        n24789) );
  INV_X1 U33304 ( .A(n31306), .ZN(n31303) );
  NAND3_X1 U33305 ( .A1(n30830), .A2(n51085), .A3(n30824), .ZN(n24783) );
  AND2_X1 U33306 ( .A1(n24783), .A2(n24784), .ZN(n24788) );
  OAI21_X1 U33307 ( .B1(n30824), .B2(n31302), .A(n30640), .ZN(n24785) );
  NAND3_X1 U33308 ( .A1(n30835), .A2(n24785), .A3(n51085), .ZN(n24787) );
  OR2_X1 U33309 ( .A1(n31306), .A2(n31300), .ZN(n30653) );
  INV_X1 U33310 ( .A(n51085), .ZN(n31294) );
  INV_X1 U33311 ( .A(n31302), .ZN(n30834) );
  NAND2_X1 U33312 ( .A1(n31301), .A2(n31306), .ZN(n30829) );
  NAND4_X1 U33313 ( .A1(n30653), .A2(n31294), .A3(n30834), .A4(n30829), .ZN(
        n24786) );
  XNOR2_X1 U33314 ( .A(n24790), .B(n25483), .ZN(n27264) );
  XNOR2_X1 U33315 ( .A(n24791), .B(n4529), .ZN(n26030) );
  XNOR2_X1 U33316 ( .A(n24792), .B(n26030), .ZN(n26439) );
  XNOR2_X1 U33317 ( .A(n27264), .B(n26439), .ZN(n24794) );
  XNOR2_X1 U33318 ( .A(n26175), .B(n24793), .ZN(n26599) );
  XNOR2_X1 U33319 ( .A(n24794), .B(n26599), .ZN(n24802) );
  XNOR2_X1 U33320 ( .A(n4754), .B(n4916), .ZN(n24796) );
  XNOR2_X1 U33321 ( .A(n24797), .B(n24796), .ZN(n24798) );
  XNOR2_X1 U33322 ( .A(n25168), .B(n24798), .ZN(n41960) );
  XNOR2_X1 U33323 ( .A(n43252), .B(n41960), .ZN(n24799) );
  XNOR2_X1 U33324 ( .A(n27477), .B(n24799), .ZN(n24800) );
  XNOR2_X1 U33325 ( .A(n25608), .B(n24800), .ZN(n24801) );
  XNOR2_X1 U33326 ( .A(n25508), .B(n44954), .ZN(n24804) );
  XNOR2_X1 U33327 ( .A(n27290), .B(n24804), .ZN(n24806) );
  XNOR2_X1 U33328 ( .A(n25268), .B(n25762), .ZN(n24805) );
  XNOR2_X1 U33329 ( .A(n24805), .B(n24806), .ZN(n25182) );
  XNOR2_X1 U33330 ( .A(n43316), .B(n42889), .ZN(n24807) );
  XNOR2_X1 U33331 ( .A(n27241), .B(n24807), .ZN(n24808) );
  XNOR2_X1 U33332 ( .A(n24808), .B(n28220), .ZN(n24809) );
  XNOR2_X1 U33333 ( .A(n24809), .B(n27439), .ZN(n24813) );
  INV_X1 U33334 ( .A(n26425), .ZN(n24811) );
  XNOR2_X1 U33335 ( .A(n24811), .B(n25351), .ZN(n24812) );
  XNOR2_X1 U33336 ( .A(n24814), .B(n25504), .ZN(n25001) );
  INV_X1 U33337 ( .A(n25001), .ZN(n24815) );
  XNOR2_X1 U33338 ( .A(n369), .B(n27447), .ZN(n24816) );
  XNOR2_X1 U33339 ( .A(n24816), .B(n27445), .ZN(n28113) );
  XNOR2_X1 U33340 ( .A(n25740), .B(n25429), .ZN(n24817) );
  XNOR2_X1 U33341 ( .A(n4589), .B(n49323), .ZN(n27387) );
  XNOR2_X1 U33342 ( .A(n24818), .B(n27387), .ZN(n42742) );
  XNOR2_X1 U33343 ( .A(n4295), .B(n3336), .ZN(n24819) );
  XNOR2_X1 U33344 ( .A(n24819), .B(n4723), .ZN(n24821) );
  XNOR2_X1 U33345 ( .A(n24821), .B(n24820), .ZN(n43674) );
  XNOR2_X1 U33346 ( .A(n43674), .B(n43691), .ZN(n24822) );
  XNOR2_X1 U33347 ( .A(n42742), .B(n24822), .ZN(n24823) );
  XNOR2_X1 U33348 ( .A(n27451), .B(n24823), .ZN(n24824) );
  XNOR2_X1 U33349 ( .A(n24825), .B(n24824), .ZN(n24826) );
  XNOR2_X1 U33350 ( .A(n749), .B(n26390), .ZN(n25218) );
  XNOR2_X1 U33351 ( .A(n26377), .B(n51415), .ZN(n24834) );
  INV_X1 U33352 ( .A(n24827), .ZN(n33807) );
  XNOR2_X1 U33353 ( .A(n33807), .B(n1336), .ZN(n43633) );
  XNOR2_X1 U33354 ( .A(n24828), .B(n4651), .ZN(n24829) );
  XNOR2_X1 U33355 ( .A(n24830), .B(n24829), .ZN(n42771) );
  XNOR2_X1 U33356 ( .A(n42771), .B(n42769), .ZN(n24831) );
  XNOR2_X1 U33357 ( .A(n43633), .B(n24831), .ZN(n24832) );
  XNOR2_X1 U33358 ( .A(n26378), .B(n24832), .ZN(n24833) );
  XNOR2_X1 U33359 ( .A(n24834), .B(n24833), .ZN(n24835) );
  XNOR2_X1 U33360 ( .A(n26547), .B(n26544), .ZN(n25569) );
  INV_X1 U33361 ( .A(n25569), .ZN(n25953) );
  XNOR2_X1 U33362 ( .A(n25953), .B(n24835), .ZN(n24836) );
  XNOR2_X1 U33363 ( .A(n26294), .B(n24836), .ZN(n24840) );
  XNOR2_X1 U33364 ( .A(n24904), .B(n24905), .ZN(n27222) );
  XNOR2_X1 U33365 ( .A(n27222), .B(n24837), .ZN(n24839) );
  XNOR2_X1 U33366 ( .A(n27226), .B(n488), .ZN(n24838) );
  XNOR2_X1 U33367 ( .A(n51441), .B(n27420), .ZN(n24841) );
  XNOR2_X1 U33368 ( .A(n24841), .B(n28371), .ZN(n28054) );
  XNOR2_X1 U33370 ( .A(n25934), .B(n28249), .ZN(n24853) );
  INV_X1 U33371 ( .A(n24843), .ZN(n24844) );
  XNOR2_X1 U33372 ( .A(n24844), .B(n33930), .ZN(n43866) );
  XNOR2_X1 U33373 ( .A(n42816), .B(n4883), .ZN(n43927) );
  XNOR2_X1 U33374 ( .A(n43863), .B(n43200), .ZN(n24845) );
  XNOR2_X1 U33375 ( .A(n43927), .B(n24845), .ZN(n24846) );
  XNOR2_X1 U33376 ( .A(n24846), .B(n42241), .ZN(n24847) );
  XNOR2_X1 U33377 ( .A(n43866), .B(n24847), .ZN(n24848) );
  XNOR2_X1 U33378 ( .A(n24849), .B(n24848), .ZN(n24851) );
  XNOR2_X1 U33379 ( .A(n24851), .B(n24850), .ZN(n24852) );
  XNOR2_X1 U33380 ( .A(n24853), .B(n24852), .ZN(n24854) );
  XNOR2_X1 U33381 ( .A(n28054), .B(n24854), .ZN(n24858) );
  XNOR2_X1 U33382 ( .A(n24855), .B(n25806), .ZN(n24857) );
  INV_X1 U33383 ( .A(n24856), .ZN(n26273) );
  INV_X1 U33385 ( .A(n30291), .ZN(n28144) );
  NOR2_X1 U33387 ( .A1(n27111), .A2(n30282), .ZN(n24859) );
  INV_X1 U33388 ( .A(n30279), .ZN(n28555) );
  XNOR2_X1 U33389 ( .A(n25385), .B(n27502), .ZN(n24860) );
  XNOR2_X1 U33390 ( .A(n24860), .B(n2125), .ZN(n24864) );
  XNOR2_X1 U33391 ( .A(n24861), .B(n4649), .ZN(n35067) );
  XNOR2_X1 U33392 ( .A(n35067), .B(n4636), .ZN(n24862) );
  XNOR2_X1 U33393 ( .A(n26530), .B(n24862), .ZN(n25155) );
  XNOR2_X1 U33394 ( .A(n26536), .B(n25155), .ZN(n24863) );
  XNOR2_X1 U33395 ( .A(n24864), .B(n24863), .ZN(n24871) );
  XNOR2_X1 U33396 ( .A(n24972), .B(n33374), .ZN(n43233) );
  XNOR2_X1 U33397 ( .A(n43233), .B(n42026), .ZN(n24865) );
  XNOR2_X1 U33398 ( .A(n28126), .B(n24865), .ZN(n24867) );
  XNOR2_X1 U33399 ( .A(n24866), .B(n24867), .ZN(n24870) );
  INV_X1 U33400 ( .A(n42721), .ZN(n41996) );
  XNOR2_X1 U33401 ( .A(n26402), .B(n41996), .ZN(n24868) );
  XNOR2_X1 U33402 ( .A(n24868), .B(n25825), .ZN(n25448) );
  INV_X1 U33403 ( .A(n25448), .ZN(n24869) );
  INV_X1 U33404 ( .A(n24872), .ZN(n24874) );
  INV_X1 U33405 ( .A(n24873), .ZN(n25231) );
  XNOR2_X1 U33406 ( .A(n25231), .B(n51121), .ZN(n25660) );
  XNOR2_X1 U33407 ( .A(n24874), .B(n25660), .ZN(n24875) );
  NAND3_X1 U33408 ( .A1(n30293), .A2(n30296), .A3(n30295), .ZN(n24876) );
  OAI21_X1 U33409 ( .B1(n30293), .B2(n30280), .A(n28560), .ZN(n24879) );
  NAND3_X1 U33410 ( .A1(n28557), .A2(n28559), .A3(n24879), .ZN(n24880) );
  INV_X1 U33412 ( .A(n30292), .ZN(n28146) );
  NAND2_X1 U33413 ( .A1(n27110), .A2(n30285), .ZN(n24883) );
  NAND2_X1 U33414 ( .A1(n28551), .A2(n30289), .ZN(n24886) );
  NAND2_X1 U33415 ( .A1(n28555), .A2(n51748), .ZN(n24885) );
  AOI21_X1 U33416 ( .B1(n24886), .B2(n24885), .A(n28560), .ZN(n24887) );
  NOR2_X1 U33417 ( .A1(n24888), .A2(n24887), .ZN(n24889) );
  XNOR2_X1 U33418 ( .A(n24891), .B(n28274), .ZN(n24899) );
  XNOR2_X1 U33419 ( .A(n24893), .B(n24892), .ZN(n43907) );
  XNOR2_X1 U33420 ( .A(n24894), .B(n4597), .ZN(n24895) );
  XNOR2_X1 U33421 ( .A(n24896), .B(n24895), .ZN(n45288) );
  XNOR2_X1 U33422 ( .A(n43907), .B(n45288), .ZN(n24897) );
  XNOR2_X1 U33423 ( .A(n27373), .B(n24897), .ZN(n24898) );
  XNOR2_X1 U33424 ( .A(n24899), .B(n24898), .ZN(n24901) );
  XNOR2_X1 U33425 ( .A(n24901), .B(n24900), .ZN(n24903) );
  XNOR2_X1 U33426 ( .A(n26556), .B(n27368), .ZN(n24902) );
  XNOR2_X1 U33427 ( .A(n24902), .B(n24903), .ZN(n24910) );
  XNOR2_X1 U33428 ( .A(n25249), .B(n24904), .ZN(n24907) );
  INV_X1 U33429 ( .A(n24905), .ZN(n24906) );
  XNOR2_X1 U33430 ( .A(n24907), .B(n24906), .ZN(n25119) );
  XNOR2_X1 U33431 ( .A(n26300), .B(n25724), .ZN(n24908) );
  XNOR2_X1 U33433 ( .A(n25119), .B(n28041), .ZN(n24909) );
  XNOR2_X1 U33434 ( .A(n24910), .B(n24909), .ZN(n24914) );
  XNOR2_X1 U33435 ( .A(n24912), .B(n24911), .ZN(n25717) );
  INV_X1 U33436 ( .A(n25717), .ZN(n24913) );
  XNOR2_X1 U33437 ( .A(n26362), .B(n51423), .ZN(n28248) );
  XNOR2_X1 U33438 ( .A(n37008), .B(n34414), .ZN(n25135) );
  XNOR2_X1 U33439 ( .A(n25683), .B(n4316), .ZN(n24917) );
  XNOR2_X1 U33440 ( .A(n25135), .B(n24917), .ZN(n24918) );
  XNOR2_X1 U33441 ( .A(n24918), .B(n39718), .ZN(n46048) );
  XNOR2_X1 U33442 ( .A(n4883), .B(n4312), .ZN(n43862) );
  XNOR2_X1 U33443 ( .A(n43862), .B(n45883), .ZN(n24920) );
  XNOR2_X1 U33444 ( .A(n24920), .B(n24919), .ZN(n44349) );
  XNOR2_X1 U33445 ( .A(n46048), .B(n44349), .ZN(n24921) );
  XNOR2_X1 U33446 ( .A(n28049), .B(n24921), .ZN(n24922) );
  XNOR2_X1 U33447 ( .A(n24924), .B(n27479), .ZN(n26254) );
  INV_X1 U33448 ( .A(n24925), .ZN(n42266) );
  INV_X1 U33449 ( .A(n28069), .ZN(n26265) );
  XNOR2_X1 U33450 ( .A(n25481), .B(n26265), .ZN(n24931) );
  XNOR2_X1 U33451 ( .A(n36941), .B(n4691), .ZN(n24927) );
  XNOR2_X1 U33452 ( .A(n25168), .B(n24927), .ZN(n41401) );
  XNOR2_X1 U33453 ( .A(n41401), .B(n24928), .ZN(n24929) );
  XNOR2_X1 U33454 ( .A(n25365), .B(n24929), .ZN(n24930) );
  XNOR2_X1 U33455 ( .A(n24931), .B(n24930), .ZN(n24935) );
  INV_X1 U33456 ( .A(n24932), .ZN(n24933) );
  XNOR2_X1 U33457 ( .A(n24933), .B(n47268), .ZN(n43728) );
  XNOR2_X1 U33458 ( .A(n27267), .B(n25604), .ZN(n24934) );
  XNOR2_X1 U33459 ( .A(n24935), .B(n24934), .ZN(n24939) );
  XNOR2_X1 U33460 ( .A(n24936), .B(n25483), .ZN(n26450) );
  XNOR2_X1 U33461 ( .A(n26600), .B(n25703), .ZN(n24937) );
  XNOR2_X1 U33462 ( .A(n26450), .B(n24937), .ZN(n24938) );
  XNOR2_X1 U33463 ( .A(n24939), .B(n24938), .ZN(n24940) );
  INV_X1 U33464 ( .A(n30248), .ZN(n29147) );
  XNOR2_X1 U33465 ( .A(n24941), .B(n4628), .ZN(n45072) );
  XNOR2_X1 U33466 ( .A(n45072), .B(n42322), .ZN(n24943) );
  XNOR2_X1 U33467 ( .A(n24942), .B(n44483), .ZN(n42314) );
  XNOR2_X1 U33468 ( .A(n24944), .B(n26581), .ZN(n24946) );
  XNOR2_X1 U33469 ( .A(n24945), .B(n24946), .ZN(n24947) );
  XNOR2_X1 U33470 ( .A(n28218), .B(n24947), .ZN(n24955) );
  XNOR2_X1 U33471 ( .A(n26160), .B(n49109), .ZN(n24948) );
  XNOR2_X1 U33472 ( .A(n27250), .B(Key[160]), .ZN(n24949) );
  XNOR2_X1 U33473 ( .A(n24950), .B(n28095), .ZN(n24953) );
  XNOR2_X1 U33474 ( .A(n25351), .B(n25762), .ZN(n24951) );
  XNOR2_X1 U33475 ( .A(n24951), .B(n26239), .ZN(n24952) );
  XNOR2_X1 U33476 ( .A(n24953), .B(n24952), .ZN(n24954) );
  XNOR2_X1 U33477 ( .A(n24956), .B(n4817), .ZN(n45256) );
  INV_X1 U33478 ( .A(n45253), .ZN(n24957) );
  XNOR2_X1 U33479 ( .A(n24957), .B(n43968), .ZN(n43835) );
  XNOR2_X1 U33480 ( .A(n4647), .B(n4641), .ZN(n24958) );
  XNOR2_X1 U33481 ( .A(n43835), .B(n24958), .ZN(n24959) );
  XNOR2_X1 U33482 ( .A(n45256), .B(n24959), .ZN(n24960) );
  XNOR2_X1 U33483 ( .A(n28427), .B(n24960), .ZN(n24961) );
  XNOR2_X1 U33484 ( .A(n24961), .B(n28104), .ZN(n24962) );
  XNOR2_X1 U33485 ( .A(n24962), .B(n25590), .ZN(n24964) );
  XNOR2_X1 U33486 ( .A(n25927), .B(n43293), .ZN(n25646) );
  XNOR2_X1 U33487 ( .A(n24964), .B(n24963), .ZN(n24967) );
  XNOR2_X1 U33488 ( .A(n24965), .B(n368), .ZN(n24966) );
  XNOR2_X1 U33489 ( .A(n26216), .B(n24967), .ZN(n24971) );
  INV_X1 U33490 ( .A(n27445), .ZN(n24968) );
  XNOR2_X1 U33491 ( .A(n27382), .B(n28106), .ZN(n24969) );
  XNOR2_X1 U33492 ( .A(n26090), .B(n24969), .ZN(n24970) );
  XNOR2_X1 U33493 ( .A(n24972), .B(n25380), .ZN(n42844) );
  XNOR2_X1 U33494 ( .A(n42844), .B(n48843), .ZN(n24973) );
  XNOR2_X1 U33495 ( .A(n41314), .B(n24973), .ZN(n24974) );
  XNOR2_X1 U33496 ( .A(n25540), .B(n24974), .ZN(n24975) );
  XNOR2_X1 U33497 ( .A(n25385), .B(n24975), .ZN(n24979) );
  XNOR2_X1 U33498 ( .A(n26530), .B(n28292), .ZN(n24977) );
  XNOR2_X1 U33499 ( .A(n25548), .B(n4653), .ZN(n26056) );
  XNOR2_X1 U33500 ( .A(n24977), .B(n26056), .ZN(n24978) );
  XNOR2_X1 U33501 ( .A(n24979), .B(n24978), .ZN(n24981) );
  XNOR2_X1 U33502 ( .A(n24981), .B(n24980), .ZN(n24983) );
  XNOR2_X1 U33503 ( .A(n26228), .B(n25444), .ZN(n26520) );
  XNOR2_X1 U33504 ( .A(n2125), .B(n25154), .ZN(n24982) );
  XNOR2_X1 U33505 ( .A(n28129), .B(n28121), .ZN(n26523) );
  NAND2_X1 U33506 ( .A1(n27957), .A2(n29159), .ZN(n29152) );
  OR2_X1 U33507 ( .A1(n29172), .A2(n29152), .ZN(n29170) );
  NAND2_X1 U33508 ( .A1(n27951), .A2(n51473), .ZN(n26488) );
  AND2_X1 U33509 ( .A1(n29170), .A2(n26488), .ZN(n24987) );
  INV_X1 U33510 ( .A(n24984), .ZN(n30249) );
  INV_X1 U33511 ( .A(n29148), .ZN(n26483) );
  NOR2_X1 U33512 ( .A1(n29174), .A2(n26483), .ZN(n24985) );
  OAI21_X1 U33513 ( .B1(n30240), .B2(n24985), .A(n29153), .ZN(n24986) );
  XNOR2_X1 U33515 ( .A(n24991), .B(n26234), .ZN(n24999) );
  INV_X1 U33516 ( .A(n28089), .ZN(n24993) );
  XNOR2_X1 U33517 ( .A(n24992), .B(n4864), .ZN(n43588) );
  XNOR2_X1 U33518 ( .A(n24993), .B(n43588), .ZN(n42551) );
  XNOR2_X1 U33519 ( .A(n33192), .B(n4486), .ZN(n44069) );
  XNOR2_X1 U33520 ( .A(n44069), .B(n31432), .ZN(n24994) );
  XNOR2_X1 U33521 ( .A(n42551), .B(n24994), .ZN(n24995) );
  XNOR2_X1 U33522 ( .A(n25501), .B(n24995), .ZN(n24996) );
  XNOR2_X1 U33523 ( .A(n25495), .B(n24996), .ZN(n24997) );
  XNOR2_X1 U33524 ( .A(n24997), .B(n23621), .ZN(n24998) );
  XNOR2_X1 U33525 ( .A(n24999), .B(n24998), .ZN(n25000) );
  XNOR2_X1 U33526 ( .A(n25001), .B(n25000), .ZN(n25007) );
  XNOR2_X1 U33527 ( .A(n26435), .B(n25003), .ZN(n25004) );
  XNOR2_X1 U33528 ( .A(n25005), .B(n25004), .ZN(n25677) );
  XNOR2_X1 U33529 ( .A(n25533), .B(n25677), .ZN(n25006) );
  XNOR2_X1 U33530 ( .A(n51648), .B(n26264), .ZN(n25008) );
  XNOR2_X1 U33531 ( .A(n25485), .B(n25008), .ZN(n25009) );
  XNOR2_X1 U33532 ( .A(n25010), .B(n25009), .ZN(n25011) );
  XNOR2_X1 U33533 ( .A(n25012), .B(n25011), .ZN(n25021) );
  XNOR2_X1 U33534 ( .A(n25883), .B(n27479), .ZN(n25712) );
  XNOR2_X1 U33535 ( .A(n33123), .B(n25013), .ZN(n44976) );
  XOR2_X1 U33536 ( .A(n4855), .B(n4836), .Z(n25014) );
  XNOR2_X1 U33537 ( .A(n44976), .B(n25014), .ZN(n25015) );
  XNOR2_X1 U33538 ( .A(n25284), .B(n33495), .ZN(n42688) );
  XNOR2_X1 U33539 ( .A(n25015), .B(n42688), .ZN(n25016) );
  XNOR2_X1 U33540 ( .A(n28352), .B(n25016), .ZN(n25017) );
  XNOR2_X1 U33541 ( .A(n25018), .B(n25610), .ZN(n25019) );
  XNOR2_X1 U33542 ( .A(n25712), .B(n25019), .ZN(n25020) );
  XNOR2_X1 U33543 ( .A(n25022), .B(n4579), .ZN(n25023) );
  XNOR2_X1 U33544 ( .A(n42083), .B(n25023), .ZN(n25024) );
  XNOR2_X1 U33545 ( .A(n43371), .B(n25024), .ZN(n25025) );
  XNOR2_X1 U33546 ( .A(n27424), .B(n25025), .ZN(n25026) );
  XNOR2_X1 U33547 ( .A(n25346), .B(n25026), .ZN(n25028) );
  XNOR2_X1 U33548 ( .A(n26565), .B(n25937), .ZN(n25027) );
  XNOR2_X1 U33549 ( .A(n25028), .B(n25027), .ZN(n25031) );
  XNOR2_X1 U33550 ( .A(n33297), .B(n45106), .ZN(n35741) );
  XNOR2_X1 U33551 ( .A(n25813), .B(n35741), .ZN(n25030) );
  XNOR2_X1 U33552 ( .A(n25030), .B(n2106), .ZN(n26277) );
  XNOR2_X1 U33553 ( .A(n25031), .B(n26277), .ZN(n25034) );
  XNOR2_X1 U33554 ( .A(n26285), .B(n25947), .ZN(n25032) );
  XNOR2_X1 U33555 ( .A(n27419), .B(n25032), .ZN(n25033) );
  XNOR2_X1 U33556 ( .A(n25033), .B(n28249), .ZN(n25695) );
  XNOR2_X1 U33557 ( .A(n25034), .B(n25695), .ZN(n25038) );
  XNOR2_X1 U33558 ( .A(n28371), .B(n25466), .ZN(n25036) );
  XNOR2_X1 U33559 ( .A(n25035), .B(n25036), .ZN(n25037) );
  XNOR2_X1 U33560 ( .A(n25038), .B(n25037), .ZN(n25421) );
  XNOR2_X1 U33561 ( .A(n25039), .B(n26544), .ZN(n26141) );
  XNOR2_X1 U33562 ( .A(n26547), .B(n26141), .ZN(n25125) );
  XNOR2_X1 U33563 ( .A(n25041), .B(n25040), .ZN(n43530) );
  XOR2_X1 U33564 ( .A(n4454), .B(n4578), .Z(n25043) );
  XNOR2_X1 U33565 ( .A(n25043), .B(n25042), .ZN(n44191) );
  XNOR2_X1 U33566 ( .A(n43530), .B(n44191), .ZN(n25044) );
  XNOR2_X1 U33567 ( .A(n25124), .B(n25044), .ZN(n25045) );
  XNOR2_X1 U33568 ( .A(n25726), .B(n25045), .ZN(n25046) );
  XNOR2_X1 U33569 ( .A(n25125), .B(n25046), .ZN(n25049) );
  XNOR2_X1 U33570 ( .A(n25798), .B(n25571), .ZN(n25048) );
  XNOR2_X1 U33571 ( .A(n25048), .B(n52163), .ZN(n25463) );
  XNOR2_X1 U33572 ( .A(n28274), .B(n4415), .ZN(n25051) );
  XNOR2_X1 U33573 ( .A(n25050), .B(n25051), .ZN(n25313) );
  NAND2_X1 U33574 ( .A1(n25053), .A2(n25052), .ZN(n25069) );
  OAI211_X1 U33575 ( .C1(n25054), .C2(n25064), .A(n25062), .B(n25061), .ZN(
        n25068) );
  NAND4_X1 U33576 ( .A1(n25058), .A2(n25057), .A3(n38626), .A4(n25056), .ZN(
        n25059) );
  OAI211_X1 U33577 ( .C1(n25062), .C2(n25061), .A(n25060), .B(n25059), .ZN(
        n25063) );
  INV_X1 U33578 ( .A(n25063), .ZN(n25067) );
  NAND3_X1 U33579 ( .A1(n25065), .A2(n38626), .A3(n25064), .ZN(n25066) );
  OAI211_X1 U33580 ( .C1(n25069), .C2(n25068), .A(n25067), .B(n25066), .ZN(
        n26302) );
  XNOR2_X1 U33581 ( .A(n26302), .B(n26377), .ZN(n25070) );
  XNOR2_X1 U33582 ( .A(n25313), .B(n25070), .ZN(n25073) );
  XNOR2_X1 U33583 ( .A(n488), .B(n25071), .ZN(n25072) );
  XNOR2_X1 U33584 ( .A(n25073), .B(n25072), .ZN(n25074) );
  NOR2_X1 U33585 ( .A1(n30263), .A2(n1708), .ZN(n29222) );
  XNOR2_X1 U33586 ( .A(n26395), .B(n28423), .ZN(n25077) );
  XNOR2_X1 U33587 ( .A(n26044), .B(n26508), .ZN(n25076) );
  XNOR2_X1 U33588 ( .A(n25077), .B(n25076), .ZN(n25083) );
  XNOR2_X1 U33589 ( .A(n25927), .B(n26210), .ZN(n25321) );
  XNOR2_X1 U33590 ( .A(n25924), .B(n4650), .ZN(n25079) );
  XNOR2_X1 U33591 ( .A(n25079), .B(n25078), .ZN(n43553) );
  XNOR2_X1 U33592 ( .A(n44220), .B(n43553), .ZN(n25080) );
  XNOR2_X1 U33593 ( .A(n25747), .B(n25080), .ZN(n25081) );
  XNOR2_X1 U33594 ( .A(n25321), .B(n25081), .ZN(n25082) );
  XNOR2_X1 U33595 ( .A(n25086), .B(n25639), .ZN(n25089) );
  XNOR2_X1 U33596 ( .A(n25088), .B(n25087), .ZN(n25600) );
  XNOR2_X1 U33598 ( .A(n25825), .B(n25161), .ZN(n25090) );
  XNOR2_X1 U33599 ( .A(n25090), .B(n25829), .ZN(n25092) );
  XNOR2_X1 U33600 ( .A(n471), .B(n25091), .ZN(n25390) );
  XNOR2_X1 U33601 ( .A(n25229), .B(n26531), .ZN(n25093) );
  XNOR2_X1 U33602 ( .A(n25093), .B(n26119), .ZN(n25544) );
  XNOR2_X1 U33603 ( .A(n25095), .B(n25094), .ZN(n44889) );
  XNOR2_X1 U33604 ( .A(n4668), .B(n4487), .ZN(n25096) );
  XNOR2_X1 U33605 ( .A(n25097), .B(n25096), .ZN(n42646) );
  XNOR2_X1 U33606 ( .A(n42646), .B(n4874), .ZN(n25098) );
  XNOR2_X1 U33607 ( .A(n44889), .B(n25098), .ZN(n25099) );
  XNOR2_X1 U33608 ( .A(n25909), .B(n25099), .ZN(n25100) );
  XNOR2_X1 U33609 ( .A(n25831), .B(n25100), .ZN(n25101) );
  XNOR2_X1 U33610 ( .A(n25101), .B(n25544), .ZN(n25102) );
  OAI22_X1 U33611 ( .A1(n29222), .A2(n8720), .B1(n29242), .B2(n30269), .ZN(
        n25105) );
  NOR2_X1 U33612 ( .A1(n30272), .A2(n1708), .ZN(n29232) );
  NAND2_X1 U33613 ( .A1(n29232), .A2(n29241), .ZN(n25417) );
  NAND2_X1 U33614 ( .A1(n27913), .A2(n25415), .ZN(n25104) );
  NAND3_X1 U33615 ( .A1(n25105), .A2(n25417), .A3(n25104), .ZN(n25113) );
  NAND2_X1 U33617 ( .A1(n25108), .A2(n25107), .ZN(n25110) );
  OR2_X1 U33618 ( .A1(n29226), .A2(n25075), .ZN(n25109) );
  XNOR2_X1 U33620 ( .A(n25115), .B(n25114), .ZN(n43784) );
  XNOR2_X1 U33621 ( .A(n43784), .B(n26541), .ZN(n25116) );
  XNOR2_X1 U33622 ( .A(n35673), .B(n25116), .ZN(n25117) );
  XNOR2_X1 U33623 ( .A(n26540), .B(n25117), .ZN(n25118) );
  XNOR2_X1 U33624 ( .A(n25118), .B(n26304), .ZN(n25120) );
  XNOR2_X1 U33625 ( .A(n25120), .B(n25119), .ZN(n25121) );
  XNOR2_X1 U33626 ( .A(n27491), .B(n25121), .ZN(n25123) );
  XNOR2_X1 U33627 ( .A(n26292), .B(n25122), .ZN(n28408) );
  XNOR2_X1 U33628 ( .A(n25123), .B(n28408), .ZN(n25126) );
  XNOR2_X1 U33629 ( .A(n28247), .B(n25127), .ZN(n25129) );
  XNOR2_X1 U33630 ( .A(n26573), .B(n25554), .ZN(n25128) );
  XNOR2_X1 U33631 ( .A(n27211), .B(n25128), .ZN(n26364) );
  XNOR2_X1 U33632 ( .A(n51119), .B(n25130), .ZN(n25139) );
  INV_X1 U33633 ( .A(n25132), .ZN(n25133) );
  XNOR2_X1 U33634 ( .A(n25133), .B(n2608), .ZN(n44135) );
  XNOR2_X1 U33635 ( .A(n25135), .B(n25134), .ZN(n43538) );
  XNOR2_X1 U33636 ( .A(n44135), .B(n43538), .ZN(n25136) );
  XNOR2_X1 U33637 ( .A(n26565), .B(n25136), .ZN(n25137) );
  XNOR2_X1 U33638 ( .A(n25141), .B(n2107), .ZN(n25566) );
  INV_X1 U33639 ( .A(n369), .ZN(n25142) );
  INV_X1 U33640 ( .A(n25145), .ZN(n25146) );
  XNOR2_X1 U33641 ( .A(n25146), .B(n42668), .ZN(n43694) );
  XNOR2_X1 U33642 ( .A(n25148), .B(n25147), .ZN(n42434) );
  XNOR2_X1 U33643 ( .A(n42434), .B(n4647), .ZN(n25149) );
  XNOR2_X1 U33644 ( .A(n43694), .B(n25149), .ZN(n25150) );
  XNOR2_X1 U33645 ( .A(n26210), .B(n25150), .ZN(n25151) );
  XNOR2_X1 U33646 ( .A(n25929), .B(n25151), .ZN(n25152) );
  XNOR2_X1 U33647 ( .A(n28129), .B(n25154), .ZN(n25157) );
  XNOR2_X1 U33648 ( .A(n471), .B(n25155), .ZN(n25156) );
  XNOR2_X1 U33649 ( .A(n25157), .B(n25156), .ZN(n25158) );
  XNOR2_X1 U33650 ( .A(n25158), .B(n25833), .ZN(n25167) );
  INV_X1 U33651 ( .A(n46126), .ZN(n35554) );
  XNOR2_X1 U33652 ( .A(n40847), .B(n48843), .ZN(n25159) );
  XNOR2_X1 U33653 ( .A(n35554), .B(n25159), .ZN(n25160) );
  XNOR2_X1 U33654 ( .A(n26529), .B(n25160), .ZN(n25162) );
  XNOR2_X1 U33655 ( .A(n25162), .B(n25161), .ZN(n25163) );
  XNOR2_X1 U33656 ( .A(n25163), .B(n25231), .ZN(n25165) );
  XNOR2_X1 U33657 ( .A(n25165), .B(n25164), .ZN(n25166) );
  XNOR2_X1 U33658 ( .A(n25169), .B(n25168), .ZN(n40305) );
  XNOR2_X1 U33659 ( .A(n25170), .B(n4855), .ZN(n25171) );
  XNOR2_X1 U33660 ( .A(n25172), .B(n25171), .ZN(n42958) );
  XNOR2_X1 U33661 ( .A(n40305), .B(n42958), .ZN(n25173) );
  XNOR2_X1 U33662 ( .A(n25174), .B(n25481), .ZN(n25175) );
  XNOR2_X1 U33663 ( .A(n26599), .B(n25175), .ZN(n25178) );
  XNOR2_X1 U33664 ( .A(n25176), .B(n27467), .ZN(n25177) );
  XNOR2_X1 U33665 ( .A(n25177), .B(n25608), .ZN(n26442) );
  XNOR2_X1 U33666 ( .A(n26442), .B(n25178), .ZN(n25180) );
  XNOR2_X1 U33667 ( .A(n25708), .B(n28352), .ZN(n25772) );
  XNOR2_X1 U33668 ( .A(n750), .B(n25772), .ZN(n26034) );
  XNOR2_X1 U33669 ( .A(n25712), .B(n26034), .ZN(n25179) );
  INV_X1 U33671 ( .A(n41924), .ZN(n33407) );
  XNOR2_X1 U33672 ( .A(n25181), .B(n25664), .ZN(n26429) );
  XNOR2_X1 U33673 ( .A(n25182), .B(n26429), .ZN(n25194) );
  XNOR2_X1 U33674 ( .A(n4676), .B(n4827), .ZN(n37239) );
  XNOR2_X1 U33675 ( .A(n37239), .B(n25183), .ZN(n42674) );
  XNOR2_X1 U33676 ( .A(n44952), .B(n42322), .ZN(n25184) );
  XNOR2_X1 U33677 ( .A(n42674), .B(n25184), .ZN(n25185) );
  XNOR2_X1 U33678 ( .A(n25493), .B(n25185), .ZN(n25186) );
  XNOR2_X1 U33679 ( .A(n28221), .B(n25186), .ZN(n25187) );
  XNOR2_X1 U33680 ( .A(n25188), .B(n25187), .ZN(n25192) );
  XNOR2_X1 U33681 ( .A(n27250), .B(n26160), .ZN(n25190) );
  INV_X1 U33682 ( .A(n26234), .ZN(n25189) );
  XNOR2_X1 U33683 ( .A(n25190), .B(n25189), .ZN(n25191) );
  XNOR2_X1 U33684 ( .A(n25192), .B(n25191), .ZN(n25193) );
  OAI21_X1 U33685 ( .B1(n28022), .B2(n30181), .A(n30312), .ZN(n25197) );
  INV_X1 U33686 ( .A(n30178), .ZN(n30183) );
  INV_X1 U33687 ( .A(n26468), .ZN(n25196) );
  NOR2_X1 U33689 ( .A1(n25199), .A2(n30306), .ZN(n25195) );
  AOI21_X1 U33690 ( .B1(n25197), .B2(n25196), .A(n25195), .ZN(n25204) );
  NAND2_X1 U33691 ( .A1(n30179), .A2(n30180), .ZN(n28032) );
  INV_X1 U33692 ( .A(n28032), .ZN(n30177) );
  NAND3_X1 U33693 ( .A1(n30177), .A2(n30306), .A3(n547), .ZN(n25202) );
  NAND3_X1 U33694 ( .A1(n29140), .A2(n28025), .A3(n1771), .ZN(n25201) );
  XNOR2_X1 U33696 ( .A(n25208), .B(n25207), .ZN(n44012) );
  XNOR2_X1 U33697 ( .A(n25210), .B(n25209), .ZN(n42562) );
  XNOR2_X1 U33698 ( .A(n42562), .B(n42995), .ZN(n25211) );
  XNOR2_X1 U33699 ( .A(n44012), .B(n25211), .ZN(n25212) );
  XNOR2_X1 U33700 ( .A(n25213), .B(n25212), .ZN(n25214) );
  XNOR2_X1 U33701 ( .A(n28103), .B(n25214), .ZN(n25216) );
  XNOR2_X1 U33702 ( .A(n25216), .B(n51502), .ZN(n25217) );
  XNOR2_X1 U33703 ( .A(n25218), .B(n25217), .ZN(n25219) );
  XNOR2_X1 U33704 ( .A(n28437), .B(n25219), .ZN(n25221) );
  XNOR2_X1 U33705 ( .A(n28391), .B(n33374), .ZN(n27348) );
  XNOR2_X1 U33706 ( .A(n25897), .B(n33845), .ZN(n25222) );
  XNOR2_X1 U33707 ( .A(n27348), .B(n25222), .ZN(n43137) );
  XNOR2_X1 U33708 ( .A(n28390), .B(n48843), .ZN(n41864) );
  XNOR2_X1 U33709 ( .A(n43137), .B(n41864), .ZN(n25223) );
  XNOR2_X1 U33710 ( .A(n28292), .B(n25223), .ZN(n25224) );
  XNOR2_X1 U33711 ( .A(n25226), .B(n25225), .ZN(n25227) );
  XNOR2_X1 U33712 ( .A(n25228), .B(n25227), .ZN(n25234) );
  XNOR2_X1 U33713 ( .A(n4177), .B(n4286), .ZN(n43130) );
  XNOR2_X1 U33714 ( .A(n25229), .B(n43130), .ZN(n25230) );
  XNOR2_X1 U33715 ( .A(n25231), .B(n25230), .ZN(n28123) );
  XNOR2_X1 U33716 ( .A(n2212), .B(n51121), .ZN(n25232) );
  XNOR2_X1 U33717 ( .A(n28123), .B(n25232), .ZN(n25233) );
  XNOR2_X1 U33718 ( .A(n25234), .B(n25233), .ZN(n28587) );
  INV_X1 U33719 ( .A(n28587), .ZN(n27121) );
  XNOR2_X1 U33720 ( .A(n4045), .B(n4637), .ZN(n25235) );
  XNOR2_X1 U33721 ( .A(n25236), .B(n25235), .ZN(n25237) );
  XNOR2_X1 U33722 ( .A(n37140), .B(n25237), .ZN(n25238) );
  XNOR2_X1 U33723 ( .A(n45310), .B(n25238), .ZN(n25239) );
  XNOR2_X1 U33724 ( .A(n25554), .B(n25239), .ZN(n25241) );
  XNOR2_X1 U33725 ( .A(n25241), .B(n25240), .ZN(n25242) );
  XNOR2_X1 U33726 ( .A(n25242), .B(n26571), .ZN(n25245) );
  XNOR2_X1 U33727 ( .A(n51441), .B(n28056), .ZN(n25244) );
  XNOR2_X1 U33728 ( .A(n25245), .B(n25244), .ZN(n25247) );
  XNOR2_X1 U33729 ( .A(n25680), .B(n28049), .ZN(n25246) );
  XNOR2_X1 U33730 ( .A(n25681), .B(n25246), .ZN(n25936) );
  XNOR2_X1 U33731 ( .A(n25247), .B(n25936), .ZN(n25248) );
  XNOR2_X1 U33732 ( .A(n27218), .B(n25806), .ZN(n28388) );
  NOR2_X1 U33733 ( .A1(n28579), .A2(n28897), .ZN(n26475) );
  INV_X1 U33734 ( .A(n25249), .ZN(n25250) );
  XNOR2_X1 U33735 ( .A(n25250), .B(n26377), .ZN(n25251) );
  XNOR2_X1 U33736 ( .A(n25251), .B(n28035), .ZN(n25253) );
  XNOR2_X1 U33737 ( .A(n25253), .B(n25252), .ZN(n25262) );
  INV_X1 U33738 ( .A(n25575), .ZN(n25254) );
  XNOR2_X1 U33739 ( .A(n25255), .B(n25254), .ZN(n36996) );
  XNOR2_X1 U33740 ( .A(n36996), .B(n49414), .ZN(n42522) );
  XNOR2_X1 U33741 ( .A(n1336), .B(n4705), .ZN(n25256) );
  XNOR2_X1 U33742 ( .A(n25718), .B(n25256), .ZN(n44057) );
  XNOR2_X1 U33743 ( .A(n42522), .B(n44057), .ZN(n25257) );
  XNOR2_X1 U33744 ( .A(n27373), .B(n25257), .ZN(n25258) );
  XNOR2_X1 U33745 ( .A(n28410), .B(n25258), .ZN(n25260) );
  XNOR2_X1 U33746 ( .A(n25260), .B(n25259), .ZN(n25261) );
  XNOR2_X1 U33747 ( .A(n25262), .B(n25261), .ZN(n25263) );
  XNOR2_X1 U33748 ( .A(n27235), .B(n25569), .ZN(n27377) );
  INV_X1 U33749 ( .A(n28907), .ZN(n26476) );
  XNOR2_X1 U33750 ( .A(n28220), .B(n25493), .ZN(n25264) );
  XNOR2_X1 U33751 ( .A(n28221), .B(n25264), .ZN(n25265) );
  XNOR2_X1 U33752 ( .A(n51484), .B(n25265), .ZN(n25266) );
  XNOR2_X1 U33753 ( .A(n25267), .B(n25266), .ZN(n25363) );
  XNOR2_X1 U33754 ( .A(n25268), .B(n26425), .ZN(n25269) );
  XNOR2_X1 U33755 ( .A(n25269), .B(n25270), .ZN(n25279) );
  XNOR2_X1 U33756 ( .A(n25501), .B(n4733), .ZN(n28093) );
  XNOR2_X1 U33757 ( .A(n26591), .B(n28093), .ZN(n25277) );
  INV_X1 U33758 ( .A(n25271), .ZN(n25272) );
  XNOR2_X1 U33759 ( .A(n25272), .B(n2601), .ZN(n41462) );
  XNOR2_X1 U33760 ( .A(n25273), .B(n4827), .ZN(n42891) );
  XNOR2_X1 U33761 ( .A(n42891), .B(n41426), .ZN(n25274) );
  XNOR2_X1 U33762 ( .A(n41462), .B(n25274), .ZN(n25275) );
  XNOR2_X1 U33763 ( .A(n26581), .B(n25275), .ZN(n25276) );
  XNOR2_X1 U33764 ( .A(n25277), .B(n25276), .ZN(n25278) );
  XNOR2_X1 U33765 ( .A(n25279), .B(n25278), .ZN(n25280) );
  XNOR2_X1 U33766 ( .A(n25280), .B(n25363), .ZN(n25297) );
  XNOR2_X1 U33767 ( .A(n25481), .B(n26600), .ZN(n25287) );
  XNOR2_X1 U33768 ( .A(n25281), .B(n26604), .ZN(n33330) );
  XNOR2_X1 U33769 ( .A(n26178), .B(n45736), .ZN(n25282) );
  XNOR2_X1 U33770 ( .A(n33330), .B(n25282), .ZN(n41873) );
  XNOR2_X1 U33771 ( .A(n4655), .B(n4818), .ZN(n25283) );
  XNOR2_X1 U33772 ( .A(n25284), .B(n25283), .ZN(n43108) );
  XNOR2_X1 U33773 ( .A(n41873), .B(n43108), .ZN(n25285) );
  XNOR2_X1 U33774 ( .A(n51749), .B(n25285), .ZN(n25286) );
  XNOR2_X1 U33775 ( .A(n25287), .B(n25286), .ZN(n25288) );
  XNOR2_X1 U33776 ( .A(n25288), .B(n26439), .ZN(n25290) );
  XNOR2_X1 U33777 ( .A(n25290), .B(n25289), .ZN(n25294) );
  XNOR2_X1 U33778 ( .A(n27479), .B(n25291), .ZN(n25292) );
  XNOR2_X1 U33779 ( .A(n25609), .B(n25610), .ZN(n27328) );
  XNOR2_X1 U33780 ( .A(n25292), .B(n27328), .ZN(n25293) );
  INV_X1 U33781 ( .A(n51118), .ZN(n27131) );
  AND2_X1 U33782 ( .A1(n28588), .A2(n27131), .ZN(n27999) );
  OAI21_X1 U33783 ( .B1(n26475), .B2(n26476), .A(n27999), .ZN(n25304) );
  NOR2_X1 U33784 ( .A1(n28579), .A2(n27119), .ZN(n25296) );
  INV_X1 U33785 ( .A(n27126), .ZN(n25295) );
  OAI21_X1 U33786 ( .B1(n25296), .B2(n25295), .A(n27128), .ZN(n25303) );
  INV_X1 U33787 ( .A(n25298), .ZN(n25301) );
  INV_X1 U33788 ( .A(n25297), .ZN(n28578) );
  NAND2_X1 U33789 ( .A1(n27132), .A2(n28578), .ZN(n27133) );
  AND2_X1 U33790 ( .A1(n27133), .A2(n27121), .ZN(n28590) );
  NAND2_X1 U33791 ( .A1(n27993), .A2(n51118), .ZN(n27123) );
  INV_X1 U33792 ( .A(n27987), .ZN(n28000) );
  AOI21_X1 U33793 ( .B1(n25298), .B2(n28578), .A(n28000), .ZN(n25299) );
  OAI211_X1 U33794 ( .C1(n27986), .C2(n25301), .A(n25300), .B(n25299), .ZN(
        n25302) );
  INV_X1 U33795 ( .A(n28579), .ZN(n27130) );
  INV_X1 U33797 ( .A(n27991), .ZN(n27129) );
  XNOR2_X1 U33798 ( .A(n26152), .B(n51416), .ZN(n25305) );
  XNOR2_X1 U33799 ( .A(n25306), .B(n25305), .ZN(n25307) );
  XNOR2_X1 U33800 ( .A(n25999), .B(n25307), .ZN(n25315) );
  XNOR2_X1 U33801 ( .A(n25308), .B(n27374), .ZN(n26148) );
  XNOR2_X1 U33802 ( .A(n25309), .B(n28266), .ZN(n45424) );
  XNOR2_X1 U33803 ( .A(n25578), .B(n2605), .ZN(n43803) );
  XNOR2_X1 U33804 ( .A(n45424), .B(n43803), .ZN(n25310) );
  XNOR2_X1 U33805 ( .A(n25724), .B(n25310), .ZN(n25311) );
  XNOR2_X1 U33806 ( .A(n26148), .B(n25311), .ZN(n25312) );
  XNOR2_X1 U33807 ( .A(n25313), .B(n25312), .ZN(n25314) );
  XNOR2_X1 U33808 ( .A(n25315), .B(n25314), .ZN(n25318) );
  XNOR2_X1 U33809 ( .A(n25319), .B(n751), .ZN(n25324) );
  XNOR2_X1 U33810 ( .A(n26044), .B(n25320), .ZN(n25742) );
  INV_X1 U33811 ( .A(n25321), .ZN(n25322) );
  XNOR2_X1 U33812 ( .A(n25742), .B(n25322), .ZN(n25323) );
  XNOR2_X1 U33813 ( .A(n34744), .B(n4723), .ZN(n43836) );
  XNOR2_X1 U33814 ( .A(n25325), .B(n4746), .ZN(n45379) );
  XNOR2_X1 U33815 ( .A(n43968), .B(n47737), .ZN(n25326) );
  XNOR2_X1 U33816 ( .A(n45379), .B(n25326), .ZN(n25327) );
  XNOR2_X1 U33817 ( .A(n43836), .B(n25327), .ZN(n25328) );
  XNOR2_X1 U33818 ( .A(n25740), .B(n25328), .ZN(n25329) );
  XNOR2_X1 U33819 ( .A(n25329), .B(n26395), .ZN(n25330) );
  XNOR2_X1 U33820 ( .A(n26393), .B(n25330), .ZN(n25331) );
  XNOR2_X1 U33821 ( .A(n27447), .B(n749), .ZN(n25332) );
  XNOR2_X1 U33822 ( .A(n25333), .B(n25332), .ZN(n25334) );
  AND2_X1 U33823 ( .A1(n29346), .A2(n30191), .ZN(n29337) );
  XNOR2_X1 U33824 ( .A(n26285), .B(n51424), .ZN(n25336) );
  XNOR2_X1 U33825 ( .A(n25336), .B(n26571), .ZN(n25337) );
  XNOR2_X1 U33826 ( .A(n25337), .B(n51380), .ZN(n26129) );
  XNOR2_X1 U33827 ( .A(n26129), .B(n25338), .ZN(n25350) );
  INV_X1 U33828 ( .A(n25937), .ZN(n25339) );
  XNOR2_X1 U33829 ( .A(n33635), .B(Key[189]), .ZN(n25340) );
  XNOR2_X1 U33830 ( .A(n25341), .B(n25340), .ZN(n25342) );
  XNOR2_X1 U33831 ( .A(n25343), .B(n25342), .ZN(n25344) );
  XNOR2_X1 U33832 ( .A(n25813), .B(n25344), .ZN(n25345) );
  XNOR2_X1 U33833 ( .A(n25346), .B(n25345), .ZN(n25347) );
  XNOR2_X1 U33834 ( .A(n28047), .B(n25347), .ZN(n25348) );
  XNOR2_X1 U33835 ( .A(n25348), .B(n27217), .ZN(n25349) );
  XNOR2_X1 U33836 ( .A(n25504), .B(n25351), .ZN(n25356) );
  XNOR2_X1 U33837 ( .A(n26159), .B(n25353), .ZN(n25510) );
  XNOR2_X1 U33838 ( .A(n25506), .B(n23621), .ZN(n25354) );
  XNOR2_X1 U33840 ( .A(n33914), .B(n4628), .ZN(n44485) );
  XNOR2_X1 U33841 ( .A(n31432), .B(n4823), .ZN(n25357) );
  XNOR2_X1 U33842 ( .A(n44485), .B(n25357), .ZN(n25358) );
  XNOR2_X1 U33843 ( .A(n25755), .B(n25358), .ZN(n25359) );
  XNOR2_X1 U33844 ( .A(n25359), .B(n25508), .ZN(n25361) );
  XNOR2_X1 U33845 ( .A(n25361), .B(n25360), .ZN(n25362) );
  XNOR2_X1 U33846 ( .A(n25363), .B(n25364), .ZN(n29343) );
  INV_X1 U33847 ( .A(n34709), .ZN(n43353) );
  XNOR2_X1 U33848 ( .A(n25775), .B(n43353), .ZN(n26177) );
  INV_X1 U33849 ( .A(n26177), .ZN(n25367) );
  XNOR2_X1 U33850 ( .A(n25367), .B(n25366), .ZN(n25368) );
  XNOR2_X1 U33851 ( .A(n25368), .B(n26450), .ZN(n25370) );
  XNOR2_X1 U33852 ( .A(n25883), .B(n25608), .ZN(n25369) );
  XNOR2_X1 U33853 ( .A(n25708), .B(n49790), .ZN(n27475) );
  INV_X1 U33854 ( .A(n25371), .ZN(n25373) );
  XNOR2_X1 U33855 ( .A(n25373), .B(n25372), .ZN(n25375) );
  XNOR2_X1 U33856 ( .A(n25375), .B(n25374), .ZN(n41742) );
  XNOR2_X1 U33857 ( .A(n25778), .B(n41742), .ZN(n25376) );
  XNOR2_X1 U33858 ( .A(n25376), .B(n26610), .ZN(n25377) );
  XNOR2_X1 U33859 ( .A(n27475), .B(n25377), .ZN(n25378) );
  XNOR2_X1 U33860 ( .A(n27467), .B(n25610), .ZN(n25893) );
  XNOR2_X1 U33861 ( .A(n25378), .B(n25893), .ZN(n25379) );
  NAND3_X1 U33863 ( .A1(n29337), .A2(n30200), .A3(n27886), .ZN(n30216) );
  INV_X1 U33864 ( .A(n30209), .ZN(n29345) );
  NAND2_X1 U33865 ( .A1(n29346), .A2(n30200), .ZN(n29344) );
  INV_X1 U33866 ( .A(n29343), .ZN(n27882) );
  NAND2_X1 U33867 ( .A1(n27882), .A2(n30191), .ZN(n29199) );
  OAI211_X1 U33868 ( .C1(n30202), .C2(n29345), .A(n29344), .B(n29199), .ZN(
        n25395) );
  XNOR2_X1 U33869 ( .A(n25380), .B(n4879), .ZN(n25381) );
  XNOR2_X1 U33870 ( .A(n25382), .B(n25381), .ZN(n43305) );
  XNOR2_X1 U33871 ( .A(n40847), .B(n4874), .ZN(n41661) );
  XNOR2_X1 U33872 ( .A(n41661), .B(n49937), .ZN(n25383) );
  XNOR2_X1 U33873 ( .A(n43305), .B(n25383), .ZN(n25384) );
  XNOR2_X1 U33874 ( .A(n25385), .B(n25384), .ZN(n25386) );
  XNOR2_X1 U33875 ( .A(n25386), .B(n51121), .ZN(n25388) );
  XNOR2_X1 U33876 ( .A(n25388), .B(n25387), .ZN(n25392) );
  XNOR2_X1 U33877 ( .A(n25445), .B(n2604), .ZN(n25389) );
  XNOR2_X1 U33878 ( .A(n2125), .B(n25389), .ZN(n25550) );
  XNOR2_X1 U33879 ( .A(n25550), .B(n25390), .ZN(n25391) );
  NAND2_X1 U33880 ( .A1(n25394), .A2(n51109), .ZN(n25402) );
  NAND2_X1 U33881 ( .A1(n25395), .A2(n29203), .ZN(n25398) );
  NAND2_X1 U33882 ( .A1(n733), .A2(n967), .ZN(n30194) );
  OAI21_X1 U33883 ( .B1(n30200), .B2(n30209), .A(n733), .ZN(n25396) );
  AOI22_X1 U33884 ( .A1(n30194), .A2(n27886), .B1(n25396), .B2(n29343), .ZN(
        n25397) );
  NAND2_X1 U33885 ( .A1(n25398), .A2(n25397), .ZN(n25401) );
  NAND2_X1 U33886 ( .A1(n27881), .A2(n733), .ZN(n25400) );
  NOR2_X1 U33887 ( .A1(n29200), .A2(n30202), .ZN(n29202) );
  NAND2_X1 U33888 ( .A1(n29202), .A2(n967), .ZN(n25399) );
  NOR2_X1 U33889 ( .A1(n32207), .A2(n32209), .ZN(n25403) );
  AOI22_X1 U33890 ( .A1(n31214), .A2(n25403), .B1(n31221), .B2(n716), .ZN(
        n25408) );
  OAI211_X1 U33892 ( .C1(n32214), .C2(n32212), .A(n5109), .B(n50981), .ZN(
        n25405) );
  NAND2_X1 U33893 ( .A1(n32209), .A2(n32212), .ZN(n31767) );
  XNOR2_X1 U33894 ( .A(n32194), .B(n32210), .ZN(n25404) );
  NAND4_X1 U33895 ( .A1(n30893), .A2(n25405), .A3(n31767), .A4(n25404), .ZN(
        n25406) );
  XNOR2_X1 U33897 ( .A(n34240), .B(n35835), .ZN(n32340) );
  OAI21_X1 U33898 ( .B1(n25415), .B2(n25411), .A(n29242), .ZN(n25414) );
  OAI21_X1 U33899 ( .B1(n30272), .B2(n25107), .A(n2158), .ZN(n25412) );
  NAND2_X1 U33900 ( .A1(n25412), .A2(n25420), .ZN(n25413) );
  AND3_X1 U33901 ( .A1(n29233), .A2(n25414), .A3(n25413), .ZN(n25852) );
  OAI21_X1 U33902 ( .B1(n1708), .B2(n30269), .A(n25415), .ZN(n25416) );
  AND2_X1 U33903 ( .A1(n25416), .A2(n25417), .ZN(n25851) );
  OAI21_X1 U33904 ( .B1(n25418), .B2(n1693), .A(n29110), .ZN(n25419) );
  OAI21_X1 U33905 ( .B1(n25420), .B2(n25419), .A(n30256), .ZN(n25422) );
  NAND2_X1 U33906 ( .A1(n52144), .A2(n6486), .ZN(n27914) );
  NAND3_X1 U33907 ( .A1(n25422), .A2(n52102), .A3(n27914), .ZN(n25854) );
  XNOR2_X1 U33908 ( .A(n369), .B(n25915), .ZN(n25423) );
  INV_X1 U33909 ( .A(n37473), .ZN(n41852) );
  XNOR2_X1 U33910 ( .A(n25747), .B(n41852), .ZN(n25424) );
  XNOR2_X1 U33911 ( .A(n25424), .B(n26044), .ZN(n25425) );
  INV_X1 U33912 ( .A(n37476), .ZN(n25427) );
  XNOR2_X1 U33913 ( .A(n25743), .B(n25426), .ZN(n42996) );
  XNOR2_X1 U33914 ( .A(n25427), .B(n42996), .ZN(n25428) );
  XNOR2_X1 U33915 ( .A(n25429), .B(n25428), .ZN(n25430) );
  XNOR2_X1 U33916 ( .A(n25917), .B(n25431), .ZN(n25432) );
  XNOR2_X1 U33917 ( .A(n27463), .B(n25432), .ZN(n25433) );
  XNOR2_X1 U33918 ( .A(n25433), .B(n25600), .ZN(n29278) );
  INV_X1 U33919 ( .A(n25434), .ZN(n25435) );
  XNOR2_X1 U33920 ( .A(n49937), .B(n4535), .ZN(n26404) );
  XNOR2_X1 U33921 ( .A(n25435), .B(n26404), .ZN(n44523) );
  XNOR2_X1 U33922 ( .A(n25436), .B(n4744), .ZN(n25437) );
  XNOR2_X1 U33923 ( .A(n25437), .B(n45051), .ZN(n42226) );
  XNOR2_X1 U33924 ( .A(n44523), .B(n42226), .ZN(n25438) );
  XNOR2_X1 U33925 ( .A(n25548), .B(n25438), .ZN(n25439) );
  XNOR2_X1 U33926 ( .A(n471), .B(n25439), .ZN(n25441) );
  XNOR2_X1 U33927 ( .A(n25821), .B(n25442), .ZN(n25443) );
  XNOR2_X1 U33928 ( .A(n25445), .B(n25444), .ZN(n25447) );
  XNOR2_X1 U33929 ( .A(n25447), .B(n25446), .ZN(n25449) );
  XNOR2_X1 U33930 ( .A(n25448), .B(n25449), .ZN(n25451) );
  XNOR2_X1 U33931 ( .A(n25450), .B(n25451), .ZN(n25452) );
  XNOR2_X1 U33932 ( .A(n25453), .B(n25452), .ZN(n29191) );
  AND2_X1 U33933 ( .A1(n29278), .A2(n29191), .ZN(n29283) );
  XNOR2_X1 U33934 ( .A(n25792), .B(n4755), .ZN(n38859) );
  XNOR2_X1 U33935 ( .A(n38859), .B(n4482), .ZN(n25454) );
  XNOR2_X1 U33936 ( .A(n43054), .B(n38626), .ZN(n31808) );
  XNOR2_X1 U33937 ( .A(n25454), .B(n31808), .ZN(n25455) );
  XNOR2_X1 U33938 ( .A(n25455), .B(n29661), .ZN(n25456) );
  XNOR2_X1 U33939 ( .A(n27374), .B(n25456), .ZN(n25459) );
  XNOR2_X1 U33940 ( .A(n25457), .B(n26378), .ZN(n25458) );
  XNOR2_X1 U33941 ( .A(n25459), .B(n25458), .ZN(n25460) );
  XNOR2_X1 U33942 ( .A(n25461), .B(n25460), .ZN(n25462) );
  XNOR2_X1 U33943 ( .A(n25464), .B(n25947), .ZN(n25465) );
  XNOR2_X1 U33946 ( .A(n25468), .B(n26358), .ZN(n37141) );
  XNOR2_X1 U33947 ( .A(n37141), .B(n4316), .ZN(n42936) );
  XNOR2_X1 U33948 ( .A(n4883), .B(n4896), .ZN(n25940) );
  XNOR2_X1 U33949 ( .A(n25940), .B(n4213), .ZN(n25469) );
  XNOR2_X1 U33950 ( .A(n25470), .B(n25469), .ZN(n40221) );
  XNOR2_X1 U33951 ( .A(n40221), .B(n4666), .ZN(n25471) );
  XNOR2_X1 U33952 ( .A(n42936), .B(n25471), .ZN(n25472) );
  XNOR2_X1 U33953 ( .A(n26573), .B(n25472), .ZN(n25473) );
  XNOR2_X1 U33954 ( .A(n25473), .B(n51667), .ZN(n25474) );
  XNOR2_X1 U33955 ( .A(n25475), .B(n25474), .ZN(n25476) );
  XNOR2_X1 U33956 ( .A(n25477), .B(n25476), .ZN(n25478) );
  NOR2_X1 U33957 ( .A1(n29183), .A2(n51116), .ZN(n25492) );
  XNOR2_X1 U33958 ( .A(n42258), .B(n44493), .ZN(n26445) );
  XNOR2_X1 U33959 ( .A(n44495), .B(n26445), .ZN(n25480) );
  XNOR2_X1 U33960 ( .A(n25481), .B(n25480), .ZN(n25482) );
  XNOR2_X1 U33961 ( .A(n25482), .B(n26610), .ZN(n25484) );
  XNOR2_X1 U33962 ( .A(n25483), .B(n4065), .ZN(n26612) );
  XNOR2_X1 U33963 ( .A(n25484), .B(n26612), .ZN(n25489) );
  XNOR2_X1 U33964 ( .A(n25775), .B(n42329), .ZN(n25612) );
  XNOR2_X1 U33965 ( .A(n25612), .B(n25485), .ZN(n25487) );
  XNOR2_X1 U33966 ( .A(n51648), .B(n27322), .ZN(n25486) );
  XNOR2_X1 U33967 ( .A(n25486), .B(n28353), .ZN(n25777) );
  XNOR2_X1 U33968 ( .A(n25487), .B(n25777), .ZN(n25488) );
  XNOR2_X1 U33969 ( .A(n25489), .B(n25488), .ZN(n25490) );
  OAI21_X1 U33970 ( .B1(n29181), .B2(n25492), .A(n377), .ZN(n25519) );
  XNOR2_X1 U33971 ( .A(n25755), .B(n25495), .ZN(n25496) );
  INV_X1 U33972 ( .A(n33749), .ZN(n25497) );
  XNOR2_X1 U33973 ( .A(n25497), .B(n48814), .ZN(n42496) );
  XNOR2_X1 U33974 ( .A(n33474), .B(n4654), .ZN(n25498) );
  XNOR2_X1 U33975 ( .A(n43766), .B(n25498), .ZN(n25499) );
  XNOR2_X1 U33976 ( .A(n42496), .B(n25499), .ZN(n25500) );
  XNOR2_X1 U33977 ( .A(n25501), .B(n25500), .ZN(n25502) );
  XNOR2_X1 U33978 ( .A(n25502), .B(n27291), .ZN(n25503) );
  XNOR2_X1 U33979 ( .A(n25352), .B(n26239), .ZN(n28083) );
  XNOR2_X1 U33980 ( .A(n28083), .B(n25505), .ZN(n25512) );
  INV_X1 U33981 ( .A(n25506), .ZN(n25507) );
  XNOR2_X1 U33982 ( .A(n25508), .B(n25507), .ZN(n25509) );
  XNOR2_X1 U33983 ( .A(n25509), .B(n25510), .ZN(n26417) );
  XNOR2_X1 U33984 ( .A(n26417), .B(n28218), .ZN(n25511) );
  OAI211_X1 U33985 ( .C1(n5656), .C2(n51116), .A(n29190), .B(n28710), .ZN(
        n25513) );
  MUX2_X1 U33986 ( .A(n25513), .B(n28708), .S(n51706), .Z(n25518) );
  NOR2_X1 U33987 ( .A1(n28715), .A2(n377), .ZN(n25515) );
  NAND2_X1 U33988 ( .A1(n29269), .A2(n27780), .ZN(n25514) );
  AND2_X1 U33989 ( .A1(n29187), .A2(n27780), .ZN(n25516) );
  XNOR2_X1 U33990 ( .A(n27289), .B(n28093), .ZN(n25527) );
  INV_X1 U33991 ( .A(n43592), .ZN(n25523) );
  XNOR2_X1 U33992 ( .A(n25521), .B(n25520), .ZN(n42710) );
  XNOR2_X1 U33993 ( .A(n42710), .B(n43586), .ZN(n25522) );
  XNOR2_X1 U33994 ( .A(n25523), .B(n25522), .ZN(n25524) );
  XNOR2_X1 U33995 ( .A(n25755), .B(n25524), .ZN(n25525) );
  XNOR2_X1 U33996 ( .A(n23621), .B(n25525), .ZN(n25526) );
  XNOR2_X1 U33997 ( .A(n25527), .B(n25526), .ZN(n25528) );
  XNOR2_X1 U33998 ( .A(n25529), .B(n25528), .ZN(n25535) );
  XNOR2_X1 U33999 ( .A(n27309), .B(n26435), .ZN(n25530) );
  XNOR2_X1 U34000 ( .A(n25530), .B(n25762), .ZN(n25531) );
  XNOR2_X1 U34001 ( .A(n28221), .B(n25664), .ZN(n26250) );
  XNOR2_X1 U34002 ( .A(n26250), .B(n25531), .ZN(n25532) );
  XNOR2_X1 U34003 ( .A(n25532), .B(n25533), .ZN(n25534) );
  XNOR2_X1 U34004 ( .A(n25534), .B(n25535), .ZN(n25603) );
  XNOR2_X1 U34005 ( .A(n45401), .B(n4286), .ZN(n25536) );
  XNOR2_X1 U34006 ( .A(n25537), .B(n25536), .ZN(n42356) );
  XNOR2_X1 U34007 ( .A(n25538), .B(n4890), .ZN(n45052) );
  XNOR2_X1 U34008 ( .A(n42356), .B(n45052), .ZN(n25539) );
  XNOR2_X1 U34009 ( .A(n25540), .B(n25539), .ZN(n25541) );
  XNOR2_X1 U34010 ( .A(n25541), .B(n25903), .ZN(n25543) );
  XNOR2_X1 U34011 ( .A(n27501), .B(n26402), .ZN(n25545) );
  XNOR2_X1 U34012 ( .A(n26053), .B(n25545), .ZN(n25546) );
  XNOR2_X1 U34013 ( .A(n2212), .B(n25546), .ZN(n27344) );
  XNOR2_X1 U34014 ( .A(n25547), .B(n27344), .ZN(n25552) );
  XNOR2_X1 U34015 ( .A(n28288), .B(n25548), .ZN(n25549) );
  XNOR2_X1 U34016 ( .A(n25549), .B(n26530), .ZN(n27347) );
  XNOR2_X1 U34017 ( .A(n27347), .B(n4781), .ZN(n25650) );
  XNOR2_X1 U34018 ( .A(n25650), .B(n25550), .ZN(n25551) );
  NAND2_X1 U34019 ( .A1(n25603), .A2(n29247), .ZN(n29120) );
  INV_X1 U34020 ( .A(n29120), .ZN(n27938) );
  XNOR2_X1 U34021 ( .A(n25691), .B(n25553), .ZN(n25950) );
  XNOR2_X1 U34022 ( .A(n27218), .B(n25950), .ZN(n25568) );
  XNOR2_X1 U34023 ( .A(n51666), .B(n25554), .ZN(n25562) );
  XNOR2_X1 U34024 ( .A(n42084), .B(n25555), .ZN(n25559) );
  XNOR2_X1 U34025 ( .A(n33733), .B(n4045), .ZN(n25556) );
  INV_X1 U34026 ( .A(n41155), .ZN(n41835) );
  XNOR2_X1 U34027 ( .A(n25556), .B(n41835), .ZN(n25557) );
  XNOR2_X1 U34028 ( .A(n25557), .B(n42102), .ZN(n25558) );
  XNOR2_X1 U34029 ( .A(n25559), .B(n25558), .ZN(n25560) );
  XNOR2_X1 U34030 ( .A(n26285), .B(n25560), .ZN(n25561) );
  XNOR2_X1 U34031 ( .A(n25562), .B(n25561), .ZN(n25564) );
  XNOR2_X1 U34032 ( .A(n26565), .B(n25947), .ZN(n25563) );
  XNOR2_X1 U34033 ( .A(n25564), .B(n26009), .ZN(n25565) );
  XNOR2_X1 U34034 ( .A(n25566), .B(n25565), .ZN(n25567) );
  XNOR2_X1 U34035 ( .A(n25570), .B(n25569), .ZN(n25802) );
  XNOR2_X1 U34036 ( .A(n25571), .B(n27222), .ZN(n25573) );
  XNOR2_X1 U34037 ( .A(n27368), .B(n27362), .ZN(n25572) );
  XNOR2_X1 U34038 ( .A(n25573), .B(n25572), .ZN(n25585) );
  XNOR2_X1 U34039 ( .A(n25798), .B(n25574), .ZN(n25583) );
  XNOR2_X1 U34040 ( .A(n25576), .B(n25575), .ZN(n44328) );
  XNOR2_X1 U34041 ( .A(n26297), .B(n4542), .ZN(n25577) );
  XNOR2_X1 U34042 ( .A(n25578), .B(n25577), .ZN(n46064) );
  XNOR2_X1 U34043 ( .A(n4597), .B(n4490), .ZN(n33652) );
  XNOR2_X1 U34044 ( .A(n46064), .B(n33652), .ZN(n25579) );
  XNOR2_X1 U34045 ( .A(n44328), .B(n25579), .ZN(n25580) );
  XNOR2_X1 U34046 ( .A(n27374), .B(n25580), .ZN(n25581) );
  XNOR2_X1 U34047 ( .A(n26300), .B(n25581), .ZN(n25582) );
  XNOR2_X1 U34048 ( .A(n25583), .B(n25582), .ZN(n25584) );
  XNOR2_X1 U34049 ( .A(n25585), .B(n25584), .ZN(n25586) );
  XNOR2_X1 U34050 ( .A(n25802), .B(n25586), .ZN(n30233) );
  XNOR2_X1 U34051 ( .A(n25927), .B(n42339), .ZN(n25587) );
  XNOR2_X1 U34052 ( .A(n25587), .B(n27177), .ZN(n25588) );
  XNOR2_X1 U34053 ( .A(n2209), .B(n25588), .ZN(n25752) );
  INV_X1 U34054 ( .A(n25589), .ZN(n25921) );
  XNOR2_X1 U34055 ( .A(n25590), .B(n25921), .ZN(n25591) );
  XNOR2_X1 U34056 ( .A(n25752), .B(n25591), .ZN(n27381) );
  XNOR2_X1 U34057 ( .A(n46097), .B(n41852), .ZN(n25592) );
  XNOR2_X1 U34058 ( .A(n27454), .B(n4624), .ZN(n44293) );
  XNOR2_X1 U34059 ( .A(n25592), .B(n44293), .ZN(n25593) );
  XNOR2_X1 U34060 ( .A(n26210), .B(n25593), .ZN(n25594) );
  XNOR2_X1 U34061 ( .A(n28311), .B(n25594), .ZN(n25597) );
  INV_X1 U34062 ( .A(n25747), .ZN(n25595) );
  XNOR2_X1 U34063 ( .A(n27451), .B(n25595), .ZN(n25596) );
  XNOR2_X1 U34064 ( .A(n25597), .B(n25596), .ZN(n25598) );
  XNOR2_X1 U34065 ( .A(n25598), .B(n28101), .ZN(n25599) );
  XNOR2_X1 U34066 ( .A(n27381), .B(n25599), .ZN(n25602) );
  INV_X1 U34067 ( .A(n25600), .ZN(n25601) );
  XNOR2_X1 U34068 ( .A(n750), .B(n25604), .ZN(n25607) );
  XNOR2_X1 U34069 ( .A(n28238), .B(n25605), .ZN(n25606) );
  XNOR2_X1 U34070 ( .A(n25607), .B(n25606), .ZN(n27314) );
  XNOR2_X1 U34071 ( .A(n25609), .B(n25608), .ZN(n25611) );
  XNOR2_X1 U34072 ( .A(n25611), .B(n25610), .ZN(n25774) );
  XNOR2_X1 U34073 ( .A(n27314), .B(n25774), .ZN(n25625) );
  INV_X1 U34074 ( .A(n25612), .ZN(n25614) );
  XNOR2_X1 U34075 ( .A(n25614), .B(n25613), .ZN(n25621) );
  XNOR2_X1 U34076 ( .A(n28069), .B(n26610), .ZN(n25619) );
  XNOR2_X1 U34077 ( .A(n25615), .B(n4691), .ZN(n45087) );
  XNOR2_X1 U34078 ( .A(n45087), .B(n25616), .ZN(n25617) );
  XNOR2_X1 U34079 ( .A(n51009), .B(n25617), .ZN(n25618) );
  XNOR2_X1 U34080 ( .A(n25619), .B(n25618), .ZN(n25620) );
  XNOR2_X1 U34081 ( .A(n25621), .B(n25620), .ZN(n25623) );
  XNOR2_X1 U34082 ( .A(n25882), .B(n27479), .ZN(n25622) );
  XNOR2_X1 U34083 ( .A(n25623), .B(n25622), .ZN(n25624) );
  XNOR2_X1 U34084 ( .A(n25625), .B(n25624), .ZN(n25626) );
  INV_X1 U34085 ( .A(n29247), .ZN(n28650) );
  OAI21_X1 U34086 ( .B1(n30233), .B2(n29252), .A(n28650), .ZN(n25627) );
  NAND2_X1 U34087 ( .A1(n29123), .A2(n29259), .ZN(n27936) );
  OAI211_X1 U34088 ( .C1(n30232), .C2(n4724), .A(n25627), .B(n27936), .ZN(
        n25628) );
  INV_X1 U34089 ( .A(n25628), .ZN(n25629) );
  NAND2_X1 U34091 ( .A1(n28658), .A2(n30226), .ZN(n30220) );
  NAND2_X1 U34092 ( .A1(n29260), .A2(n29259), .ZN(n25634) );
  OAI21_X1 U34093 ( .B1(n28658), .B2(n29120), .A(n29249), .ZN(n25631) );
  NAND2_X1 U34094 ( .A1(n25631), .A2(n29259), .ZN(n25633) );
  AND2_X1 U34095 ( .A1(n28650), .A2(n29123), .ZN(n29119) );
  OAI211_X1 U34096 ( .C1(n30220), .C2(n25634), .A(n25633), .B(n25632), .ZN(
        n25635) );
  INV_X1 U34097 ( .A(n25635), .ZN(n25849) );
  AND2_X1 U34098 ( .A1(n30226), .A2(n28650), .ZN(n30235) );
  NAND2_X1 U34099 ( .A1(n28658), .A2(n29263), .ZN(n29255) );
  NAND3_X1 U34100 ( .A1(n29264), .A2(n30226), .A3(n30232), .ZN(n25636) );
  AND2_X1 U34101 ( .A1(n25637), .A2(n25636), .ZN(n25850) );
  AND2_X1 U34102 ( .A1(n29260), .A2(n29247), .ZN(n30228) );
  XNOR2_X1 U34103 ( .A(n25915), .B(n25921), .ZN(n28319) );
  XNOR2_X1 U34104 ( .A(n26044), .B(n44909), .ZN(n26096) );
  XNOR2_X1 U34105 ( .A(n28309), .B(n25640), .ZN(n43221) );
  XNOR2_X1 U34106 ( .A(n25641), .B(n4746), .ZN(n25642) );
  XNOR2_X1 U34107 ( .A(n43221), .B(n25642), .ZN(n25643) );
  XNOR2_X1 U34108 ( .A(n25920), .B(n25643), .ZN(n25644) );
  XNOR2_X1 U34109 ( .A(n26096), .B(n25644), .ZN(n25645) );
  XNOR2_X1 U34110 ( .A(n25645), .B(n27445), .ZN(n25648) );
  XNOR2_X1 U34111 ( .A(n28311), .B(n25646), .ZN(n25647) );
  XNOR2_X1 U34112 ( .A(n25647), .B(n370), .ZN(n26051) );
  XNOR2_X1 U34113 ( .A(n25648), .B(n26051), .ZN(n25649) );
  XNOR2_X1 U34114 ( .A(n28297), .B(n25650), .ZN(n25663) );
  XNOR2_X1 U34115 ( .A(n26053), .B(n25829), .ZN(n25659) );
  INV_X1 U34116 ( .A(n25651), .ZN(n25653) );
  XNOR2_X1 U34117 ( .A(n27186), .B(n33221), .ZN(n25652) );
  XNOR2_X1 U34118 ( .A(n25653), .B(n25652), .ZN(n43621) );
  XNOR2_X1 U34119 ( .A(n2602), .B(n4826), .ZN(n25654) );
  XNOR2_X1 U34120 ( .A(n25655), .B(n25654), .ZN(n42722) );
  XNOR2_X1 U34121 ( .A(n43621), .B(n42722), .ZN(n25656) );
  XNOR2_X1 U34122 ( .A(n28287), .B(n25656), .ZN(n25657) );
  XNOR2_X1 U34123 ( .A(n25657), .B(n26529), .ZN(n25658) );
  XNOR2_X1 U34124 ( .A(n25659), .B(n25658), .ZN(n25661) );
  XNOR2_X1 U34125 ( .A(n25661), .B(n25660), .ZN(n25662) );
  XNOR2_X1 U34126 ( .A(n25663), .B(n25662), .ZN(n26083) );
  XNOR2_X1 U34127 ( .A(n25665), .B(n28223), .ZN(n25754) );
  XNOR2_X1 U34128 ( .A(n49109), .B(n4048), .ZN(n34136) );
  XNOR2_X1 U34129 ( .A(n43878), .B(n34136), .ZN(n25757) );
  XNOR2_X1 U34130 ( .A(n27297), .B(n4526), .ZN(n25666) );
  XNOR2_X1 U34131 ( .A(n25757), .B(n25666), .ZN(n25667) );
  XNOR2_X1 U34132 ( .A(n45478), .B(n25667), .ZN(n25668) );
  XNOR2_X1 U34133 ( .A(n25669), .B(n25668), .ZN(n25670) );
  XNOR2_X1 U34134 ( .A(n25670), .B(n27291), .ZN(n25671) );
  XNOR2_X1 U34135 ( .A(n24814), .B(n25671), .ZN(n25672) );
  XNOR2_X1 U34136 ( .A(n25754), .B(n25672), .ZN(n25679) );
  XNOR2_X1 U34137 ( .A(n2080), .B(n4613), .ZN(n25674) );
  XNOR2_X1 U34138 ( .A(n25673), .B(n25674), .ZN(n25676) );
  INV_X1 U34139 ( .A(n26235), .ZN(n25675) );
  XNOR2_X1 U34140 ( .A(n25675), .B(n25676), .ZN(n26021) );
  XNOR2_X1 U34141 ( .A(n26021), .B(n25677), .ZN(n25678) );
  XNOR2_X1 U34142 ( .A(n25679), .B(n25678), .ZN(n25734) );
  OR2_X1 U34143 ( .A1(n29305), .A2(n29309), .ZN(n26659) );
  XNOR2_X1 U34144 ( .A(n25681), .B(n25680), .ZN(n28369) );
  XNOR2_X1 U34145 ( .A(n25682), .B(n28049), .ZN(n25690) );
  INV_X1 U34146 ( .A(n43371), .ZN(n25684) );
  XNOR2_X1 U34147 ( .A(n25684), .B(n25683), .ZN(n35113) );
  XNOR2_X1 U34148 ( .A(n43369), .B(n25685), .ZN(n25686) );
  XNOR2_X1 U34149 ( .A(n25686), .B(n33295), .ZN(n25687) );
  XNOR2_X1 U34150 ( .A(n35113), .B(n25687), .ZN(n25688) );
  XNOR2_X1 U34151 ( .A(n51751), .B(n25688), .ZN(n25689) );
  XNOR2_X1 U34152 ( .A(n25690), .B(n25689), .ZN(n25693) );
  INV_X1 U34153 ( .A(n25691), .ZN(n25692) );
  XNOR2_X1 U34154 ( .A(n25693), .B(n25692), .ZN(n25694) );
  XNOR2_X1 U34155 ( .A(n28369), .B(n25694), .ZN(n25697) );
  INV_X1 U34156 ( .A(n25695), .ZN(n25696) );
  XNOR2_X1 U34157 ( .A(n25697), .B(n25696), .ZN(n25698) );
  XNOR2_X1 U34158 ( .A(n25700), .B(n25882), .ZN(n25701) );
  XNOR2_X1 U34159 ( .A(n25702), .B(n25701), .ZN(n25704) );
  XNOR2_X1 U34160 ( .A(n26187), .B(n25703), .ZN(n26035) );
  XNOR2_X1 U34161 ( .A(n25704), .B(n26035), .ZN(n25714) );
  INV_X1 U34162 ( .A(n33899), .ZN(n36946) );
  XNOR2_X1 U34163 ( .A(n36946), .B(n34816), .ZN(n33420) );
  XNOR2_X1 U34164 ( .A(n25705), .B(n4908), .ZN(n43605) );
  XNOR2_X1 U34165 ( .A(n43605), .B(n34232), .ZN(n25706) );
  XNOR2_X1 U34166 ( .A(n33420), .B(n25706), .ZN(n25707) );
  XNOR2_X1 U34167 ( .A(n28238), .B(n25707), .ZN(n25709) );
  XNOR2_X1 U34168 ( .A(n25709), .B(n25708), .ZN(n25710) );
  XNOR2_X1 U34169 ( .A(n25777), .B(n25710), .ZN(n25711) );
  XNOR2_X1 U34170 ( .A(n25712), .B(n25711), .ZN(n25713) );
  XNOR2_X1 U34172 ( .A(n25715), .B(n51416), .ZN(n28265) );
  XNOR2_X1 U34173 ( .A(n28265), .B(n27491), .ZN(n25716) );
  XNOR2_X1 U34174 ( .A(n25716), .B(n25717), .ZN(n25732) );
  XNOR2_X1 U34175 ( .A(n25718), .B(n27483), .ZN(n25719) );
  XNOR2_X1 U34176 ( .A(n25720), .B(n25719), .ZN(n43191) );
  XNOR2_X1 U34177 ( .A(n27364), .B(n4515), .ZN(n25721) );
  XNOR2_X1 U34178 ( .A(n25722), .B(n25721), .ZN(n42123) );
  XNOR2_X1 U34179 ( .A(n43191), .B(n42123), .ZN(n25723) );
  XNOR2_X1 U34180 ( .A(n25724), .B(n25723), .ZN(n25725) );
  XNOR2_X1 U34181 ( .A(n25726), .B(n25725), .ZN(n25728) );
  XNOR2_X1 U34182 ( .A(n25728), .B(n25727), .ZN(n25730) );
  XNOR2_X1 U34183 ( .A(n25729), .B(n25730), .ZN(n25731) );
  NAND2_X1 U34184 ( .A1(n28695), .A2(n26651), .ZN(n28701) );
  NAND2_X1 U34185 ( .A1(n29309), .A2(n26083), .ZN(n26650) );
  NAND2_X1 U34186 ( .A1(n29300), .A2(n28690), .ZN(n25733) );
  OAI21_X1 U34187 ( .B1(n28701), .B2(n28699), .A(n51517), .ZN(n25736) );
  NAND2_X1 U34189 ( .A1(n28690), .A2(n29290), .ZN(n28700) );
  AOI21_X1 U34190 ( .B1(n28700), .B2(n27844), .A(n27847), .ZN(n25735) );
  NAND2_X1 U34191 ( .A1(n31873), .A2(n31883), .ZN(n31020) );
  XNOR2_X1 U34192 ( .A(n25738), .B(n25737), .ZN(n25739) );
  XNOR2_X1 U34193 ( .A(n28311), .B(n25740), .ZN(n25741) );
  XNOR2_X1 U34194 ( .A(n25742), .B(n25741), .ZN(n25750) );
  XNOR2_X1 U34195 ( .A(n25743), .B(n4723), .ZN(n42909) );
  XNOR2_X1 U34196 ( .A(n25744), .B(n4939), .ZN(n25745) );
  XNOR2_X1 U34197 ( .A(n27390), .B(n25745), .ZN(n40758) );
  XNOR2_X1 U34198 ( .A(n42909), .B(n40758), .ZN(n25746) );
  XNOR2_X1 U34199 ( .A(n25747), .B(n25746), .ZN(n25748) );
  XNOR2_X1 U34200 ( .A(n25748), .B(n26395), .ZN(n25749) );
  XNOR2_X1 U34201 ( .A(n25750), .B(n25749), .ZN(n25751) );
  XNOR2_X1 U34202 ( .A(n27382), .B(n4800), .ZN(n25916) );
  XNOR2_X1 U34203 ( .A(n25916), .B(n26100), .ZN(n28109) );
  XNOR2_X1 U34204 ( .A(n25752), .B(n28109), .ZN(n25753) );
  INV_X1 U34205 ( .A(n25754), .ZN(n25767) );
  XNOR2_X1 U34206 ( .A(n25756), .B(n28214), .ZN(n26238) );
  XNOR2_X1 U34207 ( .A(n27299), .B(n25866), .ZN(n25758) );
  XNOR2_X1 U34208 ( .A(n25758), .B(n25757), .ZN(n43500) );
  XNOR2_X1 U34209 ( .A(n43500), .B(n44161), .ZN(n25759) );
  XNOR2_X1 U34210 ( .A(n26589), .B(n25759), .ZN(n25760) );
  XNOR2_X1 U34211 ( .A(n26238), .B(n25761), .ZN(n25765) );
  XNOR2_X1 U34212 ( .A(n25762), .B(n25763), .ZN(n25764) );
  XNOR2_X1 U34213 ( .A(n25765), .B(n25764), .ZN(n25766) );
  XNOR2_X1 U34214 ( .A(n25767), .B(n25766), .ZN(n25769) );
  XNOR2_X1 U34215 ( .A(n25769), .B(n25768), .ZN(n25789) );
  XNOR2_X1 U34217 ( .A(n750), .B(n51720), .ZN(n25773) );
  XNOR2_X1 U34218 ( .A(n25773), .B(n25772), .ZN(n26256) );
  XNOR2_X1 U34219 ( .A(n25774), .B(n26256), .ZN(n25788) );
  XNOR2_X1 U34220 ( .A(n25775), .B(n4655), .ZN(n25776) );
  XNOR2_X1 U34221 ( .A(n25776), .B(n26600), .ZN(n25886) );
  XNOR2_X1 U34222 ( .A(n25886), .B(n25777), .ZN(n25786) );
  XNOR2_X1 U34223 ( .A(n25778), .B(n4895), .ZN(n26183) );
  INV_X1 U34224 ( .A(n25779), .ZN(n25780) );
  XNOR2_X1 U34225 ( .A(n27317), .B(n25780), .ZN(n43730) );
  XNOR2_X1 U34226 ( .A(n28071), .B(n45348), .ZN(n25781) );
  XNOR2_X1 U34227 ( .A(n25781), .B(n43739), .ZN(n25782) );
  XNOR2_X1 U34228 ( .A(n43730), .B(n25782), .ZN(n25783) );
  XNOR2_X1 U34229 ( .A(n26183), .B(n25783), .ZN(n25784) );
  XNOR2_X1 U34230 ( .A(n51750), .B(n25784), .ZN(n25785) );
  XNOR2_X1 U34231 ( .A(n25786), .B(n25785), .ZN(n25787) );
  XNOR2_X2 U34232 ( .A(n25788), .B(n25787), .ZN(n26668) );
  XNOR2_X1 U34233 ( .A(n27363), .B(n25790), .ZN(n25800) );
  XNOR2_X1 U34234 ( .A(n25791), .B(n28266), .ZN(n33651) );
  XNOR2_X1 U34235 ( .A(n25793), .B(n25792), .ZN(n25794) );
  XNOR2_X1 U34236 ( .A(n33651), .B(n25794), .ZN(n40521) );
  XNOR2_X1 U34237 ( .A(n25795), .B(n2947), .ZN(n42946) );
  XNOR2_X1 U34238 ( .A(n40521), .B(n42946), .ZN(n25796) );
  XNOR2_X1 U34239 ( .A(n27232), .B(n25796), .ZN(n25797) );
  XNOR2_X1 U34240 ( .A(n25798), .B(n25797), .ZN(n25799) );
  XNOR2_X1 U34241 ( .A(n25800), .B(n25799), .ZN(n25801) );
  NAND3_X1 U34242 ( .A1(n28669), .A2(n26668), .A3(n28666), .ZN(n26666) );
  XNOR2_X1 U34243 ( .A(n25805), .B(n28246), .ZN(n25808) );
  XNOR2_X1 U34244 ( .A(n25806), .B(n25934), .ZN(n25807) );
  XNOR2_X1 U34245 ( .A(n25807), .B(n25808), .ZN(n25820) );
  XNOR2_X1 U34246 ( .A(n26285), .B(n28370), .ZN(n25815) );
  XNOR2_X1 U34247 ( .A(n28375), .B(n25939), .ZN(n25810) );
  XNOR2_X1 U34248 ( .A(n43927), .B(n2599), .ZN(n25809) );
  XNOR2_X1 U34249 ( .A(n25810), .B(n25809), .ZN(n25811) );
  XNOR2_X1 U34250 ( .A(n25811), .B(n43654), .ZN(n25812) );
  XNOR2_X1 U34251 ( .A(n25813), .B(n25812), .ZN(n25814) );
  XNOR2_X1 U34252 ( .A(n25815), .B(n25814), .ZN(n25818) );
  XNOR2_X1 U34253 ( .A(n26272), .B(n25816), .ZN(n25817) );
  XNOR2_X1 U34254 ( .A(n25818), .B(n25817), .ZN(n25819) );
  XNOR2_X1 U34255 ( .A(n51752), .B(n2125), .ZN(n25828) );
  XNOR2_X1 U34256 ( .A(n34865), .B(n4826), .ZN(n42409) );
  XNOR2_X1 U34257 ( .A(n26057), .B(n25822), .ZN(n43712) );
  XNOR2_X1 U34258 ( .A(n43712), .B(n2604), .ZN(n25823) );
  XNOR2_X1 U34259 ( .A(n42409), .B(n25823), .ZN(n25824) );
  XNOR2_X1 U34260 ( .A(n25825), .B(n25824), .ZN(n25826) );
  XNOR2_X1 U34261 ( .A(n25826), .B(n26119), .ZN(n25827) );
  XNOR2_X1 U34262 ( .A(n25828), .B(n25827), .ZN(n25830) );
  INV_X1 U34263 ( .A(n28126), .ZN(n26220) );
  XNOR2_X1 U34264 ( .A(n25829), .B(n26220), .ZN(n25907) );
  XNOR2_X1 U34265 ( .A(n25830), .B(n25907), .ZN(n25835) );
  XNOR2_X1 U34266 ( .A(n25832), .B(n25831), .ZN(n28402) );
  XNOR2_X1 U34267 ( .A(n25833), .B(n28402), .ZN(n25834) );
  NAND3_X1 U34268 ( .A1(n27859), .A2(n3124), .A3(n26671), .ZN(n25839) );
  XNOR2_X1 U34269 ( .A(n27852), .B(n28669), .ZN(n25837) );
  OAI211_X1 U34270 ( .C1(n29478), .C2(n26676), .A(n28671), .B(n25837), .ZN(
        n25838) );
  INV_X1 U34271 ( .A(n29498), .ZN(n25843) );
  OAI21_X1 U34272 ( .B1(n25843), .B2(n25842), .A(n2294), .ZN(n25845) );
  NAND2_X1 U34273 ( .A1(n27860), .A2(n28666), .ZN(n29480) );
  NAND2_X1 U34274 ( .A1(n29496), .A2(n29480), .ZN(n25844) );
  NOR2_X1 U34275 ( .A1(n31020), .A2(n28489), .ZN(n25847) );
  NAND4_X1 U34276 ( .A1(n25851), .A2(n25850), .A3(n25849), .A4(n25848), .ZN(
        n25857) );
  INV_X1 U34277 ( .A(n25852), .ZN(n25856) );
  NAND2_X1 U34278 ( .A1(n25854), .A2(n25853), .ZN(n25855) );
  NOR3_X1 U34279 ( .A1(n25857), .A2(n25856), .A3(n25855), .ZN(n25858) );
  XNOR2_X1 U34280 ( .A(n26235), .B(n25859), .ZN(n25862) );
  XNOR2_X1 U34281 ( .A(n25860), .B(n26581), .ZN(n25861) );
  XNOR2_X1 U34282 ( .A(n25862), .B(n25861), .ZN(n25863) );
  XNOR2_X1 U34283 ( .A(n25864), .B(n25863), .ZN(n25875) );
  XNOR2_X1 U34284 ( .A(n27290), .B(n25865), .ZN(n25873) );
  XNOR2_X1 U34285 ( .A(n45335), .B(n25866), .ZN(n25868) );
  XNOR2_X1 U34286 ( .A(n44952), .B(n4486), .ZN(n27434) );
  XNOR2_X1 U34287 ( .A(n27434), .B(n49109), .ZN(n45479) );
  XNOR2_X1 U34288 ( .A(n26586), .B(n4687), .ZN(n25867) );
  XNOR2_X1 U34289 ( .A(n45479), .B(n25867), .ZN(n43988) );
  XNOR2_X1 U34290 ( .A(n25868), .B(n43988), .ZN(n25869) );
  XNOR2_X1 U34291 ( .A(n25870), .B(n27291), .ZN(n25871) );
  XNOR2_X1 U34292 ( .A(n25871), .B(n27256), .ZN(n25872) );
  XNOR2_X1 U34293 ( .A(n25873), .B(n25872), .ZN(n25874) );
  INV_X1 U34294 ( .A(n44090), .ZN(n25878) );
  XOR2_X1 U34295 ( .A(n4065), .B(n4836), .Z(n25876) );
  XNOR2_X1 U34296 ( .A(n26180), .B(n25876), .ZN(n25877) );
  XNOR2_X1 U34297 ( .A(n25878), .B(n25877), .ZN(n25879) );
  XNOR2_X1 U34298 ( .A(n27272), .B(n25879), .ZN(n25880) );
  XNOR2_X1 U34299 ( .A(n25881), .B(n25880), .ZN(n25885) );
  XNOR2_X1 U34300 ( .A(n25883), .B(n25882), .ZN(n25884) );
  XNOR2_X1 U34301 ( .A(n25885), .B(n25884), .ZN(n25888) );
  XNOR2_X1 U34302 ( .A(n25888), .B(n25887), .ZN(n25895) );
  XNOR2_X1 U34303 ( .A(n28238), .B(n26264), .ZN(n25890) );
  XNOR2_X1 U34304 ( .A(n25890), .B(n25889), .ZN(n25891) );
  XNOR2_X1 U34305 ( .A(n25892), .B(n25891), .ZN(n27275) );
  XNOR2_X1 U34306 ( .A(n27275), .B(n25893), .ZN(n25894) );
  XNOR2_X1 U34307 ( .A(n25896), .B(n26228), .ZN(n25906) );
  XNOR2_X1 U34308 ( .A(n25897), .B(n32267), .ZN(n25900) );
  XNOR2_X1 U34309 ( .A(n27349), .B(n25898), .ZN(n25899) );
  XNOR2_X1 U34310 ( .A(n25900), .B(n25899), .ZN(n42580) );
  XNOR2_X1 U34311 ( .A(n25901), .B(n3481), .ZN(n44024) );
  XNOR2_X1 U34312 ( .A(n42580), .B(n44024), .ZN(n25902) );
  XNOR2_X1 U34313 ( .A(n28287), .B(n25902), .ZN(n25904) );
  XNOR2_X1 U34314 ( .A(n25903), .B(n25904), .ZN(n25905) );
  XNOR2_X1 U34315 ( .A(n25906), .B(n25905), .ZN(n25908) );
  XNOR2_X1 U34316 ( .A(n25908), .B(n25907), .ZN(n25914) );
  XNOR2_X1 U34317 ( .A(n26529), .B(n26402), .ZN(n25910) );
  XNOR2_X1 U34318 ( .A(n32856), .B(n4487), .ZN(n42575) );
  XNOR2_X1 U34319 ( .A(n25909), .B(n42575), .ZN(n27505) );
  XNOR2_X1 U34320 ( .A(n25910), .B(n27505), .ZN(n25911) );
  XNOR2_X1 U34321 ( .A(n25911), .B(n27347), .ZN(n25912) );
  XNOR2_X1 U34322 ( .A(n26055), .B(n25912), .ZN(n25913) );
  XNOR2_X2 U34323 ( .A(n25913), .B(n25914), .ZN(n29330) );
  INV_X1 U34324 ( .A(n29330), .ZN(n25975) );
  NAND2_X1 U34325 ( .A1(n51107), .A2(n25975), .ZN(n28642) );
  NAND2_X1 U34326 ( .A1(n29331), .A2(n28642), .ZN(n25967) );
  XNOR2_X1 U34327 ( .A(n25916), .B(n25915), .ZN(n25919) );
  INV_X1 U34328 ( .A(n25917), .ZN(n25918) );
  XNOR2_X1 U34329 ( .A(n26508), .B(n26100), .ZN(n25923) );
  XNOR2_X1 U34330 ( .A(n25921), .B(n25920), .ZN(n25922) );
  XNOR2_X1 U34331 ( .A(n25923), .B(n25922), .ZN(n25931) );
  XNOR2_X1 U34332 ( .A(n34744), .B(n25924), .ZN(n43121) );
  XNOR2_X1 U34333 ( .A(n25925), .B(n4076), .ZN(n41843) );
  XNOR2_X1 U34334 ( .A(n43121), .B(n41843), .ZN(n25926) );
  XNOR2_X1 U34335 ( .A(n25927), .B(n25926), .ZN(n25928) );
  XNOR2_X1 U34336 ( .A(n25929), .B(n25928), .ZN(n25930) );
  XNOR2_X1 U34337 ( .A(n25931), .B(n25930), .ZN(n25932) );
  XNOR2_X1 U34338 ( .A(n25937), .B(n28370), .ZN(n25945) );
  XNOR2_X1 U34339 ( .A(n25939), .B(n25938), .ZN(n42823) );
  XNOR2_X1 U34340 ( .A(n44043), .B(n25940), .ZN(n41156) );
  XNOR2_X1 U34341 ( .A(n41156), .B(n1224), .ZN(n25941) );
  XNOR2_X1 U34342 ( .A(n42823), .B(n25941), .ZN(n25942) );
  INV_X1 U34343 ( .A(n41183), .ZN(n26002) );
  XNOR2_X1 U34344 ( .A(n25942), .B(n26002), .ZN(n25943) );
  XNOR2_X1 U34345 ( .A(n27424), .B(n25943), .ZN(n25944) );
  XNOR2_X1 U34346 ( .A(n25945), .B(n25944), .ZN(n25949) );
  XNOR2_X1 U34347 ( .A(n25946), .B(n4431), .ZN(n25948) );
  XNOR2_X1 U34348 ( .A(n25948), .B(n25947), .ZN(n26280) );
  XNOR2_X1 U34349 ( .A(n25949), .B(n26280), .ZN(n25951) );
  XNOR2_X1 U34350 ( .A(n25951), .B(n25950), .ZN(n25952) );
  XNOR2_X1 U34351 ( .A(n25955), .B(n25954), .ZN(n25964) );
  XNOR2_X1 U34352 ( .A(n27232), .B(n4880), .ZN(n28411) );
  XNOR2_X1 U34353 ( .A(n25956), .B(n4578), .ZN(n25958) );
  XNOR2_X1 U34354 ( .A(n25958), .B(n25957), .ZN(n41818) );
  XNOR2_X1 U34355 ( .A(n25959), .B(n4325), .ZN(n43164) );
  XNOR2_X1 U34356 ( .A(n41818), .B(n43164), .ZN(n25960) );
  XNOR2_X1 U34357 ( .A(n28411), .B(n25960), .ZN(n25961) );
  XNOR2_X1 U34358 ( .A(n25962), .B(n25961), .ZN(n25963) );
  NAND3_X1 U34359 ( .A1(n25967), .A2(n52177), .A3(n29315), .ZN(n25971) );
  NAND2_X1 U34360 ( .A1(n29325), .A2(n29330), .ZN(n25968) );
  OR2_X1 U34361 ( .A1(n29331), .A2(n25968), .ZN(n27899) );
  NAND3_X1 U34363 ( .A1(n29317), .A2(n28644), .A3(n29324), .ZN(n25970) );
  INV_X1 U34364 ( .A(n29315), .ZN(n26322) );
  NAND3_X1 U34365 ( .A1(n27897), .A2(n26322), .A3(n29324), .ZN(n25969) );
  NAND2_X1 U34366 ( .A1(n29327), .A2(n29330), .ZN(n29314) );
  NOR2_X1 U34369 ( .A1(n26323), .A2(n459), .ZN(n25972) );
  AOI21_X1 U34370 ( .B1(n27805), .B2(n29317), .A(n25972), .ZN(n25979) );
  AND2_X1 U34371 ( .A1(n29332), .A2(n383), .ZN(n25974) );
  NOR2_X1 U34372 ( .A1(n29332), .A2(n28641), .ZN(n25973) );
  OAI21_X1 U34373 ( .B1(n25974), .B2(n25973), .A(n27818), .ZN(n25978) );
  OAI21_X1 U34374 ( .B1(n27808), .B2(n29324), .A(n29329), .ZN(n25976) );
  NAND2_X1 U34375 ( .A1(n25976), .A2(n29325), .ZN(n25977) );
  INV_X1 U34376 ( .A(n31879), .ZN(n25982) );
  NOR2_X1 U34377 ( .A1(n51479), .A2(n31886), .ZN(n25981) );
  INV_X1 U34378 ( .A(n31883), .ZN(n31803) );
  NOR2_X1 U34379 ( .A1(n30118), .A2(n31803), .ZN(n25980) );
  AOI22_X1 U34380 ( .A1(n25982), .A2(n25981), .B1(n31026), .B2(n25980), .ZN(
        n25985) );
  OAI21_X1 U34381 ( .B1(n51479), .B2(n52047), .A(n31798), .ZN(n25983) );
  NAND3_X1 U34382 ( .A1(n31801), .A2(n31800), .A3(n25983), .ZN(n25984) );
  INV_X1 U34383 ( .A(n42541), .ZN(n25989) );
  XNOR2_X1 U34384 ( .A(n25989), .B(n25988), .ZN(n25990) );
  XNOR2_X1 U34385 ( .A(n33566), .B(n25990), .ZN(n26353) );
  XNOR2_X1 U34386 ( .A(n27372), .B(n25991), .ZN(n26001) );
  INV_X1 U34387 ( .A(n25992), .ZN(n34300) );
  XNOR2_X1 U34388 ( .A(n25993), .B(n2606), .ZN(n43385) );
  XNOR2_X1 U34389 ( .A(n43385), .B(n34614), .ZN(n25994) );
  XNOR2_X1 U34390 ( .A(n34300), .B(n25994), .ZN(n25995) );
  XNOR2_X1 U34391 ( .A(n25996), .B(n25995), .ZN(n25997) );
  XNOR2_X1 U34392 ( .A(n28041), .B(n25997), .ZN(n25998) );
  XNOR2_X1 U34393 ( .A(n25999), .B(n25998), .ZN(n26000) );
  XNOR2_X1 U34394 ( .A(n26002), .B(n4587), .ZN(n34507) );
  XNOR2_X1 U34395 ( .A(n34507), .B(n27204), .ZN(n44557) );
  XNOR2_X1 U34396 ( .A(n45105), .B(n3367), .ZN(n26003) );
  XNOR2_X1 U34397 ( .A(n26003), .B(n41497), .ZN(n26004) );
  XNOR2_X1 U34398 ( .A(n44557), .B(n26004), .ZN(n26005) );
  XNOR2_X1 U34399 ( .A(n27196), .B(n26005), .ZN(n26006) );
  XNOR2_X1 U34400 ( .A(n26006), .B(n28048), .ZN(n26007) );
  XNOR2_X1 U34401 ( .A(n26008), .B(n26007), .ZN(n26012) );
  XNOR2_X1 U34402 ( .A(n26010), .B(n26009), .ZN(n26011) );
  XNOR2_X1 U34403 ( .A(n26011), .B(n26012), .ZN(n26015) );
  XNOR2_X1 U34404 ( .A(n26013), .B(n27217), .ZN(n26014) );
  XNOR2_X1 U34405 ( .A(n26589), .B(n43074), .ZN(n28340) );
  XNOR2_X1 U34406 ( .A(n43076), .B(n40104), .ZN(n26016) );
  XNOR2_X1 U34407 ( .A(n26159), .B(n26016), .ZN(n26017) );
  XNOR2_X1 U34408 ( .A(n28221), .B(n26017), .ZN(n26018) );
  XNOR2_X1 U34409 ( .A(n28341), .B(n27256), .ZN(n26019) );
  XNOR2_X1 U34410 ( .A(n26020), .B(n26019), .ZN(n26024) );
  INV_X1 U34413 ( .A(n35363), .ZN(n26027) );
  XNOR2_X1 U34414 ( .A(n26025), .B(n4926), .ZN(n26026) );
  XNOR2_X1 U34415 ( .A(n26027), .B(n26026), .ZN(n43821) );
  XNOR2_X1 U34416 ( .A(n43821), .B(n45463), .ZN(n26028) );
  XNOR2_X1 U34417 ( .A(n28069), .B(n26028), .ZN(n26029) );
  XNOR2_X1 U34418 ( .A(n26030), .B(n26029), .ZN(n26031) );
  XNOR2_X1 U34419 ( .A(n51750), .B(n26031), .ZN(n26033) );
  XNOR2_X1 U34420 ( .A(n26033), .B(n26032), .ZN(n26038) );
  XNOR2_X1 U34421 ( .A(n26036), .B(n26035), .ZN(n26037) );
  INV_X1 U34422 ( .A(n26207), .ZN(n26040) );
  XNOR2_X1 U34423 ( .A(n26041), .B(n26040), .ZN(n43289) );
  XNOR2_X1 U34424 ( .A(n26042), .B(n4558), .ZN(n44906) );
  XNOR2_X1 U34425 ( .A(n28303), .B(n44906), .ZN(n41598) );
  XNOR2_X1 U34426 ( .A(n43289), .B(n41598), .ZN(n26043) );
  XNOR2_X1 U34427 ( .A(n26044), .B(n26043), .ZN(n26045) );
  XNOR2_X1 U34428 ( .A(n26046), .B(n26045), .ZN(n26048) );
  XNOR2_X1 U34429 ( .A(n26048), .B(n26047), .ZN(n26050) );
  XNOR2_X1 U34431 ( .A(n51121), .B(n26222), .ZN(n26412) );
  XNOR2_X1 U34432 ( .A(n51752), .B(n26125), .ZN(n26054) );
  XNOR2_X1 U34433 ( .A(n26221), .B(n26056), .ZN(n26063) );
  INV_X1 U34434 ( .A(n26057), .ZN(n26058) );
  XNOR2_X1 U34435 ( .A(n26058), .B(n49937), .ZN(n43571) );
  XNOR2_X1 U34436 ( .A(n43571), .B(n43849), .ZN(n26059) );
  XNOR2_X1 U34437 ( .A(n26059), .B(n45406), .ZN(n26060) );
  XNOR2_X1 U34438 ( .A(n26061), .B(n26530), .ZN(n26062) );
  XNOR2_X1 U34439 ( .A(n26063), .B(n26062), .ZN(n26064) );
  NAND2_X1 U34441 ( .A1(n29439), .A2(n29447), .ZN(n26066) );
  AND2_X1 U34442 ( .A1(n27030), .A2(n26067), .ZN(n26073) );
  NOR2_X1 U34443 ( .A1(n26722), .A2(n29438), .ZN(n26070) );
  OAI21_X1 U34444 ( .B1(n26071), .B2(n26070), .A(n26068), .ZN(n26072) );
  NOR2_X1 U34446 ( .A1(n29306), .A2(n29289), .ZN(n29295) );
  INV_X1 U34447 ( .A(n27847), .ZN(n29291) );
  NAND2_X1 U34448 ( .A1(n28699), .A2(n29291), .ZN(n28689) );
  OAI22_X1 U34449 ( .A1(n28684), .A2(n28689), .B1(n29290), .B2(n28688), .ZN(
        n26074) );
  INV_X1 U34450 ( .A(n27844), .ZN(n28686) );
  OAI21_X1 U34452 ( .B1(n29308), .B2(n26083), .A(n51517), .ZN(n26076) );
  NOR2_X1 U34453 ( .A1(n28699), .A2(n27847), .ZN(n26075) );
  AOI22_X1 U34454 ( .A1(n29311), .A2(n28698), .B1(n26076), .B2(n26075), .ZN(
        n26087) );
  NOR2_X1 U34455 ( .A1(n28699), .A2(n29290), .ZN(n26078) );
  NOR2_X1 U34456 ( .A1(n26649), .A2(n26078), .ZN(n26080) );
  NAND2_X1 U34457 ( .A1(n28690), .A2(n28688), .ZN(n26079) );
  INV_X1 U34458 ( .A(n29305), .ZN(n26654) );
  NAND3_X1 U34459 ( .A1(n26654), .A2(n29289), .A3(n29308), .ZN(n26081) );
  OAI21_X1 U34460 ( .B1(n28690), .B2(n26083), .A(n29308), .ZN(n26085) );
  NAND3_X1 U34461 ( .A1(n26085), .A2(n29300), .A3(n26084), .ZN(n26086) );
  BUF_X2 U34462 ( .A(n26203), .Z(n31699) );
  XNOR2_X1 U34463 ( .A(n28106), .B(n42668), .ZN(n26089) );
  XNOR2_X1 U34464 ( .A(n26090), .B(n28423), .ZN(n26091) );
  XNOR2_X1 U34465 ( .A(n26093), .B(n26092), .ZN(n26095) );
  XNOR2_X1 U34466 ( .A(n26095), .B(n26094), .ZN(n26099) );
  INV_X1 U34467 ( .A(n26096), .ZN(n26097) );
  XNOR2_X1 U34468 ( .A(n26097), .B(n27452), .ZN(n26098) );
  XNOR2_X1 U34469 ( .A(n26098), .B(n26099), .ZN(n26110) );
  XNOR2_X1 U34470 ( .A(n26100), .B(n27177), .ZN(n26105) );
  XNOR2_X1 U34471 ( .A(n26101), .B(n4208), .ZN(n42656) );
  XNOR2_X1 U34472 ( .A(n44906), .B(n2183), .ZN(n26102) );
  XNOR2_X1 U34473 ( .A(n42656), .B(n26102), .ZN(n26103) );
  XNOR2_X1 U34474 ( .A(n28103), .B(n26103), .ZN(n26104) );
  XNOR2_X1 U34475 ( .A(n26105), .B(n26104), .ZN(n26108) );
  XNOR2_X1 U34476 ( .A(n26107), .B(n26108), .ZN(n26109) );
  XNOR2_X1 U34477 ( .A(n26110), .B(n26109), .ZN(n26111) );
  XNOR2_X1 U34478 ( .A(n26513), .B(n26111), .ZN(n29568) );
  XNOR2_X1 U34479 ( .A(n34265), .B(n4653), .ZN(n26224) );
  XNOR2_X1 U34480 ( .A(n26224), .B(n4627), .ZN(n32035) );
  XNOR2_X1 U34481 ( .A(n32035), .B(n46552), .ZN(n44233) );
  INV_X1 U34482 ( .A(n43571), .ZN(n26112) );
  XNOR2_X1 U34483 ( .A(n44233), .B(n26112), .ZN(n26113) );
  XNOR2_X1 U34484 ( .A(n26114), .B(n26113), .ZN(n26115) );
  XNOR2_X1 U34485 ( .A(n28396), .B(n26115), .ZN(n26117) );
  XNOR2_X1 U34486 ( .A(n26117), .B(n26116), .ZN(n26118) );
  XNOR2_X1 U34487 ( .A(n26118), .B(n28121), .ZN(n26123) );
  XNOR2_X1 U34488 ( .A(n26121), .B(n26120), .ZN(n26122) );
  XNOR2_X1 U34489 ( .A(n2212), .B(n51752), .ZN(n26127) );
  XNOR2_X1 U34490 ( .A(n26125), .B(n28129), .ZN(n26126) );
  XNOR2_X1 U34491 ( .A(n26129), .B(n26130), .ZN(n26139) );
  XNOR2_X1 U34492 ( .A(n26131), .B(Key[3]), .ZN(n26132) );
  XNOR2_X1 U34493 ( .A(n43746), .B(n26132), .ZN(n26133) );
  XNOR2_X1 U34494 ( .A(n27211), .B(n26134), .ZN(n26135) );
  XNOR2_X1 U34495 ( .A(n26135), .B(n26572), .ZN(n26136) );
  XNOR2_X1 U34496 ( .A(n26137), .B(n26136), .ZN(n26138) );
  XNOR2_X1 U34497 ( .A(n2605), .B(n274), .ZN(n41189) );
  XNOR2_X1 U34498 ( .A(n26378), .B(n41189), .ZN(n26140) );
  XNOR2_X1 U34499 ( .A(n26141), .B(n26140), .ZN(n26142) );
  INV_X1 U34500 ( .A(n42620), .ZN(n26145) );
  XNOR2_X1 U34501 ( .A(n34891), .B(n4597), .ZN(n26143) );
  XNOR2_X1 U34502 ( .A(n26144), .B(n26143), .ZN(n44919) );
  XNOR2_X1 U34503 ( .A(n26145), .B(n44919), .ZN(n26146) );
  XNOR2_X1 U34504 ( .A(n26147), .B(n26146), .ZN(n26149) );
  XNOR2_X1 U34505 ( .A(n26149), .B(n26148), .ZN(n26150) );
  XNOR2_X1 U34506 ( .A(n26150), .B(n28041), .ZN(n26151) );
  XNOR2_X1 U34507 ( .A(n26151), .B(n28280), .ZN(n26157) );
  XNOR2_X1 U34508 ( .A(n26152), .B(n26540), .ZN(n26153) );
  XNOR2_X1 U34509 ( .A(n26153), .B(n593), .ZN(n26154) );
  XNOR2_X1 U34510 ( .A(n26155), .B(n26154), .ZN(n26156) );
  AND2_X1 U34511 ( .A1(n26158), .A2(n27695), .ZN(n29555) );
  XNOR2_X1 U34512 ( .A(n26159), .B(n26160), .ZN(n26168) );
  XNOR2_X1 U34513 ( .A(n26418), .B(n4737), .ZN(n26161) );
  XNOR2_X1 U34514 ( .A(n26161), .B(n33199), .ZN(n26163) );
  XNOR2_X1 U34515 ( .A(n26163), .B(n26162), .ZN(n41886) );
  XNOR2_X1 U34516 ( .A(n26164), .B(n4317), .ZN(n43095) );
  XNOR2_X1 U34517 ( .A(n41886), .B(n43095), .ZN(n26165) );
  XNOR2_X1 U34518 ( .A(n26589), .B(n26165), .ZN(n26166) );
  XNOR2_X1 U34519 ( .A(n28221), .B(n26166), .ZN(n26167) );
  XNOR2_X1 U34520 ( .A(n26167), .B(n26168), .ZN(n26169) );
  XNOR2_X1 U34521 ( .A(n26170), .B(n26169), .ZN(n26172) );
  XNOR2_X1 U34522 ( .A(n26171), .B(n26172), .ZN(n26173) );
  XNOR2_X1 U34523 ( .A(n26175), .B(n26176), .ZN(n28240) );
  XNOR2_X1 U34524 ( .A(n28240), .B(n26177), .ZN(n26186) );
  XNOR2_X1 U34525 ( .A(n26178), .B(n2231), .ZN(n43510) );
  XNOR2_X1 U34526 ( .A(n43510), .B(n42258), .ZN(n26179) );
  XNOR2_X1 U34527 ( .A(n26179), .B(n46144), .ZN(n26181) );
  XNOR2_X1 U34528 ( .A(n26180), .B(n36943), .ZN(n44173) );
  XNOR2_X1 U34529 ( .A(n26181), .B(n44173), .ZN(n26182) );
  XNOR2_X1 U34530 ( .A(n28069), .B(n26182), .ZN(n26184) );
  XNOR2_X1 U34531 ( .A(n26184), .B(n26183), .ZN(n26185) );
  XNOR2_X1 U34532 ( .A(n26186), .B(n26185), .ZN(n26189) );
  XNOR2_X1 U34533 ( .A(n26187), .B(n27477), .ZN(n26188) );
  XNOR2_X1 U34534 ( .A(n26189), .B(n26188), .ZN(n26191) );
  XNOR2_X1 U34535 ( .A(n26191), .B(n26190), .ZN(n26193) );
  OAI21_X1 U34536 ( .B1(n27058), .B2(n743), .A(n27697), .ZN(n26194) );
  OAI21_X1 U34537 ( .B1(n26760), .B2(n27701), .A(n26194), .ZN(n26201) );
  INV_X1 U34538 ( .A(n27058), .ZN(n29564) );
  NOR2_X1 U34539 ( .A1(n6339), .A2(n26197), .ZN(n26195) );
  AOI22_X1 U34540 ( .A1(n29564), .A2(n26195), .B1(n29543), .B2(n29549), .ZN(
        n26200) );
  OAI21_X1 U34541 ( .B1(n26761), .B2(n27701), .A(n27697), .ZN(n26196) );
  AND2_X1 U34542 ( .A1(n29568), .A2(n29559), .ZN(n29557) );
  INV_X1 U34543 ( .A(n29555), .ZN(n26756) );
  AND2_X1 U34545 ( .A1(n29550), .A2(n51111), .ZN(n26750) );
  OAI21_X1 U34546 ( .B1(n26753), .B2(n26750), .A(n27702), .ZN(n26198) );
  NOR2_X1 U34547 ( .A1(n29085), .A2(n32130), .ZN(n26315) );
  INV_X1 U34548 ( .A(n26202), .ZN(n30814) );
  NOR2_X1 U34549 ( .A1(n30814), .A2(n26203), .ZN(n32128) );
  XNOR2_X1 U34550 ( .A(n28103), .B(n28311), .ZN(n26212) );
  INV_X1 U34551 ( .A(n26204), .ZN(n26206) );
  XNOR2_X1 U34552 ( .A(n26206), .B(n26205), .ZN(n41300) );
  XNOR2_X1 U34553 ( .A(n34742), .B(n26207), .ZN(n42859) );
  XNOR2_X1 U34554 ( .A(n42859), .B(n4932), .ZN(n26208) );
  XNOR2_X1 U34555 ( .A(n41300), .B(n26208), .ZN(n26209) );
  XNOR2_X1 U34556 ( .A(n26210), .B(n26209), .ZN(n26211) );
  XNOR2_X1 U34557 ( .A(n26212), .B(n26211), .ZN(n26213) );
  XNOR2_X1 U34558 ( .A(n28439), .B(n370), .ZN(n26215) );
  XNOR2_X1 U34559 ( .A(n26216), .B(n26217), .ZN(n26219) );
  INV_X1 U34560 ( .A(n29533), .ZN(n29513) );
  XNOR2_X1 U34561 ( .A(n26221), .B(n26220), .ZN(n27191) );
  XNOR2_X1 U34562 ( .A(n27191), .B(n26222), .ZN(n26232) );
  INV_X1 U34563 ( .A(n26223), .ZN(n33510) );
  XNOR2_X1 U34564 ( .A(n33510), .B(n4287), .ZN(n43952) );
  XNOR2_X1 U34565 ( .A(n26225), .B(n26224), .ZN(n45270) );
  XNOR2_X1 U34566 ( .A(n43952), .B(n45270), .ZN(n26226) );
  XNOR2_X1 U34567 ( .A(n27501), .B(n26226), .ZN(n26227) );
  XNOR2_X1 U34568 ( .A(n471), .B(n26227), .ZN(n26230) );
  XNOR2_X1 U34569 ( .A(n26230), .B(n26229), .ZN(n26231) );
  XNOR2_X1 U34570 ( .A(n26232), .B(n26231), .ZN(n26233) );
  XNOR2_X1 U34571 ( .A(n26235), .B(n26234), .ZN(n26236) );
  XNOR2_X1 U34572 ( .A(n26236), .B(n26237), .ZN(n26241) );
  XNOR2_X1 U34573 ( .A(n26239), .B(n26238), .ZN(n26240) );
  XNOR2_X1 U34574 ( .A(n26241), .B(n26240), .ZN(n26253) );
  XNOR2_X1 U34575 ( .A(n26243), .B(n26242), .ZN(n44385) );
  XNOR2_X1 U34576 ( .A(n26244), .B(n4845), .ZN(n46084) );
  XNOR2_X1 U34577 ( .A(n46084), .B(n4613), .ZN(n26245) );
  XNOR2_X1 U34578 ( .A(n44385), .B(n26245), .ZN(n26246) );
  XNOR2_X1 U34579 ( .A(n2080), .B(n26246), .ZN(n26247) );
  XNOR2_X1 U34580 ( .A(n26247), .B(n26581), .ZN(n26249) );
  XNOR2_X1 U34581 ( .A(n26248), .B(n26249), .ZN(n26251) );
  XNOR2_X1 U34582 ( .A(n26250), .B(n26251), .ZN(n26252) );
  INV_X1 U34583 ( .A(n26254), .ZN(n26255) );
  XNOR2_X1 U34584 ( .A(n26255), .B(n26256), .ZN(n26271) );
  XNOR2_X1 U34585 ( .A(n28232), .B(n26257), .ZN(n26258) );
  XNOR2_X1 U34586 ( .A(n26259), .B(n26258), .ZN(n45347) );
  XNOR2_X1 U34587 ( .A(n4667), .B(n4712), .ZN(n26260) );
  XNOR2_X1 U34588 ( .A(n26260), .B(n45736), .ZN(n43938) );
  XNOR2_X1 U34589 ( .A(n4926), .B(n4855), .ZN(n26261) );
  XNOR2_X1 U34590 ( .A(n43938), .B(n26261), .ZN(n26262) );
  XNOR2_X1 U34591 ( .A(n45347), .B(n26262), .ZN(n26263) );
  XNOR2_X1 U34592 ( .A(n26264), .B(n26263), .ZN(n26266) );
  XNOR2_X1 U34593 ( .A(n26266), .B(n26265), .ZN(n26267) );
  XNOR2_X1 U34594 ( .A(n26268), .B(n26267), .ZN(n26269) );
  XNOR2_X1 U34595 ( .A(n26269), .B(n27330), .ZN(n26270) );
  INV_X1 U34596 ( .A(n26288), .ZN(n26310) );
  AND2_X1 U34597 ( .A1(n28623), .A2(n26310), .ZN(n29518) );
  XNOR2_X1 U34598 ( .A(n27203), .B(n4638), .ZN(n45104) );
  XNOR2_X1 U34599 ( .A(n35376), .B(n45104), .ZN(n42369) );
  XNOR2_X1 U34600 ( .A(n51424), .B(n42369), .ZN(n26275) );
  XNOR2_X1 U34601 ( .A(n26276), .B(n26275), .ZN(n26278) );
  XNOR2_X1 U34602 ( .A(n28370), .B(n4554), .ZN(n27199) );
  XNOR2_X1 U34603 ( .A(n26279), .B(n27199), .ZN(n26282) );
  INV_X1 U34604 ( .A(n26280), .ZN(n26281) );
  XNOR2_X1 U34605 ( .A(n26282), .B(n26281), .ZN(n26283) );
  INV_X1 U34606 ( .A(Key[57]), .ZN(n48614) );
  XNOR2_X1 U34607 ( .A(n28257), .B(n48614), .ZN(n26284) );
  XNOR2_X1 U34608 ( .A(n26285), .B(n26284), .ZN(n26286) );
  XNOR2_X1 U34609 ( .A(n26287), .B(n26286), .ZN(n27430) );
  NAND2_X1 U34610 ( .A1(n29526), .A2(n28626), .ZN(n29534) );
  NAND2_X1 U34611 ( .A1(n29534), .A2(n29513), .ZN(n27800) );
  XNOR2_X1 U34612 ( .A(n26289), .B(n49414), .ZN(n41188) );
  XNOR2_X1 U34613 ( .A(n41188), .B(n4880), .ZN(n26290) );
  XNOR2_X1 U34614 ( .A(n27232), .B(n26290), .ZN(n26291) );
  XNOR2_X1 U34615 ( .A(n26292), .B(n26291), .ZN(n26293) );
  XNOR2_X1 U34616 ( .A(n26294), .B(n26293), .ZN(n28046) );
  XNOR2_X1 U34617 ( .A(n26296), .B(n26295), .ZN(n27484) );
  XNOR2_X1 U34618 ( .A(n27484), .B(n26297), .ZN(n42835) );
  XNOR2_X1 U34619 ( .A(n41223), .B(n4325), .ZN(n26298) );
  XNOR2_X1 U34620 ( .A(n42835), .B(n26298), .ZN(n26299) );
  XNOR2_X1 U34621 ( .A(n26300), .B(n26299), .ZN(n26301) );
  XNOR2_X1 U34622 ( .A(n26302), .B(n26301), .ZN(n26303) );
  XNOR2_X1 U34623 ( .A(n26304), .B(n27224), .ZN(n26305) );
  XNOR2_X1 U34624 ( .A(n26556), .B(n26305), .ZN(n27495) );
  AND2_X1 U34625 ( .A1(n28622), .A2(n51747), .ZN(n26980) );
  NAND2_X1 U34626 ( .A1(n26980), .A2(n28614), .ZN(n26983) );
  INV_X1 U34627 ( .A(n26306), .ZN(n29532) );
  INV_X1 U34628 ( .A(n28622), .ZN(n26973) );
  NAND3_X1 U34629 ( .A1(n29521), .A2(n28615), .A3(n29528), .ZN(n26307) );
  AND2_X1 U34630 ( .A1(n26983), .A2(n26307), .ZN(n26346) );
  OAI21_X1 U34631 ( .B1(n28618), .B2(n29512), .A(n29513), .ZN(n26309) );
  AND2_X1 U34632 ( .A1(n26310), .A2(n29535), .ZN(n28629) );
  OAI21_X1 U34633 ( .B1(n28629), .B2(n28623), .A(n398), .ZN(n26308) );
  NAND2_X1 U34634 ( .A1(n29505), .A2(n26310), .ZN(n26342) );
  INV_X1 U34635 ( .A(n29522), .ZN(n27797) );
  INV_X1 U34637 ( .A(n27795), .ZN(n26312) );
  NAND2_X1 U34638 ( .A1(n26700), .A2(n26312), .ZN(n26345) );
  AND2_X1 U34639 ( .A1(n28618), .A2(n29526), .ZN(n26340) );
  NAND2_X1 U34640 ( .A1(n26340), .A2(n29522), .ZN(n26313) );
  OAI211_X1 U34641 ( .C1(n26342), .C2(n27797), .A(n26345), .B(n26313), .ZN(
        n26314) );
  MUX2_X1 U34642 ( .A(n29320), .B(n29315), .S(n29330), .Z(n26318) );
  AOI21_X1 U34643 ( .B1(n51107), .B2(n52217), .A(n28641), .ZN(n26316) );
  NOR2_X1 U34644 ( .A1(n26316), .A2(n52177), .ZN(n26317) );
  NAND2_X1 U34645 ( .A1(n26318), .A2(n26317), .ZN(n26327) );
  NAND2_X1 U34646 ( .A1(n27896), .A2(n29320), .ZN(n26319) );
  INV_X1 U34647 ( .A(n29329), .ZN(n29321) );
  INV_X1 U34648 ( .A(n29331), .ZN(n29323) );
  NAND2_X1 U34649 ( .A1(n51107), .A2(n29319), .ZN(n26320) );
  AND2_X1 U34650 ( .A1(n29315), .A2(n26320), .ZN(n26321) );
  AOI22_X1 U34651 ( .A1(n26321), .A2(n27818), .B1(n27897), .B2(n28644), .ZN(
        n26326) );
  INV_X1 U34652 ( .A(n26323), .ZN(n27820) );
  OR2_X1 U34653 ( .A1(n26328), .A2(n31712), .ZN(n26352) );
  NAND4_X1 U34654 ( .A1(n28671), .A2(n26668), .A3(n26677), .A4(n26676), .ZN(
        n26333) );
  NAND3_X1 U34655 ( .A1(n2294), .A2(n26668), .A3(n25841), .ZN(n26332) );
  NAND4_X1 U34656 ( .A1(n29479), .A2(n26668), .A3(n26671), .A4(n28669), .ZN(
        n26331) );
  AND3_X1 U34657 ( .A1(n26333), .A2(n26332), .A3(n26331), .ZN(n26339) );
  AOI21_X1 U34658 ( .B1(n28674), .B2(n26334), .A(n29480), .ZN(n26337) );
  NAND2_X1 U34659 ( .A1(n28669), .A2(n28666), .ZN(n29486) );
  NAND2_X1 U34660 ( .A1(n27858), .A2(n28669), .ZN(n26335) );
  OAI21_X1 U34661 ( .B1(n29486), .B2(n25841), .A(n26335), .ZN(n26336) );
  NOR2_X1 U34662 ( .A1(n26337), .A2(n26336), .ZN(n26338) );
  MUX2_X1 U34663 ( .A(n31709), .B(n29976), .S(n31699), .Z(n26347) );
  INV_X1 U34664 ( .A(n26340), .ZN(n26341) );
  NAND2_X1 U34665 ( .A1(n26342), .A2(n26341), .ZN(n26343) );
  OAI21_X1 U34666 ( .B1(n721), .B2(n31711), .A(n26348), .ZN(n32138) );
  NAND2_X1 U34667 ( .A1(n32120), .A2(n31711), .ZN(n29973) );
  INV_X1 U34668 ( .A(n26348), .ZN(n31701) );
  NAND2_X1 U34669 ( .A1(n721), .A2(n32130), .ZN(n31706) );
  OAI21_X1 U34670 ( .B1(n31699), .B2(n31712), .A(n30814), .ZN(n26349) );
  OR2_X1 U34671 ( .A1(n26203), .A2(n32130), .ZN(n30811) );
  XNOR2_X1 U34672 ( .A(n26353), .B(n35501), .ZN(n26718) );
  XNOR2_X1 U34673 ( .A(n26355), .B(n26354), .ZN(n26367) );
  INV_X1 U34674 ( .A(n26356), .ZN(n35292) );
  XNOR2_X1 U34675 ( .A(n26358), .B(n26357), .ZN(n43649) );
  XNOR2_X1 U34676 ( .A(n43649), .B(n26359), .ZN(n26360) );
  XNOR2_X1 U34677 ( .A(n28249), .B(n26361), .ZN(n26363) );
  XNOR2_X1 U34678 ( .A(n26363), .B(n26362), .ZN(n26365) );
  XNOR2_X1 U34679 ( .A(n26365), .B(n26364), .ZN(n26366) );
  XNOR2_X1 U34680 ( .A(n26368), .B(n28267), .ZN(n42385) );
  XOR2_X1 U34681 ( .A(n2947), .B(n4542), .Z(n26369) );
  XNOR2_X1 U34682 ( .A(n26370), .B(n26369), .ZN(n45123) );
  XNOR2_X1 U34683 ( .A(n42385), .B(n45123), .ZN(n26371) );
  XNOR2_X1 U34684 ( .A(n28274), .B(n26371), .ZN(n26372) );
  XNOR2_X1 U34685 ( .A(n26374), .B(n26373), .ZN(n26382) );
  XNOR2_X1 U34686 ( .A(n26375), .B(n4755), .ZN(n26376) );
  XNOR2_X1 U34687 ( .A(n26376), .B(n26544), .ZN(n28036) );
  XNOR2_X1 U34688 ( .A(n27226), .B(n28036), .ZN(n26381) );
  XNOR2_X1 U34689 ( .A(n26378), .B(n26377), .ZN(n26379) );
  XNOR2_X1 U34690 ( .A(n27222), .B(n26379), .ZN(n26380) );
  INV_X1 U34691 ( .A(n28915), .ZN(n28931) );
  XNOR2_X1 U34692 ( .A(n26386), .B(n26385), .ZN(n45040) );
  XNOR2_X1 U34693 ( .A(n26387), .B(n4589), .ZN(n42344) );
  XNOR2_X1 U34694 ( .A(n42344), .B(n42349), .ZN(n26388) );
  XNOR2_X1 U34695 ( .A(n45040), .B(n26388), .ZN(n26389) );
  XNOR2_X1 U34696 ( .A(n26390), .B(n26389), .ZN(n26391) );
  XNOR2_X1 U34697 ( .A(n26391), .B(n28431), .ZN(n26392) );
  XNOR2_X1 U34698 ( .A(n26393), .B(n26392), .ZN(n26394) );
  XNOR2_X1 U34699 ( .A(n2209), .B(n28430), .ZN(n28100) );
  XNOR2_X1 U34700 ( .A(n26394), .B(n28100), .ZN(n26399) );
  XNOR2_X1 U34701 ( .A(n27451), .B(n28423), .ZN(n26396) );
  XNOR2_X1 U34702 ( .A(n26396), .B(n26395), .ZN(n27172) );
  XNOR2_X1 U34703 ( .A(n27172), .B(n26397), .ZN(n26398) );
  XNOR2_X1 U34704 ( .A(n26399), .B(n26398), .ZN(n26400) );
  XNOR2_X1 U34705 ( .A(n28400), .B(n26401), .ZN(n26411) );
  XNOR2_X1 U34706 ( .A(n26403), .B(n4612), .ZN(n44311) );
  XNOR2_X1 U34707 ( .A(n46122), .B(n26404), .ZN(n26405) );
  XNOR2_X1 U34708 ( .A(n44311), .B(n26405), .ZN(n26406) );
  XNOR2_X1 U34709 ( .A(n26406), .B(n46126), .ZN(n26407) );
  XNOR2_X1 U34710 ( .A(n28291), .B(n26407), .ZN(n26408) );
  XNOR2_X1 U34711 ( .A(n26409), .B(n26408), .ZN(n26410) );
  XNOR2_X1 U34712 ( .A(n26411), .B(n26410), .ZN(n26413) );
  INV_X1 U34714 ( .A(n28566), .ZN(n26416) );
  INV_X1 U34715 ( .A(n26417), .ZN(n26428) );
  XNOR2_X1 U34716 ( .A(n26418), .B(n4502), .ZN(n26422) );
  INV_X1 U34717 ( .A(n26419), .ZN(n26421) );
  XNOR2_X1 U34718 ( .A(n33474), .B(n4026), .ZN(n26420) );
  XNOR2_X1 U34719 ( .A(n26421), .B(n26420), .ZN(n41948) );
  XNOR2_X1 U34720 ( .A(n26422), .B(n41948), .ZN(n26423) );
  XNOR2_X1 U34721 ( .A(n26589), .B(n26423), .ZN(n26424) );
  XNOR2_X1 U34722 ( .A(n28213), .B(n26424), .ZN(n26426) );
  XNOR2_X1 U34723 ( .A(n26425), .B(n26426), .ZN(n26427) );
  XNOR2_X1 U34724 ( .A(n26428), .B(n26427), .ZN(n26430) );
  XNOR2_X1 U34725 ( .A(n26430), .B(n26429), .ZN(n26438) );
  XNOR2_X1 U34726 ( .A(n2080), .B(n23525), .ZN(n26433) );
  XNOR2_X1 U34727 ( .A(n26432), .B(n26433), .ZN(n26434) );
  XNOR2_X1 U34728 ( .A(n27439), .B(n26434), .ZN(n28098) );
  XNOR2_X1 U34729 ( .A(n26435), .B(n5016), .ZN(n28343) );
  XNOR2_X1 U34730 ( .A(n28098), .B(n26596), .ZN(n26437) );
  XNOR2_X1 U34731 ( .A(n26438), .B(n26437), .ZN(n26458) );
  INV_X1 U34732 ( .A(n26439), .ZN(n26440) );
  XNOR2_X1 U34733 ( .A(n26440), .B(n27325), .ZN(n26441) );
  XNOR2_X1 U34734 ( .A(n26442), .B(n26441), .ZN(n26454) );
  INV_X1 U34735 ( .A(n26443), .ZN(n26444) );
  XNOR2_X1 U34736 ( .A(n26444), .B(n4908), .ZN(n44366) );
  XNOR2_X1 U34737 ( .A(n46146), .B(n26445), .ZN(n26446) );
  XNOR2_X1 U34738 ( .A(n44366), .B(n26446), .ZN(n26447) );
  XNOR2_X1 U34739 ( .A(n26448), .B(n26447), .ZN(n26449) );
  XNOR2_X1 U34740 ( .A(n26611), .B(n26449), .ZN(n26451) );
  XNOR2_X1 U34741 ( .A(n26451), .B(n26450), .ZN(n26453) );
  AND2_X1 U34742 ( .A1(n29013), .A2(n3160), .ZN(n28201) );
  OAI211_X1 U34743 ( .C1(n28931), .C2(n51115), .A(n28571), .B(n28201), .ZN(
        n26457) );
  OR2_X1 U34744 ( .A1(n28922), .A2(n28194), .ZN(n26456) );
  NAND2_X1 U34745 ( .A1(n28919), .A2(n28923), .ZN(n28196) );
  INV_X1 U34746 ( .A(n28196), .ZN(n28203) );
  INV_X1 U34747 ( .A(n28916), .ZN(n28933) );
  NAND2_X1 U34748 ( .A1(n28933), .A2(n28926), .ZN(n28197) );
  NAND4_X1 U34749 ( .A1(n28203), .A2(n29007), .A3(n28197), .A4(n28194), .ZN(
        n28207) );
  NAND4_X1 U34750 ( .A1(n26457), .A2(n26456), .A3(n28207), .A4(n28014), .ZN(
        n26465) );
  AOI22_X1 U34751 ( .A1(n28007), .A2(n29011), .B1(n28566), .B2(n28918), .ZN(
        n26461) );
  NAND2_X1 U34752 ( .A1(n26459), .A2(n29013), .ZN(n26460) );
  NAND2_X1 U34753 ( .A1(n26461), .A2(n26460), .ZN(n26463) );
  NAND3_X1 U34754 ( .A1(n29018), .A2(n29011), .A3(n28933), .ZN(n26462) );
  AOI21_X1 U34755 ( .B1(n26463), .B2(n26462), .A(n51115), .ZN(n26464) );
  AOI22_X1 U34756 ( .A1(n30303), .A2(n739), .B1(n26466), .B2(n25199), .ZN(
        n26471) );
  OAI211_X1 U34757 ( .C1(n28025), .C2(n30163), .A(n28032), .B(n30172), .ZN(
        n26469) );
  OR2_X1 U34758 ( .A1(n27987), .A2(n28588), .ZN(n26473) );
  OAI21_X1 U34759 ( .B1(n28582), .B2(n27991), .A(n26473), .ZN(n26474) );
  AOI21_X1 U34760 ( .B1(n26475), .B2(n51118), .A(n27998), .ZN(n26481) );
  AND2_X1 U34761 ( .A1(n28587), .A2(n28578), .ZN(n27990) );
  OAI21_X1 U34762 ( .B1(n26477), .B2(n27990), .A(n26476), .ZN(n26480) );
  OR2_X1 U34763 ( .A1(n27987), .A2(n28587), .ZN(n27994) );
  NOR2_X1 U34764 ( .A1(n27994), .A2(n26478), .ZN(n28893) );
  NAND3_X1 U34765 ( .A1(n28893), .A2(n51118), .A3(n28894), .ZN(n26479) );
  OR2_X1 U34767 ( .A1(n27145), .A2(n27957), .ZN(n29169) );
  NOR2_X1 U34768 ( .A1(n29172), .A2(n26483), .ZN(n26484) );
  OAI21_X1 U34770 ( .B1(n30251), .B2(n29158), .A(n26486), .ZN(n26487) );
  INV_X1 U34771 ( .A(n26487), .ZN(n26491) );
  NAND2_X1 U34772 ( .A1(n26489), .A2(n29153), .ZN(n26490) );
  NOR2_X1 U34773 ( .A1(n31384), .A2(n30534), .ZN(n33006) );
  NAND2_X1 U34774 ( .A1(n30543), .A2(n33006), .ZN(n26634) );
  MUX2_X1 U34775 ( .A(n26501), .B(n30279), .S(n28148), .Z(n26493) );
  NOR2_X1 U34776 ( .A1(n26493), .A2(n30290), .ZN(n26497) );
  NAND2_X1 U34777 ( .A1(n27111), .A2(n26494), .ZN(n30281) );
  NAND2_X1 U34778 ( .A1(n27111), .A2(n30285), .ZN(n26495) );
  AOI21_X1 U34779 ( .B1(n30281), .B2(n30280), .A(n26495), .ZN(n26496) );
  MUX2_X1 U34780 ( .A(n26497), .B(n26496), .S(n30282), .Z(n26505) );
  NAND3_X1 U34781 ( .A1(n28147), .A2(n28560), .A3(n2881), .ZN(n26499) );
  NAND2_X1 U34782 ( .A1(n30291), .A2(n30285), .ZN(n26498) );
  NAND2_X1 U34783 ( .A1(n26500), .A2(n30295), .ZN(n28152) );
  NAND2_X1 U34784 ( .A1(n51748), .A2(n30295), .ZN(n28143) );
  INV_X1 U34785 ( .A(n28560), .ZN(n26502) );
  NOR2_X1 U34786 ( .A1(n30279), .A2(n27113), .ZN(n28546) );
  XNOR2_X1 U34787 ( .A(n26506), .B(n4886), .ZN(n44506) );
  XNOR2_X1 U34788 ( .A(n42215), .B(n44506), .ZN(n26507) );
  XNOR2_X1 U34789 ( .A(n26508), .B(n26507), .ZN(n26510) );
  XNOR2_X1 U34790 ( .A(n26510), .B(n26509), .ZN(n26511) );
  XNOR2_X1 U34791 ( .A(n26511), .B(n27446), .ZN(n26512) );
  XNOR2_X1 U34792 ( .A(n28101), .B(n26512), .ZN(n26515) );
  INV_X1 U34793 ( .A(n26513), .ZN(n26514) );
  XNOR2_X1 U34794 ( .A(n26515), .B(n26514), .ZN(n26517) );
  XNOR2_X1 U34795 ( .A(n51752), .B(n26518), .ZN(n26522) );
  INV_X1 U34796 ( .A(n26520), .ZN(n26521) );
  XNOR2_X1 U34797 ( .A(n26522), .B(n26521), .ZN(n26524) );
  XNOR2_X1 U34798 ( .A(n26524), .B(n26523), .ZN(n26539) );
  XNOR2_X1 U34799 ( .A(n41314), .B(n4874), .ZN(n36293) );
  XNOR2_X1 U34800 ( .A(n26526), .B(n26525), .ZN(n43030) );
  XNOR2_X1 U34801 ( .A(n43030), .B(n4636), .ZN(n26527) );
  XNOR2_X1 U34802 ( .A(n36293), .B(n26527), .ZN(n26528) );
  XNOR2_X1 U34803 ( .A(n26529), .B(n26528), .ZN(n26533) );
  XNOR2_X1 U34804 ( .A(n26531), .B(n26530), .ZN(n26532) );
  XNOR2_X1 U34805 ( .A(n26533), .B(n26532), .ZN(n26534) );
  XNOR2_X1 U34806 ( .A(n26534), .B(n28119), .ZN(n26537) );
  XNOR2_X1 U34807 ( .A(n26536), .B(n26535), .ZN(n28401) );
  XNOR2_X1 U34808 ( .A(n26537), .B(n28401), .ZN(n26538) );
  XNOR2_X1 U34809 ( .A(n26540), .B(n51647), .ZN(n26546) );
  INV_X1 U34810 ( .A(n44539), .ZN(n26542) );
  XNOR2_X1 U34811 ( .A(n34891), .B(n26541), .ZN(n42274) );
  XNOR2_X1 U34812 ( .A(n26542), .B(n42274), .ZN(n26543) );
  XNOR2_X1 U34813 ( .A(n26544), .B(n26543), .ZN(n26545) );
  XNOR2_X1 U34814 ( .A(n26546), .B(n26545), .ZN(n26550) );
  XNOR2_X1 U34815 ( .A(n26548), .B(n26547), .ZN(n26549) );
  XNOR2_X1 U34816 ( .A(n26550), .B(n26549), .ZN(n26554) );
  XNOR2_X1 U34817 ( .A(n27373), .B(n2082), .ZN(n26551) );
  XNOR2_X1 U34818 ( .A(n26553), .B(n52163), .ZN(n28407) );
  XNOR2_X1 U34819 ( .A(n26554), .B(n28407), .ZN(n26560) );
  XNOR2_X1 U34820 ( .A(n51057), .B(n26556), .ZN(n26557) );
  XNOR2_X1 U34821 ( .A(n26558), .B(n26557), .ZN(n26559) );
  XNOR2_X1 U34822 ( .A(n26560), .B(n26559), .ZN(n28870) );
  XNOR2_X1 U34823 ( .A(n36739), .B(n41835), .ZN(n33732) );
  XNOR2_X1 U34824 ( .A(n41156), .B(n26561), .ZN(n26562) );
  XNOR2_X1 U34825 ( .A(n33732), .B(n26562), .ZN(n26563) );
  XNOR2_X1 U34826 ( .A(n33297), .B(n33635), .ZN(n43745) );
  XNOR2_X1 U34827 ( .A(n26563), .B(n43745), .ZN(n26564) );
  XNOR2_X1 U34828 ( .A(n51751), .B(n26564), .ZN(n26566) );
  XNOR2_X1 U34829 ( .A(n26565), .B(n26566), .ZN(n26568) );
  XNOR2_X1 U34830 ( .A(n26568), .B(n51120), .ZN(n26570) );
  XNOR2_X1 U34831 ( .A(n26569), .B(n26570), .ZN(n26580) );
  XNOR2_X1 U34832 ( .A(n26572), .B(n26571), .ZN(n26577) );
  XNOR2_X1 U34833 ( .A(n26573), .B(n51423), .ZN(n26574) );
  XNOR2_X1 U34834 ( .A(n26575), .B(n26574), .ZN(n26576) );
  NAND2_X1 U34837 ( .A1(n27104), .A2(n29032), .ZN(n26616) );
  AND2_X1 U34838 ( .A1(n26619), .A2(n28882), .ZN(n28871) );
  INV_X1 U34839 ( .A(n28870), .ZN(n29028) );
  NAND2_X1 U34840 ( .A1(n28871), .A2(n28875), .ZN(n26615) );
  INV_X1 U34841 ( .A(n27290), .ZN(n26583) );
  XNOR2_X1 U34842 ( .A(n25508), .B(n23525), .ZN(n26582) );
  XNOR2_X1 U34843 ( .A(n26582), .B(n26583), .ZN(n26585) );
  XNOR2_X1 U34844 ( .A(n27242), .B(n26584), .ZN(n28226) );
  XNOR2_X1 U34845 ( .A(n26585), .B(n28226), .ZN(n26595) );
  XNOR2_X1 U34846 ( .A(n32497), .B(n33746), .ZN(n42975) );
  XNOR2_X1 U34847 ( .A(n26586), .B(n4835), .ZN(n40995) );
  XNOR2_X1 U34848 ( .A(n33199), .B(n40995), .ZN(n26587) );
  XNOR2_X1 U34849 ( .A(n42975), .B(n26587), .ZN(n26588) );
  XNOR2_X1 U34850 ( .A(n26589), .B(n26588), .ZN(n26590) );
  XNOR2_X1 U34851 ( .A(n26591), .B(n26590), .ZN(n26593) );
  XNOR2_X1 U34852 ( .A(n26593), .B(n26592), .ZN(n26594) );
  XNOR2_X1 U34853 ( .A(n26595), .B(n26594), .ZN(n26598) );
  XNOR2_X1 U34854 ( .A(n28218), .B(n26596), .ZN(n26597) );
  XNOR2_X2 U34855 ( .A(n26598), .B(n26597), .ZN(n28874) );
  XNOR2_X1 U34856 ( .A(n26599), .B(n28080), .ZN(n26609) );
  XNOR2_X1 U34857 ( .A(n36943), .B(n26601), .ZN(n26602) );
  XNOR2_X1 U34858 ( .A(n28234), .B(n26602), .ZN(n43041) );
  XNOR2_X1 U34859 ( .A(n36941), .B(n26603), .ZN(n26605) );
  XNOR2_X1 U34860 ( .A(n26605), .B(n26604), .ZN(n39537) );
  XNOR2_X1 U34861 ( .A(n43041), .B(n39537), .ZN(n26606) );
  XNOR2_X1 U34862 ( .A(n51750), .B(n26606), .ZN(n26608) );
  XNOR2_X1 U34863 ( .A(n26611), .B(n26610), .ZN(n28356) );
  XNOR2_X1 U34864 ( .A(n28356), .B(n26612), .ZN(n26613) );
  XNOR2_X1 U34865 ( .A(n28242), .B(n26613), .ZN(n26614) );
  INV_X1 U34866 ( .A(n29027), .ZN(n29034) );
  MUX2_X1 U34867 ( .A(n26616), .B(n26615), .S(n29034), .Z(n26625) );
  OAI21_X1 U34868 ( .B1(n29032), .B2(n29035), .A(n29030), .ZN(n26617) );
  NAND2_X1 U34869 ( .A1(n29045), .A2(n26617), .ZN(n26618) );
  AND2_X1 U34870 ( .A1(n27102), .A2(n26618), .ZN(n26624) );
  NAND2_X1 U34871 ( .A1(n29033), .A2(n29035), .ZN(n26620) );
  NOR2_X1 U34872 ( .A1(n28536), .A2(n26620), .ZN(n29047) );
  NAND2_X1 U34873 ( .A1(n29047), .A2(n29029), .ZN(n26623) );
  AOI21_X1 U34874 ( .B1(n28874), .B2(n28870), .A(n28155), .ZN(n26621) );
  NAND4_X1 U34875 ( .A1(n26625), .A2(n26624), .A3(n26623), .A4(n26622), .ZN(
        n26633) );
  OAI22_X1 U34876 ( .A1(n26626), .A2(n27103), .B1(n28877), .B2(n29028), .ZN(
        n26627) );
  NOR2_X1 U34877 ( .A1(n29027), .A2(n28160), .ZN(n28528) );
  AND2_X1 U34878 ( .A1(n29030), .A2(n28155), .ZN(n28880) );
  OAI21_X1 U34879 ( .B1(n26627), .B2(n28528), .A(n28880), .ZN(n26631) );
  OAI22_X1 U34880 ( .A1(n28882), .A2(n27103), .B1(n29027), .B2(n29038), .ZN(
        n26629) );
  NOR2_X1 U34881 ( .A1(n28877), .A2(n28875), .ZN(n26628) );
  OAI211_X1 U34882 ( .C1(n26629), .C2(n26628), .A(n29030), .B(n29035), .ZN(
        n26630) );
  NAND2_X1 U34883 ( .A1(n30528), .A2(n33005), .ZN(n30533) );
  NOR2_X1 U34884 ( .A1(n33005), .A2(n30534), .ZN(n31375) );
  AND2_X1 U34885 ( .A1(n31383), .A2(n30534), .ZN(n33007) );
  NAND2_X1 U34886 ( .A1(n33007), .A2(n51740), .ZN(n30529) );
  NOR2_X1 U34887 ( .A1(n33005), .A2(n51740), .ZN(n31011) );
  XNOR2_X1 U34889 ( .A(n720), .B(n31383), .ZN(n26636) );
  NAND4_X1 U34890 ( .A1(n33017), .A2(n33013), .A3(n31380), .A4(n26636), .ZN(
        n26637) );
  OAI211_X1 U34892 ( .C1(n26640), .C2(n6602), .A(n27024), .B(n27836), .ZN(
        n26641) );
  AND2_X1 U34893 ( .A1(n29439), .A2(n27040), .ZN(n26645) );
  INV_X1 U34894 ( .A(n26645), .ZN(n26642) );
  NAND2_X1 U34895 ( .A1(n26644), .A2(n26643), .ZN(n26648) );
  OR2_X1 U34896 ( .A1(n27840), .A2(n29446), .ZN(n26727) );
  NAND2_X1 U34897 ( .A1(n26645), .A2(n26723), .ZN(n26646) );
  INV_X1 U34898 ( .A(n26650), .ZN(n26652) );
  NAND3_X1 U34899 ( .A1(n26652), .A2(n26651), .A3(n51518), .ZN(n26656) );
  INV_X1 U34900 ( .A(n28688), .ZN(n26653) );
  NAND3_X1 U34901 ( .A1(n26654), .A2(n26653), .A3(n29308), .ZN(n26655) );
  NAND2_X1 U34902 ( .A1(n28695), .A2(n29294), .ZN(n29296) );
  NOR2_X1 U34903 ( .A1(n29296), .A2(n51518), .ZN(n28692) );
  NAND2_X1 U34904 ( .A1(n29308), .A2(n27844), .ZN(n26658) );
  OAI21_X1 U34905 ( .B1(n27844), .B2(n28690), .A(n29289), .ZN(n26657) );
  OAI21_X1 U34906 ( .B1(n28692), .B2(n26658), .A(n26657), .ZN(n26664) );
  INV_X1 U34907 ( .A(n26659), .ZN(n26660) );
  NAND2_X1 U34908 ( .A1(n29311), .A2(n26660), .ZN(n26663) );
  INV_X1 U34909 ( .A(n28689), .ZN(n26661) );
  OAI21_X1 U34910 ( .B1(n29295), .B2(n26661), .A(n29303), .ZN(n26662) );
  OAI211_X1 U34911 ( .C1(n29494), .C2(n26667), .A(n26666), .B(n29498), .ZN(
        n26673) );
  OAI21_X1 U34913 ( .B1(n29478), .B2(n27860), .A(n26668), .ZN(n26669) );
  OAI21_X1 U34915 ( .B1(n28674), .B2(n29480), .A(n26670), .ZN(n26672) );
  NAND3_X1 U34916 ( .A1(n25841), .A2(n51110), .A3(n28666), .ZN(n26674) );
  NAND2_X1 U34917 ( .A1(n2956), .A2(n26674), .ZN(n26675) );
  OAI21_X1 U34918 ( .B1(n26677), .B2(n26679), .A(n27863), .ZN(n26678) );
  NAND2_X1 U34919 ( .A1(n26678), .A2(n28671), .ZN(n26680) );
  INV_X1 U34920 ( .A(n26679), .ZN(n29493) );
  NAND3_X1 U34921 ( .A1(n2294), .A2(n29493), .A3(n29479), .ZN(n29500) );
  NOR2_X1 U34922 ( .A1(n26761), .A2(n29549), .ZN(n27051) );
  INV_X1 U34923 ( .A(n29546), .ZN(n29551) );
  AOI22_X1 U34924 ( .A1(n27051), .A2(n29551), .B1(n27702), .B2(n27049), .ZN(
        n26687) );
  NAND2_X1 U34925 ( .A1(n8454), .A2(n27049), .ZN(n26683) );
  OAI211_X1 U34926 ( .C1(n27058), .C2(n29559), .A(n29554), .B(n26683), .ZN(
        n26684) );
  NAND2_X1 U34927 ( .A1(n26684), .A2(n29549), .ZN(n26685) );
  NAND3_X1 U34929 ( .A1(n30580), .A2(n31033), .A3(n31815), .ZN(n26688) );
  OAI22_X1 U34930 ( .A1(n26787), .A2(n29461), .B1(n27012), .B2(n27762), .ZN(
        n26689) );
  NOR2_X1 U34931 ( .A1(n26690), .A2(n26689), .ZN(n26697) );
  INV_X1 U34932 ( .A(n29456), .ZN(n26691) );
  NAND2_X1 U34933 ( .A1(n29462), .A2(n26781), .ZN(n26693) );
  AND2_X1 U34934 ( .A1(n27765), .A2(n29467), .ZN(n27744) );
  NAND4_X1 U34935 ( .A1(n29471), .A2(n29462), .A3(n27764), .A4(n27744), .ZN(
        n26692) );
  OAI21_X1 U34936 ( .B1(n29460), .B2(n26693), .A(n26692), .ZN(n26694) );
  AOI21_X1 U34937 ( .B1(n27742), .B2(n27755), .A(n26694), .ZN(n26696) );
  NOR2_X1 U34938 ( .A1(n29460), .A2(n7973), .ZN(n27749) );
  AND2_X1 U34939 ( .A1(n27764), .A2(n29463), .ZN(n29468) );
  OAI211_X1 U34940 ( .C1(n27749), .C2(n732), .A(n29468), .B(n27015), .ZN(
        n26695) );
  NAND2_X1 U34941 ( .A1(n6059), .A2(n28626), .ZN(n26698) );
  OAI22_X1 U34942 ( .A1(n26977), .A2(n26698), .B1(n29513), .B2(n28623), .ZN(
        n26699) );
  INV_X1 U34943 ( .A(n28618), .ZN(n26979) );
  INV_X1 U34944 ( .A(n28614), .ZN(n29508) );
  NAND3_X1 U34945 ( .A1(n26979), .A2(n29531), .A3(n29515), .ZN(n26703) );
  NAND3_X1 U34946 ( .A1(n29505), .A2(n28615), .A3(n28626), .ZN(n26702) );
  NOR2_X1 U34947 ( .A1(n29508), .A2(n398), .ZN(n28628) );
  NAND3_X1 U34948 ( .A1(n26983), .A2(n29507), .A3(n28628), .ZN(n26701) );
  NOR2_X1 U34950 ( .A1(n30581), .A2(n31033), .ZN(n26706) );
  OR2_X1 U34951 ( .A1(n31816), .A2(n31821), .ZN(n26705) );
  AOI22_X1 U34952 ( .A1(n26707), .A2(n31034), .B1(n26706), .B2(n26705), .ZN(
        n26716) );
  OR2_X1 U34953 ( .A1(n31816), .A2(n31826), .ZN(n26708) );
  NOR2_X1 U34954 ( .A1(n31815), .A2(n50986), .ZN(n31827) );
  AND2_X1 U34955 ( .A1(n26710), .A2(n26709), .ZN(n26715) );
  NOR2_X1 U34956 ( .A1(n31816), .A2(n30846), .ZN(n30582) );
  INV_X1 U34957 ( .A(n26711), .ZN(n31043) );
  AND2_X1 U34958 ( .A1(n31816), .A2(n31043), .ZN(n26712) );
  AOI22_X1 U34959 ( .A1(n30579), .A2(n30582), .B1(n26712), .B2(n31038), .ZN(
        n26714) );
  XNOR2_X1 U34960 ( .A(n26718), .B(n26717), .ZN(n26719) );
  XNOR2_X1 U34961 ( .A(n32340), .B(n26719), .ZN(n27082) );
  NOR2_X1 U34962 ( .A1(n27840), .A2(n29438), .ZN(n26721) );
  INV_X1 U34963 ( .A(n27834), .ZN(n26720) );
  NAND2_X1 U34964 ( .A1(n27037), .A2(n29448), .ZN(n27842) );
  NOR2_X1 U34965 ( .A1(n26722), .A2(n27038), .ZN(n26724) );
  INV_X1 U34966 ( .A(n27840), .ZN(n27026) );
  INV_X1 U34967 ( .A(n26723), .ZN(n29444) );
  NOR2_X1 U34968 ( .A1(n26069), .A2(n29438), .ZN(n26725) );
  NOR2_X1 U34969 ( .A1(n27828), .A2(n26725), .ZN(n26728) );
  NAND2_X1 U34970 ( .A1(n29446), .A2(n747), .ZN(n27029) );
  OAI21_X1 U34971 ( .B1(n26069), .B2(n27829), .A(n27029), .ZN(n26726) );
  AND2_X1 U34972 ( .A1(n29447), .A2(n26068), .ZN(n27039) );
  AOI22_X1 U34973 ( .A1(n26728), .A2(n26727), .B1(n26726), .B2(n27039), .ZN(
        n26729) );
  INV_X1 U34974 ( .A(n31683), .ZN(n26795) );
  OR2_X1 U34975 ( .A1(n29408), .A2(n27711), .ZN(n27716) );
  AOI22_X1 U34976 ( .A1(n29428), .A2(n26989), .B1(n26985), .B2(n27711), .ZN(
        n26730) );
  MUX2_X1 U34977 ( .A(n27716), .B(n26730), .S(n27710), .Z(n26741) );
  OR2_X1 U34978 ( .A1(n26731), .A2(n51678), .ZN(n29417) );
  INV_X1 U34979 ( .A(n26733), .ZN(n26735) );
  OAI211_X1 U34980 ( .C1(n29411), .C2(n29418), .A(n27711), .B(n26905), .ZN(
        n26736) );
  INV_X1 U34981 ( .A(n26737), .ZN(n26739) );
  NOR2_X1 U34982 ( .A1(n29410), .A2(n27711), .ZN(n26738) );
  OAI21_X1 U34983 ( .B1(n26739), .B2(n26738), .A(n29426), .ZN(n26740) );
  INV_X1 U34984 ( .A(n26949), .ZN(n26877) );
  OAI21_X1 U34985 ( .B1(n26743), .B2(n26742), .A(n26877), .ZN(n26745) );
  OAI21_X1 U34986 ( .B1(n27669), .B2(n27070), .A(n27071), .ZN(n26744) );
  NAND3_X1 U34987 ( .A1(n27656), .A2(n3765), .A3(n26944), .ZN(n26749) );
  OAI22_X1 U34988 ( .A1(n27670), .A2(n27665), .B1(n27669), .B2(n26871), .ZN(
        n26746) );
  AND2_X1 U34989 ( .A1(n27662), .A2(n51117), .ZN(n27672) );
  NAND2_X1 U34990 ( .A1(n26746), .A2(n27672), .ZN(n26748) );
  NOR2_X1 U34991 ( .A1(n51117), .A2(n2642), .ZN(n26747) );
  AND2_X1 U34992 ( .A1(n2098), .A2(n31680), .ZN(n30980) );
  AND2_X1 U34993 ( .A1(n29542), .A2(n29559), .ZN(n27694) );
  INV_X1 U34994 ( .A(n27694), .ZN(n26751) );
  NOR2_X1 U34995 ( .A1(n26751), .A2(n26750), .ZN(n26752) );
  INV_X1 U34996 ( .A(n29563), .ZN(n26754) );
  OAI21_X1 U34997 ( .B1(n29542), .B2(n51111), .A(n29554), .ZN(n26755) );
  NAND2_X1 U34998 ( .A1(n26760), .A2(n29543), .ZN(n26758) );
  AND2_X1 U34999 ( .A1(n27053), .A2(n26756), .ZN(n29547) );
  NAND3_X1 U35000 ( .A1(n29547), .A2(n29557), .A3(n27056), .ZN(n26757) );
  NAND2_X1 U35001 ( .A1(n27694), .A2(n27053), .ZN(n26762) );
  NAND3_X1 U35002 ( .A1(n26763), .A2(n29556), .A3(n26762), .ZN(n26768) );
  NAND2_X1 U35003 ( .A1(n26764), .A2(n29551), .ZN(n26767) );
  NAND3_X1 U35004 ( .A1(n29551), .A2(n27695), .A3(n29564), .ZN(n26766) );
  NOR2_X1 U35005 ( .A1(n29554), .A2(n29555), .ZN(n27700) );
  NAND2_X1 U35006 ( .A1(n27700), .A2(n27697), .ZN(n26765) );
  NAND4_X1 U35007 ( .A1(n26768), .A2(n26767), .A3(n26766), .A4(n26765), .ZN(
        n26769) );
  OAI21_X1 U35008 ( .B1(n26774), .B2(n26772), .A(n27580), .ZN(n26773) );
  INV_X1 U35009 ( .A(n26774), .ZN(n27683) );
  INV_X1 U35010 ( .A(n26776), .ZN(n26778) );
  NAND2_X1 U35011 ( .A1(n27578), .A2(n27685), .ZN(n26777) );
  NAND2_X1 U35012 ( .A1(n29463), .A2(n29467), .ZN(n27759) );
  OAI21_X1 U35013 ( .B1(n29467), .B2(n29463), .A(n27759), .ZN(n26780) );
  NAND2_X1 U35014 ( .A1(n26780), .A2(n27760), .ZN(n26785) );
  NAND2_X1 U35015 ( .A1(n29471), .A2(n27765), .ZN(n27009) );
  NAND2_X1 U35016 ( .A1(n27009), .A2(n29472), .ZN(n26784) );
  AND2_X1 U35017 ( .A1(n26781), .A2(n29455), .ZN(n26783) );
  INV_X1 U35018 ( .A(n29460), .ZN(n26782) );
  AOI22_X1 U35019 ( .A1(n26785), .A2(n26784), .B1(n26783), .B2(n26782), .ZN(
        n26791) );
  INV_X1 U35020 ( .A(n29468), .ZN(n27014) );
  OAI211_X1 U35021 ( .C1(n27014), .C2(n29471), .A(n26787), .B(n26786), .ZN(
        n26789) );
  NAND2_X1 U35022 ( .A1(n26789), .A2(n27750), .ZN(n26790) );
  OAI21_X1 U35023 ( .B1(n29998), .B2(n30982), .A(n29096), .ZN(n26793) );
  INV_X1 U35024 ( .A(n30983), .ZN(n30016) );
  AOI21_X1 U35025 ( .B1(n30976), .B2(n30016), .A(n30981), .ZN(n26792) );
  AOI21_X1 U35026 ( .B1(n30980), .B2(n26793), .A(n26792), .ZN(n26799) );
  AOI21_X1 U35027 ( .B1(n708), .B2(n29998), .A(n30006), .ZN(n26794) );
  INV_X1 U35028 ( .A(n29096), .ZN(n31679) );
  AND3_X1 U35029 ( .A1(n30982), .A2(n31679), .A3(n2094), .ZN(n29999) );
  AOI21_X1 U35030 ( .B1(n26794), .B2(n30976), .A(n29999), .ZN(n26798) );
  NOR2_X1 U35031 ( .A1(n30003), .A2(n30982), .ZN(n30979) );
  NAND2_X1 U35032 ( .A1(n30979), .A2(n7598), .ZN(n30012) );
  NAND2_X1 U35033 ( .A1(n7598), .A2(n30982), .ZN(n30022) );
  NAND2_X1 U35034 ( .A1(n26796), .A2(n30974), .ZN(n26797) );
  XNOR2_X1 U35035 ( .A(n35589), .B(n4865), .ZN(n26883) );
  NAND2_X1 U35036 ( .A1(n26888), .A2(n2144), .ZN(n27733) );
  INV_X1 U35037 ( .A(n27730), .ZN(n27735) );
  NAND2_X1 U35038 ( .A1(n26891), .A2(n27623), .ZN(n26801) );
  OAI211_X1 U35039 ( .C1(n27733), .C2(n27735), .A(n26801), .B(n26800), .ZN(
        n26802) );
  INV_X1 U35040 ( .A(n26802), .ZN(n26809) );
  INV_X1 U35041 ( .A(n27728), .ZN(n27619) );
  AND2_X1 U35042 ( .A1(n26887), .A2(n26804), .ZN(n26805) );
  OAI21_X1 U35043 ( .B1(n26806), .B2(n27739), .A(n26805), .ZN(n26808) );
  OAI211_X1 U35044 ( .C1(n26891), .C2(n27623), .A(n27735), .B(n26888), .ZN(
        n26807) );
  INV_X1 U35045 ( .A(n31490), .ZN(n29841) );
  NAND2_X1 U35046 ( .A1(n26955), .A2(n27690), .ZN(n26956) );
  MUX2_X1 U35047 ( .A(n26812), .B(n26811), .S(n26810), .Z(n26822) );
  INV_X1 U35048 ( .A(n27580), .ZN(n26816) );
  NAND2_X1 U35049 ( .A1(n26817), .A2(n26816), .ZN(n26821) );
  INV_X1 U35050 ( .A(n26961), .ZN(n26827) );
  NAND3_X1 U35051 ( .A1(n26955), .A2(n26823), .A3(n26954), .ZN(n26824) );
  NAND2_X1 U35052 ( .A1(n26825), .A2(n26824), .ZN(n26826) );
  INV_X1 U35053 ( .A(n26828), .ZN(n29893) );
  INV_X1 U35054 ( .A(n30785), .ZN(n26829) );
  NAND2_X1 U35055 ( .A1(n26830), .A2(n29905), .ZN(n26838) );
  INV_X1 U35056 ( .A(n27408), .ZN(n26831) );
  OAI21_X1 U35057 ( .B1(n29904), .B2(n26831), .A(n29909), .ZN(n26837) );
  OAI21_X1 U35058 ( .B1(n26832), .B2(n29899), .A(n29895), .ZN(n27407) );
  OAI21_X1 U35059 ( .B1(n161), .B2(n29901), .A(n26833), .ZN(n26835) );
  NOR2_X1 U35060 ( .A1(n27407), .A2(n26835), .ZN(n26836) );
  OAI22_X1 U35061 ( .A1(n30751), .A2(n27558), .B1(n51697), .B2(n29915), .ZN(
        n26839) );
  AOI21_X1 U35062 ( .B1(n30766), .B2(n26840), .A(n26839), .ZN(n26847) );
  NAND2_X1 U35063 ( .A1(n51697), .A2(n30771), .ZN(n26841) );
  NAND3_X1 U35064 ( .A1(n26844), .A2(n30755), .A3(n29918), .ZN(n26846) );
  INV_X1 U35065 ( .A(n29916), .ZN(n30770) );
  INV_X1 U35066 ( .A(n26848), .ZN(n26851) );
  INV_X1 U35067 ( .A(n26849), .ZN(n26850) );
  NOR3_X1 U35068 ( .A1(n31490), .A2(n26851), .A3(n26850), .ZN(n26880) );
  MUX2_X1 U35069 ( .A(n27602), .B(n30663), .S(n27608), .Z(n26854) );
  NAND2_X1 U35070 ( .A1(n27604), .A2(n30662), .ZN(n26852) );
  OAI211_X1 U35071 ( .C1(n26854), .C2(n30669), .A(n26853), .B(n26852), .ZN(
        n26858) );
  NAND2_X1 U35072 ( .A1(n26856), .A2(n26855), .ZN(n26857) );
  NAND2_X1 U35073 ( .A1(n26858), .A2(n26857), .ZN(n26868) );
  NOR2_X1 U35074 ( .A1(n26859), .A2(n27608), .ZN(n26913) );
  INV_X1 U35075 ( .A(n26860), .ZN(n26861) );
  AOI21_X1 U35076 ( .B1(n26913), .B2(n3819), .A(n26861), .ZN(n26867) );
  NAND2_X1 U35077 ( .A1(n30658), .A2(n3819), .ZN(n26863) );
  OAI21_X1 U35078 ( .B1(n27602), .B2(n30665), .A(n27605), .ZN(n26862) );
  MUX2_X1 U35079 ( .A(n26863), .B(n26862), .S(n30661), .Z(n26866) );
  NAND2_X1 U35080 ( .A1(n26920), .A2(n26864), .ZN(n26865) );
  NAND4_X2 U35081 ( .A1(n26868), .A2(n26867), .A3(n26866), .A4(n26865), .ZN(
        n31496) );
  AND2_X1 U35082 ( .A1(n26870), .A2(n26869), .ZN(n26875) );
  INV_X1 U35083 ( .A(n26871), .ZN(n27658) );
  NAND2_X1 U35084 ( .A1(n51117), .A2(n27652), .ZN(n26872) );
  OAI211_X1 U35085 ( .C1(n27665), .C2(n26944), .A(n27658), .B(n26872), .ZN(
        n26873) );
  AOI21_X1 U35086 ( .B1(n27069), .B2(n26878), .A(n27661), .ZN(n26879) );
  OAI21_X1 U35087 ( .B1(n26880), .B2(n30110), .A(n29837), .ZN(n26881) );
  NAND2_X1 U35088 ( .A1(n30102), .A2(n31273), .ZN(n30998) );
  NAND3_X1 U35089 ( .A1(n31497), .A2(n30102), .A3(n31490), .ZN(n30990) );
  NAND2_X1 U35091 ( .A1(n26882), .A2(n29841), .ZN(n31500) );
  XNOR2_X1 U35092 ( .A(n26883), .B(n36857), .ZN(n27081) );
  INV_X1 U35093 ( .A(n27721), .ZN(n26884) );
  AND2_X1 U35094 ( .A1(n597), .A2(n27732), .ZN(n27636) );
  NAND2_X1 U35095 ( .A1(n27636), .A2(n27632), .ZN(n27628) );
  INV_X1 U35096 ( .A(n26890), .ZN(n27639) );
  NAND2_X1 U35098 ( .A1(n26886), .A2(n26885), .ZN(n26897) );
  NAND2_X1 U35099 ( .A1(n27621), .A2(n597), .ZN(n27724) );
  INV_X1 U35100 ( .A(n26887), .ZN(n27736) );
  AND3_X1 U35101 ( .A1(n27726), .A2(n27724), .A3(n26889), .ZN(n26896) );
  NAND3_X1 U35102 ( .A1(n26890), .A2(n27618), .A3(n597), .ZN(n27727) );
  NAND3_X1 U35103 ( .A1(n27641), .A2(n26891), .A3(n27720), .ZN(n26892) );
  AND2_X1 U35104 ( .A1(n27727), .A2(n26892), .ZN(n26895) );
  INV_X1 U35105 ( .A(n27733), .ZN(n27615) );
  NOR2_X1 U35106 ( .A1(n27728), .A2(n2144), .ZN(n26893) );
  OAI21_X1 U35107 ( .B1(n27615), .B2(n26893), .A(n27719), .ZN(n26894) );
  OAI21_X1 U35108 ( .B1(n7362), .B2(n51678), .A(n29422), .ZN(n26898) );
  NAND3_X1 U35109 ( .A1(n29408), .A2(n26898), .A3(n29424), .ZN(n26899) );
  NAND3_X1 U35110 ( .A1(n26900), .A2(n26899), .A3(n2115), .ZN(n26903) );
  INV_X1 U35111 ( .A(n27706), .ZN(n29420) );
  INV_X1 U35114 ( .A(n26985), .ZN(n29412) );
  OR2_X1 U35115 ( .A1(n26904), .A2(n29412), .ZN(n29432) );
  OAI21_X1 U35116 ( .B1(n27714), .B2(n27717), .A(n29411), .ZN(n26907) );
  NAND3_X1 U35117 ( .A1(n27706), .A2(n29410), .A3(n27710), .ZN(n26906) );
  NAND4_X2 U35118 ( .A1(n26908), .A2(n29432), .A3(n26907), .A4(n26906), .ZN(
        n29591) );
  INV_X1 U35119 ( .A(n26909), .ZN(n26910) );
  NOR2_X1 U35120 ( .A1(n30664), .A2(n27604), .ZN(n27610) );
  NAND2_X1 U35121 ( .A1(n26914), .A2(n3819), .ZN(n26919) );
  OAI21_X1 U35122 ( .B1(n27600), .B2(n27604), .A(n27608), .ZN(n26916) );
  INV_X1 U35123 ( .A(n27601), .ZN(n26915) );
  OAI211_X1 U35125 ( .C1(n27610), .C2(n26919), .A(n30663), .B(n26917), .ZN(
        n26923) );
  NAND2_X1 U35126 ( .A1(n30667), .A2(n27609), .ZN(n26918) );
  NAND4_X1 U35127 ( .A1(n26919), .A2(n30673), .A3(n27608), .A4(n26918), .ZN(
        n26922) );
  INV_X1 U35128 ( .A(n30661), .ZN(n30671) );
  NAND2_X1 U35129 ( .A1(n26920), .A2(n30671), .ZN(n26921) );
  NAND2_X1 U35130 ( .A1(n29591), .A2(n31110), .ZN(n31112) );
  NAND2_X1 U35131 ( .A1(n29917), .A2(n30755), .ZN(n26925) );
  INV_X1 U35132 ( .A(n30763), .ZN(n26926) );
  AOI21_X1 U35133 ( .B1(n26926), .B2(n5769), .A(n27555), .ZN(n26927) );
  OAI21_X1 U35135 ( .B1(n26929), .B2(n26930), .A(n27558), .ZN(n26931) );
  INV_X1 U35136 ( .A(n27671), .ZN(n26946) );
  NAND3_X1 U35137 ( .A1(n26933), .A2(n26946), .A3(n8290), .ZN(n26943) );
  AOI21_X1 U35138 ( .B1(n27662), .B2(n24774), .A(n748), .ZN(n26935) );
  NAND2_X1 U35139 ( .A1(n24774), .A2(n51117), .ZN(n26934) );
  OAI211_X1 U35140 ( .C1(n26945), .C2(n51117), .A(n26935), .B(n26934), .ZN(
        n26936) );
  NAND2_X1 U35141 ( .A1(n26936), .A2(n27071), .ZN(n26942) );
  NOR2_X1 U35142 ( .A1(n27671), .A2(n26937), .ZN(n26938) );
  OAI21_X1 U35143 ( .B1(n26939), .B2(n26938), .A(n27672), .ZN(n26941) );
  NAND2_X1 U35144 ( .A1(n27657), .A2(n8290), .ZN(n26953) );
  OAI21_X1 U35145 ( .B1(n26946), .B2(n27065), .A(n27068), .ZN(n26947) );
  OAI21_X1 U35146 ( .B1(n26949), .B2(n27665), .A(n26948), .ZN(n26951) );
  NAND2_X1 U35148 ( .A1(n26955), .A2(n26954), .ZN(n27688) );
  OR2_X1 U35150 ( .A1(n26960), .A2(n1484), .ZN(n27687) );
  INV_X1 U35151 ( .A(n26957), .ZN(n26958) );
  INV_X1 U35153 ( .A(n26962), .ZN(n26963) );
  OAI21_X1 U35154 ( .B1(n27577), .B2(n27678), .A(n26963), .ZN(n26965) );
  AOI21_X1 U35155 ( .B1(n6290), .B2(n27576), .A(n27685), .ZN(n26964) );
  MUX2_X1 U35156 ( .A(n26965), .B(n26964), .S(n27580), .Z(n26966) );
  INV_X1 U35157 ( .A(n31114), .ZN(n29592) );
  NAND2_X1 U35158 ( .A1(n29584), .A2(n29591), .ZN(n26968) );
  OR2_X1 U35159 ( .A1(n30941), .A2(n31112), .ZN(n31121) );
  NOR2_X1 U35160 ( .A1(n52121), .A2(n362), .ZN(n31117) );
  NAND2_X1 U35162 ( .A1(n51742), .A2(n623), .ZN(n30947) );
  NAND2_X1 U35163 ( .A1(n31115), .A2(n362), .ZN(n31105) );
  NAND4_X1 U35164 ( .A1(n29587), .A2(n29588), .A3(n30947), .A4(n31105), .ZN(
        n26971) );
  NAND2_X1 U35165 ( .A1(n29584), .A2(n362), .ZN(n30057) );
  NAND3_X1 U35167 ( .A1(n30072), .A2(n29584), .A3(n30941), .ZN(n26970) );
  MUX2_X1 U35168 ( .A(n26971), .B(n26970), .S(n29591), .Z(n26972) );
  NAND3_X1 U35169 ( .A1(n29525), .A2(n29526), .A3(n29535), .ZN(n26975) );
  AND2_X1 U35170 ( .A1(n51747), .A2(n28626), .ZN(n28617) );
  AOI22_X1 U35171 ( .A1(n29509), .A2(n28617), .B1(n26979), .B2(n29518), .ZN(
        n29506) );
  NOR2_X1 U35172 ( .A1(n29521), .A2(n29534), .ZN(n26982) );
  INV_X1 U35173 ( .A(n26980), .ZN(n29529) );
  AND2_X1 U35174 ( .A1(n29529), .A2(n29518), .ZN(n26981) );
  OAI21_X1 U35175 ( .B1(n26982), .B2(n26981), .A(n29509), .ZN(n26984) );
  INV_X1 U35176 ( .A(n26983), .ZN(n29524) );
  INV_X1 U35177 ( .A(n29521), .ZN(n29514) );
  NAND2_X1 U35178 ( .A1(n27706), .A2(n7362), .ZN(n26988) );
  INV_X1 U35179 ( .A(n26731), .ZN(n26986) );
  NAND2_X1 U35180 ( .A1(n26986), .A2(n26985), .ZN(n26987) );
  OAI211_X1 U35181 ( .C1(n26997), .C2(n26989), .A(n26988), .B(n26987), .ZN(
        n26990) );
  INV_X1 U35182 ( .A(n26990), .ZN(n27003) );
  INV_X1 U35183 ( .A(n26991), .ZN(n26992) );
  OAI22_X1 U35184 ( .A1(n29410), .A2(n2115), .B1(n26992), .B2(n27710), .ZN(
        n26993) );
  NAND2_X1 U35185 ( .A1(n26993), .A2(n29426), .ZN(n27002) );
  NAND2_X1 U35187 ( .A1(n29412), .A2(n29424), .ZN(n26995) );
  OAI211_X1 U35188 ( .C1(n26996), .C2(n29413), .A(n26995), .B(n29410), .ZN(
        n27001) );
  OAI21_X1 U35189 ( .B1(n29412), .B2(n26998), .A(n26997), .ZN(n26999) );
  NAND2_X1 U35190 ( .A1(n26999), .A2(n29410), .ZN(n27000) );
  AOI21_X1 U35191 ( .B1(n29455), .B2(n27760), .A(n27759), .ZN(n27004) );
  NAND2_X1 U35192 ( .A1(n29472), .A2(n29471), .ZN(n27017) );
  NAND2_X1 U35193 ( .A1(n27004), .A2(n27017), .ZN(n27005) );
  AND2_X1 U35194 ( .A1(n27005), .A2(n8739), .ZN(n27022) );
  INV_X1 U35195 ( .A(n29457), .ZN(n27006) );
  INV_X1 U35196 ( .A(n27007), .ZN(n27008) );
  AND2_X1 U35197 ( .A1(n29455), .A2(n27008), .ZN(n27011) );
  INV_X1 U35198 ( .A(n27009), .ZN(n27010) );
  NAND2_X1 U35199 ( .A1(n29460), .A2(n29463), .ZN(n29466) );
  NAND2_X1 U35200 ( .A1(n27012), .A2(n29457), .ZN(n27013) );
  NAND4_X1 U35201 ( .A1(n29466), .A2(n29462), .A3(n27014), .A4(n27013), .ZN(
        n27020) );
  NAND3_X1 U35202 ( .A1(n27015), .A2(n29456), .A3(n29467), .ZN(n27016) );
  NAND2_X1 U35203 ( .A1(n27017), .A2(n27016), .ZN(n27018) );
  NAND2_X1 U35204 ( .A1(n27018), .A2(n29468), .ZN(n27019) );
  NAND2_X1 U35205 ( .A1(n31347), .A2(n31340), .ZN(n27074) );
  INV_X1 U35206 ( .A(n27023), .ZN(n30051) );
  NAND4_X1 U35207 ( .A1(n27026), .A2(n6602), .A3(n26068), .A4(n27025), .ZN(
        n27027) );
  INV_X1 U35210 ( .A(n27034), .ZN(n27837) );
  MUX2_X1 U35211 ( .A(n6602), .B(n27827), .S(n29447), .Z(n27035) );
  NAND2_X1 U35212 ( .A1(n27035), .A2(n26068), .ZN(n27036) );
  OAI211_X1 U35213 ( .C1(n27037), .C2(n27837), .A(n27036), .B(n26722), .ZN(
        n27045) );
  NAND3_X1 U35214 ( .A1(n27039), .A2(n27038), .A3(n29448), .ZN(n27043) );
  NAND3_X1 U35215 ( .A1(n27039), .A2(n29444), .A3(n29441), .ZN(n27042) );
  AND3_X1 U35216 ( .A1(n27043), .A2(n27042), .A3(n27041), .ZN(n27044) );
  NAND2_X1 U35217 ( .A1(n6339), .A2(n29545), .ZN(n27050) );
  OAI22_X1 U35218 ( .A1(n29554), .A2(n27050), .B1(n29542), .B2(n27049), .ZN(
        n27052) );
  NOR2_X1 U35219 ( .A1(n27052), .A2(n27051), .ZN(n27062) );
  OR2_X1 U35220 ( .A1(n29568), .A2(n6339), .ZN(n29558) );
  NAND2_X1 U35221 ( .A1(n29546), .A2(n29558), .ZN(n27055) );
  INV_X1 U35222 ( .A(n27697), .ZN(n27054) );
  NAND3_X1 U35223 ( .A1(n27055), .A2(n27054), .A3(n27053), .ZN(n27061) );
  OAI21_X1 U35225 ( .B1(n26197), .B2(n27058), .A(n27057), .ZN(n27059) );
  NAND2_X1 U35226 ( .A1(n27059), .A2(n29563), .ZN(n27060) );
  NAND2_X1 U35228 ( .A1(n27064), .A2(n29959), .ZN(n27073) );
  INV_X1 U35229 ( .A(n27066), .ZN(n27072) );
  MUX2_X1 U35230 ( .A(n27074), .B(n27073), .S(n31339), .Z(n27080) );
  INV_X1 U35231 ( .A(n31340), .ZN(n30053) );
  INV_X1 U35232 ( .A(n31346), .ZN(n31936) );
  NAND3_X1 U35233 ( .A1(n30037), .A2(n30053), .A3(n31936), .ZN(n31342) );
  INV_X1 U35234 ( .A(n29602), .ZN(n31934) );
  AND2_X1 U35235 ( .A1(n51744), .A2(n31934), .ZN(n30034) );
  NAND2_X1 U35236 ( .A1(n51744), .A2(n29602), .ZN(n29601) );
  NAND2_X1 U35237 ( .A1(n31340), .A2(n31338), .ZN(n31933) );
  INV_X1 U35238 ( .A(n51744), .ZN(n29609) );
  NOR2_X1 U35239 ( .A1(n31933), .A2(n29609), .ZN(n31932) );
  NAND2_X1 U35240 ( .A1(n31931), .A2(n29602), .ZN(n30030) );
  OR2_X1 U35241 ( .A1(n51744), .A2(n31346), .ZN(n29599) );
  OAI21_X1 U35242 ( .B1(n30030), .B2(n29599), .A(n31935), .ZN(n27076) );
  OAI21_X1 U35243 ( .B1(n30054), .B2(n29602), .A(n27076), .ZN(n27077) );
  XNOR2_X1 U35244 ( .A(n27081), .B(n36869), .ZN(n32744) );
  XNOR2_X1 U35245 ( .A(n27082), .B(n32744), .ZN(n28479) );
  AND2_X1 U35246 ( .A1(n2201), .A2(n2815), .ZN(n30305) );
  NAND3_X1 U35247 ( .A1(n30163), .A2(n2201), .A3(n30171), .ZN(n27085) );
  NAND2_X1 U35249 ( .A1(n739), .A2(n30163), .ZN(n27083) );
  NAND4_X1 U35250 ( .A1(n28032), .A2(n30181), .A3(n29137), .A4(n27083), .ZN(
        n27084) );
  NAND4_X1 U35251 ( .A1(n28031), .A2(n28028), .A3(n27085), .A4(n27084), .ZN(
        n27088) );
  NOR2_X1 U35252 ( .A1(n27088), .A2(n27087), .ZN(n27090) );
  OAI21_X1 U35253 ( .B1(n30209), .B2(n733), .A(n29200), .ZN(n27091) );
  NAND4_X1 U35254 ( .A1(n27092), .A2(n29203), .A3(n30210), .A4(n27091), .ZN(
        n27095) );
  INV_X1 U35255 ( .A(n29200), .ZN(n27887) );
  NAND2_X1 U35256 ( .A1(n27876), .A2(n27887), .ZN(n30206) );
  AND2_X1 U35257 ( .A1(n27882), .A2(n30209), .ZN(n30197) );
  NAND2_X1 U35258 ( .A1(n30197), .A2(n29344), .ZN(n27094) );
  AND3_X1 U35259 ( .A1(n27095), .A2(n30206), .A3(n27094), .ZN(n27100) );
  INV_X1 U35260 ( .A(n27097), .ZN(n27096) );
  NAND3_X1 U35261 ( .A1(n27888), .A2(n27096), .A3(n30210), .ZN(n29353) );
  INV_X1 U35262 ( .A(n27886), .ZN(n29342) );
  NOR2_X1 U35263 ( .A1(n29203), .A2(n29342), .ZN(n27098) );
  OAI21_X1 U35264 ( .B1(n27098), .B2(n30203), .A(n30200), .ZN(n27099) );
  OR2_X1 U35265 ( .A1(n51109), .A2(n30191), .ZN(n29204) );
  NAND2_X1 U35267 ( .A1(n29034), .A2(n28536), .ZN(n27101) );
  NOR2_X1 U35268 ( .A1(n28529), .A2(n28530), .ZN(n28159) );
  OAI21_X1 U35269 ( .B1(n28159), .B2(n28879), .A(n29039), .ZN(n27109) );
  NOR2_X1 U35270 ( .A1(n28875), .A2(n28883), .ZN(n27106) );
  OAI21_X1 U35272 ( .B1(n27110), .B2(n30285), .A(n28144), .ZN(n27117) );
  AOI21_X1 U35273 ( .B1(n51748), .B2(n28548), .A(n30285), .ZN(n27112) );
  INV_X1 U35274 ( .A(n27111), .ZN(n28153) );
  OAI21_X1 U35276 ( .B1(n2195), .B2(n30295), .A(n2881), .ZN(n27114) );
  INV_X1 U35277 ( .A(n28590), .ZN(n27120) );
  NOR2_X1 U35278 ( .A1(n28584), .A2(n27120), .ZN(n27124) );
  INV_X1 U35279 ( .A(n28577), .ZN(n28895) );
  OAI21_X1 U35280 ( .B1(n28894), .B2(n27121), .A(n27987), .ZN(n27122) );
  AOI22_X1 U35281 ( .A1(n27124), .A2(n27123), .B1(n28895), .B2(n27122), .ZN(
        n27144) );
  NOR2_X1 U35282 ( .A1(n27994), .A2(n28903), .ZN(n28889) );
  INV_X1 U35283 ( .A(n28894), .ZN(n28904) );
  NOR2_X1 U35284 ( .A1(n27994), .A2(n51118), .ZN(n27127) );
  AOI22_X1 U35285 ( .A1(n28889), .A2(n28904), .B1(n27127), .B2(n27126), .ZN(
        n27143) );
  NAND3_X1 U35286 ( .A1(n27130), .A2(n27128), .A3(n27993), .ZN(n27138) );
  NAND3_X1 U35287 ( .A1(n28905), .A2(n27129), .A3(n27132), .ZN(n27137) );
  NAND3_X1 U35288 ( .A1(n27130), .A2(n28903), .A3(n28894), .ZN(n27136) );
  NOR2_X1 U35289 ( .A1(n28000), .A2(n28587), .ZN(n27134) );
  NAND4_X1 U35290 ( .A1(n27134), .A2(n28897), .A3(n27139), .A4(n27133), .ZN(
        n27135) );
  INV_X1 U35291 ( .A(n27999), .ZN(n27140) );
  NAND3_X1 U35292 ( .A1(n28908), .A2(n28905), .A3(n28894), .ZN(n27141) );
  NAND2_X1 U35294 ( .A1(n5417), .A2(n29155), .ZN(n27956) );
  OAI21_X1 U35295 ( .B1(n29152), .B2(n27145), .A(n29155), .ZN(n27148) );
  NAND3_X1 U35297 ( .A1(n5821), .A2(n5169), .A3(n27957), .ZN(n27149) );
  AND2_X1 U35298 ( .A1(n30247), .A2(n27149), .ZN(n27150) );
  NOR2_X1 U35299 ( .A1(n32500), .A2(n30877), .ZN(n27152) );
  NAND3_X1 U35300 ( .A1(n30879), .A2(n32507), .A3(n32511), .ZN(n32514) );
  AND2_X1 U35301 ( .A1(n30881), .A2(n32503), .ZN(n27154) );
  NAND2_X1 U35303 ( .A1(n32502), .A2(n31986), .ZN(n27153) );
  AND4_X1 U35304 ( .A1(n29675), .A2(n27154), .A3(n32514), .A4(n27153), .ZN(
        n27156) );
  NAND4_X1 U35305 ( .A1(n32500), .A2(n32503), .A3(n32506), .A4(n31995), .ZN(
        n27155) );
  NAND2_X1 U35309 ( .A1(n28807), .A2(n27164), .ZN(n27161) );
  NAND2_X1 U35311 ( .A1(n28810), .A2(n2169), .ZN(n27160) );
  AND2_X1 U35312 ( .A1(n29853), .A2(n27164), .ZN(n29855) );
  NAND2_X1 U35313 ( .A1(n30723), .A2(n30711), .ZN(n27165) );
  NAND3_X1 U35314 ( .A1(n28800), .A2(n28799), .A3(n27165), .ZN(n27166) );
  INV_X1 U35315 ( .A(n30723), .ZN(n27167) );
  NAND3_X1 U35316 ( .A1(n731), .A2(n27167), .A3(n29855), .ZN(n27169) );
  NAND3_X1 U35317 ( .A1(n28801), .A2(n30725), .A3(n2169), .ZN(n27168) );
  OAI21_X1 U35318 ( .B1(n30723), .B2(n2169), .A(n28810), .ZN(n27170) );
  NAND2_X1 U35319 ( .A1(n27170), .A2(n30725), .ZN(n27543) );
  NAND2_X1 U35320 ( .A1(n27588), .A2(n52218), .ZN(n27593) );
  OAI21_X1 U35321 ( .B1(n30712), .B2(n2205), .A(n27593), .ZN(n27171) );
  NAND2_X1 U35322 ( .A1(n27171), .A2(n30719), .ZN(n27544) );
  XNOR2_X1 U35323 ( .A(n28319), .B(n27172), .ZN(n27182) );
  XNOR2_X1 U35324 ( .A(n27173), .B(n46097), .ZN(n40759) );
  XNOR2_X1 U35325 ( .A(n27175), .B(n27174), .ZN(n42908) );
  XNOR2_X1 U35326 ( .A(n40759), .B(n42908), .ZN(n27176) );
  XNOR2_X1 U35327 ( .A(n27177), .B(n27176), .ZN(n27178) );
  XNOR2_X1 U35328 ( .A(n28109), .B(n27178), .ZN(n27181) );
  XNOR2_X1 U35329 ( .A(n28106), .B(n28104), .ZN(n27179) );
  XNOR2_X1 U35330 ( .A(n370), .B(n27179), .ZN(n27180) );
  XNOR2_X1 U35331 ( .A(n27184), .B(n27183), .ZN(n27278) );
  INV_X1 U35332 ( .A(n43713), .ZN(n27187) );
  XNOR2_X1 U35333 ( .A(n27186), .B(n27185), .ZN(n42408) );
  XNOR2_X1 U35334 ( .A(n27187), .B(n42408), .ZN(n27188) );
  XNOR2_X1 U35335 ( .A(n28288), .B(n27188), .ZN(n27189) );
  XNOR2_X1 U35336 ( .A(n27189), .B(n28292), .ZN(n27190) );
  XNOR2_X1 U35337 ( .A(n27190), .B(n27505), .ZN(n27192) );
  XNOR2_X1 U35338 ( .A(n27191), .B(n27192), .ZN(n27193) );
  XNOR2_X1 U35339 ( .A(n28129), .B(n51121), .ZN(n28296) );
  XNOR2_X1 U35340 ( .A(n27193), .B(n28296), .ZN(n27194) );
  NAND2_X1 U35341 ( .A1(n27278), .A2(n28971), .ZN(n29721) );
  XNOR2_X1 U35343 ( .A(n27419), .B(n27199), .ZN(n28063) );
  XNOR2_X1 U35344 ( .A(n27417), .B(n28063), .ZN(n27216) );
  XNOR2_X1 U35345 ( .A(n27200), .B(n28049), .ZN(n27202) );
  XNOR2_X1 U35346 ( .A(n27202), .B(n27201), .ZN(n27214) );
  XNOR2_X1 U35347 ( .A(n27204), .B(n27203), .ZN(n34774) );
  XNOR2_X1 U35348 ( .A(n34774), .B(n27205), .ZN(n42633) );
  INV_X1 U35349 ( .A(n37140), .ZN(n27207) );
  XNOR2_X1 U35350 ( .A(n42101), .B(n4564), .ZN(n27206) );
  XNOR2_X1 U35351 ( .A(n27207), .B(n27206), .ZN(n27208) );
  XNOR2_X1 U35352 ( .A(n42633), .B(n27208), .ZN(n27209) );
  XNOR2_X1 U35353 ( .A(n51751), .B(n27209), .ZN(n27212) );
  XNOR2_X1 U35354 ( .A(n27211), .B(n27212), .ZN(n27213) );
  XNOR2_X1 U35355 ( .A(n27214), .B(n27213), .ZN(n27215) );
  XNOR2_X1 U35356 ( .A(n27216), .B(n27215), .ZN(n27220) );
  XNOR2_X1 U35357 ( .A(n27218), .B(n27217), .ZN(n27219) );
  XNOR2_X1 U35358 ( .A(n27222), .B(n27221), .ZN(n27223) );
  XNOR2_X1 U35359 ( .A(n27224), .B(n27373), .ZN(n27225) );
  XNOR2_X1 U35360 ( .A(n27226), .B(n27227), .ZN(n28279) );
  XNOR2_X1 U35361 ( .A(n27485), .B(n27228), .ZN(n27229) );
  XNOR2_X1 U35362 ( .A(n27230), .B(n27229), .ZN(n42947) );
  XNOR2_X1 U35363 ( .A(n27483), .B(n4296), .ZN(n40520) );
  XNOR2_X1 U35364 ( .A(n42947), .B(n40520), .ZN(n27231) );
  XNOR2_X1 U35365 ( .A(n27232), .B(n27231), .ZN(n27233) );
  XNOR2_X1 U35366 ( .A(n27234), .B(n27233), .ZN(n27237) );
  INV_X1 U35367 ( .A(n27235), .ZN(n27236) );
  XNOR2_X1 U35368 ( .A(n27237), .B(n27236), .ZN(n27238) );
  XNOR2_X1 U35369 ( .A(n28279), .B(n27238), .ZN(n27239) );
  INV_X1 U35370 ( .A(n27240), .ZN(n27255) );
  XNOR2_X1 U35371 ( .A(n27241), .B(n28214), .ZN(n27243) );
  XNOR2_X1 U35372 ( .A(n27242), .B(n27243), .ZN(n27253) );
  XNOR2_X1 U35373 ( .A(n45479), .B(n2600), .ZN(n27246) );
  INV_X1 U35374 ( .A(n27244), .ZN(n27245) );
  XNOR2_X1 U35375 ( .A(n27246), .B(n27245), .ZN(n44162) );
  XNOR2_X1 U35376 ( .A(n27301), .B(n27247), .ZN(n43499) );
  XNOR2_X1 U35377 ( .A(n43499), .B(n6031), .ZN(n27248) );
  XNOR2_X1 U35378 ( .A(n44162), .B(n27248), .ZN(n27249) );
  XNOR2_X1 U35379 ( .A(n28213), .B(n27249), .ZN(n27251) );
  XNOR2_X1 U35380 ( .A(n27250), .B(n27251), .ZN(n27252) );
  XNOR2_X1 U35381 ( .A(n27253), .B(n27252), .ZN(n27254) );
  XNOR2_X1 U35382 ( .A(n27255), .B(n27254), .ZN(n27262) );
  XNOR2_X1 U35383 ( .A(n51483), .B(n27256), .ZN(n27260) );
  XNOR2_X1 U35384 ( .A(n27258), .B(n27439), .ZN(n27259) );
  XNOR2_X1 U35385 ( .A(n27260), .B(n27259), .ZN(n27261) );
  XNOR2_X1 U35386 ( .A(n27262), .B(n27261), .ZN(n27281) );
  NAND2_X1 U35387 ( .A1(n28974), .A2(n28970), .ZN(n28789) );
  XNOR2_X1 U35388 ( .A(n27325), .B(n27265), .ZN(n27266) );
  INV_X1 U35389 ( .A(n27267), .ZN(n27271) );
  XNOR2_X1 U35390 ( .A(n43727), .B(n4869), .ZN(n27268) );
  XNOR2_X1 U35391 ( .A(n42461), .B(n27268), .ZN(n27269) );
  XNOR2_X1 U35392 ( .A(n28353), .B(n27269), .ZN(n27270) );
  XNOR2_X1 U35393 ( .A(n27271), .B(n27270), .ZN(n27273) );
  XNOR2_X1 U35394 ( .A(n27272), .B(n42754), .ZN(n27465) );
  XNOR2_X1 U35395 ( .A(n27273), .B(n27465), .ZN(n27274) );
  XNOR2_X1 U35396 ( .A(n27275), .B(n27274), .ZN(n27276) );
  NAND2_X1 U35397 ( .A1(n28789), .A2(n28187), .ZN(n27277) );
  AOI21_X1 U35398 ( .B1(n29721), .B2(n29724), .A(n27277), .ZN(n27280) );
  INV_X1 U35399 ( .A(n27278), .ZN(n28793) );
  INV_X1 U35400 ( .A(n27281), .ZN(n28177) );
  NOR2_X1 U35401 ( .A1(n29715), .A2(n51342), .ZN(n27279) );
  OAI21_X1 U35402 ( .B1(n27280), .B2(n27279), .A(n28982), .ZN(n27288) );
  AND2_X1 U35403 ( .A1(n28974), .A2(n51108), .ZN(n29722) );
  INV_X1 U35404 ( .A(n28971), .ZN(n30411) );
  NAND3_X1 U35405 ( .A1(n29722), .A2(n28187), .A3(n30411), .ZN(n30405) );
  INV_X1 U35406 ( .A(n30412), .ZN(n30404) );
  NAND2_X1 U35407 ( .A1(n51108), .A2(n28796), .ZN(n28973) );
  NAND2_X1 U35408 ( .A1(n30404), .A2(n28973), .ZN(n27282) );
  AND2_X1 U35409 ( .A1(n30405), .A2(n27282), .ZN(n27287) );
  INV_X1 U35410 ( .A(n28187), .ZN(n28179) );
  NAND2_X1 U35411 ( .A1(n28182), .A2(n28974), .ZN(n27286) );
  INV_X1 U35412 ( .A(n29722), .ZN(n27283) );
  OAI21_X1 U35413 ( .B1(n28789), .B2(n28179), .A(n27283), .ZN(n27284) );
  NAND2_X1 U35414 ( .A1(n28175), .A2(n27284), .ZN(n27285) );
  NAND4_X2 U35415 ( .A1(n27288), .A2(n27287), .A3(n27285), .A4(n27286), .ZN(
        n32785) );
  OR2_X1 U35416 ( .A1(n32791), .A2(n32785), .ZN(n31863) );
  XNOR2_X1 U35417 ( .A(n27289), .B(n27290), .ZN(n27294) );
  XNOR2_X1 U35418 ( .A(n28213), .B(n43073), .ZN(n27292) );
  XNOR2_X1 U35419 ( .A(n27291), .B(n27292), .ZN(n27293) );
  XNOR2_X1 U35420 ( .A(n27294), .B(n27293), .ZN(n28347) );
  XNOR2_X1 U35421 ( .A(n23525), .B(n27295), .ZN(n27305) );
  XNOR2_X1 U35422 ( .A(n27298), .B(n27297), .ZN(n27300) );
  XNOR2_X1 U35423 ( .A(n27300), .B(n27299), .ZN(n45336) );
  XNOR2_X1 U35424 ( .A(n27301), .B(n4827), .ZN(n43986) );
  XNOR2_X1 U35425 ( .A(n45336), .B(n43986), .ZN(n27302) );
  XNOR2_X1 U35426 ( .A(n27303), .B(n27302), .ZN(n27304) );
  XNOR2_X1 U35427 ( .A(n27305), .B(n27304), .ZN(n27308) );
  XNOR2_X1 U35428 ( .A(n27439), .B(n27306), .ZN(n27307) );
  XNOR2_X1 U35429 ( .A(n27309), .B(n27310), .ZN(n27312) );
  XNOR2_X1 U35430 ( .A(n27312), .B(n27311), .ZN(n27444) );
  XNOR2_X1 U35431 ( .A(n27313), .B(n27444), .ZN(n28772) );
  INV_X1 U35432 ( .A(n27314), .ZN(n27327) );
  XNOR2_X1 U35433 ( .A(n49790), .B(n4818), .ZN(n27315) );
  XNOR2_X1 U35434 ( .A(n27316), .B(n27315), .ZN(n44088) );
  XNOR2_X1 U35435 ( .A(n27317), .B(n44088), .ZN(n27320) );
  INV_X1 U35436 ( .A(n27318), .ZN(n27319) );
  XNOR2_X1 U35437 ( .A(n27320), .B(n27319), .ZN(n27321) );
  XNOR2_X1 U35438 ( .A(n27322), .B(n27321), .ZN(n27323) );
  XNOR2_X1 U35439 ( .A(n25176), .B(n27323), .ZN(n27324) );
  XNOR2_X1 U35440 ( .A(n27325), .B(n27324), .ZN(n27326) );
  XNOR2_X1 U35441 ( .A(n27327), .B(n27326), .ZN(n27332) );
  INV_X1 U35442 ( .A(n27328), .ZN(n27329) );
  XNOR2_X1 U35443 ( .A(n27330), .B(n27329), .ZN(n27331) );
  XNOR2_X1 U35445 ( .A(n41161), .B(n41155), .ZN(n33052) );
  XNOR2_X1 U35446 ( .A(n33052), .B(n4937), .ZN(n27333) );
  XNOR2_X1 U35447 ( .A(n24916), .B(n27334), .ZN(n27338) );
  XNOR2_X1 U35448 ( .A(n24856), .B(n28246), .ZN(n27336) );
  XNOR2_X1 U35449 ( .A(n27335), .B(n27336), .ZN(n27337) );
  XNOR2_X1 U35450 ( .A(n27337), .B(n27338), .ZN(n27343) );
  INV_X1 U35451 ( .A(n27339), .ZN(n27340) );
  XNOR2_X1 U35452 ( .A(n27341), .B(n27340), .ZN(n27342) );
  INV_X1 U35453 ( .A(n27344), .ZN(n27345) );
  XNOR2_X1 U35454 ( .A(n27347), .B(n27346), .ZN(n27358) );
  INV_X1 U35455 ( .A(n27348), .ZN(n27350) );
  XNOR2_X1 U35456 ( .A(n27350), .B(n27349), .ZN(n35814) );
  XNOR2_X1 U35457 ( .A(n27351), .B(n4884), .ZN(n27352) );
  XNOR2_X1 U35458 ( .A(n35814), .B(n27352), .ZN(n44025) );
  XNOR2_X1 U35459 ( .A(n27353), .B(n4720), .ZN(n42579) );
  XNOR2_X1 U35460 ( .A(n44025), .B(n42579), .ZN(n27354) );
  XNOR2_X1 U35461 ( .A(n27356), .B(n27355), .ZN(n27357) );
  XNOR2_X1 U35462 ( .A(n27358), .B(n27357), .ZN(n27359) );
  NOR2_X1 U35463 ( .A1(n30379), .A2(n29882), .ZN(n27361) );
  NAND2_X1 U35464 ( .A1(n30375), .A2(n27361), .ZN(n30742) );
  XNOR2_X1 U35465 ( .A(n27363), .B(n27362), .ZN(n27370) );
  XNOR2_X1 U35466 ( .A(n33445), .B(n27364), .ZN(n43166) );
  XNOR2_X1 U35467 ( .A(n1336), .B(n274), .ZN(n27365) );
  XNOR2_X1 U35468 ( .A(n36994), .B(n27365), .ZN(n41817) );
  XNOR2_X1 U35469 ( .A(n41817), .B(n41567), .ZN(n27366) );
  XNOR2_X1 U35470 ( .A(n43166), .B(n27366), .ZN(n27367) );
  XNOR2_X1 U35471 ( .A(n27368), .B(n27367), .ZN(n27369) );
  XNOR2_X1 U35472 ( .A(n27370), .B(n27369), .ZN(n27371) );
  XNOR2_X1 U35473 ( .A(n27373), .B(n75), .ZN(n27375) );
  XNOR2_X1 U35474 ( .A(n27375), .B(n27374), .ZN(n27376) );
  XNOR2_X1 U35475 ( .A(n28276), .B(n27376), .ZN(n27494) );
  XNOR2_X1 U35476 ( .A(n27377), .B(n27494), .ZN(n27378) );
  INV_X1 U35477 ( .A(n27379), .ZN(n29784) );
  AND2_X1 U35478 ( .A1(n28772), .A2(n29882), .ZN(n28767) );
  NAND2_X1 U35479 ( .A1(n29784), .A2(n30374), .ZN(n29880) );
  NAND2_X1 U35480 ( .A1(n28767), .A2(n29880), .ZN(n27380) );
  INV_X1 U35482 ( .A(n30374), .ZN(n29883) );
  NAND2_X1 U35483 ( .A1(n30379), .A2(n29883), .ZN(n27400) );
  OAI22_X1 U35484 ( .A1(n30379), .A2(n29780), .B1(n28771), .B2(n52181), .ZN(
        n27399) );
  INV_X1 U35485 ( .A(n27381), .ZN(n27398) );
  XNOR2_X1 U35486 ( .A(n27450), .B(n27382), .ZN(n27383) );
  XNOR2_X1 U35487 ( .A(n27384), .B(n27383), .ZN(n27395) );
  INV_X1 U35488 ( .A(n27385), .ZN(n27386) );
  XNOR2_X1 U35489 ( .A(n27386), .B(n4517), .ZN(n41844) );
  XNOR2_X1 U35490 ( .A(n27388), .B(n27387), .ZN(n27389) );
  XNOR2_X1 U35491 ( .A(n27390), .B(n27389), .ZN(n43120) );
  XNOR2_X1 U35492 ( .A(n41844), .B(n43120), .ZN(n27391) );
  XNOR2_X1 U35493 ( .A(n27451), .B(n27391), .ZN(n27392) );
  XNOR2_X1 U35494 ( .A(n2164), .B(n27392), .ZN(n27394) );
  XNOR2_X2 U35495 ( .A(n27398), .B(n27397), .ZN(n30376) );
  NOR2_X1 U35496 ( .A1(n29780), .A2(n30376), .ZN(n30381) );
  INV_X1 U35497 ( .A(n27400), .ZN(n27401) );
  NAND2_X1 U35498 ( .A1(n30381), .A2(n27401), .ZN(n27405) );
  NOR2_X1 U35499 ( .A1(n30733), .A2(n1121), .ZN(n30366) );
  AND2_X1 U35500 ( .A1(n28772), .A2(n742), .ZN(n30740) );
  NOR2_X1 U35501 ( .A1(n29774), .A2(n30379), .ZN(n30741) );
  AOI21_X1 U35502 ( .B1(n30366), .B2(n30740), .A(n30741), .ZN(n27404) );
  INV_X1 U35503 ( .A(n30360), .ZN(n29886) );
  NOR2_X1 U35504 ( .A1(n29880), .A2(n30376), .ZN(n30731) );
  NAND2_X1 U35505 ( .A1(n30731), .A2(n30740), .ZN(n27403) );
  INV_X1 U35506 ( .A(n27407), .ZN(n27416) );
  NOR2_X1 U35507 ( .A1(n27409), .A2(n29893), .ZN(n27410) );
  NAND2_X1 U35508 ( .A1(n27411), .A2(n27410), .ZN(n27414) );
  OAI22_X1 U35509 ( .A1(n29892), .A2(n27566), .B1(n29900), .B2(n30791), .ZN(
        n27412) );
  NAND2_X1 U35510 ( .A1(n27412), .A2(n29902), .ZN(n27413) );
  NAND4_X2 U35511 ( .A1(n27415), .A2(n27416), .A3(n27414), .A4(n27413), .ZN(
        n31725) );
  XNOR2_X1 U35512 ( .A(n27417), .B(n27418), .ZN(n27429) );
  XNOR2_X1 U35513 ( .A(n27420), .B(n27421), .ZN(n27427) );
  XNOR2_X1 U35514 ( .A(n43370), .B(n43368), .ZN(n27422) );
  XNOR2_X1 U35515 ( .A(n34601), .B(n27422), .ZN(n27423) );
  XNOR2_X1 U35516 ( .A(n27424), .B(n27423), .ZN(n27425) );
  XNOR2_X1 U35517 ( .A(n27427), .B(n27426), .ZN(n27428) );
  XNOR2_X1 U35518 ( .A(n27428), .B(n27429), .ZN(n27432) );
  INV_X1 U35519 ( .A(n27430), .ZN(n27431) );
  INV_X1 U35520 ( .A(n33287), .ZN(n27436) );
  INV_X1 U35521 ( .A(n27433), .ZN(n45480) );
  XNOR2_X1 U35522 ( .A(n45480), .B(n27434), .ZN(n27435) );
  XNOR2_X1 U35523 ( .A(n27436), .B(n27435), .ZN(n27437) );
  XNOR2_X1 U35524 ( .A(n28221), .B(n27437), .ZN(n27438) );
  XNOR2_X1 U35525 ( .A(n28223), .B(n27438), .ZN(n27442) );
  XNOR2_X1 U35526 ( .A(n27440), .B(n27439), .ZN(n27441) );
  XNOR2_X1 U35527 ( .A(n27442), .B(n27441), .ZN(n27443) );
  XNOR2_X1 U35528 ( .A(n28302), .B(n27445), .ZN(n27449) );
  XNOR2_X1 U35529 ( .A(n27447), .B(n27446), .ZN(n27448) );
  XNOR2_X1 U35530 ( .A(n27451), .B(n27450), .ZN(n28107) );
  XNOR2_X1 U35531 ( .A(n28107), .B(n27452), .ZN(n27461) );
  INV_X1 U35532 ( .A(n27453), .ZN(n27455) );
  XNOR2_X1 U35533 ( .A(n27455), .B(n27454), .ZN(n43223) );
  XNOR2_X1 U35534 ( .A(n41597), .B(n4517), .ZN(n27456) );
  XNOR2_X1 U35535 ( .A(n43223), .B(n27456), .ZN(n27457) );
  XNOR2_X1 U35536 ( .A(n28427), .B(n27457), .ZN(n27458) );
  XNOR2_X1 U35537 ( .A(n370), .B(n27458), .ZN(n27460) );
  XNOR2_X1 U35538 ( .A(n27461), .B(n27460), .ZN(n27462) );
  INV_X1 U35539 ( .A(n27463), .ZN(n27464) );
  INV_X1 U35540 ( .A(n27465), .ZN(n27466) );
  XNOR2_X1 U35541 ( .A(n27467), .B(n27466), .ZN(n27468) );
  XNOR2_X1 U35542 ( .A(n27469), .B(n27468), .ZN(n27478) );
  INV_X1 U35543 ( .A(n27470), .ZN(n27471) );
  XNOR2_X1 U35544 ( .A(n27471), .B(n42755), .ZN(n27472) );
  XNOR2_X1 U35545 ( .A(n51749), .B(n27472), .ZN(n27474) );
  XNOR2_X1 U35546 ( .A(n27474), .B(n27473), .ZN(n27476) );
  XNOR2_X1 U35547 ( .A(n27477), .B(n28353), .ZN(n28230) );
  XNOR2_X1 U35548 ( .A(n27482), .B(n27481), .ZN(n27493) );
  XNOR2_X1 U35549 ( .A(n27484), .B(n27483), .ZN(n42125) );
  XNOR2_X1 U35550 ( .A(n27485), .B(n4706), .ZN(n43189) );
  XNOR2_X1 U35551 ( .A(n42769), .B(n4482), .ZN(n27486) );
  XNOR2_X1 U35552 ( .A(n43189), .B(n27486), .ZN(n27487) );
  XNOR2_X1 U35553 ( .A(n42125), .B(n27487), .ZN(n27488) );
  XNOR2_X1 U35554 ( .A(n51415), .B(n27488), .ZN(n27490) );
  XNOR2_X1 U35555 ( .A(n27491), .B(n27490), .ZN(n27492) );
  XNOR2_X1 U35556 ( .A(n27492), .B(n27493), .ZN(n27497) );
  INV_X1 U35557 ( .A(n27494), .ZN(n27496) );
  XNOR2_X1 U35558 ( .A(n42721), .B(n4618), .ZN(n27498) );
  XNOR2_X1 U35559 ( .A(n43620), .B(n27498), .ZN(n27499) );
  XNOR2_X1 U35560 ( .A(n42723), .B(n27499), .ZN(n27500) );
  XNOR2_X1 U35561 ( .A(n27501), .B(n27500), .ZN(n27503) );
  XNOR2_X1 U35562 ( .A(n27503), .B(n27502), .ZN(n27504) );
  XNOR2_X1 U35563 ( .A(n27504), .B(n28129), .ZN(n27508) );
  XNOR2_X1 U35564 ( .A(n27506), .B(n27505), .ZN(n27507) );
  XNOR2_X1 U35565 ( .A(n27508), .B(n27507), .ZN(n27510) );
  XNOR2_X1 U35566 ( .A(n27510), .B(n27509), .ZN(n27512) );
  NAND3_X1 U35567 ( .A1(n27515), .A2(n27514), .A3(n27513), .ZN(n27522) );
  NOR2_X1 U35568 ( .A1(n29868), .A2(n30434), .ZN(n28737) );
  NAND2_X1 U35570 ( .A1(n28737), .A2(n29873), .ZN(n27521) );
  NAND2_X1 U35571 ( .A1(n29867), .A2(n28333), .ZN(n30436) );
  NOR2_X1 U35572 ( .A1(n30436), .A2(n487), .ZN(n27516) );
  AOI22_X1 U35573 ( .A1(n27516), .A2(n29700), .B1(n29869), .B2(n30434), .ZN(
        n27520) );
  NAND2_X1 U35574 ( .A1(n28738), .A2(n28333), .ZN(n29698) );
  NAND2_X1 U35575 ( .A1(n486), .A2(n28333), .ZN(n27517) );
  NAND2_X1 U35576 ( .A1(n27518), .A2(n29692), .ZN(n27519) );
  NAND3_X1 U35577 ( .A1(n31863), .A2(n32778), .A3(n32286), .ZN(n27535) );
  NAND2_X1 U35578 ( .A1(n24091), .A2(n28758), .ZN(n27523) );
  MUX2_X1 U35579 ( .A(n28758), .B(n27523), .S(n30699), .Z(n27524) );
  NAND2_X1 U35580 ( .A1(n27524), .A2(n6253), .ZN(n27533) );
  AND2_X1 U35581 ( .A1(n30692), .A2(n30683), .ZN(n29932) );
  AOI21_X1 U35582 ( .B1(n30685), .B2(n30392), .A(n29932), .ZN(n27532) );
  INV_X1 U35583 ( .A(n30690), .ZN(n27526) );
  OAI21_X1 U35584 ( .B1(n30391), .B2(n27526), .A(n30398), .ZN(n27527) );
  NAND2_X1 U35585 ( .A1(n27527), .A2(n30687), .ZN(n27531) );
  NAND3_X1 U35589 ( .A1(n32787), .A2(n32151), .A3(n32788), .ZN(n27534) );
  NAND2_X1 U35590 ( .A1(n27535), .A2(n27534), .ZN(n33114) );
  NAND2_X1 U35591 ( .A1(n32157), .A2(n32785), .ZN(n32789) );
  INV_X1 U35592 ( .A(n32778), .ZN(n32149) );
  INV_X1 U35593 ( .A(n32151), .ZN(n27536) );
  NAND2_X1 U35594 ( .A1(n32149), .A2(n27536), .ZN(n32162) );
  XNOR2_X1 U35595 ( .A(n32157), .B(n32788), .ZN(n27537) );
  AOI22_X1 U35596 ( .A1(n32791), .A2(n27537), .B1(n32788), .B2(n32785), .ZN(
        n27538) );
  OAI211_X1 U35597 ( .C1(n32791), .C2(n32789), .A(n32162), .B(n27538), .ZN(
        n33115) );
  INV_X1 U35598 ( .A(n32787), .ZN(n32284) );
  NAND2_X1 U35599 ( .A1(n32284), .A2(n32785), .ZN(n32150) );
  INV_X1 U35600 ( .A(n27539), .ZN(n27540) );
  NAND3_X1 U35601 ( .A1(n4759), .A2(n27541), .A3(n27540), .ZN(n27547) );
  INV_X1 U35602 ( .A(n27542), .ZN(n27545) );
  OAI21_X1 U35603 ( .B1(n27547), .B2(n27546), .A(n32788), .ZN(n32794) );
  NAND2_X1 U35604 ( .A1(n32150), .A2(n32794), .ZN(n31862) );
  INV_X1 U35605 ( .A(n27548), .ZN(n27551) );
  INV_X1 U35606 ( .A(n27549), .ZN(n27550) );
  NAND3_X1 U35607 ( .A1(n27551), .A2(n27550), .A3(n32785), .ZN(n31864) );
  INV_X1 U35608 ( .A(n32785), .ZN(n32798) );
  NAND2_X1 U35609 ( .A1(n32798), .A2(n32788), .ZN(n31733) );
  AND2_X1 U35610 ( .A1(n31864), .A2(n31733), .ZN(n32166) );
  NOR2_X1 U35611 ( .A1(n32787), .A2(n32791), .ZN(n32163) );
  AOI21_X1 U35612 ( .B1(n32163), .B2(n32286), .A(n31725), .ZN(n27552) );
  OAI21_X1 U35613 ( .B1(n31862), .B2(n32166), .A(n27552), .ZN(n33116) );
  OAI21_X1 U35614 ( .B1(n33114), .B2(n33115), .A(n33116), .ZN(n27553) );
  NAND2_X1 U35615 ( .A1(n51696), .A2(n1676), .ZN(n27554) );
  INV_X1 U35616 ( .A(n29917), .ZN(n30759) );
  NAND2_X1 U35617 ( .A1(n30759), .A2(n30763), .ZN(n27559) );
  NAND3_X1 U35618 ( .A1(n27560), .A2(n27559), .A3(n27558), .ZN(n27563) );
  NAND3_X1 U35619 ( .A1(n30772), .A2(n30770), .A3(n738), .ZN(n27561) );
  INV_X1 U35620 ( .A(n29909), .ZN(n27564) );
  NAND3_X1 U35621 ( .A1(n30788), .A2(n27566), .A3(n23658), .ZN(n27567) );
  OAI21_X1 U35622 ( .B1(n30785), .B2(n30790), .A(n27567), .ZN(n27568) );
  NAND2_X1 U35623 ( .A1(n23658), .A2(n30795), .ZN(n27571) );
  OAI211_X1 U35624 ( .C1(n27570), .C2(n30792), .A(n30783), .B(n27571), .ZN(
        n27572) );
  OAI211_X1 U35625 ( .C1(n27574), .C2(n30795), .A(n27573), .B(n27572), .ZN(
        n27643) );
  NOR2_X2 U35626 ( .A1(n27644), .A2(n27643), .ZN(n32484) );
  OAI21_X1 U35627 ( .B1(n27686), .B2(n27685), .A(n27576), .ZN(n27691) );
  INV_X1 U35628 ( .A(n27685), .ZN(n27682) );
  OAI21_X1 U35629 ( .B1(n27579), .B2(n27682), .A(n27578), .ZN(n27586) );
  NAND2_X1 U35631 ( .A1(n27583), .A2(n27582), .ZN(n27585) );
  NAND3_X1 U35632 ( .A1(n27588), .A2(n30716), .A3(n2169), .ZN(n27589) );
  OAI211_X1 U35633 ( .C1(n28807), .C2(n30707), .A(n27590), .B(n27589), .ZN(
        n27591) );
  INV_X1 U35634 ( .A(n27591), .ZN(n27598) );
  INV_X1 U35635 ( .A(n27592), .ZN(n30713) );
  INV_X1 U35636 ( .A(n27593), .ZN(n27594) );
  NAND2_X1 U35637 ( .A1(n29850), .A2(n30725), .ZN(n27595) );
  NAND2_X1 U35638 ( .A1(n27601), .A2(n27600), .ZN(n30657) );
  OAI21_X1 U35639 ( .B1(n30677), .B2(n30673), .A(n30657), .ZN(n27603) );
  NAND2_X1 U35640 ( .A1(n27603), .A2(n27602), .ZN(n27613) );
  INV_X1 U35641 ( .A(n27608), .ZN(n30659) );
  OAI211_X1 U35642 ( .C1(n23859), .C2(n27604), .A(n30664), .B(n30659), .ZN(
        n27606) );
  INV_X1 U35643 ( .A(n27605), .ZN(n30672) );
  NAND2_X1 U35644 ( .A1(n27607), .A2(n30661), .ZN(n27612) );
  OAI211_X1 U35645 ( .C1(n32483), .C2(n32484), .A(n32472), .B(n32016), .ZN(
        n27646) );
  NAND2_X1 U35646 ( .A1(n27720), .A2(n27627), .ZN(n27614) );
  NAND3_X1 U35647 ( .A1(n27614), .A2(n27732), .A3(n27623), .ZN(n27617) );
  NAND3_X1 U35648 ( .A1(n27615), .A2(n27618), .A3(n27730), .ZN(n27616) );
  MUX2_X1 U35649 ( .A(n27619), .B(n27736), .S(n27618), .Z(n27620) );
  NAND3_X1 U35650 ( .A1(n27621), .A2(n27635), .A3(n27735), .ZN(n27626) );
  NAND4_X1 U35651 ( .A1(n27730), .A2(n27638), .A3(n22344), .A4(n27623), .ZN(
        n27625) );
  NAND2_X1 U35652 ( .A1(n27719), .A2(n27623), .ZN(n27624) );
  INV_X1 U35653 ( .A(n27627), .ZN(n27631) );
  OAI21_X1 U35655 ( .B1(n27732), .B2(n597), .A(n27632), .ZN(n27634) );
  OAI21_X1 U35656 ( .B1(n27639), .B2(n27635), .A(n27634), .ZN(n27642) );
  INV_X1 U35657 ( .A(n27636), .ZN(n27637) );
  NAND3_X1 U35658 ( .A1(n27639), .A2(n27638), .A3(n27637), .ZN(n27640) );
  XNOR2_X1 U35659 ( .A(n32027), .B(n32485), .ZN(n27645) );
  NOR2_X1 U35660 ( .A1(n27646), .A2(n27645), .ZN(n27651) );
  NAND2_X1 U35661 ( .A1(n32489), .A2(n32478), .ZN(n29626) );
  OAI211_X1 U35662 ( .C1(n29625), .C2(n32491), .A(n27647), .B(n3664), .ZN(
        n27648) );
  OAI21_X1 U35663 ( .B1(n32487), .B2(n32015), .A(n27648), .ZN(n27649) );
  NAND2_X1 U35664 ( .A1(n27649), .A2(n32484), .ZN(n27650) );
  AOI21_X1 U35665 ( .B1(n27662), .B2(n2642), .A(n27652), .ZN(n27655) );
  INV_X1 U35666 ( .A(n27659), .ZN(n27676) );
  NAND2_X1 U35667 ( .A1(n27660), .A2(n2642), .ZN(n27667) );
  OAI21_X1 U35668 ( .B1(n2642), .B2(n27662), .A(n27661), .ZN(n27664) );
  NAND2_X1 U35669 ( .A1(n27664), .A2(n51117), .ZN(n27666) );
  MUX2_X1 U35670 ( .A(n27667), .B(n27666), .S(n27665), .Z(n27675) );
  NAND2_X1 U35671 ( .A1(n27673), .A2(n27672), .ZN(n27674) );
  OAI21_X1 U35672 ( .B1(n27682), .B2(n27681), .A(n27680), .ZN(n27684) );
  INV_X1 U35673 ( .A(n27687), .ZN(n27689) );
  NAND2_X1 U35674 ( .A1(n27689), .A2(n27688), .ZN(n27692) );
  MUX2_X1 U35675 ( .A(n27692), .B(n27691), .S(n27690), .Z(n27693) );
  OAI211_X1 U35676 ( .C1(n27695), .C2(n29545), .A(n27694), .B(n29563), .ZN(
        n27696) );
  NAND2_X1 U35677 ( .A1(n29563), .A2(n29549), .ZN(n27698) );
  NOR2_X1 U35678 ( .A1(n27698), .A2(n27697), .ZN(n27699) );
  NAND2_X1 U35679 ( .A1(n29550), .A2(n6339), .ZN(n27704) );
  OAI211_X1 U35680 ( .C1(n29563), .C2(n29545), .A(n29551), .B(n27704), .ZN(
        n27705) );
  NAND2_X1 U35681 ( .A1(n30601), .A2(n29686), .ZN(n27775) );
  OR2_X1 U35682 ( .A1(n31096), .A2(n27775), .ZN(n30918) );
  NAND3_X1 U35683 ( .A1(n27707), .A2(n27706), .A3(n26731), .ZN(n27713) );
  AOI21_X1 U35684 ( .B1(n51678), .B2(n29424), .A(n29413), .ZN(n27708) );
  OAI211_X1 U35685 ( .C1(n27711), .C2(n27710), .A(n2115), .B(n27708), .ZN(
        n27712) );
  NAND2_X1 U35686 ( .A1(n27713), .A2(n27712), .ZN(n27718) );
  NAND2_X1 U35687 ( .A1(n30597), .A2(n30912), .ZN(n31090) );
  INV_X1 U35688 ( .A(n27719), .ZN(n27737) );
  OAI211_X1 U35689 ( .C1(n27724), .C2(n27737), .A(n27723), .B(n27722), .ZN(
        n27725) );
  AND2_X1 U35690 ( .A1(n27726), .A2(n27727), .ZN(n27741) );
  NAND3_X1 U35691 ( .A1(n27730), .A2(n2144), .A3(n27728), .ZN(n27731) );
  OAI21_X1 U35692 ( .B1(n27733), .B2(n27732), .A(n27731), .ZN(n27734) );
  NAND2_X1 U35693 ( .A1(n27734), .A2(n737), .ZN(n27740) );
  OAI21_X1 U35694 ( .B1(n27737), .B2(n27736), .A(n27735), .ZN(n27738) );
  OR2_X1 U35695 ( .A1(n27760), .A2(n27764), .ZN(n29465) );
  INV_X1 U35696 ( .A(n27744), .ZN(n27745) );
  INV_X1 U35697 ( .A(n27746), .ZN(n27747) );
  NOR2_X1 U35698 ( .A1(n27748), .A2(n27747), .ZN(n27770) );
  INV_X1 U35699 ( .A(n27749), .ZN(n27753) );
  NAND3_X1 U35700 ( .A1(n27751), .A2(n27760), .A3(n27015), .ZN(n27752) );
  NAND2_X1 U35701 ( .A1(n27753), .A2(n27752), .ZN(n27754) );
  NAND2_X1 U35702 ( .A1(n29461), .A2(n29469), .ZN(n27756) );
  MUX2_X1 U35703 ( .A(n27757), .B(n27756), .S(n27015), .Z(n27768) );
  NOR2_X1 U35704 ( .A1(n27759), .A2(n27758), .ZN(n27761) );
  OAI21_X1 U35705 ( .B1(n27762), .B2(n27761), .A(n27760), .ZN(n27763) );
  OAI21_X1 U35706 ( .B1(n29460), .B2(n29455), .A(n27763), .ZN(n27767) );
  NOR2_X1 U35707 ( .A1(n27765), .A2(n27764), .ZN(n27766) );
  AOI211_X1 U35708 ( .C1(n30918), .C2(n31090), .A(n30592), .B(n30607), .ZN(
        n27773) );
  NAND3_X1 U35709 ( .A1(n30592), .A2(n30912), .A3(n29686), .ZN(n30594) );
  OAI21_X1 U35710 ( .B1(n30918), .B2(n30602), .A(n30594), .ZN(n27772) );
  NOR2_X1 U35711 ( .A1(n27773), .A2(n27772), .ZN(n27779) );
  OAI21_X1 U35712 ( .B1(n30911), .B2(n30607), .A(n30590), .ZN(n27774) );
  NAND2_X1 U35713 ( .A1(n30916), .A2(n27774), .ZN(n27776) );
  NOR2_X1 U35714 ( .A1(n30593), .A2(n30601), .ZN(n31091) );
  NAND2_X1 U35715 ( .A1(n31091), .A2(n30602), .ZN(n29683) );
  NAND4_X1 U35716 ( .A1(n30598), .A2(n30607), .A3(n31096), .A4(n30601), .ZN(
        n27777) );
  XNOR2_X1 U35717 ( .A(n34128), .B(n37040), .ZN(n28478) );
  INV_X1 U35718 ( .A(n27780), .ZN(n27932) );
  OAI22_X1 U35719 ( .A1(n29186), .A2(n27780), .B1(n29191), .B2(n27783), .ZN(
        n27781) );
  OAI21_X1 U35720 ( .B1(n27782), .B2(n27932), .A(n27781), .ZN(n29277) );
  NAND2_X1 U35721 ( .A1(n51116), .A2(n27783), .ZN(n29184) );
  OAI211_X1 U35722 ( .C1(n28713), .C2(n25479), .A(n29191), .B(n29184), .ZN(
        n27784) );
  NAND2_X1 U35723 ( .A1(n28710), .A2(n29272), .ZN(n27788) );
  NAND2_X1 U35724 ( .A1(n28713), .A2(n29190), .ZN(n27786) );
  NAND2_X1 U35726 ( .A1(n27787), .A2(n29188), .ZN(n27793) );
  INV_X1 U35727 ( .A(n27788), .ZN(n27789) );
  NAND2_X1 U35728 ( .A1(n27789), .A2(n29270), .ZN(n27792) );
  NAND3_X1 U35729 ( .A1(n29188), .A2(n27930), .A3(n28711), .ZN(n27791) );
  NAND2_X1 U35730 ( .A1(n29186), .A2(n28713), .ZN(n27790) );
  AND4_X1 U35731 ( .A1(n27793), .A2(n27792), .A3(n27791), .A4(n27790), .ZN(
        n27794) );
  AOI21_X1 U35732 ( .B1(n29532), .B2(n398), .A(n29525), .ZN(n27799) );
  INV_X1 U35733 ( .A(n29534), .ZN(n27798) );
  AOI22_X1 U35734 ( .A1(n29509), .A2(n28623), .B1(n27799), .B2(n27798), .ZN(
        n27803) );
  NAND3_X1 U35735 ( .A1(n27800), .A2(n28618), .A3(n5183), .ZN(n27802) );
  NAND2_X1 U35736 ( .A1(n28628), .A2(n29532), .ZN(n27801) );
  NAND4_X2 U35737 ( .A1(n27803), .A2(n27804), .A3(n27802), .A4(n27801), .ZN(
        n31891) );
  NAND2_X1 U35738 ( .A1(n31418), .A2(n31891), .ZN(n29657) );
  INV_X1 U35739 ( .A(n27896), .ZN(n28637) );
  INV_X1 U35740 ( .A(n29314), .ZN(n28636) );
  OAI21_X1 U35742 ( .B1(n51793), .B2(n51107), .A(n29325), .ZN(n27806) );
  NAND2_X1 U35743 ( .A1(n27808), .A2(n27807), .ZN(n27889) );
  OAI21_X1 U35744 ( .B1(n29331), .B2(n52216), .A(n29319), .ZN(n27810) );
  NAND3_X1 U35745 ( .A1(n27889), .A2(n27810), .A3(n27809), .ZN(n27816) );
  NAND2_X1 U35746 ( .A1(n29324), .A2(n52217), .ZN(n27812) );
  NOR2_X1 U35747 ( .A1(n459), .A2(n29330), .ZN(n27811) );
  NAND4_X1 U35748 ( .A1(n27812), .A2(n29315), .A3(n29326), .A4(n27811), .ZN(
        n27815) );
  NAND3_X1 U35749 ( .A1(n27818), .A2(n29323), .A3(n52216), .ZN(n27814) );
  NAND2_X1 U35750 ( .A1(n27819), .A2(n27897), .ZN(n27824) );
  NAND2_X1 U35751 ( .A1(n29657), .A2(n31425), .ZN(n31423) );
  NAND2_X1 U35752 ( .A1(n27828), .A2(n27827), .ZN(n27832) );
  OAI21_X1 U35753 ( .B1(n27830), .B2(n27829), .A(n26722), .ZN(n27831) );
  NAND2_X1 U35754 ( .A1(n27835), .A2(n29441), .ZN(n27833) );
  INV_X1 U35755 ( .A(n27836), .ZN(n27838) );
  NOR2_X1 U35756 ( .A1(n27840), .A2(n29444), .ZN(n27841) );
  NOR2_X1 U35757 ( .A1(n27844), .A2(n29289), .ZN(n27846) );
  XNOR2_X1 U35758 ( .A(n26077), .B(n29291), .ZN(n27845) );
  INV_X1 U35759 ( .A(n28701), .ZN(n28683) );
  AOI22_X1 U35760 ( .A1(n27846), .A2(n29306), .B1(n27845), .B2(n28683), .ZN(
        n27851) );
  OR2_X1 U35761 ( .A1(n51518), .A2(n29294), .ZN(n29299) );
  OAI22_X1 U35762 ( .A1(n28684), .A2(n29299), .B1(n29305), .B2(n28695), .ZN(
        n27848) );
  NAND2_X1 U35763 ( .A1(n28701), .A2(n51518), .ZN(n27849) );
  NOR2_X1 U35764 ( .A1(n28688), .A2(n29294), .ZN(n28696) );
  AOI22_X1 U35765 ( .A1(n27849), .A2(n29309), .B1(n28696), .B2(n28700), .ZN(
        n27850) );
  AOI21_X1 U35766 ( .B1(n31423), .B2(n31420), .A(n31422), .ZN(n27874) );
  NOR2_X1 U35767 ( .A1(n31418), .A2(n31891), .ZN(n29991) );
  NAND2_X1 U35768 ( .A1(n29478), .A2(n6080), .ZN(n27853) );
  NAND4_X1 U35769 ( .A1(n28669), .A2(n27860), .A3(n28666), .A4(n27852), .ZN(
        n28676) );
  OAI21_X1 U35770 ( .B1(n27854), .B2(n27853), .A(n28676), .ZN(n27855) );
  INV_X1 U35771 ( .A(n27859), .ZN(n28667) );
  NAND2_X1 U35772 ( .A1(n28669), .A2(n51110), .ZN(n29485) );
  INV_X1 U35773 ( .A(n29479), .ZN(n29487) );
  NAND3_X1 U35774 ( .A1(n28671), .A2(n29494), .A3(n27856), .ZN(n27857) );
  INV_X1 U35775 ( .A(n28671), .ZN(n27861) );
  OAI211_X1 U35776 ( .C1(n29496), .C2(n27861), .A(n28672), .B(n3124), .ZN(
        n27865) );
  NAND2_X1 U35777 ( .A1(n29480), .A2(n28669), .ZN(n27862) );
  AND2_X1 U35778 ( .A1(n27863), .A2(n27862), .ZN(n27864) );
  NAND2_X1 U35779 ( .A1(n31892), .A2(n31425), .ZN(n31410) );
  AND2_X1 U35780 ( .A1(n31410), .A2(n31418), .ZN(n27870) );
  NAND2_X1 U35781 ( .A1(n31418), .A2(n31899), .ZN(n31893) );
  NAND2_X1 U35782 ( .A1(n31893), .A2(n29657), .ZN(n29990) );
  NAND2_X1 U35783 ( .A1(n31146), .A2(n31891), .ZN(n31141) );
  AOI21_X1 U35784 ( .B1(n31899), .B2(n31141), .A(n620), .ZN(n27872) );
  OR2_X1 U35785 ( .A1(n31891), .A2(n31422), .ZN(n31412) );
  OR2_X1 U35786 ( .A1(n31144), .A2(n31899), .ZN(n31137) );
  OAI21_X1 U35787 ( .B1(n31412), .B2(n31425), .A(n31137), .ZN(n27871) );
  NAND2_X1 U35788 ( .A1(n31892), .A2(n31891), .ZN(n29985) );
  OAI211_X1 U35789 ( .C1(n27872), .C2(n27871), .A(n725), .B(n29985), .ZN(
        n27873) );
  INV_X1 U35790 ( .A(n29344), .ZN(n29351) );
  NAND2_X1 U35791 ( .A1(n29202), .A2(n29351), .ZN(n27879) );
  INV_X1 U35792 ( .A(n30194), .ZN(n27875) );
  AOI21_X1 U35793 ( .B1(n27876), .B2(n27886), .A(n51109), .ZN(n27877) );
  NAND2_X1 U35794 ( .A1(n30197), .A2(n30200), .ZN(n27880) );
  MUX2_X1 U35795 ( .A(n29350), .B(n27880), .S(n30191), .Z(n27905) );
  NAND2_X1 U35796 ( .A1(n27903), .A2(n27905), .ZN(n30619) );
  XNOR2_X1 U35797 ( .A(n27882), .B(n30210), .ZN(n27883) );
  NAND2_X1 U35798 ( .A1(n30211), .A2(n29345), .ZN(n29205) );
  INV_X1 U35799 ( .A(n29204), .ZN(n30199) );
  NAND3_X1 U35800 ( .A1(n27885), .A2(n30209), .A3(n30199), .ZN(n27912) );
  NAND3_X1 U35801 ( .A1(n27888), .A2(n30210), .A3(n29200), .ZN(n27906) );
  NAND2_X1 U35802 ( .A1(n27886), .A2(n30202), .ZN(n27909) );
  NOR2_X1 U35803 ( .A1(n51793), .A2(n459), .ZN(n27891) );
  OAI21_X1 U35804 ( .B1(n29320), .B2(n27891), .A(n27890), .ZN(n27892) );
  INV_X1 U35805 ( .A(n27892), .ZN(n27893) );
  INV_X1 U35806 ( .A(n29317), .ZN(n27895) );
  OR3_X1 U35807 ( .A1(n27896), .A2(n29314), .A3(n27895), .ZN(n27900) );
  NAND2_X1 U35808 ( .A1(n27897), .A2(n29332), .ZN(n27898) );
  NAND4_X1 U35809 ( .A1(n27901), .A2(n27900), .A3(n27899), .A4(n27898), .ZN(
        n27902) );
  OR2_X1 U35810 ( .A1(n711), .A2(n32299), .ZN(n27979) );
  INV_X1 U35811 ( .A(n27903), .ZN(n27904) );
  NAND2_X1 U35812 ( .A1(n30622), .A2(n27904), .ZN(n27923) );
  INV_X1 U35813 ( .A(n27905), .ZN(n27908) );
  OR2_X1 U35814 ( .A1(n29227), .A2(n30263), .ZN(n27970) );
  OAI211_X1 U35815 ( .C1(n30268), .C2(n29240), .A(n27970), .B(n27906), .ZN(
        n27907) );
  NOR2_X1 U35816 ( .A1(n27908), .A2(n27907), .ZN(n27922) );
  INV_X1 U35818 ( .A(n27971), .ZN(n30270) );
  AND4_X1 U35820 ( .A1(n27912), .A2(n27911), .A3(n29340), .A4(n27969), .ZN(
        n27921) );
  NAND2_X1 U35821 ( .A1(n29242), .A2(n52147), .ZN(n29219) );
  INV_X1 U35822 ( .A(n27914), .ZN(n27915) );
  NAND2_X1 U35823 ( .A1(n29235), .A2(n27915), .ZN(n27916) );
  NAND2_X1 U35825 ( .A1(n27920), .A2(n27919), .ZN(n27972) );
  NAND2_X1 U35826 ( .A1(n28715), .A2(n29187), .ZN(n27926) );
  NAND2_X1 U35827 ( .A1(n27926), .A2(n27925), .ZN(n27928) );
  NAND2_X1 U35828 ( .A1(n28710), .A2(n5425), .ZN(n27927) );
  OAI211_X1 U35830 ( .C1(n29272), .C2(n29269), .A(n29283), .B(n27931), .ZN(
        n27934) );
  NAND2_X1 U35831 ( .A1(n51706), .A2(n27932), .ZN(n27933) );
  AOI21_X1 U35832 ( .B1(n27979), .B2(n32295), .A(n435), .ZN(n27984) );
  INV_X1 U35833 ( .A(n27936), .ZN(n30221) );
  NOR2_X1 U35834 ( .A1(n29247), .A2(n29263), .ZN(n27937) );
  NAND2_X1 U35835 ( .A1(n27939), .A2(n30230), .ZN(n27940) );
  NAND2_X1 U35836 ( .A1(n27940), .A2(n30234), .ZN(n27950) );
  INV_X1 U35837 ( .A(n28658), .ZN(n27941) );
  NAND2_X1 U35838 ( .A1(n30227), .A2(n27941), .ZN(n30225) );
  NAND4_X1 U35840 ( .A1(n29120), .A2(n28652), .A3(n29260), .A4(n51114), .ZN(
        n27942) );
  AND2_X1 U35841 ( .A1(n30225), .A2(n27942), .ZN(n27949) );
  INV_X1 U35842 ( .A(n29248), .ZN(n29126) );
  OAI21_X1 U35843 ( .B1(n29260), .B2(n28657), .A(n29126), .ZN(n27945) );
  NOR2_X1 U35844 ( .A1(n28650), .A2(n29263), .ZN(n27943) );
  OAI21_X1 U35845 ( .B1(n29249), .B2(n27943), .A(n29248), .ZN(n27944) );
  NAND2_X1 U35846 ( .A1(n27945), .A2(n27944), .ZN(n27948) );
  AND3_X1 U35847 ( .A1(n4724), .A2(n29123), .A3(n29247), .ZN(n28654) );
  MUX2_X1 U35848 ( .A(n28654), .B(n29119), .S(n30234), .Z(n27946) );
  NAND2_X1 U35849 ( .A1(n27946), .A2(n29251), .ZN(n27947) );
  NAND3_X1 U35850 ( .A1(n32295), .A2(n31740), .A3(n435), .ZN(n27968) );
  INV_X1 U35851 ( .A(n27951), .ZN(n27952) );
  NOR2_X1 U35852 ( .A1(n27953), .A2(n27952), .ZN(n29166) );
  NOR2_X1 U35853 ( .A1(n27953), .A2(n30251), .ZN(n27954) );
  NOR2_X1 U35854 ( .A1(n29166), .A2(n27954), .ZN(n27967) );
  OAI21_X1 U35855 ( .B1(n27955), .B2(n51473), .A(n29171), .ZN(n27966) );
  NAND3_X1 U35856 ( .A1(n29156), .A2(n29155), .A3(n52165), .ZN(n30243) );
  OAI21_X1 U35857 ( .B1(n27957), .B2(n27956), .A(n30243), .ZN(n27958) );
  NAND2_X1 U35858 ( .A1(n27958), .A2(n30249), .ZN(n27965) );
  INV_X1 U35859 ( .A(n27959), .ZN(n27963) );
  NOR2_X1 U35860 ( .A1(n27963), .A2(n27962), .ZN(n27964) );
  NAND2_X1 U35862 ( .A1(n27968), .A2(n31749), .ZN(n27983) );
  AND2_X1 U35865 ( .A1(n27971), .A2(n30268), .ZN(n27973) );
  NAND2_X1 U35866 ( .A1(n32299), .A2(n31746), .ZN(n30632) );
  NOR2_X1 U35867 ( .A1(n32299), .A2(n435), .ZN(n27975) );
  OAI211_X1 U35868 ( .C1(n711), .C2(n31746), .A(n32302), .B(n27975), .ZN(
        n27977) );
  NAND4_X1 U35869 ( .A1(n711), .A2(n4434), .A3(n31746), .A4(n31743), .ZN(
        n27976) );
  OAI211_X1 U35870 ( .C1(n31743), .C2(n30632), .A(n27977), .B(n27976), .ZN(
        n27978) );
  OAI21_X1 U35871 ( .B1(n27979), .B2(n435), .A(n30635), .ZN(n27981) );
  AOI21_X1 U35872 ( .B1(n4434), .B2(n31740), .A(n31749), .ZN(n27980) );
  NAND2_X1 U35873 ( .A1(n27981), .A2(n27980), .ZN(n27982) );
  NAND2_X1 U35874 ( .A1(n28907), .A2(n28578), .ZN(n27985) );
  AND2_X1 U35875 ( .A1(n27986), .A2(n27985), .ZN(n27989) );
  NAND2_X1 U35876 ( .A1(n27991), .A2(n27987), .ZN(n28586) );
  OAI211_X1 U35877 ( .C1(n27994), .C2(n27999), .A(n28586), .B(n28897), .ZN(
        n27988) );
  MUX2_X1 U35879 ( .A(n27989), .B(n27988), .S(n28896), .Z(n28006) );
  INV_X1 U35880 ( .A(n27990), .ZN(n27992) );
  NAND2_X1 U35881 ( .A1(n27992), .A2(n27991), .ZN(n28898) );
  NAND2_X1 U35882 ( .A1(n27993), .A2(n28000), .ZN(n28589) );
  INV_X1 U35883 ( .A(n27994), .ZN(n28583) );
  OAI211_X1 U35884 ( .C1(n27997), .C2(n28589), .A(n27996), .B(n27995), .ZN(
        n28004) );
  INV_X1 U35885 ( .A(n27998), .ZN(n28002) );
  NAND2_X1 U35886 ( .A1(n28582), .A2(n27999), .ZN(n28001) );
  AOI21_X1 U35887 ( .B1(n28002), .B2(n28001), .A(n28000), .ZN(n28003) );
  NOR2_X1 U35888 ( .A1(n28004), .A2(n28003), .ZN(n28005) );
  INV_X1 U35889 ( .A(n28926), .ZN(n29014) );
  NAND2_X1 U35890 ( .A1(n28916), .A2(n29014), .ZN(n29008) );
  INV_X1 U35891 ( .A(n28197), .ZN(n28012) );
  NAND2_X1 U35892 ( .A1(n28918), .A2(n28933), .ZN(n29016) );
  INV_X1 U35893 ( .A(n29018), .ZN(n28200) );
  INV_X1 U35894 ( .A(n28919), .ZN(n29020) );
  NOR2_X1 U35895 ( .A1(n28565), .A2(n28008), .ZN(n28011) );
  NAND2_X1 U35896 ( .A1(n28194), .A2(n29014), .ZN(n28009) );
  NAND4_X1 U35897 ( .A1(n28915), .A2(n29015), .A3(n29011), .A4(n28009), .ZN(
        n28010) );
  NAND3_X1 U35898 ( .A1(n28019), .A2(n28572), .A3(n28012), .ZN(n28013) );
  INV_X1 U35899 ( .A(n29008), .ZN(n28015) );
  NAND2_X1 U35900 ( .A1(n28197), .A2(n28923), .ZN(n28016) );
  AOI21_X1 U35901 ( .B1(n28016), .B2(n28200), .A(n29020), .ZN(n28017) );
  NAND2_X1 U35902 ( .A1(n28922), .A2(n28019), .ZN(n28569) );
  INV_X1 U35903 ( .A(n28569), .ZN(n28020) );
  INV_X1 U35904 ( .A(n30312), .ZN(n30165) );
  NAND2_X1 U35905 ( .A1(n30165), .A2(n28025), .ZN(n29133) );
  NAND2_X1 U35906 ( .A1(n28023), .A2(n28022), .ZN(n28024) );
  NAND2_X1 U35907 ( .A1(n28024), .A2(n547), .ZN(n28027) );
  NAND2_X1 U35908 ( .A1(n28025), .A2(n6084), .ZN(n28026) );
  NAND4_X1 U35909 ( .A1(n29133), .A2(n28028), .A3(n28027), .A4(n28026), .ZN(
        n28029) );
  AND2_X1 U35910 ( .A1(n30178), .A2(n30181), .ZN(n30164) );
  OAI21_X1 U35911 ( .B1(n28033), .B2(n30307), .A(n28032), .ZN(n28034) );
  XNOR2_X1 U35912 ( .A(n28036), .B(n28035), .ZN(n28044) );
  XNOR2_X1 U35913 ( .A(n44921), .B(n42619), .ZN(n28037) );
  XNOR2_X1 U35914 ( .A(n28038), .B(n28037), .ZN(n28039) );
  XNOR2_X1 U35915 ( .A(n51057), .B(n28039), .ZN(n28042) );
  XNOR2_X1 U35916 ( .A(n28042), .B(n28041), .ZN(n28043) );
  XNOR2_X1 U35917 ( .A(n28044), .B(n28043), .ZN(n28045) );
  XNOR2_X1 U35918 ( .A(n28046), .B(n28045), .ZN(n28082) );
  INV_X1 U35920 ( .A(n28047), .ZN(n28052) );
  XNOR2_X1 U35921 ( .A(n28049), .B(n28048), .ZN(n28051) );
  XNOR2_X1 U35922 ( .A(n28051), .B(n51666), .ZN(n28385) );
  XNOR2_X1 U35923 ( .A(n28052), .B(n28385), .ZN(n28053) );
  XNOR2_X1 U35924 ( .A(n28054), .B(n28053), .ZN(n28066) );
  XNOR2_X1 U35925 ( .A(n4638), .B(n4213), .ZN(n28057) );
  XNOR2_X1 U35926 ( .A(n28058), .B(n28057), .ZN(n42591) );
  XNOR2_X1 U35927 ( .A(n34601), .B(n42591), .ZN(n28059) );
  XNOR2_X1 U35928 ( .A(n28060), .B(n28059), .ZN(n28061) );
  XNOR2_X1 U35929 ( .A(n28061), .B(n28381), .ZN(n28062) );
  XNOR2_X1 U35930 ( .A(n28064), .B(n28063), .ZN(n28065) );
  XNOR2_X1 U35931 ( .A(n28066), .B(n28065), .ZN(n28965) );
  NAND2_X1 U35932 ( .A1(n29797), .A2(n28965), .ZN(n28957) );
  XNOR2_X1 U35933 ( .A(n28069), .B(n51749), .ZN(n28078) );
  XNOR2_X1 U35934 ( .A(n28070), .B(n47268), .ZN(n28072) );
  XNOR2_X1 U35935 ( .A(n28072), .B(n28071), .ZN(n28073) );
  XNOR2_X1 U35936 ( .A(n33119), .B(n28073), .ZN(n43512) );
  XNOR2_X1 U35937 ( .A(n45736), .B(n4838), .ZN(n28074) );
  XNOR2_X1 U35938 ( .A(n36854), .B(n28074), .ZN(n28075) );
  XNOR2_X1 U35939 ( .A(n35590), .B(n28075), .ZN(n44172) );
  XNOR2_X1 U35940 ( .A(n43512), .B(n44172), .ZN(n28076) );
  XNOR2_X1 U35941 ( .A(n28078), .B(n28077), .ZN(n28079) );
  INV_X1 U35942 ( .A(n28082), .ZN(n28497) );
  XNOR2_X1 U35943 ( .A(n28085), .B(n28084), .ZN(n28086) );
  XNOR2_X1 U35944 ( .A(n28087), .B(n28086), .ZN(n28088) );
  XNOR2_X1 U35945 ( .A(n28089), .B(n28088), .ZN(n43096) );
  XNOR2_X1 U35946 ( .A(n42889), .B(n28090), .ZN(n41885) );
  XNOR2_X1 U35947 ( .A(n43096), .B(n41885), .ZN(n28091) );
  XNOR2_X1 U35948 ( .A(n28220), .B(n28091), .ZN(n28092) );
  XNOR2_X1 U35949 ( .A(n28093), .B(n28092), .ZN(n28094) );
  INV_X1 U35950 ( .A(n28096), .ZN(n28097) );
  XNOR2_X1 U35951 ( .A(n28097), .B(n28098), .ZN(n28099) );
  NAND2_X1 U35952 ( .A1(n28497), .A2(n28867), .ZN(n28134) );
  XNOR2_X1 U35953 ( .A(n28101), .B(n28100), .ZN(n28112) );
  XNOR2_X1 U35954 ( .A(n37082), .B(n34575), .ZN(n44907) );
  XNOR2_X1 U35955 ( .A(n42657), .B(n44907), .ZN(n28102) );
  XNOR2_X1 U35956 ( .A(n28103), .B(n28102), .ZN(n28105) );
  XNOR2_X1 U35957 ( .A(n28105), .B(n28104), .ZN(n28108) );
  XNOR2_X1 U35958 ( .A(n28311), .B(n28106), .ZN(n28432) );
  XNOR2_X1 U35959 ( .A(n28110), .B(n28109), .ZN(n28111) );
  INV_X1 U35960 ( .A(n28113), .ZN(n28114) );
  XNOR2_X1 U35961 ( .A(n28116), .B(n28115), .ZN(n44234) );
  XNOR2_X1 U35962 ( .A(n44234), .B(n43563), .ZN(n28117) );
  XNOR2_X1 U35963 ( .A(n28396), .B(n28117), .ZN(n28118) );
  XNOR2_X1 U35964 ( .A(n28118), .B(n28291), .ZN(n28120) );
  XNOR2_X1 U35965 ( .A(n28120), .B(n28119), .ZN(n28122) );
  XNOR2_X1 U35966 ( .A(n28122), .B(n28121), .ZN(n28124) );
  XNOR2_X1 U35967 ( .A(n28124), .B(n28123), .ZN(n28133) );
  INV_X1 U35968 ( .A(n45403), .ZN(n28125) );
  XNOR2_X1 U35969 ( .A(n28126), .B(n28125), .ZN(n28128) );
  XNOR2_X1 U35970 ( .A(n28128), .B(n51121), .ZN(n28130) );
  XNOR2_X1 U35971 ( .A(n28130), .B(n28129), .ZN(n28404) );
  XNOR2_X1 U35972 ( .A(n28131), .B(n28404), .ZN(n28132) );
  AOI21_X1 U35973 ( .B1(n28507), .B2(n28134), .A(n28505), .ZN(n28137) );
  OAI21_X1 U35975 ( .B1(n29796), .B2(n5054), .A(n28508), .ZN(n28136) );
  INV_X1 U35976 ( .A(n28965), .ZN(n28138) );
  NAND3_X1 U35977 ( .A1(n28958), .A2(n5056), .A3(n28950), .ZN(n28135) );
  NAND2_X1 U35978 ( .A1(n29797), .A2(n28138), .ZN(n29794) );
  NAND2_X1 U35979 ( .A1(n28860), .A2(n28862), .ZN(n28139) );
  INV_X1 U35980 ( .A(n29796), .ZN(n29803) );
  NAND3_X1 U35981 ( .A1(n28952), .A2(n28962), .A3(n5057), .ZN(n29792) );
  INV_X1 U35982 ( .A(n28139), .ZN(n28140) );
  NAND3_X1 U35983 ( .A1(n28140), .A2(n28957), .A3(n5056), .ZN(n28141) );
  AND2_X1 U35984 ( .A1(n28963), .A2(n28141), .ZN(n28142) );
  OAI21_X1 U35986 ( .B1(n28148), .B2(n30282), .A(n28147), .ZN(n28149) );
  NAND2_X1 U35987 ( .A1(n28545), .A2(n28149), .ZN(n28150) );
  INV_X1 U35989 ( .A(n32590), .ZN(n32977) );
  AND2_X1 U35990 ( .A1(n32977), .A2(n32595), .ZN(n28166) );
  NAND2_X1 U35991 ( .A1(n28874), .A2(n28155), .ZN(n28533) );
  NAND2_X1 U35992 ( .A1(n28881), .A2(n28533), .ZN(n28156) );
  MUX2_X1 U35993 ( .A(n28881), .B(n28156), .S(n28883), .Z(n28157) );
  AND2_X1 U35994 ( .A1(n28875), .A2(n29035), .ZN(n28158) );
  OAI21_X1 U35995 ( .B1(n29047), .B2(n28159), .A(n28883), .ZN(n28162) );
  NAND3_X1 U35996 ( .A1(n29034), .A2(n28880), .A3(n28160), .ZN(n28161) );
  AND2_X1 U35997 ( .A1(n32600), .A2(n32595), .ZN(n28163) );
  AOI22_X1 U35998 ( .A1(n28166), .A2(n28164), .B1(n28163), .B2(n32988), .ZN(
        n28169) );
  NOR2_X1 U35999 ( .A1(n32595), .A2(n32990), .ZN(n28165) );
  NAND3_X1 U36001 ( .A1(n28607), .A2(n28165), .A3(n28608), .ZN(n28168) );
  NAND3_X1 U36002 ( .A1(n32601), .A2(n28166), .A3(n32600), .ZN(n28167) );
  NAND4_X1 U36003 ( .A1(n28170), .A2(n28169), .A3(n28168), .A4(n28167), .ZN(
        n28174) );
  OAI211_X1 U36004 ( .C1(n29622), .C2(n32974), .A(n28171), .B(n52046), .ZN(
        n28172) );
  OAI21_X1 U36005 ( .B1(n28607), .B2(n32987), .A(n28172), .ZN(n28173) );
  NAND2_X1 U36007 ( .A1(n28189), .A2(n28970), .ZN(n30403) );
  MUX2_X1 U36008 ( .A(n30403), .B(n28982), .S(n29719), .Z(n28176) );
  NAND2_X1 U36009 ( .A1(n28176), .A2(n28175), .ZN(n28186) );
  NAND2_X1 U36010 ( .A1(n30411), .A2(n28974), .ZN(n28792) );
  NOR2_X1 U36011 ( .A1(n28792), .A2(n29724), .ZN(n28181) );
  AOI21_X1 U36012 ( .B1(n28178), .B2(n30407), .A(n30419), .ZN(n28180) );
  OAI21_X1 U36013 ( .B1(n28181), .B2(n28180), .A(n28179), .ZN(n28185) );
  INV_X1 U36014 ( .A(n28182), .ZN(n28184) );
  INV_X1 U36015 ( .A(n29715), .ZN(n28791) );
  NAND2_X1 U36016 ( .A1(n27281), .A2(n28187), .ZN(n28797) );
  INV_X1 U36017 ( .A(n28982), .ZN(n29716) );
  OAI22_X1 U36018 ( .A1(n28970), .A2(n28797), .B1(n30412), .B2(n29716), .ZN(
        n28188) );
  NOR2_X1 U36019 ( .A1(n29719), .A2(n29724), .ZN(n30413) );
  INV_X1 U36020 ( .A(n29721), .ZN(n30421) );
  OAI21_X1 U36021 ( .B1(n28188), .B2(n30413), .A(n30421), .ZN(n28192) );
  NAND3_X1 U36022 ( .A1(n28190), .A2(n30407), .A3(n30411), .ZN(n28191) );
  NOR2_X1 U36023 ( .A1(n51115), .A2(n28923), .ZN(n28195) );
  NAND2_X1 U36024 ( .A1(n28918), .A2(n29007), .ZN(n28932) );
  OAI22_X1 U36025 ( .A1(n28195), .A2(n28194), .B1(n28932), .B2(n28916), .ZN(
        n28198) );
  NAND2_X1 U36028 ( .A1(n28201), .A2(n28915), .ZN(n28205) );
  NOR2_X1 U36029 ( .A1(n29015), .A2(n28926), .ZN(n28202) );
  NAND2_X1 U36030 ( .A1(n28203), .A2(n28202), .ZN(n28204) );
  NAND4_X1 U36031 ( .A1(n28208), .A2(n28937), .A3(n28207), .A4(n28206), .ZN(
        n28209) );
  XNOR2_X1 U36032 ( .A(n32497), .B(n28211), .ZN(n46086) );
  XNOR2_X1 U36033 ( .A(n4628), .B(n4471), .ZN(n44386) );
  XNOR2_X1 U36034 ( .A(n46086), .B(n44386), .ZN(n28212) );
  XNOR2_X1 U36035 ( .A(n28213), .B(n28212), .ZN(n28215) );
  XNOR2_X1 U36036 ( .A(n28219), .B(n28218), .ZN(n28229) );
  XNOR2_X1 U36037 ( .A(n28220), .B(n39976), .ZN(n28222) );
  XNOR2_X1 U36038 ( .A(n28221), .B(n28222), .ZN(n28225) );
  INV_X1 U36039 ( .A(n28223), .ZN(n28224) );
  XNOR2_X1 U36040 ( .A(n28224), .B(n28225), .ZN(n28228) );
  INV_X1 U36041 ( .A(n28226), .ZN(n28227) );
  XNOR2_X1 U36043 ( .A(n28231), .B(n28230), .ZN(n28244) );
  XNOR2_X1 U36044 ( .A(n28233), .B(n28232), .ZN(n28235) );
  XNOR2_X1 U36045 ( .A(n28235), .B(n28234), .ZN(n43941) );
  XNOR2_X1 U36046 ( .A(n45350), .B(n34709), .ZN(n28236) );
  XNOR2_X1 U36047 ( .A(n43941), .B(n28236), .ZN(n28237) );
  XNOR2_X1 U36048 ( .A(n28238), .B(n28237), .ZN(n28239) );
  XNOR2_X1 U36049 ( .A(n28240), .B(n28239), .ZN(n28241) );
  XNOR2_X1 U36050 ( .A(n28242), .B(n28241), .ZN(n28243) );
  XNOR2_X1 U36051 ( .A(n28243), .B(n28244), .ZN(n28245) );
  INV_X1 U36052 ( .A(n29764), .ZN(n29054) );
  XNOR2_X1 U36053 ( .A(n28250), .B(n28249), .ZN(n28261) );
  XNOR2_X1 U36054 ( .A(n42240), .B(n35107), .ZN(n42367) );
  XNOR2_X1 U36055 ( .A(n28251), .B(n42367), .ZN(n28255) );
  XNOR2_X1 U36056 ( .A(n28252), .B(n45107), .ZN(n28253) );
  XNOR2_X1 U36057 ( .A(n28253), .B(n45104), .ZN(n28254) );
  XNOR2_X1 U36058 ( .A(n28255), .B(n28254), .ZN(n28256) );
  XNOR2_X1 U36059 ( .A(n28257), .B(n28256), .ZN(n28259) );
  XNOR2_X1 U36060 ( .A(n28261), .B(n28260), .ZN(n28262) );
  XNOR2_X1 U36061 ( .A(n28265), .B(n28264), .ZN(n28278) );
  INV_X1 U36062 ( .A(n28266), .ZN(n28268) );
  XNOR2_X1 U36063 ( .A(n28268), .B(n28267), .ZN(n42833) );
  XNOR2_X1 U36064 ( .A(n41567), .B(n4752), .ZN(n28269) );
  XNOR2_X1 U36065 ( .A(n42833), .B(n28269), .ZN(n28272) );
  XNOR2_X1 U36066 ( .A(n28271), .B(n28270), .ZN(n41225) );
  XNOR2_X1 U36067 ( .A(n28272), .B(n41225), .ZN(n28273) );
  XNOR2_X1 U36068 ( .A(n28274), .B(n28273), .ZN(n28275) );
  XNOR2_X1 U36069 ( .A(n28276), .B(n28275), .ZN(n28277) );
  XNOR2_X1 U36070 ( .A(n28278), .B(n28277), .ZN(n28282) );
  INV_X1 U36071 ( .A(n28279), .ZN(n28281) );
  INV_X1 U36072 ( .A(n28283), .ZN(n28285) );
  XNOR2_X1 U36073 ( .A(n28285), .B(n28284), .ZN(n45271) );
  XNOR2_X1 U36074 ( .A(n35816), .B(n36718), .ZN(n43852) );
  XNOR2_X1 U36075 ( .A(n43852), .B(n4837), .ZN(n43951) );
  XNOR2_X1 U36076 ( .A(n45271), .B(n43951), .ZN(n28286) );
  XNOR2_X1 U36077 ( .A(n28396), .B(n28286), .ZN(n28290) );
  XNOR2_X1 U36078 ( .A(n28288), .B(n28287), .ZN(n28289) );
  XNOR2_X1 U36079 ( .A(n28290), .B(n28289), .ZN(n28294) );
  XNOR2_X1 U36080 ( .A(n28291), .B(n28292), .ZN(n28293) );
  XNOR2_X1 U36081 ( .A(n369), .B(n28302), .ZN(n28315) );
  XNOR2_X1 U36082 ( .A(n28303), .B(n36698), .ZN(n28306) );
  XNOR2_X1 U36083 ( .A(n28304), .B(n49323), .ZN(n28305) );
  XNOR2_X1 U36084 ( .A(n28306), .B(n28305), .ZN(n42861) );
  XNOR2_X1 U36085 ( .A(n28307), .B(n4650), .ZN(n28308) );
  XNOR2_X1 U36086 ( .A(n28309), .B(n28308), .ZN(n41299) );
  XNOR2_X1 U36087 ( .A(n42861), .B(n41299), .ZN(n28310) );
  XNOR2_X1 U36088 ( .A(n28311), .B(n28310), .ZN(n28313) );
  XNOR2_X1 U36089 ( .A(n28313), .B(n749), .ZN(n28314) );
  XNOR2_X1 U36090 ( .A(n28315), .B(n28314), .ZN(n28316) );
  XNOR2_X1 U36091 ( .A(n28317), .B(n28316), .ZN(n28321) );
  XNOR2_X1 U36092 ( .A(n28318), .B(n28319), .ZN(n28320) );
  NAND3_X1 U36093 ( .A1(n514), .A2(n5389), .A3(n745), .ZN(n28853) );
  NAND2_X1 U36094 ( .A1(n28787), .A2(n28853), .ZN(n28322) );
  NAND2_X1 U36095 ( .A1(n28322), .A2(n29764), .ZN(n28327) );
  OAI21_X1 U36096 ( .B1(n30348), .B2(n29764), .A(n29754), .ZN(n28324) );
  INV_X1 U36097 ( .A(n30351), .ZN(n29763) );
  NOR2_X1 U36098 ( .A1(n29062), .A2(n28849), .ZN(n28323) );
  NOR2_X1 U36099 ( .A1(n30351), .A2(n514), .ZN(n28325) );
  AND2_X1 U36100 ( .A1(n51490), .A2(n514), .ZN(n29066) );
  AOI21_X1 U36101 ( .B1(n29063), .B2(n28325), .A(n29066), .ZN(n28326) );
  NAND2_X1 U36102 ( .A1(n29692), .A2(n29703), .ZN(n29866) );
  INV_X1 U36103 ( .A(n29869), .ZN(n28328) );
  INV_X1 U36104 ( .A(n30436), .ZN(n28332) );
  NAND2_X1 U36105 ( .A1(n28329), .A2(n28328), .ZN(n28330) );
  NAND4_X1 U36106 ( .A1(n28337), .A2(n28336), .A3(n28335), .A4(n28334), .ZN(
        n28339) );
  OAI211_X1 U36107 ( .C1(n29869), .C2(n28745), .A(n29859), .B(n29698), .ZN(
        n28338) );
  NAND2_X1 U36108 ( .A1(n32175), .A2(n32960), .ZN(n32172) );
  XNOR2_X1 U36109 ( .A(n28340), .B(n40107), .ZN(n28342) );
  XNOR2_X1 U36110 ( .A(n28342), .B(n28341), .ZN(n28345) );
  XNOR2_X1 U36111 ( .A(n28345), .B(n28344), .ZN(n28346) );
  XNOR2_X1 U36112 ( .A(n28347), .B(n28346), .ZN(n28349) );
  XNOR2_X1 U36113 ( .A(n34818), .B(n34711), .ZN(n45465) );
  XNOR2_X1 U36114 ( .A(n41367), .B(n4824), .ZN(n43820) );
  XNOR2_X1 U36115 ( .A(n43820), .B(n43739), .ZN(n28350) );
  XNOR2_X1 U36116 ( .A(n45465), .B(n28350), .ZN(n28351) );
  XNOR2_X1 U36117 ( .A(n28352), .B(n28351), .ZN(n28354) );
  XNOR2_X1 U36118 ( .A(n28354), .B(n28353), .ZN(n28355) );
  XNOR2_X1 U36119 ( .A(n51749), .B(n51648), .ZN(n28360) );
  XNOR2_X1 U36120 ( .A(n28361), .B(n28360), .ZN(n28362) );
  INV_X1 U36121 ( .A(n28364), .ZN(n28365) );
  XNOR2_X1 U36122 ( .A(n28365), .B(n28366), .ZN(n28368) );
  XNOR2_X2 U36123 ( .A(n28367), .B(n28368), .ZN(n29749) );
  INV_X1 U36124 ( .A(n28369), .ZN(n28374) );
  XNOR2_X1 U36125 ( .A(n28374), .B(n28373), .ZN(n28387) );
  XNOR2_X1 U36126 ( .A(n33050), .B(n28375), .ZN(n42243) );
  XNOR2_X1 U36127 ( .A(n44044), .B(n28376), .ZN(n28377) );
  XNOR2_X1 U36128 ( .A(n42243), .B(n28377), .ZN(n28379) );
  INV_X1 U36129 ( .A(n32553), .ZN(n28378) );
  XNOR2_X1 U36130 ( .A(n28379), .B(n28378), .ZN(n28380) );
  XNOR2_X1 U36131 ( .A(n28381), .B(n28380), .ZN(n28382) );
  XNOR2_X1 U36132 ( .A(n28383), .B(n28382), .ZN(n28384) );
  XNOR2_X1 U36133 ( .A(n28385), .B(n28384), .ZN(n28386) );
  XNOR2_X1 U36134 ( .A(n28387), .B(n28386), .ZN(n28389) );
  XNOR2_X1 U36135 ( .A(n28390), .B(n3481), .ZN(n45402) );
  XNOR2_X1 U36136 ( .A(n44887), .B(n45402), .ZN(n28393) );
  INV_X1 U36137 ( .A(n28391), .ZN(n28392) );
  XNOR2_X1 U36138 ( .A(n28393), .B(n28392), .ZN(n28394) );
  XNOR2_X1 U36139 ( .A(n28394), .B(n43852), .ZN(n28395) );
  XNOR2_X1 U36140 ( .A(n28396), .B(n28395), .ZN(n28397) );
  XNOR2_X1 U36141 ( .A(n28398), .B(n28397), .ZN(n28399) );
  XNOR2_X1 U36142 ( .A(n28403), .B(n28402), .ZN(n28406) );
  INV_X1 U36143 ( .A(n28404), .ZN(n28405) );
  AND2_X1 U36144 ( .A1(n2143), .A2(n427), .ZN(n28835) );
  NAND2_X1 U36145 ( .A1(n28841), .A2(n28835), .ZN(n30454) );
  INV_X1 U36146 ( .A(n28449), .ZN(n29747) );
  XNOR2_X1 U36147 ( .A(n28408), .B(n28407), .ZN(n28422) );
  INV_X1 U36148 ( .A(n28409), .ZN(n28420) );
  XNOR2_X1 U36149 ( .A(n28410), .B(n28411), .ZN(n28418) );
  XNOR2_X1 U36150 ( .A(n28413), .B(n28412), .ZN(n43387) );
  XNOR2_X1 U36151 ( .A(n41562), .B(n41567), .ZN(n28414) );
  XNOR2_X1 U36152 ( .A(n43387), .B(n28414), .ZN(n28415) );
  XNOR2_X1 U36153 ( .A(n51646), .B(n28415), .ZN(n28417) );
  XNOR2_X1 U36154 ( .A(n28418), .B(n28417), .ZN(n28419) );
  XNOR2_X1 U36155 ( .A(n28420), .B(n28419), .ZN(n28421) );
  NAND4_X1 U36156 ( .A1(n29747), .A2(n2143), .A3(n29749), .A4(n30458), .ZN(
        n30447) );
  INV_X1 U36157 ( .A(n29749), .ZN(n28998) );
  XNOR2_X1 U36158 ( .A(n28423), .B(n28424), .ZN(n28429) );
  XNOR2_X1 U36159 ( .A(n35532), .B(n28425), .ZN(n43288) );
  XNOR2_X1 U36160 ( .A(n41597), .B(n43288), .ZN(n28426) );
  XNOR2_X1 U36161 ( .A(n28427), .B(n28426), .ZN(n28428) );
  XNOR2_X1 U36162 ( .A(n28429), .B(n28428), .ZN(n28435) );
  XNOR2_X1 U36163 ( .A(n28430), .B(n28431), .ZN(n28433) );
  XNOR2_X1 U36164 ( .A(n28432), .B(n28433), .ZN(n28434) );
  XNOR2_X1 U36165 ( .A(n28435), .B(n28434), .ZN(n28436) );
  XNOR2_X1 U36166 ( .A(n28437), .B(n28436), .ZN(n28443) );
  XNOR2_X1 U36167 ( .A(n28438), .B(n28439), .ZN(n28441) );
  INV_X1 U36168 ( .A(n25752), .ZN(n28440) );
  XNOR2_X1 U36169 ( .A(n28441), .B(n28440), .ZN(n28442) );
  XNOR2_X2 U36170 ( .A(n28443), .B(n28442), .ZN(n30461) );
  NAND2_X1 U36171 ( .A1(n28523), .A2(n51693), .ZN(n30451) );
  NAND3_X1 U36172 ( .A1(n30444), .A2(n30448), .A3(n29737), .ZN(n28444) );
  OR2_X1 U36173 ( .A1(n29747), .A2(n427), .ZN(n28995) );
  OAI21_X1 U36174 ( .B1(n29736), .B2(n2143), .A(n427), .ZN(n28446) );
  XNOR2_X1 U36175 ( .A(n30459), .B(n51692), .ZN(n28517) );
  NAND3_X1 U36176 ( .A1(n28446), .A2(n28517), .A3(n28998), .ZN(n28447) );
  OAI21_X1 U36177 ( .B1(n30448), .B2(n28995), .A(n28447), .ZN(n28448) );
  NAND2_X1 U36178 ( .A1(n28448), .A2(n29737), .ZN(n28453) );
  INV_X1 U36179 ( .A(n30442), .ZN(n28521) );
  AND2_X1 U36180 ( .A1(n2143), .A2(n30461), .ZN(n30441) );
  OAI21_X1 U36181 ( .B1(n28839), .B2(n28521), .A(n30441), .ZN(n28452) );
  INV_X1 U36182 ( .A(n28841), .ZN(n30462) );
  NOR2_X1 U36183 ( .A1(n30462), .A2(n30458), .ZN(n28827) );
  NOR2_X1 U36184 ( .A1(n28995), .A2(n29740), .ZN(n28450) );
  OAI21_X1 U36185 ( .B1(n28827), .B2(n28450), .A(n30461), .ZN(n28451) );
  NAND3_X1 U36187 ( .A1(n28866), .A2(n28865), .A3(n28862), .ZN(n28456) );
  NAND2_X1 U36188 ( .A1(n28952), .A2(n29797), .ZN(n28455) );
  OAI211_X1 U36189 ( .C1(n28950), .C2(n29800), .A(n28456), .B(n28455), .ZN(
        n28457) );
  NAND2_X1 U36190 ( .A1(n28457), .A2(n5056), .ZN(n28466) );
  INV_X1 U36191 ( .A(n28865), .ZN(n29790) );
  NAND2_X1 U36192 ( .A1(n28459), .A2(n28458), .ZN(n28461) );
  NAND2_X1 U36193 ( .A1(n28867), .A2(n28951), .ZN(n28460) );
  NAND2_X1 U36194 ( .A1(n28461), .A2(n28460), .ZN(n28465) );
  INV_X1 U36195 ( .A(n28866), .ZN(n29801) );
  NOR2_X1 U36196 ( .A1(n29801), .A2(n28501), .ZN(n28961) );
  INV_X1 U36197 ( .A(n28957), .ZN(n28462) );
  NAND2_X1 U36198 ( .A1(n28961), .A2(n28462), .ZN(n28464) );
  INV_X1 U36199 ( .A(n28501), .ZN(n29804) );
  NAND4_X2 U36200 ( .A1(n28466), .A2(n28465), .A3(n28464), .A4(n28463), .ZN(
        n32760) );
  NAND2_X1 U36202 ( .A1(n28471), .A2(n32957), .ZN(n28476) );
  AOI21_X1 U36203 ( .B1(n8390), .B2(n32765), .A(n32175), .ZN(n32772) );
  NAND2_X1 U36204 ( .A1(n32965), .A2(n32760), .ZN(n28472) );
  NAND2_X1 U36205 ( .A1(n28472), .A2(n32761), .ZN(n28473) );
  OAI211_X1 U36206 ( .C1(n8390), .C2(n32965), .A(n32772), .B(n28473), .ZN(
        n28475) );
  AND2_X1 U36207 ( .A1(n3754), .A2(n32761), .ZN(n32762) );
  AND2_X1 U36208 ( .A1(n32771), .A2(n32965), .ZN(n32529) );
  NAND3_X1 U36209 ( .A1(n32762), .A2(n32175), .A3(n32529), .ZN(n28474) );
  XNOR2_X1 U36211 ( .A(n34546), .B(n32741), .ZN(n34122) );
  XNOR2_X1 U36212 ( .A(n34720), .B(n51501), .ZN(n33775) );
  XNOR2_X1 U36213 ( .A(n28478), .B(n33775), .ZN(n35847) );
  XNOR2_X1 U36214 ( .A(n28479), .B(n35847), .ZN(n36306) );
  INV_X1 U36215 ( .A(n36306), .ZN(n36148) );
  INV_X1 U36216 ( .A(n31801), .ZN(n31791) );
  NAND2_X1 U36217 ( .A1(n51479), .A2(n31800), .ZN(n28481) );
  AND2_X1 U36218 ( .A1(n31886), .A2(n31870), .ZN(n28482) );
  NAND4_X1 U36219 ( .A1(n31803), .A2(n28482), .A3(n31876), .A4(n52047), .ZN(
        n28480) );
  OAI21_X1 U36220 ( .B1(n31791), .B2(n28481), .A(n28480), .ZN(n28485) );
  INV_X1 U36221 ( .A(n28482), .ZN(n28483) );
  NOR2_X1 U36222 ( .A1(n31020), .A2(n28483), .ZN(n28484) );
  NOR2_X1 U36223 ( .A1(n28485), .A2(n28484), .ZN(n28495) );
  NOR2_X1 U36224 ( .A1(n5912), .A2(n31876), .ZN(n30120) );
  NAND3_X1 U36225 ( .A1(n31882), .A2(n3104), .A3(n51479), .ZN(n28486) );
  OAI211_X1 U36226 ( .C1(n30120), .C2(n51479), .A(n28486), .B(n31799), .ZN(
        n28494) );
  AOI21_X1 U36228 ( .B1(n51743), .B2(n31019), .A(n31798), .ZN(n28491) );
  OR2_X1 U36229 ( .A1(n31873), .A2(n31883), .ZN(n30117) );
  NAND4_X1 U36230 ( .A1(n28491), .A2(n31882), .A3(n28490), .A4(n30117), .ZN(
        n28493) );
  AND2_X1 U36231 ( .A1(n31883), .A2(n31876), .ZN(n31792) );
  NOR2_X1 U36232 ( .A1(n31800), .A2(n52047), .ZN(n30121) );
  OAI21_X1 U36233 ( .B1(n31873), .B2(n31792), .A(n30121), .ZN(n28492) );
  MUX2_X1 U36234 ( .A(n29800), .B(n28496), .S(n29803), .Z(n28502) );
  AND2_X1 U36236 ( .A1(n28499), .A2(n28498), .ZN(n28500) );
  INV_X1 U36237 ( .A(n28952), .ZN(n28503) );
  NOR2_X1 U36238 ( .A1(n29800), .A2(n29790), .ZN(n28504) );
  INV_X1 U36239 ( .A(n28505), .ZN(n28506) );
  OAI21_X1 U36240 ( .B1(n28507), .B2(n28508), .A(n28506), .ZN(n28513) );
  AND2_X1 U36241 ( .A1(n28509), .A2(n28510), .ZN(n28512) );
  OAI211_X1 U36242 ( .C1(n28514), .C2(n28513), .A(n28512), .B(n28511), .ZN(
        n28515) );
  OAI211_X1 U36243 ( .C1(n29749), .C2(n29000), .A(n28996), .B(n28521), .ZN(
        n28520) );
  AND2_X1 U36244 ( .A1(n28521), .A2(n30461), .ZN(n29748) );
  NAND3_X1 U36245 ( .A1(n28841), .A2(n29748), .A3(n30451), .ZN(n28519) );
  NAND3_X1 U36246 ( .A1(n28998), .A2(n30458), .A3(n427), .ZN(n28524) );
  OAI211_X1 U36247 ( .C1(n28990), .C2(n30449), .A(n28526), .B(n28525), .ZN(
        n28527) );
  INV_X1 U36248 ( .A(n28528), .ZN(n29042) );
  OR2_X1 U36249 ( .A1(n28529), .A2(n28882), .ZN(n29044) );
  NAND4_X1 U36250 ( .A1(n28874), .A2(n28530), .A3(n29035), .A4(n28883), .ZN(
        n29041) );
  NAND4_X1 U36251 ( .A1(n28875), .A2(n28874), .A3(n29033), .A4(n28882), .ZN(
        n28531) );
  NAND4_X1 U36252 ( .A1(n29042), .A2(n29044), .A3(n29041), .A4(n28531), .ZN(
        n28544) );
  INV_X1 U36253 ( .A(n29045), .ZN(n28532) );
  NAND2_X1 U36254 ( .A1(n28532), .A2(n28879), .ZN(n28535) );
  NAND2_X1 U36255 ( .A1(n28533), .A2(n29038), .ZN(n28534) );
  INV_X1 U36256 ( .A(n28536), .ZN(n28537) );
  NAND3_X1 U36257 ( .A1(n28537), .A2(n29029), .A3(n28880), .ZN(n28541) );
  INV_X1 U36258 ( .A(n28875), .ZN(n28539) );
  INV_X1 U36259 ( .A(n28871), .ZN(n28538) );
  OAI211_X1 U36260 ( .C1(n28539), .C2(n29033), .A(n29039), .B(n28538), .ZN(
        n28540) );
  NOR2_X1 U36261 ( .A1(n2881), .A2(n28548), .ZN(n28549) );
  AOI22_X1 U36262 ( .A1(n28550), .A2(n28549), .B1(n30293), .B2(n30291), .ZN(
        n28553) );
  NAND3_X1 U36263 ( .A1(n30289), .A2(n28551), .A3(n28560), .ZN(n28552) );
  INV_X1 U36266 ( .A(n28559), .ZN(n28562) );
  OAI211_X1 U36267 ( .C1(n28563), .C2(n28562), .A(n28561), .B(n28560), .ZN(
        n28564) );
  NAND2_X1 U36268 ( .A1(n51115), .A2(n28566), .ZN(n28567) );
  NAND3_X1 U36269 ( .A1(n28569), .A2(n28568), .A3(n28567), .ZN(n28576) );
  OAI21_X1 U36270 ( .B1(n29020), .B2(n29007), .A(n29015), .ZN(n28570) );
  NAND2_X1 U36271 ( .A1(n28570), .A2(n28931), .ZN(n28574) );
  NAND2_X1 U36273 ( .A1(n51115), .A2(n28918), .ZN(n28934) );
  INV_X1 U36275 ( .A(n28597), .ZN(n32324) );
  NOR3_X1 U36276 ( .A1(n28896), .A2(n28907), .A3(n28577), .ZN(n28581) );
  OAI22_X1 U36277 ( .A1(n28579), .A2(n28578), .B1(n28897), .B2(n28903), .ZN(
        n28580) );
  NOR2_X1 U36278 ( .A1(n28581), .A2(n28580), .ZN(n28595) );
  AND2_X1 U36279 ( .A1(n28585), .A2(n28584), .ZN(n28594) );
  OAI211_X1 U36280 ( .C1(n28588), .C2(n28587), .A(n28586), .B(n28907), .ZN(
        n28593) );
  INV_X1 U36281 ( .A(n28589), .ZN(n28591) );
  NAND3_X1 U36282 ( .A1(n28591), .A2(n28590), .A3(n28898), .ZN(n28592) );
  AND2_X1 U36283 ( .A1(n32324), .A2(n32705), .ZN(n28596) );
  NAND2_X1 U36284 ( .A1(n28596), .A2(n52182), .ZN(n28598) );
  AND2_X1 U36285 ( .A1(n52182), .A2(n30140), .ZN(n30147) );
  XNOR2_X1 U36286 ( .A(n32327), .B(n32705), .ZN(n28599) );
  NAND2_X1 U36287 ( .A1(n28599), .A2(n31668), .ZN(n28600) );
  INV_X1 U36288 ( .A(n32705), .ZN(n29814) );
  NOR2_X1 U36289 ( .A1(n32335), .A2(n32331), .ZN(n30136) );
  NAND2_X1 U36290 ( .A1(n30136), .A2(n32325), .ZN(n28603) );
  AND2_X1 U36291 ( .A1(n52182), .A2(n32691), .ZN(n32688) );
  INV_X1 U36292 ( .A(n32332), .ZN(n31669) );
  NAND2_X1 U36293 ( .A1(n29618), .A2(n32600), .ZN(n32976) );
  NAND2_X1 U36294 ( .A1(n32976), .A2(n32977), .ZN(n28604) );
  NAND2_X1 U36295 ( .A1(n32600), .A2(n32590), .ZN(n30510) );
  OAI211_X1 U36296 ( .C1(n32988), .C2(n30510), .A(n30503), .B(n32974), .ZN(
        n28606) );
  XNOR2_X1 U36297 ( .A(n32595), .B(n32590), .ZN(n30516) );
  AOI21_X1 U36298 ( .B1(n30516), .B2(n29616), .A(n29622), .ZN(n28605) );
  NAND2_X1 U36299 ( .A1(n28606), .A2(n28605), .ZN(n28612) );
  INV_X1 U36300 ( .A(n28607), .ZN(n30517) );
  NAND2_X1 U36301 ( .A1(n32588), .A2(n30517), .ZN(n28611) );
  INV_X1 U36302 ( .A(n28608), .ZN(n28610) );
  NOR2_X1 U36303 ( .A1(n30510), .A2(n32990), .ZN(n28609) );
  NAND2_X1 U36304 ( .A1(n28610), .A2(n28609), .ZN(n32594) );
  XNOR2_X1 U36305 ( .A(n36672), .B(n4275), .ZN(n33070) );
  NAND3_X1 U36306 ( .A1(n28615), .A2(n28614), .A3(n29514), .ZN(n28621) );
  NAND2_X1 U36307 ( .A1(n28617), .A2(n28616), .ZN(n28620) );
  NAND2_X1 U36308 ( .A1(n28618), .A2(n29518), .ZN(n28619) );
  AND3_X1 U36309 ( .A1(n28621), .A2(n28620), .A3(n28619), .ZN(n28633) );
  NAND2_X1 U36310 ( .A1(n28622), .A2(n28626), .ZN(n28624) );
  AOI21_X1 U36311 ( .B1(n28624), .B2(n6059), .A(n28623), .ZN(n28625) );
  OAI21_X1 U36312 ( .B1(n29524), .B2(n28625), .A(n29509), .ZN(n28632) );
  NAND2_X1 U36313 ( .A1(n29529), .A2(n29535), .ZN(n28627) );
  OAI211_X1 U36314 ( .C1(n28628), .C2(n29519), .A(n28627), .B(n29514), .ZN(
        n28631) );
  AND2_X1 U36315 ( .A1(n398), .A2(n28629), .ZN(n29504) );
  NAND3_X1 U36316 ( .A1(n29505), .A2(n29526), .A3(n29504), .ZN(n28630) );
  NAND4_X2 U36317 ( .A1(n28633), .A2(n28631), .A3(n28632), .A4(n28630), .ZN(
        n30856) );
  NAND3_X1 U36318 ( .A1(n29323), .A2(n29330), .A3(n29315), .ZN(n28635) );
  NAND2_X1 U36319 ( .A1(n52177), .A2(n383), .ZN(n28634) );
  AND2_X1 U36320 ( .A1(n28635), .A2(n28634), .ZN(n28649) );
  AOI21_X1 U36321 ( .B1(n52177), .B2(n29325), .A(n51107), .ZN(n28640) );
  OAI21_X1 U36322 ( .B1(n29325), .B2(n29330), .A(n29332), .ZN(n28639) );
  NAND3_X1 U36323 ( .A1(n28640), .A2(n28641), .A3(n28639), .ZN(n28647) );
  INV_X1 U36324 ( .A(n28640), .ZN(n28645) );
  NAND2_X1 U36325 ( .A1(n28642), .A2(n28641), .ZN(n28643) );
  NAND3_X1 U36326 ( .A1(n28645), .A2(n28644), .A3(n28643), .ZN(n28646) );
  INV_X1 U36327 ( .A(n31637), .ZN(n28723) );
  NAND2_X1 U36328 ( .A1(n30856), .A2(n28723), .ZN(n31633) );
  NOR2_X1 U36330 ( .A1(n29125), .A2(n29260), .ZN(n29257) );
  NAND3_X1 U36332 ( .A1(n29264), .A2(n30231), .A3(n30226), .ZN(n30224) );
  AND2_X1 U36333 ( .A1(n30224), .A2(n28651), .ZN(n28665) );
  INV_X1 U36336 ( .A(n28654), .ZN(n28655) );
  AOI21_X1 U36337 ( .B1(n28656), .B2(n28655), .A(n29260), .ZN(n28661) );
  NAND3_X1 U36338 ( .A1(n29119), .A2(n51114), .A3(n30234), .ZN(n28660) );
  OAI21_X1 U36339 ( .B1(n28667), .B2(n28666), .A(n29479), .ZN(n28668) );
  NAND3_X1 U36340 ( .A1(n28668), .A2(n28671), .A3(n2533), .ZN(n28682) );
  NOR2_X1 U36341 ( .A1(n6080), .A2(n51110), .ZN(n28670) );
  OAI21_X1 U36342 ( .B1(n28671), .B2(n28670), .A(n28669), .ZN(n28673) );
  NAND3_X1 U36343 ( .A1(n28673), .A2(n29480), .A3(n28672), .ZN(n28681) );
  INV_X1 U36344 ( .A(n28674), .ZN(n28675) );
  AOI22_X1 U36345 ( .A1(n28675), .A2(n25841), .B1(n2294), .B2(n29478), .ZN(
        n28679) );
  INV_X1 U36346 ( .A(n28676), .ZN(n28677) );
  NAND2_X1 U36347 ( .A1(n29495), .A2(n28677), .ZN(n28678) );
  NAND2_X1 U36348 ( .A1(n31633), .A2(n31634), .ZN(n28721) );
  INV_X1 U36349 ( .A(n29311), .ZN(n28685) );
  OAI22_X1 U36350 ( .A1(n28685), .A2(n28684), .B1(n28699), .B2(n28683), .ZN(
        n28687) );
  OAI21_X1 U36351 ( .B1(n28690), .B2(n28689), .A(n28688), .ZN(n28691) );
  NAND3_X1 U36352 ( .A1(n28691), .A2(n28700), .A3(n26077), .ZN(n28694) );
  INV_X1 U36353 ( .A(n28692), .ZN(n28693) );
  AND2_X1 U36354 ( .A1(n28694), .A2(n28693), .ZN(n28707) );
  INV_X1 U36355 ( .A(n29295), .ZN(n28697) );
  NAND2_X1 U36356 ( .A1(n28696), .A2(n28695), .ZN(n29312) );
  AND2_X1 U36357 ( .A1(n28697), .A2(n29312), .ZN(n28706) );
  NAND2_X1 U36359 ( .A1(n28700), .A2(n28699), .ZN(n28703) );
  NAND3_X1 U36360 ( .A1(n28701), .A2(n29309), .A3(n51517), .ZN(n28702) );
  NAND4_X1 U36361 ( .A1(n28704), .A2(n29291), .A3(n28703), .A4(n28702), .ZN(
        n28705) );
  OAI22_X1 U36362 ( .A1(n28708), .A2(n28715), .B1(n29190), .B2(n29185), .ZN(
        n28709) );
  OAI21_X1 U36363 ( .B1(n29181), .B2(n28709), .A(n29192), .ZN(n28719) );
  OAI22_X1 U36364 ( .A1(n28715), .A2(n7052), .B1(n29269), .B2(n29191), .ZN(
        n28712) );
  INV_X1 U36365 ( .A(n28714), .ZN(n28716) );
  OAI211_X1 U36366 ( .C1(n28717), .C2(n28716), .A(n29191), .B(n28715), .ZN(
        n28718) );
  NAND2_X1 U36367 ( .A1(n30855), .A2(n30853), .ZN(n31622) );
  OR2_X1 U36369 ( .A1(n31624), .A2(n30854), .ZN(n30861) );
  NAND2_X1 U36370 ( .A1(n28722), .A2(n30861), .ZN(n28728) );
  INV_X1 U36371 ( .A(n30855), .ZN(n31586) );
  AND2_X1 U36374 ( .A1(n30856), .A2(n31637), .ZN(n31580) );
  NOR2_X1 U36375 ( .A1(n30856), .A2(n31637), .ZN(n30559) );
  OAI211_X1 U36376 ( .C1(n30559), .C2(n30853), .A(n28724), .B(n31586), .ZN(
        n28726) );
  NAND3_X1 U36377 ( .A1(n31632), .A2(n31631), .A3(n30853), .ZN(n28725) );
  INV_X1 U36378 ( .A(n28729), .ZN(n28730) );
  XNOR2_X1 U36379 ( .A(n28731), .B(n28730), .ZN(n28732) );
  XNOR2_X1 U36380 ( .A(n35512), .B(n28732), .ZN(n28733) );
  XNOR2_X1 U36381 ( .A(n33070), .B(n28733), .ZN(n28734) );
  XNOR2_X1 U36382 ( .A(n32757), .B(n28734), .ZN(n29102) );
  NAND3_X1 U36383 ( .A1(n29859), .A2(n487), .A3(n30434), .ZN(n28735) );
  INV_X1 U36384 ( .A(n29703), .ZN(n29863) );
  INV_X1 U36385 ( .A(n28736), .ZN(n28749) );
  INV_X1 U36386 ( .A(n28737), .ZN(n28740) );
  INV_X1 U36387 ( .A(n29692), .ZN(n29872) );
  OR2_X1 U36388 ( .A1(n29872), .A2(n28739), .ZN(n29861) );
  INV_X1 U36389 ( .A(n28741), .ZN(n28748) );
  AND3_X1 U36390 ( .A1(n30433), .A2(n51746), .A3(n487), .ZN(n28744) );
  INV_X1 U36391 ( .A(n29873), .ZN(n28742) );
  NOR2_X1 U36392 ( .A1(n28742), .A2(n30425), .ZN(n28743) );
  AOI22_X1 U36393 ( .A1(n728), .A2(n28744), .B1(n28743), .B2(n30434), .ZN(
        n28747) );
  NAND4_X2 U36394 ( .A1(n28748), .A2(n28749), .A3(n28747), .A4(n28746), .ZN(
        n32900) );
  INV_X1 U36395 ( .A(n32900), .ZN(n32916) );
  INV_X1 U36396 ( .A(n30399), .ZN(n29942) );
  OAI22_X1 U36397 ( .A1(n30392), .A2(n30694), .B1(n29942), .B2(n30387), .ZN(
        n28751) );
  INV_X1 U36398 ( .A(n29931), .ZN(n28752) );
  NAND3_X1 U36399 ( .A1(n30392), .A2(n30688), .A3(n1906), .ZN(n28755) );
  NAND2_X1 U36400 ( .A1(n28752), .A2(n30692), .ZN(n28753) );
  NOR2_X1 U36401 ( .A1(n29942), .A2(n402), .ZN(n28759) );
  AND2_X1 U36402 ( .A1(n28758), .A2(n51113), .ZN(n30384) );
  AND2_X1 U36403 ( .A1(n30386), .A2(n28761), .ZN(n28762) );
  INV_X1 U36404 ( .A(n28767), .ZN(n29776) );
  NAND2_X1 U36405 ( .A1(n29776), .A2(n29782), .ZN(n28770) );
  INV_X1 U36406 ( .A(n29880), .ZN(n28769) );
  INV_X1 U36407 ( .A(n30381), .ZN(n28768) );
  OAI211_X1 U36408 ( .C1(n2077), .C2(n28770), .A(n28769), .B(n28768), .ZN(
        n28775) );
  NAND2_X1 U36409 ( .A1(n30382), .A2(n28772), .ZN(n29881) );
  INV_X1 U36410 ( .A(n28771), .ZN(n29775) );
  AOI22_X1 U36411 ( .A1(n28773), .A2(n29775), .B1(n28772), .B2(n30376), .ZN(
        n28774) );
  AND2_X1 U36412 ( .A1(n28774), .A2(n28775), .ZN(n28776) );
  MUX2_X1 U36413 ( .A(n28779), .B(n29068), .S(n30351), .Z(n28782) );
  INV_X1 U36414 ( .A(n30340), .ZN(n29055) );
  NAND3_X1 U36415 ( .A1(n28849), .A2(n29055), .A3(n30338), .ZN(n28780) );
  NAND3_X1 U36416 ( .A1(n29063), .A2(n29060), .A3(n28780), .ZN(n28781) );
  INV_X1 U36417 ( .A(n29066), .ZN(n28784) );
  NAND2_X1 U36418 ( .A1(n28298), .A2(n7721), .ZN(n28785) );
  NOR2_X1 U36419 ( .A1(n30349), .A2(n28785), .ZN(n29758) );
  NOR2_X1 U36420 ( .A1(n28786), .A2(n29758), .ZN(n28816) );
  INV_X1 U36421 ( .A(n28787), .ZN(n29067) );
  NAND2_X1 U36422 ( .A1(n514), .A2(n745), .ZN(n29053) );
  NOR2_X1 U36423 ( .A1(n29053), .A2(n5389), .ZN(n29770) );
  INV_X1 U36424 ( .A(n30339), .ZN(n29769) );
  OAI21_X1 U36425 ( .B1(n29715), .B2(n28970), .A(n28973), .ZN(n30417) );
  NAND2_X1 U36426 ( .A1(n28793), .A2(n51108), .ZN(n29713) );
  NOR2_X1 U36427 ( .A1(n30419), .A2(n28187), .ZN(n28788) );
  AND2_X1 U36428 ( .A1(n29713), .A2(n28788), .ZN(n30416) );
  XNOR2_X1 U36429 ( .A(n28187), .B(n51108), .ZN(n28977) );
  INV_X1 U36430 ( .A(n28789), .ZN(n28790) );
  NAND3_X1 U36431 ( .A1(n28791), .A2(n28977), .A3(n28790), .ZN(n28795) );
  INV_X1 U36432 ( .A(n28797), .ZN(n29727) );
  OAI211_X1 U36433 ( .C1(n29727), .C2(n28793), .A(n28973), .B(n28792), .ZN(
        n28794) );
  OAI22_X1 U36434 ( .A1(n51108), .A2(n51342), .B1(n28797), .B2(n28796), .ZN(
        n28798) );
  INV_X1 U36435 ( .A(n29855), .ZN(n28802) );
  OAI21_X1 U36436 ( .B1(n28807), .B2(n28802), .A(n29848), .ZN(n28803) );
  NOR2_X1 U36437 ( .A1(n2169), .A2(n30711), .ZN(n28806) );
  AOI21_X1 U36438 ( .B1(n2205), .B2(n30706), .A(n30721), .ZN(n28805) );
  NAND2_X1 U36439 ( .A1(n2169), .A2(n30711), .ZN(n28804) );
  OAI211_X1 U36440 ( .C1(n28806), .C2(n30709), .A(n28805), .B(n28804), .ZN(
        n28811) );
  AND2_X1 U36441 ( .A1(n32915), .A2(n32917), .ZN(n32922) );
  NAND2_X1 U36442 ( .A1(n32900), .A2(n32908), .ZN(n30820) );
  NOR2_X1 U36443 ( .A1(n32915), .A2(n30820), .ZN(n28815) );
  INV_X1 U36444 ( .A(n28812), .ZN(n28813) );
  AOI22_X1 U36445 ( .A1(n28815), .A2(n28814), .B1(n28813), .B2(n30822), .ZN(
        n28825) );
  AND2_X1 U36446 ( .A1(n32895), .A2(n32909), .ZN(n32639) );
  NOR2_X1 U36447 ( .A1(n32634), .A2(n32633), .ZN(n28822) );
  NAND2_X1 U36448 ( .A1(n28817), .A2(n28816), .ZN(n28820) );
  INV_X1 U36449 ( .A(n28818), .ZN(n28819) );
  OAI21_X1 U36450 ( .B1(n28820), .B2(n28819), .A(n32633), .ZN(n28821) );
  AOI22_X1 U36451 ( .A1(n32639), .A2(n28822), .B1(n32907), .B2(n28821), .ZN(
        n28824) );
  INV_X1 U36453 ( .A(n28827), .ZN(n28828) );
  OR2_X1 U36454 ( .A1(n30461), .A2(n427), .ZN(n29745) );
  AOI21_X1 U36455 ( .B1(n28828), .B2(n30447), .A(n29745), .ZN(n28834) );
  AND2_X1 U36456 ( .A1(n427), .A2(n29737), .ZN(n28840) );
  OAI21_X1 U36457 ( .B1(n29749), .B2(n28523), .A(n29734), .ZN(n28830) );
  NOR2_X1 U36459 ( .A1(n28834), .A2(n28833), .ZN(n28847) );
  AOI21_X1 U36460 ( .B1(n28991), .B2(n51692), .A(n29737), .ZN(n28837) );
  MUX2_X1 U36461 ( .A(n28991), .B(n28835), .S(n30458), .Z(n28836) );
  AOI22_X1 U36462 ( .A1(n28838), .A2(n28837), .B1(n30444), .B2(n28836), .ZN(
        n28846) );
  NAND3_X1 U36463 ( .A1(n28841), .A2(n28840), .A3(n29740), .ZN(n28843) );
  AND2_X1 U36464 ( .A1(n30461), .A2(n28998), .ZN(n29741) );
  NAND2_X1 U36465 ( .A1(n29741), .A2(n29736), .ZN(n28842) );
  NAND2_X1 U36466 ( .A1(n30446), .A2(n28998), .ZN(n28844) );
  AND2_X1 U36468 ( .A1(n30348), .A2(n7721), .ZN(n29070) );
  NOR2_X1 U36469 ( .A1(n29764), .A2(n30346), .ZN(n28848) );
  OAI21_X1 U36470 ( .B1(n51490), .B2(n28848), .A(n5389), .ZN(n28850) );
  INV_X1 U36471 ( .A(n28852), .ZN(n29765) );
  NAND2_X1 U36472 ( .A1(n29765), .A2(n29063), .ZN(n28856) );
  INV_X1 U36473 ( .A(n28853), .ZN(n28854) );
  OAI21_X1 U36474 ( .B1(n28854), .B2(n29763), .A(n29760), .ZN(n28855) );
  NOR2_X1 U36475 ( .A1(n32843), .A2(n30484), .ZN(n28941) );
  AND2_X1 U36476 ( .A1(n28957), .A2(n28951), .ZN(n28859) );
  AOI22_X1 U36477 ( .A1(n28859), .A2(n28952), .B1(n28858), .B2(n28865), .ZN(
        n28869) );
  OAI21_X1 U36478 ( .B1(n28862), .B2(n28950), .A(n28860), .ZN(n28861) );
  AOI22_X1 U36479 ( .A1(n29796), .A2(n29804), .B1(n5056), .B2(n28861), .ZN(
        n28864) );
  OR2_X1 U36480 ( .A1(n28953), .A2(n5056), .ZN(n28863) );
  NAND2_X1 U36481 ( .A1(n28866), .A2(n28865), .ZN(n28955) );
  NAND4_X2 U36482 ( .A1(n28869), .A2(n28868), .A3(n28955), .A4(n29789), .ZN(
        n32386) );
  OAI21_X1 U36483 ( .B1(n28871), .B2(n28870), .A(n29035), .ZN(n28873) );
  NAND3_X1 U36484 ( .A1(n28873), .A2(n28872), .A3(n29038), .ZN(n28888) );
  NAND3_X1 U36485 ( .A1(n28875), .A2(n29035), .A3(n28874), .ZN(n28876) );
  NAND4_X1 U36486 ( .A1(n28878), .A2(n28877), .A3(n28876), .A4(n29033), .ZN(
        n28887) );
  NAND3_X1 U36487 ( .A1(n29045), .A2(n28880), .A3(n28879), .ZN(n28886) );
  INV_X1 U36488 ( .A(n28881), .ZN(n28884) );
  NAND3_X1 U36489 ( .A1(n28884), .A2(n28883), .A3(n28882), .ZN(n28885) );
  NAND4_X2 U36490 ( .A1(n28888), .A2(n28887), .A3(n28886), .A4(n28885), .ZN(
        n31910) );
  INV_X1 U36491 ( .A(n28889), .ZN(n28891) );
  OAI21_X1 U36492 ( .B1(n28891), .B2(n28904), .A(n28890), .ZN(n28892) );
  INV_X1 U36493 ( .A(n28892), .ZN(n28912) );
  INV_X1 U36494 ( .A(n28893), .ZN(n28901) );
  NAND2_X1 U36495 ( .A1(n28895), .A2(n28894), .ZN(n28900) );
  OAI21_X1 U36496 ( .B1(n28901), .B2(n28900), .A(n28899), .ZN(n28902) );
  INV_X1 U36497 ( .A(n28902), .ZN(n28911) );
  OAI22_X1 U36498 ( .A1(n28904), .A2(n28903), .B1(n28907), .B2(n27991), .ZN(
        n28906) );
  NAND2_X1 U36499 ( .A1(n28906), .A2(n28905), .ZN(n28910) );
  NAND2_X1 U36500 ( .A1(n28908), .A2(n28907), .ZN(n28909) );
  NAND4_X2 U36501 ( .A1(n28912), .A2(n28911), .A3(n28910), .A4(n28909), .ZN(
        n32841) );
  NAND2_X1 U36502 ( .A1(n32386), .A2(n31910), .ZN(n28913) );
  NAND2_X1 U36503 ( .A1(n28913), .A2(n31075), .ZN(n28914) );
  NAND3_X1 U36504 ( .A1(n28916), .A2(n29011), .A3(n29013), .ZN(n28917) );
  NAND2_X1 U36505 ( .A1(n29012), .A2(n28917), .ZN(n28921) );
  OAI22_X1 U36506 ( .A1(n51115), .A2(n28918), .B1(n29014), .B2(n28923), .ZN(
        n28920) );
  AOI21_X1 U36507 ( .B1(n28921), .B2(n29020), .A(n28920), .ZN(n28930) );
  INV_X1 U36508 ( .A(n28922), .ZN(n28925) );
  NAND2_X1 U36509 ( .A1(n28923), .A2(n29013), .ZN(n28924) );
  OAI22_X1 U36510 ( .A1(n28925), .A2(n28924), .B1(n29006), .B2(n28927), .ZN(
        n28929) );
  AOI21_X1 U36511 ( .B1(n28927), .B2(n7226), .A(n28926), .ZN(n28928) );
  OAI22_X1 U36512 ( .A1(n28930), .A2(n28929), .B1(n28928), .B2(n29020), .ZN(
        n28938) );
  AOI21_X1 U36513 ( .B1(n28932), .B2(n29020), .A(n28931), .ZN(n28989) );
  INV_X1 U36514 ( .A(n28934), .ZN(n28935) );
  NAND3_X1 U36515 ( .A1(n28935), .A2(n29007), .A3(n29006), .ZN(n28936) );
  INV_X1 U36516 ( .A(n31910), .ZN(n32840) );
  NAND3_X1 U36517 ( .A1(n32844), .A2(n32840), .A3(n32843), .ZN(n30497) );
  NOR2_X1 U36518 ( .A1(n32841), .A2(n32386), .ZN(n30483) );
  NAND3_X1 U36519 ( .A1(n31914), .A2(n32385), .A3(n30483), .ZN(n28939) );
  NAND2_X1 U36520 ( .A1(n30484), .A2(n31910), .ZN(n31078) );
  OR2_X1 U36521 ( .A1(n31078), .A2(n32385), .ZN(n32374) );
  OAI21_X1 U36522 ( .B1(n32850), .B2(n32836), .A(n32374), .ZN(n28942) );
  NAND2_X1 U36523 ( .A1(n28942), .A2(n32843), .ZN(n28944) );
  OR2_X1 U36524 ( .A1(n30484), .A2(n31910), .ZN(n32377) );
  OAI21_X1 U36526 ( .B1(n31920), .B2(n32385), .A(n30495), .ZN(n28943) );
  XNOR2_X1 U36528 ( .A(n34381), .B(n51446), .ZN(n29084) );
  OAI21_X1 U36529 ( .B1(n28948), .B2(n28957), .A(n28947), .ZN(n28949) );
  NAND2_X1 U36530 ( .A1(n28949), .A2(n29790), .ZN(n28956) );
  NAND3_X1 U36531 ( .A1(n28952), .A2(n28951), .A3(n28950), .ZN(n29791) );
  AND4_X1 U36532 ( .A1(n28956), .A2(n28955), .A3(n29791), .A4(n28954), .ZN(
        n28960) );
  INV_X1 U36533 ( .A(n28962), .ZN(n28964) );
  OAI21_X1 U36534 ( .B1(n28965), .B2(n28964), .A(n28963), .ZN(n28966) );
  NOR2_X1 U36535 ( .A1(n28967), .A2(n28966), .ZN(n28968) );
  OAI21_X1 U36536 ( .B1(n28971), .B2(n28187), .A(n30403), .ZN(n30401) );
  OAI21_X1 U36537 ( .B1(n30419), .B2(n28970), .A(n30401), .ZN(n28972) );
  NAND2_X1 U36538 ( .A1(n28971), .A2(n28974), .ZN(n29728) );
  NAND3_X1 U36539 ( .A1(n28972), .A2(n30407), .A3(n29728), .ZN(n28988) );
  INV_X1 U36540 ( .A(n28973), .ZN(n30418) );
  MUX2_X1 U36541 ( .A(n30421), .B(n30418), .S(n30404), .Z(n28976) );
  NAND2_X1 U36542 ( .A1(n28974), .A2(n28189), .ZN(n28975) );
  NAND2_X1 U36543 ( .A1(n28976), .A2(n28975), .ZN(n28987) );
  INV_X1 U36544 ( .A(n30413), .ZN(n28981) );
  INV_X1 U36545 ( .A(n28977), .ZN(n28978) );
  NAND2_X1 U36546 ( .A1(n29727), .A2(n28982), .ZN(n28984) );
  INV_X1 U36547 ( .A(n28990), .ZN(n28992) );
  OAI22_X1 U36548 ( .A1(n28992), .A2(n28996), .B1(n28991), .B2(n30448), .ZN(
        n28994) );
  INV_X1 U36549 ( .A(n30446), .ZN(n28993) );
  AOI21_X1 U36550 ( .B1(n28994), .B2(n28993), .A(n28998), .ZN(n29005) );
  INV_X1 U36552 ( .A(n28996), .ZN(n28997) );
  NAND3_X1 U36553 ( .A1(n29000), .A2(n29749), .A3(n427), .ZN(n29001) );
  NAND2_X1 U36554 ( .A1(n29001), .A2(n29737), .ZN(n29002) );
  NAND2_X1 U36555 ( .A1(n29002), .A2(n29736), .ZN(n29003) );
  OR2_X2 U36556 ( .A1(n29005), .A2(n29004), .ZN(n32876) );
  NAND3_X1 U36557 ( .A1(n29006), .A2(n29011), .A3(n29013), .ZN(n29010) );
  OAI211_X1 U36558 ( .C1(n29011), .C2(n29015), .A(n29010), .B(n29009), .ZN(
        n29022) );
  INV_X1 U36559 ( .A(n29012), .ZN(n29019) );
  AOI21_X1 U36560 ( .B1(n29015), .B2(n29014), .A(n29013), .ZN(n29017) );
  AOI22_X1 U36561 ( .A1(n29019), .A2(n29018), .B1(n29017), .B2(n29016), .ZN(
        n29021) );
  MUX2_X1 U36562 ( .A(n29022), .B(n29021), .S(n29020), .Z(n29026) );
  AND2_X2 U36563 ( .A1(n29026), .A2(n29025), .ZN(n32867) );
  NAND2_X1 U36564 ( .A1(n8544), .A2(n33030), .ZN(n31530) );
  OAI21_X1 U36565 ( .B1(n29029), .B2(n29028), .A(n29027), .ZN(n29031) );
  NAND3_X1 U36566 ( .A1(n29031), .A2(n29030), .A3(n29032), .ZN(n29037) );
  NAND3_X1 U36567 ( .A1(n29034), .A2(n29033), .A3(n29032), .ZN(n29036) );
  MUX2_X1 U36568 ( .A(n29037), .B(n29036), .S(n29035), .Z(n29050) );
  AND4_X1 U36569 ( .A1(n29043), .A2(n29042), .A3(n29041), .A4(n29040), .ZN(
        n29049) );
  INV_X1 U36570 ( .A(n29044), .ZN(n29046) );
  OAI21_X1 U36571 ( .B1(n29047), .B2(n29046), .A(n29045), .ZN(n29048) );
  AND3_X2 U36572 ( .A1(n29050), .A2(n29049), .A3(n29048), .ZN(n32874) );
  NAND2_X1 U36573 ( .A1(n30969), .A2(n32876), .ZN(n29051) );
  INV_X1 U36574 ( .A(n29053), .ZN(n30355) );
  NAND3_X1 U36575 ( .A1(n51489), .A2(n745), .A3(n29065), .ZN(n29056) );
  AOI21_X1 U36576 ( .B1(n29056), .B2(n29055), .A(n29060), .ZN(n29058) );
  NAND2_X1 U36577 ( .A1(n29069), .A2(n29056), .ZN(n29057) );
  INV_X1 U36578 ( .A(n29060), .ZN(n29768) );
  OAI22_X1 U36579 ( .A1(n29768), .A2(n29068), .B1(n30349), .B2(n29061), .ZN(
        n29064) );
  OAI21_X1 U36580 ( .B1(n29067), .B2(n29066), .A(n29065), .ZN(n29073) );
  OR2_X1 U36581 ( .A1(n29068), .A2(n5389), .ZN(n29757) );
  OAI21_X1 U36582 ( .B1(n29069), .B2(n30351), .A(n29757), .ZN(n29072) );
  OAI22_X1 U36583 ( .A1(n30339), .A2(n30338), .B1(n30349), .B2(n28300), .ZN(
        n29071) );
  NAND2_X1 U36584 ( .A1(n29074), .A2(n33026), .ZN(n29083) );
  INV_X1 U36585 ( .A(n33029), .ZN(n29075) );
  NAND2_X1 U36586 ( .A1(n33041), .A2(n32867), .ZN(n29076) );
  NAND3_X1 U36587 ( .A1(n29075), .A2(n32876), .A3(n29076), .ZN(n29082) );
  OAI211_X1 U36588 ( .C1(n30969), .C2(n32876), .A(n719), .B(n29076), .ZN(
        n29078) );
  AND2_X1 U36589 ( .A1(n29078), .A2(n29077), .ZN(n29081) );
  NAND2_X1 U36590 ( .A1(n7232), .A2(n32876), .ZN(n33036) );
  OAI21_X1 U36591 ( .B1(n33036), .B2(n719), .A(n32865), .ZN(n29079) );
  NAND3_X1 U36592 ( .A1(n29079), .A2(n32867), .A3(n33026), .ZN(n29080) );
  XNOR2_X1 U36593 ( .A(n33759), .B(n29084), .ZN(n29101) );
  OR2_X1 U36594 ( .A1(n31712), .A2(n31711), .ZN(n30816) );
  NAND2_X1 U36595 ( .A1(n32125), .A2(n31700), .ZN(n29086) );
  NAND2_X1 U36596 ( .A1(n32129), .A2(n31711), .ZN(n29092) );
  OR2_X1 U36597 ( .A1(n31700), .A2(n32130), .ZN(n32136) );
  OAI211_X1 U36598 ( .C1(n31700), .C2(n31711), .A(n721), .B(n31699), .ZN(
        n29087) );
  NAND3_X1 U36600 ( .A1(n32125), .A2(n31699), .A3(n31711), .ZN(n29089) );
  NAND2_X1 U36602 ( .A1(n30007), .A2(n51240), .ZN(n30015) );
  AND2_X1 U36603 ( .A1(n29998), .A2(n31680), .ZN(n31689) );
  NAND2_X1 U36604 ( .A1(n30022), .A2(n30983), .ZN(n29093) );
  INV_X1 U36605 ( .A(n31691), .ZN(n29095) );
  NAND3_X1 U36606 ( .A1(n29966), .A2(n29998), .A3(n29095), .ZN(n29100) );
  NOR2_X1 U36607 ( .A1(n30982), .A2(n29096), .ZN(n31675) );
  NAND2_X1 U36608 ( .A1(n30982), .A2(n29096), .ZN(n31692) );
  XNOR2_X1 U36609 ( .A(n30982), .B(n51240), .ZN(n29097) );
  AND2_X1 U36610 ( .A1(n31679), .A2(n31684), .ZN(n29967) );
  NAND3_X1 U36611 ( .A1(n29097), .A2(n29967), .A3(n30983), .ZN(n29098) );
  BUF_X2 U36612 ( .A(n35048), .Z(n34020) );
  XNOR2_X1 U36613 ( .A(n29101), .B(n34020), .ZN(n33833) );
  XNOR2_X1 U36614 ( .A(n33833), .B(n29102), .ZN(n29615) );
  OR2_X1 U36615 ( .A1(n32214), .A2(n6969), .ZN(n30892) );
  NOR2_X1 U36616 ( .A1(n30892), .A2(n32215), .ZN(n29103) );
  AND2_X1 U36617 ( .A1(n50981), .A2(n32214), .ZN(n32206) );
  AND2_X1 U36618 ( .A1(n50981), .A2(n32211), .ZN(n30888) );
  NAND2_X1 U36619 ( .A1(n29105), .A2(n30888), .ZN(n29106) );
  NAND3_X1 U36621 ( .A1(n52147), .A2(n30267), .A3(n25107), .ZN(n29112) );
  NAND2_X1 U36622 ( .A1(n29235), .A2(n29110), .ZN(n29111) );
  AOI21_X1 U36623 ( .B1(n52195), .B2(n29112), .A(n29111), .ZN(n29114) );
  INV_X1 U36624 ( .A(n29242), .ZN(n30258) );
  OAI211_X1 U36625 ( .C1(n29241), .C2(n29235), .A(n25107), .B(n30258), .ZN(
        n29116) );
  INV_X1 U36627 ( .A(n29221), .ZN(n29237) );
  MUX2_X1 U36628 ( .A(n29116), .B(n29115), .S(n29237), .Z(n29117) );
  AND3_X1 U36629 ( .A1(n5564), .A2(n625), .A3(n30267), .ZN(n29238) );
  NAND3_X1 U36630 ( .A1(n29119), .A2(n29259), .A3(n30234), .ZN(n29122) );
  OAI21_X1 U36631 ( .B1(n30231), .B2(n29260), .A(n29120), .ZN(n29121) );
  MUX2_X1 U36632 ( .A(n29122), .B(n29121), .S(n29251), .Z(n29130) );
  NAND3_X1 U36633 ( .A1(n30233), .A2(n29263), .A3(n29123), .ZN(n29124) );
  MUX2_X1 U36634 ( .A(n29125), .B(n29124), .S(n30234), .Z(n29129) );
  OAI211_X1 U36635 ( .C1(n29263), .C2(n29126), .A(n29255), .B(n30228), .ZN(
        n29128) );
  NAND2_X1 U36636 ( .A1(n30227), .A2(n30218), .ZN(n29127) );
  INV_X1 U36637 ( .A(n32066), .ZN(n32408) );
  NOR2_X1 U36638 ( .A1(n2201), .A2(n1771), .ZN(n29132) );
  OAI21_X1 U36639 ( .B1(n30183), .B2(n30171), .A(n30306), .ZN(n29131) );
  OAI21_X1 U36640 ( .B1(n30178), .B2(n1771), .A(n30304), .ZN(n29135) );
  INV_X1 U36641 ( .A(n29133), .ZN(n29134) );
  AOI22_X1 U36642 ( .A1(n29136), .A2(n29135), .B1(n29134), .B2(n30167), .ZN(
        n29145) );
  INV_X1 U36643 ( .A(n30167), .ZN(n30313) );
  INV_X1 U36644 ( .A(n29137), .ZN(n30186) );
  OAI22_X1 U36646 ( .A1(n3368), .A2(n29141), .B1(n30181), .B2(n739), .ZN(
        n29142) );
  NAND2_X1 U36647 ( .A1(n29142), .A2(n30165), .ZN(n29143) );
  INV_X1 U36648 ( .A(n29174), .ZN(n29146) );
  INV_X1 U36649 ( .A(n29152), .ZN(n29154) );
  INV_X1 U36651 ( .A(n29172), .ZN(n29173) );
  AND2_X1 U36652 ( .A1(n30249), .A2(n29155), .ZN(n29157) );
  NAND4_X1 U36654 ( .A1(n29163), .A2(n29162), .A3(n29161), .A4(n29160), .ZN(
        n29164) );
  NOR2_X1 U36655 ( .A1(n29165), .A2(n29164), .ZN(n29180) );
  INV_X1 U36656 ( .A(n29166), .ZN(n29179) );
  NAND2_X1 U36657 ( .A1(n29167), .A2(n29174), .ZN(n29168) );
  OAI21_X1 U36658 ( .B1(n29174), .B2(n30249), .A(n29173), .ZN(n29175) );
  NAND2_X1 U36659 ( .A1(n29176), .A2(n29175), .ZN(n29177) );
  BUF_X2 U36660 ( .A(n29211), .Z(n32396) );
  NOR2_X1 U36661 ( .A1(n29183), .A2(n5425), .ZN(n29280) );
  OAI21_X1 U36662 ( .B1(n29281), .B2(n29189), .A(n29188), .ZN(n29196) );
  AOI21_X1 U36663 ( .B1(n29191), .B2(n29190), .A(n51706), .ZN(n29194) );
  OAI22_X1 U36664 ( .A1(n29282), .A2(n7052), .B1(n29270), .B2(n29192), .ZN(
        n29193) );
  OAI21_X1 U36665 ( .B1(n29194), .B2(n29283), .A(n29193), .ZN(n29195) );
  NOR2_X1 U36666 ( .A1(n32066), .A2(n32401), .ZN(n32071) );
  AND2_X1 U36667 ( .A1(n29343), .A2(n30202), .ZN(n30192) );
  AOI21_X1 U36668 ( .B1(n30203), .B2(n30194), .A(n30192), .ZN(n29208) );
  AND2_X1 U36669 ( .A1(n29200), .A2(n29199), .ZN(n29201) );
  OAI21_X1 U36670 ( .B1(n29202), .B2(n29201), .A(n29351), .ZN(n29207) );
  NOR2_X1 U36671 ( .A1(n29203), .A2(n30200), .ZN(n29352) );
  INV_X1 U36672 ( .A(n29205), .ZN(n29206) );
  OAI211_X1 U36673 ( .C1(n32071), .C2(n32402), .A(n32075), .B(n32407), .ZN(
        n29210) );
  OAI21_X1 U36674 ( .B1(n31947), .B2(n31280), .A(n29210), .ZN(n29213) );
  NAND3_X1 U36675 ( .A1(n32080), .A2(n32408), .A3(n32402), .ZN(n29212) );
  OR2_X1 U36677 ( .A1(n32402), .A2(n32080), .ZN(n31289) );
  OAI211_X1 U36679 ( .C1(n32081), .C2(n31289), .A(n29214), .B(n51639), .ZN(
        n29217) );
  AND2_X1 U36680 ( .A1(n32396), .A2(n32402), .ZN(n31950) );
  XNOR2_X1 U36681 ( .A(n51519), .B(n32066), .ZN(n29215) );
  NAND3_X1 U36682 ( .A1(n31950), .A2(n714), .A3(n29215), .ZN(n29216) );
  NAND4_X2 U36683 ( .A1(n32065), .A2(n29217), .A3(n29218), .A4(n29216), .ZN(
        n35606) );
  XNOR2_X1 U36684 ( .A(n35606), .B(n36930), .ZN(n29362) );
  INV_X1 U36685 ( .A(n29219), .ZN(n29224) );
  NOR2_X1 U36686 ( .A1(n29221), .A2(n30263), .ZN(n29223) );
  INV_X1 U36687 ( .A(n29222), .ZN(n29231) );
  NAND2_X1 U36688 ( .A1(n52102), .A2(n25107), .ZN(n29225) );
  OR2_X1 U36689 ( .A1(n29226), .A2(n29225), .ZN(n29228) );
  NAND2_X1 U36690 ( .A1(n29228), .A2(n29227), .ZN(n29230) );
  NAND2_X1 U36691 ( .A1(n29228), .A2(n30263), .ZN(n29229) );
  MUX2_X1 U36692 ( .A(n30269), .B(n1708), .S(n6486), .Z(n29236) );
  OAI21_X1 U36693 ( .B1(n29236), .B2(n29235), .A(n29234), .ZN(n29246) );
  NAND2_X1 U36694 ( .A1(n29238), .A2(n29237), .ZN(n29245) );
  NAND3_X1 U36695 ( .A1(n29242), .A2(n29241), .A3(n25418), .ZN(n29243) );
  NAND3_X1 U36696 ( .A1(n29248), .A2(n30231), .A3(n29247), .ZN(n29250) );
  OAI211_X1 U36697 ( .C1(n29252), .C2(n29251), .A(n29250), .B(n29249), .ZN(
        n29253) );
  INV_X1 U36698 ( .A(n29253), .ZN(n29268) );
  INV_X1 U36699 ( .A(n30228), .ZN(n30219) );
  NOR2_X1 U36700 ( .A1(n29254), .A2(n30219), .ZN(n29258) );
  INV_X1 U36701 ( .A(n29255), .ZN(n29256) );
  OAI21_X1 U36702 ( .B1(n29258), .B2(n29257), .A(n29256), .ZN(n29267) );
  XNOR2_X1 U36703 ( .A(n29260), .B(n29259), .ZN(n29262) );
  NAND2_X1 U36704 ( .A1(n29262), .A2(n29261), .ZN(n29266) );
  NAND3_X1 U36705 ( .A1(n29264), .A2(n29263), .A3(n30218), .ZN(n29265) );
  NAND4_X2 U36706 ( .A1(n29268), .A2(n29267), .A3(n29266), .A4(n29265), .ZN(
        n32558) );
  NAND2_X1 U36707 ( .A1(n32088), .A2(n32558), .ZN(n29313) );
  OAI22_X1 U36708 ( .A1(n29272), .A2(n29271), .B1(n29270), .B2(n29269), .ZN(
        n29275) );
  INV_X1 U36709 ( .A(n29273), .ZN(n29274) );
  NOR2_X1 U36710 ( .A1(n29275), .A2(n29274), .ZN(n29276) );
  INV_X1 U36711 ( .A(n29280), .ZN(n29286) );
  INV_X1 U36712 ( .A(n29281), .ZN(n29285) );
  NAND3_X1 U36713 ( .A1(n29286), .A2(n29285), .A3(n29284), .ZN(n29287) );
  AND2_X1 U36714 ( .A1(n51517), .A2(n29308), .ZN(n29293) );
  OAI21_X1 U36715 ( .B1(n29291), .B2(n29290), .A(n29289), .ZN(n29292) );
  INV_X1 U36716 ( .A(n29296), .ZN(n29298) );
  NAND3_X1 U36717 ( .A1(n29298), .A2(n26077), .A3(n29309), .ZN(n29302) );
  INV_X1 U36718 ( .A(n29299), .ZN(n29310) );
  NAND3_X1 U36719 ( .A1(n29310), .A2(n29300), .A3(n29308), .ZN(n29301) );
  NAND3_X1 U36720 ( .A1(n29303), .A2(n29302), .A3(n29301), .ZN(n29307) );
  NOR2_X1 U36721 ( .A1(n29313), .A2(n30898), .ZN(n32111) );
  NAND2_X1 U36722 ( .A1(n31608), .A2(n32558), .ZN(n29829) );
  NOR2_X1 U36723 ( .A1(n29829), .A2(n32107), .ZN(n29336) );
  OAI22_X1 U36724 ( .A1(n29316), .A2(n29332), .B1(n29315), .B2(n29314), .ZN(
        n29318) );
  AOI22_X1 U36725 ( .A1(n29321), .A2(n29326), .B1(n29320), .B2(n29319), .ZN(
        n29335) );
  OAI211_X1 U36726 ( .C1(n29325), .C2(n29324), .A(n29323), .B(n51793), .ZN(
        n29334) );
  OAI211_X1 U36727 ( .C1(n29331), .C2(n29330), .A(n29329), .B(n29328), .ZN(
        n29333) );
  OAI21_X1 U36728 ( .B1(n32111), .B2(n29336), .A(n32089), .ZN(n29361) );
  INV_X1 U36729 ( .A(n29337), .ZN(n29341) );
  NAND2_X1 U36730 ( .A1(n735), .A2(n30209), .ZN(n30193) );
  NAND3_X1 U36731 ( .A1(n735), .A2(n733), .A3(n967), .ZN(n29338) );
  NAND3_X1 U36732 ( .A1(n30193), .A2(n30191), .A3(n29338), .ZN(n29339) );
  NAND2_X1 U36733 ( .A1(n29344), .A2(n29343), .ZN(n30213) );
  OAI21_X1 U36734 ( .B1(n29346), .B2(n29345), .A(n30213), .ZN(n29348) );
  NAND3_X1 U36735 ( .A1(n29348), .A2(n51109), .A3(n967), .ZN(n29349) );
  OAI21_X1 U36736 ( .B1(n29352), .B2(n29351), .A(n30197), .ZN(n29354) );
  AND2_X1 U36737 ( .A1(n29355), .A2(n31608), .ZN(n32576) );
  AND2_X1 U36738 ( .A1(n32107), .A2(n32558), .ZN(n30904) );
  AND2_X1 U36739 ( .A1(n32566), .A2(n32558), .ZN(n32108) );
  AOI22_X1 U36740 ( .A1(n32576), .A2(n30904), .B1(n32108), .B2(n32087), .ZN(
        n29360) );
  AND2_X1 U36741 ( .A1(n32105), .A2(n31608), .ZN(n32570) );
  AND2_X1 U36742 ( .A1(n32566), .A2(n32089), .ZN(n32573) );
  OAI21_X1 U36743 ( .B1(n32570), .B2(n624), .A(n32573), .ZN(n29359) );
  OR2_X1 U36744 ( .A1(n32566), .A2(n32560), .ZN(n29830) );
  INV_X1 U36745 ( .A(n32558), .ZN(n32574) );
  NAND2_X1 U36746 ( .A1(n32566), .A2(n32560), .ZN(n30900) );
  NAND4_X1 U36747 ( .A1(n29830), .A2(n8468), .A3(n32561), .A4(n30900), .ZN(
        n29357) );
  OAI21_X1 U36748 ( .B1(n32107), .B2(n32558), .A(n32088), .ZN(n29356) );
  NAND3_X1 U36749 ( .A1(n29357), .A2(n32096), .A3(n29356), .ZN(n29358) );
  XNOR2_X1 U36750 ( .A(n29362), .B(n34382), .ZN(n29385) );
  OR2_X1 U36751 ( .A1(n32244), .A2(n32242), .ZN(n29369) );
  NAND3_X1 U36752 ( .A1(n29369), .A2(n29363), .A3(n622), .ZN(n29368) );
  NOR2_X1 U36753 ( .A1(n32252), .A2(n31781), .ZN(n32257) );
  INV_X1 U36754 ( .A(n31240), .ZN(n32232) );
  INV_X1 U36755 ( .A(n29364), .ZN(n29365) );
  NAND3_X1 U36756 ( .A1(n29365), .A2(n32251), .A3(n32252), .ZN(n29366) );
  NAND4_X1 U36757 ( .A1(n29369), .A2(n31229), .A3(n32254), .A4(n31777), .ZN(
        n29371) );
  NAND3_X1 U36758 ( .A1(n32253), .A2(n31238), .A3(n32252), .ZN(n29370) );
  NAND2_X1 U36759 ( .A1(n30839), .A2(n32251), .ZN(n29375) );
  NAND3_X1 U36760 ( .A1(n29375), .A2(n29374), .A3(n29373), .ZN(n29376) );
  INV_X1 U36761 ( .A(n31040), .ZN(n30576) );
  NAND3_X1 U36762 ( .A1(n31039), .A2(n50986), .A3(n31826), .ZN(n29379) );
  INV_X1 U36763 ( .A(n29380), .ZN(n29383) );
  NAND2_X1 U36764 ( .A1(n31816), .A2(n31043), .ZN(n29381) );
  NAND2_X1 U36765 ( .A1(n29381), .A2(n31033), .ZN(n30852) );
  AND3_X1 U36766 ( .A1(n30592), .A2(n30912), .A3(n30911), .ZN(n29387) );
  OR2_X1 U36767 ( .A1(n30592), .A2(n30912), .ZN(n30609) );
  NOR2_X1 U36768 ( .A1(n30609), .A2(n31096), .ZN(n29386) );
  OAI211_X1 U36769 ( .C1(n30912), .C2(n29686), .A(n30593), .B(n30601), .ZN(
        n29388) );
  INV_X1 U36770 ( .A(n29388), .ZN(n29390) );
  NAND2_X1 U36771 ( .A1(n30915), .A2(n31096), .ZN(n29389) );
  AND2_X1 U36773 ( .A1(n30593), .A2(n30911), .ZN(n29392) );
  OAI21_X1 U36774 ( .B1(n30592), .B2(n30601), .A(n30602), .ZN(n29391) );
  NAND3_X1 U36775 ( .A1(n30590), .A2(n29391), .A3(n29686), .ZN(n29395) );
  XNOR2_X1 U36776 ( .A(n30599), .B(n30597), .ZN(n29393) );
  NAND2_X1 U36777 ( .A1(n29393), .A2(n29392), .ZN(n29394) );
  AND2_X1 U36778 ( .A1(n31302), .A2(n31300), .ZN(n29653) );
  OAI21_X1 U36779 ( .B1(n29653), .B2(n51086), .A(n31303), .ZN(n29397) );
  INV_X1 U36780 ( .A(n30829), .ZN(n29396) );
  NAND3_X1 U36781 ( .A1(n30834), .A2(n29396), .A3(n31300), .ZN(n30648) );
  OAI211_X1 U36782 ( .C1(n30652), .C2(n29398), .A(n29397), .B(n30648), .ZN(
        n29399) );
  NAND2_X1 U36783 ( .A1(n29399), .A2(n30824), .ZN(n29406) );
  NAND2_X1 U36784 ( .A1(n31298), .A2(n30649), .ZN(n29401) );
  NAND2_X1 U36785 ( .A1(n30640), .A2(n31300), .ZN(n29400) );
  MUX2_X1 U36786 ( .A(n29401), .B(n29400), .S(n51086), .Z(n29405) );
  OAI211_X1 U36787 ( .C1(n51085), .C2(n29403), .A(n29402), .B(n30647), .ZN(
        n29404) );
  XNOR2_X1 U36788 ( .A(n35059), .B(n36847), .ZN(n29583) );
  INV_X1 U36789 ( .A(n29407), .ZN(n29409) );
  NAND2_X1 U36790 ( .A1(n29409), .A2(n29408), .ZN(n29416) );
  NAND2_X1 U36791 ( .A1(n29411), .A2(n29410), .ZN(n29415) );
  AOI21_X1 U36792 ( .B1(n29416), .B2(n29415), .A(n29414), .ZN(n29436) );
  INV_X1 U36793 ( .A(n29417), .ZN(n29430) );
  AND2_X1 U36794 ( .A1(n29419), .A2(n29418), .ZN(n29425) );
  OAI211_X1 U36795 ( .C1(n29430), .C2(n29425), .A(n29424), .B(n29423), .ZN(
        n29434) );
  OAI21_X1 U36796 ( .B1(n29430), .B2(n29429), .A(n29428), .ZN(n29433) );
  NAND4_X1 U36797 ( .A1(n29434), .A2(n29433), .A3(n29432), .A4(n29431), .ZN(
        n29435) );
  NOR2_X1 U36798 ( .A1(n29447), .A2(n29438), .ZN(n29440) );
  XNOR2_X1 U36799 ( .A(n2213), .B(n430), .ZN(n29445) );
  NAND2_X1 U36800 ( .A1(n29445), .A2(n29444), .ZN(n29451) );
  NAND4_X1 U36801 ( .A1(n29452), .A2(n29451), .A3(n29450), .A4(n29449), .ZN(
        n29453) );
  NOR2_X1 U36802 ( .A1(n30924), .A2(n29642), .ZN(n29577) );
  NAND2_X1 U36803 ( .A1(n29458), .A2(n29457), .ZN(n29477) );
  OAI22_X1 U36804 ( .A1(n29462), .A2(n29461), .B1(n29460), .B2(n29459), .ZN(
        n29464) );
  NAND3_X1 U36805 ( .A1(n29466), .A2(n29472), .A3(n29465), .ZN(n29476) );
  NAND3_X1 U36806 ( .A1(n29471), .A2(n29468), .A3(n29467), .ZN(n29473) );
  INV_X1 U36807 ( .A(n29469), .ZN(n29470) );
  OAI22_X1 U36808 ( .A1(n29473), .A2(n29472), .B1(n29471), .B2(n29470), .ZN(
        n29474) );
  INV_X1 U36809 ( .A(n29474), .ZN(n29475) );
  AND2_X1 U36810 ( .A1(n29479), .A2(n29478), .ZN(n29482) );
  INV_X1 U36811 ( .A(n29480), .ZN(n29481) );
  AOI22_X1 U36812 ( .A1(n29495), .A2(n29482), .B1(n29496), .B2(n29481), .ZN(
        n29483) );
  INV_X1 U36813 ( .A(n29489), .ZN(n29492) );
  NAND2_X1 U36814 ( .A1(n29489), .A2(n51110), .ZN(n29490) );
  OAI211_X1 U36815 ( .C1(n29492), .C2(n29491), .A(n29490), .B(n2956), .ZN(
        n29502) );
  OAI21_X1 U36816 ( .B1(n29495), .B2(n29494), .A(n29493), .ZN(n29499) );
  NAND3_X1 U36817 ( .A1(n2294), .A2(n29496), .A3(n26676), .ZN(n29497) );
  AND4_X1 U36818 ( .A1(n29499), .A2(n29500), .A3(n29498), .A4(n29497), .ZN(
        n29501) );
  NAND2_X1 U36819 ( .A1(n30924), .A2(n29642), .ZN(n31068) );
  OAI211_X1 U36820 ( .C1(n29577), .C2(n3099), .A(n31513), .B(n31068), .ZN(
        n29575) );
  NAND3_X1 U36821 ( .A1(n29521), .A2(n29507), .A3(n29528), .ZN(n29511) );
  NAND3_X1 U36822 ( .A1(n29509), .A2(n29508), .A3(n29514), .ZN(n29510) );
  NAND2_X1 U36823 ( .A1(n29511), .A2(n29510), .ZN(n29517) );
  OAI22_X1 U36824 ( .A1(n29515), .A2(n29514), .B1(n29513), .B2(n29512), .ZN(
        n29516) );
  NOR2_X1 U36825 ( .A1(n29517), .A2(n29516), .ZN(n29540) );
  OAI21_X1 U36826 ( .B1(n29521), .B2(n729), .A(n29520), .ZN(n29523) );
  OAI21_X1 U36827 ( .B1(n29524), .B2(n29523), .A(n29522), .ZN(n29539) );
  OAI21_X1 U36828 ( .B1(n398), .B2(n29526), .A(n29525), .ZN(n29527) );
  OAI21_X1 U36829 ( .B1(n29529), .B2(n29528), .A(n29527), .ZN(n29530) );
  OAI21_X1 U36830 ( .B1(n29534), .B2(n398), .A(n6059), .ZN(n29536) );
  NAND3_X1 U36831 ( .A1(n29543), .A2(n29542), .A3(n743), .ZN(n29544) );
  NAND2_X1 U36832 ( .A1(n29548), .A2(n29547), .ZN(n29572) );
  NAND3_X1 U36833 ( .A1(n29551), .A2(n29550), .A3(n29549), .ZN(n29553) );
  NAND3_X1 U36834 ( .A1(n29557), .A2(n29556), .A3(n29555), .ZN(n29562) );
  INV_X1 U36835 ( .A(n29558), .ZN(n29560) );
  NAND3_X1 U36836 ( .A1(n29560), .A2(n29564), .A3(n29559), .ZN(n29561) );
  AND2_X1 U36837 ( .A1(n29561), .A2(n29562), .ZN(n29571) );
  NAND2_X1 U36838 ( .A1(n29564), .A2(n29563), .ZN(n29566) );
  OAI211_X1 U36839 ( .C1(n6339), .C2(n29567), .A(n29566), .B(n29565), .ZN(
        n29569) );
  NAND2_X1 U36840 ( .A1(n29569), .A2(n8454), .ZN(n29570) );
  NAND3_X1 U36841 ( .A1(n30936), .A2(n31510), .A3(n3099), .ZN(n29574) );
  AND2_X1 U36842 ( .A1(n30931), .A2(n31512), .ZN(n30091) );
  NAND3_X1 U36843 ( .A1(n30091), .A2(n3099), .A3(n31513), .ZN(n29573) );
  AND3_X1 U36844 ( .A1(n29575), .A2(n29574), .A3(n29573), .ZN(n29582) );
  INV_X1 U36845 ( .A(n30931), .ZN(n31517) );
  NAND2_X1 U36846 ( .A1(n30935), .A2(n31517), .ZN(n31515) );
  OR2_X1 U36847 ( .A1(n31512), .A2(n29642), .ZN(n31516) );
  NAND2_X1 U36848 ( .A1(n31515), .A2(n31516), .ZN(n29576) );
  NAND2_X1 U36849 ( .A1(n29577), .A2(n3099), .ZN(n31050) );
  NAND3_X1 U36850 ( .A1(n30082), .A2(n30925), .A3(n30930), .ZN(n29578) );
  NAND2_X1 U36851 ( .A1(n31050), .A2(n29578), .ZN(n29579) );
  NAND2_X1 U36852 ( .A1(n29579), .A2(n30931), .ZN(n29581) );
  NAND2_X1 U36853 ( .A1(n3099), .A2(n30925), .ZN(n30929) );
  INV_X1 U36854 ( .A(n31512), .ZN(n29641) );
  XNOR2_X1 U36855 ( .A(n37066), .B(n29583), .ZN(n34146) );
  NAND3_X1 U36856 ( .A1(n31122), .A2(n31116), .A3(n30940), .ZN(n31125) );
  AND2_X1 U36857 ( .A1(n30058), .A2(n362), .ZN(n29953) );
  NAND3_X1 U36858 ( .A1(n29953), .A2(n29592), .A3(n31115), .ZN(n30066) );
  OAI21_X1 U36860 ( .B1(n30943), .B2(n29591), .A(n7957), .ZN(n29585) );
  NAND2_X1 U36861 ( .A1(n30073), .A2(n7957), .ZN(n29586) );
  OAI22_X1 U36862 ( .A1(n29587), .A2(n623), .B1(n30941), .B2(n29586), .ZN(
        n29590) );
  NAND3_X1 U36863 ( .A1(n29588), .A2(n31106), .A3(n52121), .ZN(n29589) );
  NAND2_X1 U36864 ( .A1(n29590), .A2(n29589), .ZN(n29596) );
  NAND3_X1 U36865 ( .A1(n29592), .A2(n31106), .A3(n31116), .ZN(n29594) );
  NAND2_X1 U36866 ( .A1(n29592), .A2(n29591), .ZN(n29593) );
  MUX2_X1 U36867 ( .A(n29594), .B(n29593), .S(n30057), .Z(n29595) );
  NOR2_X1 U36868 ( .A1(n31931), .A2(n30043), .ZN(n30031) );
  OAI21_X1 U36869 ( .B1(n51744), .B2(n29602), .A(n31338), .ZN(n29598) );
  NOR2_X1 U36870 ( .A1(n30037), .A2(n29598), .ZN(n29600) );
  AOI22_X1 U36871 ( .A1(n30031), .A2(n31333), .B1(n29600), .B2(n29599), .ZN(
        n29612) );
  NAND2_X1 U36872 ( .A1(n30037), .A2(n30051), .ZN(n29604) );
  INV_X1 U36873 ( .A(n29601), .ZN(n29603) );
  AND2_X1 U36874 ( .A1(n31346), .A2(n29602), .ZN(n31938) );
  AOI22_X1 U36875 ( .A1(n29604), .A2(n29603), .B1(n31938), .B2(n30053), .ZN(
        n29611) );
  INV_X1 U36876 ( .A(n29959), .ZN(n29605) );
  NAND2_X1 U36877 ( .A1(n30033), .A2(n29605), .ZN(n29610) );
  INV_X1 U36878 ( .A(n31933), .ZN(n29606) );
  AOI21_X1 U36879 ( .B1(n29606), .B2(n29609), .A(n31936), .ZN(n29608) );
  XNOR2_X1 U36880 ( .A(n34146), .B(n51664), .ZN(n29613) );
  XNOR2_X1 U36881 ( .A(n35517), .B(n29613), .ZN(n29614) );
  XNOR2_X1 U36882 ( .A(n29615), .B(n29614), .ZN(n38547) );
  NAND2_X1 U36883 ( .A1(n36148), .A2(n38547), .ZN(n38228) );
  OAI21_X1 U36884 ( .B1(n32986), .B2(n712), .A(n32981), .ZN(n29620) );
  OAI21_X1 U36885 ( .B1(n32983), .B2(n29618), .A(n29617), .ZN(n29619) );
  NOR2_X1 U36886 ( .A1(n29621), .A2(n32600), .ZN(n32598) );
  NAND2_X1 U36887 ( .A1(n32598), .A2(n29622), .ZN(n32589) );
  AND2_X1 U36888 ( .A1(n32491), .A2(n32478), .ZN(n31208) );
  INV_X1 U36889 ( .A(n31208), .ZN(n29623) );
  OAI21_X1 U36890 ( .B1(n32489), .B2(n32487), .A(n29623), .ZN(n29624) );
  INV_X1 U36892 ( .A(n32028), .ZN(n31006) );
  NAND2_X1 U36893 ( .A1(n29624), .A2(n31006), .ZN(n29632) );
  AND2_X1 U36894 ( .A1(n29627), .A2(n29626), .ZN(n29631) );
  INV_X1 U36895 ( .A(n32015), .ZN(n31204) );
  NAND2_X1 U36896 ( .A1(n32485), .A2(n32473), .ZN(n31201) );
  NAND2_X1 U36897 ( .A1(n31201), .A2(n32478), .ZN(n32476) );
  OAI21_X1 U36898 ( .B1(n32484), .B2(n32478), .A(n32476), .ZN(n29628) );
  NAND2_X1 U36899 ( .A1(n31204), .A2(n29628), .ZN(n29630) );
  INV_X1 U36900 ( .A(n32027), .ZN(n32479) );
  NOR2_X1 U36901 ( .A1(n32479), .A2(n32484), .ZN(n31206) );
  OAI21_X1 U36902 ( .B1(n32483), .B2(n32472), .A(n31206), .ZN(n29629) );
  NAND4_X2 U36903 ( .A1(n29632), .A2(n29630), .A3(n29631), .A4(n29629), .ZN(
        n34896) );
  XNOR2_X1 U36904 ( .A(n35124), .B(n34896), .ZN(n29640) );
  AND2_X1 U36905 ( .A1(n33005), .A2(n51740), .ZN(n31387) );
  AND2_X1 U36906 ( .A1(n31384), .A2(n720), .ZN(n33014) );
  NAND2_X1 U36907 ( .A1(n31387), .A2(n33014), .ZN(n30540) );
  AND2_X1 U36908 ( .A1(n30540), .A2(n33009), .ZN(n29639) );
  NAND3_X1 U36909 ( .A1(n33017), .A2(n31011), .A3(n3487), .ZN(n29634) );
  OAI21_X1 U36910 ( .B1(n31379), .B2(n51740), .A(n33005), .ZN(n29636) );
  NAND2_X1 U36911 ( .A1(n33004), .A2(n29636), .ZN(n29637) );
  XNOR2_X1 U36912 ( .A(n32644), .B(n4880), .ZN(n33439) );
  XNOR2_X1 U36913 ( .A(n29640), .B(n33439), .ZN(n29670) );
  NAND2_X1 U36914 ( .A1(n31058), .A2(n30931), .ZN(n31061) );
  AOI21_X1 U36915 ( .B1(n31061), .B2(n31509), .A(n30082), .ZN(n29649) );
  NOR2_X1 U36916 ( .A1(n29643), .A2(n30931), .ZN(n31054) );
  INV_X1 U36917 ( .A(n31054), .ZN(n29647) );
  NAND2_X1 U36918 ( .A1(n30931), .A2(n30930), .ZN(n30085) );
  INV_X1 U36919 ( .A(n30929), .ZN(n30092) );
  NAND2_X1 U36920 ( .A1(n29644), .A2(n30092), .ZN(n29646) );
  INV_X1 U36921 ( .A(n30924), .ZN(n31056) );
  NOR2_X1 U36922 ( .A1(n31056), .A2(n30931), .ZN(n31052) );
  INV_X1 U36923 ( .A(n31052), .ZN(n29645) );
  NAND2_X1 U36924 ( .A1(n30640), .A2(n30649), .ZN(n29651) );
  NOR2_X1 U36925 ( .A1(n31311), .A2(n51085), .ZN(n30643) );
  NOR2_X1 U36928 ( .A1(n31302), .A2(n31303), .ZN(n31315) );
  INV_X1 U36929 ( .A(n31315), .ZN(n29654) );
  INV_X1 U36930 ( .A(n31891), .ZN(n29655) );
  OR2_X1 U36931 ( .A1(n31141), .A2(n31425), .ZN(n31143) );
  INV_X1 U36932 ( .A(n31143), .ZN(n29656) );
  OAI21_X1 U36933 ( .B1(n29992), .B2(n725), .A(n29656), .ZN(n29659) );
  AND2_X1 U36934 ( .A1(n31422), .A2(n31425), .ZN(n31898) );
  INV_X1 U36935 ( .A(n29657), .ZN(n29984) );
  OAI21_X1 U36936 ( .B1(n29995), .B2(n31898), .A(n29984), .ZN(n29658) );
  INV_X1 U36937 ( .A(n29661), .ZN(n29666) );
  XNOR2_X1 U36938 ( .A(n29662), .B(n1326), .ZN(n29663) );
  XNOR2_X1 U36939 ( .A(n29664), .B(n29663), .ZN(n29665) );
  XNOR2_X1 U36940 ( .A(n29666), .B(n29665), .ZN(n29667) );
  XNOR2_X1 U36941 ( .A(n34156), .B(n29667), .ZN(n29668) );
  XNOR2_X1 U36942 ( .A(n36873), .B(n29668), .ZN(n29669) );
  XNOR2_X1 U36943 ( .A(n29670), .B(n29669), .ZN(n29824) );
  AND2_X1 U36944 ( .A1(n30879), .A2(n32503), .ZN(n30878) );
  OAI21_X1 U36945 ( .B1(n30881), .B2(n30882), .A(n31987), .ZN(n29671) );
  NOR2_X1 U36946 ( .A1(n30878), .A2(n29671), .ZN(n29681) );
  INV_X1 U36947 ( .A(n32506), .ZN(n29672) );
  NOR2_X1 U36948 ( .A1(n32509), .A2(n7897), .ZN(n31191) );
  AND2_X1 U36949 ( .A1(n31995), .A2(n32004), .ZN(n29673) );
  AOI22_X1 U36950 ( .A1(n29672), .A2(n31191), .B1(n707), .B2(n29673), .ZN(
        n29680) );
  INV_X1 U36951 ( .A(n29673), .ZN(n29674) );
  NAND3_X1 U36952 ( .A1(n31191), .A2(n29674), .A3(n30877), .ZN(n29679) );
  INV_X1 U36953 ( .A(n29675), .ZN(n29676) );
  OAI21_X1 U36954 ( .B1(n29677), .B2(n32503), .A(n29676), .ZN(n29678) );
  INV_X1 U36955 ( .A(n30591), .ZN(n29682) );
  OR2_X1 U36956 ( .A1(n29683), .A2(n29682), .ZN(n29689) );
  NOR3_X1 U36957 ( .A1(n31096), .A2(n29684), .A3(n30592), .ZN(n29685) );
  NAND2_X1 U36958 ( .A1(n31096), .A2(n30592), .ZN(n30910) );
  NAND3_X1 U36959 ( .A1(n29687), .A2(n30593), .A3(n30590), .ZN(n29688) );
  XNOR2_X1 U36960 ( .A(n36766), .B(n46062), .ZN(n29823) );
  OAI21_X1 U36961 ( .B1(n29872), .B2(n30436), .A(n29691), .ZN(n29696) );
  NAND3_X1 U36962 ( .A1(n29859), .A2(n51746), .A3(n29703), .ZN(n29693) );
  NAND2_X1 U36963 ( .A1(n29694), .A2(n29693), .ZN(n29695) );
  AOI21_X1 U36964 ( .B1(n29697), .B2(n29696), .A(n29695), .ZN(n29712) );
  MUX2_X1 U36965 ( .A(n29698), .B(n29703), .S(n51746), .Z(n29699) );
  NAND2_X1 U36966 ( .A1(n29699), .A2(n486), .ZN(n29701) );
  AOI22_X1 U36967 ( .A1(n29702), .A2(n29869), .B1(n29701), .B2(n29700), .ZN(
        n29711) );
  NOR2_X1 U36968 ( .A1(n29703), .A2(n30429), .ZN(n29705) );
  NOR2_X1 U36969 ( .A1(n30429), .A2(n6770), .ZN(n29704) );
  INV_X1 U36971 ( .A(n29862), .ZN(n29708) );
  AOI22_X1 U36972 ( .A1(n29873), .A2(n29708), .B1(n29707), .B2(n29706), .ZN(
        n29709) );
  INV_X1 U36973 ( .A(n29713), .ZN(n30415) );
  MUX2_X1 U36974 ( .A(n30415), .B(n29717), .S(n28187), .Z(n29726) );
  NAND2_X1 U36975 ( .A1(n30407), .A2(n51108), .ZN(n29720) );
  AOI21_X1 U36976 ( .B1(n29721), .B2(n29720), .A(n51342), .ZN(n29723) );
  OR2_X1 U36977 ( .A1(n29723), .A2(n29722), .ZN(n29725) );
  OAI21_X1 U36978 ( .B1(n29726), .B2(n29725), .A(n29724), .ZN(n29732) );
  NAND2_X1 U36979 ( .A1(n29728), .A2(n29727), .ZN(n29729) );
  OAI22_X1 U36980 ( .A1(n29729), .A2(n30401), .B1(n30419), .B2(n30407), .ZN(
        n29730) );
  INV_X1 U36981 ( .A(n29730), .ZN(n29731) );
  NAND2_X1 U36982 ( .A1(n29736), .A2(n427), .ZN(n29733) );
  NAND2_X1 U36983 ( .A1(n29747), .A2(n2143), .ZN(n29739) );
  NAND2_X1 U36984 ( .A1(n29736), .A2(n51692), .ZN(n29738) );
  NAND4_X1 U36985 ( .A1(n29739), .A2(n29738), .A3(n29749), .A4(n29737), .ZN(
        n29743) );
  INV_X1 U36986 ( .A(n29745), .ZN(n29746) );
  NAND2_X1 U36987 ( .A1(n29748), .A2(n29747), .ZN(n29751) );
  NAND3_X1 U36988 ( .A1(n8747), .A2(n30461), .A3(n29749), .ZN(n29750) );
  NAND2_X1 U36989 ( .A1(n30349), .A2(n29754), .ZN(n29755) );
  NAND2_X1 U36990 ( .A1(n29755), .A2(n28300), .ZN(n29756) );
  INV_X1 U36991 ( .A(n29758), .ZN(n29762) );
  INV_X1 U36992 ( .A(n28300), .ZN(n29759) );
  OAI22_X1 U36993 ( .A1(n29765), .A2(n29764), .B1(n29763), .B2(n30354), .ZN(
        n29766) );
  NAND3_X1 U36994 ( .A1(n29769), .A2(n30340), .A3(n29768), .ZN(n29772) );
  INV_X1 U36995 ( .A(n29770), .ZN(n29771) );
  INV_X1 U36996 ( .A(n32725), .ZN(n32458) );
  INV_X1 U36997 ( .A(n30733), .ZN(n30746) );
  INV_X1 U36998 ( .A(n29774), .ZN(n30370) );
  NAND2_X1 U36999 ( .A1(n30733), .A2(n30379), .ZN(n30369) );
  OAI211_X1 U37000 ( .C1(n30746), .C2(n30370), .A(n30734), .B(n30369), .ZN(
        n29778) );
  OAI211_X1 U37001 ( .C1(n29776), .C2(n29784), .A(n29775), .B(n1121), .ZN(
        n29777) );
  AND2_X1 U37002 ( .A1(n29778), .A2(n29777), .ZN(n29787) );
  NAND2_X1 U37003 ( .A1(n30375), .A2(n30370), .ZN(n30747) );
  INV_X1 U37004 ( .A(n30747), .ZN(n29779) );
  NAND2_X1 U37005 ( .A1(n1121), .A2(n30382), .ZN(n29884) );
  INV_X1 U37006 ( .A(n29780), .ZN(n29781) );
  NAND2_X1 U37007 ( .A1(n29781), .A2(n29880), .ZN(n30736) );
  OAI21_X1 U37008 ( .B1(n27379), .B2(n29782), .A(n30374), .ZN(n29783) );
  OAI211_X1 U37009 ( .C1(n742), .C2(n29784), .A(n29783), .B(n52181), .ZN(
        n30377) );
  INV_X1 U37010 ( .A(n30377), .ZN(n29785) );
  INV_X1 U37011 ( .A(n32716), .ZN(n32729) );
  NAND2_X1 U37012 ( .A1(n32458), .A2(n32729), .ZN(n29788) );
  NAND2_X1 U37013 ( .A1(n32714), .A2(n29788), .ZN(n29813) );
  INV_X1 U37014 ( .A(n5054), .ZN(n29795) );
  OAI21_X1 U37015 ( .B1(n29796), .B2(n29795), .A(n29794), .ZN(n29799) );
  NAND2_X1 U37016 ( .A1(n29799), .A2(n29798), .ZN(n29807) );
  OAI21_X1 U37017 ( .B1(n29802), .B2(n29801), .A(n29800), .ZN(n29805) );
  NAND3_X1 U37018 ( .A1(n29805), .A2(n29804), .A3(n5057), .ZN(n29806) );
  NAND3_X2 U37019 ( .A1(n8738), .A2(n29807), .A3(n29806), .ZN(n32719) );
  AND2_X1 U37020 ( .A1(n32724), .A2(n32732), .ZN(n32312) );
  OAI21_X1 U37021 ( .B1(n32318), .B2(n32312), .A(n31644), .ZN(n29812) );
  XNOR2_X1 U37022 ( .A(n32719), .B(n32463), .ZN(n29808) );
  NAND2_X1 U37023 ( .A1(n29808), .A2(n32724), .ZN(n29809) );
  AOI21_X1 U37025 ( .B1(n32731), .B2(n29809), .A(n32464), .ZN(n29811) );
  NAND2_X1 U37026 ( .A1(n32716), .A2(n32719), .ZN(n31969) );
  NOR2_X1 U37027 ( .A1(n31969), .A2(n32732), .ZN(n31646) );
  NAND2_X1 U37028 ( .A1(n31646), .A2(n32725), .ZN(n29810) );
  NAND2_X1 U37030 ( .A1(n29814), .A2(n30140), .ZN(n32692) );
  OR2_X1 U37031 ( .A1(n32684), .A2(n31658), .ZN(n32706) );
  AOI22_X1 U37034 ( .A1(n29816), .A2(n32706), .B1(n30144), .B2(n30140), .ZN(
        n29822) );
  NAND2_X1 U37035 ( .A1(n32684), .A2(n32324), .ZN(n29817) );
  NAND4_X1 U37036 ( .A1(n29817), .A2(n30140), .A3(n32327), .A4(n32705), .ZN(
        n29818) );
  NAND2_X1 U37037 ( .A1(n31658), .A2(n32684), .ZN(n32700) );
  AND2_X1 U37038 ( .A1(n32700), .A2(n29818), .ZN(n29821) );
  NAND2_X1 U37039 ( .A1(n30144), .A2(n32327), .ZN(n32687) );
  INV_X1 U37040 ( .A(n32335), .ZN(n29819) );
  OAI21_X1 U37041 ( .B1(n29819), .B2(n32325), .A(n32333), .ZN(n29820) );
  XNOR2_X1 U37043 ( .A(n29823), .B(n460), .ZN(n35772) );
  XNOR2_X1 U37044 ( .A(n35772), .B(n29824), .ZN(n29983) );
  INV_X1 U37046 ( .A(n33159), .ZN(n29825) );
  OAI21_X1 U37047 ( .B1(n31950), .B2(n31290), .A(n32081), .ZN(n33162) );
  NAND3_X1 U37048 ( .A1(n7430), .A2(n32071), .A3(n32407), .ZN(n33152) );
  NAND2_X1 U37050 ( .A1(n33154), .A2(n33155), .ZN(n29826) );
  NAND2_X1 U37051 ( .A1(n31580), .A2(n30854), .ZN(n29827) );
  INV_X1 U37052 ( .A(n30856), .ZN(n31577) );
  NAND2_X1 U37053 ( .A1(n51545), .A2(n30856), .ZN(n31629) );
  INV_X1 U37054 ( .A(n30549), .ZN(n29828) );
  NAND2_X1 U37055 ( .A1(n30898), .A2(n29829), .ZN(n29832) );
  INV_X1 U37056 ( .A(n29830), .ZN(n29831) );
  NAND2_X1 U37057 ( .A1(n29832), .A2(n29831), .ZN(n29836) );
  NAND3_X1 U37058 ( .A1(n32114), .A2(n32104), .A3(n32089), .ZN(n29835) );
  OAI211_X1 U37059 ( .C1(n30904), .C2(n32560), .A(n32561), .B(n32087), .ZN(
        n29833) );
  NOR2_X1 U37060 ( .A1(n854), .A2(n32105), .ZN(n32571) );
  NAND2_X1 U37061 ( .A1(n29833), .A2(n32571), .ZN(n29834) );
  NAND2_X1 U37062 ( .A1(n32088), .A2(n32107), .ZN(n32568) );
  XNOR2_X1 U37064 ( .A(n35133), .B(n36999), .ZN(n29949) );
  NAND2_X1 U37065 ( .A1(n31489), .A2(n31484), .ZN(n30109) );
  INV_X1 U37066 ( .A(n30106), .ZN(n30994) );
  NOR2_X1 U37067 ( .A1(n30102), .A2(n31496), .ZN(n30097) );
  INV_X1 U37068 ( .A(n29837), .ZN(n31499) );
  NAND2_X1 U37069 ( .A1(n30097), .A2(n31499), .ZN(n29838) );
  OAI211_X1 U37070 ( .C1(n30109), .C2(n30994), .A(n31266), .B(n29838), .ZN(
        n29839) );
  INV_X1 U37071 ( .A(n29839), .ZN(n29847) );
  NOR2_X1 U37072 ( .A1(n31497), .A2(n1472), .ZN(n31483) );
  INV_X1 U37073 ( .A(n30109), .ZN(n31498) );
  NAND2_X1 U37074 ( .A1(n31483), .A2(n31498), .ZN(n29845) );
  NAND3_X1 U37075 ( .A1(n3224), .A2(n29841), .A3(n31489), .ZN(n29842) );
  NAND2_X1 U37076 ( .A1(n29842), .A2(n30102), .ZN(n29843) );
  NAND2_X1 U37077 ( .A1(n29843), .A2(n31497), .ZN(n29844) );
  NOR2_X1 U37078 ( .A1(n29848), .A2(n30716), .ZN(n29849) );
  OAI21_X1 U37079 ( .B1(n29850), .B2(n29849), .A(n29853), .ZN(n29858) );
  NOR2_X1 U37080 ( .A1(n30705), .A2(n29851), .ZN(n29852) );
  AOI22_X1 U37081 ( .A1(n29852), .A2(n30709), .B1(n30721), .B2(n2205), .ZN(
        n29857) );
  AOI21_X1 U37082 ( .B1(n29853), .B2(n30721), .A(n30706), .ZN(n29854) );
  NAND3_X1 U37083 ( .A1(n30719), .A2(n29855), .A3(n30712), .ZN(n29856) );
  NAND2_X1 U37084 ( .A1(n29859), .A2(n30434), .ZN(n29860) );
  AND3_X1 U37085 ( .A1(n29862), .A2(n29861), .A3(n29860), .ZN(n29879) );
  INV_X1 U37086 ( .A(n30429), .ZN(n29865) );
  AOI22_X1 U37087 ( .A1(n29875), .A2(n29865), .B1(n728), .B2(n29864), .ZN(
        n29878) );
  INV_X1 U37088 ( .A(n29866), .ZN(n29871) );
  NOR2_X1 U37089 ( .A1(n29868), .A2(n29867), .ZN(n29870) );
  OAI21_X1 U37090 ( .B1(n29871), .B2(n29870), .A(n29869), .ZN(n29877) );
  NOR2_X1 U37091 ( .A1(n29872), .A2(n30434), .ZN(n29874) );
  OAI21_X1 U37092 ( .B1(n29875), .B2(n29874), .A(n29873), .ZN(n29876) );
  INV_X1 U37093 ( .A(n30375), .ZN(n30737) );
  AOI21_X1 U37094 ( .B1(n30364), .B2(n30379), .A(n30380), .ZN(n29891) );
  AND3_X1 U37095 ( .A1(n30382), .A2(n30379), .A3(n29883), .ZN(n29885) );
  OAI211_X1 U37096 ( .C1(n30731), .C2(n29885), .A(n30740), .B(n29884), .ZN(
        n29889) );
  OAI21_X1 U37097 ( .B1(n29887), .B2(n29886), .A(n30375), .ZN(n29888) );
  INV_X1 U37098 ( .A(n32438), .ZN(n31320) );
  NAND2_X1 U37099 ( .A1(n29892), .A2(n29905), .ZN(n29894) );
  AOI21_X1 U37100 ( .B1(n29895), .B2(n29894), .A(n29893), .ZN(n29898) );
  NOR2_X1 U37101 ( .A1(n29898), .A2(n29897), .ZN(n29914) );
  OAI222_X1 U37102 ( .A1(n30785), .A2(n30783), .B1(n29901), .B2(n29900), .C1(
        n29899), .C2(n30794), .ZN(n29903) );
  AOI22_X1 U37103 ( .A1(n29904), .A2(n30791), .B1(n29903), .B2(n29902), .ZN(
        n29913) );
  XNOR2_X1 U37104 ( .A(n30785), .B(n29905), .ZN(n29906) );
  INV_X1 U37105 ( .A(n29907), .ZN(n30782) );
  OAI21_X1 U37106 ( .B1(n29910), .B2(n30792), .A(n29909), .ZN(n29911) );
  NAND2_X1 U37107 ( .A1(n31320), .A2(n32439), .ZN(n32436) );
  NAND2_X1 U37108 ( .A1(n32056), .A2(n32439), .ZN(n32352) );
  AND2_X1 U37109 ( .A1(n29920), .A2(n29919), .ZN(n29929) );
  NAND2_X1 U37110 ( .A1(n29922), .A2(n29921), .ZN(n30777) );
  NOR2_X1 U37111 ( .A1(n29924), .A2(n8377), .ZN(n29925) );
  OAI21_X1 U37112 ( .B1(n51696), .B2(n29925), .A(n30758), .ZN(n29927) );
  NAND2_X1 U37113 ( .A1(n30768), .A2(n30771), .ZN(n30760) );
  NOR2_X1 U37114 ( .A1(n30760), .A2(n738), .ZN(n29926) );
  OR2_X1 U37115 ( .A1(n29931), .A2(n402), .ZN(n30682) );
  OAI211_X1 U37117 ( .C1(n30687), .C2(n29933), .A(n29932), .B(n30389), .ZN(
        n29934) );
  OAI211_X1 U37118 ( .C1(n30682), .C2(n29936), .A(n29935), .B(n29934), .ZN(
        n29937) );
  INV_X1 U37119 ( .A(n29937), .ZN(n29947) );
  NOR2_X1 U37120 ( .A1(n29938), .A2(n24091), .ZN(n29939) );
  AOI22_X1 U37121 ( .A1(n30690), .A2(n29939), .B1(n30392), .B2(n30688), .ZN(
        n29946) );
  MUX2_X1 U37122 ( .A(n29940), .B(n30683), .S(n30696), .Z(n29941) );
  NAND2_X1 U37123 ( .A1(n29941), .A2(n30394), .ZN(n29945) );
  NAND2_X1 U37124 ( .A1(n29942), .A2(n30690), .ZN(n29944) );
  INV_X1 U37125 ( .A(n32051), .ZN(n31326) );
  AND2_X1 U37126 ( .A1(n32356), .A2(n32439), .ZN(n31323) );
  NOR2_X1 U37127 ( .A1(n31955), .A2(n32056), .ZN(n32455) );
  NAND2_X1 U37128 ( .A1(n32345), .A2(n32438), .ZN(n32044) );
  NOR2_X1 U37129 ( .A1(n32044), .A2(n718), .ZN(n31321) );
  NAND2_X1 U37130 ( .A1(n31321), .A2(n32351), .ZN(n29948) );
  XNOR2_X1 U37131 ( .A(n29949), .B(n52221), .ZN(n35486) );
  INV_X1 U37132 ( .A(n31121), .ZN(n29952) );
  OAI21_X1 U37133 ( .B1(n29950), .B2(n31106), .A(n30941), .ZN(n29951) );
  OAI211_X1 U37134 ( .C1(n29952), .C2(n30073), .A(n29951), .B(n623), .ZN(
        n29957) );
  INV_X1 U37135 ( .A(n29953), .ZN(n31123) );
  INV_X1 U37136 ( .A(n31105), .ZN(n29954) );
  OAI21_X1 U37137 ( .B1(n30943), .B2(n29954), .A(n30070), .ZN(n29956) );
  NAND2_X1 U37138 ( .A1(n30072), .A2(n31111), .ZN(n29955) );
  NOR2_X1 U37139 ( .A1(n31931), .A2(n31346), .ZN(n29958) );
  NOR2_X1 U37140 ( .A1(n2354), .A2(n29958), .ZN(n29965) );
  NOR2_X1 U37141 ( .A1(n30051), .A2(n51744), .ZN(n30038) );
  OAI21_X1 U37142 ( .B1(n2906), .B2(n31938), .A(n30038), .ZN(n29964) );
  OAI21_X1 U37143 ( .B1(n30038), .B2(n30037), .A(n29959), .ZN(n31331) );
  NAND2_X1 U37144 ( .A1(n30053), .A2(n31338), .ZN(n30029) );
  INV_X1 U37145 ( .A(n30029), .ZN(n29960) );
  NAND2_X1 U37146 ( .A1(n31331), .A2(n29960), .ZN(n29963) );
  NAND2_X1 U37147 ( .A1(n31938), .A2(n31338), .ZN(n29961) );
  NAND4_X1 U37148 ( .A1(n31339), .A2(n30053), .A3(n29961), .A4(n5682), .ZN(
        n29962) );
  AOI21_X1 U37149 ( .B1(n2098), .B2(n51240), .A(n31690), .ZN(n29971) );
  INV_X1 U37150 ( .A(n29967), .ZN(n29968) );
  OAI211_X1 U37151 ( .C1(n708), .C2(n29968), .A(n31676), .B(n2098), .ZN(n29970) );
  INV_X1 U37152 ( .A(n30974), .ZN(n31687) );
  OAI21_X1 U37153 ( .B1(n31682), .B2(n31687), .A(n30013), .ZN(n29969) );
  INV_X1 U37154 ( .A(n29973), .ZN(n29974) );
  AND2_X1 U37155 ( .A1(n32125), .A2(n32130), .ZN(n30818) );
  OAI21_X1 U37156 ( .B1(n30818), .B2(n32119), .A(n32131), .ZN(n29980) );
  NAND3_X1 U37157 ( .A1(n29976), .A2(n29975), .A3(n31699), .ZN(n29977) );
  OAI21_X1 U37158 ( .B1(n31701), .B2(n32128), .A(n29977), .ZN(n29979) );
  AND2_X1 U37159 ( .A1(n31708), .A2(n32130), .ZN(n31710) );
  NAND2_X1 U37160 ( .A1(n31701), .A2(n31710), .ZN(n29978) );
  XNOR2_X1 U37162 ( .A(n35283), .B(n35678), .ZN(n35128) );
  XNOR2_X1 U37163 ( .A(n35128), .B(n35486), .ZN(n29982) );
  MUX2_X1 U37164 ( .A(n38228), .B(n36148), .S(n38558), .Z(n31353) );
  NOR2_X1 U37165 ( .A1(n31425), .A2(n31422), .ZN(n31149) );
  OAI211_X1 U37166 ( .C1(n31149), .C2(n31899), .A(n29984), .B(n31151), .ZN(
        n29987) );
  NAND4_X1 U37167 ( .A1(n29985), .A2(n31146), .A3(n31413), .A4(n725), .ZN(
        n29986) );
  NAND2_X1 U37168 ( .A1(n29987), .A2(n29986), .ZN(n29988) );
  INV_X1 U37169 ( .A(n29990), .ZN(n31895) );
  NAND3_X1 U37170 ( .A1(n31895), .A2(n31898), .A3(n31892), .ZN(n29997) );
  OAI21_X1 U37171 ( .B1(n29991), .B2(n31425), .A(n31413), .ZN(n29993) );
  INV_X1 U37172 ( .A(n31690), .ZN(n30002) );
  OAI211_X1 U37173 ( .C1(n30007), .C2(n31680), .A(n31691), .B(n29998), .ZN(
        n30001) );
  INV_X1 U37174 ( .A(n29999), .ZN(n30000) );
  OAI211_X1 U37175 ( .C1(n31684), .C2(n30002), .A(n30001), .B(n30000), .ZN(
        n30011) );
  INV_X1 U37176 ( .A(n30003), .ZN(n30005) );
  OAI21_X1 U37177 ( .B1(n30005), .B2(n30004), .A(n31687), .ZN(n30009) );
  NAND2_X1 U37178 ( .A1(n30009), .A2(n30008), .ZN(n30010) );
  NOR2_X1 U37179 ( .A1(n30011), .A2(n30010), .ZN(n30028) );
  NOR2_X1 U37180 ( .A1(n30016), .A2(n30014), .ZN(n30020) );
  INV_X1 U37181 ( .A(n30015), .ZN(n30019) );
  NOR2_X1 U37182 ( .A1(n30975), .A2(n30016), .ZN(n30018) );
  INV_X1 U37183 ( .A(n30978), .ZN(n30017) );
  AOI22_X1 U37184 ( .A1(n30020), .A2(n30019), .B1(n30018), .B2(n30017), .ZN(
        n30026) );
  INV_X1 U37185 ( .A(n30979), .ZN(n30021) );
  NAND2_X1 U37186 ( .A1(n30024), .A2(n30023), .ZN(n30025) );
  XNOR2_X1 U37187 ( .A(n51739), .B(n33218), .ZN(n30078) );
  NOR2_X1 U37188 ( .A1(n30030), .A2(n30029), .ZN(n31344) );
  INV_X1 U37189 ( .A(n30031), .ZN(n30032) );
  OAI21_X1 U37190 ( .B1(n30054), .B2(n31333), .A(n30032), .ZN(n30042) );
  INV_X1 U37191 ( .A(n30034), .ZN(n30035) );
  NOR2_X1 U37192 ( .A1(n30036), .A2(n30035), .ZN(n30041) );
  NAND3_X1 U37193 ( .A1(n30038), .A2(n30053), .A3(n30037), .ZN(n30039) );
  NAND3_X1 U37194 ( .A1(n31935), .A2(n31346), .A3(n30039), .ZN(n30040) );
  OAI22_X1 U37195 ( .A1(n31344), .A2(n30042), .B1(n30041), .B2(n30040), .ZN(
        n30056) );
  XNOR2_X1 U37196 ( .A(n30051), .B(n51744), .ZN(n30046) );
  AND2_X1 U37197 ( .A1(n31340), .A2(n31934), .ZN(n30045) );
  NAND2_X1 U37198 ( .A1(n31346), .A2(n31338), .ZN(n30044) );
  NAND4_X1 U37199 ( .A1(n30046), .A2(n31931), .A3(n30045), .A4(n30044), .ZN(
        n30049) );
  AOI21_X1 U37200 ( .B1(n30052), .B2(n30051), .A(n30050), .ZN(n30055) );
  NOR2_X1 U37201 ( .A1(n51744), .A2(n31934), .ZN(n31336) );
  INV_X1 U37202 ( .A(n30057), .ZN(n30063) );
  NAND2_X1 U37204 ( .A1(n30073), .A2(n30058), .ZN(n30060) );
  NOR2_X1 U37205 ( .A1(n31106), .A2(n362), .ZN(n30059) );
  NAND4_X1 U37206 ( .A1(n30060), .A2(n30947), .A3(n30059), .A4(n52121), .ZN(
        n30061) );
  AND3_X1 U37207 ( .A1(n30062), .A2(n30944), .A3(n30061), .ZN(n30068) );
  MUX2_X1 U37208 ( .A(n30063), .B(n30946), .S(n31116), .Z(n30064) );
  INV_X1 U37209 ( .A(n30064), .ZN(n30067) );
  NAND4_X1 U37210 ( .A1(n31117), .A2(n30073), .A3(n30058), .A4(n623), .ZN(
        n30065) );
  INV_X1 U37211 ( .A(n30943), .ZN(n31104) );
  INV_X1 U37212 ( .A(n30941), .ZN(n30069) );
  NAND2_X1 U37213 ( .A1(n31106), .A2(n7658), .ZN(n30949) );
  NOR2_X2 U37216 ( .A1(n30077), .A2(n30076), .ZN(n35334) );
  XNOR2_X1 U37217 ( .A(n37108), .B(n35334), .ZN(n33983) );
  XNOR2_X1 U37218 ( .A(n33983), .B(n30078), .ZN(n30116) );
  INV_X1 U37219 ( .A(n30082), .ZN(n31518) );
  OAI211_X1 U37220 ( .C1(n31055), .C2(n31067), .A(n31051), .B(n30931), .ZN(
        n30089) );
  NAND2_X1 U37221 ( .A1(n31058), .A2(n31513), .ZN(n31523) );
  NAND2_X1 U37222 ( .A1(n30936), .A2(n31510), .ZN(n30084) );
  AND4_X1 U37223 ( .A1(n31523), .A2(n30084), .A3(n30927), .A4(n30083), .ZN(
        n30088) );
  INV_X1 U37224 ( .A(n30085), .ZN(n30086) );
  NAND3_X1 U37225 ( .A1(n30086), .A2(n30929), .A3(n31512), .ZN(n30087) );
  INV_X1 U37226 ( .A(n30091), .ZN(n31066) );
  NAND2_X1 U37228 ( .A1(n30936), .A2(n30925), .ZN(n30093) );
  MUX2_X1 U37229 ( .A(n30094), .B(n30093), .S(n30935), .Z(n30095) );
  INV_X1 U37230 ( .A(n30097), .ZN(n30099) );
  OAI211_X1 U37231 ( .C1(n30109), .C2(n30099), .A(n30098), .B(n31488), .ZN(
        n30101) );
  NAND2_X1 U37232 ( .A1(n31481), .A2(n31497), .ZN(n30100) );
  NAND2_X1 U37233 ( .A1(n30101), .A2(n30100), .ZN(n30115) );
  AND2_X1 U37234 ( .A1(n31496), .A2(n31490), .ZN(n31264) );
  INV_X1 U37235 ( .A(n31264), .ZN(n31487) );
  NOR2_X1 U37236 ( .A1(n31496), .A2(n31490), .ZN(n31502) );
  AND2_X1 U37237 ( .A1(n31496), .A2(n31489), .ZN(n30996) );
  OAI21_X1 U37238 ( .B1(n30996), .B2(n30104), .A(n31488), .ZN(n30105) );
  NAND3_X1 U37239 ( .A1(n30106), .A2(n31497), .A3(n31490), .ZN(n30108) );
  AND3_X1 U37240 ( .A1(n30993), .A2(n30108), .A3(n30107), .ZN(n30113) );
  XNOR2_X1 U37241 ( .A(n3224), .B(n31497), .ZN(n30111) );
  NAND4_X1 U37242 ( .A1(n30111), .A2(n31490), .A3(n30110), .A4(n30109), .ZN(
        n30112) );
  XNOR2_X1 U37243 ( .A(n30116), .B(n2168), .ZN(n31966) );
  INV_X1 U37244 ( .A(n30118), .ZN(n31021) );
  OAI211_X1 U37245 ( .C1(n31800), .C2(n30120), .A(n31801), .B(n51479), .ZN(
        n30123) );
  NAND3_X1 U37246 ( .A1(n31874), .A2(n31799), .A3(n30121), .ZN(n30122) );
  NAND3_X1 U37247 ( .A1(n31799), .A2(n51479), .A3(n52047), .ZN(n30128) );
  NAND2_X1 U37248 ( .A1(n30125), .A2(n31803), .ZN(n30126) );
  OAI211_X1 U37249 ( .C1(n31882), .C2(n30128), .A(n30127), .B(n30126), .ZN(
        n30129) );
  NOR2_X1 U37250 ( .A1(n30130), .A2(n30129), .ZN(n30131) );
  OR2_X1 U37251 ( .A1(n52182), .A2(n32684), .ZN(n32328) );
  NAND2_X1 U37252 ( .A1(n32333), .A2(n52182), .ZN(n30135) );
  NAND2_X1 U37253 ( .A1(n32684), .A2(n32327), .ZN(n30133) );
  NAND2_X1 U37254 ( .A1(n30133), .A2(n30140), .ZN(n30134) );
  NAND4_X1 U37255 ( .A1(n32328), .A2(n32324), .A3(n30135), .A4(n30134), .ZN(
        n30139) );
  INV_X1 U37256 ( .A(n30136), .ZN(n30138) );
  OR2_X1 U37257 ( .A1(n32700), .A2(n32705), .ZN(n30137) );
  AND3_X1 U37258 ( .A1(n30138), .A2(n30139), .A3(n30137), .ZN(n30158) );
  NOR2_X1 U37259 ( .A1(n32684), .A2(n32691), .ZN(n32708) );
  NOR2_X1 U37260 ( .A1(n32684), .A2(n32705), .ZN(n30142) );
  NAND2_X1 U37261 ( .A1(n52301), .A2(n30140), .ZN(n30152) );
  OAI211_X1 U37262 ( .C1(n32708), .C2(n30142), .A(n30141), .B(n30152), .ZN(
        n30146) );
  AND2_X1 U37263 ( .A1(n30145), .A2(n30146), .ZN(n30157) );
  OR2_X1 U37264 ( .A1(n32684), .A2(n32327), .ZN(n32690) );
  NAND2_X1 U37265 ( .A1(n32690), .A2(n32332), .ZN(n30154) );
  INV_X1 U37266 ( .A(n30154), .ZN(n30151) );
  INV_X1 U37267 ( .A(n30147), .ZN(n30149) );
  INV_X1 U37268 ( .A(n32331), .ZN(n30148) );
  NOR2_X1 U37269 ( .A1(n30149), .A2(n30148), .ZN(n30150) );
  NAND2_X1 U37270 ( .A1(n30151), .A2(n30150), .ZN(n30156) );
  INV_X1 U37271 ( .A(n30152), .ZN(n30153) );
  NAND3_X1 U37272 ( .A1(n30154), .A2(n30153), .A3(n32324), .ZN(n30155) );
  NOR2_X1 U37273 ( .A1(n30159), .A2(n2201), .ZN(n30162) );
  INV_X1 U37274 ( .A(n30160), .ZN(n30161) );
  NAND2_X1 U37275 ( .A1(n30164), .A2(n30163), .ZN(n30311) );
  NAND3_X1 U37276 ( .A1(n30167), .A2(n30165), .A3(n30314), .ZN(n30166) );
  AND3_X1 U37277 ( .A1(n30317), .A2(n30311), .A3(n30166), .ZN(n30190) );
  XNOR2_X1 U37278 ( .A(n30167), .B(n30181), .ZN(n30170) );
  AND2_X1 U37279 ( .A1(n30168), .A2(n30183), .ZN(n30169) );
  NAND2_X1 U37281 ( .A1(n30175), .A2(n30178), .ZN(n30319) );
  OAI21_X1 U37282 ( .B1(n6084), .B2(n30178), .A(n30181), .ZN(n30187) );
  NAND2_X1 U37283 ( .A1(n30181), .A2(n2201), .ZN(n30185) );
  OAI21_X1 U37284 ( .B1(n30183), .B2(n30182), .A(n25199), .ZN(n30184) );
  NAND4_X1 U37285 ( .A1(n30187), .A2(n30186), .A3(n30185), .A4(n30184), .ZN(
        n30188) );
  AND2_X1 U37286 ( .A1(n30310), .A2(n30188), .ZN(n30189) );
  NAND2_X1 U37287 ( .A1(n30197), .A2(n30191), .ZN(n30196) );
  NAND2_X1 U37288 ( .A1(n30193), .A2(n30192), .ZN(n30195) );
  MUX2_X1 U37289 ( .A(n30196), .B(n30195), .S(n30194), .Z(n30205) );
  INV_X1 U37290 ( .A(n30197), .ZN(n30198) );
  OAI211_X1 U37291 ( .C1(n30203), .C2(n30202), .A(n30201), .B(n30200), .ZN(
        n30204) );
  AND2_X1 U37292 ( .A1(n30205), .A2(n30204), .ZN(n30217) );
  NAND3_X1 U37293 ( .A1(n30211), .A2(n30210), .A3(n30209), .ZN(n30212) );
  NAND2_X1 U37294 ( .A1(n30213), .A2(n30212), .ZN(n30214) );
  NAND2_X1 U37295 ( .A1(n30214), .A2(n1871), .ZN(n30215) );
  NAND2_X1 U37296 ( .A1(n30222), .A2(n30221), .ZN(n30239) );
  AND3_X1 U37297 ( .A1(n30224), .A2(n30225), .A3(n30223), .ZN(n30238) );
  NAND3_X1 U37298 ( .A1(n30228), .A2(n30227), .A3(n30226), .ZN(n30229) );
  AND2_X1 U37299 ( .A1(n30230), .A2(n30229), .ZN(n30237) );
  NAND2_X1 U37300 ( .A1(n30242), .A2(n52165), .ZN(n30255) );
  INV_X1 U37301 ( .A(n30243), .ZN(n30246) );
  OAI21_X1 U37302 ( .B1(n30246), .B2(n30245), .A(n5417), .ZN(n30254) );
  OAI21_X1 U37303 ( .B1(n30249), .B2(n52165), .A(n626), .ZN(n30250) );
  NAND2_X1 U37304 ( .A1(n30251), .A2(n30250), .ZN(n30252) );
  AND2_X1 U37305 ( .A1(n32608), .A2(n31558), .ZN(n31158) );
  NOR2_X1 U37306 ( .A1(n51106), .A2(n32608), .ZN(n31564) );
  INV_X1 U37307 ( .A(n30257), .ZN(n30261) );
  NAND2_X1 U37308 ( .A1(n30258), .A2(n25075), .ZN(n30260) );
  NAND3_X1 U37309 ( .A1(n52195), .A2(n2158), .A3(n52102), .ZN(n30259) );
  OAI22_X1 U37311 ( .A1(n25418), .A2(n52195), .B1(n30263), .B2(n25107), .ZN(
        n30266) );
  MUX2_X1 U37313 ( .A(n30269), .B(n30268), .S(n30267), .Z(n30271) );
  NAND2_X1 U37314 ( .A1(n30271), .A2(n30270), .ZN(n30276) );
  INV_X1 U37315 ( .A(n30272), .ZN(n30274) );
  NAND2_X1 U37316 ( .A1(n30274), .A2(n52147), .ZN(n30275) );
  NAND3_X1 U37318 ( .A1(n30281), .A2(n30280), .A3(n30279), .ZN(n30288) );
  AOI21_X1 U37319 ( .B1(n2881), .B2(n30283), .A(n30282), .ZN(n30287) );
  NAND2_X1 U37320 ( .A1(n51748), .A2(n30285), .ZN(n30286) );
  NAND2_X1 U37321 ( .A1(n30290), .A2(n30289), .ZN(n30300) );
  OAI21_X1 U37322 ( .B1(n30292), .B2(n2110), .A(n30291), .ZN(n30294) );
  NAND2_X1 U37323 ( .A1(n30294), .A2(n30293), .ZN(n30298) );
  NAND3_X1 U37324 ( .A1(n51748), .A2(n30296), .A3(n30295), .ZN(n30297) );
  INV_X1 U37325 ( .A(n30302), .ZN(n30321) );
  NAND3_X1 U37326 ( .A1(n30304), .A2(n30303), .A3(n1771), .ZN(n30309) );
  NAND3_X1 U37327 ( .A1(n30307), .A2(n30306), .A3(n30305), .ZN(n30308) );
  AND3_X1 U37328 ( .A1(n30310), .A2(n30309), .A3(n30308), .ZN(n30318) );
  OAI21_X1 U37329 ( .B1(n30313), .B2(n30312), .A(n30311), .ZN(n30315) );
  NAND2_X1 U37330 ( .A1(n30315), .A2(n30314), .ZN(n30316) );
  NAND4_X1 U37331 ( .A1(n30319), .A2(n30318), .A3(n30317), .A4(n30316), .ZN(
        n30320) );
  OAI21_X1 U37332 ( .B1(n30321), .B2(n30320), .A(n31558), .ZN(n31462) );
  AND2_X1 U37336 ( .A1(n30323), .A2(n30324), .ZN(n30335) );
  INV_X1 U37337 ( .A(n31462), .ZN(n31470) );
  NOR3_X1 U37338 ( .A1(n32608), .A2(n32616), .A3(n31558), .ZN(n30326) );
  NAND2_X1 U37339 ( .A1(n32609), .A2(n31466), .ZN(n32610) );
  INV_X1 U37340 ( .A(n32610), .ZN(n30325) );
  OAI21_X1 U37341 ( .B1(n31470), .B2(n30326), .A(n30325), .ZN(n30329) );
  AND4_X1 U37342 ( .A1(n32620), .A2(n31466), .A3(n7626), .A4(n7625), .ZN(
        n30327) );
  AND2_X1 U37343 ( .A1(n31466), .A2(n31558), .ZN(n31461) );
  AOI22_X1 U37344 ( .A1(n30327), .A2(n51106), .B1(n31461), .B2(n32608), .ZN(
        n30328) );
  AND3_X1 U37345 ( .A1(n30328), .A2(n30329), .A3(n31160), .ZN(n30334) );
  NAND2_X1 U37346 ( .A1(n51106), .A2(n32608), .ZN(n31161) );
  INV_X1 U37347 ( .A(n31161), .ZN(n30332) );
  NAND2_X1 U37348 ( .A1(n30330), .A2(n32616), .ZN(n30331) );
  OAI211_X1 U37349 ( .C1(n30332), .C2(n31566), .A(n30331), .B(n31159), .ZN(
        n30333) );
  XNOR2_X1 U37350 ( .A(n34760), .B(n35070), .ZN(n30337) );
  OAI22_X1 U37351 ( .A1(n30339), .A2(n28300), .B1(n30349), .B2(n30338), .ZN(
        n30341) );
  NAND2_X1 U37352 ( .A1(n30341), .A2(n30340), .ZN(n30359) );
  AND2_X1 U37353 ( .A1(n51489), .A2(n7721), .ZN(n30347) );
  NAND2_X1 U37354 ( .A1(n30347), .A2(n514), .ZN(n30353) );
  NAND2_X1 U37355 ( .A1(n30347), .A2(n30346), .ZN(n30352) );
  NAND2_X1 U37356 ( .A1(n30349), .A2(n30348), .ZN(n30350) );
  NAND4_X1 U37357 ( .A1(n30353), .A2(n30352), .A3(n30351), .A4(n30350), .ZN(
        n30357) );
  AOI22_X1 U37358 ( .A1(n29063), .A2(n5389), .B1(n30355), .B2(n30354), .ZN(
        n30356) );
  NAND4_X2 U37359 ( .A1(n30359), .A2(n30358), .A3(n30357), .A4(n30356), .ZN(
        n31401) );
  MUX2_X1 U37360 ( .A(n30733), .B(n30360), .S(n30382), .Z(n30362) );
  AOI21_X1 U37361 ( .B1(n30362), .B2(n1121), .A(n30361), .ZN(n30363) );
  AOI21_X1 U37362 ( .B1(n30365), .B2(n30364), .A(n30363), .ZN(n30373) );
  INV_X1 U37363 ( .A(n30366), .ZN(n30368) );
  NAND2_X1 U37364 ( .A1(n30733), .A2(n30370), .ZN(n30367) );
  NAND3_X1 U37365 ( .A1(n30734), .A2(n30370), .A3(n30369), .ZN(n30371) );
  NAND2_X1 U37366 ( .A1(n30375), .A2(n30374), .ZN(n30378) );
  MUX2_X1 U37367 ( .A(n30381), .B(n30380), .S(n30379), .Z(n30383) );
  NAND3_X1 U37368 ( .A1(n30384), .A2(n30687), .A3(n30389), .ZN(n30385) );
  AND2_X1 U37369 ( .A1(n30389), .A2(n24091), .ZN(n30390) );
  AND2_X1 U37370 ( .A1(n30683), .A2(n51113), .ZN(n30695) );
  NOR2_X1 U37371 ( .A1(n30692), .A2(n30393), .ZN(n30395) );
  NOR2_X1 U37372 ( .A1(n30401), .A2(n30419), .ZN(n30402) );
  NAND2_X1 U37373 ( .A1(n30402), .A2(n28793), .ZN(n30410) );
  NAND2_X1 U37374 ( .A1(n30406), .A2(n30405), .ZN(n30408) );
  NAND2_X1 U37375 ( .A1(n30408), .A2(n30407), .ZN(n30409) );
  NAND2_X1 U37376 ( .A1(n30412), .A2(n30411), .ZN(n30414) );
  AOI21_X1 U37377 ( .B1(n30415), .B2(n30414), .A(n30413), .ZN(n30423) );
  NAND2_X1 U37378 ( .A1(n30417), .A2(n30416), .ZN(n30422) );
  INV_X1 U37379 ( .A(n31401), .ZN(n32821) );
  OAI21_X1 U37380 ( .B1(n31401), .B2(n32823), .A(n32415), .ZN(n30470) );
  AND2_X1 U37381 ( .A1(n486), .A2(n30425), .ZN(n30435) );
  OAI22_X1 U37382 ( .A1(n30435), .A2(n30434), .B1(n30433), .B2(n51746), .ZN(
        n30438) );
  INV_X1 U37383 ( .A(n32428), .ZN(n30440) );
  AND2_X1 U37384 ( .A1(n32424), .A2(n30440), .ZN(n30469) );
  INV_X1 U37385 ( .A(n30441), .ZN(n30443) );
  NOR2_X1 U37386 ( .A1(n30443), .A2(n427), .ZN(n30445) );
  OAI21_X1 U37387 ( .B1(n30446), .B2(n30445), .A(n30444), .ZN(n30468) );
  OAI21_X1 U37388 ( .B1(n30449), .B2(n30448), .A(n30447), .ZN(n30450) );
  INV_X1 U37389 ( .A(n30450), .ZN(n30467) );
  AND2_X1 U37391 ( .A1(n30453), .A2(n30454), .ZN(n30466) );
  NOR2_X1 U37392 ( .A1(n30461), .A2(n51693), .ZN(n30456) );
  OAI21_X1 U37393 ( .B1(n2143), .B2(n30458), .A(n28521), .ZN(n30460) );
  AOI21_X1 U37394 ( .B1(n30462), .B2(n30461), .A(n30460), .ZN(n30463) );
  INV_X1 U37396 ( .A(n32828), .ZN(n32421) );
  NOR2_X1 U37397 ( .A1(n32420), .A2(n31401), .ZN(n30471) );
  NAND2_X1 U37398 ( .A1(n32421), .A2(n30471), .ZN(n31258) );
  INV_X1 U37401 ( .A(n32825), .ZN(n31404) );
  AOI21_X1 U37402 ( .B1(n30473), .B2(n32428), .A(n31398), .ZN(n30475) );
  OAI211_X1 U37403 ( .C1(n31404), .C2(n32429), .A(n30475), .B(n30474), .ZN(
        n30476) );
  OAI21_X1 U37404 ( .B1(n32829), .B2(n30477), .A(n30476), .ZN(n30480) );
  NAND2_X1 U37405 ( .A1(n51618), .A2(n31398), .ZN(n31249) );
  INV_X1 U37406 ( .A(n31249), .ZN(n30478) );
  NAND3_X1 U37407 ( .A1(n31397), .A2(n32821), .A3(n30478), .ZN(n30479) );
  NOR2_X1 U37408 ( .A1(n31075), .A2(n32386), .ZN(n30481) );
  INV_X1 U37409 ( .A(n32850), .ZN(n30496) );
  MUX2_X1 U37410 ( .A(n30481), .B(n30496), .S(n32841), .Z(n30489) );
  AOI21_X1 U37411 ( .B1(n32379), .B2(n32386), .A(n31911), .ZN(n30482) );
  OAI21_X1 U37412 ( .B1(n30482), .B2(n32841), .A(n31914), .ZN(n30488) );
  INV_X1 U37413 ( .A(n30483), .ZN(n30486) );
  XNOR2_X1 U37414 ( .A(n30484), .B(n31910), .ZN(n30485) );
  OAI21_X1 U37415 ( .B1(n30486), .B2(n30485), .A(n31911), .ZN(n30487) );
  OAI211_X1 U37416 ( .C1(n30489), .C2(n31914), .A(n30488), .B(n30487), .ZN(
        n30494) );
  NOR2_X1 U37417 ( .A1(n32389), .A2(n32381), .ZN(n30490) );
  NOR2_X1 U37418 ( .A1(n31920), .A2(n30490), .ZN(n30493) );
  NAND4_X1 U37419 ( .A1(n30494), .A2(n30493), .A3(n30492), .A4(n30491), .ZN(
        n30500) );
  NOR2_X1 U37420 ( .A1(n32852), .A2(n32385), .ZN(n31083) );
  INV_X1 U37421 ( .A(n31083), .ZN(n30498) );
  AOI21_X1 U37422 ( .B1(n30498), .B2(n30497), .A(n30496), .ZN(n30499) );
  XNOR2_X1 U37423 ( .A(n30501), .B(n37111), .ZN(n33851) );
  XNOR2_X1 U37424 ( .A(n31966), .B(n33851), .ZN(n30810) );
  NOR2_X1 U37425 ( .A1(n32988), .A2(n2984), .ZN(n32975) );
  AND3_X1 U37426 ( .A1(n32980), .A2(n30505), .A3(n30504), .ZN(n30524) );
  INV_X1 U37427 ( .A(n30506), .ZN(n30507) );
  NAND3_X1 U37428 ( .A1(n32983), .A2(n30507), .A3(n32974), .ZN(n30509) );
  AND2_X1 U37429 ( .A1(n30509), .A2(n30508), .ZN(n30523) );
  NAND2_X1 U37430 ( .A1(n32988), .A2(n32590), .ZN(n30511) );
  NAND2_X1 U37431 ( .A1(n30511), .A2(n30510), .ZN(n30514) );
  NAND2_X1 U37432 ( .A1(n32988), .A2(n712), .ZN(n30512) );
  OAI22_X1 U37433 ( .A1(n32989), .A2(n30514), .B1(n30513), .B2(n30512), .ZN(
        n30515) );
  NAND2_X1 U37434 ( .A1(n30515), .A2(n32990), .ZN(n30522) );
  NAND2_X1 U37435 ( .A1(n30518), .A2(n32586), .ZN(n30520) );
  NAND2_X1 U37436 ( .A1(n30520), .A2(n30519), .ZN(n30521) );
  XNOR2_X1 U37437 ( .A(n30526), .B(n30525), .ZN(n30527) );
  XNOR2_X1 U37438 ( .A(n32860), .B(n30527), .ZN(n30569) );
  NOR2_X1 U37440 ( .A1(n33002), .A2(n33005), .ZN(n33008) );
  INV_X1 U37441 ( .A(n30528), .ZN(n30537) );
  NAND4_X1 U37442 ( .A1(n33008), .A2(n33017), .A3(n30537), .A4(n30543), .ZN(
        n30530) );
  OAI211_X1 U37443 ( .C1(n31384), .C2(n30531), .A(n30530), .B(n30529), .ZN(
        n30532) );
  INV_X1 U37444 ( .A(n30532), .ZN(n30548) );
  INV_X1 U37445 ( .A(n30533), .ZN(n30536) );
  AND4_X1 U37446 ( .A1(n33002), .A2(n3241), .A3(n33005), .A4(n30534), .ZN(
        n30535) );
  OAI21_X1 U37447 ( .B1(n30536), .B2(n30535), .A(n33017), .ZN(n30547) );
  NOR2_X1 U37448 ( .A1(n33019), .A2(n33017), .ZN(n30541) );
  NAND4_X1 U37450 ( .A1(n30541), .A2(n30540), .A3(n30539), .A4(n30538), .ZN(
        n30546) );
  NAND2_X1 U37451 ( .A1(n30542), .A2(n31385), .ZN(n31014) );
  INV_X1 U37452 ( .A(n31014), .ZN(n33003) );
  INV_X1 U37453 ( .A(n30543), .ZN(n31388) );
  AND4_X1 U37454 ( .A1(n33017), .A2(n31388), .A3(n33014), .A4(n33005), .ZN(
        n30544) );
  NOR2_X1 U37455 ( .A1(n33003), .A2(n30544), .ZN(n30545) );
  AOI21_X1 U37457 ( .B1(n51545), .B2(n30855), .A(n31624), .ZN(n30552) );
  INV_X1 U37458 ( .A(n31580), .ZN(n30551) );
  OR2_X1 U37459 ( .A1(n30552), .A2(n30551), .ZN(n30556) );
  INV_X1 U37460 ( .A(n31639), .ZN(n30553) );
  INV_X1 U37461 ( .A(n30558), .ZN(n31576) );
  OAI211_X1 U37462 ( .C1(n30553), .C2(n31576), .A(n31586), .B(n31625), .ZN(
        n30555) );
  OAI211_X1 U37463 ( .C1(n30559), .C2(n31631), .A(n31632), .B(n30853), .ZN(
        n30554) );
  NAND4_X1 U37464 ( .A1(n30557), .A2(n30556), .A3(n30555), .A4(n30554), .ZN(
        n30568) );
  NAND2_X1 U37465 ( .A1(n30558), .A2(n30854), .ZN(n30560) );
  NAND4_X1 U37466 ( .A1(n30560), .A2(n30559), .A3(n30855), .A4(n30861), .ZN(
        n30566) );
  AND2_X1 U37467 ( .A1(n31631), .A2(n30856), .ZN(n30562) );
  NAND2_X1 U37468 ( .A1(n30853), .A2(n31624), .ZN(n30561) );
  OAI211_X1 U37469 ( .C1(n51545), .C2(n30855), .A(n30562), .B(n30561), .ZN(
        n30565) );
  AND2_X1 U37470 ( .A1(n30853), .A2(n31638), .ZN(n30563) );
  NAND4_X1 U37471 ( .A1(n31586), .A2(n30563), .A3(n30854), .A4(n30856), .ZN(
        n30564) );
  NAND3_X1 U37472 ( .A1(n30566), .A2(n30565), .A3(n30564), .ZN(n30567) );
  XNOR2_X1 U37473 ( .A(n30569), .B(n33085), .ZN(n30618) );
  INV_X1 U37474 ( .A(n31029), .ZN(n30570) );
  AND2_X1 U37475 ( .A1(n31821), .A2(n30846), .ZN(n30848) );
  NOR3_X1 U37476 ( .A1(n30572), .A2(n30571), .A3(n31816), .ZN(n30574) );
  NAND2_X1 U37477 ( .A1(n31816), .A2(n31039), .ZN(n31822) );
  AND2_X1 U37478 ( .A1(n50986), .A2(n31815), .ZN(n31829) );
  NOR2_X1 U37479 ( .A1(n30574), .A2(n30573), .ZN(n30588) );
  NOR2_X1 U37480 ( .A1(n30577), .A2(n31816), .ZN(n30578) );
  AOI22_X1 U37481 ( .A1(n31830), .A2(n30579), .B1(n30578), .B2(n31038), .ZN(
        n30587) );
  INV_X1 U37483 ( .A(n31827), .ZN(n30850) );
  OAI21_X1 U37484 ( .B1(n31033), .B2(n30846), .A(n31816), .ZN(n30583) );
  NAND4_X1 U37485 ( .A1(n2486), .A2(n30585), .A3(n30584), .A4(n30583), .ZN(
        n30586) );
  XNOR2_X1 U37486 ( .A(n2204), .B(n4487), .ZN(n30617) );
  MUX2_X1 U37487 ( .A(n30918), .B(n30590), .S(n31087), .Z(n30616) );
  AND2_X1 U37488 ( .A1(n30592), .A2(n30593), .ZN(n30913) );
  NAND3_X1 U37489 ( .A1(n30913), .A2(n30599), .A3(n31086), .ZN(n30596) );
  AOI21_X1 U37490 ( .B1(n31087), .B2(n30599), .A(n30609), .ZN(n30606) );
  OAI21_X1 U37491 ( .B1(n31088), .B2(n30601), .A(n30600), .ZN(n30604) );
  NOR2_X1 U37492 ( .A1(n30607), .A2(n30602), .ZN(n30603) );
  NAND2_X1 U37493 ( .A1(n30608), .A2(n30607), .ZN(n30612) );
  INV_X1 U37494 ( .A(n30609), .ZN(n30610) );
  NAND2_X1 U37495 ( .A1(n31093), .A2(n30610), .ZN(n30611) );
  MUX2_X1 U37496 ( .A(n30612), .B(n30611), .S(n31086), .Z(n30613) );
  XNOR2_X1 U37497 ( .A(n30617), .B(n37113), .ZN(n35627) );
  XNOR2_X1 U37498 ( .A(n30618), .B(n35627), .ZN(n30808) );
  INV_X1 U37499 ( .A(n32302), .ZN(n30629) );
  INV_X1 U37500 ( .A(n30619), .ZN(n30621) );
  INV_X1 U37501 ( .A(n30623), .ZN(n30620) );
  NAND2_X1 U37502 ( .A1(n30621), .A2(n30620), .ZN(n30625) );
  OR2_X1 U37503 ( .A1(n30623), .A2(n30622), .ZN(n30624) );
  NAND2_X1 U37504 ( .A1(n7383), .A2(n31749), .ZN(n30630) );
  INV_X1 U37505 ( .A(n30630), .ZN(n30626) );
  NAND4_X1 U37506 ( .A1(n30635), .A2(n30626), .A3(n31369), .A4(n31366), .ZN(
        n30628) );
  OAI21_X1 U37508 ( .B1(n31849), .B2(n711), .A(n31742), .ZN(n30627) );
  NAND3_X1 U37509 ( .A1(n711), .A2(n7383), .A3(n31746), .ZN(n32301) );
  OAI21_X1 U37510 ( .B1(n31743), .B2(n31369), .A(n32301), .ZN(n30631) );
  NAND3_X1 U37511 ( .A1(n30631), .A2(n31740), .A3(n30630), .ZN(n30638) );
  INV_X1 U37512 ( .A(n30632), .ZN(n31368) );
  NOR2_X1 U37514 ( .A1(n4299), .A2(n31740), .ZN(n30633) );
  OR2_X1 U37516 ( .A1(n32295), .A2(n31749), .ZN(n30634) );
  OAI211_X1 U37517 ( .C1(n32301), .C2(n386), .A(n32297), .B(n30634), .ZN(
        n30637) );
  NAND2_X1 U37518 ( .A1(n32299), .A2(n386), .ZN(n31744) );
  INV_X1 U37519 ( .A(n31312), .ZN(n30639) );
  OAI211_X1 U37520 ( .C1(n31294), .C2(n30824), .A(n30639), .B(n30647), .ZN(
        n30641) );
  INV_X1 U37521 ( .A(n30643), .ZN(n30831) );
  NAND2_X1 U37522 ( .A1(n51086), .A2(n30644), .ZN(n30645) );
  NAND2_X1 U37523 ( .A1(n30645), .A2(n31303), .ZN(n30646) );
  AND2_X1 U37524 ( .A1(n31302), .A2(n51086), .ZN(n30650) );
  AND2_X1 U37525 ( .A1(n31301), .A2(n31300), .ZN(n30651) );
  AOI22_X1 U37526 ( .A1(n30650), .A2(n30651), .B1(n30649), .B2(n51085), .ZN(
        n30656) );
  INV_X1 U37527 ( .A(n30653), .ZN(n30654) );
  NAND4_X1 U37528 ( .A1(n30654), .A2(n30825), .A3(n4607), .A4(n51085), .ZN(
        n30655) );
  INV_X1 U37529 ( .A(n30657), .ZN(n30660) );
  OAI21_X1 U37530 ( .B1(n30660), .B2(n30659), .A(n30658), .ZN(n30681) );
  OAI21_X1 U37531 ( .B1(n30663), .B2(n30662), .A(n30661), .ZN(n30666) );
  NAND3_X1 U37532 ( .A1(n30666), .A2(n30665), .A3(n30664), .ZN(n30675) );
  NAND2_X1 U37533 ( .A1(n23859), .A2(n30667), .ZN(n30668) );
  OAI211_X1 U37534 ( .C1(n30671), .C2(n30670), .A(n30669), .B(n30668), .ZN(
        n30674) );
  NAND4_X1 U37535 ( .A1(n30675), .A2(n30674), .A3(n30673), .A4(n30672), .ZN(
        n30679) );
  INV_X1 U37536 ( .A(n30682), .ZN(n30686) );
  NOR2_X1 U37537 ( .A1(n30694), .A2(n30683), .ZN(n30684) );
  AOI21_X1 U37538 ( .B1(n30686), .B2(n30685), .A(n30684), .ZN(n30704) );
  MUX2_X1 U37539 ( .A(n51257), .B(n30688), .S(n30687), .Z(n30691) );
  NAND2_X1 U37540 ( .A1(n30691), .A2(n30690), .ZN(n30703) );
  NAND2_X1 U37541 ( .A1(n24091), .A2(n30692), .ZN(n30693) );
  NAND2_X1 U37542 ( .A1(n30697), .A2(n30696), .ZN(n30702) );
  NAND2_X1 U37543 ( .A1(n30700), .A2(n28758), .ZN(n30701) );
  NOR2_X1 U37544 ( .A1(n31452), .A2(n32665), .ZN(n31447) );
  OAI21_X1 U37545 ( .B1(n30707), .B2(n30706), .A(n30705), .ZN(n30708) );
  AND2_X1 U37546 ( .A1(n30711), .A2(n30712), .ZN(n30714) );
  AOI21_X1 U37547 ( .B1(n30715), .B2(n30714), .A(n30713), .ZN(n30729) );
  NAND2_X1 U37548 ( .A1(n30722), .A2(n2205), .ZN(n30720) );
  OAI22_X1 U37549 ( .A1(n30724), .A2(n30723), .B1(n30722), .B2(n30721), .ZN(
        n30726) );
  NAND2_X1 U37550 ( .A1(n30726), .A2(n30725), .ZN(n30727) );
  AOI21_X1 U37554 ( .B1(n30748), .B2(n30747), .A(n30746), .ZN(n30749) );
  NOR2_X1 U37555 ( .A1(n30759), .A2(n30758), .ZN(n30762) );
  INV_X1 U37556 ( .A(n30760), .ZN(n30761) );
  NAND3_X1 U37557 ( .A1(n30764), .A2(n738), .A3(n30763), .ZN(n30765) );
  OAI21_X1 U37558 ( .B1(n30770), .B2(n30769), .A(n30768), .ZN(n30775) );
  NOR2_X1 U37559 ( .A1(n30772), .A2(n30771), .ZN(n30774) );
  OAI21_X1 U37560 ( .B1(n30775), .B2(n30774), .A(n30773), .ZN(n30776) );
  NAND3_X1 U37561 ( .A1(n30778), .A2(n30777), .A3(n30776), .ZN(n30779) );
  MUX2_X1 U37562 ( .A(n31540), .B(n31450), .S(n31169), .Z(n30801) );
  NOR2_X1 U37563 ( .A1(n30782), .A2(n30781), .ZN(n30787) );
  NOR2_X1 U37564 ( .A1(n23658), .A2(n30792), .ZN(n30784) );
  NAND2_X1 U37565 ( .A1(n30789), .A2(n30788), .ZN(n30797) );
  NOR2_X1 U37566 ( .A1(n30791), .A2(n30790), .ZN(n30793) );
  NAND3_X1 U37567 ( .A1(n27570), .A2(n30795), .A3(n30794), .ZN(n30796) );
  NOR2_X1 U37568 ( .A1(n31454), .A2(n31452), .ZN(n30805) );
  AOI21_X1 U37569 ( .B1(n382), .B2(n32665), .A(n31538), .ZN(n30799) );
  NAND2_X1 U37570 ( .A1(n31452), .A2(n32665), .ZN(n30962) );
  INV_X1 U37571 ( .A(n30962), .ZN(n32662) );
  NOR2_X1 U37572 ( .A1(n31454), .A2(n31546), .ZN(n31539) );
  NAND3_X1 U37573 ( .A1(n31539), .A2(n31538), .A3(n32665), .ZN(n30804) );
  NAND2_X1 U37574 ( .A1(n32663), .A2(n30962), .ZN(n30803) );
  MUX2_X1 U37575 ( .A(n30804), .B(n30803), .S(n381), .Z(n30807) );
  NAND2_X1 U37576 ( .A1(n31539), .A2(n31538), .ZN(n30967) );
  INV_X1 U37578 ( .A(n30805), .ZN(n31536) );
  NAND2_X1 U37579 ( .A1(n382), .A2(n31452), .ZN(n32666) );
  XNOR2_X1 U37581 ( .A(n35065), .B(n35237), .ZN(n34263) );
  XNOR2_X1 U37582 ( .A(n34263), .B(n30808), .ZN(n30809) );
  INV_X1 U37583 ( .A(n30811), .ZN(n32126) );
  INV_X1 U37584 ( .A(n31709), .ZN(n30812) );
  INV_X1 U37585 ( .A(n31699), .ZN(n32137) );
  NAND4_X1 U37586 ( .A1(n31706), .A2(n32137), .A3(n32125), .A4(n31711), .ZN(
        n30813) );
  NAND2_X1 U37587 ( .A1(n31706), .A2(n32118), .ZN(n30815) );
  INV_X1 U37588 ( .A(n32120), .ZN(n31714) );
  OAI21_X1 U37589 ( .B1(n30818), .B2(n30815), .A(n31714), .ZN(n30819) );
  INV_X1 U37590 ( .A(n30816), .ZN(n30817) );
  NAND2_X1 U37591 ( .A1(n30818), .A2(n30817), .ZN(n32135) );
  NOR2_X1 U37592 ( .A1(n30820), .A2(n32909), .ZN(n30821) );
  AND2_X1 U37593 ( .A1(n32895), .A2(n32916), .ZN(n32548) );
  INV_X1 U37594 ( .A(n32917), .ZN(n32901) );
  NAND4_X1 U37595 ( .A1(n32548), .A2(n32915), .A3(n32894), .A4(n32901), .ZN(
        n30823) );
  NOR2_X1 U37596 ( .A1(n31312), .A2(n30824), .ZN(n30827) );
  NAND2_X1 U37597 ( .A1(n31294), .A2(n31306), .ZN(n30832) );
  INV_X1 U37598 ( .A(n30825), .ZN(n30826) );
  AOI22_X1 U37599 ( .A1(n31313), .A2(n30827), .B1(n30832), .B2(n30826), .ZN(
        n30838) );
  OAI211_X1 U37600 ( .C1(n30834), .C2(n30833), .A(n30832), .B(n30831), .ZN(
        n30836) );
  NAND2_X1 U37601 ( .A1(n30836), .A2(n30835), .ZN(n30837) );
  AOI22_X1 U37602 ( .A1(n32225), .A2(n32226), .B1(n32253), .B2(n32251), .ZN(
        n30844) );
  NAND2_X1 U37603 ( .A1(n32252), .A2(n32254), .ZN(n30840) );
  NAND2_X1 U37604 ( .A1(n30840), .A2(n32230), .ZN(n30841) );
  NAND2_X1 U37605 ( .A1(n30841), .A2(n31238), .ZN(n30843) );
  OR2_X1 U37607 ( .A1(n32243), .A2(n32252), .ZN(n31779) );
  OAI211_X1 U37608 ( .C1(n32231), .C2(n31781), .A(n31779), .B(n31240), .ZN(
        n30842) );
  AND2_X1 U37609 ( .A1(n31816), .A2(n30846), .ZN(n31820) );
  INV_X1 U37610 ( .A(n31829), .ZN(n30847) );
  NOR2_X1 U37611 ( .A1(n31630), .A2(n30853), .ZN(n30859) );
  NOR2_X1 U37612 ( .A1(n31583), .A2(n30855), .ZN(n30858) );
  AOI22_X1 U37613 ( .A1(n30859), .A2(n30858), .B1(n30857), .B2(n30856), .ZN(
        n30865) );
  INV_X1 U37614 ( .A(n31636), .ZN(n31585) );
  NAND2_X1 U37615 ( .A1(n30860), .A2(n31585), .ZN(n30863) );
  NAND2_X1 U37616 ( .A1(n31636), .A2(n30861), .ZN(n31641) );
  NAND2_X1 U37617 ( .A1(n31641), .A2(n31640), .ZN(n30862) );
  INV_X1 U37618 ( .A(n31466), .ZN(n31557) );
  AOI21_X1 U37619 ( .B1(n31557), .B2(n32608), .A(n51471), .ZN(n30866) );
  NAND2_X1 U37620 ( .A1(n51471), .A2(n31466), .ZN(n31565) );
  NOR2_X1 U37621 ( .A1(n31565), .A2(n32609), .ZN(n31563) );
  NAND3_X1 U37622 ( .A1(n31564), .A2(n31563), .A3(n31558), .ZN(n30870) );
  NAND2_X1 U37623 ( .A1(n31557), .A2(n32616), .ZN(n30868) );
  OR2_X1 U37624 ( .A1(n32617), .A2(n30868), .ZN(n30869) );
  NAND3_X1 U37625 ( .A1(n30872), .A2(n7897), .A3(n30877), .ZN(n30876) );
  AND2_X1 U37629 ( .A1(n30876), .A2(n32003), .ZN(n30885) );
  NAND2_X1 U37630 ( .A1(n30878), .A2(n8722), .ZN(n30884) );
  INV_X1 U37631 ( .A(n32500), .ZN(n32009) );
  INV_X1 U37632 ( .A(n30879), .ZN(n30880) );
  OAI211_X1 U37633 ( .C1(n32009), .C2(n31995), .A(n30880), .B(n51105), .ZN(
        n30883) );
  XNOR2_X1 U37634 ( .A(n32310), .B(n35345), .ZN(n35804) );
  XNOR2_X1 U37635 ( .A(n35804), .B(n36983), .ZN(n30886) );
  XNOR2_X1 U37636 ( .A(n30887), .B(n30886), .ZN(n30959) );
  NAND2_X1 U37637 ( .A1(n31764), .A2(n30893), .ZN(n30890) );
  INV_X1 U37638 ( .A(n30888), .ZN(n31770) );
  NAND2_X1 U37640 ( .A1(n30891), .A2(n32194), .ZN(n30897) );
  INV_X1 U37641 ( .A(n30892), .ZN(n31225) );
  AOI21_X1 U37642 ( .B1(n5109), .B2(n32194), .A(n50981), .ZN(n30895) );
  INV_X1 U37643 ( .A(n32197), .ZN(n30894) );
  AOI22_X1 U37644 ( .A1(n31225), .A2(n30895), .B1(n30894), .B2(n30893), .ZN(
        n30896) );
  INV_X1 U37645 ( .A(n32207), .ZN(n32193) );
  INV_X1 U37646 ( .A(n32114), .ZN(n31609) );
  INV_X1 U37647 ( .A(n32087), .ZN(n32102) );
  INV_X1 U37648 ( .A(n30898), .ZN(n30899) );
  AOI22_X1 U37649 ( .A1(n31609), .A2(n32102), .B1(n30899), .B2(n30901), .ZN(
        n32557) );
  OR2_X1 U37650 ( .A1(n32107), .A2(n32574), .ZN(n32095) );
  NOR2_X1 U37651 ( .A1(n32095), .A2(n32561), .ZN(n30903) );
  NOR2_X1 U37652 ( .A1(n30900), .A2(n32105), .ZN(n31607) );
  NOR2_X1 U37653 ( .A1(n32106), .A2(n32566), .ZN(n30902) );
  AOI22_X1 U37654 ( .A1(n30903), .A2(n31607), .B1(n30902), .B2(n30901), .ZN(
        n30908) );
  OAI211_X1 U37655 ( .C1(n624), .C2(n32566), .A(n32105), .B(n32089), .ZN(
        n30906) );
  INV_X1 U37656 ( .A(n30904), .ZN(n30905) );
  MUX2_X1 U37657 ( .A(n30906), .B(n30905), .S(n32561), .Z(n30907) );
  AND3_X1 U37658 ( .A1(n32557), .A2(n30908), .A3(n30907), .ZN(n33097) );
  AOI22_X1 U37659 ( .A1(n30914), .A2(n31093), .B1(n30913), .B2(n30912), .ZN(
        n30922) );
  INV_X1 U37660 ( .A(n30915), .ZN(n30917) );
  OAI21_X1 U37661 ( .B1(n30917), .B2(n31086), .A(n30916), .ZN(n30921) );
  INV_X1 U37662 ( .A(n30918), .ZN(n30919) );
  NAND3_X1 U37663 ( .A1(n30919), .A2(n31087), .A3(n31094), .ZN(n30920) );
  NAND2_X1 U37664 ( .A1(n30925), .A2(n30924), .ZN(n30928) );
  NAND4_X1 U37665 ( .A1(n30928), .A2(n31517), .A3(n3099), .A4(n31512), .ZN(
        n30926) );
  INV_X1 U37666 ( .A(n31061), .ZN(n30933) );
  NAND2_X1 U37667 ( .A1(n30929), .A2(n30928), .ZN(n30932) );
  OR2_X1 U37668 ( .A1(n30931), .A2(n30930), .ZN(n30934) );
  OAI21_X1 U37669 ( .B1(n30933), .B2(n30932), .A(n30934), .ZN(n30938) );
  NAND3_X1 U37671 ( .A1(n30936), .A2(n31519), .A3(n30935), .ZN(n30937) );
  XNOR2_X1 U37672 ( .A(n32337), .B(n31923), .ZN(n33226) );
  OAI211_X1 U37673 ( .C1(n31122), .C2(n30943), .A(n30942), .B(n30941), .ZN(
        n30945) );
  NAND2_X1 U37675 ( .A1(n30946), .A2(n31117), .ZN(n30951) );
  INV_X1 U37676 ( .A(n30947), .ZN(n30948) );
  NAND2_X1 U37677 ( .A1(n30949), .A2(n30948), .ZN(n30950) );
  AOI21_X1 U37678 ( .B1(n30951), .B2(n30950), .A(n31116), .ZN(n30952) );
  XNOR2_X1 U37679 ( .A(n30953), .B(n4589), .ZN(n30954) );
  XNOR2_X1 U37680 ( .A(n44220), .B(n30954), .ZN(n30955) );
  XNOR2_X1 U37681 ( .A(n35536), .B(n30955), .ZN(n30956) );
  XNOR2_X1 U37682 ( .A(n33226), .B(n30956), .ZN(n30957) );
  XNOR2_X1 U37683 ( .A(n34051), .B(n30957), .ZN(n30958) );
  XNOR2_X1 U37684 ( .A(n30959), .B(n30958), .ZN(n31018) );
  NAND2_X1 U37685 ( .A1(n31454), .A2(n31452), .ZN(n31541) );
  NOR2_X1 U37686 ( .A1(n31546), .A2(n31544), .ZN(n30960) );
  AND2_X1 U37687 ( .A1(n31541), .A2(n30960), .ZN(n30961) );
  OAI21_X1 U37688 ( .B1(n31168), .B2(n30961), .A(n382), .ZN(n30966) );
  NAND3_X1 U37689 ( .A1(n31166), .A2(n31541), .A3(n30962), .ZN(n30963) );
  OAI21_X1 U37690 ( .B1(n30964), .B2(n30963), .A(n31549), .ZN(n30965) );
  XNOR2_X1 U37691 ( .A(n2129), .B(n2183), .ZN(n32280) );
  OAI21_X1 U37693 ( .B1(n30975), .B2(n708), .A(n30974), .ZN(n30977) );
  NAND2_X1 U37694 ( .A1(n30980), .A2(n30979), .ZN(n30988) );
  OAI21_X1 U37695 ( .B1(n30982), .B2(n31680), .A(n30981), .ZN(n30985) );
  NAND3_X1 U37696 ( .A1(n30985), .A2(n51240), .A3(n30983), .ZN(n30987) );
  NAND2_X1 U37697 ( .A1(n31687), .A2(n30004), .ZN(n30986) );
  XNOR2_X1 U37698 ( .A(n34446), .B(n32280), .ZN(n31017) );
  INV_X1 U37699 ( .A(n30990), .ZN(n30991) );
  INV_X1 U37700 ( .A(n30999), .ZN(n30995) );
  OAI21_X1 U37701 ( .B1(n30995), .B2(n30994), .A(n30993), .ZN(n31275) );
  NAND3_X1 U37702 ( .A1(n30999), .A2(n31484), .A3(n30998), .ZN(n31000) );
  OAI21_X1 U37703 ( .B1(n32472), .B2(n32485), .A(n32027), .ZN(n31207) );
  NAND2_X1 U37704 ( .A1(n31208), .A2(n31207), .ZN(n31009) );
  NOR2_X1 U37705 ( .A1(n32486), .A2(n32484), .ZN(n31209) );
  NAND2_X1 U37706 ( .A1(n32478), .A2(n32025), .ZN(n31005) );
  NAND3_X1 U37707 ( .A1(n32491), .A2(n31209), .A3(n31005), .ZN(n31004) );
  INV_X1 U37708 ( .A(n31005), .ZN(n31007) );
  OAI21_X1 U37709 ( .B1(n31007), .B2(n31006), .A(n32479), .ZN(n31008) );
  XNOR2_X1 U37710 ( .A(n35085), .B(n35088), .ZN(n31015) );
  INV_X1 U37712 ( .A(n31011), .ZN(n31013) );
  XNOR2_X1 U37713 ( .A(n31015), .B(n35086), .ZN(n31016) );
  XNOR2_X1 U37714 ( .A(n31017), .B(n31016), .ZN(n36788) );
  OR2_X1 U37715 ( .A1(n31020), .A2(n31799), .ZN(n31023) );
  NAND2_X1 U37716 ( .A1(n31021), .A2(n31792), .ZN(n31022) );
  AND2_X1 U37717 ( .A1(n52047), .A2(n31870), .ZN(n31025) );
  NAND2_X1 U37719 ( .A1(n31029), .A2(n31827), .ZN(n31032) );
  NAND3_X1 U37720 ( .A1(n31034), .A2(n31033), .A3(n31829), .ZN(n31035) );
  AND2_X1 U37721 ( .A1(n31036), .A2(n31035), .ZN(n31048) );
  NOR2_X1 U37722 ( .A1(n31821), .A2(n50986), .ZN(n31037) );
  OAI21_X1 U37723 ( .B1(n31038), .B2(n31037), .A(n31820), .ZN(n31047) );
  OAI21_X1 U37724 ( .B1(n31041), .B2(n50986), .A(n31039), .ZN(n31045) );
  NAND2_X1 U37725 ( .A1(n31045), .A2(n31044), .ZN(n31046) );
  INV_X1 U37726 ( .A(n31050), .ZN(n31053) );
  OAI21_X1 U37727 ( .B1(n31053), .B2(n31052), .A(n31051), .ZN(n31064) );
  NAND2_X1 U37728 ( .A1(n31054), .A2(n31513), .ZN(n31522) );
  OAI21_X1 U37729 ( .B1(n31057), .B2(n31056), .A(n31517), .ZN(n31060) );
  NAND2_X1 U37730 ( .A1(n31058), .A2(n31067), .ZN(n31059) );
  NAND4_X1 U37731 ( .A1(n31062), .A2(n31061), .A3(n31060), .A4(n31059), .ZN(
        n31063) );
  AND3_X1 U37732 ( .A1(n31064), .A2(n31522), .A3(n31063), .ZN(n31072) );
  OAI21_X1 U37733 ( .B1(n31068), .B2(n31067), .A(n31066), .ZN(n31069) );
  NAND2_X1 U37735 ( .A1(n32841), .A2(n32386), .ZN(n31073) );
  INV_X1 U37736 ( .A(n31078), .ZN(n32838) );
  NAND2_X1 U37738 ( .A1(n32846), .A2(n32851), .ZN(n31077) );
  INV_X1 U37739 ( .A(n32377), .ZN(n31074) );
  AOI21_X1 U37740 ( .B1(n31075), .B2(n32843), .A(n31074), .ZN(n31076) );
  NAND2_X1 U37741 ( .A1(n31077), .A2(n31076), .ZN(n31081) );
  NAND2_X1 U37742 ( .A1(n32843), .A2(n31911), .ZN(n32378) );
  AOI21_X1 U37743 ( .B1(n32378), .B2(n31078), .A(n32389), .ZN(n31079) );
  NOR2_X1 U37744 ( .A1(n31079), .A2(n31920), .ZN(n31080) );
  MUX2_X1 U37745 ( .A(n31081), .B(n31080), .S(n713), .Z(n31085) );
  NAND3_X1 U37746 ( .A1(n31914), .A2(n713), .A3(n32838), .ZN(n32373) );
  AND2_X1 U37747 ( .A1(n32850), .A2(n32843), .ZN(n31082) );
  NAND2_X1 U37748 ( .A1(n31083), .A2(n32389), .ZN(n31084) );
  OR2_X1 U37749 ( .A1(n31091), .A2(n31090), .ZN(n31092) );
  INV_X1 U37750 ( .A(n31093), .ZN(n31095) );
  OAI211_X1 U37751 ( .C1(n31097), .C2(n31096), .A(n31095), .B(n31094), .ZN(
        n31101) );
  OAI21_X1 U37752 ( .B1(n31099), .B2(n31098), .A(n31097), .ZN(n31100) );
  XNOR2_X1 U37753 ( .A(n31103), .B(n35296), .ZN(n35474) );
  OAI21_X1 U37754 ( .B1(n52121), .B2(n623), .A(n31104), .ZN(n31107) );
  AOI21_X1 U37755 ( .B1(n31107), .B2(n31106), .A(n31105), .ZN(n31108) );
  NAND3_X1 U37756 ( .A1(n31111), .A2(n31117), .A3(n623), .ZN(n31120) );
  NAND3_X1 U37757 ( .A1(n7093), .A2(n52121), .A3(n7658), .ZN(n31119) );
  NAND3_X1 U37758 ( .A1(n31117), .A2(n31116), .A3(n31115), .ZN(n31118) );
  AND3_X1 U37759 ( .A1(n31120), .A2(n31119), .A3(n31118), .ZN(n31127) );
  OAI21_X1 U37760 ( .B1(n31123), .B2(n31122), .A(n31121), .ZN(n31124) );
  INV_X1 U37761 ( .A(n31124), .ZN(n31126) );
  XNOR2_X1 U37762 ( .A(n31129), .B(n4565), .ZN(n31130) );
  XNOR2_X1 U37763 ( .A(n31131), .B(n31130), .ZN(n31133) );
  INV_X1 U37764 ( .A(n45105), .ZN(n31132) );
  XNOR2_X1 U37765 ( .A(n31133), .B(n31132), .ZN(n31134) );
  XNOR2_X1 U37766 ( .A(n31135), .B(n31134), .ZN(n31136) );
  XNOR2_X1 U37767 ( .A(n34163), .B(n31136), .ZN(n31153) );
  NAND2_X1 U37768 ( .A1(n31420), .A2(n31137), .ZN(n31139) );
  OR2_X1 U37771 ( .A1(n31141), .A2(n717), .ZN(n31142) );
  INV_X1 U37772 ( .A(n31144), .ZN(n31414) );
  AOI21_X1 U37773 ( .B1(n31414), .B2(n31899), .A(n31425), .ZN(n31148) );
  NAND3_X1 U37774 ( .A1(n31425), .A2(n31422), .A3(n31899), .ZN(n31145) );
  OAI211_X1 U37775 ( .C1(n31422), .C2(n31899), .A(n31145), .B(n31892), .ZN(
        n31147) );
  XNOR2_X1 U37776 ( .A(n35656), .B(n31153), .ZN(n31187) );
  AND2_X1 U37777 ( .A1(n31466), .A2(n32616), .ZN(n31465) );
  NAND2_X1 U37778 ( .A1(n32617), .A2(n31465), .ZN(n31555) );
  AND3_X1 U37781 ( .A1(n31157), .A2(n31555), .A3(n31156), .ZN(n31164) );
  MUX2_X1 U37782 ( .A(n31159), .B(n31475), .S(n31466), .Z(n31163) );
  NOR2_X1 U37783 ( .A1(n31166), .A2(n31165), .ZN(n31167) );
  OAI21_X1 U37784 ( .B1(n31168), .B2(n31549), .A(n31167), .ZN(n31186) );
  INV_X1 U37785 ( .A(n31454), .ZN(n31171) );
  AOI21_X1 U37786 ( .B1(n3847), .B2(n31452), .A(n31170), .ZN(n31175) );
  NAND2_X1 U37787 ( .A1(n31172), .A2(n31455), .ZN(n31174) );
  AND2_X1 U37788 ( .A1(n382), .A2(n31538), .ZN(n31181) );
  NAND2_X1 U37789 ( .A1(n32669), .A2(n31181), .ZN(n31173) );
  NAND4_X1 U37790 ( .A1(n31176), .A2(n31175), .A3(n31174), .A4(n31173), .ZN(
        n31185) );
  NAND2_X1 U37791 ( .A1(n31546), .A2(n31177), .ZN(n31178) );
  AND2_X1 U37792 ( .A1(n31179), .A2(n31178), .ZN(n31184) );
  NOR2_X1 U37793 ( .A1(n382), .A2(n31452), .ZN(n32671) );
  NAND2_X1 U37795 ( .A1(n31188), .A2(n32001), .ZN(n32516) );
  NAND2_X1 U37796 ( .A1(n7667), .A2(n32503), .ZN(n32510) );
  OAI21_X1 U37797 ( .B1(n31991), .B2(n32503), .A(n32510), .ZN(n31189) );
  NOR2_X1 U37798 ( .A1(n32507), .A2(n31995), .ZN(n32501) );
  NAND2_X1 U37799 ( .A1(n31189), .A2(n32501), .ZN(n31190) );
  NAND2_X1 U37800 ( .A1(n32516), .A2(n31190), .ZN(n31200) );
  NOR2_X1 U37801 ( .A1(n32506), .A2(n32511), .ZN(n31193) );
  OAI21_X1 U37802 ( .B1(n31193), .B2(n31192), .A(n31191), .ZN(n31199) );
  OR2_X1 U37803 ( .A1(n31995), .A2(n32004), .ZN(n32504) );
  NAND4_X1 U37804 ( .A1(n32504), .A2(n32508), .A3(n32503), .A4(n31194), .ZN(
        n31198) );
  NOR2_X1 U37805 ( .A1(n32004), .A2(n32503), .ZN(n32512) );
  OAI21_X1 U37806 ( .B1(n31993), .B2(n32512), .A(n31986), .ZN(n31197) );
  INV_X1 U37807 ( .A(n31194), .ZN(n31195) );
  NOR2_X1 U37808 ( .A1(n31201), .A2(n32478), .ZN(n32477) );
  OAI21_X1 U37809 ( .B1(n32478), .B2(n32487), .A(n32025), .ZN(n31202) );
  AOI22_X1 U37810 ( .A1(n31204), .A2(n32477), .B1(n31203), .B2(n31202), .ZN(
        n31213) );
  OAI21_X1 U37811 ( .B1(n31206), .B2(n32492), .A(n32028), .ZN(n31212) );
  NAND2_X1 U37812 ( .A1(n32025), .A2(n32473), .ZN(n32480) );
  OAI211_X1 U37813 ( .C1(n31209), .C2(n32480), .A(n31208), .B(n31207), .ZN(
        n31211) );
  XNOR2_X1 U37815 ( .A(n33142), .B(n33306), .ZN(n33252) );
  NOR2_X1 U37816 ( .A1(n31215), .A2(n6969), .ZN(n31217) );
  NAND2_X1 U37817 ( .A1(n31215), .A2(n31218), .ZN(n31216) );
  NOR2_X1 U37818 ( .A1(n31218), .A2(n32212), .ZN(n31220) );
  AOI22_X1 U37819 ( .A1(n32204), .A2(n31220), .B1(n31219), .B2(n31763), .ZN(
        n31227) );
  NAND2_X1 U37820 ( .A1(n50981), .A2(n32215), .ZN(n31223) );
  OAI211_X1 U37821 ( .C1(n31225), .C2(n32210), .A(n31763), .B(n32211), .ZN(
        n31226) );
  INV_X1 U37822 ( .A(n31229), .ZN(n31230) );
  NAND2_X1 U37823 ( .A1(n31230), .A2(n32244), .ZN(n31234) );
  AND2_X1 U37824 ( .A1(n32242), .A2(n32244), .ZN(n32256) );
  NAND2_X1 U37825 ( .A1(n32257), .A2(n32256), .ZN(n31233) );
  INV_X1 U37826 ( .A(n32247), .ZN(n31231) );
  NAND2_X1 U37827 ( .A1(n31231), .A2(n31781), .ZN(n31232) );
  NAND4_X1 U37828 ( .A1(n31234), .A2(n31788), .A3(n31233), .A4(n31232), .ZN(
        n31235) );
  NAND2_X1 U37829 ( .A1(n31235), .A2(n32254), .ZN(n31248) );
  OAI21_X1 U37830 ( .B1(n32230), .B2(n31783), .A(n31236), .ZN(n31237) );
  INV_X1 U37831 ( .A(n31237), .ZN(n31247) );
  AOI21_X1 U37832 ( .B1(n32246), .B2(n32243), .A(n622), .ZN(n31243) );
  INV_X1 U37833 ( .A(n31238), .ZN(n31239) );
  NAND3_X1 U37834 ( .A1(n31239), .A2(n32243), .A3(n32242), .ZN(n31242) );
  NAND4_X1 U37835 ( .A1(n31243), .A2(n31242), .A3(n31241), .A4(n31240), .ZN(
        n31246) );
  NAND3_X1 U37836 ( .A1(n32225), .A2(n31244), .A3(n32226), .ZN(n31245) );
  XNOR2_X1 U37837 ( .A(n35745), .B(n34503), .ZN(n31674) );
  XNOR2_X1 U37838 ( .A(n31674), .B(n33252), .ZN(n36832) );
  NOR2_X1 U37839 ( .A1(n7409), .A2(n31904), .ZN(n32827) );
  NAND2_X1 U37840 ( .A1(n32827), .A2(n32825), .ZN(n31251) );
  NAND3_X1 U37841 ( .A1(n31252), .A2(n31251), .A3(n31250), .ZN(n31256) );
  NAND2_X1 U37842 ( .A1(n32429), .A2(n32829), .ZN(n31254) );
  NAND2_X1 U37843 ( .A1(n32424), .A2(n31904), .ZN(n31253) );
  NOR2_X1 U37844 ( .A1(n31256), .A2(n31255), .ZN(n31263) );
  NAND2_X1 U37845 ( .A1(n32830), .A2(n32829), .ZN(n32814) );
  OAI21_X1 U37846 ( .B1(n32819), .B2(n32420), .A(n32828), .ZN(n31257) );
  NAND2_X1 U37847 ( .A1(n32814), .A2(n31257), .ZN(n31259) );
  NOR2_X1 U37848 ( .A1(n32829), .A2(n32420), .ZN(n32416) );
  OAI21_X1 U37849 ( .B1(n32823), .B2(n32821), .A(n32416), .ZN(n31261) );
  NAND2_X1 U37850 ( .A1(n31264), .A2(n31488), .ZN(n31268) );
  AND2_X1 U37851 ( .A1(n31266), .A2(n31265), .ZN(n31267) );
  OAI211_X1 U37852 ( .C1(n31488), .C2(n31273), .A(n31484), .B(n31490), .ZN(
        n31274) );
  NAND2_X1 U37853 ( .A1(n31275), .A2(n31274), .ZN(n31277) );
  NOR2_X1 U37854 ( .A1(n31284), .A2(n32066), .ZN(n31281) );
  OAI21_X1 U37855 ( .B1(n51639), .B2(n32409), .A(n31282), .ZN(n31283) );
  OAI211_X1 U37856 ( .C1(n32080), .C2(n51519), .A(n31286), .B(n32407), .ZN(
        n31287) );
  INV_X1 U37857 ( .A(n31289), .ZN(n31291) );
  AND2_X1 U37858 ( .A1(n32407), .A2(n32402), .ZN(n32070) );
  OAI21_X1 U37859 ( .B1(n31291), .B2(n32070), .A(n31290), .ZN(n31292) );
  OAI211_X1 U37860 ( .C1(n31302), .C2(n31311), .A(n31294), .B(n31300), .ZN(
        n31295) );
  NAND2_X1 U37861 ( .A1(n31296), .A2(n31295), .ZN(n31319) );
  MUX2_X1 U37862 ( .A(n31298), .B(n31297), .S(n51086), .Z(n31299) );
  INV_X1 U37863 ( .A(n31299), .ZN(n31318) );
  OR2_X1 U37864 ( .A1(n51086), .A2(n31300), .ZN(n31304) );
  NAND4_X1 U37865 ( .A1(n31304), .A2(n31303), .A3(n31302), .A4(n4607), .ZN(
        n31310) );
  INV_X1 U37866 ( .A(n31305), .ZN(n31308) );
  NAND3_X1 U37867 ( .A1(n31308), .A2(n51086), .A3(n31306), .ZN(n31309) );
  AND2_X1 U37868 ( .A1(n31310), .A2(n31309), .ZN(n31317) );
  NOR2_X1 U37869 ( .A1(n31312), .A2(n31311), .ZN(n31314) );
  OAI21_X1 U37870 ( .B1(n31315), .B2(n31314), .A(n31313), .ZN(n31316) );
  NAND2_X1 U37871 ( .A1(n32345), .A2(n32439), .ZN(n32444) );
  OAI21_X1 U37872 ( .B1(n31322), .B2(n31321), .A(n32440), .ZN(n31330) );
  NAND2_X1 U37873 ( .A1(n32056), .A2(n32438), .ZN(n31953) );
  NAND2_X1 U37874 ( .A1(n32057), .A2(n31953), .ZN(n31324) );
  NAND2_X1 U37875 ( .A1(n31959), .A2(n31324), .ZN(n31329) );
  OAI22_X1 U37876 ( .A1(n32042), .A2(n32051), .B1(n32047), .B2(n32439), .ZN(
        n31325) );
  NAND2_X1 U37877 ( .A1(n31325), .A2(n718), .ZN(n31328) );
  OR2_X1 U37878 ( .A1(n32352), .A2(n31326), .ZN(n31327) );
  XNOR2_X1 U37879 ( .A(n35115), .B(n36829), .ZN(n31350) );
  INV_X1 U37880 ( .A(n31333), .ZN(n31335) );
  AOI21_X1 U37881 ( .B1(n31336), .B2(n31335), .A(n31334), .ZN(n31337) );
  NAND2_X1 U37882 ( .A1(n31942), .A2(n31337), .ZN(n31349) );
  NAND2_X1 U37883 ( .A1(n31346), .A2(n31340), .ZN(n31341) );
  NAND3_X1 U37884 ( .A1(n31343), .A2(n31342), .A3(n31341), .ZN(n31345) );
  OAI21_X1 U37885 ( .B1(n31345), .B2(n31344), .A(n5682), .ZN(n31348) );
  XNOR2_X1 U37886 ( .A(n31350), .B(n37137), .ZN(n33263) );
  OR2_X1 U37887 ( .A1(n38552), .A2(n36141), .ZN(n36147) );
  NAND3_X1 U37889 ( .A1(n6734), .A2(n38558), .A3(n38213), .ZN(n31352) );
  INV_X1 U37890 ( .A(n31354), .ZN(n31362) );
  NOR2_X1 U37892 ( .A1(n38542), .A2(n31357), .ZN(n31361) );
  INV_X1 U37893 ( .A(n38550), .ZN(n36142) );
  NAND3_X1 U37894 ( .A1(n35170), .A2(n35178), .A3(n36305), .ZN(n31359) );
  OAI21_X1 U37895 ( .B1(n31845), .B2(n386), .A(n32297), .ZN(n31365) );
  OAI211_X1 U37896 ( .C1(n4299), .C2(n32299), .A(n31743), .B(n31369), .ZN(
        n31364) );
  NAND2_X1 U37897 ( .A1(n31747), .A2(n32295), .ZN(n31363) );
  NOR2_X1 U37898 ( .A1(n711), .A2(n386), .ZN(n31367) );
  NAND2_X1 U37899 ( .A1(n711), .A2(n31369), .ZN(n31371) );
  OAI21_X1 U37900 ( .B1(n32303), .B2(n31740), .A(n31369), .ZN(n31370) );
  INV_X1 U37901 ( .A(n31742), .ZN(n31855) );
  NAND4_X1 U37902 ( .A1(n31371), .A2(n31370), .A3(n31855), .A4(n31749), .ZN(
        n31373) );
  OAI21_X1 U37903 ( .B1(n32300), .B2(n31749), .A(n31846), .ZN(n31372) );
  INV_X1 U37904 ( .A(n31375), .ZN(n31378) );
  INV_X1 U37905 ( .A(n33006), .ZN(n31376) );
  XNOR2_X1 U37906 ( .A(n33017), .B(n31379), .ZN(n31382) );
  NOR2_X1 U37907 ( .A1(n33006), .A2(n31380), .ZN(n31381) );
  NAND2_X1 U37908 ( .A1(n31382), .A2(n31381), .ZN(n31390) );
  OAI211_X1 U37910 ( .C1(n33017), .C2(n31388), .A(n31387), .B(n8260), .ZN(
        n31389) );
  NAND3_X1 U37911 ( .A1(n31904), .A2(n31398), .A3(n32420), .ZN(n31393) );
  OAI211_X1 U37912 ( .C1(n32426), .C2(n31394), .A(n31393), .B(n31392), .ZN(
        n31396) );
  NOR2_X1 U37914 ( .A1(n31396), .A2(n8749), .ZN(n31408) );
  MUX2_X1 U37915 ( .A(n31400), .B(n31399), .S(n31398), .Z(n31407) );
  NOR2_X1 U37916 ( .A1(n32830), .A2(n31401), .ZN(n32423) );
  INV_X1 U37917 ( .A(n32424), .ZN(n31403) );
  NAND2_X1 U37918 ( .A1(n32423), .A2(n31405), .ZN(n31406) );
  NAND3_X2 U37919 ( .A1(n31408), .A2(n31407), .A3(n31406), .ZN(n35778) );
  XNOR2_X2 U37920 ( .A(n35778), .B(n51447), .ZN(n34739) );
  XNOR2_X1 U37921 ( .A(n34143), .B(n34739), .ZN(n31430) );
  NAND2_X1 U37922 ( .A1(n31414), .A2(n31892), .ZN(n31411) );
  NAND2_X1 U37923 ( .A1(n725), .A2(n31891), .ZN(n31409) );
  OAI22_X1 U37924 ( .A1(n31420), .A2(n31411), .B1(n31410), .B2(n31409), .ZN(
        n31417) );
  OAI211_X1 U37925 ( .C1(n31414), .C2(n31413), .A(n725), .B(n31412), .ZN(
        n31416) );
  NAND3_X1 U37926 ( .A1(n31414), .A2(n31413), .A3(n31425), .ZN(n31415) );
  NAND3_X1 U37927 ( .A1(n31898), .A2(n31419), .A3(n31418), .ZN(n31428) );
  OAI211_X1 U37928 ( .C1(n31423), .C2(n31422), .A(n31421), .B(n31420), .ZN(
        n31427) );
  XNOR2_X1 U37929 ( .A(n36932), .B(n33911), .ZN(n33751) );
  XNOR2_X1 U37930 ( .A(n33753), .B(n37065), .ZN(n36674) );
  XNOR2_X1 U37931 ( .A(n36674), .B(n33751), .ZN(n31429) );
  XNOR2_X1 U37932 ( .A(n31430), .B(n31429), .ZN(n31439) );
  XNOR2_X1 U37933 ( .A(n35512), .B(n4526), .ZN(n33473) );
  XNOR2_X1 U37934 ( .A(n31431), .B(n5016), .ZN(n31433) );
  XNOR2_X1 U37935 ( .A(n31433), .B(n31432), .ZN(n31434) );
  XNOR2_X1 U37936 ( .A(n31434), .B(n32520), .ZN(n31435) );
  XNOR2_X1 U37937 ( .A(n33914), .B(n31435), .ZN(n31436) );
  XNOR2_X1 U37938 ( .A(n33473), .B(n31436), .ZN(n31437) );
  XNOR2_X1 U37939 ( .A(n34146), .B(n31437), .ZN(n31438) );
  XNOR2_X1 U37940 ( .A(n31439), .B(n31438), .ZN(n31508) );
  NAND2_X1 U37941 ( .A1(n31440), .A2(n32663), .ZN(n31442) );
  NAND3_X1 U37942 ( .A1(n31546), .A2(n382), .A3(n32665), .ZN(n31441) );
  NAND3_X1 U37943 ( .A1(n31445), .A2(n31536), .A3(n31444), .ZN(n31446) );
  AND2_X1 U37945 ( .A1(n31546), .A2(n31447), .ZN(n31451) );
  INV_X1 U37946 ( .A(n31448), .ZN(n31449) );
  NAND3_X1 U37948 ( .A1(n31547), .A2(n31452), .A3(n31546), .ZN(n31453) );
  OAI21_X1 U37949 ( .B1(n31549), .B2(n31454), .A(n31453), .ZN(n31456) );
  NAND2_X1 U37950 ( .A1(n31456), .A2(n31455), .ZN(n31457) );
  XNOR2_X1 U37952 ( .A(n36669), .B(n34141), .ZN(n33908) );
  INV_X1 U37953 ( .A(n31461), .ZN(n31464) );
  NAND2_X1 U37954 ( .A1(n31462), .A2(n31557), .ZN(n31472) );
  NAND2_X1 U37955 ( .A1(n31472), .A2(n31463), .ZN(n32613) );
  MUX2_X1 U37956 ( .A(n31464), .B(n32613), .S(n31566), .Z(n31480) );
  NAND2_X1 U37957 ( .A1(n31465), .A2(n32609), .ZN(n31560) );
  INV_X1 U37958 ( .A(n31560), .ZN(n31469) );
  AND2_X1 U37959 ( .A1(n51106), .A2(n7626), .ZN(n31468) );
  XNOR2_X1 U37960 ( .A(n31466), .B(n51471), .ZN(n31467) );
  AOI22_X1 U37961 ( .A1(n31469), .A2(n51106), .B1(n31468), .B2(n31467), .ZN(
        n31479) );
  OAI211_X1 U37962 ( .C1(n32617), .C2(n31470), .A(n32622), .B(n7626), .ZN(
        n31474) );
  NAND3_X1 U37963 ( .A1(n31472), .A2(n31471), .A3(n32616), .ZN(n31473) );
  AND2_X1 U37964 ( .A1(n31474), .A2(n31473), .ZN(n31478) );
  INV_X1 U37965 ( .A(n31475), .ZN(n31476) );
  NAND3_X1 U37966 ( .A1(n31476), .A2(n32609), .A3(n32616), .ZN(n31477) );
  XNOR2_X1 U37967 ( .A(n33908), .B(n34829), .ZN(n33583) );
  NAND2_X1 U37968 ( .A1(n31481), .A2(n31490), .ZN(n31486) );
  INV_X1 U37969 ( .A(n31481), .ZN(n31482) );
  MUX2_X1 U37970 ( .A(n31486), .B(n31485), .S(n31484), .Z(n31506) );
  AOI21_X1 U37971 ( .B1(n31497), .B2(n31492), .A(n31491), .ZN(n31493) );
  NOR2_X1 U37973 ( .A1(n31497), .A2(n31496), .ZN(n31501) );
  OAI21_X1 U37974 ( .B1(n31499), .B2(n31498), .A(n31501), .ZN(n31504) );
  OAI21_X1 U37975 ( .B1(n31502), .B2(n31501), .A(n31500), .ZN(n31503) );
  XNOR2_X1 U37977 ( .A(n51663), .B(n34553), .ZN(n31507) );
  XNOR2_X1 U37978 ( .A(n31507), .B(n33583), .ZN(n34476) );
  AND2_X1 U37979 ( .A1(n3099), .A2(n31512), .ZN(n31514) );
  INV_X1 U37980 ( .A(n31515), .ZN(n31521) );
  INV_X1 U37981 ( .A(n33026), .ZN(n33035) );
  NAND4_X1 U37982 ( .A1(n31528), .A2(n33028), .A3(n31527), .A4(n31526), .ZN(
        n31535) );
  OAI211_X1 U37983 ( .C1(n32867), .C2(n32876), .A(n33041), .B(n719), .ZN(
        n31532) );
  NAND2_X1 U37984 ( .A1(n32879), .A2(n32867), .ZN(n33025) );
  NAND2_X1 U37985 ( .A1(n33025), .A2(n33026), .ZN(n31529) );
  NAND4_X1 U37986 ( .A1(n32645), .A2(n32874), .A3(n8544), .A4(n31529), .ZN(
        n31531) );
  OAI211_X1 U37987 ( .C1(n31533), .C2(n31532), .A(n31531), .B(n31530), .ZN(
        n31534) );
  NAND2_X1 U37988 ( .A1(n31537), .A2(n31536), .ZN(n31552) );
  OR2_X1 U37989 ( .A1(n31539), .A2(n31538), .ZN(n31543) );
  INV_X1 U37990 ( .A(n31541), .ZN(n31542) );
  NOR2_X1 U37991 ( .A1(n381), .A2(n2011), .ZN(n31548) );
  AND2_X1 U37992 ( .A1(n31554), .A2(n31555), .ZN(n31572) );
  AOI22_X1 U37993 ( .A1(n31564), .A2(n31563), .B1(n31562), .B2(n31561), .ZN(
        n31571) );
  INV_X1 U37994 ( .A(n31565), .ZN(n31568) );
  INV_X1 U37995 ( .A(n34128), .ZN(n31574) );
  XNOR2_X1 U37996 ( .A(n33489), .B(n34810), .ZN(n31620) );
  AOI22_X1 U37997 ( .A1(n31631), .A2(n31632), .B1(n31576), .B2(n31625), .ZN(
        n31593) );
  AOI21_X1 U37998 ( .B1(n31636), .B2(n31577), .A(n31637), .ZN(n31592) );
  NOR2_X1 U38000 ( .A1(n31636), .A2(n31583), .ZN(n31589) );
  AOI21_X1 U38001 ( .B1(n31586), .B2(n31585), .A(n31584), .ZN(n31588) );
  OAI21_X1 U38002 ( .B1(n31589), .B2(n31588), .A(n31587), .ZN(n31590) );
  XNOR2_X1 U38003 ( .A(n31595), .B(n31594), .ZN(n31596) );
  XNOR2_X1 U38004 ( .A(n51413), .B(n31596), .ZN(n31597) );
  XNOR2_X1 U38005 ( .A(n376), .B(n31597), .ZN(n31598) );
  XNOR2_X1 U38006 ( .A(n37256), .B(n31598), .ZN(n31618) );
  NAND2_X1 U38007 ( .A1(n32540), .A2(n32900), .ZN(n32632) );
  OAI21_X1 U38008 ( .B1(n32894), .B2(n32632), .A(n32631), .ZN(n31599) );
  NAND2_X1 U38009 ( .A1(n31603), .A2(n32916), .ZN(n31601) );
  OAI21_X1 U38010 ( .B1(n32900), .B2(n32908), .A(n32915), .ZN(n31600) );
  NAND2_X1 U38011 ( .A1(n6269), .A2(n32915), .ZN(n31602) );
  NAND4_X1 U38012 ( .A1(n32918), .A2(n31602), .A3(n32540), .A4(n32894), .ZN(
        n31605) );
  OAI211_X1 U38013 ( .C1(n32894), .C2(n32634), .A(n31603), .B(n32901), .ZN(
        n31604) );
  OAI21_X1 U38014 ( .B1(n32561), .B2(n32107), .A(n8468), .ZN(n31606) );
  AOI22_X1 U38015 ( .A1(n31607), .A2(n31606), .B1(n32573), .B2(n32105), .ZN(
        n31617) );
  NAND2_X1 U38016 ( .A1(n624), .A2(n31608), .ZN(n32575) );
  INV_X1 U38017 ( .A(n32575), .ZN(n32091) );
  XNOR2_X1 U38018 ( .A(n31608), .B(n32560), .ZN(n31612) );
  OAI211_X1 U38019 ( .C1(n31612), .C2(n32558), .A(n31611), .B(n32575), .ZN(
        n31615) );
  NOR2_X1 U38020 ( .A1(n32561), .A2(n32566), .ZN(n32097) );
  OAI21_X1 U38021 ( .B1(n624), .B2(n32105), .A(n32095), .ZN(n31613) );
  XNOR2_X1 U38025 ( .A(n33335), .B(n34535), .ZN(n37251) );
  XNOR2_X1 U38026 ( .A(n37251), .B(n31618), .ZN(n31619) );
  INV_X1 U38027 ( .A(n31622), .ZN(n31623) );
  OAI21_X1 U38028 ( .B1(n31625), .B2(n31624), .A(n31623), .ZN(n31628) );
  INV_X1 U38029 ( .A(n31626), .ZN(n31627) );
  INV_X1 U38030 ( .A(n31633), .ZN(n31635) );
  OAI21_X1 U38031 ( .B1(n31636), .B2(n31635), .A(n31634), .ZN(n31642) );
  NOR2_X1 U38032 ( .A1(n32725), .A2(n32719), .ZN(n31643) );
  AOI22_X1 U38033 ( .A1(n32714), .A2(n32315), .B1(n31643), .B2(n32312), .ZN(
        n31654) );
  NAND2_X1 U38034 ( .A1(n32731), .A2(n2359), .ZN(n31653) );
  NOR2_X1 U38036 ( .A1(n32716), .A2(n32463), .ZN(n31968) );
  INV_X1 U38037 ( .A(n31968), .ZN(n31647) );
  NAND3_X1 U38038 ( .A1(n31648), .A2(n31647), .A3(n32720), .ZN(n31651) );
  INV_X1 U38039 ( .A(n32312), .ZN(n31650) );
  NAND2_X1 U38040 ( .A1(n31968), .A2(n32732), .ZN(n31649) );
  NAND4_X1 U38041 ( .A1(n31651), .A2(n32318), .A3(n31650), .A4(n31649), .ZN(
        n31652) );
  XNOR2_X1 U38042 ( .A(n36747), .B(n44046), .ZN(n31655) );
  XNOR2_X1 U38043 ( .A(n31655), .B(n33938), .ZN(n31656) );
  XNOR2_X1 U38044 ( .A(n31657), .B(n31656), .ZN(n34522) );
  AOI21_X1 U38045 ( .B1(n31659), .B2(n31658), .A(n32705), .ZN(n31662) );
  NOR2_X1 U38046 ( .A1(n32700), .A2(n31660), .ZN(n31661) );
  INV_X1 U38047 ( .A(n32700), .ZN(n31663) );
  NOR2_X1 U38048 ( .A1(n31663), .A2(n32708), .ZN(n31664) );
  OR2_X1 U38049 ( .A1(n31665), .A2(n31664), .ZN(n31672) );
  OAI211_X1 U38050 ( .C1(n32327), .C2(n32324), .A(n32688), .B(n31666), .ZN(
        n31667) );
  OAI211_X1 U38052 ( .C1(n32688), .C2(n31669), .A(n31668), .B(n1988), .ZN(
        n31670) );
  XNOR2_X1 U38053 ( .A(n34605), .B(n35115), .ZN(n33728) );
  OAI21_X1 U38054 ( .B1(n31675), .B2(n2094), .A(n2237), .ZN(n31678) );
  NAND3_X1 U38055 ( .A1(n31676), .A2(n2098), .A3(n31675), .ZN(n31677) );
  AND2_X1 U38056 ( .A1(n31678), .A2(n31677), .ZN(n31698) );
  AND2_X1 U38057 ( .A1(n31680), .A2(n31679), .ZN(n31681) );
  OAI21_X1 U38058 ( .B1(n31682), .B2(n31681), .A(n7598), .ZN(n31688) );
  NAND4_X1 U38059 ( .A1(n31688), .A2(n31687), .A3(n31686), .A4(n31685), .ZN(
        n31697) );
  AOI22_X1 U38060 ( .A1(n2098), .A2(n31690), .B1(n31689), .B2(n7598), .ZN(
        n31696) );
  INV_X1 U38061 ( .A(n31692), .ZN(n31694) );
  XNOR2_X1 U38062 ( .A(n35471), .B(n37023), .ZN(n33925) );
  NAND2_X1 U38063 ( .A1(n32118), .A2(n31699), .ZN(n31703) );
  NAND2_X1 U38064 ( .A1(n31711), .A2(n31700), .ZN(n32124) );
  MUX2_X1 U38065 ( .A(n31703), .B(n31702), .S(n31701), .Z(n31717) );
  NAND2_X1 U38066 ( .A1(n31706), .A2(n31708), .ZN(n31704) );
  OAI211_X1 U38067 ( .C1(n31706), .C2(n31705), .A(n31704), .B(n32125), .ZN(
        n31707) );
  INV_X1 U38068 ( .A(n31710), .ZN(n31715) );
  NAND2_X1 U38069 ( .A1(n31712), .A2(n31711), .ZN(n31713) );
  AOI21_X1 U38070 ( .B1(n31715), .B2(n31714), .A(n31713), .ZN(n31716) );
  XNOR2_X1 U38071 ( .A(n34163), .B(n34169), .ZN(n31722) );
  XNOR2_X1 U38072 ( .A(n35108), .B(n2117), .ZN(n31718) );
  XNOR2_X1 U38073 ( .A(n31719), .B(n31718), .ZN(n31720) );
  XNOR2_X1 U38074 ( .A(n33142), .B(n31720), .ZN(n31721) );
  XNOR2_X1 U38075 ( .A(n31722), .B(n31721), .ZN(n31723) );
  XNOR2_X1 U38076 ( .A(n31723), .B(n50982), .ZN(n31760) );
  INV_X1 U38077 ( .A(n32788), .ZN(n31724) );
  NOR2_X1 U38079 ( .A1(n31725), .A2(n32784), .ZN(n32797) );
  NAND2_X1 U38080 ( .A1(n32797), .A2(n32785), .ZN(n32282) );
  INV_X1 U38081 ( .A(n32282), .ZN(n31729) );
  INV_X1 U38082 ( .A(n31725), .ZN(n32793) );
  AND2_X1 U38083 ( .A1(n32794), .A2(n31727), .ZN(n31728) );
  INV_X1 U38084 ( .A(n32150), .ZN(n32287) );
  OAI211_X1 U38085 ( .C1(n32782), .C2(n31729), .A(n31728), .B(n32287), .ZN(
        n31738) );
  INV_X1 U38086 ( .A(n31864), .ZN(n32158) );
  NAND2_X1 U38087 ( .A1(n31725), .A2(n32784), .ZN(n31730) );
  NOR2_X1 U38088 ( .A1(n31730), .A2(n32788), .ZN(n31731) );
  AOI22_X1 U38089 ( .A1(n32778), .A2(n32158), .B1(n31863), .B2(n31731), .ZN(
        n31737) );
  NOR2_X1 U38090 ( .A1(n31733), .A2(n32157), .ZN(n31732) );
  INV_X1 U38091 ( .A(n32791), .ZN(n32780) );
  AOI22_X1 U38092 ( .A1(n32778), .A2(n31732), .B1(n32780), .B2(n32797), .ZN(
        n31736) );
  INV_X1 U38093 ( .A(n31733), .ZN(n31734) );
  OAI21_X1 U38094 ( .B1(n31734), .B2(n31725), .A(n32163), .ZN(n31735) );
  INV_X1 U38095 ( .A(n42419), .ZN(n31739) );
  XNOR2_X1 U38096 ( .A(n34604), .B(n31739), .ZN(n31759) );
  NOR2_X1 U38097 ( .A1(n32299), .A2(n31740), .ZN(n31741) );
  NOR2_X1 U38098 ( .A1(n4434), .A2(n31746), .ZN(n31853) );
  AND2_X1 U38099 ( .A1(n31749), .A2(n435), .ZN(n31750) );
  AOI22_X1 U38100 ( .A1(n32300), .A2(n31741), .B1(n31853), .B2(n31750), .ZN(
        n31758) );
  INV_X1 U38101 ( .A(n31744), .ZN(n31844) );
  AOI22_X1 U38102 ( .A1(n31742), .A2(n31849), .B1(n31844), .B2(n32295), .ZN(
        n32305) );
  NOR2_X1 U38103 ( .A1(n31744), .A2(n31743), .ZN(n31745) );
  NAND2_X1 U38105 ( .A1(n31749), .A2(n386), .ZN(n31752) );
  INV_X1 U38106 ( .A(n31750), .ZN(n31751) );
  OAI22_X1 U38107 ( .A1(n711), .A2(n31752), .B1(n31751), .B2(n32295), .ZN(
        n31754) );
  XNOR2_X1 U38108 ( .A(n37304), .B(n31759), .ZN(n33262) );
  XNOR2_X1 U38109 ( .A(n31760), .B(n33262), .ZN(n31761) );
  XNOR2_X1 U38110 ( .A(n33925), .B(n31761), .ZN(n31762) );
  BUF_X2 U38111 ( .A(n35017), .Z(n36338) );
  NAND2_X1 U38112 ( .A1(n31767), .A2(n50981), .ZN(n31766) );
  XNOR2_X1 U38113 ( .A(n32194), .B(n6969), .ZN(n31765) );
  NOR2_X1 U38114 ( .A1(n31766), .A2(n31765), .ZN(n31775) );
  OAI22_X1 U38115 ( .A1(n31770), .A2(n32197), .B1(n50980), .B2(n31767), .ZN(
        n31773) );
  NOR2_X1 U38116 ( .A1(n31769), .A2(n6969), .ZN(n31772) );
  NAND3_X1 U38117 ( .A1(n31770), .A2(n32215), .A3(n32204), .ZN(n31771) );
  INV_X1 U38119 ( .A(n31779), .ZN(n31780) );
  NAND2_X1 U38120 ( .A1(n32252), .A2(n31781), .ZN(n31782) );
  NOR2_X1 U38121 ( .A1(n32246), .A2(n32251), .ZN(n31784) );
  AOI21_X1 U38122 ( .B1(n31785), .B2(n32231), .A(n31784), .ZN(n31786) );
  OAI211_X1 U38123 ( .C1(n32225), .C2(n31788), .A(n31787), .B(n31786), .ZN(
        n35768) );
  XNOR2_X1 U38124 ( .A(n36758), .B(n35768), .ZN(n34888) );
  XNOR2_X1 U38125 ( .A(n34888), .B(n51366), .ZN(n31814) );
  NAND2_X1 U38126 ( .A1(n31798), .A2(n52047), .ZN(n31790) );
  OAI21_X1 U38127 ( .B1(n31791), .B2(n31790), .A(n31789), .ZN(n31796) );
  INV_X1 U38128 ( .A(n31792), .ZN(n31794) );
  NOR2_X1 U38129 ( .A1(n31796), .A2(n31795), .ZN(n31806) );
  INV_X1 U38130 ( .A(n31797), .ZN(n31878) );
  NAND3_X1 U38131 ( .A1(n31878), .A2(n31799), .A3(n31798), .ZN(n31805) );
  XNOR2_X1 U38132 ( .A(n52047), .B(n31800), .ZN(n31802) );
  OAI21_X1 U38133 ( .B1(n31803), .B2(n31802), .A(n31801), .ZN(n31804) );
  INV_X1 U38134 ( .A(n31807), .ZN(n31809) );
  XNOR2_X1 U38135 ( .A(n31809), .B(n31808), .ZN(n31810) );
  XNOR2_X1 U38136 ( .A(n37318), .B(n31810), .ZN(n31811) );
  XNOR2_X1 U38137 ( .A(n32628), .B(n32644), .ZN(n36761) );
  XNOR2_X1 U38138 ( .A(n31812), .B(n36761), .ZN(n31813) );
  XNOR2_X1 U38139 ( .A(n31814), .B(n31813), .ZN(n31842) );
  OAI21_X1 U38140 ( .B1(n31816), .B2(n31821), .A(n31815), .ZN(n31818) );
  AOI22_X1 U38141 ( .A1(n31820), .A2(n31819), .B1(n31818), .B2(n31817), .ZN(
        n31834) );
  INV_X1 U38142 ( .A(n31820), .ZN(n31824) );
  OAI21_X1 U38143 ( .B1(n31824), .B2(n31823), .A(n31822), .ZN(n31825) );
  INV_X1 U38144 ( .A(n31825), .ZN(n31833) );
  OAI21_X1 U38145 ( .B1(n31830), .B2(n31829), .A(n31828), .ZN(n31831) );
  AND2_X1 U38146 ( .A1(n32960), .A2(n32760), .ZN(n32767) );
  MUX2_X1 U38147 ( .A(n32767), .B(n32762), .S(n32771), .Z(n31838) );
  NAND2_X1 U38149 ( .A1(n32175), .A2(n32965), .ZN(n32759) );
  INV_X1 U38150 ( .A(n32767), .ZN(n32532) );
  NOR2_X1 U38151 ( .A1(n32532), .A2(n32962), .ZN(n32773) );
  AND2_X1 U38152 ( .A1(n32965), .A2(n32957), .ZN(n32966) );
  NOR2_X1 U38153 ( .A1(n3303), .A2(n32765), .ZN(n31836) );
  OAI21_X1 U38154 ( .B1(n32773), .B2(n31836), .A(n32175), .ZN(n31837) );
  XNOR2_X1 U38155 ( .A(n31839), .B(n35124), .ZN(n31841) );
  INV_X1 U38156 ( .A(n35283), .ZN(n31840) );
  XNOR2_X1 U38157 ( .A(n31840), .B(n31841), .ZN(n33539) );
  OAI21_X1 U38158 ( .B1(n32300), .B2(n31844), .A(n31843), .ZN(n31861) );
  INV_X1 U38159 ( .A(n31845), .ZN(n31848) );
  NAND2_X1 U38160 ( .A1(n32302), .A2(n31846), .ZN(n31847) );
  AND2_X1 U38161 ( .A1(n31848), .A2(n31847), .ZN(n31860) );
  INV_X1 U38162 ( .A(n31849), .ZN(n31852) );
  INV_X1 U38163 ( .A(n32295), .ZN(n31851) );
  NAND3_X1 U38164 ( .A1(n31852), .A2(n31851), .A3(n435), .ZN(n31859) );
  INV_X1 U38165 ( .A(n31853), .ZN(n31856) );
  NAND2_X1 U38167 ( .A1(n31857), .A2(n32302), .ZN(n31858) );
  NOR2_X1 U38168 ( .A1(n32157), .A2(n31725), .ZN(n32164) );
  NAND2_X1 U38169 ( .A1(n31862), .A2(n32164), .ZN(n31868) );
  INV_X1 U38171 ( .A(n31865), .ZN(n31867) );
  OAI21_X1 U38172 ( .B1(n32787), .B2(n31725), .A(n32784), .ZN(n32779) );
  OR2_X1 U38173 ( .A1(n32782), .A2(n32779), .ZN(n31866) );
  XNOR2_X1 U38174 ( .A(n34359), .B(n34294), .ZN(n35685) );
  XNOR2_X1 U38175 ( .A(n36766), .B(n35685), .ZN(n33668) );
  NAND2_X1 U38176 ( .A1(n35017), .A2(n38142), .ZN(n38136) );
  INV_X1 U38177 ( .A(n38142), .ZN(n36337) );
  XNOR2_X1 U38179 ( .A(n35345), .B(n34841), .ZN(n35227) );
  NOR3_X1 U38180 ( .A1(n5912), .A2(n31886), .A3(n31870), .ZN(n31872) );
  AND2_X1 U38181 ( .A1(n31873), .A2(n31872), .ZN(n31875) );
  AOI22_X1 U38182 ( .A1(n31877), .A2(n31876), .B1(n31875), .B2(n31874), .ZN(
        n31890) );
  NAND3_X1 U38183 ( .A1(n31879), .A2(n31878), .A3(n31886), .ZN(n31889) );
  NAND2_X1 U38184 ( .A1(n31881), .A2(n31880), .ZN(n31888) );
  NAND2_X1 U38185 ( .A1(n31882), .A2(n31019), .ZN(n31884) );
  OAI211_X1 U38186 ( .C1(n31886), .C2(n31885), .A(n31884), .B(n51479), .ZN(
        n31887) );
  XNOR2_X1 U38187 ( .A(n35227), .B(n35635), .ZN(n37285) );
  NAND4_X1 U38188 ( .A1(n31893), .A2(n620), .A3(n31892), .A4(n31891), .ZN(
        n31894) );
  OAI21_X1 U38189 ( .B1(n31895), .B2(n31149), .A(n31894), .ZN(n31896) );
  NOR2_X1 U38190 ( .A1(n31897), .A2(n31896), .ZN(n31901) );
  XNOR2_X1 U38191 ( .A(n37285), .B(n33395), .ZN(n31924) );
  INV_X1 U38192 ( .A(n32822), .ZN(n31902) );
  NOR2_X1 U38193 ( .A1(n32830), .A2(n31902), .ZN(n31907) );
  OAI22_X1 U38195 ( .A1(n32823), .A2(n51630), .B1(n31904), .B2(n32420), .ZN(
        n31906) );
  NOR2_X1 U38196 ( .A1(n31907), .A2(n31906), .ZN(n31908) );
  AOI21_X1 U38197 ( .B1(n32852), .B2(n32374), .A(n32389), .ZN(n31916) );
  XNOR2_X1 U38198 ( .A(n31911), .B(n31910), .ZN(n31913) );
  NAND2_X1 U38199 ( .A1(n32381), .A2(n32840), .ZN(n31912) );
  AND4_X1 U38200 ( .A1(n31914), .A2(n31913), .A3(n32389), .A4(n31912), .ZN(
        n31915) );
  NOR2_X1 U38201 ( .A1(n31916), .A2(n31915), .ZN(n31922) );
  NOR2_X1 U38202 ( .A1(n32843), .A2(n32386), .ZN(n32837) );
  INV_X1 U38203 ( .A(n32837), .ZN(n31919) );
  INV_X1 U38204 ( .A(n32844), .ZN(n31918) );
  NAND2_X1 U38205 ( .A1(n32389), .A2(n32850), .ZN(n31917) );
  OAI211_X1 U38206 ( .C1(n31920), .C2(n31919), .A(n31918), .B(n31917), .ZN(
        n31921) );
  AND2_X1 U38207 ( .A1(n31922), .A2(n31921), .ZN(n34116) );
  XNOR2_X1 U38208 ( .A(n31923), .B(n34116), .ZN(n33397) );
  XNOR2_X1 U38209 ( .A(n33397), .B(n34433), .ZN(n35637) );
  XNOR2_X1 U38210 ( .A(n31924), .B(n35637), .ZN(n31965) );
  XNOR2_X1 U38211 ( .A(n41272), .B(n47737), .ZN(n31925) );
  XNOR2_X1 U38212 ( .A(n31926), .B(n31925), .ZN(n31927) );
  XNOR2_X1 U38213 ( .A(n31928), .B(n31927), .ZN(n31929) );
  XNOR2_X1 U38214 ( .A(n35088), .B(n31929), .ZN(n31930) );
  XNOR2_X1 U38215 ( .A(n31930), .B(n35085), .ZN(n31946) );
  NOR2_X1 U38216 ( .A1(n31932), .A2(n31931), .ZN(n31944) );
  OAI21_X1 U38217 ( .B1(n31935), .B2(n31934), .A(n31933), .ZN(n31937) );
  NAND2_X1 U38218 ( .A1(n31937), .A2(n31936), .ZN(n31943) );
  INV_X1 U38219 ( .A(n31938), .ZN(n31939) );
  NAND3_X1 U38220 ( .A1(n31334), .A2(n5682), .A3(n31939), .ZN(n31941) );
  XNOR2_X1 U38221 ( .A(n35544), .B(n35536), .ZN(n32292) );
  INV_X1 U38222 ( .A(n32292), .ZN(n31945) );
  XNOR2_X1 U38223 ( .A(n31946), .B(n31945), .ZN(n31963) );
  INV_X1 U38224 ( .A(n31947), .ZN(n32063) );
  NOR2_X1 U38225 ( .A1(n32396), .A2(n51520), .ZN(n32410) );
  OAI21_X1 U38226 ( .B1(n8253), .B2(n32063), .A(n32410), .ZN(n31952) );
  NAND2_X1 U38227 ( .A1(n32411), .A2(n32080), .ZN(n31951) );
  INV_X1 U38228 ( .A(n32081), .ZN(n31948) );
  NAND2_X1 U38229 ( .A1(n31948), .A2(n32074), .ZN(n31949) );
  INV_X1 U38230 ( .A(n31953), .ZN(n31958) );
  NAND2_X1 U38231 ( .A1(n31955), .A2(n31954), .ZN(n31957) );
  INV_X1 U38232 ( .A(n31959), .ZN(n31962) );
  INV_X1 U38233 ( .A(n32347), .ZN(n31960) );
  NOR3_X1 U38234 ( .A1(n31960), .A2(n32345), .A3(n718), .ZN(n31961) );
  XNOR2_X1 U38235 ( .A(n31963), .B(n34109), .ZN(n31964) );
  INV_X1 U38237 ( .A(n31967), .ZN(n31985) );
  NAND3_X1 U38238 ( .A1(n32458), .A2(n31968), .A3(n32719), .ZN(n32321) );
  AND2_X1 U38239 ( .A1(n32725), .A2(n32732), .ZN(n32313) );
  INV_X1 U38240 ( .A(n31969), .ZN(n31970) );
  NAND2_X1 U38241 ( .A1(n31970), .A2(n32732), .ZN(n32722) );
  AND3_X1 U38242 ( .A1(n31971), .A2(n32321), .A3(n32722), .ZN(n31984) );
  INV_X1 U38243 ( .A(n32718), .ZN(n31973) );
  AOI21_X1 U38244 ( .B1(n32720), .B2(n32725), .A(n32315), .ZN(n31972) );
  INV_X1 U38245 ( .A(n32318), .ZN(n32730) );
  NOR2_X1 U38247 ( .A1(n32315), .A2(n32720), .ZN(n32460) );
  INV_X1 U38248 ( .A(n32460), .ZN(n31975) );
  OAI21_X1 U38249 ( .B1(n32311), .B2(n32719), .A(n31648), .ZN(n31974) );
  NAND4_X1 U38250 ( .A1(n31975), .A2(n2483), .A3(n31974), .A4(n32458), .ZN(
        n31982) );
  NAND4_X1 U38251 ( .A1(n31648), .A2(n32316), .A3(n32724), .A4(n32716), .ZN(
        n31979) );
  INV_X1 U38252 ( .A(n32465), .ZN(n31976) );
  NAND2_X1 U38253 ( .A1(n32720), .A2(n31976), .ZN(n31978) );
  OAI211_X1 U38255 ( .C1(n32715), .C2(n31979), .A(n31978), .B(n31977), .ZN(
        n31980) );
  INV_X1 U38256 ( .A(n31980), .ZN(n31981) );
  XNOR2_X1 U38257 ( .A(n33703), .B(n31985), .ZN(n33383) );
  NAND2_X1 U38258 ( .A1(n31986), .A2(n32503), .ZN(n31988) );
  NAND2_X1 U38259 ( .A1(n31992), .A2(n32511), .ZN(n31998) );
  OAI211_X1 U38260 ( .C1(n31996), .C2(n32508), .A(n31995), .B(n31994), .ZN(
        n31997) );
  AOI22_X1 U38261 ( .A1(n32000), .A2(n31999), .B1(n31998), .B2(n31997), .ZN(
        n32012) );
  NAND3_X1 U38262 ( .A1(n32001), .A2(n32508), .A3(n32509), .ZN(n32002) );
  AND2_X1 U38263 ( .A1(n32003), .A2(n32002), .ZN(n32011) );
  OAI211_X1 U38264 ( .C1(n7897), .C2(n32004), .A(n32508), .B(n32507), .ZN(
        n32006) );
  INV_X1 U38265 ( .A(n32006), .ZN(n32008) );
  AOI22_X1 U38266 ( .A1(n8722), .A2(n32009), .B1(n32008), .B2(n32007), .ZN(
        n32010) );
  NAND4_X2 U38267 ( .A1(n32012), .A2(n32010), .A3(n32011), .A4(n32013), .ZN(
        n36812) );
  AOI21_X1 U38269 ( .B1(n32017), .B2(n32025), .A(n32016), .ZN(n32018) );
  NAND2_X1 U38270 ( .A1(n32486), .A2(n32472), .ZN(n32020) );
  NAND4_X1 U38271 ( .A1(n32021), .A2(n32484), .A3(n32478), .A4(n32020), .ZN(
        n32022) );
  AND2_X1 U38272 ( .A1(n32023), .A2(n32022), .ZN(n32033) );
  OAI21_X1 U38273 ( .B1(n32487), .B2(n32485), .A(n32025), .ZN(n32026) );
  AOI21_X1 U38274 ( .B1(n709), .B2(n32489), .A(n32028), .ZN(n32029) );
  NAND2_X1 U38275 ( .A1(n32030), .A2(n32029), .ZN(n32031) );
  NAND4_X2 U38276 ( .A1(n32034), .A2(n32032), .A3(n32031), .A4(n32033), .ZN(
        n34455) );
  XNOR2_X2 U38277 ( .A(n36812), .B(n34455), .ZN(n37095) );
  XNOR2_X1 U38278 ( .A(n33383), .B(n37095), .ZN(n34770) );
  XNOR2_X1 U38279 ( .A(n32860), .B(n37113), .ZN(n36731) );
  INV_X1 U38280 ( .A(n32935), .ZN(n34453) );
  XNOR2_X1 U38281 ( .A(n32035), .B(n32267), .ZN(n32036) );
  XNOR2_X1 U38282 ( .A(n32037), .B(n32036), .ZN(n32038) );
  XNOR2_X1 U38283 ( .A(n34453), .B(n32038), .ZN(n32039) );
  XNOR2_X1 U38284 ( .A(n36731), .B(n32039), .ZN(n32040) );
  INV_X1 U38285 ( .A(n32044), .ZN(n32045) );
  NAND3_X1 U38287 ( .A1(n32045), .A2(n3703), .A3(n32056), .ZN(n32046) );
  AOI21_X1 U38288 ( .B1(n32046), .B2(n32436), .A(n32351), .ZN(n32050) );
  NOR2_X1 U38289 ( .A1(n32050), .A2(n32049), .ZN(n32060) );
  NOR2_X1 U38290 ( .A1(n32056), .A2(n32438), .ZN(n32446) );
  NAND2_X1 U38291 ( .A1(n32446), .A2(n32051), .ZN(n32449) );
  INV_X1 U38292 ( .A(n32452), .ZN(n32054) );
  NAND2_X1 U38293 ( .A1(n32438), .A2(n32356), .ZN(n32053) );
  NAND2_X1 U38294 ( .A1(n32056), .A2(n32453), .ZN(n32052) );
  NAND4_X1 U38295 ( .A1(n32054), .A2(n32440), .A3(n32053), .A4(n32052), .ZN(
        n32055) );
  AND2_X1 U38296 ( .A1(n32449), .A2(n32055), .ZN(n32059) );
  AND2_X1 U38299 ( .A1(n32407), .A2(n32066), .ZN(n32399) );
  INV_X1 U38300 ( .A(n32399), .ZN(n32068) );
  INV_X1 U38301 ( .A(n32398), .ZN(n32067) );
  INV_X1 U38302 ( .A(n32070), .ZN(n32073) );
  OAI21_X1 U38303 ( .B1(n32074), .B2(n32073), .A(n32072), .ZN(n32079) );
  NAND2_X1 U38304 ( .A1(n714), .A2(n7430), .ZN(n32077) );
  NAND3_X1 U38305 ( .A1(n32396), .A2(n32408), .A3(n51519), .ZN(n32076) );
  OAI22_X1 U38306 ( .A1(n32077), .A2(n32076), .B1(n32075), .B2(n32396), .ZN(
        n32078) );
  NOR2_X1 U38307 ( .A1(n32079), .A2(n32078), .ZN(n32084) );
  OAI21_X1 U38308 ( .B1(n32081), .B2(n32080), .A(n51638), .ZN(n32082) );
  XNOR2_X1 U38309 ( .A(n35618), .B(n36807), .ZN(n33607) );
  NOR2_X1 U38310 ( .A1(n32107), .A2(n32560), .ZN(n32103) );
  XNOR2_X1 U38311 ( .A(n32105), .B(n32558), .ZN(n32092) );
  OAI21_X1 U38312 ( .B1(n8468), .B2(n32089), .A(n854), .ZN(n32090) );
  XNOR2_X1 U38313 ( .A(n32566), .B(n32560), .ZN(n32094) );
  INV_X1 U38314 ( .A(n32103), .ZN(n32093) );
  NAND4_X1 U38315 ( .A1(n32094), .A2(n32093), .A3(n32096), .A4(n32561), .ZN(
        n32099) );
  INV_X1 U38316 ( .A(n32095), .ZN(n32569) );
  NAND4_X1 U38317 ( .A1(n32101), .A2(n32100), .A3(n32099), .A4(n32098), .ZN(
        n32117) );
  AOI21_X1 U38318 ( .B1(n32104), .B2(n32103), .A(n32102), .ZN(n32115) );
  NAND4_X1 U38319 ( .A1(n32106), .A2(n32105), .A3(n32574), .A4(n32566), .ZN(
        n32110) );
  NAND2_X1 U38320 ( .A1(n32108), .A2(n32107), .ZN(n32109) );
  AND2_X1 U38321 ( .A1(n32109), .A2(n32110), .ZN(n32113) );
  INV_X1 U38322 ( .A(n32111), .ZN(n32112) );
  OAI211_X1 U38323 ( .C1(n32115), .C2(n32114), .A(n32113), .B(n32112), .ZN(
        n32116) );
  NOR2_X1 U38324 ( .A1(n32118), .A2(n32130), .ZN(n32121) );
  AOI22_X1 U38325 ( .A1(n32121), .A2(n32120), .B1(n32119), .B2(n32118), .ZN(
        n32123) );
  NOR2_X1 U38326 ( .A1(n32125), .A2(n32124), .ZN(n32127) );
  INV_X1 U38327 ( .A(n32129), .ZN(n32133) );
  INV_X1 U38328 ( .A(n34275), .ZN(n32142) );
  XNOR2_X1 U38329 ( .A(n33607), .B(n32142), .ZN(n33359) );
  NAND2_X1 U38330 ( .A1(n36338), .A2(n36340), .ZN(n36328) );
  NAND2_X1 U38331 ( .A1(n36328), .A2(n35010), .ZN(n32143) );
  OAI21_X1 U38332 ( .B1(n38131), .B2(n32143), .A(n38148), .ZN(n32147) );
  NAND2_X1 U38333 ( .A1(n38132), .A2(n38142), .ZN(n38064) );
  NOR2_X1 U38334 ( .A1(n38064), .A2(n35010), .ZN(n32144) );
  AOI22_X1 U38335 ( .A1(n32144), .A2(n36336), .B1(n36338), .B2(n38146), .ZN(
        n32146) );
  NAND3_X1 U38336 ( .A1(n38058), .A2(n611), .A3(n36167), .ZN(n32145) );
  NAND2_X1 U38337 ( .A1(n51012), .A2(n41150), .ZN(n41144) );
  XNOR2_X1 U38338 ( .A(n33711), .B(n36805), .ZN(n32171) );
  OR2_X1 U38339 ( .A1(n32788), .A2(n32785), .ZN(n32160) );
  OAI21_X1 U38340 ( .B1(n32149), .B2(n32160), .A(n32777), .ZN(n32156) );
  NAND2_X1 U38341 ( .A1(n32785), .A2(n31725), .ZN(n32153) );
  AOI21_X1 U38342 ( .B1(n32780), .B2(n32153), .A(n32152), .ZN(n32154) );
  AOI22_X1 U38343 ( .A1(n32780), .A2(n32156), .B1(n32155), .B2(n32154), .ZN(
        n32170) );
  OAI21_X1 U38344 ( .B1(n32794), .B2(n32164), .A(n32282), .ZN(n32159) );
  AOI22_X1 U38345 ( .A1(n32159), .A2(n32284), .B1(n32158), .B2(n32157), .ZN(
        n32169) );
  INV_X1 U38346 ( .A(n32160), .ZN(n32161) );
  NAND3_X1 U38347 ( .A1(n32162), .A2(n32161), .A3(n32284), .ZN(n32168) );
  INV_X1 U38348 ( .A(n32163), .ZN(n32165) );
  XNOR2_X1 U38350 ( .A(n32171), .B(n36811), .ZN(n34037) );
  XNOR2_X1 U38351 ( .A(n35331), .B(n4720), .ZN(n34454) );
  NAND2_X1 U38352 ( .A1(n32175), .A2(n32760), .ZN(n32955) );
  NOR2_X1 U38353 ( .A1(n32955), .A2(n32771), .ZN(n32174) );
  NOR2_X1 U38354 ( .A1(n32172), .A2(n32957), .ZN(n32173) );
  MUX2_X1 U38355 ( .A(n32174), .B(n32173), .S(n32962), .Z(n32181) );
  OAI21_X1 U38356 ( .B1(n32770), .B2(n32957), .A(n3035), .ZN(n32180) );
  INV_X1 U38357 ( .A(n32955), .ZN(n32176) );
  NAND3_X1 U38359 ( .A1(n32176), .A2(n32771), .A3(n32956), .ZN(n32177) );
  NAND2_X1 U38360 ( .A1(n32960), .A2(n32766), .ZN(n32186) );
  NAND3_X1 U38361 ( .A1(n8390), .A2(n32771), .A3(n32761), .ZN(n32184) );
  INV_X1 U38362 ( .A(n32762), .ZN(n32183) );
  NAND2_X1 U38363 ( .A1(n32184), .A2(n32183), .ZN(n32185) );
  INV_X1 U38364 ( .A(n3811), .ZN(n32963) );
  NAND2_X1 U38365 ( .A1(n32185), .A2(n32963), .ZN(n32189) );
  INV_X1 U38366 ( .A(n32186), .ZN(n32187) );
  NAND2_X1 U38367 ( .A1(n32187), .A2(n32957), .ZN(n32188) );
  XNOR2_X1 U38368 ( .A(n33983), .B(n37097), .ZN(n35825) );
  XNOR2_X1 U38369 ( .A(n703), .B(n36812), .ZN(n32224) );
  AOI22_X1 U38370 ( .A1(n5110), .A2(n51103), .B1(n32214), .B2(n32194), .ZN(
        n32198) );
  NAND3_X1 U38371 ( .A1(n51103), .A2(n32194), .A3(n32211), .ZN(n32195) );
  OAI211_X1 U38372 ( .C1(n32198), .C2(n32197), .A(n32196), .B(n32195), .ZN(
        n32200) );
  NOR2_X1 U38373 ( .A1(n32201), .A2(n5109), .ZN(n32205) );
  INV_X1 U38374 ( .A(n32202), .ZN(n32203) );
  AOI22_X1 U38375 ( .A1(n32206), .A2(n32205), .B1(n32204), .B2(n32203), .ZN(
        n32222) );
  NAND2_X1 U38376 ( .A1(n32208), .A2(n32207), .ZN(n32221) );
  AOI21_X1 U38377 ( .B1(n32214), .B2(n5109), .A(n32209), .ZN(n32219) );
  NAND2_X1 U38378 ( .A1(n32211), .A2(n32210), .ZN(n32213) );
  AOI22_X1 U38379 ( .A1(n32214), .A2(n32215), .B1(n32213), .B2(n32212), .ZN(
        n32217) );
  OAI211_X1 U38380 ( .C1(n32219), .C2(n51103), .A(n32217), .B(n32216), .ZN(
        n32220) );
  XNOR2_X1 U38381 ( .A(n33848), .B(n37113), .ZN(n32223) );
  XNOR2_X1 U38382 ( .A(n34455), .B(n32935), .ZN(n32264) );
  INV_X1 U38383 ( .A(n32231), .ZN(n32241) );
  NOR2_X1 U38384 ( .A1(n32241), .A2(n32237), .ZN(n32229) );
  INV_X1 U38385 ( .A(n32257), .ZN(n32228) );
  AOI22_X1 U38386 ( .A1(n32229), .A2(n32228), .B1(n32227), .B2(n32226), .ZN(
        n32262) );
  INV_X1 U38387 ( .A(n32230), .ZN(n32240) );
  OAI211_X1 U38388 ( .C1(n32237), .C2(n32236), .A(n32235), .B(n32234), .ZN(
        n32238) );
  NAND3_X1 U38389 ( .A1(n32241), .A2(n32240), .A3(n32239), .ZN(n32250) );
  NOR2_X1 U38390 ( .A1(n1037), .A2(n32242), .ZN(n32248) );
  NAND2_X1 U38391 ( .A1(n32252), .A2(n32244), .ZN(n32245) );
  NAND4_X1 U38392 ( .A1(n32248), .A2(n32247), .A3(n32246), .A4(n32245), .ZN(
        n32249) );
  AND2_X1 U38393 ( .A1(n32250), .A2(n32249), .ZN(n32261) );
  OAI21_X1 U38394 ( .B1(n32255), .B2(n32254), .A(n32253), .ZN(n32259) );
  AND2_X1 U38395 ( .A1(n32259), .A2(n32258), .ZN(n32260) );
  XNOR2_X1 U38396 ( .A(n33973), .B(n48843), .ZN(n32263) );
  XNOR2_X1 U38397 ( .A(n32264), .B(n32263), .ZN(n32265) );
  XNOR2_X1 U38398 ( .A(n32268), .B(n32267), .ZN(n32269) );
  XNOR2_X1 U38399 ( .A(n32270), .B(n32269), .ZN(n32271) );
  XNOR2_X1 U38400 ( .A(n51739), .B(n32271), .ZN(n32272) );
  XNOR2_X1 U38401 ( .A(n33213), .B(n32274), .ZN(n32275) );
  INV_X1 U38402 ( .A(n34971), .ZN(n35026) );
  XNOR2_X1 U38403 ( .A(n32277), .B(n32276), .ZN(n32278) );
  XNOR2_X1 U38404 ( .A(n34841), .B(n32278), .ZN(n32279) );
  XNOR2_X1 U38405 ( .A(n33722), .B(n47737), .ZN(n33630) );
  XNOR2_X1 U38406 ( .A(n32279), .B(n33630), .ZN(n32281) );
  XNOR2_X1 U38407 ( .A(n32281), .B(n32280), .ZN(n32293) );
  NAND2_X1 U38408 ( .A1(n32286), .A2(n32788), .ZN(n32290) );
  INV_X1 U38409 ( .A(n32794), .ZN(n32283) );
  AOI22_X1 U38410 ( .A1(n32285), .A2(n32284), .B1(n32283), .B2(n32785), .ZN(
        n32289) );
  OAI211_X1 U38412 ( .C1(n32287), .C2(n32793), .A(n32782), .B(n32795), .ZN(
        n32288) );
  XNOR2_X1 U38414 ( .A(n37292), .B(n35088), .ZN(n33398) );
  XNOR2_X1 U38415 ( .A(n33398), .B(n32292), .ZN(n33966) );
  XNOR2_X1 U38416 ( .A(n32293), .B(n33966), .ZN(n32339) );
  NAND2_X1 U38417 ( .A1(n32297), .A2(n32294), .ZN(n32296) );
  AOI22_X1 U38418 ( .A1(n32298), .A2(n32297), .B1(n32296), .B2(n32295), .ZN(
        n32308) );
  NAND2_X1 U38419 ( .A1(n32300), .A2(n32299), .ZN(n32307) );
  INV_X1 U38420 ( .A(n32301), .ZN(n32304) );
  NAND3_X1 U38421 ( .A1(n32304), .A2(n32303), .A3(n32302), .ZN(n32306) );
  XNOR2_X1 U38422 ( .A(n33343), .B(n35633), .ZN(n32309) );
  XNOR2_X1 U38423 ( .A(n32309), .B(n34753), .ZN(n33235) );
  XNOR2_X1 U38424 ( .A(n32310), .B(n49429), .ZN(n37089) );
  XNOR2_X1 U38425 ( .A(n37089), .B(n34041), .ZN(n33101) );
  AOI22_X1 U38427 ( .A1(n32314), .A2(n32313), .B1(n32312), .B2(n32719), .ZN(
        n32323) );
  OAI21_X1 U38428 ( .B1(n32316), .B2(n32716), .A(n32315), .ZN(n32317) );
  OAI21_X1 U38429 ( .B1(n32318), .B2(n32317), .A(n32718), .ZN(n32322) );
  OAI21_X1 U38430 ( .B1(n32729), .B2(n32724), .A(n32457), .ZN(n32319) );
  NAND2_X1 U38431 ( .A1(n32715), .A2(n32319), .ZN(n32320) );
  INV_X1 U38432 ( .A(n32694), .ZN(n32685) );
  INV_X1 U38433 ( .A(n32328), .ZN(n32330) );
  XNOR2_X1 U38434 ( .A(n32691), .B(n32705), .ZN(n32329) );
  OAI211_X1 U38435 ( .C1(n32685), .C2(n32691), .A(n32330), .B(n32329), .ZN(
        n32336) );
  INV_X1 U38436 ( .A(n32333), .ZN(n32334) );
  INV_X1 U38437 ( .A(n36364), .ZN(n36362) );
  INV_X1 U38438 ( .A(n32340), .ZN(n32367) );
  XNOR2_X1 U38439 ( .A(n32342), .B(n32341), .ZN(n32343) );
  XNOR2_X1 U38440 ( .A(n36685), .B(n32343), .ZN(n32365) );
  XNOR2_X1 U38441 ( .A(n32438), .B(n32345), .ZN(n32344) );
  NAND3_X1 U38442 ( .A1(n32344), .A2(n32056), .A3(n32440), .ZN(n32350) );
  OAI21_X1 U38443 ( .B1(n32438), .B2(n32356), .A(n3703), .ZN(n32346) );
  NAND3_X1 U38444 ( .A1(n32359), .A2(n32347), .A3(n32056), .ZN(n32348) );
  INV_X1 U38446 ( .A(n32352), .ZN(n32354) );
  NOR2_X1 U38447 ( .A1(n32440), .A2(n32356), .ZN(n32353) );
  AOI22_X1 U38448 ( .A1(n32446), .A2(n32355), .B1(n32354), .B2(n32353), .ZN(
        n32363) );
  AND2_X1 U38449 ( .A1(n718), .A2(n32439), .ZN(n32358) );
  AND3_X1 U38450 ( .A1(n32438), .A2(n32440), .A3(n32356), .ZN(n32357) );
  NAND2_X1 U38452 ( .A1(n32360), .A2(n3703), .ZN(n32361) );
  XNOR2_X1 U38453 ( .A(n37261), .B(n4855), .ZN(n33902) );
  XNOR2_X1 U38454 ( .A(n32365), .B(n33902), .ZN(n32366) );
  XNOR2_X1 U38455 ( .A(n32367), .B(n32366), .ZN(n32371) );
  INV_X1 U38456 ( .A(n34400), .ZN(n32368) );
  XNOR2_X1 U38457 ( .A(n37252), .B(n32368), .ZN(n32369) );
  XNOR2_X1 U38458 ( .A(n34128), .B(n32369), .ZN(n32370) );
  XNOR2_X1 U38459 ( .A(n32371), .B(n32370), .ZN(n32434) );
  XNOR2_X1 U38460 ( .A(n32372), .B(n36869), .ZN(n33763) );
  INV_X1 U38461 ( .A(n32373), .ZN(n32376) );
  NOR2_X1 U38462 ( .A1(n32376), .A2(n32375), .ZN(n32393) );
  OAI21_X1 U38463 ( .B1(n32378), .B2(n32377), .A(n32389), .ZN(n32384) );
  NAND2_X1 U38464 ( .A1(n32380), .A2(n32843), .ZN(n32382) );
  NAND3_X1 U38465 ( .A1(n32382), .A2(n32841), .A3(n32381), .ZN(n32383) );
  NAND2_X1 U38466 ( .A1(n32384), .A2(n32383), .ZN(n32392) );
  NOR2_X1 U38467 ( .A1(n32844), .A2(n32843), .ZN(n32388) );
  MUX2_X1 U38468 ( .A(n32386), .B(n32385), .S(n32841), .Z(n32387) );
  NAND2_X1 U38469 ( .A1(n32388), .A2(n32387), .ZN(n32391) );
  NAND3_X1 U38470 ( .A1(n32837), .A2(n32389), .A3(n32844), .ZN(n32390) );
  XNOR2_X1 U38471 ( .A(n35829), .B(n375), .ZN(n34492) );
  NAND2_X1 U38472 ( .A1(n32396), .A2(n51520), .ZN(n32397) );
  NAND2_X1 U38473 ( .A1(n32400), .A2(n32399), .ZN(n32406) );
  AND2_X1 U38474 ( .A1(n32402), .A2(n51519), .ZN(n32403) );
  OAI211_X1 U38475 ( .C1(n32404), .C2(n32403), .A(n32408), .B(n32407), .ZN(
        n32405) );
  XNOR2_X1 U38476 ( .A(n34492), .B(n34811), .ZN(n32432) );
  BUF_X2 U38477 ( .A(n33566), .Z(n36939) );
  NAND2_X1 U38478 ( .A1(n8536), .A2(n32829), .ZN(n32419) );
  INV_X1 U38479 ( .A(n32415), .ZN(n32418) );
  AOI22_X1 U38480 ( .A1(n32419), .A2(n32418), .B1(n32417), .B2(n32416), .ZN(
        n32431) );
  NOR2_X1 U38481 ( .A1(n32421), .A2(n32420), .ZN(n32422) );
  OAI211_X1 U38482 ( .C1(n32423), .C2(n32827), .A(n32422), .B(n32426), .ZN(
        n32430) );
  XNOR2_X1 U38483 ( .A(n36939), .B(n35830), .ZN(n34824) );
  XNOR2_X1 U38484 ( .A(n32432), .B(n34824), .ZN(n37053) );
  XNOR2_X1 U38485 ( .A(n37053), .B(n33763), .ZN(n32433) );
  OAI211_X1 U38486 ( .C1(n32444), .C2(n718), .A(n32443), .B(n32442), .ZN(
        n32450) );
  NAND3_X1 U38487 ( .A1(n32447), .A2(n32446), .A3(n723), .ZN(n32448) );
  NOR2_X1 U38488 ( .A1(n32452), .A2(n718), .ZN(n32454) );
  OAI21_X1 U38489 ( .B1(n32455), .B2(n32454), .A(n32453), .ZN(n32456) );
  NOR2_X1 U38490 ( .A1(n32458), .A2(n32457), .ZN(n32459) );
  AOI22_X1 U38491 ( .A1(n32725), .A2(n32460), .B1(n32459), .B2(n31648), .ZN(
        n32470) );
  NAND3_X1 U38492 ( .A1(n32725), .A2(n32719), .A3(n32463), .ZN(n32461) );
  OAI211_X1 U38493 ( .C1(n32725), .C2(n32463), .A(n32462), .B(n32461), .ZN(
        n32469) );
  INV_X1 U38496 ( .A(n32471), .ZN(n32494) );
  INV_X1 U38497 ( .A(n32474), .ZN(n32475) );
  AOI22_X1 U38498 ( .A1(n32477), .A2(n32486), .B1(n32476), .B2(n32475), .ZN(
        n32493) );
  NOR2_X1 U38499 ( .A1(n32479), .A2(n32478), .ZN(n32482) );
  NAND2_X1 U38500 ( .A1(n32486), .A2(n32485), .ZN(n32488) );
  XNOR2_X1 U38502 ( .A(n32495), .B(n5016), .ZN(n32496) );
  XNOR2_X1 U38503 ( .A(n32497), .B(n32496), .ZN(n32498) );
  XNOR2_X1 U38504 ( .A(n34835), .B(n32498), .ZN(n32499) );
  XNOR2_X1 U38505 ( .A(n32499), .B(n37067), .ZN(n32519) );
  NAND2_X1 U38506 ( .A1(n32501), .A2(n32500), .ZN(n32505) );
  AOI21_X1 U38507 ( .B1(n32511), .B2(n32509), .A(n32508), .ZN(n32513) );
  XNOR2_X1 U38508 ( .A(n33911), .B(n36672), .ZN(n32517) );
  XNOR2_X1 U38509 ( .A(n33470), .B(n32517), .ZN(n32518) );
  XNOR2_X1 U38510 ( .A(n32519), .B(n32518), .ZN(n32522) );
  XNOR2_X1 U38511 ( .A(n34382), .B(n32520), .ZN(n32755) );
  XNOR2_X1 U38512 ( .A(n34020), .B(n32755), .ZN(n32521) );
  XNOR2_X1 U38513 ( .A(n32522), .B(n32521), .ZN(n32523) );
  XNOR2_X1 U38514 ( .A(n34012), .B(n32523), .ZN(n32678) );
  NAND2_X1 U38515 ( .A1(n38002), .A2(n5872), .ZN(n38188) );
  OAI21_X1 U38516 ( .B1(n32967), .B2(n32524), .A(n32763), .ZN(n32526) );
  NOR2_X1 U38518 ( .A1(n32771), .A2(n32960), .ZN(n32528) );
  AND2_X1 U38519 ( .A1(n32766), .A2(n32760), .ZN(n32527) );
  OAI21_X1 U38520 ( .B1(n32956), .B2(n32528), .A(n32527), .ZN(n32531) );
  AND2_X1 U38521 ( .A1(n32761), .A2(n32960), .ZN(n32958) );
  NAND2_X1 U38522 ( .A1(n32529), .A2(n32958), .ZN(n32530) );
  NOR2_X1 U38523 ( .A1(n32532), .A2(n32957), .ZN(n32534) );
  AND2_X1 U38524 ( .A1(n32766), .A2(n32965), .ZN(n32535) );
  OAI21_X1 U38525 ( .B1(n32967), .B2(n32535), .A(n32761), .ZN(n32536) );
  XNOR2_X1 U38526 ( .A(n34503), .B(n34413), .ZN(n34247) );
  OAI211_X1 U38527 ( .C1(n32633), .C2(n32909), .A(n32895), .B(n32540), .ZN(
        n32541) );
  NOR2_X1 U38528 ( .A1(n32634), .A2(n32916), .ZN(n32542) );
  AOI22_X1 U38529 ( .A1(n32636), .A2(n32547), .B1(n32639), .B2(n32542), .ZN(
        n32550) );
  NOR2_X1 U38530 ( .A1(n32900), .A2(n32909), .ZN(n32543) );
  NAND2_X1 U38531 ( .A1(n32634), .A2(n32895), .ZN(n32546) );
  OAI211_X1 U38532 ( .C1(n32548), .C2(n32634), .A(n32547), .B(n32546), .ZN(
        n32549) );
  XNOR2_X1 U38533 ( .A(n42102), .B(n1224), .ZN(n32552) );
  XNOR2_X1 U38534 ( .A(n32553), .B(n32552), .ZN(n32554) );
  XNOR2_X1 U38535 ( .A(n32554), .B(n42592), .ZN(n32555) );
  XNOR2_X1 U38536 ( .A(n37303), .B(n32555), .ZN(n32556) );
  XNOR2_X1 U38537 ( .A(n34247), .B(n32556), .ZN(n32584) );
  INV_X1 U38538 ( .A(n32557), .ZN(n32563) );
  OAI211_X1 U38539 ( .C1(n32561), .C2(n32560), .A(n854), .B(n32558), .ZN(
        n32562) );
  NAND2_X1 U38540 ( .A1(n32563), .A2(n32562), .ZN(n32582) );
  INV_X1 U38541 ( .A(n32570), .ZN(n32564) );
  NAND2_X1 U38542 ( .A1(n32565), .A2(n32564), .ZN(n32567) );
  NAND2_X1 U38543 ( .A1(n32567), .A2(n32566), .ZN(n32581) );
  INV_X1 U38544 ( .A(n32568), .ZN(n32572) );
  AOI22_X1 U38545 ( .A1(n32572), .A2(n32571), .B1(n32570), .B2(n32569), .ZN(
        n32580) );
  NAND3_X1 U38546 ( .A1(n32575), .A2(n32574), .A3(n32573), .ZN(n32578) );
  INV_X1 U38547 ( .A(n32576), .ZN(n32577) );
  AND2_X1 U38548 ( .A1(n32578), .A2(n32577), .ZN(n32579) );
  XNOR2_X1 U38550 ( .A(n32584), .B(n32583), .ZN(n32585) );
  XNOR2_X1 U38551 ( .A(n51493), .B(n35105), .ZN(n35659) );
  INV_X1 U38552 ( .A(n32976), .ZN(n32591) );
  INV_X1 U38553 ( .A(n32989), .ZN(n32592) );
  NAND3_X1 U38554 ( .A1(n32592), .A2(n32591), .A3(n32590), .ZN(n32593) );
  AND2_X1 U38555 ( .A1(n32594), .A2(n32593), .ZN(n32604) );
  OAI21_X1 U38556 ( .B1(n32597), .B2(n32596), .A(n32595), .ZN(n32603) );
  INV_X1 U38557 ( .A(n32598), .ZN(n32599) );
  OAI211_X1 U38558 ( .C1(n32601), .C2(n32600), .A(n32599), .B(n32987), .ZN(
        n32602) );
  XNOR2_X1 U38559 ( .A(n33142), .B(n517), .ZN(n32605) );
  XNOR2_X2 U38561 ( .A(n32607), .B(n34611), .ZN(n38005) );
  XNOR2_X1 U38562 ( .A(n36764), .B(n34896), .ZN(n32626) );
  NAND2_X1 U38563 ( .A1(n32609), .A2(n32608), .ZN(n32612) );
  NAND2_X1 U38564 ( .A1(n32610), .A2(n32616), .ZN(n32611) );
  AOI21_X1 U38565 ( .B1(n32613), .B2(n32612), .A(n32611), .ZN(n32625) );
  INV_X1 U38566 ( .A(n32614), .ZN(n32615) );
  XNOR2_X1 U38567 ( .A(n32628), .B(n32627), .ZN(n34889) );
  XNOR2_X1 U38568 ( .A(n34369), .B(n4639), .ZN(n34157) );
  NOR2_X1 U38569 ( .A1(n32915), .A2(n32895), .ZN(n32629) );
  OAI21_X1 U38570 ( .B1(n32922), .B2(n32629), .A(n32899), .ZN(n32643) );
  NAND2_X1 U38571 ( .A1(n32634), .A2(n32894), .ZN(n32630) );
  AND2_X1 U38572 ( .A1(n32631), .A2(n32630), .ZN(n32642) );
  AND2_X1 U38573 ( .A1(n32908), .A2(n32632), .ZN(n32637) );
  AND2_X1 U38574 ( .A1(n32634), .A2(n32633), .ZN(n32635) );
  AOI22_X1 U38575 ( .A1(n32637), .A2(n32636), .B1(n32899), .B2(n32635), .ZN(
        n32641) );
  XNOR2_X1 U38577 ( .A(n37324), .B(n36999), .ZN(n33953) );
  XNOR2_X1 U38578 ( .A(n33953), .B(n35678), .ZN(n32654) );
  OAI21_X1 U38579 ( .B1(n32865), .B2(n33041), .A(n32645), .ZN(n32646) );
  NAND3_X1 U38581 ( .A1(n32646), .A2(n32882), .A3(n32868), .ZN(n32653) );
  AND2_X1 U38582 ( .A1(n32882), .A2(n32876), .ZN(n33024) );
  INV_X1 U38583 ( .A(n32887), .ZN(n32648) );
  OAI21_X1 U38584 ( .B1(n8544), .B2(n33024), .A(n32648), .ZN(n32647) );
  OAI211_X1 U38585 ( .C1(n719), .C2(n8544), .A(n32647), .B(n33041), .ZN(n32652) );
  NAND2_X1 U38586 ( .A1(n5498), .A2(n33035), .ZN(n32651) );
  NAND2_X1 U38587 ( .A1(n33026), .A2(n32876), .ZN(n32886) );
  NOR2_X1 U38588 ( .A1(n32886), .A2(n32648), .ZN(n32649) );
  NOR2_X1 U38589 ( .A1(n32649), .A2(n32877), .ZN(n32650) );
  XNOR2_X1 U38590 ( .A(n32654), .B(n34625), .ZN(n37130) );
  XNOR2_X1 U38591 ( .A(n32655), .B(n37130), .ZN(n32677) );
  INV_X1 U38592 ( .A(n37318), .ZN(n32656) );
  XNOR2_X1 U38593 ( .A(n32658), .B(n32657), .ZN(n32659) );
  OAI21_X1 U38594 ( .B1(n32664), .B2(n32663), .A(n32662), .ZN(n32670) );
  NAND3_X1 U38595 ( .A1(n32667), .A2(n32666), .A3(n32665), .ZN(n32668) );
  XNOR2_X1 U38596 ( .A(n32673), .B(n33943), .ZN(n32674) );
  XNOR2_X1 U38597 ( .A(n36766), .B(n32674), .ZN(n32675) );
  XNOR2_X1 U38598 ( .A(n35136), .B(n32675), .ZN(n32676) );
  XNOR2_X1 U38599 ( .A(n32677), .B(n32676), .ZN(n36359) );
  NAND3_X1 U38600 ( .A1(n38001), .A2(n36359), .A3(n35028), .ZN(n38179) );
  NAND2_X1 U38601 ( .A1(n38006), .A2(n35028), .ZN(n38012) );
  OR2_X1 U38602 ( .A1(n38014), .A2(n38012), .ZN(n38178) );
  NAND2_X1 U38603 ( .A1(n38184), .A2(n36362), .ZN(n38024) );
  NOR2_X1 U38605 ( .A1(n38190), .A2(n38188), .ZN(n38000) );
  INV_X1 U38606 ( .A(n38005), .ZN(n38019) );
  OAI21_X1 U38608 ( .B1(n38000), .B2(n32679), .A(n38192), .ZN(n32683) );
  NOR2_X1 U38609 ( .A1(n37997), .A2(n5872), .ZN(n38185) );
  NAND2_X1 U38610 ( .A1(n38019), .A2(n34971), .ZN(n36361) );
  OAI21_X1 U38611 ( .B1(n36364), .B2(n38018), .A(n38015), .ZN(n32680) );
  NOR2_X1 U38612 ( .A1(n36361), .A2(n32680), .ZN(n32681) );
  NOR2_X1 U38613 ( .A1(n38185), .A2(n32681), .ZN(n32682) );
  NAND2_X1 U38614 ( .A1(n32685), .A2(n1988), .ZN(n32686) );
  AND2_X1 U38615 ( .A1(n32687), .A2(n32686), .ZN(n32713) );
  INV_X1 U38616 ( .A(n32688), .ZN(n32689) );
  NOR2_X1 U38617 ( .A1(n32689), .A2(n32705), .ZN(n32698) );
  INV_X1 U38618 ( .A(n32690), .ZN(n32697) );
  NAND2_X1 U38619 ( .A1(n32705), .A2(n32691), .ZN(n32693) );
  NAND2_X1 U38620 ( .A1(n32694), .A2(n32693), .ZN(n32695) );
  AOI22_X1 U38621 ( .A1(n32698), .A2(n32697), .B1(n32696), .B2(n32695), .ZN(
        n32712) );
  INV_X1 U38622 ( .A(n32699), .ZN(n32703) );
  OAI21_X1 U38623 ( .B1(n32704), .B2(n52182), .A(n32700), .ZN(n32702) );
  NAND2_X1 U38624 ( .A1(n32703), .A2(n32702), .ZN(n32711) );
  INV_X1 U38625 ( .A(n32704), .ZN(n32709) );
  OAI211_X1 U38626 ( .C1(n32709), .C2(n32708), .A(n32707), .B(n32706), .ZN(
        n32710) );
  OAI211_X1 U38627 ( .C1(n32720), .C2(n32719), .A(n32718), .B(n32717), .ZN(
        n32723) );
  AND3_X1 U38628 ( .A1(n32723), .A2(n32722), .A3(n32721), .ZN(n32735) );
  INV_X1 U38629 ( .A(n34491), .ZN(n33502) );
  XNOR2_X1 U38630 ( .A(n51702), .B(n35501), .ZN(n33764) );
  XNOR2_X1 U38631 ( .A(n33889), .B(n35833), .ZN(n35493) );
  XNOR2_X1 U38632 ( .A(n35493), .B(n32737), .ZN(n32748) );
  XNOR2_X1 U38633 ( .A(n43252), .B(n32738), .ZN(n32739) );
  XNOR2_X1 U38634 ( .A(n34400), .B(n32739), .ZN(n32740) );
  XNOR2_X1 U38635 ( .A(n32740), .B(n37252), .ZN(n32743) );
  INV_X1 U38636 ( .A(n32741), .ZN(n35588) );
  XNOR2_X1 U38637 ( .A(n35588), .B(n47268), .ZN(n32742) );
  XNOR2_X1 U38638 ( .A(n32743), .B(n35033), .ZN(n32746) );
  INV_X1 U38639 ( .A(n32744), .ZN(n32745) );
  XNOR2_X1 U38640 ( .A(n32746), .B(n32745), .ZN(n32747) );
  XNOR2_X1 U38641 ( .A(n34219), .B(n33759), .ZN(n32750) );
  XNOR2_X1 U38642 ( .A(n36932), .B(n4676), .ZN(n32749) );
  XNOR2_X1 U38643 ( .A(n32750), .B(n32749), .ZN(n35612) );
  XNOR2_X1 U38644 ( .A(n35048), .B(n33470), .ZN(n33078) );
  INV_X1 U38645 ( .A(n33078), .ZN(n32751) );
  XNOR2_X1 U38646 ( .A(n32752), .B(n40104), .ZN(n32753) );
  XNOR2_X1 U38647 ( .A(n52117), .B(n32753), .ZN(n32754) );
  XNOR2_X1 U38648 ( .A(n32755), .B(n32754), .ZN(n32756) );
  XNOR2_X1 U38649 ( .A(n32757), .B(n32756), .ZN(n32758) );
  XNOR2_X1 U38650 ( .A(n37063), .B(n33194), .ZN(n32802) );
  NAND3_X1 U38651 ( .A1(n32763), .A2(n32762), .A3(n3035), .ZN(n32764) );
  NOR2_X1 U38652 ( .A1(n32964), .A2(n32962), .ZN(n32769) );
  AND2_X1 U38653 ( .A1(n3754), .A2(n32960), .ZN(n32768) );
  AOI22_X1 U38654 ( .A1(n32769), .A2(n32768), .B1(n32767), .B2(n32766), .ZN(
        n32776) );
  OAI21_X1 U38655 ( .B1(n32773), .B2(n32772), .A(n32771), .ZN(n32774) );
  OAI21_X1 U38656 ( .B1(n32779), .B2(n32778), .A(n32777), .ZN(n32781) );
  NAND2_X1 U38657 ( .A1(n32781), .A2(n32780), .ZN(n32800) );
  NAND3_X1 U38658 ( .A1(n32785), .A2(n32788), .A3(n32784), .ZN(n32786) );
  NOR2_X1 U38659 ( .A1(n32787), .A2(n32786), .ZN(n32792) );
  AND2_X1 U38660 ( .A1(n32788), .A2(n31725), .ZN(n32790) );
  NAND2_X1 U38661 ( .A1(n32794), .A2(n32793), .ZN(n32796) );
  XNOR2_X1 U38662 ( .A(n33550), .B(n34156), .ZN(n35478) );
  XNOR2_X1 U38663 ( .A(n35478), .B(n33942), .ZN(n32805) );
  XNOR2_X1 U38664 ( .A(n36761), .B(n35283), .ZN(n32804) );
  XNOR2_X1 U38665 ( .A(n32804), .B(n32805), .ZN(n32813) );
  XNOR2_X1 U38666 ( .A(n32807), .B(n32806), .ZN(n32808) );
  XNOR2_X1 U38667 ( .A(n35683), .B(n32808), .ZN(n32809) );
  XNOR2_X1 U38668 ( .A(n35124), .B(n32809), .ZN(n32810) );
  XNOR2_X1 U38669 ( .A(n32811), .B(n32810), .ZN(n32812) );
  XNOR2_X1 U38670 ( .A(n32812), .B(n32813), .ZN(n32855) );
  INV_X1 U38671 ( .A(n32814), .ZN(n32818) );
  AOI21_X1 U38672 ( .B1(n32816), .B2(n51618), .A(n32821), .ZN(n32817) );
  NAND2_X1 U38673 ( .A1(n32818), .A2(n32817), .ZN(n32835) );
  INV_X1 U38674 ( .A(n32819), .ZN(n32820) );
  NAND2_X1 U38675 ( .A1(n32824), .A2(n32823), .ZN(n32826) );
  NAND2_X1 U38676 ( .A1(n32826), .A2(n32825), .ZN(n32834) );
  INV_X1 U38677 ( .A(n32827), .ZN(n32833) );
  OAI21_X1 U38678 ( .B1(n32830), .B2(n32829), .A(n32828), .ZN(n32832) );
  NAND2_X1 U38679 ( .A1(n32841), .A2(n32840), .ZN(n32842) );
  NAND2_X1 U38680 ( .A1(n32843), .A2(n32842), .ZN(n32845) );
  NAND2_X1 U38681 ( .A1(n32845), .A2(n32844), .ZN(n32847) );
  NAND4_X1 U38682 ( .A1(n32849), .A2(n32848), .A3(n32847), .A4(n32846), .ZN(
        n32854) );
  AOI21_X1 U38683 ( .B1(n32852), .B2(n32851), .A(n32850), .ZN(n32853) );
  AND2_X1 U38684 ( .A1(n38570), .A2(n38561), .ZN(n33060) );
  INV_X1 U38685 ( .A(n32856), .ZN(n32857) );
  XNOR2_X1 U38686 ( .A(n703), .B(n32857), .ZN(n32858) );
  XNOR2_X1 U38687 ( .A(n37113), .B(n32858), .ZN(n36808) );
  XNOR2_X1 U38688 ( .A(n35325), .B(n32859), .ZN(n33515) );
  INV_X1 U38689 ( .A(n32860), .ZN(n33372) );
  XNOR2_X1 U38690 ( .A(n33515), .B(n33372), .ZN(n33707) );
  INV_X1 U38691 ( .A(n32870), .ZN(n32861) );
  OAI21_X1 U38692 ( .B1(n32861), .B2(n32867), .A(n33026), .ZN(n32864) );
  NOR3_X1 U38693 ( .A1(n33026), .A2(n33041), .A3(n719), .ZN(n32862) );
  OAI211_X1 U38694 ( .C1(n32865), .C2(n32864), .A(n33032), .B(n32863), .ZN(
        n32866) );
  INV_X1 U38695 ( .A(n32866), .ZN(n32893) );
  OR2_X1 U38696 ( .A1(n33026), .A2(n32867), .ZN(n32869) );
  NOR2_X1 U38697 ( .A1(n32869), .A2(n33034), .ZN(n32873) );
  NOR2_X1 U38699 ( .A1(n32870), .A2(n32869), .ZN(n32871) );
  NAND4_X1 U38701 ( .A1(n8544), .A2(n33034), .A3(n32874), .A4(n719), .ZN(
        n32875) );
  INV_X1 U38702 ( .A(n32877), .ZN(n33039) );
  AOI21_X1 U38703 ( .B1(n32875), .B2(n33039), .A(n32882), .ZN(n32881) );
  NOR2_X1 U38704 ( .A1(n32881), .A2(n32880), .ZN(n32891) );
  NAND2_X1 U38705 ( .A1(n33026), .A2(n32882), .ZN(n32884) );
  OAI21_X1 U38706 ( .B1(n32885), .B2(n32884), .A(n32883), .ZN(n32889) );
  OAI21_X1 U38707 ( .B1(n32887), .B2(n32886), .A(n8544), .ZN(n32888) );
  NAND2_X1 U38708 ( .A1(n32889), .A2(n32888), .ZN(n32890) );
  AND3_X1 U38710 ( .A1(n32895), .A2(n32900), .A3(n32909), .ZN(n32897) );
  NAND4_X1 U38711 ( .A1(n32899), .A2(n6269), .A3(n32915), .A4(n32909), .ZN(
        n32903) );
  NAND4_X1 U38712 ( .A1(n32901), .A2(n32915), .A3(n6269), .A4(n32900), .ZN(
        n32902) );
  NAND2_X1 U38713 ( .A1(n32903), .A2(n32902), .ZN(n32904) );
  OR2_X1 U38714 ( .A1(n32909), .A2(n32908), .ZN(n32910) );
  AOI21_X1 U38715 ( .B1(n32911), .B2(n32910), .A(n32915), .ZN(n32914) );
  NOR2_X1 U38716 ( .A1(n32918), .A2(n32912), .ZN(n32913) );
  NOR2_X1 U38717 ( .A1(n32914), .A2(n32913), .ZN(n32926) );
  INV_X1 U38718 ( .A(n32919), .ZN(n32920) );
  NAND2_X1 U38719 ( .A1(n32921), .A2(n32920), .ZN(n32925) );
  XNOR2_X1 U38720 ( .A(n51497), .B(n34275), .ZN(n32928) );
  XNOR2_X1 U38721 ( .A(n32928), .B(n33608), .ZN(n33095) );
  XNOR2_X1 U38722 ( .A(n32929), .B(n37108), .ZN(n34101) );
  INV_X1 U38723 ( .A(n32930), .ZN(n32931) );
  XNOR2_X1 U38724 ( .A(n32931), .B(n4653), .ZN(n32932) );
  XNOR2_X1 U38725 ( .A(n35070), .B(n32932), .ZN(n32933) );
  XNOR2_X1 U38726 ( .A(n32934), .B(n32933), .ZN(n32936) );
  XNOR2_X2 U38727 ( .A(n33848), .B(n32935), .ZN(n37096) );
  XNOR2_X1 U38728 ( .A(n37096), .B(n32936), .ZN(n32937) );
  XNOR2_X1 U38729 ( .A(n34101), .B(n32937), .ZN(n32938) );
  XNOR2_X1 U38730 ( .A(n42339), .B(n4589), .ZN(n32939) );
  XNOR2_X1 U38731 ( .A(n32940), .B(n32939), .ZN(n32942) );
  XNOR2_X1 U38732 ( .A(n32942), .B(n32941), .ZN(n32945) );
  OAI21_X1 U38733 ( .B1(n32943), .B2(n32944), .A(n32945), .ZN(n32950) );
  INV_X1 U38734 ( .A(n32943), .ZN(n32948) );
  INV_X1 U38735 ( .A(n32944), .ZN(n32947) );
  INV_X1 U38736 ( .A(n32945), .ZN(n32946) );
  NAND3_X1 U38737 ( .A1(n32948), .A2(n32947), .A3(n32946), .ZN(n32949) );
  NAND2_X1 U38738 ( .A1(n32950), .A2(n32949), .ZN(n32951) );
  XNOR2_X1 U38739 ( .A(n34841), .B(n32951), .ZN(n32953) );
  XNOR2_X1 U38740 ( .A(n32953), .B(n33386), .ZN(n32954) );
  XNOR2_X1 U38741 ( .A(n33343), .B(n35543), .ZN(n34052) );
  XNOR2_X1 U38742 ( .A(n32954), .B(n34052), .ZN(n32973) );
  NAND2_X1 U38743 ( .A1(n32955), .A2(n32964), .ZN(n32959) );
  INV_X1 U38744 ( .A(n32956), .ZN(n32968) );
  AOI22_X1 U38745 ( .A1(n32959), .A2(n32968), .B1(n32958), .B2(n32957), .ZN(
        n32972) );
  NAND4_X1 U38746 ( .A1(n32963), .A2(n32962), .A3(n32961), .A4(n32960), .ZN(
        n32971) );
  NAND3_X1 U38747 ( .A1(n2473), .A2(n32965), .A3(n32964), .ZN(n32970) );
  OAI21_X1 U38748 ( .B1(n32968), .B2(n32967), .A(n32966), .ZN(n32969) );
  NAND4_X2 U38749 ( .A1(n32972), .A2(n32969), .A3(n32970), .A4(n32971), .ZN(
        n37086) );
  XNOR2_X1 U38750 ( .A(n32973), .B(n36714), .ZN(n33001) );
  XNOR2_X1 U38751 ( .A(n35086), .B(n35085), .ZN(n36704) );
  NAND2_X1 U38752 ( .A1(n32975), .A2(n32974), .ZN(n32979) );
  INV_X1 U38753 ( .A(n32981), .ZN(n32982) );
  NOR2_X1 U38754 ( .A1(n32983), .A2(n32982), .ZN(n32984) );
  NAND2_X1 U38755 ( .A1(n32987), .A2(n32986), .ZN(n32993) );
  OAI211_X1 U38756 ( .C1(n52046), .C2(n32990), .A(n32989), .B(n32988), .ZN(
        n32992) );
  XNOR2_X1 U38757 ( .A(n32996), .B(n35537), .ZN(n35090) );
  XNOR2_X1 U38758 ( .A(n36704), .B(n35090), .ZN(n32999) );
  XNOR2_X1 U38759 ( .A(n35095), .B(n32997), .ZN(n33526) );
  INV_X1 U38760 ( .A(n31923), .ZN(n35080) );
  XNOR2_X1 U38761 ( .A(n33526), .B(n35080), .ZN(n33111) );
  INV_X1 U38762 ( .A(n33111), .ZN(n32998) );
  XNOR2_X1 U38763 ( .A(n32999), .B(n32998), .ZN(n33000) );
  INV_X1 U38764 ( .A(n35104), .ZN(n33046) );
  NAND2_X1 U38765 ( .A1(n33003), .A2(n33002), .ZN(n33012) );
  AOI22_X1 U38766 ( .A1(n33008), .A2(n33007), .B1(n33006), .B2(n33005), .ZN(
        n33010) );
  INV_X1 U38767 ( .A(n33024), .ZN(n33040) );
  INV_X1 U38768 ( .A(n33025), .ZN(n33027) );
  NAND2_X1 U38769 ( .A1(n33030), .A2(n33041), .ZN(n33031) );
  NAND2_X1 U38770 ( .A1(n33032), .A2(n33031), .ZN(n33033) );
  NAND2_X1 U38771 ( .A1(n33033), .A2(n33034), .ZN(n33045) );
  XNOR2_X1 U38772 ( .A(n33034), .B(n33041), .ZN(n33038) );
  OAI211_X1 U38773 ( .C1(n33038), .C2(n719), .A(n8544), .B(n33037), .ZN(n33044) );
  OAI21_X1 U38774 ( .B1(n33041), .B2(n33040), .A(n33039), .ZN(n33042) );
  NAND2_X1 U38775 ( .A1(n5498), .A2(n33042), .ZN(n33043) );
  XNOR2_X1 U38776 ( .A(n35285), .B(n33046), .ZN(n33645) );
  XNOR2_X1 U38777 ( .A(n35105), .B(n35115), .ZN(n33047) );
  XNOR2_X1 U38778 ( .A(n33047), .B(n33938), .ZN(n33048) );
  XNOR2_X1 U38779 ( .A(n34163), .B(n35468), .ZN(n33267) );
  XNOR2_X1 U38780 ( .A(n33050), .B(n33049), .ZN(n33051) );
  XNOR2_X1 U38781 ( .A(n33052), .B(n33051), .ZN(n33054) );
  XNOR2_X1 U38782 ( .A(n33054), .B(n33053), .ZN(n33055) );
  XNOR2_X1 U38783 ( .A(n2131), .B(n33055), .ZN(n33056) );
  INV_X1 U38784 ( .A(n36832), .ZN(n37133) );
  NAND3_X1 U38785 ( .A1(n33062), .A2(n38561), .A3(n6869), .ZN(n33058) );
  INV_X1 U38786 ( .A(n38200), .ZN(n36098) );
  AND2_X1 U38787 ( .A1(n591), .A2(n36098), .ZN(n36106) );
  AOI22_X1 U38788 ( .A1(n33060), .A2(n38566), .B1(n33059), .B2(n36106), .ZN(
        n33066) );
  INV_X1 U38789 ( .A(n38575), .ZN(n35151) );
  NAND3_X1 U38790 ( .A1(n38565), .A2(n7759), .A3(n38201), .ZN(n33061) );
  NAND2_X1 U38791 ( .A1(n33063), .A2(n38196), .ZN(n33065) );
  NAND3_X1 U38792 ( .A1(n38567), .A2(n38576), .A3(n38204), .ZN(n35713) );
  NAND2_X1 U38793 ( .A1(n33067), .A2(n38561), .ZN(n35706) );
  AOI21_X1 U38794 ( .B1(n36104), .B2(n6869), .A(n35706), .ZN(n33068) );
  XNOR2_X1 U38795 ( .A(n34141), .B(n5016), .ZN(n35513) );
  XNOR2_X1 U38796 ( .A(n35513), .B(n33070), .ZN(n33076) );
  XNOR2_X1 U38797 ( .A(n33072), .B(n33071), .ZN(n33073) );
  XNOR2_X1 U38798 ( .A(n52117), .B(n33073), .ZN(n33074) );
  XNOR2_X1 U38799 ( .A(n33074), .B(n34553), .ZN(n33075) );
  XNOR2_X1 U38800 ( .A(n33076), .B(n33075), .ZN(n33080) );
  XNOR2_X1 U38801 ( .A(n36930), .B(n37067), .ZN(n33077) );
  XNOR2_X1 U38802 ( .A(n33077), .B(n34219), .ZN(n36677) );
  XNOR2_X1 U38803 ( .A(n36677), .B(n33078), .ZN(n33079) );
  XNOR2_X1 U38804 ( .A(n33080), .B(n33079), .ZN(n33083) );
  XNOR2_X1 U38805 ( .A(n35265), .B(n42297), .ZN(n33081) );
  XNOR2_X1 U38806 ( .A(n33081), .B(n51664), .ZN(n33082) );
  XNOR2_X1 U38807 ( .A(n34230), .B(n33083), .ZN(n33174) );
  XNOR2_X1 U38808 ( .A(n37095), .B(n37096), .ZN(n33084) );
  XNOR2_X1 U38809 ( .A(n34343), .B(n33084), .ZN(n33094) );
  XNOR2_X1 U38810 ( .A(n34760), .B(n35334), .ZN(n36971) );
  XNOR2_X1 U38811 ( .A(n36971), .B(n33085), .ZN(n33092) );
  INV_X1 U38812 ( .A(n36293), .ZN(n33088) );
  XNOR2_X1 U38813 ( .A(n33086), .B(n48843), .ZN(n33087) );
  XNOR2_X1 U38814 ( .A(n33088), .B(n33087), .ZN(n33089) );
  XNOR2_X1 U38815 ( .A(n703), .B(n33089), .ZN(n33090) );
  XNOR2_X1 U38816 ( .A(n37113), .B(n33090), .ZN(n33091) );
  XNOR2_X1 U38817 ( .A(n33092), .B(n33091), .ZN(n33093) );
  XNOR2_X1 U38818 ( .A(n33094), .B(n33093), .ZN(n33096) );
  INV_X1 U38819 ( .A(n33097), .ZN(n34842) );
  XNOR2_X1 U38820 ( .A(n34842), .B(n36792), .ZN(n33099) );
  XNOR2_X1 U38821 ( .A(n2129), .B(n35633), .ZN(n33098) );
  XNOR2_X1 U38822 ( .A(n33099), .B(n33098), .ZN(n33100) );
  XNOR2_X1 U38823 ( .A(n33101), .B(n33100), .ZN(n33102) );
  XNOR2_X1 U38824 ( .A(n33102), .B(n36714), .ZN(n33113) );
  XNOR2_X1 U38825 ( .A(n35536), .B(n44015), .ZN(n33103) );
  XNOR2_X1 U38826 ( .A(n33103), .B(n35537), .ZN(n37079) );
  XNOR2_X1 U38827 ( .A(n42339), .B(n34742), .ZN(n33106) );
  XNOR2_X1 U38828 ( .A(n33106), .B(n33105), .ZN(n33107) );
  XNOR2_X1 U38829 ( .A(n36981), .B(n33107), .ZN(n33108) );
  XNOR2_X1 U38830 ( .A(n33109), .B(n33108), .ZN(n33110) );
  XNOR2_X1 U38831 ( .A(n37079), .B(n33110), .ZN(n33112) );
  XNOR2_X1 U38832 ( .A(n34491), .B(n33893), .ZN(n33117) );
  XNOR2_X1 U38833 ( .A(n33578), .B(n33117), .ZN(n34724) );
  XNOR2_X1 U38834 ( .A(n36940), .B(n36681), .ZN(n33118) );
  XNOR2_X1 U38835 ( .A(n34238), .B(n33118), .ZN(n33129) );
  INV_X1 U38836 ( .A(n33119), .ZN(n33125) );
  XNOR2_X1 U38837 ( .A(n4908), .B(n49790), .ZN(n33120) );
  XNOR2_X1 U38838 ( .A(n33121), .B(n33120), .ZN(n33122) );
  XNOR2_X1 U38839 ( .A(n33123), .B(n33122), .ZN(n33124) );
  XNOR2_X1 U38840 ( .A(n33125), .B(n33124), .ZN(n33126) );
  XNOR2_X1 U38841 ( .A(n35835), .B(n33126), .ZN(n33127) );
  XNOR2_X1 U38842 ( .A(n33127), .B(n35501), .ZN(n33128) );
  XNOR2_X1 U38843 ( .A(n35833), .B(n33131), .ZN(n33132) );
  XNOR2_X1 U38844 ( .A(n33132), .B(n51413), .ZN(n33133) );
  XNOR2_X1 U38845 ( .A(n34719), .B(n35372), .ZN(n33134) );
  OAI22_X1 U38846 ( .A1(n38037), .A2(n38031), .B1(n36383), .B2(n35156), .ZN(
        n33150) );
  XNOR2_X1 U38847 ( .A(n34503), .B(n42240), .ZN(n33253) );
  INV_X1 U38848 ( .A(n42824), .ZN(n33138) );
  XNOR2_X1 U38849 ( .A(n33136), .B(n43202), .ZN(n33137) );
  XNOR2_X1 U38850 ( .A(n33138), .B(n33137), .ZN(n33139) );
  XNOR2_X1 U38851 ( .A(n34412), .B(n33139), .ZN(n33140) );
  XNOR2_X1 U38852 ( .A(n33140), .B(n33253), .ZN(n33141) );
  XNOR2_X1 U38853 ( .A(n35748), .B(n37303), .ZN(n34082) );
  XNOR2_X1 U38854 ( .A(n33141), .B(n34082), .ZN(n33144) );
  XNOR2_X1 U38855 ( .A(n33142), .B(n36829), .ZN(n34248) );
  XNOR2_X1 U38856 ( .A(n36746), .B(n34248), .ZN(n33143) );
  XNOR2_X1 U38857 ( .A(n33144), .B(n33143), .ZN(n33147) );
  INV_X1 U38858 ( .A(n34169), .ZN(n35106) );
  XNOR2_X1 U38860 ( .A(n37017), .B(n33729), .ZN(n33146) );
  XNOR2_X1 U38861 ( .A(n33147), .B(n33146), .ZN(n33149) );
  XNOR2_X1 U38862 ( .A(n33149), .B(n33148), .ZN(n33173) );
  AOI21_X1 U38863 ( .B1(n36383), .B2(n38043), .A(n38029), .ZN(n36370) );
  XNOR2_X1 U38864 ( .A(n35136), .B(n34305), .ZN(n33171) );
  AND2_X1 U38865 ( .A1(n51639), .A2(n33152), .ZN(n33163) );
  INV_X1 U38868 ( .A(n33157), .ZN(n33158) );
  NAND2_X1 U38869 ( .A1(n33159), .A2(n33158), .ZN(n33160) );
  XNOR2_X1 U38870 ( .A(n33164), .B(n1326), .ZN(n33165) );
  XNOR2_X1 U38871 ( .A(n33166), .B(n33165), .ZN(n33167) );
  XNOR2_X1 U38872 ( .A(n36998), .B(n33167), .ZN(n33168) );
  XNOR2_X1 U38873 ( .A(n34359), .B(n33168), .ZN(n33169) );
  XNOR2_X1 U38874 ( .A(n52220), .B(n33169), .ZN(n33170) );
  NAND2_X1 U38875 ( .A1(n35154), .A2(n34945), .ZN(n33172) );
  NAND2_X1 U38876 ( .A1(n36370), .A2(n33172), .ZN(n33177) );
  NAND2_X1 U38877 ( .A1(n34945), .A2(n38040), .ZN(n34208) );
  INV_X1 U38878 ( .A(n33173), .ZN(n38034) );
  AOI22_X1 U38879 ( .A1(n38036), .A2(n36376), .B1(n36381), .B2(n36372), .ZN(
        n33176) );
  INV_X1 U38880 ( .A(n38029), .ZN(n35157) );
  NAND3_X1 U38881 ( .A1(n38612), .A2(n682), .A3(n51012), .ZN(n38618) );
  NAND3_X1 U38883 ( .A1(n40382), .A2(n40385), .A3(n51012), .ZN(n33178) );
  XNOR2_X1 U38884 ( .A(n376), .B(n33893), .ZN(n33179) );
  XNOR2_X1 U38886 ( .A(n36858), .B(n33179), .ZN(n33186) );
  INV_X1 U38887 ( .A(n33180), .ZN(n33183) );
  XNOR2_X1 U38888 ( .A(n42327), .B(n33181), .ZN(n33182) );
  XNOR2_X1 U38889 ( .A(n33183), .B(n33182), .ZN(n33184) );
  XNOR2_X1 U38890 ( .A(n37261), .B(n33184), .ZN(n33185) );
  XNOR2_X1 U38891 ( .A(n33889), .B(n35255), .ZN(n34000) );
  XNOR2_X1 U38892 ( .A(n33187), .B(n36869), .ZN(n33189) );
  XNOR2_X1 U38893 ( .A(n33189), .B(n33188), .ZN(n35032) );
  XNOR2_X1 U38894 ( .A(n36669), .B(n34553), .ZN(n33190) );
  XNOR2_X1 U38895 ( .A(n33191), .B(n34555), .ZN(n35775) );
  XNOR2_X1 U38896 ( .A(n52117), .B(n33192), .ZN(n33193) );
  XNOR2_X1 U38897 ( .A(n33194), .B(n33193), .ZN(n33910) );
  XNOR2_X1 U38898 ( .A(n33195), .B(n34381), .ZN(n33196) );
  XNOR2_X1 U38899 ( .A(n33196), .B(n33759), .ZN(n33198) );
  INV_X1 U38900 ( .A(n34020), .ZN(n33197) );
  XNOR2_X1 U38901 ( .A(n33197), .B(n33198), .ZN(n36845) );
  XNOR2_X1 U38902 ( .A(n33200), .B(n33199), .ZN(n33203) );
  INV_X1 U38903 ( .A(n33201), .ZN(n33202) );
  XNOR2_X1 U38904 ( .A(n33203), .B(n33202), .ZN(n33204) );
  XNOR2_X1 U38905 ( .A(n34835), .B(n33204), .ZN(n33205) );
  XNOR2_X1 U38906 ( .A(n33205), .B(n37067), .ZN(n33207) );
  XNOR2_X1 U38907 ( .A(n33470), .B(n33473), .ZN(n33206) );
  XNOR2_X1 U38908 ( .A(n33207), .B(n33206), .ZN(n33208) );
  XNOR2_X1 U38909 ( .A(n36845), .B(n33208), .ZN(n33209) );
  NAND2_X1 U38910 ( .A1(n34187), .A2(n34189), .ZN(n38092) );
  XNOR2_X1 U38911 ( .A(n35237), .B(n34760), .ZN(n33210) );
  XNOR2_X1 U38912 ( .A(n33212), .B(n33211), .ZN(n35808) );
  INV_X1 U38913 ( .A(n33213), .ZN(n33214) );
  XNOR2_X1 U38914 ( .A(n33214), .B(n35808), .ZN(n33225) );
  XNOR2_X1 U38915 ( .A(n33216), .B(n33215), .ZN(n33217) );
  XNOR2_X1 U38916 ( .A(n33219), .B(n33218), .ZN(n33220) );
  XNOR2_X1 U38917 ( .A(n51495), .B(n33220), .ZN(n33223) );
  XNOR2_X1 U38918 ( .A(n36722), .B(n33221), .ZN(n35238) );
  XNOR2_X1 U38919 ( .A(n2168), .B(n35238), .ZN(n33222) );
  XNOR2_X1 U38920 ( .A(n33223), .B(n33222), .ZN(n33224) );
  INV_X1 U38921 ( .A(n33226), .ZN(n33227) );
  XNOR2_X1 U38922 ( .A(n34433), .B(n33227), .ZN(n33234) );
  XNOR2_X1 U38923 ( .A(n33228), .B(n4800), .ZN(n33229) );
  XNOR2_X1 U38924 ( .A(n33230), .B(n33229), .ZN(n33231) );
  XNOR2_X1 U38925 ( .A(n35543), .B(n33231), .ZN(n33232) );
  XNOR2_X1 U38926 ( .A(n33232), .B(n34842), .ZN(n33233) );
  XNOR2_X1 U38927 ( .A(n33234), .B(n33233), .ZN(n33236) );
  INV_X1 U38928 ( .A(n33235), .ZN(n34848) );
  XNOR2_X1 U38929 ( .A(n34848), .B(n33236), .ZN(n33239) );
  XNOR2_X1 U38930 ( .A(n34446), .B(n36704), .ZN(n34110) );
  INV_X1 U38931 ( .A(n34572), .ZN(n33237) );
  XNOR2_X1 U38932 ( .A(n33237), .B(n33398), .ZN(n34357) );
  XNOR2_X1 U38933 ( .A(n34357), .B(n34110), .ZN(n33238) );
  NAND2_X1 U38934 ( .A1(n36632), .A2(n34958), .ZN(n38086) );
  OAI22_X1 U38935 ( .A1(n36640), .A2(n38086), .B1(n34184), .B2(n1360), .ZN(
        n33270) );
  INV_X1 U38936 ( .A(n35136), .ZN(n33240) );
  XNOR2_X1 U38937 ( .A(n34294), .B(n33943), .ZN(n33450) );
  XNOR2_X1 U38938 ( .A(n33450), .B(n35128), .ZN(n33250) );
  INV_X1 U38939 ( .A(n35133), .ZN(n33241) );
  XNOR2_X1 U38940 ( .A(n33241), .B(n52219), .ZN(n33311) );
  XNOR2_X1 U38941 ( .A(n43054), .B(n4578), .ZN(n33243) );
  XNOR2_X1 U38942 ( .A(n33243), .B(n33242), .ZN(n33244) );
  XNOR2_X1 U38943 ( .A(n33245), .B(n33244), .ZN(n33246) );
  XNOR2_X1 U38944 ( .A(n34896), .B(n33246), .ZN(n33247) );
  XNOR2_X1 U38945 ( .A(n36992), .B(n33247), .ZN(n33248) );
  XNOR2_X1 U38946 ( .A(n33311), .B(n33248), .ZN(n33249) );
  XNOR2_X1 U38947 ( .A(n33250), .B(n33249), .ZN(n33251) );
  XNOR2_X1 U38948 ( .A(n35386), .B(n33253), .ZN(n33261) );
  INV_X1 U38949 ( .A(n33254), .ZN(n33257) );
  XNOR2_X1 U38950 ( .A(n34080), .B(n4739), .ZN(n33255) );
  XNOR2_X1 U38951 ( .A(n41497), .B(n33255), .ZN(n33256) );
  XNOR2_X1 U38952 ( .A(n33257), .B(n33256), .ZN(n33258) );
  XNOR2_X1 U38953 ( .A(n36747), .B(n33258), .ZN(n33259) );
  XNOR2_X1 U38954 ( .A(n33259), .B(n33145), .ZN(n33260) );
  XNOR2_X1 U38955 ( .A(n33261), .B(n33260), .ZN(n33265) );
  XNOR2_X1 U38956 ( .A(n33263), .B(n33262), .ZN(n33264) );
  XNOR2_X1 U38957 ( .A(n33265), .B(n33264), .ZN(n33269) );
  XNOR2_X1 U38958 ( .A(n34412), .B(n37303), .ZN(n33266) );
  XNOR2_X1 U38959 ( .A(n34608), .B(n33266), .ZN(n34175) );
  XNOR2_X1 U38960 ( .A(n34175), .B(n33267), .ZN(n33926) );
  XNOR2_X1 U38961 ( .A(n33926), .B(n35756), .ZN(n33268) );
  AND2_X1 U38962 ( .A1(n36628), .A2(n50984), .ZN(n36317) );
  NAND2_X1 U38963 ( .A1(n36312), .A2(n50984), .ZN(n34960) );
  AND2_X1 U38964 ( .A1(n34193), .A2(n36312), .ZN(n34199) );
  OAI211_X1 U38965 ( .C1(n36313), .C2(n695), .A(n36629), .B(n38094), .ZN(
        n33272) );
  INV_X1 U38966 ( .A(n33272), .ZN(n33273) );
  OAI21_X1 U38967 ( .B1(n34186), .B2(n34199), .A(n33273), .ZN(n33276) );
  NOR2_X1 U38969 ( .A1(n36320), .A2(n33274), .ZN(n38076) );
  INV_X1 U38971 ( .A(n36627), .ZN(n38082) );
  NAND2_X1 U38972 ( .A1(n38082), .A2(n36313), .ZN(n34190) );
  OAI21_X1 U38973 ( .B1(n38076), .B2(n36642), .A(n34190), .ZN(n33275) );
  NAND2_X1 U38974 ( .A1(n51012), .A2(n40377), .ZN(n38621) );
  NAND2_X1 U38975 ( .A1(n39843), .A2(n38621), .ZN(n33280) );
  INV_X1 U38976 ( .A(n39830), .ZN(n41152) );
  OAI21_X1 U38977 ( .B1(n39839), .B2(n1931), .A(n40385), .ZN(n33279) );
  AND2_X1 U38978 ( .A1(n39835), .A2(n39834), .ZN(n33278) );
  AOI22_X1 U38979 ( .A1(n33280), .A2(n41152), .B1(n33279), .B2(n33278), .ZN(
        n33284) );
  NOR2_X1 U38981 ( .A1(n41150), .A2(n40388), .ZN(n38622) );
  AND2_X1 U38982 ( .A1(n40377), .A2(n41150), .ZN(n37838) );
  NAND2_X1 U38983 ( .A1(n37838), .A2(n41143), .ZN(n33281) );
  AND2_X1 U38984 ( .A1(n37833), .A2(n33281), .ZN(n33283) );
  XNOR2_X1 U38985 ( .A(n34471), .B(n36931), .ZN(n34567) );
  XNOR2_X1 U38986 ( .A(n33285), .B(n4803), .ZN(n33286) );
  XNOR2_X1 U38987 ( .A(n33287), .B(n33286), .ZN(n33288) );
  XNOR2_X1 U38988 ( .A(n37062), .B(n33288), .ZN(n33289) );
  XNOR2_X1 U38989 ( .A(n33759), .B(n33289), .ZN(n33291) );
  XNOR2_X1 U38990 ( .A(n35606), .B(n33911), .ZN(n33290) );
  XNOR2_X1 U38991 ( .A(n33291), .B(n33290), .ZN(n33292) );
  XNOR2_X1 U38992 ( .A(n34567), .B(n33292), .ZN(n33293) );
  XNOR2_X1 U38993 ( .A(n34143), .B(n34555), .ZN(n35045) );
  XNOR2_X1 U38994 ( .A(n35045), .B(n34839), .ZN(n33294) );
  XNOR2_X1 U38995 ( .A(n33295), .B(n4157), .ZN(n41499) );
  XNOR2_X1 U38996 ( .A(n41499), .B(n33296), .ZN(n33298) );
  XNOR2_X1 U38997 ( .A(n33297), .B(n33429), .ZN(n44555) );
  XNOR2_X1 U38998 ( .A(n33298), .B(n44555), .ZN(n33300) );
  XNOR2_X1 U38999 ( .A(n33300), .B(n33299), .ZN(n33301) );
  XNOR2_X1 U39000 ( .A(n34169), .B(n33301), .ZN(n33302) );
  XNOR2_X1 U39001 ( .A(n34078), .B(n33302), .ZN(n33304) );
  XNOR2_X1 U39002 ( .A(n33303), .B(n35383), .ZN(n33537) );
  XNOR2_X1 U39003 ( .A(n34881), .B(n35289), .ZN(n33307) );
  XNOR2_X1 U39004 ( .A(n2131), .B(n33307), .ZN(n34782) );
  XNOR2_X1 U39005 ( .A(n35748), .B(n37304), .ZN(n36819) );
  XNOR2_X1 U39006 ( .A(n34782), .B(n36819), .ZN(n33308) );
  XNOR2_X1 U39007 ( .A(n50983), .B(n517), .ZN(n35476) );
  XNOR2_X1 U39008 ( .A(n35476), .B(n33308), .ZN(n33309) );
  XNOR2_X2 U39009 ( .A(n33310), .B(n33309), .ZN(n37496) );
  INV_X1 U39010 ( .A(n4415), .ZN(n47244) );
  XNOR2_X1 U39011 ( .A(n33311), .B(n33312), .ZN(n33323) );
  XNOR2_X1 U39012 ( .A(n33549), .B(n34156), .ZN(n33313) );
  XNOR2_X1 U39013 ( .A(n33314), .B(n33313), .ZN(n33321) );
  INV_X1 U39014 ( .A(n33315), .ZN(n33317) );
  XNOR2_X1 U39015 ( .A(n33317), .B(n33316), .ZN(n33318) );
  XNOR2_X1 U39016 ( .A(n35683), .B(n33318), .ZN(n33319) );
  XNOR2_X1 U39017 ( .A(n33319), .B(n36991), .ZN(n33320) );
  XNOR2_X1 U39018 ( .A(n33321), .B(n33320), .ZN(n33322) );
  XNOR2_X1 U39019 ( .A(n33323), .B(n33322), .ZN(n33324) );
  XNOR2_X1 U39020 ( .A(n34812), .B(n33566), .ZN(n34133) );
  XNOR2_X1 U39021 ( .A(n34133), .B(n35830), .ZN(n33325) );
  INV_X1 U39022 ( .A(n34492), .ZN(n34823) );
  XNOR2_X1 U39024 ( .A(n33326), .B(n36855), .ZN(n33333) );
  XNOR2_X1 U39025 ( .A(n34711), .B(n42460), .ZN(n33328) );
  XNOR2_X1 U39026 ( .A(n33567), .B(n4529), .ZN(n33327) );
  XNOR2_X1 U39027 ( .A(n33328), .B(n33327), .ZN(n33329) );
  XNOR2_X1 U39028 ( .A(n33330), .B(n33329), .ZN(n33331) );
  XNOR2_X1 U39029 ( .A(n35588), .B(n33331), .ZN(n33332) );
  XNOR2_X1 U39030 ( .A(n33333), .B(n33332), .ZN(n33334) );
  XNOR2_X1 U39032 ( .A(n33335), .B(n619), .ZN(n33338) );
  XNOR2_X1 U39033 ( .A(n33338), .B(n33337), .ZN(n36956) );
  INV_X1 U39034 ( .A(n36956), .ZN(n33339) );
  XNOR2_X1 U39035 ( .A(n33340), .B(n33339), .ZN(n33342) );
  XNOR2_X1 U39036 ( .A(n34720), .B(n37040), .ZN(n36868) );
  XNOR2_X1 U39037 ( .A(n36868), .B(n34128), .ZN(n34552) );
  INV_X1 U39038 ( .A(n34552), .ZN(n33341) );
  XNOR2_X1 U39041 ( .A(n33343), .B(n4909), .ZN(n33344) );
  INV_X1 U39042 ( .A(n44909), .ZN(n33349) );
  XNOR2_X1 U39043 ( .A(n43293), .B(n2183), .ZN(n33345) );
  XNOR2_X1 U39044 ( .A(n33387), .B(n33345), .ZN(n33347) );
  XNOR2_X1 U39045 ( .A(n33347), .B(n33346), .ZN(n33348) );
  XNOR2_X1 U39046 ( .A(n33349), .B(n33348), .ZN(n33350) );
  XNOR2_X1 U39047 ( .A(n37086), .B(n33350), .ZN(n33351) );
  XNOR2_X1 U39048 ( .A(n35544), .B(n33351), .ZN(n33353) );
  XNOR2_X1 U39049 ( .A(n33353), .B(n33352), .ZN(n33354) );
  XNOR2_X1 U39050 ( .A(n36703), .B(n35095), .ZN(n33864) );
  XNOR2_X1 U39051 ( .A(n51449), .B(n35086), .ZN(n34858) );
  INV_X1 U39052 ( .A(n37091), .ZN(n33355) );
  XNOR2_X1 U39053 ( .A(n33355), .B(n34858), .ZN(n33356) );
  XNOR2_X1 U39054 ( .A(n36812), .B(n35334), .ZN(n33357) );
  XNOR2_X1 U39055 ( .A(n33357), .B(n37108), .ZN(n33358) );
  XNOR2_X1 U39056 ( .A(n37097), .B(n33358), .ZN(n35561) );
  XNOR2_X1 U39057 ( .A(n33359), .B(n35561), .ZN(n33369) );
  INV_X1 U39058 ( .A(n34760), .ZN(n33360) );
  XNOR2_X1 U39059 ( .A(n33362), .B(n33361), .ZN(n33363) );
  XNOR2_X1 U39060 ( .A(n35075), .B(n33363), .ZN(n33364) );
  XNOR2_X1 U39061 ( .A(n33702), .B(n33711), .ZN(n33365) );
  XNOR2_X1 U39062 ( .A(n33365), .B(n36811), .ZN(n33366) );
  XNOR2_X1 U39063 ( .A(n33382), .B(n33366), .ZN(n37100) );
  XNOR2_X1 U39064 ( .A(n33367), .B(n37100), .ZN(n33368) );
  NAND2_X1 U39066 ( .A1(n37750), .A2(n37496), .ZN(n36242) );
  NAND2_X1 U39067 ( .A1(n37750), .A2(n37759), .ZN(n37502) );
  NAND2_X1 U39068 ( .A1(n37496), .A2(n36251), .ZN(n36244) );
  XNOR2_X1 U39069 ( .A(n51445), .B(n34869), .ZN(n33371) );
  XNOR2_X1 U39070 ( .A(n35325), .B(n33372), .ZN(n33379) );
  INV_X1 U39071 ( .A(n33373), .ZN(n33376) );
  XNOR2_X1 U39072 ( .A(n33374), .B(n1354), .ZN(n33375) );
  XNOR2_X1 U39073 ( .A(n33376), .B(n33375), .ZN(n33377) );
  XNOR2_X1 U39074 ( .A(n33973), .B(n33377), .ZN(n33378) );
  XNOR2_X1 U39075 ( .A(n33379), .B(n33378), .ZN(n33380) );
  XNOR2_X1 U39076 ( .A(n33711), .B(n36811), .ZN(n33605) );
  XNOR2_X1 U39077 ( .A(n52197), .B(n36960), .ZN(n33384) );
  XNOR2_X1 U39078 ( .A(n515), .B(n35635), .ZN(n36988) );
  XNOR2_X1 U39079 ( .A(n33387), .B(n4647), .ZN(n33389) );
  XNOR2_X1 U39080 ( .A(n33389), .B(n33388), .ZN(n33390) );
  XNOR2_X1 U39081 ( .A(n33391), .B(n33390), .ZN(n33392) );
  XNOR2_X1 U39082 ( .A(n35537), .B(n33392), .ZN(n33393) );
  INV_X1 U39083 ( .A(n36703), .ZN(n34351) );
  XNOR2_X1 U39084 ( .A(n33393), .B(n34351), .ZN(n33394) );
  XNOR2_X1 U39085 ( .A(n36988), .B(n33394), .ZN(n33396) );
  XNOR2_X1 U39086 ( .A(n33396), .B(n33718), .ZN(n33401) );
  XNOR2_X1 U39087 ( .A(n52119), .B(n35534), .ZN(n33399) );
  XNOR2_X1 U39088 ( .A(n36796), .B(n33399), .ZN(n33400) );
  XNOR2_X1 U39089 ( .A(n33401), .B(n33400), .ZN(n36196) );
  INV_X1 U39090 ( .A(n36196), .ZN(n33456) );
  XNOR2_X1 U39091 ( .A(n34141), .B(n37241), .ZN(n33402) );
  XNOR2_X1 U39092 ( .A(n33402), .B(n52148), .ZN(n33403) );
  XNOR2_X1 U39093 ( .A(n33403), .B(n51472), .ZN(n36935) );
  INV_X1 U39094 ( .A(n33404), .ZN(n33405) );
  XNOR2_X1 U39095 ( .A(n34835), .B(n33405), .ZN(n33831) );
  XNOR2_X1 U39096 ( .A(n33406), .B(n49109), .ZN(n33408) );
  XNOR2_X1 U39097 ( .A(n33408), .B(n33407), .ZN(n33409) );
  XNOR2_X1 U39098 ( .A(n33753), .B(n33409), .ZN(n33410) );
  XNOR2_X1 U39099 ( .A(n33831), .B(n33410), .ZN(n33411) );
  XNOR2_X1 U39100 ( .A(n34471), .B(n34739), .ZN(n33413) );
  XNOR2_X1 U39101 ( .A(n33470), .B(n34219), .ZN(n33412) );
  XNOR2_X1 U39102 ( .A(n33413), .B(n33412), .ZN(n34389) );
  INV_X1 U39103 ( .A(n34389), .ZN(n33414) );
  INV_X1 U39105 ( .A(n39350), .ZN(n34692) );
  INV_X1 U39106 ( .A(n34238), .ZN(n33416) );
  XNOR2_X1 U39107 ( .A(n36856), .B(n33416), .ZN(n34394) );
  XNOR2_X1 U39108 ( .A(n376), .B(n36939), .ZN(n33417) );
  XNOR2_X1 U39109 ( .A(n33417), .B(n35830), .ZN(n33765) );
  XNOR2_X1 U39110 ( .A(n34394), .B(n33765), .ZN(n33418) );
  INV_X1 U39111 ( .A(n33420), .ZN(n33421) );
  XNOR2_X1 U39112 ( .A(n33421), .B(n4897), .ZN(n42757) );
  XNOR2_X1 U39113 ( .A(n42757), .B(n33422), .ZN(n33423) );
  XNOR2_X1 U39114 ( .A(n37045), .B(n33423), .ZN(n33424) );
  XNOR2_X1 U39115 ( .A(n33902), .B(n33424), .ZN(n33425) );
  XNOR2_X1 U39116 ( .A(n33425), .B(n51702), .ZN(n33426) );
  INV_X1 U39117 ( .A(n33427), .ZN(n33454) );
  XNOR2_X1 U39118 ( .A(n37019), .B(n33740), .ZN(n33428) );
  XNOR2_X1 U39119 ( .A(n33430), .B(n33429), .ZN(n33431) );
  XNOR2_X1 U39120 ( .A(n33432), .B(n33431), .ZN(n33433) );
  XNOR2_X1 U39121 ( .A(n33434), .B(n35464), .ZN(n33435) );
  XNOR2_X1 U39122 ( .A(n37324), .B(n34156), .ZN(n33437) );
  XNOR2_X1 U39123 ( .A(n35133), .B(n33437), .ZN(n33438) );
  XNOR2_X1 U39124 ( .A(n33540), .B(n33438), .ZN(n33441) );
  XNOR2_X1 U39125 ( .A(n36999), .B(n34361), .ZN(n33664) );
  XNOR2_X1 U39126 ( .A(n33439), .B(n33664), .ZN(n33440) );
  XNOR2_X1 U39127 ( .A(n33441), .B(n33440), .ZN(n33683) );
  INV_X1 U39128 ( .A(n35761), .ZN(n37319) );
  XNOR2_X1 U39129 ( .A(n33549), .B(n37319), .ZN(n33448) );
  XNOR2_X1 U39130 ( .A(n33443), .B(n33442), .ZN(n33444) );
  XNOR2_X1 U39131 ( .A(n33445), .B(n33444), .ZN(n33446) );
  XNOR2_X1 U39132 ( .A(n33806), .B(n33446), .ZN(n33447) );
  XNOR2_X1 U39133 ( .A(n33448), .B(n33447), .ZN(n33449) );
  XNOR2_X1 U39134 ( .A(n33450), .B(n33449), .ZN(n33452) );
  XNOR2_X1 U39135 ( .A(n701), .B(n35283), .ZN(n34372) );
  INV_X1 U39136 ( .A(n34372), .ZN(n33451) );
  AND2_X1 U39137 ( .A1(n37774), .A2(n36200), .ZN(n39348) );
  OAI211_X1 U39138 ( .C1(n33454), .C2(n39349), .A(n33453), .B(n39348), .ZN(
        n33455) );
  NAND2_X1 U39139 ( .A1(n36186), .A2(n36189), .ZN(n33458) );
  INV_X1 U39140 ( .A(n39342), .ZN(n36191) );
  AOI21_X1 U39142 ( .B1(n39347), .B2(n36199), .A(n37778), .ZN(n33460) );
  NAND2_X1 U39143 ( .A1(n37775), .A2(n36196), .ZN(n35943) );
  INV_X1 U39144 ( .A(n37780), .ZN(n33457) );
  OAI21_X1 U39145 ( .B1(n35943), .B2(n52054), .A(n33457), .ZN(n34684) );
  NAND3_X1 U39146 ( .A1(n34684), .A2(n37782), .A3(n33458), .ZN(n33459) );
  OAI211_X1 U39147 ( .C1(n36199), .C2(n36196), .A(n37775), .B(n39340), .ZN(
        n36202) );
  NAND2_X1 U39148 ( .A1(n39347), .A2(n33461), .ZN(n34691) );
  INV_X1 U39149 ( .A(n37781), .ZN(n33462) );
  NAND3_X1 U39150 ( .A1(n33464), .A2(n39340), .A3(n39351), .ZN(n33465) );
  XNOR2_X1 U39151 ( .A(n34829), .B(n34555), .ZN(n36844) );
  INV_X1 U39152 ( .A(n33467), .ZN(n33468) );
  XNOR2_X1 U39153 ( .A(n35522), .B(n33468), .ZN(n33469) );
  XNOR2_X1 U39154 ( .A(n33469), .B(n34219), .ZN(n33471) );
  XNOR2_X1 U39155 ( .A(n51463), .B(n33471), .ZN(n33472) );
  XNOR2_X1 U39156 ( .A(n34466), .B(n37066), .ZN(n35049) );
  XNOR2_X1 U39157 ( .A(n35049), .B(n33473), .ZN(n33483) );
  XOR2_X1 U39158 ( .A(n4486), .B(n4823), .Z(n33475) );
  XNOR2_X1 U39159 ( .A(n33475), .B(n33474), .ZN(n33476) );
  XNOR2_X1 U39160 ( .A(n34377), .B(n33476), .ZN(n33479) );
  INV_X1 U39161 ( .A(n33477), .ZN(n33478) );
  XNOR2_X1 U39162 ( .A(n33479), .B(n33478), .ZN(n33480) );
  XNOR2_X1 U39163 ( .A(n34381), .B(n33480), .ZN(n33481) );
  XNOR2_X1 U39164 ( .A(n33481), .B(n34141), .ZN(n33482) );
  XNOR2_X1 U39165 ( .A(n33483), .B(n33482), .ZN(n33486) );
  INV_X1 U39166 ( .A(n33751), .ZN(n33484) );
  XNOR2_X1 U39167 ( .A(n33486), .B(n33485), .ZN(n33487) );
  INV_X1 U39168 ( .A(n33489), .ZN(n33892) );
  INV_X1 U39169 ( .A(n33490), .ZN(n33491) );
  XNOR2_X1 U39170 ( .A(n37262), .B(n33491), .ZN(n35250) );
  INV_X1 U39171 ( .A(n35250), .ZN(n33492) );
  XNOR2_X1 U39172 ( .A(n34720), .B(n33492), .ZN(n33493) );
  XNOR2_X1 U39173 ( .A(n33892), .B(n33493), .ZN(n33505) );
  XNOR2_X1 U39174 ( .A(n4529), .B(n45736), .ZN(n33494) );
  XNOR2_X1 U39175 ( .A(n33495), .B(n33494), .ZN(n33496) );
  XNOR2_X1 U39176 ( .A(n35036), .B(n33496), .ZN(n33497) );
  XNOR2_X1 U39177 ( .A(n35503), .B(n33497), .ZN(n33498) );
  XNOR2_X1 U39178 ( .A(n704), .B(n33498), .ZN(n33499) );
  XNOR2_X1 U39179 ( .A(n33764), .B(n33499), .ZN(n33504) );
  XNOR2_X1 U39180 ( .A(n34546), .B(n376), .ZN(n33501) );
  XNOR2_X1 U39181 ( .A(n35829), .B(n2230), .ZN(n33500) );
  XNOR2_X1 U39182 ( .A(n33501), .B(n33500), .ZN(n33503) );
  XNOR2_X1 U39183 ( .A(n33503), .B(n33502), .ZN(n34405) );
  XNOR2_X1 U39185 ( .A(n37096), .B(n34275), .ZN(n33507) );
  XNOR2_X1 U39186 ( .A(n37269), .B(n703), .ZN(n33506) );
  XNOR2_X1 U39187 ( .A(n33507), .B(n33506), .ZN(n35232) );
  XNOR2_X1 U39188 ( .A(n37277), .B(n35333), .ZN(n34342) );
  XNOR2_X1 U39189 ( .A(n33508), .B(n49937), .ZN(n33509) );
  XNOR2_X1 U39190 ( .A(n33510), .B(n33509), .ZN(n33511) );
  XNOR2_X1 U39191 ( .A(n37108), .B(n33511), .ZN(n33512) );
  XNOR2_X1 U39192 ( .A(n36807), .B(n33512), .ZN(n33513) );
  XNOR2_X1 U39193 ( .A(n34342), .B(n33513), .ZN(n33514) );
  XNOR2_X1 U39194 ( .A(n35232), .B(n33514), .ZN(n33518) );
  XNOR2_X1 U39195 ( .A(n34594), .B(n4837), .ZN(n33618) );
  INV_X1 U39196 ( .A(n4636), .ZN(n47802) );
  XNOR2_X1 U39197 ( .A(n33711), .B(n47802), .ZN(n35619) );
  XNOR2_X1 U39198 ( .A(n33515), .B(n35619), .ZN(n33516) );
  XNOR2_X1 U39199 ( .A(n33517), .B(n33516), .ZN(n35551) );
  XNOR2_X1 U39200 ( .A(n33722), .B(n34842), .ZN(n35096) );
  XNOR2_X1 U39201 ( .A(n34446), .B(n35096), .ZN(n33524) );
  XNOR2_X1 U39202 ( .A(n33520), .B(n33519), .ZN(n33521) );
  XNOR2_X1 U39203 ( .A(n35224), .B(n33521), .ZN(n33522) );
  XNOR2_X1 U39204 ( .A(n35534), .B(n33522), .ZN(n33523) );
  XNOR2_X1 U39205 ( .A(n33524), .B(n33523), .ZN(n33525) );
  XNOR2_X1 U39206 ( .A(n33525), .B(n36714), .ZN(n33528) );
  INV_X1 U39207 ( .A(n34350), .ZN(n35649) );
  XNOR2_X1 U39208 ( .A(n36988), .B(n35649), .ZN(n33527) );
  XNOR2_X1 U39209 ( .A(n33528), .B(n33527), .ZN(n37519) );
  XNOR2_X1 U39210 ( .A(Key[189]), .B(n4587), .ZN(n43647) );
  XNOR2_X1 U39211 ( .A(n33529), .B(n43647), .ZN(n33530) );
  XNOR2_X1 U39212 ( .A(n33530), .B(n43150), .ZN(n33531) );
  XNOR2_X1 U39213 ( .A(n33531), .B(n45105), .ZN(n33532) );
  XNOR2_X1 U39214 ( .A(n45310), .B(n33532), .ZN(n33533) );
  XNOR2_X1 U39215 ( .A(n36818), .B(n33533), .ZN(n33534) );
  XNOR2_X1 U39216 ( .A(n33534), .B(n37023), .ZN(n33536) );
  XNOR2_X1 U39217 ( .A(n518), .B(n34883), .ZN(n33535) );
  XNOR2_X1 U39218 ( .A(n33536), .B(n33535), .ZN(n33538) );
  INV_X1 U39219 ( .A(n33539), .ZN(n33946) );
  XNOR2_X1 U39220 ( .A(n33543), .B(n4847), .ZN(n33544) );
  XNOR2_X1 U39221 ( .A(n33545), .B(n33544), .ZN(n33546) );
  XNOR2_X1 U39222 ( .A(n35762), .B(n33546), .ZN(n33547) );
  XNOR2_X1 U39223 ( .A(n33547), .B(n51366), .ZN(n33548) );
  XNOR2_X1 U39224 ( .A(n51422), .B(n33548), .ZN(n33553) );
  XNOR2_X1 U39225 ( .A(n34360), .B(n35483), .ZN(n33551) );
  XNOR2_X1 U39226 ( .A(n37001), .B(n33551), .ZN(n33552) );
  XNOR2_X1 U39227 ( .A(n33553), .B(n33552), .ZN(n33554) );
  XNOR2_X2 U39228 ( .A(n33555), .B(n33554), .ZN(n38494) );
  NOR3_X1 U39229 ( .A1(n37387), .A2(n618), .A3(n37384), .ZN(n33556) );
  NAND3_X1 U39230 ( .A1(n37520), .A2(n38496), .A3(n33556), .ZN(n33557) );
  NAND3_X1 U39231 ( .A1(n35953), .A2(n38495), .A3(n37384), .ZN(n37518) );
  AND2_X1 U39232 ( .A1(n37521), .A2(n37520), .ZN(n35577) );
  NAND3_X1 U39233 ( .A1(n38495), .A2(n38494), .A3(n38496), .ZN(n37531) );
  INV_X1 U39234 ( .A(n37531), .ZN(n33561) );
  NAND2_X1 U39235 ( .A1(n37385), .A2(n618), .ZN(n35949) );
  AOI21_X1 U39236 ( .B1(n37531), .B2(n35950), .A(n35949), .ZN(n33560) );
  OAI21_X1 U39237 ( .B1(n35577), .B2(n33561), .A(n33560), .ZN(n33564) );
  NOR2_X1 U39238 ( .A1(n35951), .A2(n38496), .ZN(n37394) );
  OAI21_X1 U39240 ( .B1(n37394), .B2(n35571), .A(n35578), .ZN(n33563) );
  INV_X1 U39241 ( .A(n41403), .ZN(n33570) );
  XNOR2_X1 U39242 ( .A(n33568), .B(n33567), .ZN(n33569) );
  XNOR2_X1 U39243 ( .A(n33570), .B(n33569), .ZN(n33571) );
  XNOR2_X1 U39244 ( .A(n34546), .B(n33571), .ZN(n33572) );
  XNOR2_X1 U39245 ( .A(n376), .B(n36855), .ZN(n33573) );
  XNOR2_X1 U39246 ( .A(n34240), .B(n33573), .ZN(n33574) );
  XNOR2_X1 U39247 ( .A(n33575), .B(n33574), .ZN(n33577) );
  XNOR2_X1 U39248 ( .A(n35830), .B(n34400), .ZN(n34132) );
  XNOR2_X1 U39249 ( .A(n34535), .B(n34132), .ZN(n33576) );
  XNOR2_X1 U39250 ( .A(n33577), .B(n33576), .ZN(n33582) );
  XNOR2_X1 U39251 ( .A(n33578), .B(n51702), .ZN(n33581) );
  XNOR2_X1 U39252 ( .A(n35503), .B(n619), .ZN(n33579) );
  XNOR2_X1 U39253 ( .A(n704), .B(n33579), .ZN(n33580) );
  INV_X1 U39254 ( .A(n33583), .ZN(n33584) );
  XNOR2_X1 U39256 ( .A(n34382), .B(n49109), .ZN(n34221) );
  XNOR2_X1 U39257 ( .A(n34143), .B(n34221), .ZN(n33587) );
  XNOR2_X1 U39258 ( .A(n34381), .B(n37241), .ZN(n33586) );
  INV_X1 U39259 ( .A(n33911), .ZN(n33585) );
  XNOR2_X1 U39260 ( .A(n33586), .B(n33585), .ZN(n35514) );
  XNOR2_X1 U39261 ( .A(n33587), .B(n35514), .ZN(n33602) );
  INV_X1 U39262 ( .A(n33588), .ZN(n33593) );
  XNOR2_X1 U39263 ( .A(n33589), .B(n5016), .ZN(n33591) );
  INV_X1 U39264 ( .A(n43985), .ZN(n33590) );
  XNOR2_X1 U39265 ( .A(n33591), .B(n33590), .ZN(n33592) );
  XNOR2_X1 U39266 ( .A(n33593), .B(n33592), .ZN(n33594) );
  XNOR2_X1 U39267 ( .A(n35606), .B(n33594), .ZN(n33596) );
  XNOR2_X1 U39268 ( .A(n36841), .B(n35609), .ZN(n33595) );
  XNOR2_X1 U39269 ( .A(n33596), .B(n33595), .ZN(n33600) );
  XNOR2_X1 U39270 ( .A(n36931), .B(n51446), .ZN(n33598) );
  XNOR2_X1 U39271 ( .A(n35522), .B(n35512), .ZN(n33597) );
  XNOR2_X1 U39272 ( .A(n33598), .B(n33597), .ZN(n33599) );
  XNOR2_X1 U39273 ( .A(n33600), .B(n33599), .ZN(n33601) );
  XNOR2_X1 U39274 ( .A(n33602), .B(n33601), .ZN(n33603) );
  OR2_X1 U39275 ( .A1(n37406), .A2(n51418), .ZN(n36268) );
  XNOR2_X1 U39276 ( .A(n36805), .B(n1354), .ZN(n33604) );
  XNOR2_X1 U39277 ( .A(n33605), .B(n33604), .ZN(n33606) );
  XNOR2_X1 U39278 ( .A(n33607), .B(n33606), .ZN(n34461) );
  INV_X1 U39279 ( .A(n36812), .ZN(n33609) );
  XNOR2_X1 U39280 ( .A(n33610), .B(n35810), .ZN(n36727) );
  XNOR2_X1 U39281 ( .A(n34461), .B(n36727), .ZN(n33620) );
  XNOR2_X1 U39282 ( .A(n33612), .B(n33611), .ZN(n33613) );
  XNOR2_X1 U39283 ( .A(n35070), .B(n33613), .ZN(n33615) );
  XNOR2_X1 U39284 ( .A(n33702), .B(n2204), .ZN(n33614) );
  XNOR2_X1 U39285 ( .A(n33615), .B(n33614), .ZN(n33616) );
  XNOR2_X1 U39286 ( .A(n33617), .B(n33618), .ZN(n34264) );
  NAND2_X1 U39287 ( .A1(n36268), .A2(n34676), .ZN(n33676) );
  XNOR2_X1 U39288 ( .A(n37079), .B(n34754), .ZN(n33623) );
  INV_X1 U39289 ( .A(n34446), .ZN(n33621) );
  XNOR2_X1 U39290 ( .A(n33621), .B(n34433), .ZN(n33622) );
  XNOR2_X1 U39291 ( .A(n33623), .B(n33622), .ZN(n33624) );
  XNOR2_X1 U39292 ( .A(n33624), .B(n33718), .ZN(n33633) );
  XNOR2_X1 U39293 ( .A(n33625), .B(n43968), .ZN(n33626) );
  XNOR2_X1 U39294 ( .A(n33627), .B(n33626), .ZN(n33628) );
  XNOR2_X1 U39295 ( .A(n36792), .B(n33628), .ZN(n33629) );
  XNOR2_X1 U39296 ( .A(n33630), .B(n33629), .ZN(n33631) );
  XNOR2_X1 U39297 ( .A(n36988), .B(n33631), .ZN(n33632) );
  XNOR2_X1 U39298 ( .A(n33633), .B(n33632), .ZN(n33648) );
  XNOR2_X1 U39299 ( .A(n37304), .B(n33145), .ZN(n33634) );
  XNOR2_X1 U39300 ( .A(n33634), .B(n34078), .ZN(n33644) );
  XNOR2_X1 U39301 ( .A(n34169), .B(n2131), .ZN(n33642) );
  XNOR2_X1 U39302 ( .A(n33635), .B(n4045), .ZN(n33636) );
  XNOR2_X1 U39303 ( .A(n45105), .B(n33636), .ZN(n33637) );
  XNOR2_X1 U39304 ( .A(n42243), .B(n33637), .ZN(n33639) );
  XNOR2_X1 U39305 ( .A(n33639), .B(n33638), .ZN(n33640) );
  XNOR2_X1 U39306 ( .A(n35745), .B(n33640), .ZN(n33641) );
  XNOR2_X1 U39307 ( .A(n33642), .B(n33641), .ZN(n33643) );
  INV_X1 U39308 ( .A(n33645), .ZN(n33646) );
  XNOR2_X1 U39309 ( .A(n37019), .B(n33646), .ZN(n33647) );
  NOR2_X1 U39310 ( .A1(n37553), .A2(n37560), .ZN(n33672) );
  NAND2_X1 U39311 ( .A1(n37545), .A2(n37544), .ZN(n37397) );
  INV_X1 U39312 ( .A(n33651), .ZN(n33657) );
  XNOR2_X1 U39313 ( .A(n33653), .B(n33652), .ZN(n33654) );
  XNOR2_X1 U39314 ( .A(n33655), .B(n33654), .ZN(n33656) );
  XNOR2_X1 U39315 ( .A(n33657), .B(n33656), .ZN(n33658) );
  XNOR2_X1 U39316 ( .A(n34369), .B(n33658), .ZN(n33659) );
  XNOR2_X1 U39317 ( .A(n35124), .B(n33659), .ZN(n33661) );
  INV_X1 U39318 ( .A(n35477), .ZN(n33660) );
  XNOR2_X1 U39319 ( .A(n33660), .B(n33661), .ZN(n33662) );
  XNOR2_X1 U39320 ( .A(n35680), .B(n33662), .ZN(n33667) );
  XNOR2_X1 U39321 ( .A(n36991), .B(n35483), .ZN(n33663) );
  XNOR2_X1 U39322 ( .A(n35488), .B(n33663), .ZN(n34626) );
  XNOR2_X1 U39324 ( .A(n33664), .B(n37324), .ZN(n35403) );
  XNOR2_X1 U39326 ( .A(n33667), .B(n33666), .ZN(n33670) );
  INV_X1 U39327 ( .A(n33668), .ZN(n33669) );
  INV_X1 U39328 ( .A(n36272), .ZN(n37561) );
  NAND4_X1 U39329 ( .A1(n34676), .A2(n37399), .A3(n37561), .A4(n37557), .ZN(
        n33671) );
  NAND4_X1 U39330 ( .A1(n33672), .A2(n525), .A3(n37397), .A4(n33671), .ZN(
        n33673) );
  OAI211_X1 U39331 ( .C1(n36281), .C2(n33674), .A(n33673), .B(n37533), .ZN(
        n33682) );
  INV_X1 U39332 ( .A(n36268), .ZN(n37547) );
  NAND2_X1 U39333 ( .A1(n37547), .A2(n37557), .ZN(n33675) );
  NAND2_X1 U39334 ( .A1(n33676), .A2(n33675), .ZN(n33680) );
  NAND2_X1 U39335 ( .A1(n37545), .A2(n37560), .ZN(n36269) );
  OAI211_X1 U39336 ( .C1(n36272), .C2(n37560), .A(n37399), .B(n37543), .ZN(
        n33677) );
  NOR2_X1 U39337 ( .A1(n33678), .A2(n33677), .ZN(n33679) );
  NAND2_X1 U39338 ( .A1(n36272), .A2(n37560), .ZN(n34681) );
  MUX2_X1 U39339 ( .A(n33680), .B(n33679), .S(n34681), .Z(n33681) );
  NAND3_X1 U39340 ( .A1(n43667), .A2(n51950), .A3(n40632), .ZN(n33882) );
  INV_X1 U39341 ( .A(n33683), .ZN(n33695) );
  XNOR2_X1 U39342 ( .A(n36758), .B(n41223), .ZN(n33685) );
  INV_X1 U39343 ( .A(n35762), .ZN(n33684) );
  XNOR2_X1 U39344 ( .A(n33685), .B(n33684), .ZN(n33688) );
  XNOR2_X1 U39345 ( .A(n34622), .B(n36881), .ZN(n33687) );
  XNOR2_X1 U39346 ( .A(n33688), .B(n33687), .ZN(n34161) );
  XNOR2_X1 U39347 ( .A(n33690), .B(n33689), .ZN(n33691) );
  XNOR2_X1 U39348 ( .A(n33692), .B(n36991), .ZN(n33693) );
  XNOR2_X1 U39349 ( .A(n34620), .B(n37325), .ZN(n35668) );
  XNOR2_X1 U39350 ( .A(n33693), .B(n35668), .ZN(n33694) );
  INV_X1 U39351 ( .A(n33780), .ZN(n37587) );
  INV_X1 U39352 ( .A(n33696), .ZN(n33700) );
  XNOR2_X1 U39353 ( .A(n48843), .B(n46552), .ZN(n33697) );
  XNOR2_X1 U39354 ( .A(n33698), .B(n33697), .ZN(n33699) );
  XNOR2_X1 U39355 ( .A(n33700), .B(n33699), .ZN(n33701) );
  XNOR2_X1 U39356 ( .A(n33702), .B(n33701), .ZN(n33704) );
  XNOR2_X1 U39357 ( .A(n33704), .B(n35625), .ZN(n33705) );
  XNOR2_X1 U39358 ( .A(n33707), .B(n37111), .ZN(n33708) );
  XNOR2_X1 U39359 ( .A(n37113), .B(n2204), .ZN(n33710) );
  XNOR2_X1 U39360 ( .A(n37095), .B(n33710), .ZN(n33853) );
  INV_X1 U39361 ( .A(n33853), .ZN(n35326) );
  XNOR2_X1 U39362 ( .A(n33711), .B(n41660), .ZN(n33712) );
  XNOR2_X1 U39363 ( .A(n33712), .B(n36811), .ZN(n34341) );
  INV_X1 U39364 ( .A(n34341), .ZN(n33713) );
  XNOR2_X1 U39365 ( .A(n35326), .B(n33713), .ZN(n33714) );
  XNOR2_X1 U39366 ( .A(n35534), .B(n34446), .ZN(n33715) );
  XNOR2_X1 U39367 ( .A(n33715), .B(n34754), .ZN(n33717) );
  XNOR2_X1 U39368 ( .A(n36704), .B(n34753), .ZN(n33716) );
  XNOR2_X1 U39369 ( .A(n33717), .B(n33716), .ZN(n35349) );
  XNOR2_X1 U39370 ( .A(n33720), .B(n33719), .ZN(n33721) );
  XNOR2_X1 U39371 ( .A(n33722), .B(n33721), .ZN(n33723) );
  XNOR2_X1 U39372 ( .A(n33723), .B(n35633), .ZN(n33724) );
  XNOR2_X1 U39373 ( .A(n33726), .B(n33725), .ZN(n33727) );
  XNOR2_X1 U39374 ( .A(n35387), .B(n35386), .ZN(n33730) );
  XNOR2_X1 U39375 ( .A(n33730), .B(n33729), .ZN(n35662) );
  INV_X1 U39376 ( .A(n33731), .ZN(n33738) );
  INV_X1 U39377 ( .A(n33732), .ZN(n33736) );
  XNOR2_X1 U39378 ( .A(n33734), .B(n33733), .ZN(n33735) );
  XNOR2_X1 U39379 ( .A(n33736), .B(n33735), .ZN(n33737) );
  XNOR2_X1 U39380 ( .A(n33738), .B(n33737), .ZN(n33739) );
  XNOR2_X1 U39381 ( .A(n37017), .B(n33739), .ZN(n33741) );
  XNOR2_X1 U39382 ( .A(n33741), .B(n33740), .ZN(n33742) );
  XNOR2_X1 U39383 ( .A(n33742), .B(n35662), .ZN(n33743) );
  INV_X1 U39384 ( .A(n34726), .ZN(n33744) );
  XNOR2_X1 U39385 ( .A(n34567), .B(n33744), .ZN(n37071) );
  XNOR2_X1 U39386 ( .A(n33745), .B(n49109), .ZN(n33747) );
  XNOR2_X1 U39387 ( .A(n33747), .B(n33746), .ZN(n33748) );
  XNOR2_X1 U39388 ( .A(n33749), .B(n33748), .ZN(n33750) );
  XNOR2_X1 U39389 ( .A(n34141), .B(n33750), .ZN(n33752) );
  XNOR2_X1 U39390 ( .A(n33752), .B(n33751), .ZN(n33755) );
  XNOR2_X1 U39391 ( .A(n35778), .B(n33753), .ZN(n33754) );
  XNOR2_X1 U39392 ( .A(n33755), .B(n33754), .ZN(n33756) );
  XNOR2_X1 U39393 ( .A(n37071), .B(n33756), .ZN(n33762) );
  XNOR2_X1 U39394 ( .A(n37067), .B(n35609), .ZN(n33757) );
  XNOR2_X1 U39395 ( .A(n33757), .B(n34219), .ZN(n33758) );
  XNOR2_X1 U39396 ( .A(n33758), .B(n34555), .ZN(n34737) );
  INV_X1 U39397 ( .A(n34381), .ZN(n33760) );
  XNOR2_X1 U39398 ( .A(n33759), .B(n33760), .ZN(n34474) );
  INV_X1 U39399 ( .A(n34474), .ZN(n35790) );
  XNOR2_X1 U39400 ( .A(n35790), .B(n34020), .ZN(n35351) );
  INV_X1 U39401 ( .A(n35351), .ZN(n33761) );
  INV_X1 U39402 ( .A(n33763), .ZN(n33767) );
  XNOR2_X1 U39403 ( .A(n33764), .B(n33765), .ZN(n33766) );
  XNOR2_X1 U39404 ( .A(n33767), .B(n33766), .ZN(n33777) );
  INV_X1 U39405 ( .A(n33768), .ZN(n33770) );
  XNOR2_X1 U39406 ( .A(n33770), .B(n33769), .ZN(n33771) );
  XNOR2_X1 U39407 ( .A(n35589), .B(n33771), .ZN(n33772) );
  XNOR2_X1 U39408 ( .A(n33772), .B(n37252), .ZN(n33774) );
  XNOR2_X1 U39409 ( .A(n35595), .B(n619), .ZN(n33773) );
  XNOR2_X1 U39410 ( .A(n33774), .B(n33773), .ZN(n33776) );
  INV_X1 U39411 ( .A(n33778), .ZN(n37596) );
  NAND3_X1 U39412 ( .A1(n36233), .A2(n35458), .A3(n35452), .ZN(n33779) );
  NOR2_X1 U39413 ( .A1(n35457), .A2(n37593), .ZN(n33781) );
  OAI21_X1 U39414 ( .B1(n37379), .B2(n33781), .A(n37597), .ZN(n33782) );
  NAND2_X1 U39415 ( .A1(n37592), .A2(n37378), .ZN(n33783) );
  NAND2_X1 U39416 ( .A1(n33784), .A2(n33783), .ZN(n33785) );
  INV_X1 U39417 ( .A(n34514), .ZN(n33788) );
  XNOR2_X1 U39418 ( .A(n33788), .B(n35105), .ZN(n33789) );
  XNOR2_X1 U39419 ( .A(n33790), .B(n33789), .ZN(n36821) );
  XNOR2_X1 U39420 ( .A(n34425), .B(n33791), .ZN(n33799) );
  XNOR2_X1 U39421 ( .A(n41496), .B(n4940), .ZN(n33792) );
  XNOR2_X1 U39422 ( .A(n33793), .B(n33792), .ZN(n33794) );
  XNOR2_X1 U39423 ( .A(n33795), .B(n33794), .ZN(n33796) );
  XNOR2_X1 U39424 ( .A(n35468), .B(n33796), .ZN(n33797) );
  XNOR2_X1 U39425 ( .A(n35386), .B(n33797), .ZN(n33798) );
  XNOR2_X1 U39426 ( .A(n33799), .B(n33798), .ZN(n33800) );
  XNOR2_X1 U39427 ( .A(n33800), .B(n36821), .ZN(n33805) );
  INV_X1 U39428 ( .A(n35745), .ZN(n33801) );
  XNOR2_X1 U39429 ( .A(n37017), .B(n33801), .ZN(n33802) );
  XNOR2_X1 U39430 ( .A(n33803), .B(n33802), .ZN(n34786) );
  INV_X1 U39431 ( .A(n34786), .ZN(n33804) );
  XNOR2_X1 U39432 ( .A(n33804), .B(n33805), .ZN(n33871) );
  XNOR2_X1 U39433 ( .A(n34296), .B(n35124), .ZN(n37119) );
  XNOR2_X1 U39434 ( .A(n33808), .B(n49414), .ZN(n33809) );
  XNOR2_X1 U39435 ( .A(n24827), .B(n33809), .ZN(n33810) );
  XNOR2_X1 U39436 ( .A(n36999), .B(n33810), .ZN(n33811) );
  XNOR2_X1 U39437 ( .A(n33943), .B(n33811), .ZN(n33812) );
  XNOR2_X1 U39438 ( .A(n37119), .B(n33812), .ZN(n33813) );
  XNOR2_X1 U39439 ( .A(n34625), .B(n34294), .ZN(n33814) );
  NAND2_X1 U39440 ( .A1(n39479), .A2(n37804), .ZN(n39475) );
  XNOR2_X1 U39441 ( .A(n36939), .B(n34400), .ZN(n33816) );
  XNOR2_X1 U39442 ( .A(n33816), .B(n36681), .ZN(n33817) );
  XNOR2_X1 U39444 ( .A(n33818), .B(n33894), .ZN(n33819) );
  XNOR2_X1 U39445 ( .A(n33820), .B(n33819), .ZN(n33827) );
  INV_X1 U39446 ( .A(n33821), .ZN(n33823) );
  XNOR2_X1 U39447 ( .A(n33823), .B(n33822), .ZN(n33824) );
  XNOR2_X1 U39448 ( .A(n35255), .B(n33824), .ZN(n33825) );
  XNOR2_X1 U39449 ( .A(n33902), .B(n33825), .ZN(n33826) );
  XNOR2_X1 U39450 ( .A(n36858), .B(n51702), .ZN(n35249) );
  XNOR2_X1 U39451 ( .A(n35372), .B(n35249), .ZN(n33828) );
  XNOR2_X1 U39452 ( .A(n37062), .B(n34141), .ZN(n33830) );
  XNOR2_X1 U39453 ( .A(n33830), .B(n52148), .ZN(n34556) );
  XNOR2_X1 U39454 ( .A(n37243), .B(n33831), .ZN(n33832) );
  XNOR2_X1 U39455 ( .A(n33832), .B(n34556), .ZN(n33834) );
  XNOR2_X1 U39456 ( .A(n33834), .B(n33833), .ZN(n33842) );
  XNOR2_X1 U39457 ( .A(n35606), .B(n47679), .ZN(n33835) );
  XOR2_X1 U39458 ( .A(n4613), .B(n48814), .Z(n33836) );
  XNOR2_X1 U39459 ( .A(n33837), .B(n33836), .ZN(n33838) );
  XNOR2_X1 U39460 ( .A(n36934), .B(n33839), .ZN(n33840) );
  XNOR2_X1 U39461 ( .A(n33840), .B(n34737), .ZN(n33841) );
  XNOR2_X1 U39462 ( .A(n4537), .B(n4826), .ZN(n33843) );
  XNOR2_X1 U39463 ( .A(n2604), .B(n33843), .ZN(n33844) );
  XNOR2_X1 U39464 ( .A(n33845), .B(n33844), .ZN(n33846) );
  XNOR2_X1 U39465 ( .A(n41663), .B(n33846), .ZN(n33847) );
  XNOR2_X1 U39466 ( .A(n33973), .B(n33847), .ZN(n33849) );
  XNOR2_X1 U39467 ( .A(n33849), .B(n33848), .ZN(n33850) );
  XNOR2_X1 U39468 ( .A(n33853), .B(n34337), .ZN(n34102) );
  XNOR2_X1 U39469 ( .A(n33854), .B(n47401), .ZN(n33855) );
  XNOR2_X1 U39470 ( .A(n33856), .B(n33855), .ZN(n33857) );
  XNOR2_X1 U39471 ( .A(n35543), .B(n33858), .ZN(n33859) );
  XNOR2_X1 U39472 ( .A(n33859), .B(n34753), .ZN(n33861) );
  XNOR2_X1 U39473 ( .A(n33861), .B(n33860), .ZN(n33866) );
  XNOR2_X1 U39474 ( .A(n33864), .B(n33863), .ZN(n34120) );
  INV_X1 U39475 ( .A(n34120), .ZN(n33865) );
  XNOR2_X1 U39477 ( .A(n35632), .B(n37292), .ZN(n33867) );
  XNOR2_X1 U39478 ( .A(n34572), .B(n33867), .ZN(n34755) );
  XNOR2_X1 U39479 ( .A(n34110), .B(n34755), .ZN(n33868) );
  NOR2_X1 U39480 ( .A1(n39475), .A2(n473), .ZN(n34700) );
  OAI21_X1 U39481 ( .B1(n34700), .B2(n39471), .A(n37798), .ZN(n33875) );
  NAND2_X1 U39484 ( .A1(n34698), .A2(n39481), .ZN(n33874) );
  INV_X1 U39485 ( .A(n37798), .ZN(n38974) );
  NAND2_X1 U39486 ( .A1(n39474), .A2(n1075), .ZN(n33872) );
  OAI211_X1 U39487 ( .C1(n38974), .C2(n37802), .A(n39484), .B(n33872), .ZN(
        n33873) );
  NAND4_X1 U39488 ( .A1(n38988), .A2(n33875), .A3(n33874), .A4(n33873), .ZN(
        n33879) );
  NAND2_X1 U39489 ( .A1(n37802), .A2(n2177), .ZN(n36205) );
  NAND2_X1 U39490 ( .A1(n39474), .A2(n7159), .ZN(n33876) );
  NAND2_X1 U39491 ( .A1(n36205), .A2(n33876), .ZN(n33877) );
  NAND3_X1 U39492 ( .A1(n38815), .A2(n43669), .A3(n41796), .ZN(n33881) );
  INV_X1 U39493 ( .A(n38805), .ZN(n41802) );
  NAND3_X1 U39494 ( .A1(n41802), .A2(n51684), .A3(n51734), .ZN(n33880) );
  AND3_X1 U39495 ( .A1(n33882), .A2(n33881), .A3(n33880), .ZN(n33888) );
  OAI211_X1 U39497 ( .C1(n41794), .C2(n43669), .A(n51950), .B(n43665), .ZN(
        n33887) );
  NAND2_X1 U39498 ( .A1(n33883), .A2(n41794), .ZN(n33886) );
  AOI21_X1 U39499 ( .B1(n40639), .B2(n51734), .A(n51684), .ZN(n33884) );
  XNOR2_X1 U39500 ( .A(n33890), .B(n33889), .ZN(n33891) );
  XNOR2_X1 U39501 ( .A(n33892), .B(n33891), .ZN(n33907) );
  XNOR2_X1 U39502 ( .A(n33893), .B(n35255), .ZN(n34393) );
  XNOR2_X1 U39503 ( .A(n33894), .B(n4926), .ZN(n33895) );
  XNOR2_X1 U39504 ( .A(n34393), .B(n33895), .ZN(n34134) );
  INV_X1 U39505 ( .A(n33896), .ZN(n33898) );
  XNOR2_X1 U39506 ( .A(n33898), .B(n33897), .ZN(n33900) );
  XNOR2_X1 U39507 ( .A(n33900), .B(n33899), .ZN(n33901) );
  XNOR2_X1 U39508 ( .A(n34811), .B(n33901), .ZN(n33903) );
  XNOR2_X1 U39509 ( .A(n33903), .B(n33902), .ZN(n33904) );
  XNOR2_X1 U39510 ( .A(n33904), .B(n34824), .ZN(n33905) );
  XNOR2_X1 U39511 ( .A(n34134), .B(n33905), .ZN(n33906) );
  XNOR2_X1 U39512 ( .A(n33907), .B(n33906), .ZN(n34987) );
  INV_X1 U39513 ( .A(n34987), .ZN(n33994) );
  XNOR2_X1 U39514 ( .A(n33908), .B(n35265), .ZN(n33909) );
  XNOR2_X1 U39515 ( .A(n33909), .B(n51663), .ZN(n34387) );
  XNOR2_X1 U39516 ( .A(n34387), .B(n33910), .ZN(n33924) );
  XNOR2_X1 U39517 ( .A(n33911), .B(n36930), .ZN(n33913) );
  XNOR2_X1 U39518 ( .A(n34835), .B(n36841), .ZN(n33912) );
  XNOR2_X1 U39519 ( .A(n33913), .B(n33912), .ZN(n33921) );
  INV_X1 U39520 ( .A(n33914), .ZN(n33917) );
  XNOR2_X1 U39521 ( .A(n33915), .B(n49109), .ZN(n33916) );
  XNOR2_X1 U39522 ( .A(n33917), .B(n33916), .ZN(n33918) );
  XNOR2_X1 U39523 ( .A(n35606), .B(n33918), .ZN(n33919) );
  XNOR2_X1 U39524 ( .A(n33919), .B(n34553), .ZN(n33920) );
  XNOR2_X1 U39525 ( .A(n33921), .B(n33920), .ZN(n33922) );
  XNOR2_X1 U39526 ( .A(n37072), .B(n34739), .ZN(n36851) );
  XNOR2_X1 U39527 ( .A(n36851), .B(n33922), .ZN(n33923) );
  INV_X1 U39528 ( .A(n33925), .ZN(n33928) );
  INV_X1 U39529 ( .A(n33926), .ZN(n33927) );
  XNOR2_X1 U39530 ( .A(n36829), .B(n34881), .ZN(n33929) );
  XNOR2_X1 U39531 ( .A(n33929), .B(n33145), .ZN(n37021) );
  XNOR2_X1 U39532 ( .A(n33931), .B(n33930), .ZN(n33932) );
  XNOR2_X1 U39533 ( .A(n33933), .B(n33932), .ZN(n33936) );
  INV_X1 U39534 ( .A(n33934), .ZN(n33935) );
  XNOR2_X1 U39535 ( .A(n33936), .B(n33935), .ZN(n33937) );
  XNOR2_X1 U39536 ( .A(n33938), .B(n33937), .ZN(n33939) );
  XNOR2_X1 U39537 ( .A(n34604), .B(n36747), .ZN(n35753) );
  XNOR2_X1 U39538 ( .A(n33939), .B(n35753), .ZN(n33940) );
  XNOR2_X1 U39539 ( .A(n52221), .B(n33942), .ZN(n33944) );
  XNOR2_X1 U39540 ( .A(n36998), .B(n3383), .ZN(n36760) );
  XNOR2_X1 U39541 ( .A(n36760), .B(n33943), .ZN(n34898) );
  XNOR2_X1 U39542 ( .A(n33944), .B(n34898), .ZN(n33945) );
  XNOR2_X1 U39543 ( .A(n33946), .B(n33945), .ZN(n33957) );
  XNOR2_X1 U39544 ( .A(n34156), .B(n52071), .ZN(n33947) );
  XNOR2_X1 U39545 ( .A(n34896), .B(n33947), .ZN(n33948) );
  XNOR2_X1 U39546 ( .A(n34294), .B(n33948), .ZN(n34489) );
  XNOR2_X1 U39547 ( .A(n33949), .B(n35672), .ZN(n33950) );
  XNOR2_X1 U39548 ( .A(n33951), .B(n33950), .ZN(n33952) );
  XNOR2_X1 U39549 ( .A(n36992), .B(n33952), .ZN(n33954) );
  XNOR2_X1 U39550 ( .A(n33954), .B(n33953), .ZN(n33955) );
  XNOR2_X1 U39551 ( .A(n34489), .B(n33955), .ZN(n33956) );
  XNOR2_X1 U39552 ( .A(n33957), .B(n33956), .ZN(n37983) );
  AND2_X1 U39553 ( .A1(n594), .A2(n37987), .ZN(n36517) );
  NAND2_X1 U39554 ( .A1(n36519), .A2(n36517), .ZN(n36349) );
  AND2_X1 U39555 ( .A1(n5711), .A2(n37983), .ZN(n36077) );
  NAND2_X1 U39556 ( .A1(n36077), .A2(n37976), .ZN(n36073) );
  XNOR2_X1 U39558 ( .A(n33958), .B(n34433), .ZN(n35229) );
  XNOR2_X1 U39559 ( .A(n33960), .B(n33959), .ZN(n33961) );
  XNOR2_X1 U39560 ( .A(n35800), .B(n33961), .ZN(n33962) );
  XNOR2_X1 U39561 ( .A(n33963), .B(n33962), .ZN(n33964) );
  XNOR2_X1 U39562 ( .A(n34052), .B(n33964), .ZN(n33965) );
  XNOR2_X1 U39563 ( .A(n33965), .B(n35229), .ZN(n33971) );
  INV_X1 U39564 ( .A(n33966), .ZN(n33969) );
  XNOR2_X1 U39565 ( .A(n35632), .B(n47401), .ZN(n33967) );
  XNOR2_X1 U39566 ( .A(n515), .B(n34288), .ZN(n33968) );
  XNOR2_X1 U39567 ( .A(n33969), .B(n33968), .ZN(n33970) );
  XNOR2_X1 U39568 ( .A(n33971), .B(n33970), .ZN(n33995) );
  INV_X1 U39569 ( .A(n33995), .ZN(n37974) );
  XNOR2_X1 U39570 ( .A(n36811), .B(n4177), .ZN(n35822) );
  INV_X1 U39571 ( .A(n33973), .ZN(n33974) );
  XNOR2_X1 U39572 ( .A(n33974), .B(n34760), .ZN(n34862) );
  INV_X1 U39573 ( .A(n34862), .ZN(n33975) );
  XNOR2_X1 U39574 ( .A(n35822), .B(n33975), .ZN(n33976) );
  XNOR2_X1 U39575 ( .A(n34455), .B(n35618), .ZN(n34588) );
  XNOR2_X1 U39576 ( .A(n33976), .B(n34588), .ZN(n33985) );
  INV_X1 U39577 ( .A(n43564), .ZN(n33978) );
  XNOR2_X1 U39578 ( .A(n33978), .B(n33977), .ZN(n33979) );
  XNOR2_X1 U39579 ( .A(n51739), .B(n33979), .ZN(n33980) );
  XNOR2_X1 U39580 ( .A(n2168), .B(n33980), .ZN(n33982) );
  XNOR2_X1 U39581 ( .A(n51495), .B(n33982), .ZN(n33984) );
  XNOR2_X1 U39582 ( .A(n33985), .B(n33984), .ZN(n33992) );
  INV_X1 U39583 ( .A(n33986), .ZN(n33987) );
  XNOR2_X1 U39584 ( .A(n35331), .B(n33987), .ZN(n33988) );
  XNOR2_X1 U39585 ( .A(n33990), .B(n33989), .ZN(n35552) );
  XNOR2_X1 U39586 ( .A(n52197), .B(n35552), .ZN(n33991) );
  XNOR2_X1 U39587 ( .A(n33992), .B(n33991), .ZN(n34984) );
  INV_X1 U39588 ( .A(n34984), .ZN(n37988) );
  AND2_X1 U39589 ( .A1(n37975), .A2(n37987), .ZN(n33993) );
  NAND2_X1 U39590 ( .A1(n37988), .A2(n594), .ZN(n37982) );
  INV_X1 U39591 ( .A(n37982), .ZN(n37979) );
  AOI21_X1 U39592 ( .B1(n37991), .B2(n33993), .A(n37979), .ZN(n33998) );
  MUX2_X1 U39593 ( .A(n36518), .B(n37977), .S(n37980), .Z(n33996) );
  OAI21_X1 U39594 ( .B1(n33996), .B2(n37988), .A(n36080), .ZN(n33997) );
  XNOR2_X1 U39595 ( .A(n33999), .B(n34000), .ZN(n34011) );
  INV_X1 U39596 ( .A(n34001), .ZN(n35031) );
  INV_X1 U39597 ( .A(n34002), .ZN(n34005) );
  XNOR2_X1 U39598 ( .A(n34003), .B(n4908), .ZN(n34004) );
  XNOR2_X1 U39599 ( .A(n34005), .B(n34004), .ZN(n34006) );
  XNOR2_X1 U39600 ( .A(n37261), .B(n34006), .ZN(n34007) );
  XNOR2_X1 U39601 ( .A(n34007), .B(n619), .ZN(n34008) );
  XNOR2_X1 U39602 ( .A(n34008), .B(n36869), .ZN(n34009) );
  XNOR2_X1 U39603 ( .A(n35031), .B(n34009), .ZN(n34010) );
  XNOR2_X1 U39604 ( .A(n34011), .B(n34010), .ZN(n34089) );
  XNOR2_X1 U39606 ( .A(n36930), .B(n52148), .ZN(n34013) );
  XNOR2_X1 U39607 ( .A(n34216), .B(n4654), .ZN(n34014) );
  XNOR2_X1 U39608 ( .A(n34015), .B(n34014), .ZN(n34016) );
  XNOR2_X1 U39609 ( .A(n37062), .B(n34016), .ZN(n34017) );
  XNOR2_X1 U39610 ( .A(n34219), .B(n34017), .ZN(n34018) );
  XNOR2_X1 U39611 ( .A(n34019), .B(n34018), .ZN(n34022) );
  BUF_X2 U39613 ( .A(n34056), .Z(n36547) );
  XNOR2_X1 U39614 ( .A(n36722), .B(n34455), .ZN(n35809) );
  XNOR2_X1 U39615 ( .A(n35809), .B(n34862), .ZN(n34025) );
  XNOR2_X1 U39616 ( .A(n34025), .B(n34026), .ZN(n34036) );
  XNOR2_X1 U39617 ( .A(n33702), .B(n34869), .ZN(n34033) );
  XNOR2_X1 U39618 ( .A(n34028), .B(n34027), .ZN(n34029) );
  XNOR2_X1 U39619 ( .A(n34030), .B(n34029), .ZN(n34031) );
  XNOR2_X1 U39620 ( .A(n51739), .B(n34031), .ZN(n34032) );
  XNOR2_X1 U39621 ( .A(n34033), .B(n34032), .ZN(n34034) );
  XNOR2_X1 U39622 ( .A(n35627), .B(n34034), .ZN(n34035) );
  XNOR2_X1 U39623 ( .A(n34036), .B(n34035), .ZN(n34038) );
  XNOR2_X1 U39624 ( .A(n35825), .B(n34037), .ZN(n34873) );
  XNOR2_X1 U39625 ( .A(n34038), .B(n34873), .ZN(n34084) );
  XNOR2_X1 U39626 ( .A(n2129), .B(n35800), .ZN(n34039) );
  XNOR2_X1 U39627 ( .A(n34039), .B(n34351), .ZN(n34280) );
  XNOR2_X1 U39628 ( .A(n34041), .B(n34040), .ZN(n34042) );
  XNOR2_X1 U39629 ( .A(n34280), .B(n34042), .ZN(n34045) );
  XNOR2_X1 U39630 ( .A(n34044), .B(n34045), .ZN(n34055) );
  XNOR2_X1 U39631 ( .A(n34047), .B(n34046), .ZN(n34048) );
  XNOR2_X1 U39632 ( .A(n37086), .B(n34048), .ZN(n34049) );
  XNOR2_X1 U39633 ( .A(n35095), .B(n34049), .ZN(n34050) );
  XNOR2_X1 U39634 ( .A(n34051), .B(n34050), .ZN(n34053) );
  XNOR2_X1 U39635 ( .A(n34052), .B(n34053), .ZN(n34054) );
  NAND2_X1 U39636 ( .A1(n34084), .A2(n37969), .ZN(n36540) );
  INV_X1 U39637 ( .A(n34056), .ZN(n34090) );
  INV_X1 U39638 ( .A(n34057), .ZN(n44196) );
  XNOR2_X1 U39639 ( .A(n34891), .B(n4755), .ZN(n34058) );
  XNOR2_X1 U39640 ( .A(n34059), .B(n34058), .ZN(n34060) );
  XNOR2_X1 U39641 ( .A(n44196), .B(n34060), .ZN(n34061) );
  XNOR2_X1 U39642 ( .A(n35768), .B(n34061), .ZN(n34062) );
  XNOR2_X1 U39643 ( .A(n34063), .B(n34062), .ZN(n34064) );
  XNOR2_X1 U39644 ( .A(n34064), .B(n34294), .ZN(n34066) );
  XNOR2_X1 U39645 ( .A(n36873), .B(n36760), .ZN(n34065) );
  XNOR2_X1 U39646 ( .A(n34066), .B(n34065), .ZN(n34070) );
  XNOR2_X1 U39647 ( .A(n35482), .B(n52220), .ZN(n34068) );
  INV_X1 U39648 ( .A(n37323), .ZN(n34067) );
  XNOR2_X1 U39649 ( .A(n34068), .B(n34067), .ZN(n34364) );
  XNOR2_X1 U39650 ( .A(n34881), .B(n35105), .ZN(n34076) );
  INV_X1 U39651 ( .A(n34071), .ZN(n34073) );
  XNOR2_X1 U39652 ( .A(n34073), .B(n34072), .ZN(n34074) );
  XNOR2_X1 U39653 ( .A(n35468), .B(n34074), .ZN(n34075) );
  XNOR2_X1 U39654 ( .A(n34076), .B(n34075), .ZN(n34077) );
  XNOR2_X1 U39655 ( .A(n34078), .B(n35753), .ZN(n34260) );
  INV_X1 U39656 ( .A(n34260), .ZN(n34079) );
  XNOR2_X1 U39657 ( .A(n34169), .B(n34080), .ZN(n34081) );
  XNOR2_X1 U39658 ( .A(n34082), .B(n34081), .ZN(n34251) );
  INV_X1 U39659 ( .A(n34611), .ZN(n34083) );
  INV_X1 U39660 ( .A(n34084), .ZN(n36545) );
  NOR2_X1 U39661 ( .A1(n36547), .A2(n36027), .ZN(n34085) );
  NAND2_X1 U39662 ( .A1(n36553), .A2(n34085), .ZN(n37961) );
  OAI21_X1 U39663 ( .B1(n37962), .B2(n51077), .A(n37961), .ZN(n34087) );
  NAND2_X1 U39665 ( .A1(n36545), .A2(n699), .ZN(n36550) );
  AND2_X1 U39666 ( .A1(n36027), .A2(n36545), .ZN(n34997) );
  INV_X1 U39667 ( .A(n34997), .ZN(n36549) );
  NAND2_X1 U39668 ( .A1(n36542), .A2(n36549), .ZN(n34086) );
  NAND2_X1 U39669 ( .A1(n36029), .A2(n52156), .ZN(n34661) );
  INV_X1 U39670 ( .A(n34661), .ZN(n34088) );
  AND2_X1 U39671 ( .A1(n36027), .A2(n51077), .ZN(n36548) );
  OAI21_X1 U39672 ( .B1(n34090), .B2(n34088), .A(n36548), .ZN(n34091) );
  INV_X1 U39673 ( .A(n36540), .ZN(n37965) );
  AND2_X1 U39674 ( .A1(n36552), .A2(n51077), .ZN(n34093) );
  INV_X1 U39675 ( .A(n36553), .ZN(n34993) );
  NOR2_X1 U39676 ( .A1(n37964), .A2(n36550), .ZN(n34092) );
  NAND2_X1 U39677 ( .A1(n37964), .A2(n36027), .ZN(n36037) );
  AND2_X1 U39678 ( .A1(n36539), .A2(n699), .ZN(n36034) );
  NAND2_X1 U39679 ( .A1(n7117), .A2(n40341), .ZN(n34322) );
  INV_X1 U39680 ( .A(n34095), .ZN(n34098) );
  XNOR2_X1 U39681 ( .A(n34096), .B(n4177), .ZN(n34097) );
  XNOR2_X1 U39682 ( .A(n34098), .B(n34097), .ZN(n34099) );
  XNOR2_X1 U39683 ( .A(n36811), .B(n34099), .ZN(n34100) );
  XNOR2_X1 U39684 ( .A(n34101), .B(n34100), .ZN(n34103) );
  XNOR2_X1 U39685 ( .A(n34103), .B(n34102), .ZN(n34108) );
  INV_X1 U39686 ( .A(n34594), .ZN(n34331) );
  XNOR2_X1 U39687 ( .A(n34331), .B(n37277), .ZN(n34106) );
  XNOR2_X1 U39688 ( .A(n34104), .B(n35625), .ZN(n34105) );
  XNOR2_X1 U39689 ( .A(n34106), .B(n34105), .ZN(n34458) );
  XNOR2_X1 U39690 ( .A(n34263), .B(n34458), .ZN(n34107) );
  INV_X1 U39691 ( .A(n34357), .ZN(n34111) );
  INV_X1 U39692 ( .A(n42657), .ZN(n34114) );
  XNOR2_X1 U39693 ( .A(n34114), .B(n34113), .ZN(n34115) );
  XNOR2_X1 U39694 ( .A(n37086), .B(n34115), .ZN(n34117) );
  XNOR2_X1 U39695 ( .A(n34117), .B(n36701), .ZN(n34118) );
  XNOR2_X1 U39696 ( .A(n34288), .B(n34118), .ZN(n34119) );
  NAND2_X1 U39697 ( .A1(n36575), .A2(n36015), .ZN(n36495) );
  INV_X1 U39698 ( .A(n36495), .ZN(n36569) );
  INV_X1 U39699 ( .A(n34121), .ZN(n34545) );
  XNOR2_X1 U39700 ( .A(n36685), .B(n34545), .ZN(n34123) );
  XNOR2_X1 U39701 ( .A(n51501), .B(n34123), .ZN(n34499) );
  XNOR2_X1 U39702 ( .A(n35372), .B(n34499), .ZN(n34131) );
  INV_X1 U39703 ( .A(n34124), .ZN(n34126) );
  XNOR2_X1 U39704 ( .A(n34126), .B(n34125), .ZN(n34127) );
  XNOR2_X1 U39705 ( .A(n34491), .B(n34127), .ZN(n34129) );
  XNOR2_X1 U39706 ( .A(n34128), .B(n34129), .ZN(n34130) );
  XNOR2_X1 U39707 ( .A(n34132), .B(n34133), .ZN(n34244) );
  XNOR2_X1 U39708 ( .A(n34134), .B(n34244), .ZN(n34135) );
  NAND2_X1 U39709 ( .A1(n36569), .A2(n36571), .ZN(n36482) );
  XNOR2_X1 U39710 ( .A(n43314), .B(n34136), .ZN(n34137) );
  XNOR2_X1 U39711 ( .A(n45478), .B(n34137), .ZN(n34138) );
  XNOR2_X1 U39712 ( .A(n37062), .B(n34138), .ZN(n34139) );
  XNOR2_X1 U39713 ( .A(n52148), .B(n34139), .ZN(n34140) );
  XNOR2_X1 U39714 ( .A(n35778), .B(n4687), .ZN(n34469) );
  XNOR2_X1 U39715 ( .A(n34140), .B(n34469), .ZN(n34145) );
  XNOR2_X1 U39716 ( .A(n34141), .B(n34382), .ZN(n34142) );
  XNOR2_X1 U39717 ( .A(n34143), .B(n34142), .ZN(n34144) );
  XNOR2_X1 U39718 ( .A(n34144), .B(n34145), .ZN(n34148) );
  XNOR2_X1 U39719 ( .A(n36934), .B(n34146), .ZN(n34147) );
  XNOR2_X1 U39720 ( .A(n34148), .B(n34147), .ZN(n34150) );
  XNOR2_X1 U39721 ( .A(n35351), .B(n37237), .ZN(n34149) );
  INV_X1 U39723 ( .A(n36488), .ZN(n36562) );
  XNOR2_X1 U39724 ( .A(n37323), .B(n35764), .ZN(n34152) );
  XNOR2_X1 U39725 ( .A(n36764), .B(n34620), .ZN(n34484) );
  XNOR2_X1 U39726 ( .A(n34484), .B(n52219), .ZN(n34151) );
  XNOR2_X1 U39727 ( .A(n34153), .B(n36999), .ZN(n35126) );
  XNOR2_X1 U39728 ( .A(n44539), .B(n34154), .ZN(n34155) );
  XNOR2_X1 U39729 ( .A(n34156), .B(n34155), .ZN(n34158) );
  XNOR2_X1 U39730 ( .A(n34158), .B(n34157), .ZN(n34159) );
  XNOR2_X1 U39731 ( .A(n35126), .B(n34159), .ZN(n34160) );
  XNOR2_X1 U39732 ( .A(n34605), .B(n34163), .ZN(n34164) );
  XNOR2_X1 U39733 ( .A(n35386), .B(n34164), .ZN(n34172) );
  INV_X1 U39734 ( .A(n34165), .ZN(n34167) );
  XNOR2_X1 U39735 ( .A(n34167), .B(n34166), .ZN(n34168) );
  XNOR2_X1 U39736 ( .A(n34169), .B(n34168), .ZN(n34170) );
  XNOR2_X1 U39737 ( .A(n33303), .B(n34170), .ZN(n34171) );
  XNOR2_X1 U39738 ( .A(n34172), .B(n34171), .ZN(n34174) );
  XNOR2_X1 U39739 ( .A(n34425), .B(n34247), .ZN(n34173) );
  XNOR2_X1 U39740 ( .A(n34174), .B(n34173), .ZN(n34178) );
  INV_X1 U39741 ( .A(n35120), .ZN(n34177) );
  XNOR2_X1 U39742 ( .A(n34175), .B(n35296), .ZN(n34176) );
  INV_X1 U39743 ( .A(n36567), .ZN(n36492) );
  AND2_X1 U39744 ( .A1(n36493), .A2(n36567), .ZN(n36474) );
  OAI21_X1 U39745 ( .B1(n36572), .B2(n36474), .A(n36558), .ZN(n34179) );
  NAND3_X1 U39746 ( .A1(n36482), .A2(n36014), .A3(n34179), .ZN(n34180) );
  NAND2_X1 U39747 ( .A1(n34180), .A2(n36490), .ZN(n34183) );
  INV_X1 U39748 ( .A(n36561), .ZN(n34181) );
  NOR2_X1 U39749 ( .A1(n36570), .A2(n4246), .ZN(n36471) );
  INV_X1 U39751 ( .A(n35315), .ZN(n36576) );
  OR2_X1 U39752 ( .A1(n36472), .A2(n36495), .ZN(n35313) );
  INV_X1 U39753 ( .A(n35311), .ZN(n36019) );
  NAND2_X1 U39754 ( .A1(n36493), .A2(n63), .ZN(n34182) );
  NOR2_X1 U39755 ( .A1(n4246), .A2(n34182), .ZN(n36560) );
  NAND2_X1 U39756 ( .A1(n36639), .A2(n34184), .ZN(n34185) );
  NAND2_X1 U39757 ( .A1(n34188), .A2(n38073), .ZN(n34202) );
  INV_X1 U39758 ( .A(n36635), .ZN(n34194) );
  AND2_X1 U39759 ( .A1(n34189), .A2(n36313), .ZN(n38075) );
  OAI21_X1 U39760 ( .B1(n34194), .B2(n38075), .A(n34190), .ZN(n34191) );
  AND2_X1 U39761 ( .A1(n36628), .A2(n38094), .ZN(n34192) );
  NAND3_X1 U39762 ( .A1(n34191), .A2(n34192), .A3(n38086), .ZN(n34201) );
  AOI21_X1 U39763 ( .B1(n34192), .B2(n34963), .A(n38086), .ZN(n34196) );
  AND3_X1 U39764 ( .A1(n36313), .A2(n36312), .A3(n50984), .ZN(n36319) );
  INV_X1 U39765 ( .A(n34197), .ZN(n34198) );
  NOR2_X1 U39766 ( .A1(n52101), .A2(n40327), .ZN(n37868) );
  INV_X1 U39767 ( .A(n37868), .ZN(n34321) );
  INV_X1 U39768 ( .A(n36381), .ZN(n38038) );
  OAI21_X1 U39769 ( .B1(n38038), .B2(n36376), .A(n35157), .ZN(n34205) );
  AND2_X1 U39770 ( .A1(n36372), .A2(n35155), .ZN(n36380) );
  NOR2_X1 U39771 ( .A1(n35156), .A2(n38040), .ZN(n34203) );
  OAI21_X1 U39772 ( .B1(n34203), .B2(n35154), .A(n38027), .ZN(n34204) );
  INV_X1 U39773 ( .A(n35162), .ZN(n38028) );
  AOI22_X1 U39774 ( .A1(n34205), .A2(n36380), .B1(n34204), .B2(n38028), .ZN(
        n34214) );
  NOR2_X1 U39775 ( .A1(n38031), .A2(n34948), .ZN(n34944) );
  OAI21_X1 U39776 ( .B1(n36381), .B2(n35157), .A(n34944), .ZN(n34213) );
  NAND2_X1 U39777 ( .A1(n35156), .A2(n34945), .ZN(n34206) );
  NOR2_X1 U39778 ( .A1(n34207), .A2(n34206), .ZN(n36369) );
  NOR2_X1 U39779 ( .A1(n34948), .A2(n34208), .ZN(n34209) );
  OAI21_X1 U39780 ( .B1(n36369), .B2(n34209), .A(n38043), .ZN(n34212) );
  INV_X1 U39781 ( .A(n36383), .ZN(n34939) );
  NAND3_X1 U39782 ( .A1(n34939), .A2(n36381), .A3(n35159), .ZN(n34211) );
  XNOR2_X1 U39783 ( .A(n34216), .B(n34215), .ZN(n34217) );
  XNOR2_X1 U39784 ( .A(n34217), .B(n43267), .ZN(n34218) );
  XNOR2_X1 U39785 ( .A(n37065), .B(n34218), .ZN(n34220) );
  XNOR2_X1 U39786 ( .A(n34219), .B(n34220), .ZN(n34222) );
  XNOR2_X1 U39787 ( .A(n34222), .B(n34221), .ZN(n34228) );
  XNOR2_X1 U39788 ( .A(n36669), .B(n34381), .ZN(n34226) );
  INV_X1 U39789 ( .A(n35059), .ZN(n34224) );
  XNOR2_X1 U39790 ( .A(n34224), .B(n36841), .ZN(n34225) );
  XNOR2_X1 U39791 ( .A(n34226), .B(n34225), .ZN(n34227) );
  XNOR2_X1 U39792 ( .A(n34228), .B(n34227), .ZN(n34229) );
  XNOR2_X1 U39793 ( .A(n34233), .B(n34232), .ZN(n43607) );
  XNOR2_X1 U39794 ( .A(n34234), .B(n4788), .ZN(n34235) );
  XNOR2_X1 U39795 ( .A(n43607), .B(n34235), .ZN(n34236) );
  XNOR2_X1 U39796 ( .A(n34546), .B(n34236), .ZN(n34237) );
  XNOR2_X1 U39797 ( .A(n34238), .B(n34237), .ZN(n34241) );
  INV_X1 U39798 ( .A(n35841), .ZN(n34239) );
  XNOR2_X1 U39799 ( .A(n34240), .B(n34239), .ZN(n34498) );
  XNOR2_X1 U39800 ( .A(n34241), .B(n34498), .ZN(n34242) );
  XNOR2_X1 U39801 ( .A(n34724), .B(n34242), .ZN(n34246) );
  XNOR2_X1 U39802 ( .A(n34533), .B(n35255), .ZN(n36692) );
  XNOR2_X1 U39803 ( .A(n36692), .B(n704), .ZN(n34243) );
  XNOR2_X1 U39804 ( .A(n34244), .B(n34243), .ZN(n34245) );
  XNOR2_X1 U39805 ( .A(n34246), .B(n34245), .ZN(n34649) );
  XNOR2_X1 U39806 ( .A(n35471), .B(n36818), .ZN(n34250) );
  XNOR2_X1 U39807 ( .A(n34247), .B(n34248), .ZN(n34249) );
  XNOR2_X1 U39808 ( .A(n34252), .B(n42816), .ZN(n34253) );
  XNOR2_X1 U39809 ( .A(n34254), .B(n34253), .ZN(n34256) );
  XNOR2_X1 U39810 ( .A(n34256), .B(n34255), .ZN(n34257) );
  XNOR2_X1 U39811 ( .A(n35115), .B(n34257), .ZN(n34258) );
  XNOR2_X1 U39812 ( .A(n34258), .B(n36748), .ZN(n34259) );
  XNOR2_X1 U39813 ( .A(n35285), .B(n34259), .ZN(n34261) );
  XNOR2_X1 U39814 ( .A(n34261), .B(n34260), .ZN(n34262) );
  XNOR2_X1 U39815 ( .A(n34264), .B(n34263), .ZN(n34274) );
  XNOR2_X1 U39816 ( .A(n34266), .B(n34265), .ZN(n34267) );
  XNOR2_X1 U39817 ( .A(n34268), .B(n34267), .ZN(n34269) );
  XNOR2_X1 U39818 ( .A(n37113), .B(n34269), .ZN(n34270) );
  XNOR2_X1 U39819 ( .A(n36811), .B(n34270), .ZN(n34271) );
  XNOR2_X1 U39820 ( .A(n34272), .B(n34271), .ZN(n34273) );
  XNOR2_X1 U39821 ( .A(n34273), .B(n34274), .ZN(n34278) );
  INV_X1 U39822 ( .A(n36807), .ZN(n34276) );
  XNOR2_X1 U39823 ( .A(n51497), .B(n34276), .ZN(n34277) );
  XNOR2_X1 U39824 ( .A(n34277), .B(n35077), .ZN(n34771) );
  XNOR2_X1 U39825 ( .A(n35080), .B(n35537), .ZN(n34279) );
  XNOR2_X1 U39826 ( .A(n51449), .B(n34279), .ZN(n34281) );
  XNOR2_X1 U39827 ( .A(n34281), .B(n34280), .ZN(n34282) );
  XNOR2_X1 U39828 ( .A(n34282), .B(n36714), .ZN(n34293) );
  INV_X1 U39829 ( .A(n43694), .ZN(n34285) );
  XNOR2_X1 U39830 ( .A(n34283), .B(n43702), .ZN(n34284) );
  XNOR2_X1 U39831 ( .A(n34285), .B(n34284), .ZN(n34286) );
  XNOR2_X1 U39832 ( .A(n35536), .B(n34286), .ZN(n34287) );
  XNOR2_X1 U39833 ( .A(n34572), .B(n34287), .ZN(n34289) );
  XNOR2_X1 U39834 ( .A(n34288), .B(n34289), .ZN(n34291) );
  INV_X1 U39835 ( .A(n43293), .ZN(n43220) );
  XNOR2_X1 U39836 ( .A(n35095), .B(n43220), .ZN(n36707) );
  XNOR2_X1 U39837 ( .A(n37081), .B(n35085), .ZN(n34579) );
  XNOR2_X1 U39838 ( .A(n36707), .B(n34579), .ZN(n34290) );
  XNOR2_X1 U39839 ( .A(n34291), .B(n34290), .ZN(n34292) );
  NAND2_X1 U39840 ( .A1(n6276), .A2(n51015), .ZN(n36062) );
  INV_X1 U39841 ( .A(n36614), .ZN(n36066) );
  NAND2_X1 U39842 ( .A1(n36062), .A2(n36428), .ZN(n36622) );
  NAND2_X1 U39843 ( .A1(n36622), .A2(n36606), .ZN(n34309) );
  INV_X1 U39844 ( .A(n34896), .ZN(n34295) );
  XNOR2_X1 U39845 ( .A(n34296), .B(n34295), .ZN(n35278) );
  XOR2_X1 U39846 ( .A(n4665), .B(n4578), .Z(n34297) );
  XNOR2_X1 U39847 ( .A(n34298), .B(n34297), .ZN(n34299) );
  XNOR2_X1 U39848 ( .A(n34300), .B(n34299), .ZN(n34301) );
  XNOR2_X1 U39849 ( .A(n34369), .B(n34301), .ZN(n34302) );
  XNOR2_X1 U39850 ( .A(n34302), .B(n35483), .ZN(n34303) );
  XNOR2_X1 U39851 ( .A(n35126), .B(n34303), .ZN(n34304) );
  INV_X1 U39852 ( .A(n35404), .ZN(n34306) );
  XNOR2_X1 U39853 ( .A(n34306), .B(n34305), .ZN(n34307) );
  AOI21_X1 U39854 ( .B1(n36623), .B2(n34309), .A(n36427), .ZN(n34318) );
  INV_X1 U39855 ( .A(n51715), .ZN(n34650) );
  AND2_X1 U39856 ( .A1(n36428), .A2(n51015), .ZN(n34931) );
  INV_X1 U39857 ( .A(n34931), .ZN(n34310) );
  NAND2_X1 U39858 ( .A1(n34311), .A2(n34310), .ZN(n34312) );
  NAND2_X1 U39859 ( .A1(n34312), .A2(n34930), .ZN(n34316) );
  NAND2_X1 U39860 ( .A1(n34313), .A2(n36428), .ZN(n34314) );
  OAI211_X1 U39861 ( .C1(n36606), .C2(n34648), .A(n34314), .B(n36604), .ZN(
        n34315) );
  NAND2_X1 U39862 ( .A1(n34316), .A2(n34315), .ZN(n34317) );
  NAND2_X1 U39863 ( .A1(n40328), .A2(n52101), .ZN(n34319) );
  NAND3_X1 U39864 ( .A1(n34319), .A2(n40330), .A3(n40340), .ZN(n34320) );
  INV_X1 U39865 ( .A(n34323), .ZN(n34329) );
  AND2_X1 U39866 ( .A1(n40327), .A2(n40330), .ZN(n40335) );
  OAI21_X1 U39867 ( .B1(n40335), .B2(n40340), .A(n34324), .ZN(n34328) );
  NAND2_X1 U39868 ( .A1(n40341), .A2(n40330), .ZN(n38851) );
  INV_X1 U39869 ( .A(n38851), .ZN(n34325) );
  NAND2_X1 U39870 ( .A1(n39857), .A2(n40338), .ZN(n37869) );
  INV_X1 U39871 ( .A(n37869), .ZN(n39640) );
  NAND2_X1 U39872 ( .A1(n39855), .A2(n40327), .ZN(n37862) );
  NAND4_X1 U39873 ( .A1(n40337), .A2(n39640), .A3(n52101), .A4(n37862), .ZN(
        n34326) );
  XNOR2_X1 U39874 ( .A(n46128), .B(n4618), .ZN(n34330) );
  XNOR2_X1 U39875 ( .A(n34333), .B(n34332), .ZN(n34334) );
  XNOR2_X1 U39876 ( .A(n51739), .B(n34334), .ZN(n34335) );
  XNOR2_X1 U39877 ( .A(n34336), .B(n34335), .ZN(n34338) );
  XNOR2_X1 U39878 ( .A(n34337), .B(n34338), .ZN(n34340) );
  XNOR2_X1 U39879 ( .A(n37269), .B(n35334), .ZN(n34339) );
  XNOR2_X1 U39880 ( .A(n34339), .B(n37096), .ZN(n36800) );
  XNOR2_X1 U39881 ( .A(n34346), .B(n34345), .ZN(n34347) );
  XNOR2_X1 U39882 ( .A(n35536), .B(n34347), .ZN(n34348) );
  XNOR2_X1 U39883 ( .A(n34434), .B(n34348), .ZN(n34349) );
  XNOR2_X1 U39884 ( .A(n34350), .B(n34349), .ZN(n34354) );
  XNOR2_X1 U39885 ( .A(n37086), .B(n34844), .ZN(n34352) );
  XNOR2_X1 U39886 ( .A(n34352), .B(n34351), .ZN(n34353) );
  XNOR2_X1 U39887 ( .A(n34353), .B(n35534), .ZN(n36975) );
  XNOR2_X1 U39888 ( .A(n34354), .B(n36975), .ZN(n34358) );
  XNOR2_X1 U39889 ( .A(n36981), .B(n4817), .ZN(n36793) );
  XNOR2_X1 U39890 ( .A(n37081), .B(n36793), .ZN(n34356) );
  XNOR2_X1 U39891 ( .A(n515), .B(n34356), .ZN(n36713) );
  XNOR2_X1 U39893 ( .A(n37324), .B(n34361), .ZN(n34482) );
  XNOR2_X1 U39894 ( .A(n35669), .B(n34482), .ZN(n34362) );
  XNOR2_X1 U39895 ( .A(n36993), .B(n34362), .ZN(n34363) );
  XNOR2_X1 U39896 ( .A(n34363), .B(n34364), .ZN(n34375) );
  INV_X1 U39897 ( .A(n34365), .ZN(n34367) );
  XNOR2_X1 U39898 ( .A(n34367), .B(n34366), .ZN(n34368) );
  XNOR2_X1 U39899 ( .A(n34369), .B(n34368), .ZN(n34370) );
  XNOR2_X1 U39900 ( .A(n34370), .B(n35483), .ZN(n34371) );
  XNOR2_X1 U39901 ( .A(n35680), .B(n34371), .ZN(n34373) );
  XNOR2_X1 U39902 ( .A(n34373), .B(n34372), .ZN(n34374) );
  XNOR2_X1 U39903 ( .A(n34375), .B(n34374), .ZN(n35215) );
  INV_X1 U39904 ( .A(n34376), .ZN(n34559) );
  XNOR2_X1 U39905 ( .A(n34559), .B(n34377), .ZN(n34378) );
  XNOR2_X1 U39906 ( .A(n34379), .B(n34378), .ZN(n34380) );
  XNOR2_X1 U39907 ( .A(n34381), .B(n34380), .ZN(n34383) );
  XNOR2_X1 U39908 ( .A(n34383), .B(n34382), .ZN(n34384) );
  XNOR2_X1 U39909 ( .A(n52117), .B(n1341), .ZN(n34385) );
  XNOR2_X1 U39910 ( .A(n34466), .B(n34385), .ZN(n35358) );
  XNOR2_X1 U39911 ( .A(n34386), .B(n35358), .ZN(n34388) );
  XNOR2_X1 U39912 ( .A(n34387), .B(n34388), .ZN(n34390) );
  NAND3_X1 U39913 ( .A1(n36454), .A2(n36590), .A3(n35879), .ZN(n34391) );
  NAND3_X1 U39914 ( .A1(n35214), .A2(n36457), .A3(n34391), .ZN(n34409) );
  XNOR2_X1 U39915 ( .A(n34393), .B(n51702), .ZN(n34395) );
  XNOR2_X1 U39916 ( .A(n36940), .B(n4836), .ZN(n35366) );
  XNOR2_X1 U39917 ( .A(n35501), .B(n35830), .ZN(n34396) );
  XNOR2_X1 U39918 ( .A(n35366), .B(n34396), .ZN(n34404) );
  XNOR2_X1 U39919 ( .A(n34398), .B(n34397), .ZN(n34399) );
  XNOR2_X1 U39920 ( .A(n34400), .B(n34399), .ZN(n34401) );
  XNOR2_X1 U39921 ( .A(n34402), .B(n34401), .ZN(n34403) );
  XNOR2_X1 U39922 ( .A(n34403), .B(n34404), .ZN(n34406) );
  XNOR2_X1 U39923 ( .A(n34406), .B(n34405), .ZN(n34407) );
  AND2_X1 U39925 ( .A1(n35209), .A2(n34409), .ZN(n34428) );
  INV_X1 U39928 ( .A(n36585), .ZN(n36048) );
  XNOR2_X1 U39929 ( .A(n2131), .B(n34412), .ZN(n34418) );
  XNOR2_X1 U39930 ( .A(n42083), .B(n34414), .ZN(n34415) );
  XNOR2_X1 U39931 ( .A(n44135), .B(n34415), .ZN(n34416) );
  XNOR2_X1 U39932 ( .A(n34504), .B(n34416), .ZN(n34417) );
  XNOR2_X1 U39933 ( .A(n34418), .B(n34417), .ZN(n34419) );
  INV_X1 U39934 ( .A(n4666), .ZN(n34420) );
  XNOR2_X1 U39935 ( .A(n34514), .B(n34420), .ZN(n35374) );
  XNOR2_X1 U39936 ( .A(n34421), .B(n35374), .ZN(n34422) );
  XNOR2_X1 U39937 ( .A(n34423), .B(n34422), .ZN(n34427) );
  XNOR2_X1 U39938 ( .A(n36748), .B(n34424), .ZN(n34426) );
  XNOR2_X1 U39939 ( .A(n34425), .B(n34426), .ZN(n34607) );
  NAND2_X1 U39940 ( .A1(n36595), .A2(n35215), .ZN(n35204) );
  INV_X1 U39941 ( .A(n35204), .ZN(n35212) );
  NAND4_X1 U39942 ( .A1(n35212), .A2(n36590), .A3(n36459), .A4(n36050), .ZN(
        n34431) );
  NOR2_X1 U39943 ( .A1(n36462), .A2(n36050), .ZN(n35217) );
  INV_X1 U39944 ( .A(n35217), .ZN(n36600) );
  OR2_X1 U39945 ( .A1(n35880), .A2(n36045), .ZN(n36580) );
  INV_X1 U39946 ( .A(n36595), .ZN(n34429) );
  INV_X1 U39948 ( .A(n36592), .ZN(n36046) );
  NAND3_X1 U39949 ( .A1(n36581), .A2(n34429), .A3(n36046), .ZN(n34430) );
  XNOR2_X1 U39951 ( .A(n34433), .B(n36701), .ZN(n34438) );
  XNOR2_X1 U39952 ( .A(n34436), .B(n34435), .ZN(n34437) );
  XNOR2_X1 U39953 ( .A(n34440), .B(n34439), .ZN(n34441) );
  XNOR2_X1 U39954 ( .A(n51449), .B(n34441), .ZN(n34444) );
  XNOR2_X1 U39955 ( .A(n43702), .B(n4589), .ZN(n34442) );
  XNOR2_X1 U39956 ( .A(n35536), .B(n34442), .ZN(n34443) );
  XNOR2_X1 U39957 ( .A(n34443), .B(n35537), .ZN(n35648) );
  XNOR2_X1 U39958 ( .A(n34444), .B(n35648), .ZN(n34445) );
  XNOR2_X1 U39959 ( .A(n34569), .B(n34445), .ZN(n34449) );
  XNOR2_X1 U39960 ( .A(n34446), .B(n35086), .ZN(n34447) );
  XNOR2_X1 U39961 ( .A(n36714), .B(n34447), .ZN(n35230) );
  XNOR2_X1 U39962 ( .A(n34451), .B(n34450), .ZN(n34452) );
  XNOR2_X1 U39963 ( .A(n34455), .B(n35333), .ZN(n34456) );
  XNOR2_X1 U39964 ( .A(n51739), .B(n2204), .ZN(n35557) );
  XNOR2_X1 U39965 ( .A(n34456), .B(n35557), .ZN(n34457) );
  INV_X1 U39967 ( .A(n34462), .ZN(n34464) );
  XNOR2_X1 U39968 ( .A(n34464), .B(n34463), .ZN(n34465) );
  XNOR2_X1 U39969 ( .A(n35059), .B(n34465), .ZN(n34467) );
  XNOR2_X1 U39970 ( .A(n34466), .B(n34467), .ZN(n34468) );
  XNOR2_X1 U39971 ( .A(n34469), .B(n34468), .ZN(n34473) );
  XNOR2_X1 U39972 ( .A(n4737), .B(n4518), .ZN(n34470) );
  XNOR2_X1 U39973 ( .A(n35522), .B(n34470), .ZN(n35779) );
  XNOR2_X1 U39974 ( .A(n34471), .B(n35779), .ZN(n34472) );
  XNOR2_X1 U39975 ( .A(n34473), .B(n34472), .ZN(n34475) );
  XNOR2_X1 U39976 ( .A(n36680), .B(n34475), .ZN(n34478) );
  INV_X1 U39977 ( .A(n34476), .ZN(n34477) );
  XNOR2_X1 U39979 ( .A(n34480), .B(n34479), .ZN(n34481) );
  XNOR2_X1 U39980 ( .A(n35762), .B(n34481), .ZN(n34483) );
  XNOR2_X1 U39981 ( .A(n34483), .B(n34482), .ZN(n34486) );
  XNOR2_X1 U39982 ( .A(n34484), .B(n36766), .ZN(n34485) );
  XNOR2_X1 U39983 ( .A(n34486), .B(n34485), .ZN(n34487) );
  XNOR2_X1 U39984 ( .A(n35669), .B(n460), .ZN(n34488) );
  XNOR2_X1 U39985 ( .A(n34489), .B(n34488), .ZN(n34490) );
  XNOR2_X1 U39986 ( .A(n33335), .B(n34492), .ZN(n34493) );
  XNOR2_X1 U39987 ( .A(n34493), .B(n34535), .ZN(n35600) );
  XNOR2_X1 U39988 ( .A(n35600), .B(n35260), .ZN(n34502) );
  XNOR2_X1 U39989 ( .A(n34495), .B(n34494), .ZN(n34496) );
  XNOR2_X1 U39990 ( .A(n35830), .B(n34496), .ZN(n34497) );
  XNOR2_X1 U39991 ( .A(n34498), .B(n34497), .ZN(n34500) );
  XNOR2_X1 U39992 ( .A(n34500), .B(n34499), .ZN(n34501) );
  INV_X1 U39993 ( .A(n34529), .ZN(n38271) );
  XNOR2_X1 U39994 ( .A(n35289), .B(n34503), .ZN(n34506) );
  INV_X1 U39995 ( .A(n34504), .ZN(n35752) );
  XNOR2_X1 U39996 ( .A(n35752), .B(n34604), .ZN(n34505) );
  XNOR2_X1 U39997 ( .A(n34505), .B(n34506), .ZN(n34517) );
  INV_X1 U39998 ( .A(n34507), .ZN(n34512) );
  XNOR2_X1 U39999 ( .A(n34508), .B(n4940), .ZN(n34509) );
  XNOR2_X1 U40000 ( .A(n34509), .B(n42816), .ZN(n34510) );
  XNOR2_X1 U40001 ( .A(n34510), .B(n41828), .ZN(n34511) );
  XNOR2_X1 U40002 ( .A(n34512), .B(n34511), .ZN(n34513) );
  XNOR2_X1 U40003 ( .A(n37303), .B(n34513), .ZN(n34515) );
  XNOR2_X1 U40004 ( .A(n34514), .B(n34515), .ZN(n34516) );
  XNOR2_X1 U40005 ( .A(n34517), .B(n34516), .ZN(n34518) );
  XNOR2_X1 U40006 ( .A(n34518), .B(n35296), .ZN(n34521) );
  XNOR2_X1 U40007 ( .A(n33303), .B(n34519), .ZN(n34520) );
  XNOR2_X1 U40008 ( .A(n35471), .B(n34520), .ZN(n36751) );
  XNOR2_X1 U40009 ( .A(n34521), .B(n36751), .ZN(n34523) );
  INV_X1 U40010 ( .A(n34522), .ZN(n35664) );
  NAND3_X1 U40011 ( .A1(n37617), .A2(n38272), .A3(n38279), .ZN(n34524) );
  NAND2_X1 U40012 ( .A1(n2123), .A2(n38270), .ZN(n37623) );
  NAND4_X1 U40013 ( .A1(n34524), .A2(n2120), .A3(n613), .A4(n35866), .ZN(
        n34526) );
  XNOR2_X1 U40014 ( .A(n34529), .B(n38282), .ZN(n34525) );
  INV_X1 U40015 ( .A(n35416), .ZN(n37620) );
  OR2_X1 U40016 ( .A1(n37617), .A2(n37623), .ZN(n35420) );
  INV_X1 U40017 ( .A(n35420), .ZN(n37631) );
  OAI22_X1 U40018 ( .A1(n38290), .A2(n51339), .B1(n37629), .B2(n38270), .ZN(
        n34527) );
  OAI21_X1 U40019 ( .B1(n37631), .B2(n34527), .A(n38292), .ZN(n34531) );
  NAND2_X1 U40020 ( .A1(n38277), .A2(n38270), .ZN(n38288) );
  MUX2_X1 U40021 ( .A(n37630), .B(n38288), .S(n36436), .Z(n34530) );
  XNOR2_X1 U40022 ( .A(n34533), .B(n2203), .ZN(n34534) );
  XNOR2_X1 U40023 ( .A(n34534), .B(n619), .ZN(n37052) );
  XNOR2_X1 U40024 ( .A(n34535), .B(n37052), .ZN(n34543) );
  XNOR2_X1 U40025 ( .A(n35841), .B(n35830), .ZN(n34541) );
  INV_X1 U40026 ( .A(n34536), .ZN(n34538) );
  XNOR2_X1 U40027 ( .A(n42329), .B(n35251), .ZN(n34537) );
  XNOR2_X1 U40028 ( .A(n34538), .B(n34537), .ZN(n34539) );
  XNOR2_X1 U40029 ( .A(n35254), .B(n34539), .ZN(n34540) );
  XNOR2_X1 U40030 ( .A(n34541), .B(n34540), .ZN(n34542) );
  XNOR2_X1 U40031 ( .A(n34543), .B(n34542), .ZN(n34550) );
  XNOR2_X1 U40032 ( .A(n376), .B(n34545), .ZN(n34548) );
  XOR2_X1 U40033 ( .A(n34546), .B(n35829), .Z(n34547) );
  XNOR2_X1 U40034 ( .A(n34548), .B(n34547), .ZN(n34549) );
  XNOR2_X1 U40036 ( .A(n34550), .B(n35494), .ZN(n34551) );
  XNOR2_X1 U40037 ( .A(n34551), .B(n34552), .ZN(n34628) );
  XNOR2_X1 U40038 ( .A(n33195), .B(n34553), .ZN(n34554) );
  XNOR2_X1 U40039 ( .A(n34556), .B(n34557), .ZN(n34566) );
  XNOR2_X1 U40040 ( .A(n34559), .B(n34558), .ZN(n34561) );
  INV_X1 U40041 ( .A(n43768), .ZN(n34560) );
  XNOR2_X1 U40042 ( .A(n34561), .B(n34560), .ZN(n34562) );
  XNOR2_X1 U40043 ( .A(n37065), .B(n34562), .ZN(n34563) );
  XNOR2_X1 U40044 ( .A(n35778), .B(n34563), .ZN(n34564) );
  XNOR2_X1 U40045 ( .A(n35514), .B(n34564), .ZN(n34565) );
  XNOR2_X1 U40046 ( .A(n34567), .B(n34839), .ZN(n34568) );
  NAND2_X1 U40047 ( .A1(n34628), .A2(n37636), .ZN(n36000) );
  XNOR2_X1 U40048 ( .A(n36981), .B(n34570), .ZN(n34571) );
  XNOR2_X1 U40049 ( .A(n35224), .B(n34571), .ZN(n34573) );
  XNOR2_X1 U40050 ( .A(n34573), .B(n34572), .ZN(n34574) );
  XNOR2_X1 U40051 ( .A(n37288), .B(n34575), .ZN(n36976) );
  XNOR2_X1 U40052 ( .A(n36976), .B(n43968), .ZN(n34576) );
  XNOR2_X1 U40053 ( .A(n37476), .B(n34576), .ZN(n34577) );
  XNOR2_X1 U40054 ( .A(n35537), .B(n34577), .ZN(n34578) );
  XNOR2_X1 U40055 ( .A(n34579), .B(n34578), .ZN(n34580) );
  XNOR2_X1 U40056 ( .A(n34580), .B(n34754), .ZN(n34581) );
  XNOR2_X1 U40057 ( .A(n35549), .B(n34581), .ZN(n34582) );
  INV_X1 U40058 ( .A(n34584), .ZN(n34600) );
  XNOR2_X1 U40059 ( .A(n51445), .B(n35237), .ZN(n34586) );
  XNOR2_X1 U40060 ( .A(n37113), .B(n35625), .ZN(n34585) );
  XNOR2_X1 U40061 ( .A(n34586), .B(n34585), .ZN(n34587) );
  XNOR2_X1 U40062 ( .A(n34588), .B(n34587), .ZN(n34598) );
  INV_X1 U40063 ( .A(n34589), .ZN(n34592) );
  XNOR2_X1 U40064 ( .A(n34590), .B(n4537), .ZN(n34591) );
  XNOR2_X1 U40065 ( .A(n34592), .B(n34591), .ZN(n34593) );
  XNOR2_X1 U40066 ( .A(n33702), .B(n34593), .ZN(n34595) );
  XNOR2_X1 U40067 ( .A(n34594), .B(n34595), .ZN(n34596) );
  XNOR2_X1 U40068 ( .A(n34598), .B(n34597), .ZN(n34599) );
  INV_X1 U40069 ( .A(n34601), .ZN(n41479) );
  XNOR2_X1 U40070 ( .A(n34602), .B(n41479), .ZN(n34603) );
  XNOR2_X1 U40071 ( .A(n35752), .B(n34605), .ZN(n36817) );
  XNOR2_X1 U40072 ( .A(n35285), .B(n34609), .ZN(n34610) );
  INV_X1 U40074 ( .A(n34613), .ZN(n34618) );
  XNOR2_X1 U40075 ( .A(n34614), .B(n4755), .ZN(n34615) );
  XNOR2_X1 U40076 ( .A(n34616), .B(n34615), .ZN(n34617) );
  XNOR2_X1 U40077 ( .A(n34618), .B(n34617), .ZN(n34619) );
  XNOR2_X1 U40078 ( .A(n34620), .B(n34619), .ZN(n34621) );
  XNOR2_X1 U40079 ( .A(n34622), .B(n34621), .ZN(n34623) );
  XNOR2_X1 U40080 ( .A(n35133), .B(n37324), .ZN(n34624) );
  XNOR2_X1 U40081 ( .A(n34624), .B(n52221), .ZN(n35760) );
  XNOR2_X1 U40082 ( .A(n34626), .B(n35490), .ZN(n34627) );
  OAI22_X1 U40083 ( .A1(n35728), .A2(n36405), .B1(n36410), .B2(n34632), .ZN(
        n34639) );
  INV_X1 U40084 ( .A(n34628), .ZN(n37647) );
  NAND2_X1 U40085 ( .A1(n37647), .A2(n37636), .ZN(n35736) );
  INV_X1 U40086 ( .A(n35728), .ZN(n36402) );
  AND2_X1 U40087 ( .A1(n36405), .A2(n37646), .ZN(n36397) );
  OAI21_X1 U40088 ( .B1(n35736), .B2(n36402), .A(n36397), .ZN(n34638) );
  INV_X1 U40089 ( .A(n37636), .ZN(n35732) );
  INV_X1 U40090 ( .A(n36396), .ZN(n34630) );
  NAND2_X1 U40091 ( .A1(n51334), .A2(n36414), .ZN(n35194) );
  INV_X1 U40092 ( .A(n35194), .ZN(n34631) );
  NAND2_X1 U40093 ( .A1(n34631), .A2(n36410), .ZN(n34636) );
  AOI21_X1 U40094 ( .B1(n37647), .B2(n35728), .A(n51334), .ZN(n34634) );
  NAND2_X1 U40095 ( .A1(n37637), .A2(n35732), .ZN(n34633) );
  NAND2_X1 U40096 ( .A1(n51324), .A2(n36557), .ZN(n36494) );
  AOI22_X1 U40097 ( .A1(n36561), .A2(n36494), .B1(n36565), .B2(n458), .ZN(
        n34644) );
  NAND2_X1 U40098 ( .A1(n34641), .A2(n36567), .ZN(n34643) );
  NAND3_X1 U40099 ( .A1(n36558), .A2(n36565), .A3(n36492), .ZN(n34642) );
  NAND2_X1 U40100 ( .A1(n39712), .A2(n41079), .ZN(n39141) );
  NAND3_X1 U40101 ( .A1(n34928), .A2(n698), .A3(n34656), .ZN(n34646) );
  NAND2_X1 U40102 ( .A1(n36614), .A2(n34656), .ZN(n36424) );
  NAND2_X1 U40103 ( .A1(n51717), .A2(n34649), .ZN(n36420) );
  AND2_X1 U40104 ( .A1(n36420), .A2(n51015), .ZN(n36058) );
  NOR2_X1 U40105 ( .A1(n36424), .A2(n36058), .ZN(n34647) );
  NAND2_X1 U40106 ( .A1(n34650), .A2(n36430), .ZN(n36057) );
  NAND2_X1 U40107 ( .A1(n34650), .A2(n34649), .ZN(n36610) );
  NAND2_X1 U40108 ( .A1(n36606), .A2(n36610), .ZN(n34927) );
  AND2_X1 U40109 ( .A1(n34656), .A2(n36428), .ZN(n36618) );
  NAND2_X1 U40110 ( .A1(n36618), .A2(n36430), .ZN(n34651) );
  OAI22_X1 U40111 ( .A1(n34651), .A2(n36062), .B1(n36611), .B2(n51015), .ZN(
        n34652) );
  AOI21_X1 U40112 ( .B1(n34929), .B2(n34927), .A(n34652), .ZN(n34658) );
  NAND3_X1 U40113 ( .A1(n34930), .A2(n36428), .A3(n36067), .ZN(n34654) );
  INV_X1 U40114 ( .A(n36425), .ZN(n36065) );
  NAND2_X1 U40115 ( .A1(n34923), .A2(n36426), .ZN(n34657) );
  NOR2_X1 U40116 ( .A1(n39141), .A2(n41083), .ZN(n34666) );
  NAND2_X1 U40117 ( .A1(n41082), .A2(n8316), .ZN(n38866) );
  NAND2_X1 U40118 ( .A1(n37965), .A2(n36552), .ZN(n34663) );
  INV_X1 U40119 ( .A(n34663), .ZN(n34659) );
  NAND2_X1 U40120 ( .A1(n34659), .A2(n36542), .ZN(n34660) );
  AND2_X1 U40121 ( .A1(n41085), .A2(n38866), .ZN(n34665) );
  NAND2_X1 U40122 ( .A1(n38870), .A2(n41082), .ZN(n39709) );
  NAND3_X1 U40123 ( .A1(n34668), .A2(n41077), .A3(n34667), .ZN(n34673) );
  INV_X1 U40124 ( .A(n41084), .ZN(n38869) );
  AND2_X1 U40125 ( .A1(n41083), .A2(n39712), .ZN(n39145) );
  OAI21_X1 U40126 ( .B1(n34669), .B2(n41088), .A(n39145), .ZN(n34672) );
  NAND2_X1 U40127 ( .A1(n38869), .A2(n39713), .ZN(n38362) );
  INV_X1 U40128 ( .A(n38362), .ZN(n34670) );
  NOR2_X1 U40129 ( .A1(n41082), .A2(n41079), .ZN(n38871) );
  NAND2_X1 U40130 ( .A1(n34670), .A2(n38871), .ZN(n34671) );
  INV_X1 U40131 ( .A(n37560), .ZN(n35927) );
  NAND2_X1 U40132 ( .A1(n37561), .A2(n35927), .ZN(n34682) );
  NOR2_X1 U40133 ( .A1(n37550), .A2(n34682), .ZN(n34674) );
  NOR2_X1 U40134 ( .A1(n37544), .A2(n36272), .ZN(n34675) );
  AND2_X1 U40135 ( .A1(n37545), .A2(n37557), .ZN(n37404) );
  AOI22_X1 U40136 ( .A1(n37554), .A2(n34675), .B1(n37404), .B2(n36268), .ZN(
        n34679) );
  AND2_X1 U40137 ( .A1(n34676), .A2(n37399), .ZN(n36265) );
  NOR2_X1 U40138 ( .A1(n37557), .A2(n5784), .ZN(n34677) );
  AND2_X1 U40139 ( .A1(n35927), .A2(n36272), .ZN(n37410) );
  OAI211_X1 U40140 ( .C1(n36265), .C2(n34677), .A(n37410), .B(n37397), .ZN(
        n34678) );
  INV_X1 U40141 ( .A(n34681), .ZN(n37535) );
  NAND3_X1 U40142 ( .A1(n37554), .A2(n37535), .A3(n5784), .ZN(n37548) );
  INV_X1 U40143 ( .A(n34682), .ZN(n37558) );
  OAI21_X1 U40144 ( .B1(n37535), .B2(n37558), .A(n37539), .ZN(n34683) );
  AND2_X1 U40145 ( .A1(n36186), .A2(n37774), .ZN(n34685) );
  NOR2_X1 U40146 ( .A1(n2089), .A2(n39342), .ZN(n37779) );
  INV_X1 U40148 ( .A(n39349), .ZN(n34686) );
  OAI22_X1 U40149 ( .A1(n34686), .A2(n36189), .B1(n36191), .B2(n37775), .ZN(
        n34689) );
  AOI21_X1 U40150 ( .B1(n35943), .B2(n36200), .A(n37774), .ZN(n34688) );
  NAND2_X1 U40151 ( .A1(n36186), .A2(n36200), .ZN(n34687) );
  AND2_X1 U40152 ( .A1(n35939), .A2(n37774), .ZN(n36188) );
  NAND2_X1 U40153 ( .A1(n34691), .A2(n39348), .ZN(n34694) );
  AND2_X1 U40154 ( .A1(n34692), .A2(n36200), .ZN(n37783) );
  NAND2_X1 U40155 ( .A1(n37780), .A2(n37783), .ZN(n39345) );
  NAND2_X1 U40156 ( .A1(n39345), .A2(n37782), .ZN(n34693) );
  NAND3_X1 U40157 ( .A1(n34694), .A2(n34693), .A3(n36197), .ZN(n34695) );
  NAND2_X1 U40158 ( .A1(n41985), .A2(n41647), .ZN(n41098) );
  OAI21_X1 U40159 ( .B1(n38979), .B2(n34700), .A(n2177), .ZN(n34708) );
  OAI22_X1 U40160 ( .A1(n39473), .A2(n34701), .B1(n37809), .B2(n39472), .ZN(
        n34702) );
  NOR2_X1 U40161 ( .A1(n39485), .A2(n34702), .ZN(n34707) );
  NOR2_X1 U40162 ( .A1(n39479), .A2(n1075), .ZN(n34703) );
  OAI211_X1 U40163 ( .C1(n39484), .C2(n34703), .A(n39481), .B(n39478), .ZN(
        n36208) );
  INV_X1 U40164 ( .A(n37800), .ZN(n34705) );
  NOR2_X1 U40165 ( .A1(n2177), .A2(n39472), .ZN(n34704) );
  OAI21_X1 U40166 ( .B1(n34705), .B2(n34704), .A(n39471), .ZN(n34706) );
  INV_X1 U40168 ( .A(n41650), .ZN(n41096) );
  NOR2_X1 U40169 ( .A1(n41098), .A2(n6938), .ZN(n40622) );
  XNOR2_X1 U40170 ( .A(n36856), .B(n704), .ZN(n34718) );
  XNOR2_X1 U40171 ( .A(n34710), .B(n34709), .ZN(n34712) );
  XNOR2_X1 U40172 ( .A(n34712), .B(n34711), .ZN(n34714) );
  XNOR2_X1 U40173 ( .A(n34714), .B(n34713), .ZN(n34715) );
  XNOR2_X1 U40174 ( .A(n35588), .B(n34715), .ZN(n34716) );
  XNOR2_X1 U40175 ( .A(n34716), .B(n36939), .ZN(n34717) );
  XNOR2_X1 U40176 ( .A(n34718), .B(n34717), .ZN(n34723) );
  XNOR2_X1 U40177 ( .A(n35587), .B(n34721), .ZN(n34722) );
  XNOR2_X1 U40178 ( .A(n34722), .B(n34723), .ZN(n34725) );
  INV_X1 U40179 ( .A(n34724), .ZN(n35369) );
  XNOR2_X1 U40180 ( .A(n34729), .B(n34728), .ZN(n34730) );
  XNOR2_X1 U40181 ( .A(n34731), .B(n34730), .ZN(n34732) );
  XNOR2_X1 U40182 ( .A(n37062), .B(n34732), .ZN(n34733) );
  XNOR2_X1 U40183 ( .A(n33759), .B(n34733), .ZN(n34734) );
  XNOR2_X1 U40184 ( .A(n34734), .B(n51472), .ZN(n34735) );
  XNOR2_X1 U40187 ( .A(n35086), .B(n35536), .ZN(n34741) );
  XNOR2_X1 U40188 ( .A(n34741), .B(n35537), .ZN(n35803) );
  XNOR2_X1 U40189 ( .A(n35095), .B(n34842), .ZN(n34748) );
  XNOR2_X1 U40190 ( .A(n34743), .B(n34742), .ZN(n34745) );
  XNOR2_X1 U40191 ( .A(n34745), .B(n34744), .ZN(n34746) );
  XNOR2_X1 U40192 ( .A(n2129), .B(n34746), .ZN(n34747) );
  XNOR2_X1 U40193 ( .A(n34748), .B(n34747), .ZN(n34749) );
  XNOR2_X1 U40194 ( .A(n35803), .B(n34749), .ZN(n34752) );
  XNOR2_X1 U40195 ( .A(n35345), .B(n36701), .ZN(n34750) );
  XNOR2_X1 U40196 ( .A(n34750), .B(n35633), .ZN(n34751) );
  XNOR2_X1 U40197 ( .A(n34751), .B(n51449), .ZN(n36787) );
  XNOR2_X1 U40198 ( .A(n34752), .B(n36787), .ZN(n34758) );
  XNOR2_X1 U40199 ( .A(n34754), .B(n34753), .ZN(n34756) );
  XNOR2_X1 U40200 ( .A(n34756), .B(n34755), .ZN(n34757) );
  INV_X1 U40201 ( .A(n39438), .ZN(n37720) );
  XNOR2_X1 U40202 ( .A(n35075), .B(n34760), .ZN(n34767) );
  XNOR2_X1 U40203 ( .A(n34761), .B(n35067), .ZN(n34764) );
  INV_X1 U40204 ( .A(n34762), .ZN(n34763) );
  XNOR2_X1 U40205 ( .A(n34764), .B(n34763), .ZN(n34765) );
  XNOR2_X1 U40206 ( .A(n36805), .B(n34765), .ZN(n34766) );
  XNOR2_X1 U40207 ( .A(n34767), .B(n34766), .ZN(n34768) );
  AND2_X1 U40208 ( .A1(n39028), .A2(n39438), .ZN(n39034) );
  NAND2_X1 U40209 ( .A1(n39034), .A2(n34800), .ZN(n36896) );
  XNOR2_X1 U40210 ( .A(n34774), .B(n34773), .ZN(n34775) );
  XNOR2_X1 U40211 ( .A(n34776), .B(n34775), .ZN(n34777) );
  XNOR2_X1 U40212 ( .A(n36829), .B(n34777), .ZN(n34778) );
  XNOR2_X1 U40213 ( .A(n35656), .B(n34778), .ZN(n34781) );
  INV_X1 U40214 ( .A(n37008), .ZN(n34779) );
  XNOR2_X1 U40215 ( .A(n34875), .B(n34781), .ZN(n34783) );
  XNOR2_X1 U40216 ( .A(n34783), .B(n34782), .ZN(n34784) );
  XNOR2_X1 U40217 ( .A(n34784), .B(n36751), .ZN(n34785) );
  XNOR2_X1 U40218 ( .A(n35482), .B(n36999), .ZN(n34787) );
  XNOR2_X1 U40219 ( .A(n34888), .B(n34787), .ZN(n34788) );
  XNOR2_X1 U40220 ( .A(n34789), .B(n34891), .ZN(n34792) );
  INV_X1 U40221 ( .A(n34790), .ZN(n34791) );
  XNOR2_X1 U40222 ( .A(n34792), .B(n34791), .ZN(n34793) );
  XNOR2_X1 U40223 ( .A(n35683), .B(n34793), .ZN(n34794) );
  XNOR2_X1 U40224 ( .A(n35133), .B(n34794), .ZN(n34795) );
  XNOR2_X1 U40225 ( .A(n37001), .B(n34795), .ZN(n34796) );
  NAND2_X1 U40226 ( .A1(n37716), .A2(n39437), .ZN(n34805) );
  AND2_X1 U40227 ( .A1(n39035), .A2(n36901), .ZN(n36260) );
  NAND2_X1 U40228 ( .A1(n467), .A2(n37720), .ZN(n36912) );
  AOI21_X1 U40229 ( .B1(n36260), .B2(n36259), .A(n36912), .ZN(n34799) );
  NAND2_X1 U40230 ( .A1(n39453), .A2(n51737), .ZN(n34798) );
  NAND2_X1 U40231 ( .A1(n34806), .A2(n39438), .ZN(n36895) );
  INV_X1 U40232 ( .A(n36895), .ZN(n36907) );
  OAI21_X1 U40233 ( .B1(n36907), .B2(n36901), .A(n39453), .ZN(n34797) );
  INV_X1 U40234 ( .A(n39034), .ZN(n39462) );
  NOR2_X1 U40235 ( .A1(n39462), .A2(n51737), .ZN(n39443) );
  INV_X1 U40236 ( .A(n39448), .ZN(n39463) );
  NAND3_X1 U40237 ( .A1(n39443), .A2(n39463), .A3(n39035), .ZN(n34803) );
  NOR2_X1 U40238 ( .A1(n37722), .A2(n51737), .ZN(n34801) );
  AND2_X1 U40239 ( .A1(n34806), .A2(n37720), .ZN(n36903) );
  AOI22_X1 U40240 ( .A1(n34801), .A2(n39441), .B1(n39442), .B2(n36903), .ZN(
        n34802) );
  AOI21_X1 U40241 ( .B1(n39448), .B2(n39032), .A(n39452), .ZN(n37719) );
  NAND2_X1 U40242 ( .A1(n34806), .A2(n39464), .ZN(n34807) );
  MUX2_X1 U40243 ( .A(n37719), .B(n36254), .S(n39438), .Z(n34808) );
  INV_X2 U40244 ( .A(n41645), .ZN(n41977) );
  XNOR2_X1 U40245 ( .A(n34811), .B(n45736), .ZN(n34813) );
  XNOR2_X1 U40246 ( .A(n34813), .B(n51413), .ZN(n34814) );
  XNOR2_X1 U40247 ( .A(n35254), .B(n37045), .ZN(n34815) );
  XNOR2_X1 U40249 ( .A(n44495), .B(n34816), .ZN(n34817) );
  XNOR2_X1 U40250 ( .A(n34818), .B(n34817), .ZN(n34819) );
  XNOR2_X1 U40251 ( .A(n37261), .B(n34819), .ZN(n34820) );
  XNOR2_X1 U40252 ( .A(n34820), .B(n36681), .ZN(n34821) );
  XNOR2_X1 U40254 ( .A(n34823), .B(n34824), .ZN(n35371) );
  INV_X1 U40255 ( .A(n35371), .ZN(n34825) );
  XNOR2_X1 U40256 ( .A(n34826), .B(n34825), .ZN(n34827) );
  INV_X1 U40257 ( .A(n34830), .ZN(n34832) );
  XNOR2_X1 U40258 ( .A(n42549), .B(n43586), .ZN(n34831) );
  XNOR2_X1 U40259 ( .A(n34832), .B(n34831), .ZN(n34833) );
  XNOR2_X1 U40260 ( .A(n37241), .B(n34833), .ZN(n34834) );
  XNOR2_X1 U40261 ( .A(n33195), .B(n34834), .ZN(n34837) );
  XNOR2_X1 U40262 ( .A(n34835), .B(n35609), .ZN(n34836) );
  XNOR2_X1 U40263 ( .A(n34837), .B(n34836), .ZN(n34838) );
  XNOR2_X1 U40264 ( .A(n34839), .B(n35350), .ZN(n34840) );
  XNOR2_X1 U40265 ( .A(n34841), .B(n4558), .ZN(n34843) );
  XNOR2_X1 U40266 ( .A(n34843), .B(n8135), .ZN(n36709) );
  XNOR2_X1 U40267 ( .A(n35095), .B(n2129), .ZN(n34846) );
  XNOR2_X1 U40268 ( .A(n35537), .B(n37292), .ZN(n34845) );
  XNOR2_X1 U40269 ( .A(n34846), .B(n34845), .ZN(n34847) );
  XNOR2_X1 U40270 ( .A(n36709), .B(n34847), .ZN(n34849) );
  INV_X1 U40271 ( .A(n34850), .ZN(n34853) );
  XNOR2_X1 U40272 ( .A(n34851), .B(n43702), .ZN(n34852) );
  XNOR2_X1 U40273 ( .A(n34853), .B(n34852), .ZN(n34854) );
  XNOR2_X1 U40274 ( .A(n37081), .B(n34854), .ZN(n34855) );
  XNOR2_X1 U40275 ( .A(n34857), .B(n34856), .ZN(n34859) );
  XNOR2_X1 U40276 ( .A(n34859), .B(n34858), .ZN(n34860) );
  XNOR2_X1 U40277 ( .A(n35240), .B(n4653), .ZN(n34861) );
  XNOR2_X1 U40278 ( .A(n37095), .B(n34861), .ZN(n36963) );
  INV_X1 U40279 ( .A(n36963), .ZN(n34864) );
  INV_X1 U40280 ( .A(n34865), .ZN(n34867) );
  XNOR2_X1 U40281 ( .A(n34867), .B(n34866), .ZN(n34868) );
  XNOR2_X1 U40282 ( .A(n34869), .B(n34868), .ZN(n34870) );
  XNOR2_X1 U40283 ( .A(n36807), .B(n34870), .ZN(n34871) );
  XNOR2_X1 U40284 ( .A(n37111), .B(n34871), .ZN(n34872) );
  INV_X1 U40285 ( .A(n34875), .ZN(n34876) );
  XNOR2_X1 U40286 ( .A(n35476), .B(n34877), .ZN(n34886) );
  XNOR2_X1 U40287 ( .A(n34878), .B(n36739), .ZN(n34879) );
  XNOR2_X1 U40288 ( .A(n34879), .B(n44555), .ZN(n34880) );
  XNOR2_X1 U40289 ( .A(n34881), .B(n34880), .ZN(n34882) );
  XNOR2_X1 U40290 ( .A(n35747), .B(n34882), .ZN(n34884) );
  XNOR2_X1 U40291 ( .A(n34884), .B(n34883), .ZN(n34885) );
  XNOR2_X1 U40292 ( .A(n34886), .B(n34885), .ZN(n34887) );
  XNOR2_X1 U40293 ( .A(n35120), .B(n36748), .ZN(n37151) );
  XNOR2_X1 U40294 ( .A(n35761), .B(n34888), .ZN(n37120) );
  XNOR2_X1 U40295 ( .A(n37120), .B(n34889), .ZN(n37003) );
  XNOR2_X1 U40296 ( .A(n35680), .B(n460), .ZN(n34890) );
  XNOR2_X1 U40297 ( .A(n37003), .B(n34890), .ZN(n34902) );
  XNOR2_X1 U40298 ( .A(n34892), .B(n34891), .ZN(n34894) );
  XNOR2_X1 U40299 ( .A(n34894), .B(n34893), .ZN(n34895) );
  XNOR2_X1 U40300 ( .A(n34896), .B(n34895), .ZN(n34897) );
  XNOR2_X1 U40301 ( .A(n37001), .B(n34897), .ZN(n34899) );
  XNOR2_X1 U40302 ( .A(n34899), .B(n34898), .ZN(n34900) );
  XNOR2_X1 U40303 ( .A(n37130), .B(n34900), .ZN(n34901) );
  XNOR2_X2 U40304 ( .A(n34901), .B(n34902), .ZN(n39395) );
  AND3_X1 U40305 ( .A1(n3577), .A2(n39003), .A3(n39395), .ZN(n34903) );
  INV_X1 U40306 ( .A(n34905), .ZN(n39400) );
  INV_X1 U40308 ( .A(n39397), .ZN(n39402) );
  NAND2_X1 U40309 ( .A1(n34906), .A2(n38998), .ZN(n37894) );
  INV_X1 U40310 ( .A(n39395), .ZN(n38999) );
  OAI211_X1 U40311 ( .C1(n38999), .C2(n3735), .A(n34909), .B(n39399), .ZN(
        n34910) );
  NAND2_X1 U40312 ( .A1(n41642), .A2(n41646), .ZN(n34917) );
  NAND2_X1 U40313 ( .A1(n41977), .A2(n34917), .ZN(n34919) );
  AOI22_X1 U40314 ( .A1(n37762), .A2(n36248), .B1(n37510), .B2(n35923), .ZN(
        n34916) );
  NAND3_X1 U40315 ( .A1(n36248), .A2(n37499), .A3(n36251), .ZN(n34912) );
  INV_X1 U40316 ( .A(n37502), .ZN(n34913) );
  NAND4_X1 U40317 ( .A1(n36240), .A2(n37749), .A3(n34913), .A4(n37757), .ZN(
        n34915) );
  XNOR2_X1 U40318 ( .A(n40617), .B(n41647), .ZN(n34918) );
  AND2_X1 U40319 ( .A1(n41104), .A2(n34917), .ZN(n41101) );
  INV_X1 U40320 ( .A(n41975), .ZN(n41103) );
  OAI21_X1 U40321 ( .B1(n41650), .B2(n41646), .A(n6940), .ZN(n34920) );
  INV_X1 U40322 ( .A(n41647), .ZN(n40608) );
  NAND2_X1 U40323 ( .A1(n41650), .A2(n41646), .ZN(n40615) );
  INV_X1 U40324 ( .A(n36426), .ZN(n34921) );
  NOR2_X1 U40325 ( .A1(n36062), .A2(n34921), .ZN(n34922) );
  INV_X1 U40326 ( .A(n34924), .ZN(n34926) );
  NAND2_X1 U40327 ( .A1(n51717), .A2(n36427), .ZN(n34925) );
  INV_X1 U40328 ( .A(n34930), .ZN(n34933) );
  NAND2_X1 U40329 ( .A1(n36420), .A2(n36427), .ZN(n34932) );
  NAND4_X1 U40330 ( .A1(n34933), .A2(n34932), .A3(n34931), .A4(n36057), .ZN(
        n34934) );
  NOR2_X1 U40331 ( .A1(n36065), .A2(n36420), .ZN(n36603) );
  NOR2_X1 U40332 ( .A1(n36609), .A2(n36604), .ZN(n34935) );
  OAI21_X1 U40333 ( .B1(n36603), .B2(n34935), .A(n36426), .ZN(n34936) );
  OAI211_X1 U40334 ( .C1(n36376), .C2(n34938), .A(n36375), .B(n34937), .ZN(
        n34942) );
  NAND3_X1 U40336 ( .A1(n38031), .A2(n36381), .A3(n35159), .ZN(n34940) );
  AND3_X1 U40337 ( .A1(n34941), .A2(n34942), .A3(n34940), .ZN(n34957) );
  OAI21_X1 U40338 ( .B1(n38043), .B2(n38037), .A(n38038), .ZN(n34943) );
  NOR2_X1 U40340 ( .A1(n38030), .A2(n38040), .ZN(n36382) );
  AOI22_X1 U40341 ( .A1(n34944), .A2(n34943), .B1(n36382), .B2(n38037), .ZN(
        n34956) );
  NOR2_X1 U40342 ( .A1(n38031), .A2(n35157), .ZN(n38044) );
  NAND2_X1 U40343 ( .A1(n38034), .A2(n34945), .ZN(n35160) );
  NOR2_X1 U40344 ( .A1(n36376), .A2(n35160), .ZN(n34946) );
  AOI22_X1 U40345 ( .A1(n38044), .A2(n34947), .B1(n36371), .B2(n34946), .ZN(
        n34955) );
  NAND2_X1 U40346 ( .A1(n34948), .A2(n38043), .ZN(n34952) );
  INV_X1 U40347 ( .A(n38036), .ZN(n34951) );
  OAI211_X1 U40348 ( .C1(n34952), .C2(n34951), .A(n34950), .B(n34949), .ZN(
        n34953) );
  INV_X1 U40349 ( .A(n34953), .ZN(n34954) );
  NOR2_X1 U40350 ( .A1(n41049), .A2(n6392), .ZN(n38389) );
  NAND2_X1 U40352 ( .A1(n34959), .A2(n38082), .ZN(n34968) );
  INV_X1 U40353 ( .A(n36317), .ZN(n34961) );
  OAI21_X1 U40354 ( .B1(n36640), .B2(n34961), .A(n36641), .ZN(n34962) );
  NAND2_X1 U40355 ( .A1(n34962), .A2(n36629), .ZN(n34967) );
  NAND3_X1 U40356 ( .A1(n36639), .A2(n38073), .A3(n34963), .ZN(n34966) );
  OAI21_X1 U40357 ( .B1(n36635), .B2(n36312), .A(n38094), .ZN(n34964) );
  NAND2_X1 U40358 ( .A1(n34964), .A2(n36632), .ZN(n34965) );
  OR2_X1 U40360 ( .A1(n38389), .A2(n41057), .ZN(n38391) );
  NOR2_X1 U40361 ( .A1(n37997), .A2(n35028), .ZN(n36358) );
  OAI21_X1 U40362 ( .B1(n36358), .B2(n34969), .A(n38177), .ZN(n34979) );
  INV_X1 U40363 ( .A(n37997), .ZN(n35027) );
  NAND2_X1 U40366 ( .A1(n38015), .A2(n36364), .ZN(n34973) );
  AOI21_X1 U40367 ( .B1(n34971), .B2(n38002), .A(n38018), .ZN(n34972) );
  AOI21_X1 U40368 ( .B1(n34973), .B2(n34972), .A(n38019), .ZN(n34974) );
  NAND2_X1 U40370 ( .A1(n34984), .A2(n36518), .ZN(n36516) );
  INV_X1 U40371 ( .A(n36516), .ZN(n36525) );
  INV_X1 U40372 ( .A(n37975), .ZN(n36530) );
  NAND3_X1 U40373 ( .A1(n36525), .A2(n37980), .A3(n36530), .ZN(n34983) );
  NAND3_X1 U40374 ( .A1(n37991), .A2(n36351), .A3(n36522), .ZN(n34981) );
  NAND3_X1 U40375 ( .A1(n37991), .A2(n594), .A3(n37975), .ZN(n34980) );
  OAI22_X1 U40376 ( .A1(n34985), .A2(n37974), .B1(n34984), .B2(n36080), .ZN(
        n34986) );
  NAND2_X1 U40377 ( .A1(n34987), .A2(n37976), .ZN(n36524) );
  INV_X1 U40380 ( .A(n36077), .ZN(n36353) );
  OAI21_X1 U40381 ( .B1(n36516), .B2(n37980), .A(n36353), .ZN(n34989) );
  NAND2_X1 U40382 ( .A1(n34989), .A2(n36351), .ZN(n36348) );
  NAND2_X1 U40383 ( .A1(n40512), .A2(n41063), .ZN(n39601) );
  AND2_X1 U40384 ( .A1(n34993), .A2(n37957), .ZN(n35002) );
  OAI21_X1 U40385 ( .B1(n51909), .B2(n36027), .A(n36542), .ZN(n35001) );
  NAND2_X1 U40386 ( .A1(n37965), .A2(n36547), .ZN(n34992) );
  INV_X1 U40387 ( .A(n36552), .ZN(n34994) );
  NAND2_X1 U40388 ( .A1(n34994), .A2(n8016), .ZN(n34996) );
  NAND2_X1 U40389 ( .A1(n34997), .A2(n51077), .ZN(n34998) );
  NAND2_X1 U40390 ( .A1(n6392), .A2(n40502), .ZN(n41047) );
  NAND2_X1 U40391 ( .A1(n41047), .A2(n41057), .ZN(n35003) );
  OR2_X1 U40393 ( .A1(n40513), .A2(n41047), .ZN(n40508) );
  NAND3_X1 U40394 ( .A1(n39131), .A2(n41065), .A3(n41057), .ZN(n35005) );
  XNOR2_X1 U40395 ( .A(n41065), .B(n41063), .ZN(n35006) );
  OAI211_X1 U40396 ( .C1(n41066), .C2(n35006), .A(n39129), .B(n41064), .ZN(
        n35007) );
  NOR2_X1 U40397 ( .A1(n38053), .A2(n36338), .ZN(n36344) );
  INV_X1 U40398 ( .A(n36336), .ZN(n38065) );
  AND2_X1 U40399 ( .A1(n38054), .A2(n38146), .ZN(n35011) );
  AOI22_X1 U40400 ( .A1(n36344), .A2(n38065), .B1(n35011), .B2(n38058), .ZN(
        n35022) );
  XNOR2_X1 U40401 ( .A(n38055), .B(n36338), .ZN(n35012) );
  NAND2_X1 U40402 ( .A1(n5443), .A2(n36340), .ZN(n38063) );
  INV_X1 U40403 ( .A(n38063), .ZN(n36330) );
  AND2_X1 U40404 ( .A1(n36340), .A2(n36337), .ZN(n38147) );
  NAND4_X1 U40405 ( .A1(n36167), .A2(n38050), .A3(n38147), .A4(n38145), .ZN(
        n35013) );
  AND2_X1 U40406 ( .A1(n35014), .A2(n35013), .ZN(n35021) );
  INV_X1 U40407 ( .A(n36167), .ZN(n35015) );
  NAND3_X1 U40408 ( .A1(n36325), .A2(n36338), .A3(n36336), .ZN(n35016) );
  AND2_X1 U40409 ( .A1(n38052), .A2(n35016), .ZN(n35020) );
  NAND2_X1 U40410 ( .A1(n51522), .A2(n38142), .ZN(n36335) );
  OAI21_X1 U40411 ( .B1(n38055), .B2(n38145), .A(n36335), .ZN(n35018) );
  OAI211_X1 U40412 ( .C1(n36342), .C2(n38136), .A(n38144), .B(n35018), .ZN(
        n35019) );
  INV_X1 U40413 ( .A(n38001), .ZN(n38016) );
  OAI211_X1 U40414 ( .C1(n36359), .C2(n38016), .A(n37997), .B(n35023), .ZN(
        n35024) );
  INV_X1 U40415 ( .A(n38173), .ZN(n35025) );
  OAI211_X1 U40416 ( .C1(n38005), .C2(n35028), .A(n38001), .B(n38006), .ZN(
        n35029) );
  XNOR2_X1 U40417 ( .A(n35032), .B(n35031), .ZN(n35044) );
  XNOR2_X1 U40418 ( .A(n35586), .B(n35033), .ZN(n35042) );
  XNOR2_X1 U40419 ( .A(n37262), .B(n35034), .ZN(n37047) );
  XNOR2_X1 U40420 ( .A(n35036), .B(n35035), .ZN(n35037) );
  XNOR2_X1 U40421 ( .A(n35038), .B(n35037), .ZN(n35039) );
  XNOR2_X1 U40422 ( .A(n35833), .B(n35039), .ZN(n35040) );
  XNOR2_X1 U40423 ( .A(n37047), .B(n35040), .ZN(n35041) );
  XNOR2_X1 U40424 ( .A(n35042), .B(n35041), .ZN(n35043) );
  INV_X1 U40425 ( .A(n35045), .ZN(n35046) );
  XNOR2_X1 U40426 ( .A(n35046), .B(n35350), .ZN(n35064) );
  XNOR2_X1 U40427 ( .A(n35047), .B(n35048), .ZN(n35051) );
  INV_X1 U40428 ( .A(n35049), .ZN(n35050) );
  XNOR2_X1 U40429 ( .A(n35051), .B(n35050), .ZN(n35614) );
  XNOR2_X1 U40430 ( .A(n36932), .B(n35052), .ZN(n35054) );
  XNOR2_X1 U40431 ( .A(n35054), .B(n33759), .ZN(n37236) );
  INV_X1 U40432 ( .A(n35055), .ZN(n35057) );
  XNOR2_X1 U40433 ( .A(n35057), .B(n35056), .ZN(n35058) );
  XNOR2_X1 U40434 ( .A(n35059), .B(n35058), .ZN(n35060) );
  XNOR2_X1 U40435 ( .A(n37063), .B(n35060), .ZN(n35061) );
  XNOR2_X1 U40436 ( .A(n35061), .B(n37236), .ZN(n35062) );
  XNOR2_X1 U40437 ( .A(n35062), .B(n35614), .ZN(n35063) );
  XNOR2_X1 U40438 ( .A(n35326), .B(n35066), .ZN(n35074) );
  XNOR2_X1 U40439 ( .A(n35068), .B(n35067), .ZN(n35069) );
  XNOR2_X1 U40440 ( .A(n35325), .B(n35069), .ZN(n35071) );
  XNOR2_X1 U40441 ( .A(n35070), .B(n4890), .ZN(n37094) );
  XNOR2_X1 U40442 ( .A(n35071), .B(n37094), .ZN(n35072) );
  XNOR2_X1 U40443 ( .A(n35074), .B(n35073), .ZN(n35079) );
  XNOR2_X1 U40444 ( .A(n35075), .B(n37108), .ZN(n37270) );
  XNOR2_X1 U40445 ( .A(n37270), .B(n35333), .ZN(n35076) );
  XNOR2_X1 U40446 ( .A(n35077), .B(n35076), .ZN(n35630) );
  XNOR2_X1 U40447 ( .A(n35544), .B(n35080), .ZN(n35084) );
  XNOR2_X1 U40448 ( .A(n35081), .B(n37082), .ZN(n35082) );
  XNOR2_X1 U40449 ( .A(n35345), .B(n35082), .ZN(n35083) );
  XNOR2_X1 U40450 ( .A(n35084), .B(n35083), .ZN(n35087) );
  XNOR2_X1 U40451 ( .A(n35087), .B(n37284), .ZN(n35092) );
  XNOR2_X1 U40452 ( .A(n35800), .B(n35088), .ZN(n35089) );
  XNOR2_X1 U40453 ( .A(n35089), .B(n36792), .ZN(n37078) );
  XNOR2_X1 U40454 ( .A(n35090), .B(n37078), .ZN(n35091) );
  XNOR2_X1 U40455 ( .A(n35091), .B(n35092), .ZN(n35101) );
  INV_X1 U40456 ( .A(n35093), .ZN(n35094) );
  XNOR2_X1 U40457 ( .A(n35095), .B(n35094), .ZN(n35226) );
  INV_X1 U40458 ( .A(n35226), .ZN(n35098) );
  INV_X1 U40459 ( .A(n35096), .ZN(n35097) );
  XNOR2_X1 U40460 ( .A(n35098), .B(n35097), .ZN(n35099) );
  XNOR2_X1 U40461 ( .A(n37091), .B(n35099), .ZN(n35100) );
  XNOR2_X1 U40462 ( .A(n35101), .B(n35100), .ZN(n38483) );
  INV_X1 U40463 ( .A(n38483), .ZN(n38480) );
  NAND2_X1 U40464 ( .A1(n35102), .A2(n38480), .ZN(n38473) );
  INV_X1 U40465 ( .A(n38468), .ZN(n37417) );
  NAND2_X1 U40466 ( .A1(n37414), .A2(n38471), .ZN(n38111) );
  NAND2_X1 U40467 ( .A1(n37415), .A2(n38111), .ZN(n37422) );
  OAI211_X1 U40468 ( .C1(n38119), .C2(n38473), .A(n38118), .B(n37422), .ZN(
        n35139) );
  XNOR2_X1 U40469 ( .A(n35106), .B(n35105), .ZN(n35117) );
  XNOR2_X1 U40470 ( .A(n35107), .B(n4739), .ZN(n35109) );
  XNOR2_X1 U40471 ( .A(n35109), .B(n35108), .ZN(n35111) );
  XNOR2_X1 U40472 ( .A(n35111), .B(n35110), .ZN(n35112) );
  XNOR2_X1 U40473 ( .A(n35113), .B(n35112), .ZN(n35114) );
  XNOR2_X1 U40474 ( .A(n35115), .B(n35114), .ZN(n35116) );
  XNOR2_X1 U40475 ( .A(n35117), .B(n35116), .ZN(n35118) );
  INV_X1 U40476 ( .A(n35464), .ZN(n35121) );
  XNOR2_X1 U40477 ( .A(n35121), .B(n518), .ZN(n35122) );
  XNOR2_X1 U40479 ( .A(n35482), .B(n35124), .ZN(n35125) );
  INV_X1 U40480 ( .A(n35488), .ZN(n35667) );
  XNOR2_X1 U40481 ( .A(n35667), .B(n35125), .ZN(n35127) );
  XNOR2_X1 U40482 ( .A(n35127), .B(n35126), .ZN(n35129) );
  XNOR2_X1 U40483 ( .A(n35129), .B(n35128), .ZN(n35138) );
  XNOR2_X1 U40484 ( .A(n44921), .B(n35130), .ZN(n35131) );
  XNOR2_X1 U40485 ( .A(n35683), .B(n35131), .ZN(n35132) );
  XNOR2_X1 U40486 ( .A(n35133), .B(n35132), .ZN(n35134) );
  XNOR2_X1 U40487 ( .A(n35134), .B(n35669), .ZN(n35135) );
  XNOR2_X1 U40488 ( .A(n35136), .B(n35135), .ZN(n35137) );
  NOR2_X1 U40491 ( .A1(n8509), .A2(n38471), .ZN(n35140) );
  AOI22_X1 U40492 ( .A1(n35141), .A2(n38485), .B1(n38481), .B2(n35140), .ZN(
        n35145) );
  AND2_X1 U40493 ( .A1(n38481), .A2(n6637), .ZN(n38122) );
  NAND2_X1 U40494 ( .A1(n38122), .A2(n37414), .ZN(n35142) );
  MUX2_X1 U40495 ( .A(n38484), .B(n35142), .S(n38473), .Z(n35143) );
  AND2_X1 U40496 ( .A1(n33062), .A2(n38201), .ZN(n38573) );
  AND2_X1 U40497 ( .A1(n38196), .A2(n38201), .ZN(n35146) );
  NAND2_X1 U40498 ( .A1(n38570), .A2(n38576), .ZN(n35147) );
  INV_X1 U40499 ( .A(n38204), .ZN(n35150) );
  NAND3_X1 U40500 ( .A1(n36106), .A2(n1764), .A3(n38204), .ZN(n35148) );
  INV_X1 U40501 ( .A(n35706), .ZN(n38560) );
  NAND3_X1 U40502 ( .A1(n38567), .A2(n38560), .A3(n38565), .ZN(n35702) );
  OAI21_X1 U40503 ( .B1(n36103), .B2(n35706), .A(n35702), .ZN(n35149) );
  INV_X1 U40504 ( .A(n35149), .ZN(n35152) );
  NOR2_X1 U40505 ( .A1(n36383), .A2(n614), .ZN(n35153) );
  AOI22_X1 U40506 ( .A1(n35153), .A2(n35159), .B1(n38036), .B2(n38037), .ZN(
        n35167) );
  INV_X1 U40507 ( .A(n36372), .ZN(n35154) );
  OAI21_X1 U40508 ( .B1(n35156), .B2(n35155), .A(n38027), .ZN(n35158) );
  AOI22_X1 U40509 ( .A1(n36384), .A2(n35158), .B1(n36380), .B2(n35157), .ZN(
        n35166) );
  INV_X1 U40510 ( .A(n35159), .ZN(n35161) );
  NOR2_X1 U40511 ( .A1(n35161), .A2(n35160), .ZN(n38042) );
  INV_X1 U40512 ( .A(n36376), .ZN(n38039) );
  OAI21_X1 U40513 ( .B1(n35162), .B2(n35161), .A(n38039), .ZN(n35163) );
  INV_X1 U40514 ( .A(n38031), .ZN(n36377) );
  OAI21_X1 U40515 ( .B1(n38042), .B2(n35163), .A(n36377), .ZN(n35165) );
  NAND3_X1 U40516 ( .A1(n38042), .A2(n36375), .A3(n38039), .ZN(n35164) );
  NAND2_X1 U40517 ( .A1(n40417), .A2(n41275), .ZN(n35168) );
  OAI22_X1 U40518 ( .A1(n35168), .A2(n52192), .B1(n40417), .B2(n41275), .ZN(
        n35184) );
  INV_X1 U40519 ( .A(n35169), .ZN(n38551) );
  INV_X1 U40521 ( .A(n35170), .ZN(n35180) );
  NOR2_X1 U40523 ( .A1(n38553), .A2(n38550), .ZN(n35174) );
  NOR2_X1 U40524 ( .A1(n38552), .A2(n38558), .ZN(n35172) );
  NOR2_X1 U40525 ( .A1(n38226), .A2(n35175), .ZN(n35176) );
  AOI21_X1 U40526 ( .B1(n35177), .B2(n38214), .A(n35176), .ZN(n35182) );
  NOR2_X1 U40527 ( .A1(n35179), .A2(n36141), .ZN(n36307) );
  NAND2_X1 U40528 ( .A1(n35180), .A2(n36307), .ZN(n35181) );
  AOI22_X1 U40529 ( .A1(n35185), .A2(n397), .B1(n35184), .B2(n39115), .ZN(
        n35193) );
  OR2_X1 U40530 ( .A1(n41029), .A2(n41276), .ZN(n40410) );
  NAND2_X1 U40531 ( .A1(n41293), .A2(n41292), .ZN(n41282) );
  NAND2_X1 U40532 ( .A1(n52192), .A2(n41276), .ZN(n40418) );
  OAI211_X1 U40533 ( .C1(n397), .C2(n40410), .A(n41282), .B(n40418), .ZN(
        n35186) );
  NAND2_X1 U40534 ( .A1(n35186), .A2(n41286), .ZN(n35192) );
  AND2_X1 U40535 ( .A1(n41029), .A2(n41039), .ZN(n41033) );
  AOI21_X1 U40536 ( .B1(n41039), .B2(n52192), .A(n41276), .ZN(n35187) );
  NOR2_X1 U40537 ( .A1(n41033), .A2(n35187), .ZN(n35189) );
  OR2_X1 U40538 ( .A1(n41039), .A2(n41292), .ZN(n35188) );
  NAND4_X1 U40539 ( .A1(n35189), .A2(n41274), .A3(n40422), .A4(n35188), .ZN(
        n35191) );
  INV_X1 U40540 ( .A(n41282), .ZN(n39121) );
  OAI21_X1 U40541 ( .B1(n41033), .B2(n41276), .A(n39121), .ZN(n35190) );
  NAND4_X2 U40542 ( .A1(n35193), .A2(n35192), .A3(n35191), .A4(n35190), .ZN(
        n43623) );
  XNOR2_X1 U40543 ( .A(n45279), .B(n45415), .ZN(n44318) );
  XNOR2_X1 U40544 ( .A(n44318), .B(n42353), .ZN(n42734) );
  NAND2_X1 U40545 ( .A1(n37645), .A2(n35728), .ZN(n35201) );
  NAND3_X1 U40546 ( .A1(n35736), .A2(n37637), .A3(n37649), .ZN(n35195) );
  NAND2_X1 U40547 ( .A1(n35195), .A2(n35194), .ZN(n35197) );
  NAND3_X1 U40548 ( .A1(n36000), .A2(n34632), .A3(n37646), .ZN(n35196) );
  NAND2_X1 U40549 ( .A1(n35197), .A2(n35196), .ZN(n35200) );
  NAND2_X1 U40550 ( .A1(n36414), .A2(n36410), .ZN(n36403) );
  NAND3_X1 U40551 ( .A1(n35201), .A2(n35200), .A3(n35199), .ZN(n35202) );
  OR2_X1 U40552 ( .A1(n35880), .A2(n36047), .ZN(n36056) );
  INV_X1 U40553 ( .A(n35880), .ZN(n35871) );
  NAND3_X1 U40554 ( .A1(n35871), .A2(n36462), .A3(n36595), .ZN(n35206) );
  OAI211_X1 U40555 ( .C1(n36052), .C2(n3927), .A(n36454), .B(n35879), .ZN(
        n35208) );
  OAI21_X1 U40556 ( .B1(n35214), .B2(n35209), .A(n35208), .ZN(n35211) );
  NOR2_X1 U40557 ( .A1(n36592), .A2(n36458), .ZN(n35210) );
  NOR2_X1 U40558 ( .A1(n36462), .A2(n36595), .ZN(n35213) );
  AOI22_X1 U40559 ( .A1(n35213), .A2(n36046), .B1(n35212), .B2(n35881), .ZN(
        n35219) );
  NOR2_X1 U40560 ( .A1(n35214), .A2(n36589), .ZN(n35216) );
  OAI21_X1 U40561 ( .B1(n35217), .B2(n35216), .A(n36591), .ZN(n35218) );
  INV_X1 U40562 ( .A(n35220), .ZN(n35222) );
  XNOR2_X1 U40563 ( .A(n35222), .B(n35221), .ZN(n35223) );
  XNOR2_X1 U40564 ( .A(n35224), .B(n35223), .ZN(n35225) );
  XNOR2_X1 U40565 ( .A(n35226), .B(n35225), .ZN(n35228) );
  XNOR2_X1 U40566 ( .A(n35227), .B(n35633), .ZN(n37077) );
  INV_X1 U40567 ( .A(n51497), .ZN(n35231) );
  XNOR2_X1 U40569 ( .A(n36730), .B(n35232), .ZN(n35245) );
  INV_X1 U40570 ( .A(n44889), .ZN(n35235) );
  XNOR2_X1 U40571 ( .A(n35233), .B(n4826), .ZN(n35234) );
  XNOR2_X1 U40572 ( .A(n35235), .B(n35234), .ZN(n35236) );
  XNOR2_X1 U40573 ( .A(n35237), .B(n35236), .ZN(n35239) );
  XNOR2_X1 U40574 ( .A(n35239), .B(n35238), .ZN(n35242) );
  XNOR2_X1 U40575 ( .A(n37114), .B(n37108), .ZN(n35241) );
  XNOR2_X1 U40576 ( .A(n35242), .B(n35241), .ZN(n35243) );
  XNOR2_X1 U40577 ( .A(n36959), .B(n35243), .ZN(n35244) );
  NAND2_X1 U40578 ( .A1(n38259), .A2(n51360), .ZN(n37224) );
  XNOR2_X1 U40579 ( .A(n35829), .B(n35589), .ZN(n35246) );
  XNOR2_X1 U40580 ( .A(n35246), .B(n36857), .ZN(n35248) );
  XNOR2_X1 U40581 ( .A(n37040), .B(n35250), .ZN(n35258) );
  XNOR2_X1 U40582 ( .A(n35252), .B(n35251), .ZN(n35253) );
  XNOR2_X1 U40583 ( .A(n35254), .B(n35253), .ZN(n35256) );
  XNOR2_X1 U40584 ( .A(n35255), .B(n45463), .ZN(n35842) );
  XNOR2_X1 U40585 ( .A(n35256), .B(n35842), .ZN(n35257) );
  XNOR2_X1 U40586 ( .A(n35258), .B(n35257), .ZN(n35259) );
  XNOR2_X1 U40588 ( .A(n33195), .B(n52148), .ZN(n35264) );
  XNOR2_X1 U40589 ( .A(n40107), .B(n35261), .ZN(n35262) );
  XNOR2_X1 U40590 ( .A(n37066), .B(n35262), .ZN(n35263) );
  XNOR2_X1 U40591 ( .A(n35264), .B(n35263), .ZN(n35267) );
  XNOR2_X1 U40592 ( .A(n35265), .B(n37243), .ZN(n35266) );
  XNOR2_X1 U40593 ( .A(n35762), .B(n35683), .ZN(n35275) );
  XNOR2_X1 U40594 ( .A(n35270), .B(n4706), .ZN(n35271) );
  XNOR2_X1 U40595 ( .A(n35272), .B(n35271), .ZN(n35273) );
  XNOR2_X1 U40596 ( .A(n35275), .B(n35274), .ZN(n35277) );
  XNOR2_X1 U40597 ( .A(n35277), .B(n35276), .ZN(n35279) );
  XNOR2_X1 U40598 ( .A(n35278), .B(n35279), .ZN(n35281) );
  XNOR2_X1 U40599 ( .A(n35281), .B(n35280), .ZN(n35284) );
  XNOR2_X1 U40600 ( .A(n35283), .B(n37329), .ZN(n37005) );
  INV_X1 U40601 ( .A(n35304), .ZN(n35305) );
  INV_X1 U40602 ( .A(n35285), .ZN(n37136) );
  XNOR2_X1 U40603 ( .A(n37136), .B(n35286), .ZN(n35288) );
  INV_X1 U40604 ( .A(n517), .ZN(n35287) );
  XNOR2_X1 U40605 ( .A(n35288), .B(n35287), .ZN(n37311) );
  XNOR2_X1 U40606 ( .A(n35289), .B(n36747), .ZN(n35295) );
  XNOR2_X1 U40607 ( .A(n35290), .B(n1224), .ZN(n35291) );
  XNOR2_X1 U40608 ( .A(n35292), .B(n35291), .ZN(n35293) );
  XNOR2_X1 U40609 ( .A(n35295), .B(n35294), .ZN(n35297) );
  XNOR2_X1 U40610 ( .A(n35297), .B(n35296), .ZN(n35298) );
  XNOR2_X1 U40611 ( .A(n37311), .B(n35298), .ZN(n35299) );
  INV_X1 U40612 ( .A(n38258), .ZN(n35310) );
  NAND3_X1 U40613 ( .A1(n37219), .A2(n68), .A3(n38630), .ZN(n35300) );
  AND2_X1 U40614 ( .A1(n38627), .A2(n35300), .ZN(n35301) );
  NAND2_X1 U40617 ( .A1(n68), .A2(n35310), .ZN(n37680) );
  INV_X1 U40618 ( .A(n38259), .ZN(n38628) );
  NAND2_X1 U40619 ( .A1(n38640), .A2(n38641), .ZN(n35307) );
  OAI211_X1 U40620 ( .C1(n37689), .C2(n38635), .A(n38252), .B(n38630), .ZN(
        n35306) );
  OAI211_X1 U40621 ( .C1(n35308), .C2(n37680), .A(n35307), .B(n35306), .ZN(
        n35309) );
  INV_X1 U40622 ( .A(n35309), .ZN(n35432) );
  NAND2_X1 U40623 ( .A1(n35311), .A2(n36558), .ZN(n35312) );
  AND2_X1 U40624 ( .A1(n35313), .A2(n35312), .ZN(n35324) );
  OAI21_X1 U40625 ( .B1(n35314), .B2(n36565), .A(n36491), .ZN(n35316) );
  AND2_X1 U40626 ( .A1(n36480), .A2(n35316), .ZN(n35323) );
  INV_X1 U40627 ( .A(n36494), .ZN(n36559) );
  INV_X1 U40628 ( .A(n36558), .ZN(n35317) );
  OAI211_X1 U40629 ( .C1(n36559), .C2(n458), .A(n36557), .B(n35317), .ZN(
        n35318) );
  NAND2_X1 U40630 ( .A1(n35318), .A2(n36572), .ZN(n35322) );
  NAND2_X1 U40631 ( .A1(n458), .A2(n36493), .ZN(n36568) );
  NOR2_X1 U40632 ( .A1(n36568), .A2(n51324), .ZN(n36566) );
  OAI21_X1 U40633 ( .B1(n36566), .B2(n35320), .A(n36492), .ZN(n35321) );
  XNOR2_X1 U40634 ( .A(n35325), .B(n37269), .ZN(n35811) );
  XNOR2_X1 U40635 ( .A(n35326), .B(n35811), .ZN(n35327) );
  XNOR2_X1 U40636 ( .A(n35328), .B(n1354), .ZN(n35329) );
  XNOR2_X1 U40637 ( .A(n40849), .B(n35329), .ZN(n35330) );
  XNOR2_X1 U40638 ( .A(n35331), .B(n35330), .ZN(n35332) );
  XNOR2_X1 U40639 ( .A(n37114), .B(n35332), .ZN(n35336) );
  XNOR2_X1 U40640 ( .A(n35333), .B(n35334), .ZN(n35335) );
  XNOR2_X1 U40641 ( .A(n35336), .B(n35335), .ZN(n35338) );
  XNOR2_X1 U40642 ( .A(n35338), .B(n35337), .ZN(n35339) );
  XNOR2_X1 U40643 ( .A(n35340), .B(n43691), .ZN(n35341) );
  XNOR2_X1 U40644 ( .A(n35342), .B(n35341), .ZN(n35343) );
  XNOR2_X1 U40645 ( .A(n36981), .B(n35343), .ZN(n35344) );
  XNOR2_X1 U40646 ( .A(n35344), .B(n35537), .ZN(n35347) );
  INV_X1 U40647 ( .A(n35352), .ZN(n35354) );
  XNOR2_X1 U40648 ( .A(n35354), .B(n35353), .ZN(n35355) );
  XNOR2_X1 U40649 ( .A(n37067), .B(n35355), .ZN(n35356) );
  XNOR2_X1 U40650 ( .A(n35265), .B(n35356), .ZN(n35357) );
  XNOR2_X1 U40651 ( .A(n35358), .B(n35357), .ZN(n35359) );
  NOR2_X1 U40652 ( .A1(n38338), .A2(n37665), .ZN(n37673) );
  XNOR2_X1 U40653 ( .A(n36856), .B(n36858), .ZN(n35368) );
  XNOR2_X1 U40654 ( .A(n35361), .B(n4934), .ZN(n35362) );
  XNOR2_X1 U40655 ( .A(n35363), .B(n35362), .ZN(n35364) );
  XNOR2_X1 U40656 ( .A(n35589), .B(n35364), .ZN(n35365) );
  XNOR2_X1 U40657 ( .A(n35366), .B(n35365), .ZN(n35367) );
  XNOR2_X1 U40658 ( .A(n35368), .B(n35367), .ZN(n35370) );
  XNOR2_X1 U40659 ( .A(n35371), .B(n35372), .ZN(n35373) );
  NOR2_X1 U40661 ( .A1(n35889), .A2(n36468), .ZN(n35390) );
  INV_X1 U40662 ( .A(n35374), .ZN(n35375) );
  XNOR2_X1 U40663 ( .A(n37136), .B(n35375), .ZN(n37024) );
  INV_X1 U40664 ( .A(n35376), .ZN(n35379) );
  XNOR2_X1 U40665 ( .A(n35377), .B(n4883), .ZN(n35378) );
  XNOR2_X1 U40666 ( .A(n35379), .B(n35378), .ZN(n35381) );
  XNOR2_X1 U40667 ( .A(n35381), .B(n35380), .ZN(n35382) );
  XNOR2_X1 U40668 ( .A(n35383), .B(n35382), .ZN(n35384) );
  XNOR2_X1 U40669 ( .A(n37024), .B(n35384), .ZN(n35389) );
  XNOR2_X1 U40670 ( .A(n35745), .B(n4793), .ZN(n35385) );
  XNOR2_X1 U40671 ( .A(n35386), .B(n35385), .ZN(n35388) );
  INV_X1 U40672 ( .A(n35387), .ZN(n35475) );
  XNOR2_X1 U40673 ( .A(n35388), .B(n35475), .ZN(n37309) );
  XNOR2_X1 U40674 ( .A(n35391), .B(n35669), .ZN(n35400) );
  INV_X1 U40675 ( .A(n35392), .ZN(n35395) );
  XNOR2_X1 U40676 ( .A(n35393), .B(n49414), .ZN(n35394) );
  XNOR2_X1 U40677 ( .A(n35395), .B(n35394), .ZN(n35396) );
  XNOR2_X1 U40678 ( .A(n37325), .B(n35396), .ZN(n35397) );
  XNOR2_X1 U40679 ( .A(n52220), .B(n35397), .ZN(n35399) );
  XNOR2_X1 U40680 ( .A(n35400), .B(n35399), .ZN(n35401) );
  NAND2_X1 U40681 ( .A1(n37670), .A2(n38329), .ZN(n37188) );
  NOR2_X1 U40682 ( .A1(n37188), .A2(n37190), .ZN(n37669) );
  INV_X1 U40683 ( .A(n35406), .ZN(n37191) );
  NOR2_X1 U40684 ( .A1(n37664), .A2(n37670), .ZN(n35408) );
  AOI21_X1 U40685 ( .B1(n37669), .B2(n35894), .A(n35408), .ZN(n35413) );
  NAND3_X1 U40686 ( .A1(n35893), .A2(n38337), .A3(n37188), .ZN(n35412) );
  AND2_X1 U40687 ( .A1(n40014), .A2(n39097), .ZN(n39995) );
  AOI22_X1 U40688 ( .A1(n35415), .A2(n38284), .B1(n38292), .B2(n38282), .ZN(
        n35421) );
  NOR2_X1 U40689 ( .A1(n35416), .A2(n38279), .ZN(n36440) );
  NAND2_X1 U40690 ( .A1(n36440), .A2(n38291), .ZN(n35419) );
  NAND4_X1 U40691 ( .A1(n35417), .A2(n613), .A3(n37617), .A4(n38275), .ZN(
        n35418) );
  NAND4_X1 U40692 ( .A1(n35421), .A2(n35420), .A3(n35419), .A4(n35418), .ZN(
        n35428) );
  AOI21_X1 U40693 ( .B1(n51339), .B2(n38275), .A(n38270), .ZN(n35422) );
  OAI211_X1 U40694 ( .C1(n38271), .C2(n38270), .A(n37629), .B(n37624), .ZN(
        n35423) );
  OAI211_X1 U40695 ( .C1(n37618), .C2(n35424), .A(n35423), .B(n37623), .ZN(
        n35425) );
  AOI21_X1 U40696 ( .B1(n35426), .B2(n38279), .A(n35425), .ZN(n35427) );
  INV_X1 U40697 ( .A(n40003), .ZN(n39668) );
  INV_X1 U40698 ( .A(n35429), .ZN(n35430) );
  OR2_X1 U40699 ( .A1(n35432), .A2(n39667), .ZN(n35433) );
  AND2_X1 U40700 ( .A1(n39097), .A2(n39667), .ZN(n38429) );
  NAND2_X1 U40701 ( .A1(n38429), .A2(n39098), .ZN(n40008) );
  NAND2_X1 U40702 ( .A1(n39099), .A2(n40003), .ZN(n35436) );
  MUX2_X1 U40703 ( .A(n35437), .B(n35436), .S(n40015), .Z(n35438) );
  NAND2_X1 U40704 ( .A1(n37415), .A2(n38119), .ZN(n35440) );
  AND2_X1 U40705 ( .A1(n35441), .A2(n35440), .ZN(n35450) );
  OAI21_X1 U40706 ( .B1(n38468), .B2(n38464), .A(n38481), .ZN(n35444) );
  AND2_X1 U40707 ( .A1(n1950), .A2(n38484), .ZN(n35443) );
  NOR2_X1 U40708 ( .A1(n38108), .A2(n37416), .ZN(n37426) );
  INV_X1 U40709 ( .A(n38478), .ZN(n35445) );
  OAI21_X1 U40711 ( .B1(n37414), .B2(n38475), .A(n6637), .ZN(n35446) );
  INV_X1 U40713 ( .A(n37598), .ZN(n35977) );
  NAND2_X1 U40714 ( .A1(n35977), .A2(n37376), .ZN(n35456) );
  OR2_X1 U40715 ( .A1(n37585), .A2(n37596), .ZN(n35979) );
  NAND3_X1 U40716 ( .A1(n35979), .A2(n35980), .A3(n37587), .ZN(n35455) );
  INV_X1 U40718 ( .A(n36222), .ZN(n37364) );
  NAND3_X1 U40719 ( .A1(n37591), .A2(n37587), .A3(n37371), .ZN(n35451) );
  NAND3_X1 U40720 ( .A1(n37376), .A2(n37592), .A3(n37585), .ZN(n37368) );
  NAND3_X1 U40721 ( .A1(n37586), .A2(n37592), .A3(n37377), .ZN(n36228) );
  OAI22_X1 U40722 ( .A1(n37379), .A2(n37593), .B1(n37378), .B2(n37372), .ZN(
        n35459) );
  AND2_X1 U40723 ( .A1(n35458), .A2(n36232), .ZN(n37382) );
  NAND2_X1 U40724 ( .A1(n35459), .A2(n37382), .ZN(n35461) );
  NAND2_X1 U40725 ( .A1(n36231), .A2(n35973), .ZN(n35460) );
  NAND3_X1 U40726 ( .A1(n36228), .A2(n35461), .A3(n35460), .ZN(n35462) );
  XNOR2_X1 U40727 ( .A(n36819), .B(n35464), .ZN(n35473) );
  XNOR2_X1 U40728 ( .A(n35466), .B(n35465), .ZN(n35467) );
  XNOR2_X1 U40729 ( .A(n35468), .B(n35467), .ZN(n35469) );
  XNOR2_X1 U40730 ( .A(n35469), .B(n37015), .ZN(n35470) );
  XNOR2_X1 U40731 ( .A(n51493), .B(n35470), .ZN(n35472) );
  XNOR2_X1 U40732 ( .A(n35476), .B(n35475), .ZN(n35758) );
  XNOR2_X1 U40733 ( .A(n35480), .B(n35479), .ZN(n35481) );
  XNOR2_X1 U40734 ( .A(n35482), .B(n35481), .ZN(n35484) );
  XNOR2_X1 U40735 ( .A(n35484), .B(n35483), .ZN(n35485) );
  XNOR2_X1 U40736 ( .A(n35487), .B(n35486), .ZN(n35492) );
  XNOR2_X1 U40737 ( .A(n35488), .B(n35668), .ZN(n35489) );
  XNOR2_X1 U40738 ( .A(n35490), .B(n35489), .ZN(n35491) );
  INV_X1 U40739 ( .A(n35493), .ZN(n35495) );
  XNOR2_X1 U40740 ( .A(n35495), .B(n35494), .ZN(n35508) );
  XNOR2_X1 U40742 ( .A(n35497), .B(n4923), .ZN(n35498) );
  XNOR2_X1 U40743 ( .A(n35499), .B(n35498), .ZN(n35500) );
  XNOR2_X1 U40744 ( .A(n36855), .B(n35500), .ZN(n35502) );
  XNOR2_X1 U40745 ( .A(n35502), .B(n35501), .ZN(n35504) );
  XNOR2_X1 U40746 ( .A(n35503), .B(n35589), .ZN(n35837) );
  XNOR2_X1 U40749 ( .A(n35508), .B(n35507), .ZN(n35531) );
  XNOR2_X1 U40750 ( .A(n36671), .B(n35509), .ZN(n35511) );
  BUF_X2 U40751 ( .A(n35510), .Z(n37243) );
  XNOR2_X1 U40752 ( .A(n37243), .B(n35511), .ZN(n35788) );
  XNOR2_X1 U40753 ( .A(n35512), .B(n4687), .ZN(n35607) );
  XNOR2_X1 U40754 ( .A(n35513), .B(n35607), .ZN(n35515) );
  INV_X1 U40755 ( .A(n35517), .ZN(n35527) );
  XNOR2_X1 U40756 ( .A(n37067), .B(n35778), .ZN(n35525) );
  XNOR2_X1 U40757 ( .A(n35518), .B(n48814), .ZN(n35519) );
  XNOR2_X1 U40758 ( .A(n35520), .B(n35519), .ZN(n35521) );
  XNOR2_X1 U40759 ( .A(n35522), .B(n35521), .ZN(n35523) );
  XNOR2_X1 U40760 ( .A(n35525), .B(n35524), .ZN(n35526) );
  XNOR2_X1 U40761 ( .A(n35527), .B(n35526), .ZN(n35528) );
  XNOR2_X2 U40762 ( .A(n35528), .B(n35529), .ZN(n37489) );
  NAND2_X1 U40763 ( .A1(n35531), .A2(n37489), .ZN(n38530) );
  INV_X1 U40764 ( .A(n38530), .ZN(n38512) );
  OAI22_X1 U40767 ( .A1(n35960), .A2(n38535), .B1(n37437), .B2(n35966), .ZN(
        n35550) );
  XNOR2_X1 U40768 ( .A(n37081), .B(n35533), .ZN(n35535) );
  XNOR2_X1 U40769 ( .A(n35534), .B(n35535), .ZN(n35806) );
  XNOR2_X1 U40770 ( .A(n36792), .B(n35536), .ZN(n35538) );
  XNOR2_X1 U40771 ( .A(n35538), .B(n35537), .ZN(n37296) );
  XNOR2_X1 U40772 ( .A(n35539), .B(n47737), .ZN(n35540) );
  XNOR2_X1 U40773 ( .A(n35541), .B(n35540), .ZN(n35542) );
  XNOR2_X1 U40774 ( .A(n35543), .B(n35542), .ZN(n35545) );
  INV_X1 U40775 ( .A(n35544), .ZN(n35645) );
  XNOR2_X1 U40776 ( .A(n35545), .B(n35645), .ZN(n35547) );
  XNOR2_X1 U40777 ( .A(n35547), .B(n35546), .ZN(n35548) );
  NAND2_X1 U40778 ( .A1(n35550), .A2(n36161), .ZN(n35570) );
  INV_X1 U40779 ( .A(n35551), .ZN(n35565) );
  INV_X1 U40780 ( .A(n35552), .ZN(n35560) );
  XNOR2_X1 U40781 ( .A(n35554), .B(n35553), .ZN(n35555) );
  XNOR2_X1 U40782 ( .A(n35625), .B(n35555), .ZN(n35556) );
  INV_X1 U40785 ( .A(n35561), .ZN(n35562) );
  AOI21_X1 U40786 ( .B1(n38529), .B2(n51411), .A(n37442), .ZN(n35566) );
  NOR2_X1 U40787 ( .A1(n38522), .A2(n51363), .ZN(n35567) );
  AND2_X1 U40788 ( .A1(n35567), .A2(n37442), .ZN(n37483) );
  AOI22_X1 U40790 ( .A1(n37483), .A2(n38517), .B1(n37442), .B2(n51411), .ZN(
        n35569) );
  OAI21_X1 U40791 ( .B1(n37437), .B2(n617), .A(n37490), .ZN(n37436) );
  NOR2_X1 U40792 ( .A1(n37436), .A2(n38535), .ZN(n35568) );
  NAND2_X1 U40793 ( .A1(n51735), .A2(n35568), .ZN(n38538) );
  INV_X1 U40795 ( .A(n35571), .ZN(n35572) );
  INV_X1 U40796 ( .A(n38493), .ZN(n38506) );
  NAND2_X1 U40797 ( .A1(n37531), .A2(n37520), .ZN(n38502) );
  NOR2_X1 U40798 ( .A1(n35951), .A2(n38504), .ZN(n35575) );
  AOI22_X1 U40799 ( .A1(n35577), .A2(n35576), .B1(n38502), .B2(n35575), .ZN(
        n35584) );
  NOR2_X1 U40800 ( .A1(n37521), .A2(n38494), .ZN(n35582) );
  OAI21_X1 U40801 ( .B1(n37520), .B2(n37384), .A(n38504), .ZN(n35581) );
  NAND2_X1 U40803 ( .A1(n35579), .A2(n35949), .ZN(n35580) );
  OAI211_X1 U40804 ( .C1(n35582), .C2(n35581), .A(n35580), .B(n35951), .ZN(
        n35583) );
  XNOR2_X1 U40806 ( .A(n35589), .B(n35588), .ZN(n37253) );
  XNOR2_X1 U40807 ( .A(n37047), .B(n37253), .ZN(n35597) );
  XNOR2_X1 U40808 ( .A(n35590), .B(n4865), .ZN(n35591) );
  XNOR2_X1 U40809 ( .A(n35592), .B(n35591), .ZN(n35593) );
  XNOR2_X1 U40810 ( .A(n36939), .B(n35593), .ZN(n35594) );
  XNOR2_X1 U40811 ( .A(n35595), .B(n35594), .ZN(n35596) );
  XNOR2_X1 U40812 ( .A(n35597), .B(n35596), .ZN(n35598) );
  XNOR2_X1 U40813 ( .A(n35599), .B(n35598), .ZN(n35602) );
  INV_X1 U40814 ( .A(n35600), .ZN(n35601) );
  INV_X1 U40815 ( .A(n35603), .ZN(n37249) );
  XNOR2_X1 U40816 ( .A(n43076), .B(n35604), .ZN(n35605) );
  XNOR2_X1 U40817 ( .A(n35606), .B(n35605), .ZN(n35608) );
  XNOR2_X1 U40818 ( .A(n35608), .B(n35607), .ZN(n35611) );
  XNOR2_X1 U40819 ( .A(n35778), .B(n35609), .ZN(n35610) );
  XNOR2_X1 U40820 ( .A(n35611), .B(n35610), .ZN(n35613) );
  XNOR2_X1 U40821 ( .A(n35612), .B(n35613), .ZN(n35616) );
  INV_X1 U40822 ( .A(n35614), .ZN(n35615) );
  XNOR2_X1 U40823 ( .A(n35616), .B(n35615), .ZN(n35617) );
  INV_X1 U40824 ( .A(n38589), .ZN(n38156) );
  XNOR2_X1 U40825 ( .A(n35623), .B(n35622), .ZN(n35624) );
  XNOR2_X1 U40826 ( .A(n35625), .B(n35624), .ZN(n35626) );
  XNOR2_X1 U40827 ( .A(n36807), .B(n35626), .ZN(n35628) );
  XNOR2_X1 U40828 ( .A(n35627), .B(n35628), .ZN(n35629) );
  XNOR2_X1 U40829 ( .A(n35632), .B(n35633), .ZN(n35634) );
  XNOR2_X1 U40830 ( .A(n35635), .B(n35634), .ZN(n35636) );
  XNOR2_X1 U40831 ( .A(n35636), .B(n37284), .ZN(n35639) );
  INV_X1 U40832 ( .A(n35637), .ZN(n35638) );
  XNOR2_X1 U40833 ( .A(n35639), .B(n35638), .ZN(n35652) );
  INV_X1 U40834 ( .A(n35640), .ZN(n35643) );
  XNOR2_X1 U40835 ( .A(n35641), .B(n43691), .ZN(n35642) );
  XNOR2_X1 U40836 ( .A(n35643), .B(n35642), .ZN(n35644) );
  XNOR2_X1 U40837 ( .A(n35646), .B(n35645), .ZN(n35647) );
  XNOR2_X1 U40838 ( .A(n35648), .B(n35647), .ZN(n35650) );
  XNOR2_X1 U40839 ( .A(n35650), .B(n35649), .ZN(n35651) );
  XNOR2_X2 U40840 ( .A(n35652), .B(n35651), .ZN(n38599) );
  INV_X1 U40841 ( .A(n38599), .ZN(n38159) );
  INV_X1 U40843 ( .A(n37580), .ZN(n38167) );
  XNOR2_X1 U40844 ( .A(n35653), .B(n4605), .ZN(n35655) );
  XNOR2_X1 U40845 ( .A(n35656), .B(n35657), .ZN(n35658) );
  XNOR2_X1 U40846 ( .A(n35658), .B(n518), .ZN(n35661) );
  INV_X1 U40847 ( .A(n35659), .ZN(n35660) );
  XNOR2_X1 U40848 ( .A(n35660), .B(n35661), .ZN(n35663) );
  XNOR2_X1 U40849 ( .A(n35663), .B(n35662), .ZN(n35665) );
  XNOR2_X1 U40851 ( .A(n35669), .B(n35668), .ZN(n35670) );
  XNOR2_X1 U40852 ( .A(n35671), .B(n35670), .ZN(n35682) );
  XNOR2_X1 U40853 ( .A(n35673), .B(n35672), .ZN(n42476) );
  XNOR2_X1 U40854 ( .A(n35674), .B(n4931), .ZN(n35675) );
  XNOR2_X1 U40855 ( .A(n42476), .B(n35675), .ZN(n35676) );
  XNOR2_X1 U40856 ( .A(n36999), .B(n35676), .ZN(n35677) );
  XNOR2_X1 U40857 ( .A(n51366), .B(n35677), .ZN(n35679) );
  XNOR2_X1 U40858 ( .A(n35680), .B(n35679), .ZN(n35681) );
  XNOR2_X1 U40859 ( .A(n35682), .B(n35681), .ZN(n35686) );
  XNOR2_X1 U40860 ( .A(n36766), .B(n35683), .ZN(n35684) );
  XNOR2_X1 U40861 ( .A(n35685), .B(n35684), .ZN(n37331) );
  INV_X1 U40862 ( .A(n35693), .ZN(n38164) );
  NAND4_X1 U40863 ( .A1(n38584), .A2(n38166), .A3(n38592), .A4(n38164), .ZN(
        n35687) );
  AND2_X1 U40864 ( .A1(n35688), .A2(n35687), .ZN(n35699) );
  OAI21_X1 U40865 ( .B1(n37580), .B2(n38165), .A(n37569), .ZN(n35689) );
  NAND3_X1 U40866 ( .A1(n35689), .A2(n38593), .A3(n38589), .ZN(n35692) );
  NOR2_X1 U40867 ( .A1(n37448), .A2(n38165), .ZN(n37577) );
  INV_X1 U40868 ( .A(n37577), .ZN(n35691) );
  INV_X1 U40869 ( .A(n38590), .ZN(n36132) );
  AND2_X1 U40870 ( .A1(n38592), .A2(n38159), .ZN(n37576) );
  NAND2_X1 U40871 ( .A1(n36133), .A2(n38585), .ZN(n35694) );
  OR2_X1 U40872 ( .A1(n37569), .A2(n35694), .ZN(n37579) );
  NOR2_X1 U40873 ( .A1(n52159), .A2(n40556), .ZN(n35700) );
  NAND2_X1 U40874 ( .A1(n40146), .A2(n35700), .ZN(n35725) );
  AND2_X1 U40876 ( .A1(n40558), .A2(n4951), .ZN(n35719) );
  INV_X1 U40877 ( .A(n38573), .ZN(n35705) );
  INV_X1 U40878 ( .A(n38205), .ZN(n35701) );
  OAI211_X1 U40879 ( .C1(n689), .C2(n35705), .A(n35702), .B(n35701), .ZN(
        n35703) );
  NAND2_X1 U40880 ( .A1(n35703), .A2(n38204), .ZN(n35717) );
  INV_X1 U40881 ( .A(n35704), .ZN(n35710) );
  AND2_X1 U40883 ( .A1(n35706), .A2(n481), .ZN(n35708) );
  INV_X1 U40884 ( .A(n38567), .ZN(n38571) );
  OAI21_X1 U40885 ( .B1(n38201), .B2(n591), .A(n38571), .ZN(n35707) );
  AOI22_X1 U40886 ( .A1(n35710), .A2(n35709), .B1(n35708), .B2(n35707), .ZN(
        n35716) );
  INV_X1 U40887 ( .A(n36103), .ZN(n35712) );
  NOR2_X1 U40888 ( .A1(n35712), .A2(n35711), .ZN(n35714) );
  NAND2_X1 U40889 ( .A1(n40316), .A2(n40565), .ZN(n40157) );
  INV_X1 U40890 ( .A(n40157), .ZN(n40571) );
  OAI21_X1 U40891 ( .B1(n39653), .B2(n4951), .A(n40151), .ZN(n35720) );
  NAND2_X1 U40892 ( .A1(n35720), .A2(n40559), .ZN(n35724) );
  OAI21_X1 U40893 ( .B1(n40316), .B2(n40565), .A(n40558), .ZN(n35721) );
  OAI21_X1 U40894 ( .B1(n40315), .B2(n40556), .A(n35721), .ZN(n35722) );
  NAND2_X1 U40895 ( .A1(n35722), .A2(n40311), .ZN(n35723) );
  NAND3_X1 U40896 ( .A1(n34632), .A2(n37648), .A3(n37636), .ZN(n36404) );
  NAND4_X1 U40897 ( .A1(n36404), .A2(n5588), .A3(n36410), .A4(n36402), .ZN(
        n35727) );
  NAND2_X1 U40898 ( .A1(n37640), .A2(n34632), .ZN(n35730) );
  NAND2_X1 U40899 ( .A1(n2141), .A2(n35728), .ZN(n35729) );
  NAND4_X1 U40900 ( .A1(n35730), .A2(n35729), .A3(n37646), .A4(n36404), .ZN(
        n35731) );
  INV_X1 U40901 ( .A(n36397), .ZN(n35733) );
  NOR2_X1 U40902 ( .A1(n35733), .A2(n5590), .ZN(n35735) );
  NOR2_X1 U40903 ( .A1(n35733), .A2(n37643), .ZN(n35734) );
  AOI22_X1 U40904 ( .A1(n37644), .A2(n35735), .B1(n35734), .B2(n36398), .ZN(
        n35738) );
  NAND2_X1 U40905 ( .A1(n36398), .A2(n36410), .ZN(n36002) );
  XNOR2_X1 U40906 ( .A(n35741), .B(n4431), .ZN(n35742) );
  XNOR2_X1 U40907 ( .A(n35743), .B(n35742), .ZN(n35744) );
  XNOR2_X1 U40908 ( .A(n35745), .B(n35744), .ZN(n35746) );
  XNOR2_X1 U40909 ( .A(n35748), .B(n35749), .ZN(n35750) );
  XNOR2_X1 U40911 ( .A(n37307), .B(n35753), .ZN(n35754) );
  XNOR2_X1 U40912 ( .A(n35755), .B(n35754), .ZN(n35757) );
  XNOR2_X1 U40913 ( .A(n35757), .B(n35756), .ZN(n35759) );
  XNOR2_X1 U40914 ( .A(n35761), .B(n35762), .ZN(n35763) );
  XNOR2_X1 U40915 ( .A(n35764), .B(n35763), .ZN(n35771) );
  XNOR2_X1 U40916 ( .A(n35766), .B(n35765), .ZN(n35767) );
  XNOR2_X1 U40917 ( .A(n52071), .B(n35767), .ZN(n35769) );
  XNOR2_X1 U40918 ( .A(n35769), .B(n37325), .ZN(n35770) );
  XNOR2_X1 U40919 ( .A(n35771), .B(n35770), .ZN(n35773) );
  XNOR2_X1 U40920 ( .A(n35773), .B(n35772), .ZN(n35774) );
  INV_X1 U40921 ( .A(n35775), .ZN(n35787) );
  XNOR2_X1 U40922 ( .A(n51447), .B(n43878), .ZN(n35777) );
  XNOR2_X1 U40923 ( .A(n35778), .B(n35777), .ZN(n37244) );
  INV_X1 U40924 ( .A(n35779), .ZN(n35784) );
  XNOR2_X1 U40925 ( .A(n35781), .B(n35780), .ZN(n35782) );
  XNOR2_X1 U40926 ( .A(n36841), .B(n35782), .ZN(n35783) );
  XNOR2_X1 U40927 ( .A(n35784), .B(n35783), .ZN(n35785) );
  XNOR2_X1 U40928 ( .A(n37244), .B(n35785), .ZN(n35786) );
  XNOR2_X1 U40929 ( .A(n35787), .B(n35786), .ZN(n35794) );
  INV_X1 U40930 ( .A(n35788), .ZN(n35792) );
  XNOR2_X1 U40931 ( .A(n37241), .B(n36672), .ZN(n35789) );
  XNOR2_X1 U40932 ( .A(n35790), .B(n35789), .ZN(n37074) );
  INV_X1 U40933 ( .A(n37074), .ZN(n35791) );
  XNOR2_X1 U40934 ( .A(n35792), .B(n35791), .ZN(n35793) );
  XNOR2_X1 U40935 ( .A(n35794), .B(n35793), .ZN(n35849) );
  INV_X1 U40937 ( .A(n35795), .ZN(n35797) );
  XNOR2_X1 U40938 ( .A(n35797), .B(n35796), .ZN(n35799) );
  XNOR2_X1 U40939 ( .A(n35801), .B(n36703), .ZN(n35802) );
  XNOR2_X1 U40940 ( .A(n35804), .B(n37294), .ZN(n35805) );
  INV_X1 U40941 ( .A(n35808), .ZN(n36801) );
  XNOR2_X1 U40942 ( .A(n35810), .B(n35809), .ZN(n35812) );
  XNOR2_X1 U40943 ( .A(n35812), .B(n35811), .ZN(n35813) );
  XNOR2_X1 U40944 ( .A(n36801), .B(n35813), .ZN(n35827) );
  INV_X1 U40945 ( .A(n35814), .ZN(n35819) );
  XNOR2_X1 U40946 ( .A(n44887), .B(n35815), .ZN(n35817) );
  XNOR2_X1 U40947 ( .A(n35817), .B(n35816), .ZN(n35818) );
  XNOR2_X1 U40948 ( .A(n35819), .B(n35818), .ZN(n35820) );
  XNOR2_X1 U40949 ( .A(n703), .B(n35821), .ZN(n35823) );
  XNOR2_X1 U40950 ( .A(n35823), .B(n35822), .ZN(n35824) );
  XNOR2_X1 U40951 ( .A(n35825), .B(n35824), .ZN(n35826) );
  XNOR2_X1 U40952 ( .A(n35827), .B(n35826), .ZN(n35828) );
  INV_X1 U40953 ( .A(n35828), .ZN(n39291) );
  XNOR2_X1 U40954 ( .A(n35830), .B(n35829), .ZN(n36865) );
  XNOR2_X1 U40955 ( .A(n37045), .B(n35831), .ZN(n35832) );
  INV_X1 U40956 ( .A(n35833), .ZN(n35834) );
  XNOR2_X1 U40957 ( .A(n35835), .B(n35834), .ZN(n37039) );
  INV_X1 U40958 ( .A(n37039), .ZN(n35836) );
  XNOR2_X1 U40959 ( .A(n35836), .B(n35837), .ZN(n35845) );
  XNOR2_X1 U40960 ( .A(n35839), .B(n35838), .ZN(n35840) );
  XNOR2_X1 U40961 ( .A(n35841), .B(n35840), .ZN(n35843) );
  XNOR2_X1 U40962 ( .A(n35843), .B(n35842), .ZN(n35844) );
  XNOR2_X1 U40963 ( .A(n35845), .B(n35844), .ZN(n35846) );
  XNOR2_X1 U40964 ( .A(n37250), .B(n35846), .ZN(n35848) );
  XNOR2_X1 U40965 ( .A(n35848), .B(n35847), .ZN(n38731) );
  INV_X1 U40966 ( .A(n38731), .ZN(n39289) );
  INV_X1 U40967 ( .A(n35849), .ZN(n39290) );
  INV_X1 U40969 ( .A(n38314), .ZN(n38734) );
  INV_X1 U40970 ( .A(n39293), .ZN(n38716) );
  OAI21_X1 U40971 ( .B1(n38734), .B2(n39289), .A(n38716), .ZN(n35851) );
  NOR2_X1 U40972 ( .A1(n38313), .A2(n38722), .ZN(n35852) );
  NOR2_X1 U40974 ( .A1(n35854), .A2(n35853), .ZN(n35855) );
  NOR2_X1 U40975 ( .A1(n8077), .A2(n37654), .ZN(n38715) );
  NAND2_X1 U40976 ( .A1(n38715), .A2(n38314), .ZN(n39314) );
  INV_X1 U40977 ( .A(n38321), .ZN(n35857) );
  NAND2_X1 U40978 ( .A1(n35857), .A2(n38721), .ZN(n35858) );
  OAI21_X1 U40979 ( .B1(n38272), .B2(n38282), .A(n36436), .ZN(n35861) );
  NAND2_X1 U40980 ( .A1(n37628), .A2(n35861), .ZN(n35865) );
  NAND2_X1 U40981 ( .A1(n37624), .A2(n38276), .ZN(n35864) );
  OAI211_X1 U40982 ( .C1(n38276), .C2(n37624), .A(n38284), .B(n37623), .ZN(
        n35863) );
  NAND3_X1 U40983 ( .A1(n37627), .A2(n38283), .A3(n38272), .ZN(n35862) );
  AND2_X1 U40985 ( .A1(n37617), .A2(n38272), .ZN(n37616) );
  INV_X1 U40986 ( .A(n37616), .ZN(n35868) );
  NAND2_X1 U40987 ( .A1(n613), .A2(n37624), .ZN(n35867) );
  OAI22_X1 U40988 ( .A1(n35868), .A2(n35867), .B1(n38282), .B2(n35866), .ZN(
        n35869) );
  NAND3_X1 U40989 ( .A1(n36054), .A2(n35871), .A3(n36595), .ZN(n36598) );
  INV_X1 U40990 ( .A(n36056), .ZN(n35876) );
  OAI21_X1 U40991 ( .B1(n35876), .B2(n35875), .A(n35874), .ZN(n35885) );
  NAND2_X1 U40992 ( .A1(n36047), .A2(n36045), .ZN(n35877) );
  NAND3_X1 U40993 ( .A1(n35878), .A2(n36591), .A3(n35877), .ZN(n35884) );
  OR2_X1 U40994 ( .A1(n35880), .A2(n35879), .ZN(n36450) );
  INV_X1 U40995 ( .A(n36450), .ZN(n35882) );
  OAI21_X1 U40996 ( .B1(n35882), .B2(n36585), .A(n35881), .ZN(n35883) );
  NAND2_X1 U40997 ( .A1(n39912), .A2(n38445), .ZN(n38438) );
  NOR2_X1 U40998 ( .A1(n38335), .A2(n38330), .ZN(n35888) );
  INV_X1 U40999 ( .A(n38322), .ZN(n38336) );
  NAND2_X1 U41000 ( .A1(n38328), .A2(n2514), .ZN(n35891) );
  NOR2_X1 U41001 ( .A1(n35892), .A2(n35891), .ZN(n35898) );
  INV_X1 U41002 ( .A(n35894), .ZN(n38334) );
  INV_X1 U41003 ( .A(n38346), .ZN(n35896) );
  NAND2_X1 U41004 ( .A1(n38337), .A2(n37670), .ZN(n35895) );
  NAND2_X1 U41005 ( .A1(n38438), .A2(n39907), .ZN(n39781) );
  INV_X1 U41006 ( .A(n37689), .ZN(n35899) );
  INV_X1 U41007 ( .A(n37680), .ZN(n38255) );
  NAND2_X1 U41008 ( .A1(n38257), .A2(n2188), .ZN(n37682) );
  AOI22_X1 U41009 ( .A1(n51360), .A2(n38252), .B1(n38264), .B2(n38637), .ZN(
        n35902) );
  INV_X1 U41010 ( .A(n38640), .ZN(n38261) );
  NAND3_X1 U41011 ( .A1(n38261), .A2(n38629), .A3(n37689), .ZN(n35901) );
  NAND2_X1 U41012 ( .A1(n39908), .A2(n38448), .ZN(n35905) );
  NAND2_X1 U41013 ( .A1(n35905), .A2(n37356), .ZN(n35906) );
  AND2_X1 U41014 ( .A1(n39789), .A2(n51377), .ZN(n35908) );
  OAI21_X1 U41015 ( .B1(n39912), .B2(n38448), .A(n39899), .ZN(n35907) );
  NOR2_X1 U41016 ( .A1(n38455), .A2(n39907), .ZN(n39787) );
  AOI22_X1 U41017 ( .A1(n35908), .A2(n35907), .B1(n39787), .B2(n39908), .ZN(
        n35912) );
  AND2_X1 U41018 ( .A1(n39907), .A2(n37356), .ZN(n39910) );
  NAND3_X1 U41019 ( .A1(n39910), .A2(n39915), .A3(n39912), .ZN(n35911) );
  XNOR2_X1 U41020 ( .A(n39907), .B(n51377), .ZN(n35909) );
  OR2_X1 U41021 ( .A1(n39912), .A2(n39899), .ZN(n39916) );
  INV_X1 U41022 ( .A(n39916), .ZN(n38441) );
  OAI21_X1 U41023 ( .B1(n35909), .B2(n38441), .A(n38440), .ZN(n35910) );
  AND2_X1 U41024 ( .A1(n37757), .A2(n37759), .ZN(n36252) );
  NAND3_X1 U41025 ( .A1(n37766), .A2(n36252), .A3(n37765), .ZN(n35916) );
  NOR2_X1 U41026 ( .A1(n36248), .A2(n37745), .ZN(n35918) );
  AOI21_X1 U41027 ( .B1(n37750), .B2(n37765), .A(n37759), .ZN(n35917) );
  OAI21_X1 U41028 ( .B1(n37749), .B2(n35918), .A(n35917), .ZN(n35920) );
  NAND2_X1 U41030 ( .A1(n35921), .A2(n37757), .ZN(n35922) );
  INV_X1 U41031 ( .A(n36252), .ZN(n36241) );
  NAND2_X1 U41032 ( .A1(n35923), .A2(n36251), .ZN(n37748) );
  INV_X1 U41033 ( .A(n37559), .ZN(n35932) );
  NAND2_X1 U41034 ( .A1(n37558), .A2(n37543), .ZN(n35931) );
  NOR2_X1 U41035 ( .A1(n37399), .A2(n37557), .ZN(n35928) );
  AOI22_X1 U41036 ( .A1(n35928), .A2(n37410), .B1(n37538), .B2(n34676), .ZN(
        n35930) );
  XNOR2_X1 U41037 ( .A(n37538), .B(n525), .ZN(n35935) );
  NAND2_X1 U41038 ( .A1(n37544), .A2(n36272), .ZN(n35933) );
  OAI21_X1 U41039 ( .B1(n525), .B2(n35933), .A(n36268), .ZN(n35934) );
  OAI21_X1 U41040 ( .B1(n35935), .B2(n34676), .A(n35934), .ZN(n35936) );
  NAND3_X1 U41042 ( .A1(n39335), .A2(n36186), .A3(n39342), .ZN(n35938) );
  NAND2_X1 U41043 ( .A1(n35939), .A2(n36200), .ZN(n37773) );
  AOI21_X1 U41044 ( .B1(n35939), .B2(n52054), .A(n36200), .ZN(n35940) );
  NAND3_X1 U41045 ( .A1(n36186), .A2(n36200), .A3(n36189), .ZN(n35941) );
  OAI21_X1 U41046 ( .B1(n36199), .B2(n35942), .A(n39342), .ZN(n35944) );
  INV_X1 U41047 ( .A(n35943), .ZN(n39343) );
  NAND2_X1 U41048 ( .A1(n35944), .A2(n39343), .ZN(n35945) );
  AND2_X1 U41049 ( .A1(n42209), .A2(n41938), .ZN(n40247) );
  INV_X1 U41050 ( .A(n40247), .ZN(n38925) );
  INV_X1 U41051 ( .A(n37517), .ZN(n38503) );
  OR2_X1 U41052 ( .A1(n38503), .A2(n35949), .ZN(n37523) );
  INV_X1 U41053 ( .A(n37523), .ZN(n35947) );
  NAND3_X1 U41054 ( .A1(n35948), .A2(n35947), .A3(n38504), .ZN(n35959) );
  NOR2_X1 U41055 ( .A1(n35950), .A2(n35949), .ZN(n37529) );
  OAI22_X1 U41056 ( .A1(n37521), .A2(n37386), .B1(n35951), .B2(n38495), .ZN(
        n35952) );
  AOI21_X1 U41057 ( .B1(n37527), .B2(n37529), .A(n35952), .ZN(n35958) );
  NAND2_X1 U41058 ( .A1(n35954), .A2(n35953), .ZN(n35957) );
  NAND2_X1 U41059 ( .A1(n35955), .A2(n38496), .ZN(n35956) );
  OR2_X1 U41060 ( .A1(n36159), .A2(n38512), .ZN(n38533) );
  INV_X1 U41061 ( .A(n38533), .ZN(n35961) );
  AND2_X1 U41062 ( .A1(n38530), .A2(n37438), .ZN(n35962) );
  AOI22_X1 U41063 ( .A1(n37437), .A2(n37483), .B1(n37491), .B2(n35962), .ZN(
        n35964) );
  AND2_X1 U41064 ( .A1(n37442), .A2(n38522), .ZN(n38532) );
  NAND3_X1 U41065 ( .A1(n37491), .A2(n38528), .A3(n38530), .ZN(n36155) );
  INV_X1 U41066 ( .A(n38513), .ZN(n37432) );
  NAND2_X1 U41067 ( .A1(n37432), .A2(n37480), .ZN(n35968) );
  OR2_X1 U41068 ( .A1(n35966), .A2(n37489), .ZN(n37445) );
  INV_X1 U41069 ( .A(n37445), .ZN(n35967) );
  AOI21_X1 U41071 ( .B1(n36234), .B2(n35971), .A(n37591), .ZN(n35976) );
  NAND2_X1 U41072 ( .A1(n37372), .A2(n35973), .ZN(n35972) );
  NAND2_X1 U41074 ( .A1(n37366), .A2(n35974), .ZN(n35975) );
  NOR2_X1 U41075 ( .A1(n35976), .A2(n35975), .ZN(n35988) );
  OAI22_X1 U41076 ( .A1(n35977), .A2(n37596), .B1(n37378), .B2(n37594), .ZN(
        n35978) );
  NOR2_X1 U41077 ( .A1(n36225), .A2(n37377), .ZN(n35982) );
  INV_X1 U41078 ( .A(n35979), .ZN(n35981) );
  OR2_X1 U41079 ( .A1(n36222), .A2(n37371), .ZN(n37381) );
  NAND2_X1 U41080 ( .A1(n37592), .A2(n694), .ZN(n35983) );
  AND2_X1 U41082 ( .A1(n37591), .A2(n37585), .ZN(n35984) );
  NAND2_X1 U41083 ( .A1(n35985), .A2(n35984), .ZN(n35986) );
  NAND4_X1 U41084 ( .A1(n41939), .A2(n680), .A3(n40249), .A4(n42201), .ZN(
        n38926) );
  NOR2_X1 U41085 ( .A1(n40250), .A2(n42201), .ZN(n38921) );
  INV_X1 U41086 ( .A(n38921), .ZN(n35989) );
  NAND3_X1 U41087 ( .A1(n35989), .A2(n41939), .A3(n41927), .ZN(n35991) );
  NAND2_X1 U41089 ( .A1(n37824), .A2(n41925), .ZN(n35990) );
  INV_X1 U41090 ( .A(n42201), .ZN(n39543) );
  NOR2_X1 U41091 ( .A1(n41927), .A2(n42201), .ZN(n38931) );
  NAND2_X1 U41092 ( .A1(n42209), .A2(n42201), .ZN(n35992) );
  NAND2_X1 U41093 ( .A1(n35992), .A2(n40250), .ZN(n35995) );
  OAI211_X1 U41094 ( .C1(n38931), .C2(n35995), .A(n35994), .B(n35993), .ZN(
        n35996) );
  XNOR2_X1 U41095 ( .A(n43575), .B(n43238), .ZN(n36298) );
  NAND3_X1 U41096 ( .A1(n51334), .A2(n37636), .A3(n36410), .ZN(n36408) );
  NAND2_X1 U41097 ( .A1(n35997), .A2(n36396), .ZN(n36009) );
  INV_X1 U41098 ( .A(n36400), .ZN(n35999) );
  NOR2_X1 U41099 ( .A1(n37640), .A2(n36401), .ZN(n35998) );
  NOR2_X1 U41100 ( .A1(n35999), .A2(n35998), .ZN(n36008) );
  OAI21_X1 U41101 ( .B1(n36402), .B2(n36000), .A(n36004), .ZN(n36003) );
  NAND2_X1 U41102 ( .A1(n37636), .A2(n37646), .ZN(n36411) );
  AOI21_X1 U41103 ( .B1(n36411), .B2(n37632), .A(n36402), .ZN(n36001) );
  INV_X1 U41104 ( .A(n36004), .ZN(n36005) );
  NAND2_X1 U41105 ( .A1(n36005), .A2(n36397), .ZN(n36006) );
  INV_X1 U41106 ( .A(n36490), .ZN(n36475) );
  NAND2_X1 U41107 ( .A1(n36560), .A2(n36475), .ZN(n36011) );
  AOI22_X1 U41108 ( .A1(n36471), .A2(n36571), .B1(n36491), .B2(n36559), .ZN(
        n36010) );
  MUX2_X1 U41109 ( .A(n36011), .B(n36010), .S(n36492), .Z(n36026) );
  NAND2_X1 U41110 ( .A1(n458), .A2(n36473), .ZN(n36021) );
  INV_X1 U41111 ( .A(n36021), .ZN(n36012) );
  AND2_X1 U41112 ( .A1(n36014), .A2(n36013), .ZN(n36025) );
  NAND2_X1 U41113 ( .A1(n2086), .A2(n36493), .ZN(n36016) );
  OAI22_X1 U41114 ( .A1(n36495), .A2(n36016), .B1(n36557), .B2(n36576), .ZN(
        n36017) );
  AOI21_X1 U41115 ( .B1(n36019), .B2(n36018), .A(n36017), .ZN(n36024) );
  NAND2_X1 U41117 ( .A1(n36495), .A2(n36021), .ZN(n36022) );
  OAI211_X1 U41118 ( .C1(n36498), .C2(n36022), .A(n36567), .B(n36494), .ZN(
        n36023) );
  INV_X1 U41119 ( .A(n37964), .ZN(n36031) );
  AOI21_X1 U41120 ( .B1(n36553), .B2(n36029), .A(n6218), .ZN(n36030) );
  AND2_X1 U41121 ( .A1(n37964), .A2(n51077), .ZN(n36033) );
  NOR2_X1 U41122 ( .A1(n36540), .A2(n37957), .ZN(n36032) );
  AOI22_X1 U41123 ( .A1(n36034), .A2(n36033), .B1(n36032), .B2(n36031), .ZN(
        n36042) );
  NAND2_X1 U41124 ( .A1(n36539), .A2(n6218), .ZN(n36036) );
  AOI21_X1 U41125 ( .B1(n36037), .B2(n36036), .A(n51077), .ZN(n36038) );
  OR2_X1 U41126 ( .A1(n36038), .A2(n36550), .ZN(n36041) );
  NAND2_X1 U41127 ( .A1(n36039), .A2(n36548), .ZN(n36040) );
  NOR2_X1 U41128 ( .A1(n40194), .A2(n40120), .ZN(n38780) );
  NOR2_X1 U41129 ( .A1(n36462), .A2(n36051), .ZN(n36461) );
  NAND2_X1 U41130 ( .A1(n36047), .A2(n696), .ZN(n36451) );
  OAI211_X1 U41131 ( .C1(n36054), .C2(n36051), .A(n36048), .B(n36451), .ZN(
        n36049) );
  OAI21_X1 U41132 ( .B1(n36052), .B2(n36051), .A(n36050), .ZN(n36053) );
  NAND2_X1 U41133 ( .A1(n36054), .A2(n36053), .ZN(n36055) );
  INV_X1 U41134 ( .A(n36058), .ZN(n36061) );
  NAND3_X1 U41135 ( .A1(n36058), .A2(n36616), .A3(n36057), .ZN(n36059) );
  OAI211_X1 U41136 ( .C1(n36424), .C2(n36061), .A(n36060), .B(n36059), .ZN(
        n36072) );
  INV_X1 U41137 ( .A(n36062), .ZN(n36063) );
  NAND3_X1 U41138 ( .A1(n36063), .A2(n36427), .A3(n36610), .ZN(n36070) );
  NAND3_X1 U41139 ( .A1(n36066), .A2(n36065), .A3(n36064), .ZN(n36069) );
  NAND2_X1 U41140 ( .A1(n36426), .A2(n36067), .ZN(n36068) );
  NAND4_X1 U41141 ( .A1(n36070), .A2(n36069), .A3(n36611), .A4(n36068), .ZN(
        n36071) );
  NAND2_X1 U41142 ( .A1(n51352), .A2(n584), .ZN(n38380) );
  INV_X1 U41143 ( .A(n38380), .ZN(n40126) );
  NAND2_X1 U41144 ( .A1(n36073), .A2(n37990), .ZN(n36076) );
  NAND2_X1 U41145 ( .A1(n37985), .A2(n36518), .ZN(n36074) );
  AND4_X1 U41146 ( .A1(n36522), .A2(n36516), .A3(n37975), .A4(n36074), .ZN(
        n36075) );
  AOI21_X1 U41147 ( .B1(n36076), .B2(n36525), .A(n36075), .ZN(n36091) );
  NAND3_X1 U41148 ( .A1(n37991), .A2(n36077), .A3(n36524), .ZN(n36078) );
  AND2_X1 U41149 ( .A1(n36079), .A2(n36078), .ZN(n36090) );
  NAND2_X1 U41150 ( .A1(n37988), .A2(n37976), .ZN(n36081) );
  AND2_X1 U41151 ( .A1(n507), .A2(n584), .ZN(n36085) );
  NAND2_X1 U41152 ( .A1(n40125), .A2(n40110), .ZN(n38769) );
  AND2_X1 U41153 ( .A1(n40119), .A2(n584), .ZN(n36084) );
  NOR2_X1 U41154 ( .A1(n40125), .A2(n584), .ZN(n40114) );
  NAND2_X1 U41156 ( .A1(n36086), .A2(n37975), .ZN(n36089) );
  NAND3_X1 U41157 ( .A1(n36087), .A2(n37977), .A3(n37975), .ZN(n36088) );
  OAI21_X1 U41159 ( .B1(n38781), .B2(n38782), .A(n36094), .ZN(n36092) );
  NAND2_X1 U41160 ( .A1(n36092), .A2(n40120), .ZN(n36093) );
  INV_X1 U41161 ( .A(n40121), .ZN(n40203) );
  AND2_X1 U41162 ( .A1(n40121), .A2(n2153), .ZN(n38777) );
  INV_X1 U41163 ( .A(n40125), .ZN(n40204) );
  NOR2_X1 U41164 ( .A1(n38562), .A2(n33062), .ZN(n38199) );
  NOR2_X1 U41165 ( .A1(n38204), .A2(n38569), .ZN(n36097) );
  NAND2_X1 U41166 ( .A1(n38576), .A2(n481), .ZN(n36102) );
  NAND3_X1 U41167 ( .A1(n38567), .A2(n38201), .A3(n481), .ZN(n36101) );
  NAND2_X1 U41168 ( .A1(n36098), .A2(n38201), .ZN(n36099) );
  NAND4_X1 U41169 ( .A1(n38570), .A2(n33062), .A3(n7759), .A4(n36099), .ZN(
        n36100) );
  AND4_X1 U41170 ( .A1(n36103), .A2(n36102), .A3(n36101), .A4(n36100), .ZN(
        n36110) );
  NAND2_X1 U41171 ( .A1(n36104), .A2(n38560), .ZN(n36109) );
  NAND2_X1 U41172 ( .A1(n36107), .A2(n36106), .ZN(n36108) );
  NOR2_X1 U41174 ( .A1(n38468), .A2(n36112), .ZN(n38115) );
  NAND2_X1 U41175 ( .A1(n38477), .A2(n38475), .ZN(n38465) );
  INV_X1 U41176 ( .A(n38465), .ZN(n38125) );
  AOI21_X1 U41177 ( .B1(n38115), .B2(n38467), .A(n38125), .ZN(n36113) );
  XNOR2_X1 U41178 ( .A(n38468), .B(n38475), .ZN(n36114) );
  NOR2_X1 U41179 ( .A1(n36115), .A2(n37420), .ZN(n38476) );
  NAND2_X1 U41180 ( .A1(n38476), .A2(n38478), .ZN(n36116) );
  INV_X1 U41181 ( .A(n38126), .ZN(n36119) );
  NAND2_X1 U41182 ( .A1(n38116), .A2(n38471), .ZN(n36118) );
  NAND2_X1 U41183 ( .A1(n36119), .A2(n36118), .ZN(n36120) );
  OAI21_X1 U41185 ( .B1(n38153), .B2(n38152), .A(n38166), .ZN(n36121) );
  OR2_X1 U41186 ( .A1(n36137), .A2(n38590), .ZN(n38155) );
  NAND2_X1 U41187 ( .A1(n37580), .A2(n38164), .ZN(n38157) );
  NOR2_X1 U41188 ( .A1(n36124), .A2(n38157), .ZN(n36125) );
  INV_X1 U41189 ( .A(n38158), .ZN(n36128) );
  NAND2_X1 U41190 ( .A1(n52104), .A2(n38599), .ZN(n36127) );
  NAND3_X1 U41191 ( .A1(n36127), .A2(n51429), .A3(n36133), .ZN(n36126) );
  OAI211_X1 U41192 ( .C1(n36128), .C2(n36127), .A(n36126), .B(n38585), .ZN(
        n36129) );
  OR2_X1 U41193 ( .A1(n37453), .A2(n38590), .ZN(n37572) );
  OAI21_X1 U41194 ( .B1(n37571), .B2(n37448), .A(n37572), .ZN(n36136) );
  NAND2_X1 U41195 ( .A1(n36132), .A2(n38152), .ZN(n36135) );
  NAND3_X1 U41196 ( .A1(n52104), .A2(n36133), .A3(n38585), .ZN(n37450) );
  OAI211_X1 U41197 ( .C1(n38152), .C2(n38585), .A(n38166), .B(n37450), .ZN(
        n36134) );
  OR2_X1 U41199 ( .A1(n38582), .A2(n38599), .ZN(n36138) );
  NOR2_X1 U41201 ( .A1(n39499), .A2(n51430), .ZN(n41209) );
  OAI21_X1 U41202 ( .B1(n38228), .B2(n5846), .A(n36141), .ZN(n36145) );
  OAI21_X1 U41203 ( .B1(n36142), .B2(n31355), .A(n35175), .ZN(n36143) );
  OAI21_X1 U41204 ( .B1(n36145), .B2(n36144), .A(n36143), .ZN(n36154) );
  INV_X1 U41205 ( .A(n38213), .ZN(n38548) );
  NOR2_X1 U41206 ( .A1(n38548), .A2(n38221), .ZN(n36146) );
  AOI22_X1 U41207 ( .A1(n36146), .A2(n38214), .B1(n38549), .B2(n38226), .ZN(
        n36153) );
  INV_X1 U41208 ( .A(n36147), .ZN(n36149) );
  NAND2_X1 U41209 ( .A1(n36149), .A2(n36148), .ZN(n36152) );
  OAI21_X1 U41210 ( .B1(n38226), .B2(n51738), .A(n35175), .ZN(n36150) );
  OAI211_X1 U41211 ( .C1(n38558), .C2(n38226), .A(n38553), .B(n36150), .ZN(
        n36151) );
  NAND3_X1 U41212 ( .A1(n51735), .A2(n38528), .A3(n38517), .ZN(n38523) );
  NAND3_X1 U41214 ( .A1(n51735), .A2(n38517), .A3(n37480), .ZN(n36165) );
  NAND3_X1 U41215 ( .A1(n51411), .A2(n51363), .A3(n37489), .ZN(n36156) );
  NAND2_X1 U41216 ( .A1(n37480), .A2(n36156), .ZN(n36157) );
  OAI21_X1 U41217 ( .B1(n51487), .B2(n38514), .A(n8315), .ZN(n36158) );
  NAND3_X1 U41218 ( .A1(n36158), .A2(n38518), .A3(n38517), .ZN(n36163) );
  NAND2_X1 U41219 ( .A1(n37442), .A2(n37489), .ZN(n36160) );
  OAI211_X1 U41220 ( .C1(n38517), .C2(n36161), .A(n36160), .B(n38515), .ZN(
        n36162) );
  INV_X1 U41221 ( .A(n36335), .ZN(n36343) );
  AOI22_X1 U41222 ( .A1(n36343), .A2(n36325), .B1(n36342), .B2(n38054), .ZN(
        n36173) );
  INV_X1 U41223 ( .A(n38067), .ZN(n36170) );
  NAND3_X1 U41224 ( .A1(n36170), .A2(n36325), .A3(n38050), .ZN(n38061) );
  AND2_X1 U41225 ( .A1(n5443), .A2(n38057), .ZN(n38137) );
  INV_X1 U41226 ( .A(n38137), .ZN(n36168) );
  NAND4_X1 U41227 ( .A1(n36169), .A2(n38132), .A3(n38050), .A4(n36168), .ZN(
        n36172) );
  NAND3_X1 U41228 ( .A1(n36170), .A2(n36330), .A3(n51522), .ZN(n36171) );
  NAND4_X1 U41229 ( .A1(n36173), .A2(n38061), .A3(n36172), .A4(n36171), .ZN(
        n36178) );
  INV_X1 U41230 ( .A(n36329), .ZN(n36174) );
  NAND2_X1 U41231 ( .A1(n36174), .A2(n36330), .ZN(n36176) );
  NAND2_X1 U41232 ( .A1(n611), .A2(n38050), .ZN(n36175) );
  AOI21_X1 U41233 ( .B1(n36176), .B2(n36175), .A(n38136), .ZN(n36177) );
  OR2_X2 U41234 ( .A1(n36178), .A2(n36177), .ZN(n41207) );
  OAI21_X1 U41235 ( .B1(n41209), .B2(n36179), .A(n41210), .ZN(n36185) );
  AND2_X1 U41236 ( .A1(n685), .A2(n40029), .ZN(n41196) );
  AND2_X1 U41238 ( .A1(n41206), .A2(n41205), .ZN(n36184) );
  NAND2_X1 U41239 ( .A1(n51052), .A2(n41207), .ZN(n40665) );
  AND2_X1 U41240 ( .A1(n41212), .A2(n40029), .ZN(n39505) );
  OAI211_X1 U41241 ( .C1(n39502), .C2(n7955), .A(n36180), .B(n39505), .ZN(
        n36183) );
  AND2_X1 U41242 ( .A1(n41195), .A2(n41212), .ZN(n40184) );
  OR2_X1 U41243 ( .A1(n41211), .A2(n40029), .ZN(n40033) );
  OAI21_X1 U41244 ( .B1(n40033), .B2(n41210), .A(n51052), .ZN(n36181) );
  AND2_X1 U41245 ( .A1(n51052), .A2(n41195), .ZN(n40028) );
  AOI22_X1 U41246 ( .A1(n40184), .A2(n36181), .B1(n40028), .B2(n5060), .ZN(
        n36182) );
  XNOR2_X1 U41247 ( .A(n51101), .B(n44240), .ZN(n36296) );
  INV_X1 U41248 ( .A(n37773), .ZN(n36187) );
  NAND3_X1 U41249 ( .A1(n36187), .A2(n36189), .A3(n36186), .ZN(n36194) );
  INV_X1 U41250 ( .A(n36188), .ZN(n36193) );
  OAI21_X1 U41251 ( .B1(n37782), .B2(n36189), .A(n37775), .ZN(n36190) );
  NAND2_X1 U41252 ( .A1(n36191), .A2(n36190), .ZN(n36192) );
  NAND4_X1 U41253 ( .A1(n36195), .A2(n36194), .A3(n36193), .A4(n36192), .ZN(
        n42055) );
  NAND2_X1 U41254 ( .A1(n39349), .A2(n39348), .ZN(n36198) );
  AOI21_X1 U41255 ( .B1(n36198), .B2(n36197), .A(n36196), .ZN(n42056) );
  INV_X1 U41256 ( .A(n36199), .ZN(n36201) );
  NAND2_X1 U41257 ( .A1(n39334), .A2(n39338), .ZN(n42057) );
  INV_X1 U41258 ( .A(n36202), .ZN(n36203) );
  NOR2_X1 U41259 ( .A1(n42057), .A2(n36203), .ZN(n36204) );
  NAND3_X1 U41260 ( .A1(n37809), .A2(n473), .A3(n37805), .ZN(n37801) );
  NAND2_X1 U41261 ( .A1(n39473), .A2(n37801), .ZN(n36206) );
  INV_X1 U41262 ( .A(n39484), .ZN(n36207) );
  NAND2_X1 U41263 ( .A1(n39481), .A2(n36215), .ZN(n38980) );
  NAND2_X1 U41265 ( .A1(n36211), .A2(n36210), .ZN(n36221) );
  INV_X1 U41266 ( .A(n39481), .ZN(n38982) );
  NAND2_X1 U41267 ( .A1(n39481), .A2(n36216), .ZN(n38971) );
  OAI211_X1 U41268 ( .C1(n36215), .C2(n36214), .A(n38981), .B(n39488), .ZN(
        n36219) );
  NAND4_X1 U41269 ( .A1(n39486), .A2(n36216), .A3(n37805), .A4(n39478), .ZN(
        n36217) );
  INV_X1 U41270 ( .A(n36223), .ZN(n36230) );
  INV_X1 U41271 ( .A(n37597), .ZN(n36224) );
  NOR2_X1 U41272 ( .A1(n36225), .A2(n36224), .ZN(n36226) );
  AOI22_X1 U41273 ( .A1(n690), .A2(n36227), .B1(n36226), .B2(n37598), .ZN(
        n36229) );
  OAI21_X1 U41274 ( .B1(n37597), .B2(n36231), .A(n37376), .ZN(n36235) );
  NAND3_X1 U41275 ( .A1(n36235), .A2(n36234), .A3(n37367), .ZN(n36236) );
  NAND2_X1 U41276 ( .A1(n36236), .A2(n37377), .ZN(n36237) );
  INV_X1 U41277 ( .A(n36242), .ZN(n36243) );
  OAI211_X1 U41278 ( .C1(n37507), .C2(n36244), .A(n36243), .B(n37501), .ZN(
        n36245) );
  INV_X1 U41279 ( .A(n37748), .ZN(n37511) );
  INV_X1 U41280 ( .A(n36247), .ZN(n37760) );
  NAND2_X1 U41281 ( .A1(n37747), .A2(n37757), .ZN(n36250) );
  AOI21_X1 U41282 ( .B1(n37757), .B2(n36251), .A(n36248), .ZN(n36249) );
  NAND4_X1 U41283 ( .A1(n36252), .A2(n37764), .A3(n37753), .A4(n36251), .ZN(
        n36253) );
  NAND2_X1 U41285 ( .A1(n39464), .A2(n51737), .ZN(n39445) );
  INV_X1 U41286 ( .A(n39445), .ZN(n36909) );
  NAND3_X1 U41287 ( .A1(n39034), .A2(n36909), .A3(n39453), .ZN(n36906) );
  NAND3_X1 U41288 ( .A1(n36907), .A2(n39448), .A3(n39032), .ZN(n36256) );
  AOI21_X1 U41291 ( .B1(n36909), .B2(n36259), .A(n39441), .ZN(n36262) );
  NAND2_X1 U41292 ( .A1(n36260), .A2(n34800), .ZN(n36261) );
  INV_X1 U41293 ( .A(n36903), .ZN(n39461) );
  MUX2_X1 U41294 ( .A(n36262), .B(n36261), .S(n39461), .Z(n36263) );
  NAND2_X1 U41295 ( .A1(n36265), .A2(n36272), .ZN(n36280) );
  OAI211_X1 U41296 ( .C1(n36269), .C2(n37544), .A(n36268), .B(n36267), .ZN(
        n36271) );
  INV_X1 U41297 ( .A(n37410), .ZN(n36270) );
  AOI21_X1 U41299 ( .B1(n37406), .B2(n37560), .A(n36272), .ZN(n36274) );
  OAI21_X1 U41300 ( .B1(n37547), .B2(n36274), .A(n34676), .ZN(n36275) );
  XNOR2_X1 U41302 ( .A(n37399), .B(n37543), .ZN(n36277) );
  NAND3_X1 U41303 ( .A1(n36277), .A2(n37406), .A3(n37558), .ZN(n36278) );
  AND2_X1 U41304 ( .A1(n42062), .A2(n480), .ZN(n36285) );
  INV_X1 U41305 ( .A(n480), .ZN(n41480) );
  NOR2_X1 U41306 ( .A1(n686), .A2(n42061), .ZN(n36282) );
  NOR2_X1 U41307 ( .A1(n36282), .A2(n42049), .ZN(n36283) );
  INV_X1 U41309 ( .A(n40294), .ZN(n39064) );
  NAND2_X1 U41310 ( .A1(n36282), .A2(n42441), .ZN(n40287) );
  INV_X1 U41311 ( .A(n36284), .ZN(n36289) );
  NAND2_X1 U41312 ( .A1(n686), .A2(n42061), .ZN(n42043) );
  AOI22_X1 U41313 ( .A1(n40051), .A2(n42043), .B1(n36286), .B2(n36285), .ZN(
        n36287) );
  XNOR2_X1 U41314 ( .A(n36291), .B(n2603), .ZN(n36292) );
  XNOR2_X1 U41315 ( .A(n36293), .B(n36292), .ZN(n36294) );
  XNOR2_X1 U41316 ( .A(n43954), .B(n36294), .ZN(n36295) );
  XNOR2_X1 U41317 ( .A(n36296), .B(n36295), .ZN(n36297) );
  XNOR2_X1 U41318 ( .A(n36298), .B(n36297), .ZN(n37353) );
  AOI22_X1 U41319 ( .A1(n38228), .A2(n5846), .B1(n38541), .B2(n51524), .ZN(
        n36304) );
  INV_X1 U41320 ( .A(n36300), .ZN(n36303) );
  NAND3_X1 U41321 ( .A1(n36305), .A2(n38544), .A3(n38549), .ZN(n36302) );
  OAI21_X1 U41322 ( .B1(n38550), .B2(n31355), .A(n38217), .ZN(n36301) );
  OAI211_X1 U41323 ( .C1(n36304), .C2(n36303), .A(n36302), .B(n36301), .ZN(
        n36311) );
  NAND2_X1 U41324 ( .A1(n36307), .A2(n51524), .ZN(n36308) );
  INV_X1 U41325 ( .A(n36320), .ZN(n36314) );
  OAI22_X1 U41326 ( .A1(n36314), .A2(n50984), .B1(n36313), .B2(n36312), .ZN(
        n36316) );
  INV_X1 U41327 ( .A(n38086), .ZN(n38083) );
  NAND2_X1 U41328 ( .A1(n38083), .A2(n38073), .ZN(n36315) );
  MUX2_X1 U41329 ( .A(n36316), .B(n36315), .S(n38082), .Z(n36324) );
  NAND2_X1 U41330 ( .A1(n36318), .A2(n36317), .ZN(n36323) );
  INV_X1 U41331 ( .A(n36319), .ZN(n36633) );
  NAND2_X1 U41332 ( .A1(n36321), .A2(n38094), .ZN(n36322) );
  INV_X1 U41333 ( .A(n38052), .ZN(n36327) );
  OAI21_X1 U41334 ( .B1(n36327), .B2(n36326), .A(n38058), .ZN(n36334) );
  NAND3_X1 U41335 ( .A1(n38131), .A2(n38148), .A3(n38142), .ZN(n36333) );
  OAI21_X1 U41336 ( .B1(n38050), .B2(n38142), .A(n38145), .ZN(n36331) );
  NAND2_X1 U41337 ( .A1(n36331), .A2(n36330), .ZN(n36332) );
  OAI211_X1 U41338 ( .C1(n38057), .C2(n38135), .A(n36338), .B(n36337), .ZN(
        n36339) );
  NAND4_X1 U41339 ( .A1(n36341), .A2(n38142), .A3(n38137), .A4(n38145), .ZN(
        n36347) );
  NAND3_X1 U41340 ( .A1(n38058), .A2(n36342), .A3(n38050), .ZN(n36346) );
  NAND2_X1 U41341 ( .A1(n36344), .A2(n36343), .ZN(n36345) );
  MUX2_X1 U41342 ( .A(n37991), .B(n36525), .S(n37990), .Z(n36350) );
  NOR2_X1 U41343 ( .A1(n36350), .A2(n36533), .ZN(n36357) );
  INV_X1 U41344 ( .A(n36524), .ZN(n36532) );
  OAI21_X1 U41345 ( .B1(n36353), .B2(n36532), .A(n36529), .ZN(n36352) );
  NAND2_X1 U41346 ( .A1(n36352), .A2(n37991), .ZN(n36356) );
  INV_X1 U41347 ( .A(n36522), .ZN(n36354) );
  NAND4_X1 U41348 ( .A1(n37977), .A2(n36354), .A3(n36524), .A4(n36353), .ZN(
        n36355) );
  INV_X1 U41349 ( .A(n36358), .ZN(n36363) );
  NAND3_X1 U41350 ( .A1(n38001), .A2(n36359), .A3(n38015), .ZN(n36360) );
  OAI211_X1 U41351 ( .C1(n36363), .C2(n36362), .A(n36361), .B(n36360), .ZN(
        n36368) );
  MUX2_X1 U41352 ( .A(n38189), .B(n38177), .S(n38005), .Z(n36367) );
  INV_X1 U41353 ( .A(n38190), .ZN(n36365) );
  NAND3_X1 U41354 ( .A1(n38173), .A2(n38189), .A3(n38012), .ZN(n36366) );
  NAND2_X1 U41355 ( .A1(n39768), .A2(n39160), .ZN(n41430) );
  OAI22_X1 U41356 ( .A1(n36373), .A2(n36376), .B1(n38029), .B2(n36372), .ZN(
        n36374) );
  NAND3_X1 U41357 ( .A1(n36375), .A2(n38043), .A3(n38029), .ZN(n36378) );
  INV_X1 U41358 ( .A(n36382), .ZN(n36387) );
  NOR2_X1 U41359 ( .A1(n36383), .A2(n38043), .ZN(n36385) );
  NOR2_X1 U41360 ( .A1(n36385), .A2(n36384), .ZN(n36386) );
  NAND2_X1 U41361 ( .A1(n39767), .A2(n5983), .ZN(n41447) );
  NAND2_X1 U41362 ( .A1(n40644), .A2(n41447), .ZN(n36391) );
  NAND2_X1 U41363 ( .A1(n39767), .A2(n41446), .ZN(n41434) );
  NOR2_X1 U41364 ( .A1(n41434), .A2(n40655), .ZN(n36389) );
  AND2_X1 U41365 ( .A1(n39768), .A2(n40651), .ZN(n38912) );
  MUX2_X1 U41366 ( .A(n40652), .B(n8759), .S(n40655), .Z(n36392) );
  NAND3_X1 U41367 ( .A1(n36398), .A2(n36397), .A3(n36396), .ZN(n36399) );
  AND2_X1 U41368 ( .A1(n36400), .A2(n36399), .ZN(n36419) );
  INV_X1 U41369 ( .A(n36401), .ZN(n37638) );
  NAND3_X1 U41370 ( .A1(n36404), .A2(n36403), .A3(n36402), .ZN(n36407) );
  NAND2_X1 U41371 ( .A1(n36407), .A2(n36406), .ZN(n36409) );
  NAND4_X1 U41372 ( .A1(n37644), .A2(n37648), .A3(n36410), .A4(n37649), .ZN(
        n36417) );
  INV_X1 U41373 ( .A(n36411), .ZN(n36412) );
  OAI21_X1 U41374 ( .B1(n5588), .B2(n5590), .A(n36412), .ZN(n36413) );
  OAI21_X1 U41375 ( .B1(n37640), .B2(n37646), .A(n36413), .ZN(n36415) );
  NOR2_X1 U41377 ( .A1(n36610), .A2(n51015), .ZN(n36615) );
  OAI211_X1 U41378 ( .C1(n36426), .C2(n51716), .A(n36421), .B(n36420), .ZN(
        n36423) );
  NAND2_X1 U41379 ( .A1(n36618), .A2(n51717), .ZN(n36422) );
  OAI211_X1 U41380 ( .C1(n36424), .C2(n36615), .A(n36423), .B(n36422), .ZN(
        n36434) );
  OAI21_X1 U41381 ( .B1(n36426), .B2(n36606), .A(n36425), .ZN(n36432) );
  INV_X1 U41382 ( .A(n36610), .ZN(n36431) );
  NOR2_X1 U41383 ( .A1(n38279), .A2(n38276), .ZN(n36437) );
  NAND2_X1 U41384 ( .A1(n38286), .A2(n36437), .ZN(n36444) );
  INV_X1 U41385 ( .A(n37617), .ZN(n38289) );
  AOI22_X1 U41386 ( .A1(n37627), .A2(n38289), .B1(n38292), .B2(n36436), .ZN(
        n36443) );
  NOR2_X1 U41387 ( .A1(n51339), .A2(n37624), .ZN(n36438) );
  AOI22_X1 U41388 ( .A1(n37627), .A2(n36438), .B1(n2120), .B2(n37629), .ZN(
        n36442) );
  NAND2_X1 U41389 ( .A1(n36440), .A2(n36439), .ZN(n36441) );
  NAND4_X1 U41390 ( .A1(n36444), .A2(n36443), .A3(n36442), .A4(n36441), .ZN(
        n36447) );
  NAND2_X1 U41391 ( .A1(n38276), .A2(n38275), .ZN(n37619) );
  NOR2_X1 U41392 ( .A1(n36445), .A2(n37619), .ZN(n36446) );
  NOR2_X1 U41393 ( .A1(n36449), .A2(n36592), .ZN(n36583) );
  OAI21_X1 U41394 ( .B1(n1692), .B2(n36451), .A(n36450), .ZN(n36453) );
  NOR2_X1 U41396 ( .A1(n36454), .A2(n36459), .ZN(n36455) );
  NOR2_X1 U41397 ( .A1(n36456), .A2(n36455), .ZN(n36465) );
  OAI21_X1 U41398 ( .B1(n36459), .B2(n36458), .A(n36457), .ZN(n36460) );
  OAI21_X1 U41399 ( .B1(n36461), .B2(n36460), .A(n36585), .ZN(n36464) );
  INV_X1 U41400 ( .A(n36462), .ZN(n36597) );
  NAND3_X1 U41401 ( .A1(n36600), .A2(n36591), .A3(n36597), .ZN(n36463) );
  OAI21_X1 U41403 ( .B1(n37664), .B2(n6614), .A(n37663), .ZN(n36467) );
  AOI22_X1 U41404 ( .A1(n37669), .A2(n37665), .B1(n38322), .B2(n38337), .ZN(
        n36469) );
  NAND2_X1 U41405 ( .A1(n38838), .A2(n52095), .ZN(n38830) );
  AND2_X1 U41406 ( .A1(n36470), .A2(n39938), .ZN(n36503) );
  AND2_X1 U41408 ( .A1(n63), .A2(n458), .ZN(n36484) );
  NAND3_X1 U41409 ( .A1(n36484), .A2(n36475), .A3(n36473), .ZN(n36477) );
  NAND3_X1 U41410 ( .A1(n36558), .A2(n36475), .A3(n36474), .ZN(n36476) );
  OAI21_X1 U41411 ( .B1(n36482), .B2(n36481), .A(n36480), .ZN(n36483) );
  INV_X1 U41412 ( .A(n36483), .ZN(n36501) );
  NAND2_X1 U41413 ( .A1(n36484), .A2(n36567), .ZN(n36487) );
  NAND4_X1 U41414 ( .A1(n36490), .A2(n36488), .A3(n63), .A4(n36567), .ZN(
        n36486) );
  AND2_X1 U41415 ( .A1(n36493), .A2(n36492), .ZN(n36496) );
  NOR2_X1 U41416 ( .A1(n36495), .A2(n36494), .ZN(n36497) );
  OAI21_X1 U41417 ( .B1(n36498), .B2(n36497), .A(n36496), .ZN(n36499) );
  OAI21_X1 U41418 ( .B1(n36504), .B2(n36503), .A(n39943), .ZN(n36515) );
  NAND2_X1 U41419 ( .A1(n575), .A2(n39938), .ZN(n36506) );
  OAI21_X1 U41420 ( .B1(n39112), .B2(n36506), .A(n36505), .ZN(n36507) );
  NAND2_X1 U41421 ( .A1(n36507), .A2(n39937), .ZN(n36514) );
  OAI211_X1 U41422 ( .C1(n52095), .C2(n39938), .A(n36508), .B(n52073), .ZN(
        n36513) );
  NAND2_X1 U41423 ( .A1(n39955), .A2(n39754), .ZN(n39761) );
  INV_X1 U41424 ( .A(n39761), .ZN(n36511) );
  NAND2_X1 U41425 ( .A1(n39751), .A2(n52094), .ZN(n39953) );
  INV_X1 U41426 ( .A(n39953), .ZN(n36510) );
  NAND3_X1 U41427 ( .A1(n36511), .A2(n36510), .A3(n39943), .ZN(n36512) );
  XNOR2_X1 U41428 ( .A(n43950), .B(n52096), .ZN(n36664) );
  NAND2_X1 U41429 ( .A1(n36535), .A2(n36524), .ZN(n36523) );
  NAND2_X1 U41430 ( .A1(n36529), .A2(n594), .ZN(n37986) );
  AOI21_X1 U41431 ( .B1(n37977), .B2(n36530), .A(n37986), .ZN(n36538) );
  OAI21_X1 U41432 ( .B1(n36532), .B2(n37987), .A(n36531), .ZN(n36537) );
  NAND3_X1 U41433 ( .A1(n36542), .A2(n36541), .A3(n6218), .ZN(n36543) );
  NAND3_X1 U41435 ( .A1(n36548), .A2(n36547), .A3(n37969), .ZN(n36556) );
  OAI211_X1 U41436 ( .C1(n37957), .C2(n7851), .A(n36550), .B(n36549), .ZN(
        n36551) );
  NAND2_X1 U41437 ( .A1(n36551), .A2(n37963), .ZN(n36555) );
  NAND3_X1 U41438 ( .A1(n36553), .A2(n6218), .A3(n36552), .ZN(n36554) );
  INV_X1 U41439 ( .A(n39682), .ZN(n39683) );
  NAND2_X1 U41440 ( .A1(n36558), .A2(n36557), .ZN(n36564) );
  AOI22_X1 U41441 ( .A1(n36562), .A2(n36561), .B1(n36560), .B2(n36559), .ZN(
        n36563) );
  MUX2_X1 U41442 ( .A(n36564), .B(n36563), .S(n36567), .Z(n36579) );
  NOR2_X1 U41443 ( .A1(n36566), .A2(n36565), .ZN(n36578) );
  MUX2_X1 U41444 ( .A(n36569), .B(n36568), .S(n36567), .Z(n36577) );
  INV_X1 U41445 ( .A(n36570), .ZN(n36573) );
  NAND4_X1 U41446 ( .A1(n36573), .A2(n36572), .A3(n36571), .A4(n458), .ZN(
        n36574) );
  NAND2_X1 U41447 ( .A1(n39683), .A2(n39674), .ZN(n36663) );
  INV_X1 U41448 ( .A(n36580), .ZN(n36582) );
  INV_X1 U41450 ( .A(n36584), .ZN(n36588) );
  NOR2_X1 U41451 ( .A1(n36586), .A2(n36585), .ZN(n36587) );
  NOR2_X1 U41453 ( .A1(n36590), .A2(n36589), .ZN(n36596) );
  NAND2_X1 U41454 ( .A1(n36593), .A2(n36592), .ZN(n36594) );
  OAI211_X1 U41455 ( .C1(n36597), .C2(n36596), .A(n36595), .B(n36594), .ZN(
        n36599) );
  INV_X1 U41456 ( .A(n36603), .ZN(n36608) );
  NAND2_X1 U41457 ( .A1(n36606), .A2(n36604), .ZN(n36605) );
  OAI211_X1 U41458 ( .C1(n698), .C2(n36606), .A(n36605), .B(n36618), .ZN(
        n36607) );
  AND2_X1 U41459 ( .A1(n36608), .A2(n36607), .ZN(n36626) );
  AND2_X1 U41460 ( .A1(n36610), .A2(n36609), .ZN(n36613) );
  AOI22_X1 U41462 ( .A1(n36615), .A2(n36614), .B1(n36613), .B2(n36612), .ZN(
        n36625) );
  NAND2_X1 U41463 ( .A1(n36617), .A2(n36616), .ZN(n36620) );
  INV_X1 U41464 ( .A(n36618), .ZN(n36619) );
  NAND4_X1 U41465 ( .A1(n36622), .A2(n51716), .A3(n36620), .A4(n36619), .ZN(
        n36624) );
  NAND2_X1 U41466 ( .A1(n40684), .A2(n40676), .ZN(n39680) );
  MUX2_X1 U41468 ( .A(n39680), .B(n39931), .S(n39929), .Z(n36662) );
  NAND2_X1 U41469 ( .A1(n36627), .A2(n36632), .ZN(n38071) );
  NAND2_X1 U41470 ( .A1(n38071), .A2(n36629), .ZN(n36630) );
  AOI22_X1 U41471 ( .A1(n36635), .A2(n36634), .B1(n50984), .B2(n36633), .ZN(
        n36636) );
  NAND2_X1 U41472 ( .A1(n36637), .A2(n36636), .ZN(n36648) );
  NAND2_X1 U41473 ( .A1(n36640), .A2(n36639), .ZN(n36645) );
  INV_X1 U41474 ( .A(n36641), .ZN(n36643) );
  OAI21_X1 U41475 ( .B1(n36643), .B2(n38082), .A(n36642), .ZN(n36644) );
  NOR2_X1 U41476 ( .A1(n39674), .A2(n40683), .ZN(n40693) );
  AND2_X1 U41477 ( .A1(n51022), .A2(n40689), .ZN(n39684) );
  NAND3_X1 U41478 ( .A1(n40693), .A2(n39684), .A3(n40684), .ZN(n36657) );
  AND2_X1 U41479 ( .A1(n39674), .A2(n40683), .ZN(n40677) );
  OAI211_X1 U41482 ( .C1(n39673), .C2(n36649), .A(n36653), .B(n40684), .ZN(
        n36654) );
  NAND2_X1 U41483 ( .A1(n40677), .A2(n36654), .ZN(n36656) );
  NAND2_X1 U41484 ( .A1(n40685), .A2(n40684), .ZN(n38415) );
  AND2_X1 U41485 ( .A1(n40683), .A2(n40689), .ZN(n40682) );
  NAND2_X1 U41486 ( .A1(n38415), .A2(n40682), .ZN(n36655) );
  INV_X1 U41487 ( .A(n40684), .ZN(n40692) );
  NAND2_X1 U41488 ( .A1(n40692), .A2(n38401), .ZN(n38409) );
  NAND2_X1 U41489 ( .A1(n38409), .A2(n40675), .ZN(n36659) );
  NAND3_X1 U41490 ( .A1(n38404), .A2(n40685), .A3(n39929), .ZN(n36658) );
  INV_X1 U41491 ( .A(n40677), .ZN(n39672) );
  NAND4_X1 U41492 ( .A1(n36659), .A2(n39673), .A3(n36658), .A4(n39672), .ZN(
        n36660) );
  XNOR2_X1 U41493 ( .A(n36664), .B(n51099), .ZN(n37352) );
  INV_X1 U41494 ( .A(n36665), .ZN(n36666) );
  XNOR2_X1 U41495 ( .A(n36667), .B(n36666), .ZN(n36668) );
  XNOR2_X1 U41496 ( .A(n36847), .B(n36668), .ZN(n36670) );
  XNOR2_X1 U41497 ( .A(n36670), .B(n52148), .ZN(n36676) );
  XNOR2_X1 U41498 ( .A(n36672), .B(n36671), .ZN(n36673) );
  XNOR2_X1 U41499 ( .A(n36673), .B(n36674), .ZN(n36675) );
  XNOR2_X1 U41500 ( .A(n36675), .B(n36676), .ZN(n36678) );
  XNOR2_X1 U41501 ( .A(n31573), .B(n36681), .ZN(n36952) );
  XNOR2_X1 U41502 ( .A(n36952), .B(n37039), .ZN(n36689) );
  XNOR2_X1 U41503 ( .A(n36855), .B(n36940), .ZN(n36687) );
  XNOR2_X1 U41504 ( .A(n36683), .B(n36682), .ZN(n36684) );
  XNOR2_X1 U41505 ( .A(n36685), .B(n36684), .ZN(n36686) );
  XNOR2_X1 U41506 ( .A(n36687), .B(n36686), .ZN(n36688) );
  XNOR2_X1 U41507 ( .A(n36689), .B(n36688), .ZN(n36690) );
  XNOR2_X1 U41508 ( .A(n36690), .B(n2322), .ZN(n36696) );
  INV_X1 U41509 ( .A(n36691), .ZN(n36694) );
  XNOR2_X1 U41510 ( .A(n36856), .B(n36692), .ZN(n36693) );
  XNOR2_X1 U41511 ( .A(n36694), .B(n36693), .ZN(n36695) );
  INV_X1 U41512 ( .A(n36697), .ZN(n36699) );
  XNOR2_X1 U41513 ( .A(n36699), .B(n36698), .ZN(n36700) );
  XNOR2_X1 U41514 ( .A(n36704), .B(n36705), .ZN(n36706) );
  XNOR2_X1 U41515 ( .A(n36706), .B(n37296), .ZN(n36712) );
  INV_X1 U41516 ( .A(n36707), .ZN(n36708) );
  XNOR2_X1 U41517 ( .A(n36708), .B(n37089), .ZN(n36710) );
  XNOR2_X1 U41518 ( .A(n36710), .B(n36709), .ZN(n36711) );
  XNOR2_X1 U41519 ( .A(n36712), .B(n36711), .ZN(n36716) );
  XNOR2_X1 U41520 ( .A(n36714), .B(n36713), .ZN(n36715) );
  INV_X1 U41522 ( .A(n39007), .ZN(n39268) );
  NAND2_X1 U41523 ( .A1(n39270), .A2(n39268), .ZN(n39015) );
  INV_X1 U41524 ( .A(n39269), .ZN(n39265) );
  XNOR2_X1 U41525 ( .A(n36718), .B(n36717), .ZN(n36719) );
  XNOR2_X1 U41526 ( .A(n36720), .B(n36719), .ZN(n36721) );
  XNOR2_X1 U41527 ( .A(n36722), .B(n36721), .ZN(n36725) );
  INV_X1 U41528 ( .A(n36723), .ZN(n36724) );
  XNOR2_X1 U41529 ( .A(n36725), .B(n36724), .ZN(n36726) );
  XNOR2_X1 U41530 ( .A(n36962), .B(n36726), .ZN(n36729) );
  INV_X1 U41531 ( .A(n36727), .ZN(n36728) );
  XNOR2_X1 U41532 ( .A(n36728), .B(n36729), .ZN(n36736) );
  INV_X1 U41533 ( .A(n36730), .ZN(n36734) );
  INV_X1 U41534 ( .A(n36731), .ZN(n36732) );
  XNOR2_X1 U41535 ( .A(n36971), .B(n36732), .ZN(n36733) );
  XNOR2_X1 U41536 ( .A(n36734), .B(n36733), .ZN(n36735) );
  XNOR2_X1 U41537 ( .A(n36736), .B(n36735), .ZN(n36771) );
  INV_X1 U41538 ( .A(n39264), .ZN(n37942) );
  XNOR2_X1 U41539 ( .A(n36737), .B(n4451), .ZN(n36826) );
  XNOR2_X1 U41540 ( .A(n36739), .B(n36738), .ZN(n36740) );
  XNOR2_X1 U41541 ( .A(n36826), .B(n36740), .ZN(n36743) );
  INV_X1 U41542 ( .A(n36741), .ZN(n36742) );
  XNOR2_X1 U41543 ( .A(n36743), .B(n36742), .ZN(n36744) );
  XNOR2_X1 U41544 ( .A(n37304), .B(n36744), .ZN(n36745) );
  XNOR2_X1 U41545 ( .A(n36746), .B(n36745), .ZN(n36750) );
  XNOR2_X1 U41546 ( .A(n36748), .B(n36747), .ZN(n36749) );
  XNOR2_X1 U41547 ( .A(n36750), .B(n36749), .ZN(n36752) );
  XNOR2_X1 U41548 ( .A(n36751), .B(n36752), .ZN(n36753) );
  XNOR2_X1 U41549 ( .A(n36756), .B(n2605), .ZN(n36757) );
  XNOR2_X1 U41550 ( .A(n36758), .B(n36757), .ZN(n36759) );
  XNOR2_X1 U41551 ( .A(n36761), .B(n36760), .ZN(n36762) );
  XNOR2_X1 U41552 ( .A(n36763), .B(n36762), .ZN(n36768) );
  XNOR2_X1 U41553 ( .A(n36764), .B(n37318), .ZN(n36765) );
  XNOR2_X1 U41554 ( .A(n36766), .B(n36765), .ZN(n36767) );
  XNOR2_X1 U41555 ( .A(n36767), .B(n36881), .ZN(n37129) );
  XNOR2_X1 U41556 ( .A(n36768), .B(n37129), .ZN(n36769) );
  INV_X1 U41557 ( .A(n39284), .ZN(n36770) );
  AND2_X1 U41558 ( .A1(n39262), .A2(n39273), .ZN(n37202) );
  AND2_X1 U41559 ( .A1(n8480), .A2(n39019), .ZN(n39280) );
  OAI21_X1 U41560 ( .B1(n39285), .B2(n37202), .A(n39280), .ZN(n36773) );
  AOI21_X1 U41561 ( .B1(n36774), .B2(n36773), .A(n551), .ZN(n36777) );
  NAND2_X1 U41562 ( .A1(n39266), .A2(n39264), .ZN(n39020) );
  OAI21_X1 U41563 ( .B1(n39020), .B2(n39263), .A(n36775), .ZN(n36776) );
  INV_X1 U41564 ( .A(n39285), .ZN(n39012) );
  NAND2_X1 U41565 ( .A1(n39262), .A2(n36781), .ZN(n36778) );
  NOR2_X1 U41566 ( .A1(n39282), .A2(n36781), .ZN(n36782) );
  MUX2_X1 U41567 ( .A(n39265), .B(n36779), .S(n8429), .Z(n36783) );
  AND2_X1 U41568 ( .A1(n39014), .A2(n39268), .ZN(n39274) );
  OAI21_X1 U41569 ( .B1(n36783), .B2(n551), .A(n39274), .ZN(n36784) );
  XNOR2_X1 U41570 ( .A(n36788), .B(n36787), .ZN(n36799) );
  INV_X1 U41571 ( .A(n42215), .ZN(n36790) );
  XNOR2_X1 U41572 ( .A(n36790), .B(n36789), .ZN(n36791) );
  XNOR2_X1 U41573 ( .A(n36792), .B(n36791), .ZN(n36794) );
  XNOR2_X1 U41574 ( .A(n36794), .B(n36793), .ZN(n36795) );
  XNOR2_X1 U41575 ( .A(n36795), .B(n37294), .ZN(n36797) );
  XNOR2_X1 U41576 ( .A(n36797), .B(n36796), .ZN(n36798) );
  INV_X1 U41577 ( .A(n39410), .ZN(n38946) );
  XNOR2_X1 U41578 ( .A(n36801), .B(n36800), .ZN(n36816) );
  XNOR2_X1 U41579 ( .A(n36803), .B(n36802), .ZN(n36804) );
  XNOR2_X1 U41580 ( .A(n36805), .B(n36804), .ZN(n36806) );
  XNOR2_X1 U41581 ( .A(n36807), .B(n36806), .ZN(n36810) );
  INV_X1 U41582 ( .A(n36808), .ZN(n36809) );
  XNOR2_X1 U41583 ( .A(n36809), .B(n36810), .ZN(n36814) );
  XNOR2_X1 U41584 ( .A(n36812), .B(n36811), .ZN(n37278) );
  XNOR2_X1 U41585 ( .A(n2598), .B(n37278), .ZN(n36813) );
  XOR2_X1 U41586 ( .A(n36814), .B(n36813), .Z(n36815) );
  XNOR2_X1 U41589 ( .A(n36822), .B(n36821), .ZN(n36834) );
  XNOR2_X1 U41590 ( .A(n36824), .B(n36823), .ZN(n45441) );
  XNOR2_X1 U41591 ( .A(n45104), .B(n37138), .ZN(n36825) );
  XNOR2_X1 U41592 ( .A(n36826), .B(n36825), .ZN(n36827) );
  XNOR2_X1 U41593 ( .A(n45441), .B(n36827), .ZN(n36828) );
  XNOR2_X1 U41594 ( .A(n36829), .B(n36828), .ZN(n36830) );
  XNOR2_X1 U41595 ( .A(n36830), .B(n33145), .ZN(n36831) );
  XNOR2_X1 U41596 ( .A(n50983), .B(n36831), .ZN(n36833) );
  MUX2_X1 U41597 ( .A(n39423), .B(n39410), .S(n38953), .Z(n36835) );
  NOR2_X1 U41598 ( .A1(n36835), .A2(n39430), .ZN(n36894) );
  INV_X1 U41599 ( .A(n36836), .ZN(n36839) );
  XNOR2_X1 U41600 ( .A(n36837), .B(n42889), .ZN(n36838) );
  XNOR2_X1 U41601 ( .A(n36839), .B(n36838), .ZN(n36840) );
  XNOR2_X1 U41602 ( .A(n37062), .B(n36840), .ZN(n36842) );
  XNOR2_X1 U41603 ( .A(n36842), .B(n52138), .ZN(n36843) );
  XNOR2_X1 U41604 ( .A(n52117), .B(n37067), .ZN(n36849) );
  XNOR2_X1 U41605 ( .A(n36849), .B(n37243), .ZN(n36850) );
  XNOR2_X1 U41606 ( .A(n36851), .B(n36850), .ZN(n36937) );
  INV_X1 U41607 ( .A(n36937), .ZN(n36852) );
  XNOR2_X1 U41608 ( .A(n36855), .B(n36854), .ZN(n37264) );
  XNOR2_X1 U41609 ( .A(n36858), .B(n36857), .ZN(n37051) );
  INV_X1 U41610 ( .A(n36859), .ZN(n36860) );
  XNOR2_X1 U41611 ( .A(n36860), .B(n4529), .ZN(n36862) );
  XNOR2_X1 U41612 ( .A(n36862), .B(n36861), .ZN(n36863) );
  XNOR2_X1 U41613 ( .A(n36940), .B(n36863), .ZN(n36864) );
  XNOR2_X1 U41614 ( .A(n36951), .B(n36864), .ZN(n36866) );
  XNOR2_X1 U41615 ( .A(n36865), .B(n36866), .ZN(n36867) );
  INV_X1 U41616 ( .A(n36868), .ZN(n36871) );
  XNOR2_X1 U41617 ( .A(n36869), .B(n704), .ZN(n36870) );
  XNOR2_X1 U41618 ( .A(n36871), .B(n36870), .ZN(n36872) );
  XNOR2_X1 U41619 ( .A(n36875), .B(n36874), .ZN(n36884) );
  XNOR2_X1 U41620 ( .A(n36876), .B(n4578), .ZN(n36877) );
  XNOR2_X1 U41621 ( .A(n36878), .B(n36877), .ZN(n36879) );
  XNOR2_X1 U41622 ( .A(n36880), .B(n36879), .ZN(n36882) );
  XNOR2_X1 U41623 ( .A(n36882), .B(n460), .ZN(n36883) );
  XNOR2_X1 U41624 ( .A(n36884), .B(n36883), .ZN(n36886) );
  AND2_X1 U41625 ( .A1(n38937), .A2(n38940), .ZN(n39211) );
  INV_X1 U41626 ( .A(n37907), .ZN(n38938) );
  NAND3_X1 U41627 ( .A1(n39207), .A2(n38938), .A3(n38940), .ZN(n36891) );
  NAND2_X1 U41628 ( .A1(n38953), .A2(n39430), .ZN(n36890) );
  INV_X1 U41629 ( .A(n38940), .ZN(n38950) );
  NOR2_X1 U41630 ( .A1(n36895), .A2(n39464), .ZN(n39030) );
  INV_X1 U41631 ( .A(n39030), .ZN(n36897) );
  NAND2_X1 U41632 ( .A1(n36897), .A2(n36896), .ZN(n36900) );
  NAND2_X1 U41633 ( .A1(n39444), .A2(n36901), .ZN(n36899) );
  NAND3_X1 U41634 ( .A1(n36900), .A2(n39453), .A3(n36899), .ZN(n36916) );
  NAND2_X1 U41635 ( .A1(n467), .A2(n36901), .ZN(n39031) );
  INV_X1 U41636 ( .A(n39031), .ZN(n36902) );
  NAND3_X1 U41637 ( .A1(n36902), .A2(n39438), .A3(n39036), .ZN(n36905) );
  NAND2_X1 U41638 ( .A1(n36903), .A2(n39032), .ZN(n36904) );
  AND3_X1 U41639 ( .A1(n36906), .A2(n36905), .A3(n36904), .ZN(n36915) );
  NAND3_X1 U41640 ( .A1(n36907), .A2(n39026), .A3(n39453), .ZN(n36911) );
  NAND2_X1 U41641 ( .A1(n34800), .A2(n39438), .ZN(n36908) );
  NAND4_X1 U41642 ( .A1(n39461), .A2(n36909), .A3(n39036), .A4(n36908), .ZN(
        n36910) );
  AND2_X1 U41643 ( .A1(n36911), .A2(n36910), .ZN(n36914) );
  INV_X1 U41644 ( .A(n36912), .ZN(n39454) );
  NAND2_X1 U41645 ( .A1(n37719), .A2(n39454), .ZN(n36913) );
  NAND2_X1 U41646 ( .A1(n37740), .A2(n39395), .ZN(n37735) );
  XNOR2_X1 U41647 ( .A(n3735), .B(n38998), .ZN(n36919) );
  NOR2_X1 U41648 ( .A1(n39003), .A2(n37731), .ZN(n36918) );
  AOI22_X1 U41649 ( .A1(n37890), .A2(n37739), .B1(n36919), .B2(n36918), .ZN(
        n36925) );
  NAND2_X1 U41650 ( .A1(n39003), .A2(n37885), .ZN(n36920) );
  NAND3_X1 U41651 ( .A1(n3577), .A2(n38998), .A3(n51474), .ZN(n39396) );
  OAI21_X1 U41652 ( .B1(n37894), .B2(n36920), .A(n39396), .ZN(n36921) );
  INV_X1 U41653 ( .A(n36921), .ZN(n36924) );
  INV_X1 U41654 ( .A(n37894), .ZN(n39394) );
  NAND2_X1 U41655 ( .A1(n39399), .A2(n38999), .ZN(n36922) );
  OAI211_X1 U41656 ( .C1(n39394), .C2(n39400), .A(n39402), .B(n36922), .ZN(
        n36923) );
  XOR2_X1 U41657 ( .A(n48814), .B(n5016), .Z(n36926) );
  XNOR2_X1 U41658 ( .A(n41949), .B(n36926), .ZN(n36927) );
  XNOR2_X1 U41659 ( .A(n36928), .B(n36927), .ZN(n36929) );
  XNOR2_X1 U41660 ( .A(n36932), .B(n33195), .ZN(n36933) );
  XNOR2_X1 U41661 ( .A(n36935), .B(n36936), .ZN(n36938) );
  XNOR2_X1 U41662 ( .A(n36940), .B(n36939), .ZN(n36950) );
  XNOR2_X1 U41663 ( .A(n36941), .B(n2203), .ZN(n36942) );
  XNOR2_X1 U41664 ( .A(n36943), .B(n36942), .ZN(n36944) );
  XNOR2_X1 U41665 ( .A(n36945), .B(n36944), .ZN(n36947) );
  XNOR2_X1 U41666 ( .A(n36947), .B(n36946), .ZN(n36948) );
  XNOR2_X1 U41667 ( .A(n37045), .B(n36948), .ZN(n36949) );
  XNOR2_X1 U41668 ( .A(n36954), .B(n36953), .ZN(n36958) );
  XNOR2_X1 U41669 ( .A(n36956), .B(n36955), .ZN(n36957) );
  XNOR2_X1 U41670 ( .A(n36958), .B(n36957), .ZN(n39195) );
  INV_X1 U41671 ( .A(n36959), .ZN(n36961) );
  XNOR2_X1 U41672 ( .A(n36962), .B(n36963), .ZN(n36974) );
  XNOR2_X1 U41673 ( .A(n36964), .B(n4636), .ZN(n36965) );
  XNOR2_X1 U41674 ( .A(n36966), .B(n36965), .ZN(n36967) );
  XNOR2_X1 U41675 ( .A(n36968), .B(n36967), .ZN(n36969) );
  XNOR2_X1 U41676 ( .A(n33702), .B(n36969), .ZN(n36970) );
  INV_X1 U41677 ( .A(n36971), .ZN(n36972) );
  INV_X1 U41678 ( .A(n36975), .ZN(n37286) );
  XNOR2_X1 U41679 ( .A(n36977), .B(n36976), .ZN(n36978) );
  XNOR2_X1 U41680 ( .A(n36979), .B(n36978), .ZN(n36980) );
  XNOR2_X1 U41681 ( .A(n36981), .B(n36980), .ZN(n36982) );
  XNOR2_X1 U41682 ( .A(n36983), .B(n36982), .ZN(n36984) );
  XNOR2_X1 U41683 ( .A(n37078), .B(n36984), .ZN(n36985) );
  XNOR2_X1 U41684 ( .A(n36985), .B(n37286), .ZN(n36990) );
  XNOR2_X1 U41685 ( .A(n36988), .B(n36987), .ZN(n36989) );
  NAND2_X1 U41686 ( .A1(n37881), .A2(n37790), .ZN(n37882) );
  NOR2_X1 U41687 ( .A1(n39192), .A2(n37882), .ZN(n39359) );
  XNOR2_X1 U41688 ( .A(n36992), .B(n36991), .ZN(n37126) );
  XNOR2_X1 U41689 ( .A(n36994), .B(n42769), .ZN(n36995) );
  XNOR2_X1 U41690 ( .A(n36996), .B(n36995), .ZN(n36997) );
  XNOR2_X1 U41691 ( .A(n36998), .B(n36997), .ZN(n37000) );
  XNOR2_X1 U41692 ( .A(n37004), .B(n37003), .ZN(n37007) );
  INV_X1 U41693 ( .A(n37005), .ZN(n37006) );
  XNOR2_X2 U41694 ( .A(n37007), .B(n37006), .ZN(n39377) );
  XNOR2_X1 U41695 ( .A(n37138), .B(n37008), .ZN(n37011) );
  XNOR2_X1 U41696 ( .A(n37009), .B(n4431), .ZN(n37010) );
  XNOR2_X1 U41697 ( .A(n37011), .B(n37010), .ZN(n37012) );
  XNOR2_X1 U41698 ( .A(n37013), .B(n37012), .ZN(n37014) );
  XNOR2_X1 U41699 ( .A(n37015), .B(n37014), .ZN(n37016) );
  XNOR2_X1 U41700 ( .A(n37017), .B(n37016), .ZN(n37018) );
  XNOR2_X1 U41701 ( .A(n37021), .B(n50982), .ZN(n37022) );
  XNOR2_X1 U41702 ( .A(n37024), .B(n37023), .ZN(n37025) );
  NOR2_X1 U41704 ( .A1(n39388), .A2(n51322), .ZN(n37026) );
  NOR2_X1 U41705 ( .A1(n39359), .A2(n37026), .ZN(n37030) );
  NOR2_X1 U41706 ( .A1(n37033), .A2(n51322), .ZN(n39366) );
  OR2_X1 U41708 ( .A1(n51102), .A2(n39195), .ZN(n39360) );
  OAI211_X1 U41709 ( .C1(n39366), .C2(n39361), .A(n38963), .B(n39360), .ZN(
        n37029) );
  INV_X1 U41710 ( .A(n39388), .ZN(n39198) );
  NAND3_X1 U41711 ( .A1(n39198), .A2(n38962), .A3(n39360), .ZN(n37028) );
  NAND3_X1 U41712 ( .A1(n39376), .A2(n39378), .A3(n39194), .ZN(n37027) );
  OAI21_X1 U41713 ( .B1(n39360), .B2(n37033), .A(n38966), .ZN(n37036) );
  NAND2_X1 U41714 ( .A1(n41735), .A2(n41113), .ZN(n41115) );
  NAND2_X1 U41715 ( .A1(n41111), .A2(n41268), .ZN(n40477) );
  INV_X1 U41716 ( .A(n39191), .ZN(n37035) );
  OAI21_X1 U41717 ( .B1(n37036), .B2(n37035), .A(n39369), .ZN(n37038) );
  NAND2_X1 U41718 ( .A1(n37038), .A2(n37037), .ZN(n37169) );
  XNOR2_X1 U41719 ( .A(n37041), .B(n37040), .ZN(n37050) );
  XNOR2_X1 U41720 ( .A(n37043), .B(n37042), .ZN(n37044) );
  XNOR2_X1 U41721 ( .A(n37045), .B(n37044), .ZN(n37046) );
  XNOR2_X1 U41722 ( .A(n37048), .B(n37047), .ZN(n37049) );
  XNOR2_X1 U41723 ( .A(n37050), .B(n37049), .ZN(n37057) );
  XNOR2_X1 U41724 ( .A(n37052), .B(n37051), .ZN(n37055) );
  INV_X1 U41725 ( .A(n37053), .ZN(n37054) );
  XNOR2_X1 U41726 ( .A(n37054), .B(n37055), .ZN(n37056) );
  XNOR2_X1 U41727 ( .A(n37058), .B(n43878), .ZN(n37059) );
  XNOR2_X1 U41728 ( .A(n37060), .B(n37059), .ZN(n37061) );
  XNOR2_X1 U41729 ( .A(n37062), .B(n37061), .ZN(n37064) );
  XNOR2_X1 U41730 ( .A(n37064), .B(n37063), .ZN(n37069) );
  XNOR2_X1 U41731 ( .A(n37066), .B(n37065), .ZN(n37068) );
  XNOR2_X1 U41732 ( .A(n37068), .B(n37067), .ZN(n37235) );
  XNOR2_X1 U41733 ( .A(n37235), .B(n37069), .ZN(n37070) );
  XNOR2_X1 U41734 ( .A(n37071), .B(n37070), .ZN(n37076) );
  XNOR2_X1 U41735 ( .A(n37072), .B(n37243), .ZN(n37073) );
  XNOR2_X1 U41736 ( .A(n37074), .B(n37073), .ZN(n37075) );
  XNOR2_X1 U41737 ( .A(n37079), .B(n37078), .ZN(n37080) );
  XNOR2_X1 U41738 ( .A(n37082), .B(n4295), .ZN(n37083) );
  XNOR2_X1 U41739 ( .A(n37084), .B(n37083), .ZN(n37085) );
  XNOR2_X1 U41740 ( .A(n37086), .B(n37085), .ZN(n37087) );
  XNOR2_X1 U41741 ( .A(n37088), .B(n37087), .ZN(n37090) );
  XNOR2_X1 U41742 ( .A(n37090), .B(n37089), .ZN(n37092) );
  XNOR2_X1 U41743 ( .A(n37091), .B(n37092), .ZN(n37093) );
  NAND2_X1 U41744 ( .A1(n38662), .A2(n39184), .ZN(n39173) );
  XNOR2_X1 U41745 ( .A(n37095), .B(n37094), .ZN(n37099) );
  XNOR2_X1 U41746 ( .A(n37097), .B(n37096), .ZN(n37098) );
  XNOR2_X1 U41747 ( .A(n37098), .B(n37099), .ZN(n37101) );
  XNOR2_X1 U41748 ( .A(n37101), .B(n37100), .ZN(n37118) );
  INV_X1 U41749 ( .A(n37102), .ZN(n37106) );
  XNOR2_X1 U41750 ( .A(n37104), .B(n37103), .ZN(n37105) );
  XNOR2_X1 U41751 ( .A(n37106), .B(n37105), .ZN(n37107) );
  XNOR2_X1 U41752 ( .A(n37108), .B(n37109), .ZN(n37110) );
  XNOR2_X1 U41753 ( .A(n37111), .B(n37110), .ZN(n37116) );
  XNOR2_X1 U41754 ( .A(n37113), .B(n51739), .ZN(n37115) );
  XNOR2_X1 U41755 ( .A(n37114), .B(n37115), .ZN(n37272) );
  XNOR2_X1 U41756 ( .A(n37272), .B(n37116), .ZN(n37117) );
  XNOR2_X2 U41757 ( .A(n37118), .B(n37117), .ZN(n38659) );
  XNOR2_X1 U41758 ( .A(n37120), .B(n37119), .ZN(n37128) );
  INV_X1 U41759 ( .A(n37121), .ZN(n37124) );
  XNOR2_X1 U41760 ( .A(n37122), .B(n274), .ZN(n37123) );
  XNOR2_X1 U41761 ( .A(n37124), .B(n37123), .ZN(n37125) );
  XNOR2_X1 U41762 ( .A(n37126), .B(n37125), .ZN(n37127) );
  XNOR2_X1 U41763 ( .A(n37128), .B(n37127), .ZN(n37132) );
  XNOR2_X1 U41764 ( .A(n37129), .B(n37130), .ZN(n37131) );
  AOI21_X1 U41765 ( .B1(n700), .B2(n37209), .A(n38241), .ZN(n37153) );
  XNOR2_X1 U41766 ( .A(n37133), .B(n37134), .ZN(n37150) );
  XNOR2_X1 U41767 ( .A(n37136), .B(n518), .ZN(n37148) );
  XNOR2_X1 U41768 ( .A(n37138), .B(n43368), .ZN(n37139) );
  XNOR2_X1 U41769 ( .A(n37140), .B(n37139), .ZN(n37143) );
  INV_X1 U41770 ( .A(n37141), .ZN(n37142) );
  XNOR2_X1 U41771 ( .A(n37143), .B(n37142), .ZN(n37144) );
  XNOR2_X1 U41772 ( .A(n33145), .B(n37144), .ZN(n37145) );
  XNOR2_X1 U41773 ( .A(n37146), .B(n37145), .ZN(n37147) );
  XNOR2_X1 U41774 ( .A(n37148), .B(n37147), .ZN(n37149) );
  XNOR2_X1 U41775 ( .A(n37149), .B(n37150), .ZN(n37152) );
  INV_X1 U41776 ( .A(n38241), .ZN(n37928) );
  NAND2_X1 U41777 ( .A1(n38659), .A2(n39184), .ZN(n39167) );
  NAND2_X1 U41778 ( .A1(n38659), .A2(n37209), .ZN(n37155) );
  NAND4_X1 U41779 ( .A1(n39167), .A2(n37927), .A3(n38241), .A4(n37155), .ZN(
        n37156) );
  NAND3_X1 U41780 ( .A1(n37157), .A2(n39182), .A3(n37156), .ZN(n37163) );
  AND2_X1 U41781 ( .A1(n38664), .A2(n38241), .ZN(n39179) );
  NAND3_X1 U41782 ( .A1(n37210), .A2(n39179), .A3(n38667), .ZN(n38248) );
  INV_X1 U41783 ( .A(n39167), .ZN(n38246) );
  NAND2_X1 U41784 ( .A1(n39183), .A2(n38246), .ZN(n37162) );
  AND2_X1 U41785 ( .A1(n37928), .A2(n37158), .ZN(n37925) );
  INV_X1 U41786 ( .A(n37925), .ZN(n37160) );
  NAND2_X1 U41787 ( .A1(n38670), .A2(n37927), .ZN(n37159) );
  NAND4_X1 U41788 ( .A1(n38663), .A2(n39169), .A3(n37160), .A4(n37159), .ZN(
        n37161) );
  NAND4_X2 U41789 ( .A1(n37163), .A2(n38248), .A3(n37162), .A4(n37161), .ZN(
        n41123) );
  NAND2_X1 U41790 ( .A1(n37034), .A2(n41123), .ZN(n37164) );
  OR2_X1 U41791 ( .A1(n37169), .A2(n37164), .ZN(n39594) );
  NOR2_X1 U41792 ( .A1(n39594), .A2(n41735), .ZN(n41729) );
  AND2_X1 U41793 ( .A1(n41268), .A2(n41123), .ZN(n40479) );
  AOI22_X1 U41794 ( .A1(n41729), .A2(n41110), .B1(n40479), .B2(n40486), .ZN(
        n37175) );
  NAND2_X1 U41795 ( .A1(n41263), .A2(n41268), .ZN(n40485) );
  OAI22_X1 U41796 ( .A1(n40485), .A2(n39598), .B1(n40476), .B2(n41256), .ZN(
        n37167) );
  NOR2_X1 U41797 ( .A1(n41735), .A2(n41123), .ZN(n37165) );
  NAND2_X1 U41798 ( .A1(n41110), .A2(n37165), .ZN(n41126) );
  NOR2_X1 U41799 ( .A1(n41257), .A2(n41126), .ZN(n37166) );
  NOR2_X1 U41800 ( .A1(n37167), .A2(n37166), .ZN(n37174) );
  NOR2_X1 U41801 ( .A1(n37169), .A2(n37168), .ZN(n37170) );
  XNOR2_X1 U41802 ( .A(n37170), .B(n41265), .ZN(n37172) );
  AND2_X1 U41803 ( .A1(n41110), .A2(n41735), .ZN(n41727) );
  OAI21_X1 U41804 ( .B1(n37172), .B2(n37171), .A(n41727), .ZN(n37173) );
  NOR2_X1 U41806 ( .A1(n38728), .A2(n39299), .ZN(n37177) );
  OAI21_X1 U41807 ( .B1(n37177), .B2(n38732), .A(n38317), .ZN(n37181) );
  NAND3_X1 U41808 ( .A1(n38720), .A2(n38313), .A3(n39299), .ZN(n37180) );
  NAND3_X1 U41810 ( .A1(n38314), .A2(n38727), .A3(n39300), .ZN(n37178) );
  NAND2_X1 U41812 ( .A1(n38313), .A2(n38727), .ZN(n37183) );
  NAND2_X1 U41813 ( .A1(n39311), .A2(n39293), .ZN(n37184) );
  MUX2_X1 U41814 ( .A(n37184), .B(n39291), .S(n39302), .Z(n37185) );
  OAI21_X1 U41815 ( .B1(n37188), .B2(n3257), .A(n37187), .ZN(n37189) );
  NAND3_X1 U41816 ( .A1(n3257), .A2(n37190), .A3(n6614), .ZN(n37192) );
  NAND3_X1 U41817 ( .A1(n38322), .A2(n38323), .A3(n38334), .ZN(n37193) );
  NOR2_X1 U41818 ( .A1(n38338), .A2(n38330), .ZN(n38347) );
  NOR2_X1 U41819 ( .A1(n6615), .A2(n38337), .ZN(n37194) );
  NOR2_X1 U41820 ( .A1(n38347), .A2(n37194), .ZN(n37196) );
  NAND2_X1 U41821 ( .A1(n40456), .A2(n40453), .ZN(n38368) );
  AND3_X1 U41822 ( .A1(n39264), .A2(n39270), .A3(n39263), .ZN(n37199) );
  AOI22_X1 U41823 ( .A1(n37199), .A2(n37198), .B1(n37941), .B2(n8480), .ZN(
        n37208) );
  NOR2_X1 U41824 ( .A1(n39284), .A2(n39262), .ZN(n37201) );
  INV_X1 U41825 ( .A(n37202), .ZN(n37203) );
  MUX2_X1 U41826 ( .A(n39282), .B(n39012), .S(n39271), .Z(n37205) );
  NAND2_X1 U41827 ( .A1(n38666), .A2(n38670), .ZN(n38679) );
  NAND2_X1 U41828 ( .A1(n700), .A2(n37928), .ZN(n39172) );
  AND2_X1 U41829 ( .A1(n39176), .A2(n39172), .ZN(n37212) );
  OAI21_X1 U41830 ( .B1(n37209), .B2(n38664), .A(n39169), .ZN(n37211) );
  AOI22_X1 U41831 ( .A1(n38679), .A2(n37212), .B1(n37211), .B2(n37210), .ZN(
        n37217) );
  NAND2_X1 U41832 ( .A1(n39179), .A2(n38659), .ZN(n37216) );
  OAI22_X1 U41833 ( .A1(n39182), .A2(n38662), .B1(n38677), .B2(n39176), .ZN(
        n37213) );
  INV_X1 U41835 ( .A(n38237), .ZN(n38672) );
  NAND2_X1 U41836 ( .A1(n37213), .A2(n38672), .ZN(n37215) );
  NOR2_X1 U41837 ( .A1(n39167), .A2(n51496), .ZN(n39171) );
  NAND2_X1 U41838 ( .A1(n39171), .A2(n37927), .ZN(n37214) );
  OAI21_X1 U41839 ( .B1(n38368), .B2(n40447), .A(n39979), .ZN(n37344) );
  INV_X1 U41840 ( .A(n40456), .ZN(n40436) );
  NAND2_X1 U41841 ( .A1(n40447), .A2(n40436), .ZN(n37343) );
  INV_X1 U41842 ( .A(n38632), .ZN(n37686) );
  AOI22_X1 U41843 ( .A1(n38641), .A2(n37688), .B1(n37219), .B2(n197), .ZN(
        n37220) );
  NAND2_X1 U41844 ( .A1(n37686), .A2(n37220), .ZN(n37223) );
  NAND3_X1 U41846 ( .A1(n37688), .A2(n38252), .A3(n37224), .ZN(n37221) );
  AOI21_X1 U41848 ( .B1(n38629), .B2(n37223), .A(n37222), .ZN(n37234) );
  NOR2_X1 U41849 ( .A1(n37688), .A2(n37224), .ZN(n38631) );
  OAI21_X1 U41850 ( .B1(n37677), .B2(n38631), .A(n38255), .ZN(n37233) );
  NOR2_X1 U41851 ( .A1(n38640), .A2(n35310), .ZN(n38265) );
  NOR2_X1 U41852 ( .A1(n37224), .A2(n5989), .ZN(n37227) );
  INV_X1 U41853 ( .A(n38641), .ZN(n37225) );
  OAI22_X1 U41854 ( .A1(n38262), .A2(n38257), .B1(n37225), .B2(n38637), .ZN(
        n37226) );
  AND2_X1 U41855 ( .A1(n68), .A2(n2188), .ZN(n38636) );
  INV_X1 U41856 ( .A(n37688), .ZN(n37229) );
  MUX2_X1 U41857 ( .A(n37229), .B(n37228), .S(n68), .Z(n37230) );
  OAI21_X1 U41858 ( .B1(n37230), .B2(n35310), .A(n37689), .ZN(n37231) );
  NOR2_X1 U41859 ( .A1(n37345), .A2(n40456), .ZN(n38370) );
  XNOR2_X1 U41860 ( .A(n37235), .B(n37236), .ZN(n37238) );
  XNOR2_X1 U41861 ( .A(n37238), .B(n37237), .ZN(n37247) );
  XNOR2_X1 U41862 ( .A(n43592), .B(n37239), .ZN(n37240) );
  XNOR2_X1 U41863 ( .A(n37241), .B(n37240), .ZN(n37242) );
  XNOR2_X1 U41864 ( .A(n37243), .B(n37242), .ZN(n37245) );
  XNOR2_X1 U41865 ( .A(n37245), .B(n37244), .ZN(n37246) );
  XNOR2_X1 U41866 ( .A(n37247), .B(n37246), .ZN(n37248) );
  XNOR2_X1 U41868 ( .A(n37252), .B(n619), .ZN(n37254) );
  XNOR2_X1 U41869 ( .A(n37254), .B(n37253), .ZN(n37255) );
  XNOR2_X1 U41870 ( .A(n37256), .B(n37255), .ZN(n37267) );
  INV_X1 U41871 ( .A(n37257), .ZN(n37259) );
  XNOR2_X1 U41872 ( .A(n37259), .B(n37258), .ZN(n37260) );
  XNOR2_X1 U41873 ( .A(n37261), .B(n37260), .ZN(n37263) );
  XNOR2_X1 U41874 ( .A(n37262), .B(n37263), .ZN(n37265) );
  XNOR2_X1 U41875 ( .A(n37265), .B(n37264), .ZN(n37266) );
  XNOR2_X1 U41876 ( .A(n37267), .B(n37266), .ZN(n37268) );
  XNOR2_X1 U41877 ( .A(n37269), .B(n37270), .ZN(n37271) );
  XNOR2_X1 U41878 ( .A(n37271), .B(n37272), .ZN(n37281) );
  XNOR2_X1 U41879 ( .A(n42918), .B(n37273), .ZN(n37274) );
  XNOR2_X1 U41880 ( .A(n37275), .B(n37274), .ZN(n37276) );
  XOR2_X1 U41882 ( .A(n37280), .B(n37281), .Z(n37282) );
  NAND2_X1 U41883 ( .A1(n38706), .A2(n51507), .ZN(n37912) );
  XNOR2_X1 U41884 ( .A(n37285), .B(n37284), .ZN(n37287) );
  XNOR2_X1 U41885 ( .A(n37289), .B(n37288), .ZN(n37290) );
  XNOR2_X1 U41886 ( .A(n37293), .B(n37292), .ZN(n37295) );
  XNOR2_X1 U41887 ( .A(n37295), .B(n37294), .ZN(n37297) );
  XNOR2_X1 U41888 ( .A(n37297), .B(n37296), .ZN(n37298) );
  XNOR2_X1 U41890 ( .A(n37299), .B(n4885), .ZN(n37300) );
  XNOR2_X1 U41891 ( .A(n37301), .B(n37300), .ZN(n37302) );
  XNOR2_X1 U41892 ( .A(n37303), .B(n37302), .ZN(n37305) );
  XNOR2_X1 U41893 ( .A(n37304), .B(n37305), .ZN(n37306) );
  XNOR2_X1 U41894 ( .A(n37307), .B(n37306), .ZN(n37308) );
  XNOR2_X1 U41895 ( .A(n37314), .B(n49414), .ZN(n37315) );
  XNOR2_X1 U41896 ( .A(n37316), .B(n37315), .ZN(n37317) );
  XNOR2_X1 U41897 ( .A(n37319), .B(n37318), .ZN(n37320) );
  XNOR2_X1 U41900 ( .A(n37325), .B(n37324), .ZN(n37326) );
  XNOR2_X1 U41901 ( .A(n37328), .B(n37327), .ZN(n37330) );
  XNOR2_X1 U41902 ( .A(n37330), .B(n37329), .ZN(n37333) );
  INV_X1 U41903 ( .A(n37331), .ZN(n37332) );
  NAND2_X1 U41905 ( .A1(n39236), .A2(n38704), .ZN(n37334) );
  OAI211_X1 U41906 ( .C1(n37912), .C2(n39236), .A(n37335), .B(n37334), .ZN(
        n37339) );
  INV_X1 U41907 ( .A(n39221), .ZN(n37702) );
  NAND2_X1 U41908 ( .A1(n37911), .A2(n51507), .ZN(n39232) );
  NAND3_X1 U41909 ( .A1(n37702), .A2(n38706), .A3(n39232), .ZN(n37338) );
  NOR2_X1 U41910 ( .A1(n37916), .A2(n51508), .ZN(n39239) );
  INV_X1 U41911 ( .A(n38706), .ZN(n37336) );
  NAND2_X1 U41912 ( .A1(n39239), .A2(n37336), .ZN(n37337) );
  NOR2_X1 U41913 ( .A1(n39233), .A2(n51508), .ZN(n38301) );
  NOR2_X1 U41914 ( .A1(n37911), .A2(n51063), .ZN(n37341) );
  INV_X1 U41915 ( .A(n38303), .ZN(n37701) );
  NAND2_X1 U41916 ( .A1(n38701), .A2(n37283), .ZN(n38298) );
  INV_X1 U41917 ( .A(n38298), .ZN(n37340) );
  NAND3_X1 U41918 ( .A1(n38704), .A2(n6343), .A3(n51736), .ZN(n39242) );
  AOI22_X1 U41919 ( .A1(n37344), .A2(n37343), .B1(n38370), .B2(n39978), .ZN(
        n37351) );
  NAND2_X1 U41921 ( .A1(n37345), .A2(n40456), .ZN(n40402) );
  NOR2_X1 U41922 ( .A1(n6851), .A2(n40403), .ZN(n37346) );
  NOR2_X1 U41923 ( .A1(n40402), .A2(n37346), .ZN(n37347) );
  OAI21_X1 U41924 ( .B1(n39741), .B2(n40446), .A(n37347), .ZN(n37349) );
  NAND3_X1 U41925 ( .A1(n39990), .A2(n40404), .A3(n40456), .ZN(n37348) );
  XNOR2_X1 U41927 ( .A(n37352), .B(n608), .ZN(n43029) );
  XNOR2_X1 U41928 ( .A(n37353), .B(n43029), .ZN(n37354) );
  NAND2_X1 U41929 ( .A1(n38448), .A2(n37356), .ZN(n37355) );
  MUX2_X1 U41930 ( .A(n37355), .B(n39789), .S(n39908), .Z(n37358) );
  NAND2_X1 U41932 ( .A1(n39782), .A2(n51377), .ZN(n38446) );
  INV_X1 U41933 ( .A(n38446), .ZN(n37357) );
  NAND2_X1 U41934 ( .A1(n39562), .A2(n38445), .ZN(n37359) );
  NAND2_X1 U41935 ( .A1(n37363), .A2(n37362), .ZN(n45382) );
  NAND2_X1 U41936 ( .A1(n37364), .A2(n37377), .ZN(n37365) );
  NAND2_X1 U41937 ( .A1(n37368), .A2(n37367), .ZN(n37369) );
  OAI211_X1 U41938 ( .C1(n37373), .C2(n37591), .A(n690), .B(n37585), .ZN(
        n37374) );
  AND2_X1 U41939 ( .A1(n37375), .A2(n37374), .ZN(n40061) );
  INV_X1 U41940 ( .A(n431), .ZN(n40585) );
  AND2_X1 U41941 ( .A1(n37384), .A2(n37516), .ZN(n37388) );
  INV_X1 U41942 ( .A(n37520), .ZN(n37528) );
  NAND2_X1 U41943 ( .A1(n37528), .A2(n38505), .ZN(n37391) );
  INV_X1 U41944 ( .A(n37521), .ZN(n37389) );
  OAI21_X1 U41945 ( .B1(n37389), .B2(n38494), .A(n38505), .ZN(n37390) );
  NAND2_X1 U41946 ( .A1(n38490), .A2(n37394), .ZN(n37395) );
  NAND3_X1 U41947 ( .A1(n37554), .A2(n37410), .A3(n37396), .ZN(n37402) );
  INV_X1 U41948 ( .A(n37397), .ZN(n37398) );
  NAND3_X1 U41949 ( .A1(n37398), .A2(n37410), .A3(n37557), .ZN(n37401) );
  NAND2_X1 U41950 ( .A1(n37535), .A2(n37399), .ZN(n37400) );
  OR2_X1 U41951 ( .A1(n37403), .A2(n37553), .ZN(n37409) );
  INV_X1 U41952 ( .A(n37404), .ZN(n37534) );
  MUX2_X1 U41953 ( .A(n37409), .B(n37534), .S(n37547), .Z(n37413) );
  NAND2_X1 U41954 ( .A1(n37405), .A2(n525), .ZN(n37408) );
  OAI22_X1 U41955 ( .A1(n37553), .A2(n37557), .B1(n37545), .B2(n37406), .ZN(
        n37407) );
  AND2_X1 U41956 ( .A1(n37561), .A2(n37560), .ZN(n37552) );
  AOI22_X1 U41957 ( .A1(n37408), .A2(n37535), .B1(n37407), .B2(n37552), .ZN(
        n37412) );
  INV_X1 U41958 ( .A(n37409), .ZN(n37411) );
  NAND2_X1 U41959 ( .A1(n37411), .A2(n37410), .ZN(n37541) );
  INV_X1 U41960 ( .A(n38110), .ZN(n37419) );
  OAI21_X1 U41961 ( .B1(n38119), .B2(n38485), .A(n37417), .ZN(n37418) );
  NOR2_X1 U41962 ( .A1(n37420), .A2(n38471), .ZN(n37421) );
  INV_X1 U41963 ( .A(n38473), .ZN(n38107) );
  AOI22_X1 U41964 ( .A1(n37415), .A2(n37421), .B1(n38107), .B2(n38484), .ZN(
        n37429) );
  INV_X1 U41965 ( .A(n37422), .ZN(n37424) );
  NOR2_X1 U41966 ( .A1(n38108), .A2(n38471), .ZN(n37423) );
  OAI21_X1 U41967 ( .B1(n37424), .B2(n37423), .A(n38116), .ZN(n37428) );
  NAND2_X1 U41968 ( .A1(n37426), .A2(n37425), .ZN(n37427) );
  NOR2_X1 U41969 ( .A1(n38513), .A2(n37489), .ZN(n38520) );
  OAI211_X1 U41970 ( .C1(n38520), .C2(n37431), .A(n38517), .B(n51411), .ZN(
        n37447) );
  NAND2_X1 U41971 ( .A1(n38521), .A2(n38522), .ZN(n37435) );
  INV_X1 U41972 ( .A(n38517), .ZN(n37485) );
  INV_X1 U41973 ( .A(n37436), .ZN(n37443) );
  NAND3_X1 U41974 ( .A1(n37438), .A2(n51363), .A3(n37437), .ZN(n37441) );
  NAND3_X1 U41975 ( .A1(n38522), .A2(n38514), .A3(n37439), .ZN(n37440) );
  NAND4_X1 U41976 ( .A1(n37443), .A2(n37442), .A3(n37441), .A4(n37440), .ZN(
        n37444) );
  INV_X1 U41977 ( .A(n38596), .ZN(n37449) );
  AOI22_X1 U41978 ( .A1(n37449), .A2(n38165), .B1(n693), .B2(n51429), .ZN(
        n37459) );
  NAND2_X1 U41979 ( .A1(n37568), .A2(n37450), .ZN(n37451) );
  NAND2_X1 U41980 ( .A1(n37451), .A2(n38153), .ZN(n37458) );
  OAI22_X1 U41981 ( .A1(n37453), .A2(n38589), .B1(n37452), .B2(n38584), .ZN(
        n37454) );
  NAND2_X1 U41982 ( .A1(n37454), .A2(n37576), .ZN(n37457) );
  NAND2_X1 U41983 ( .A1(n38592), .A2(n38585), .ZN(n37455) );
  OAI211_X1 U41984 ( .C1(n38153), .C2(n38593), .A(n37455), .B(n38584), .ZN(
        n37456) );
  NOR2_X1 U41985 ( .A1(n40774), .A2(n426), .ZN(n39801) );
  XNOR2_X1 U41986 ( .A(n40776), .B(n426), .ZN(n37460) );
  INV_X1 U41987 ( .A(n40590), .ZN(n37461) );
  NOR2_X1 U41988 ( .A1(n432), .A2(n40768), .ZN(n39802) );
  AOI22_X1 U41989 ( .A1(n37461), .A2(n39802), .B1(n40600), .B2(n40786), .ZN(
        n37463) );
  AND2_X1 U41990 ( .A1(n40768), .A2(n40775), .ZN(n40073) );
  AND2_X1 U41991 ( .A1(n431), .A2(n40777), .ZN(n40787) );
  NOR3_X1 U41992 ( .A1(n40768), .A2(n40775), .A3(n426), .ZN(n37462) );
  XNOR2_X1 U41993 ( .A(n43123), .B(n51371), .ZN(n37479) );
  NOR2_X1 U41994 ( .A1(n37468), .A2(n40556), .ZN(n40552) );
  INV_X1 U41995 ( .A(n40559), .ZN(n37465) );
  AOI22_X1 U41997 ( .A1(n40552), .A2(n40154), .B1(n37466), .B2(n40558), .ZN(
        n37472) );
  NOR2_X1 U41998 ( .A1(n40573), .A2(n40567), .ZN(n37467) );
  NOR2_X1 U41999 ( .A1(n40556), .A2(n40558), .ZN(n40147) );
  AOI22_X1 U42000 ( .A1(n37467), .A2(n40154), .B1(n2597), .B2(n40147), .ZN(
        n37471) );
  INV_X1 U42001 ( .A(n40556), .ZN(n40156) );
  AND2_X1 U42002 ( .A1(n40558), .A2(n40316), .ZN(n40148) );
  NAND3_X1 U42003 ( .A1(n40148), .A2(n40567), .A3(n52159), .ZN(n37470) );
  XNOR2_X1 U42004 ( .A(n37474), .B(n37473), .ZN(n37475) );
  XNOR2_X1 U42005 ( .A(n37476), .B(n37475), .ZN(n37477) );
  XNOR2_X1 U42006 ( .A(n43225), .B(n37477), .ZN(n37478) );
  XNOR2_X1 U42007 ( .A(n37479), .B(n37478), .ZN(n37832) );
  NAND2_X1 U42008 ( .A1(n38532), .A2(n38515), .ZN(n37482) );
  OAI22_X1 U42009 ( .A1(n37491), .A2(n51411), .B1(n51487), .B2(n51363), .ZN(
        n37481) );
  MUX2_X1 U42010 ( .A(n37482), .B(n37481), .S(n37480), .Z(n37495) );
  NAND2_X1 U42011 ( .A1(n37483), .A2(n38535), .ZN(n37487) );
  NAND2_X1 U42012 ( .A1(n37485), .A2(n51411), .ZN(n37486) );
  AOI22_X1 U42014 ( .A1(n51735), .A2(n37489), .B1(n38528), .B2(n51487), .ZN(
        n37493) );
  NAND3_X1 U42015 ( .A1(n37491), .A2(n37490), .A3(n38514), .ZN(n37492) );
  NAND2_X1 U42017 ( .A1(n37497), .A2(n37496), .ZN(n37506) );
  OAI211_X1 U42018 ( .C1(n37500), .C2(n37499), .A(n37498), .B(n37756), .ZN(
        n37505) );
  NAND3_X1 U42019 ( .A1(n37766), .A2(n37510), .A3(n37764), .ZN(n37768) );
  NAND2_X1 U42020 ( .A1(n37749), .A2(n37511), .ZN(n37509) );
  NAND2_X1 U42021 ( .A1(n37507), .A2(n37762), .ZN(n37508) );
  NAND3_X1 U42022 ( .A1(n37511), .A2(n37510), .A3(n37753), .ZN(n37512) );
  NAND4_X1 U42023 ( .A1(n37521), .A2(n37520), .A3(n38494), .A4(n618), .ZN(
        n37522) );
  NAND2_X1 U42024 ( .A1(n37529), .A2(n37528), .ZN(n37530) );
  INV_X1 U42025 ( .A(n37533), .ZN(n37537) );
  NOR2_X1 U42026 ( .A1(n3164), .A2(n37534), .ZN(n37536) );
  OAI21_X1 U42027 ( .B1(n37537), .B2(n37536), .A(n37535), .ZN(n37542) );
  NOR2_X1 U42028 ( .A1(n37544), .A2(n37543), .ZN(n37546) );
  OAI211_X1 U42029 ( .C1(n37547), .C2(n37546), .A(n37545), .B(n37552), .ZN(
        n37549) );
  AND2_X1 U42030 ( .A1(n37549), .A2(n37548), .ZN(n37567) );
  NAND3_X1 U42031 ( .A1(n37554), .A2(n37553), .A3(n37552), .ZN(n37555) );
  AND2_X1 U42032 ( .A1(n37556), .A2(n37555), .ZN(n37566) );
  NAND3_X1 U42033 ( .A1(n37559), .A2(n37558), .A3(n37557), .ZN(n37565) );
  OAI21_X1 U42034 ( .B1(n37396), .B2(n37561), .A(n37560), .ZN(n37563) );
  NAND2_X1 U42035 ( .A1(n37563), .A2(n37562), .ZN(n37564) );
  INV_X1 U42036 ( .A(n37572), .ZN(n37575) );
  INV_X1 U42037 ( .A(n37568), .ZN(n37570) );
  OAI21_X1 U42038 ( .B1(n37570), .B2(n37569), .A(n38596), .ZN(n37574) );
  AOI21_X1 U42039 ( .B1(n37572), .B2(n38585), .A(n37571), .ZN(n37573) );
  OAI21_X1 U42040 ( .B1(n37575), .B2(n37574), .A(n37573), .ZN(n37584) );
  INV_X1 U42041 ( .A(n38582), .ZN(n37578) );
  INV_X1 U42042 ( .A(n38584), .ZN(n38591) );
  OAI21_X1 U42043 ( .B1(n38591), .B2(n37580), .A(n37579), .ZN(n37581) );
  INV_X1 U42044 ( .A(n37581), .ZN(n37583) );
  NAND2_X1 U42045 ( .A1(n37586), .A2(n37585), .ZN(n37589) );
  MUX2_X1 U42046 ( .A(n37589), .B(n37588), .S(n37587), .Z(n37602) );
  AOI22_X1 U42047 ( .A1(n37592), .A2(n37590), .B1(n37591), .B2(n694), .ZN(
        n37601) );
  OAI21_X1 U42048 ( .B1(n37595), .B2(n694), .A(n37594), .ZN(n37600) );
  NAND3_X1 U42049 ( .A1(n37598), .A2(n37597), .A3(n37596), .ZN(n37599) );
  NAND2_X1 U42050 ( .A1(n43325), .A2(n43327), .ZN(n37603) );
  OAI22_X1 U42053 ( .A1(n37609), .A2(n37604), .B1(n37603), .B2(n40800), .ZN(
        n37608) );
  NAND3_X1 U42054 ( .A1(n43325), .A2(n37605), .A3(n40807), .ZN(n37606) );
  NOR2_X1 U42055 ( .A1(n37608), .A2(n37607), .ZN(n37615) );
  INV_X1 U42056 ( .A(n37609), .ZN(n38755) );
  NAND2_X1 U42057 ( .A1(n38764), .A2(n51358), .ZN(n39614) );
  AOI21_X1 U42058 ( .B1(n38755), .B2(n39576), .A(n37610), .ZN(n37614) );
  NAND2_X1 U42059 ( .A1(n43328), .A2(n43327), .ZN(n41020) );
  AND2_X1 U42060 ( .A1(n5911), .A2(n39576), .ZN(n38765) );
  NAND2_X1 U42061 ( .A1(n38765), .A2(n41008), .ZN(n37612) );
  AND2_X1 U42062 ( .A1(n39576), .A2(n43327), .ZN(n40799) );
  INV_X1 U42063 ( .A(n40799), .ZN(n37611) );
  MUX2_X1 U42064 ( .A(n37612), .B(n37611), .S(n7000), .Z(n37613) );
  NAND4_X1 U42065 ( .A1(n37616), .A2(n37624), .A3(n38277), .A4(n613), .ZN(
        n37622) );
  OAI21_X1 U42066 ( .B1(n37617), .B2(n38275), .A(n38279), .ZN(n37621) );
  INV_X1 U42068 ( .A(n37632), .ZN(n37634) );
  NAND2_X1 U42069 ( .A1(n37634), .A2(n5590), .ZN(n37652) );
  OAI21_X1 U42070 ( .B1(n37637), .B2(n37636), .A(n37635), .ZN(n37642) );
  OAI21_X1 U42071 ( .B1(n37640), .B2(n37639), .A(n37638), .ZN(n37641) );
  OAI211_X2 U42072 ( .C1(n37653), .C2(n37652), .A(n37651), .B(n37650), .ZN(
        n40838) );
  AND2_X1 U42073 ( .A1(n40838), .A2(n51990), .ZN(n40143) );
  MUX2_X1 U42075 ( .A(n38314), .B(n39291), .S(n39302), .Z(n37655) );
  AND2_X1 U42076 ( .A1(n38728), .A2(n38313), .ZN(n39308) );
  AOI22_X1 U42077 ( .A1(n38720), .A2(n39291), .B1(n39308), .B2(n39293), .ZN(
        n37662) );
  INV_X1 U42078 ( .A(n38310), .ZN(n37657) );
  NAND2_X1 U42079 ( .A1(n37657), .A2(n39288), .ZN(n37661) );
  INV_X1 U42080 ( .A(n39300), .ZN(n37658) );
  NAND3_X1 U42081 ( .A1(n2436), .A2(n37659), .A3(n37658), .ZN(n37660) );
  INV_X1 U42082 ( .A(n38337), .ZN(n37671) );
  NOR2_X1 U42084 ( .A1(n38338), .A2(n38341), .ZN(n37672) );
  AOI22_X1 U42085 ( .A1(n37672), .A2(n37671), .B1(n37670), .B2(n38341), .ZN(
        n37675) );
  INV_X1 U42086 ( .A(n40820), .ZN(n39697) );
  NAND2_X1 U42087 ( .A1(n37677), .A2(n38629), .ZN(n37694) );
  NAND3_X1 U42088 ( .A1(n38640), .A2(n38629), .A3(n35305), .ZN(n37678) );
  OAI21_X1 U42089 ( .B1(n38633), .B2(n5990), .A(n37678), .ZN(n37679) );
  INV_X1 U42090 ( .A(n37679), .ZN(n37693) );
  INV_X1 U42091 ( .A(n38629), .ZN(n37681) );
  NAND4_X1 U42092 ( .A1(n37683), .A2(n37682), .A3(n38630), .A4(n37681), .ZN(
        n37687) );
  INV_X1 U42093 ( .A(n38262), .ZN(n37684) );
  NAND3_X1 U42094 ( .A1(n37684), .A2(n2188), .A3(n38641), .ZN(n37685) );
  AND3_X1 U42095 ( .A1(n37687), .A2(n37686), .A3(n37685), .ZN(n37692) );
  NOR2_X1 U42096 ( .A1(n37688), .A2(n2188), .ZN(n37690) );
  OAI21_X1 U42097 ( .B1(n38265), .B2(n37690), .A(n37689), .ZN(n37691) );
  NAND4_X2 U42098 ( .A1(n37692), .A2(n37694), .A3(n37693), .A4(n37691), .ZN(
        n40818) );
  INV_X1 U42099 ( .A(n40818), .ZN(n39512) );
  INV_X1 U42101 ( .A(n39233), .ZN(n37910) );
  NAND3_X1 U42103 ( .A1(n38699), .A2(n38700), .A3(n37910), .ZN(n37700) );
  INV_X1 U42104 ( .A(n39242), .ZN(n37698) );
  OAI211_X1 U42105 ( .C1(n39245), .C2(n37698), .A(n37697), .B(n39243), .ZN(
        n37699) );
  AND2_X1 U42106 ( .A1(n51508), .A2(n3874), .ZN(n38299) );
  NAND3_X1 U42107 ( .A1(n38299), .A2(n39245), .A3(n39240), .ZN(n37703) );
  INV_X1 U42108 ( .A(n39695), .ZN(n40828) );
  OAI21_X1 U42109 ( .B1(n40815), .B2(n40817), .A(n40828), .ZN(n37706) );
  NAND3_X1 U42110 ( .A1(n39693), .A2(n39512), .A3(n37706), .ZN(n37707) );
  OR2_X1 U42111 ( .A1(n40838), .A2(n40823), .ZN(n39689) );
  AND2_X1 U42112 ( .A1(n39077), .A2(n40818), .ZN(n40840) );
  INV_X1 U42113 ( .A(n40840), .ZN(n37709) );
  OAI21_X1 U42114 ( .B1(n39689), .B2(n37709), .A(n40822), .ZN(n37710) );
  OR2_X1 U42115 ( .A1(n40838), .A2(n40822), .ZN(n39691) );
  NOR2_X1 U42116 ( .A1(n40815), .A2(n40822), .ZN(n39513) );
  NOR2_X1 U42117 ( .A1(n51455), .A2(n40818), .ZN(n37712) );
  NOR2_X1 U42118 ( .A1(n51455), .A2(n40815), .ZN(n37711) );
  NAND2_X1 U42119 ( .A1(n40822), .A2(n52151), .ZN(n40836) );
  INV_X1 U42120 ( .A(n40836), .ZN(n40133) );
  AOI22_X1 U42121 ( .A1(n39513), .A2(n37712), .B1(n37711), .B2(n40133), .ZN(
        n37714) );
  NAND2_X1 U42123 ( .A1(n39071), .A2(n40831), .ZN(n37713) );
  INV_X1 U42125 ( .A(n37716), .ZN(n37717) );
  NAND3_X1 U42126 ( .A1(n37717), .A2(n51737), .A3(n39030), .ZN(n37725) );
  AOI22_X1 U42127 ( .A1(n39443), .A2(n39448), .B1(n467), .B2(n51389), .ZN(
        n37724) );
  NOR2_X1 U42128 ( .A1(n39445), .A2(n39036), .ZN(n37718) );
  OAI21_X1 U42129 ( .B1(n37719), .B2(n37718), .A(n39438), .ZN(n37723) );
  NAND2_X1 U42130 ( .A1(n467), .A2(n51737), .ZN(n39467) );
  OAI21_X1 U42131 ( .B1(n37894), .B2(n39393), .A(n37726), .ZN(n37727) );
  NAND2_X1 U42132 ( .A1(n37727), .A2(n39003), .ZN(n37729) );
  AOI21_X1 U42133 ( .B1(n37730), .B2(n37892), .A(n39395), .ZN(n37728) );
  NAND2_X1 U42134 ( .A1(n37729), .A2(n37728), .ZN(n37734) );
  NAND2_X1 U42135 ( .A1(n38999), .A2(n3735), .ZN(n37893) );
  NAND2_X1 U42136 ( .A1(n39393), .A2(n37893), .ZN(n37736) );
  AOI21_X1 U42137 ( .B1(n37736), .B2(n37739), .A(n39003), .ZN(n37737) );
  NAND3_X1 U42138 ( .A1(n39005), .A2(n37739), .A3(n39407), .ZN(n37742) );
  NAND2_X1 U42139 ( .A1(n39406), .A2(n39004), .ZN(n37741) );
  OAI22_X1 U42140 ( .A1(n37749), .A2(n37748), .B1(n37747), .B2(n37746), .ZN(
        n37755) );
  AOI21_X1 U42141 ( .B1(n37753), .B2(n37752), .A(n37751), .ZN(n37754) );
  NOR2_X1 U42142 ( .A1(n37755), .A2(n37754), .ZN(n37772) );
  NAND2_X1 U42143 ( .A1(n37765), .A2(n37756), .ZN(n37758) );
  OAI211_X1 U42144 ( .C1(n3650), .C2(n37759), .A(n37758), .B(n37757), .ZN(
        n37761) );
  NAND3_X1 U42145 ( .A1(n37766), .A2(n37765), .A3(n37764), .ZN(n37767) );
  OAI211_X1 U42148 ( .C1(n37780), .C2(n37774), .A(n37773), .B(n39342), .ZN(
        n37777) );
  NAND3_X1 U42149 ( .A1(n37779), .A2(n37782), .A3(n37778), .ZN(n37785) );
  OAI211_X1 U42150 ( .C1(n37783), .C2(n37782), .A(n37781), .B(n37780), .ZN(
        n37784) );
  NOR2_X1 U42151 ( .A1(n39194), .A2(n39388), .ZN(n39358) );
  NAND2_X1 U42152 ( .A1(n39358), .A2(n39361), .ZN(n37797) );
  OAI21_X1 U42153 ( .B1(n37790), .B2(n39195), .A(n37881), .ZN(n37786) );
  NAND2_X1 U42154 ( .A1(n37786), .A2(n51322), .ZN(n37788) );
  AND2_X1 U42155 ( .A1(n39377), .A2(n39195), .ZN(n37878) );
  AND2_X1 U42156 ( .A1(n38962), .A2(n39369), .ZN(n37787) );
  AOI22_X1 U42157 ( .A1(n39381), .A2(n37788), .B1(n37878), .B2(n37787), .ZN(
        n37796) );
  OAI21_X1 U42158 ( .B1(n39379), .B2(n39388), .A(n39189), .ZN(n37789) );
  NAND2_X1 U42159 ( .A1(n37789), .A2(n39380), .ZN(n37795) );
  NAND3_X1 U42160 ( .A1(n39377), .A2(n37790), .A3(n39369), .ZN(n37791) );
  NAND3_X1 U42161 ( .A1(n39367), .A2(n37791), .A3(n39377), .ZN(n37793) );
  NAND2_X1 U42162 ( .A1(n37791), .A2(n37882), .ZN(n37792) );
  NAND3_X1 U42163 ( .A1(n37793), .A2(n39360), .A3(n37792), .ZN(n37794) );
  NAND2_X1 U42164 ( .A1(n42132), .A2(n42154), .ZN(n40257) );
  INV_X1 U42165 ( .A(n37815), .ZN(n42157) );
  OR2_X1 U42167 ( .A1(n39475), .A2(n1075), .ZN(n38977) );
  NAND3_X1 U42168 ( .A1(n37803), .A2(n39479), .A3(n37802), .ZN(n37814) );
  OAI21_X1 U42169 ( .B1(n37810), .B2(n37805), .A(n37804), .ZN(n37808) );
  OAI211_X1 U42170 ( .C1(n2177), .C2(n7159), .A(n473), .B(n37806), .ZN(n37807)
         );
  NAND2_X1 U42171 ( .A1(n37808), .A2(n37807), .ZN(n37812) );
  NAND3_X1 U42172 ( .A1(n37812), .A2(n39472), .A3(n37811), .ZN(n37813) );
  AND2_X1 U42174 ( .A1(n42154), .A2(n51375), .ZN(n40262) );
  NAND2_X1 U42175 ( .A1(n40262), .A2(n52092), .ZN(n42141) );
  OAI211_X1 U42176 ( .C1(n40257), .C2(n52092), .A(n37816), .B(n42141), .ZN(
        n37817) );
  INV_X1 U42177 ( .A(n37817), .ZN(n37821) );
  NOR2_X1 U42178 ( .A1(n42148), .A2(n42145), .ZN(n37819) );
  NOR2_X1 U42179 ( .A1(n42136), .A2(n51375), .ZN(n37818) );
  AND2_X1 U42180 ( .A1(n42136), .A2(n42131), .ZN(n42158) );
  OAI21_X1 U42181 ( .B1(n42132), .B2(n42154), .A(n42144), .ZN(n37820) );
  INV_X1 U42182 ( .A(n41925), .ZN(n39541) );
  INV_X1 U42183 ( .A(n38928), .ZN(n37823) );
  AND2_X1 U42184 ( .A1(n42209), .A2(n40249), .ZN(n41928) );
  OAI21_X1 U42185 ( .B1(n39541), .B2(n6578), .A(n41928), .ZN(n37822) );
  OAI21_X1 U42186 ( .B1(n39541), .B2(n37823), .A(n37822), .ZN(n37826) );
  INV_X1 U42187 ( .A(n42206), .ZN(n37825) );
  OR2_X1 U42188 ( .A1(n38921), .A2(n41938), .ZN(n42208) );
  OAI21_X1 U42189 ( .B1(n42205), .B2(n40249), .A(n6617), .ZN(n42207) );
  NAND3_X1 U42190 ( .A1(n42208), .A2(n42209), .A3(n42207), .ZN(n37830) );
  NAND2_X1 U42191 ( .A1(n41939), .A2(n42205), .ZN(n39542) );
  INV_X1 U42192 ( .A(n39542), .ZN(n37827) );
  INV_X1 U42193 ( .A(n42202), .ZN(n37828) );
  INV_X1 U42194 ( .A(n41942), .ZN(n42203) );
  NAND4_X1 U42195 ( .A1(n37828), .A2(n42203), .A3(n41939), .A4(n39543), .ZN(
        n37829) );
  XNOR2_X1 U42196 ( .A(n44207), .B(n43698), .ZN(n37831) );
  NAND2_X1 U42197 ( .A1(n677), .A2(n52083), .ZN(n37834) );
  MUX2_X1 U42198 ( .A(n7977), .B(n37834), .S(n51012), .Z(n37836) );
  NOR2_X1 U42199 ( .A1(n37836), .A2(n218), .ZN(n37837) );
  NAND2_X1 U42200 ( .A1(n40380), .A2(n41146), .ZN(n37841) );
  NAND3_X1 U42201 ( .A1(n39842), .A2(n38612), .A3(n41150), .ZN(n37840) );
  NAND3_X1 U42202 ( .A1(n38612), .A2(n51012), .A3(n40388), .ZN(n37839) );
  NAND2_X1 U42203 ( .A1(n37838), .A2(n40388), .ZN(n38616) );
  NAND4_X1 U42204 ( .A1(n37841), .A2(n37840), .A3(n37839), .A4(n38616), .ZN(
        n37842) );
  NAND2_X1 U42205 ( .A1(n39103), .A2(n39097), .ZN(n37846) );
  AOI21_X1 U42206 ( .B1(n37843), .B2(n37846), .A(n39995), .ZN(n37845) );
  NAND2_X1 U42207 ( .A1(n40003), .A2(n39097), .ZN(n39104) );
  AOI21_X1 U42208 ( .B1(n37848), .B2(n6740), .A(n39104), .ZN(n37844) );
  NAND2_X1 U42209 ( .A1(n39663), .A2(n51297), .ZN(n37855) );
  OAI21_X1 U42210 ( .B1(n39099), .B2(n39668), .A(n38429), .ZN(n37854) );
  NAND2_X1 U42211 ( .A1(n39097), .A2(n51297), .ZN(n37850) );
  INV_X1 U42212 ( .A(n37846), .ZN(n37847) );
  NAND2_X1 U42213 ( .A1(n37847), .A2(n39101), .ZN(n38418) );
  AND2_X1 U42214 ( .A1(n39103), .A2(n38428), .ZN(n40005) );
  INV_X1 U42215 ( .A(n37848), .ZN(n39662) );
  NAND2_X1 U42216 ( .A1(n40005), .A2(n39662), .ZN(n37849) );
  OAI211_X1 U42217 ( .C1(n40000), .C2(n37850), .A(n38418), .B(n37849), .ZN(
        n37851) );
  INV_X1 U42218 ( .A(n37851), .ZN(n37853) );
  INV_X1 U42219 ( .A(n40014), .ZN(n38424) );
  NAND3_X1 U42220 ( .A1(n6884), .A2(n38424), .A3(n40003), .ZN(n37852) );
  NAND4_X1 U42221 ( .A1(n37855), .A2(n37854), .A3(n37853), .A4(n37852), .ZN(
        n40757) );
  NOR2_X1 U42222 ( .A1(n39943), .A2(n39754), .ZN(n38832) );
  NOR2_X1 U42223 ( .A1(n575), .A2(n39938), .ZN(n37856) );
  NAND3_X1 U42224 ( .A1(n39751), .A2(n39943), .A3(n39754), .ZN(n37857) );
  AND2_X1 U42225 ( .A1(n39112), .A2(n37857), .ZN(n41603) );
  NAND2_X1 U42226 ( .A1(n41607), .A2(n41603), .ZN(n37861) );
  XNOR2_X1 U42227 ( .A(n39938), .B(n52095), .ZN(n37858) );
  OAI21_X1 U42229 ( .B1(n39943), .B2(n37858), .A(n38837), .ZN(n41606) );
  MUX2_X1 U42230 ( .A(n684), .B(n575), .S(n39754), .Z(n37860) );
  NAND4_X1 U42231 ( .A1(n39943), .A2(n39751), .A3(n575), .A4(n39942), .ZN(
        n37859) );
  OAI211_X1 U42232 ( .C1(n37860), .C2(n39943), .A(n39955), .B(n37859), .ZN(
        n41604) );
  NOR2_X1 U42234 ( .A1(n40327), .A2(n40340), .ZN(n38843) );
  NOR2_X1 U42235 ( .A1(n37862), .A2(n40338), .ZN(n37863) );
  NOR2_X1 U42236 ( .A1(n40341), .A2(n52101), .ZN(n39862) );
  AOI22_X1 U42237 ( .A1(n37864), .A2(n38843), .B1(n37863), .B2(n39862), .ZN(
        n37875) );
  NAND2_X1 U42238 ( .A1(n40328), .A2(n40327), .ZN(n39856) );
  NOR2_X1 U42239 ( .A1(n39856), .A2(n37865), .ZN(n37866) );
  OAI21_X1 U42240 ( .B1(n37868), .B2(n40330), .A(n37867), .ZN(n37873) );
  NAND2_X1 U42241 ( .A1(n37869), .A2(n40327), .ZN(n37871) );
  NAND2_X1 U42242 ( .A1(n7117), .A2(n40328), .ZN(n37870) );
  XNOR2_X1 U42244 ( .A(n37876), .B(n45252), .ZN(n45376) );
  OAI21_X1 U42246 ( .B1(n39376), .B2(n37878), .A(n38962), .ZN(n37879) );
  OAI211_X1 U42247 ( .C1(n39361), .C2(n38963), .A(n37879), .B(n39189), .ZN(
        n37880) );
  INV_X1 U42248 ( .A(n39381), .ZN(n39193) );
  AOI22_X1 U42249 ( .A1(n51872), .A2(n39198), .B1(n39379), .B2(n39361), .ZN(
        n37883) );
  NAND2_X1 U42251 ( .A1(n39390), .A2(n51322), .ZN(n38960) );
  OAI211_X1 U42252 ( .C1(n38966), .C2(n39193), .A(n37883), .B(n38960), .ZN(
        n40939) );
  INV_X1 U42253 ( .A(n38997), .ZN(n37887) );
  OAI21_X1 U42254 ( .B1(n37894), .B2(n37885), .A(n39401), .ZN(n37886) );
  OAI211_X1 U42255 ( .C1(n37887), .C2(n39005), .A(n39003), .B(n37886), .ZN(
        n37899) );
  NAND2_X1 U42256 ( .A1(n37891), .A2(n37890), .ZN(n37898) );
  NOR2_X1 U42257 ( .A1(n38991), .A2(n37895), .ZN(n37896) );
  NOR2_X1 U42258 ( .A1(n41544), .A2(n41535), .ZN(n40228) );
  INV_X1 U42259 ( .A(n39426), .ZN(n39411) );
  NAND2_X1 U42260 ( .A1(n37900), .A2(n39410), .ZN(n39206) );
  NAND2_X1 U42261 ( .A1(n38953), .A2(n38940), .ZN(n39210) );
  INV_X1 U42262 ( .A(n39206), .ZN(n38952) );
  NAND2_X1 U42263 ( .A1(n38943), .A2(n38952), .ZN(n37904) );
  OAI22_X1 U42264 ( .A1(n39417), .A2(n37901), .B1(n37907), .B2(n38941), .ZN(
        n37902) );
  NAND2_X1 U42265 ( .A1(n37902), .A2(n39207), .ZN(n37903) );
  NAND4_X1 U42266 ( .A1(n37905), .A2(n37904), .A3(n39421), .A4(n37903), .ZN(
        n37909) );
  NAND2_X1 U42267 ( .A1(n39422), .A2(n39430), .ZN(n37906) );
  NAND2_X1 U42268 ( .A1(n37907), .A2(n38941), .ZN(n39213) );
  OAI21_X1 U42269 ( .B1(n39234), .B2(n39221), .A(n51508), .ZN(n37914) );
  AND2_X1 U42270 ( .A1(n37911), .A2(n51063), .ZN(n38696) );
  NAND3_X1 U42271 ( .A1(n37912), .A2(n38696), .A3(n39246), .ZN(n37913) );
  NOR2_X1 U42272 ( .A1(n37916), .A2(n39243), .ZN(n37918) );
  AOI22_X1 U42273 ( .A1(n38696), .A2(n37918), .B1(n39236), .B2(n37917), .ZN(
        n37920) );
  INV_X1 U42274 ( .A(n39236), .ZN(n38697) );
  NAND3_X1 U42275 ( .A1(n38697), .A2(n38706), .A3(n39245), .ZN(n37919) );
  XNOR2_X1 U42276 ( .A(n41554), .B(n52120), .ZN(n37949) );
  NAND3_X1 U42277 ( .A1(n38659), .A2(n420), .A3(n37924), .ZN(n37921) );
  MUX2_X1 U42278 ( .A(n38662), .B(n38667), .S(n39167), .Z(n37922) );
  NAND2_X1 U42279 ( .A1(n37922), .A2(n39179), .ZN(n37936) );
  OAI21_X1 U42280 ( .B1(n38667), .B2(n37928), .A(n38670), .ZN(n37923) );
  NAND2_X1 U42281 ( .A1(n37923), .A2(n38672), .ZN(n37935) );
  NAND3_X1 U42282 ( .A1(n38672), .A2(n37928), .A3(n38245), .ZN(n37933) );
  AND2_X1 U42283 ( .A1(n37924), .A2(n39184), .ZN(n37926) );
  NAND4_X1 U42284 ( .A1(n37926), .A2(n37925), .A3(n38670), .A4(n700), .ZN(
        n37932) );
  INV_X1 U42285 ( .A(n37926), .ZN(n37930) );
  NOR2_X1 U42286 ( .A1(n51496), .A2(n37927), .ZN(n37929) );
  AND3_X1 U42287 ( .A1(n37933), .A2(n37932), .A3(n37931), .ZN(n37934) );
  INV_X1 U42288 ( .A(n38667), .ZN(n38239) );
  NAND2_X1 U42289 ( .A1(n38246), .A2(n38239), .ZN(n37937) );
  AOI21_X1 U42290 ( .B1(n38658), .B2(n37937), .A(n39182), .ZN(n37938) );
  NAND2_X1 U42291 ( .A1(n41540), .A2(n40989), .ZN(n37948) );
  OAI22_X1 U42292 ( .A1(n36779), .A2(n39284), .B1(n8480), .B2(n39263), .ZN(
        n37939) );
  NAND3_X1 U42293 ( .A1(n37939), .A2(n39007), .A3(n39269), .ZN(n37946) );
  NOR2_X1 U42294 ( .A1(n39258), .A2(n39262), .ZN(n37940) );
  AOI21_X1 U42295 ( .B1(n37941), .B2(n39266), .A(n37940), .ZN(n37945) );
  NOR2_X1 U42296 ( .A1(n37942), .A2(n551), .ZN(n38684) );
  OAI21_X1 U42297 ( .B1(n39258), .B2(n39007), .A(n39262), .ZN(n37944) );
  AND2_X1 U42298 ( .A1(n41524), .A2(n41539), .ZN(n41551) );
  NAND2_X1 U42299 ( .A1(n41551), .A2(n52120), .ZN(n37947) );
  NAND4_X1 U42300 ( .A1(n40228), .A2(n37949), .A3(n37948), .A4(n37947), .ZN(
        n37955) );
  NAND3_X1 U42301 ( .A1(n41544), .A2(n41554), .A3(n41394), .ZN(n37950) );
  OAI211_X1 U42302 ( .C1(n37951), .C2(n41544), .A(n52120), .B(n37950), .ZN(
        n37954) );
  NAND2_X1 U42303 ( .A1(n41395), .A2(n40986), .ZN(n40941) );
  NOR2_X1 U42304 ( .A1(n40941), .A2(n40943), .ZN(n41537) );
  NOR2_X1 U42305 ( .A1(n41556), .A2(n41537), .ZN(n37953) );
  NAND3_X1 U42307 ( .A1(n41554), .A2(n41526), .A3(n40989), .ZN(n37952) );
  NOR2_X1 U42308 ( .A1(n37957), .A2(n37956), .ZN(n37958) );
  OAI21_X1 U42309 ( .B1(n37959), .B2(n37958), .A(n8016), .ZN(n37973) );
  AND2_X1 U42310 ( .A1(n37966), .A2(n37967), .ZN(n37971) );
  NOR2_X1 U42311 ( .A1(n37975), .A2(n37974), .ZN(n37978) );
  AOI22_X1 U42312 ( .A1(n37979), .A2(n37978), .B1(n37977), .B2(n37976), .ZN(
        n37995) );
  OAI21_X1 U42313 ( .B1(n37981), .B2(n37990), .A(n37980), .ZN(n37984) );
  NAND3_X1 U42314 ( .A1(n37984), .A2(n37983), .A3(n37982), .ZN(n37994) );
  NAND3_X1 U42315 ( .A1(n37986), .A2(n37991), .A3(n37985), .ZN(n37993) );
  NAND2_X1 U42316 ( .A1(n37988), .A2(n37987), .ZN(n37989) );
  OAI211_X1 U42317 ( .C1(n37991), .C2(n594), .A(n37990), .B(n37989), .ZN(
        n37992) );
  OAI21_X1 U42318 ( .B1(n37997), .B2(n37996), .A(n38189), .ZN(n37999) );
  INV_X1 U42319 ( .A(n38188), .ZN(n38174) );
  OAI21_X1 U42320 ( .B1(n37997), .B2(n38174), .A(n38014), .ZN(n37998) );
  OAI21_X1 U42321 ( .B1(n38000), .B2(n37999), .A(n37998), .ZN(n38011) );
  NAND3_X1 U42322 ( .A1(n38173), .A2(n38002), .A3(n38001), .ZN(n38176) );
  INV_X1 U42323 ( .A(n38178), .ZN(n38003) );
  OAI21_X1 U42324 ( .B1(n38004), .B2(n38003), .A(n38173), .ZN(n38010) );
  OAI21_X1 U42325 ( .B1(n38007), .B2(n38006), .A(n38005), .ZN(n38008) );
  NAND2_X1 U42326 ( .A1(n38008), .A2(n38192), .ZN(n38009) );
  INV_X1 U42328 ( .A(n38192), .ZN(n38013) );
  INV_X1 U42329 ( .A(n38177), .ZN(n38017) );
  OAI22_X1 U42330 ( .A1(n5872), .A2(n38017), .B1(n38016), .B2(n38015), .ZN(
        n38021) );
  NOR2_X1 U42331 ( .A1(n38019), .A2(n38018), .ZN(n38020) );
  OAI21_X1 U42332 ( .B1(n38022), .B2(n38021), .A(n38020), .ZN(n38023) );
  OAI21_X1 U42333 ( .B1(n38024), .B2(n38190), .A(n38023), .ZN(n38025) );
  NAND2_X1 U42334 ( .A1(n38030), .A2(n38029), .ZN(n38032) );
  MUX2_X1 U42335 ( .A(n38033), .B(n38032), .S(n38031), .Z(n38048) );
  NOR2_X1 U42336 ( .A1(n38038), .A2(n38037), .ZN(n38041) );
  OAI211_X1 U42337 ( .C1(n38042), .C2(n38041), .A(n38040), .B(n38039), .ZN(
        n38046) );
  NAND2_X1 U42338 ( .A1(n38044), .A2(n38043), .ZN(n38045) );
  NOR2_X1 U42339 ( .A1(n40269), .A2(n40909), .ZN(n40094) );
  NAND2_X1 U42340 ( .A1(n5072), .A2(n40094), .ZN(n38049) );
  NAND2_X1 U42341 ( .A1(n40269), .A2(n40909), .ZN(n40892) );
  OAI211_X1 U42342 ( .C1(n40893), .C2(n40274), .A(n38049), .B(n40892), .ZN(
        n38101) );
  OAI211_X1 U42343 ( .C1(n38057), .C2(n38146), .A(n38056), .B(n38055), .ZN(
        n38059) );
  NAND2_X1 U42344 ( .A1(n38059), .A2(n38058), .ZN(n38060) );
  AND2_X1 U42345 ( .A1(n38061), .A2(n38060), .ZN(n38070) );
  NAND2_X1 U42346 ( .A1(n31621), .A2(n38142), .ZN(n38062) );
  OAI22_X1 U42347 ( .A1(n38065), .A2(n38064), .B1(n38063), .B2(n38062), .ZN(
        n38066) );
  NAND2_X1 U42348 ( .A1(n38066), .A2(n38145), .ZN(n38069) );
  OR2_X1 U42349 ( .A1(n38067), .A2(n38146), .ZN(n38134) );
  INV_X1 U42350 ( .A(n38134), .ZN(n38068) );
  NAND2_X1 U42351 ( .A1(n38072), .A2(n38071), .ZN(n38074) );
  NAND2_X1 U42352 ( .A1(n38074), .A2(n38073), .ZN(n38100) );
  INV_X1 U42353 ( .A(n38075), .ZN(n38088) );
  NAND2_X1 U42354 ( .A1(n1360), .A2(n38088), .ZN(n38080) );
  NAND3_X1 U42355 ( .A1(n38086), .A2(n38092), .A3(n50984), .ZN(n38079) );
  INV_X1 U42356 ( .A(n38076), .ZN(n38077) );
  OAI211_X1 U42357 ( .C1(n38080), .C2(n38079), .A(n38078), .B(n38077), .ZN(
        n38081) );
  INV_X1 U42358 ( .A(n38081), .ZN(n38099) );
  NAND2_X1 U42359 ( .A1(n38083), .A2(n38082), .ZN(n38091) );
  NAND2_X1 U42360 ( .A1(n695), .A2(n50984), .ZN(n38085) );
  NOR2_X1 U42361 ( .A1(n38086), .A2(n38085), .ZN(n38090) );
  AOI22_X1 U42363 ( .A1(n38091), .A2(n38090), .B1(n38089), .B2(n38092), .ZN(
        n38098) );
  INV_X1 U42364 ( .A(n38091), .ZN(n38096) );
  NOR2_X1 U42365 ( .A1(n38093), .A2(n38092), .ZN(n38095) );
  OAI21_X1 U42366 ( .B1(n38096), .B2(n38095), .A(n38094), .ZN(n38097) );
  NAND2_X1 U42367 ( .A1(n5072), .A2(n2223), .ZN(n40098) );
  NAND3_X1 U42369 ( .A1(n40098), .A2(n40906), .A3(n40901), .ZN(n38102) );
  AND2_X1 U42370 ( .A1(n40910), .A2(n40269), .ZN(n40897) );
  NAND2_X1 U42371 ( .A1(n40897), .A2(n2224), .ZN(n40083) );
  NOR2_X1 U42372 ( .A1(n40903), .A2(n2224), .ZN(n38794) );
  NOR2_X1 U42373 ( .A1(n40271), .A2(n40909), .ZN(n40268) );
  OAI21_X1 U42374 ( .B1(n38794), .B2(n40269), .A(n40268), .ZN(n38105) );
  NOR2_X1 U42375 ( .A1(n40087), .A2(n40903), .ZN(n40267) );
  NAND2_X1 U42376 ( .A1(n40267), .A2(n40901), .ZN(n38104) );
  AOI22_X1 U42377 ( .A1(n38107), .A2(n38485), .B1(n38468), .B2(n38116), .ZN(
        n38114) );
  NOR2_X1 U42378 ( .A1(n38108), .A2(n6637), .ZN(n38109) );
  INV_X1 U42379 ( .A(n38111), .ZN(n38112) );
  MUX2_X1 U42380 ( .A(n38114), .B(n38113), .S(n38112), .Z(n38130) );
  NAND2_X1 U42381 ( .A1(n38115), .A2(n38119), .ZN(n38121) );
  INV_X1 U42382 ( .A(n38116), .ZN(n38117) );
  OAI22_X1 U42383 ( .A1(n38471), .A2(n38473), .B1(n36115), .B2(n38478), .ZN(
        n38124) );
  NOR2_X1 U42384 ( .A1(n38484), .A2(n38477), .ZN(n38123) );
  OAI21_X1 U42385 ( .B1(n38124), .B2(n38123), .A(n38122), .ZN(n38128) );
  OAI21_X1 U42386 ( .B1(n38126), .B2(n38125), .A(n38480), .ZN(n38127) );
  NAND3_X1 U42387 ( .A1(n38137), .A2(n38132), .A3(n38145), .ZN(n38133) );
  INV_X1 U42388 ( .A(n38136), .ZN(n38139) );
  AND3_X1 U42389 ( .A1(n38139), .A2(n38138), .A3(n38137), .ZN(n38140) );
  NOR2_X1 U42390 ( .A1(n38141), .A2(n38140), .ZN(n38151) );
  NAND2_X1 U42391 ( .A1(n38146), .A2(n38142), .ZN(n38143) );
  NAND3_X1 U42392 ( .A1(n38147), .A2(n38146), .A3(n38145), .ZN(n38149) );
  NAND3_X1 U42393 ( .A1(n693), .A2(n38153), .A3(n38152), .ZN(n38154) );
  AND2_X1 U42394 ( .A1(n38155), .A2(n38154), .ZN(n38171) );
  NAND2_X1 U42395 ( .A1(n38157), .A2(n38156), .ZN(n38163) );
  NAND2_X1 U42396 ( .A1(n38158), .A2(n38164), .ZN(n38162) );
  NAND4_X1 U42397 ( .A1(n38163), .A2(n38166), .A3(n38162), .A4(n38161), .ZN(
        n38170) );
  NAND2_X1 U42398 ( .A1(n38165), .A2(n38164), .ZN(n38583) );
  OR2_X1 U42399 ( .A1(n38583), .A2(n38166), .ZN(n38581) );
  INV_X1 U42400 ( .A(n38581), .ZN(n38168) );
  OAI21_X1 U42401 ( .B1(n38168), .B2(n38591), .A(n38167), .ZN(n38169) );
  AOI21_X1 U42403 ( .B1(n38176), .B2(n38175), .A(n38174), .ZN(n38183) );
  NAND4_X1 U42404 ( .A1(n38181), .A2(n38180), .A3(n38179), .A4(n38178), .ZN(
        n38182) );
  INV_X1 U42405 ( .A(n38184), .ZN(n38187) );
  INV_X1 U42406 ( .A(n38185), .ZN(n38186) );
  OAI21_X1 U42407 ( .B1(n38187), .B2(n38190), .A(n38186), .ZN(n38193) );
  AOI21_X1 U42408 ( .B1(n38193), .B2(n38192), .A(n38191), .ZN(n38194) );
  NAND2_X1 U42410 ( .A1(n38195), .A2(n7759), .ZN(n38209) );
  NOR2_X1 U42411 ( .A1(n38196), .A2(n38200), .ZN(n38197) );
  AOI22_X1 U42412 ( .A1(n38199), .A2(n38566), .B1(n38198), .B2(n38197), .ZN(
        n38208) );
  OAI211_X1 U42413 ( .C1(n6869), .C2(n38201), .A(n33062), .B(n38200), .ZN(
        n38202) );
  INV_X1 U42414 ( .A(n38202), .ZN(n38203) );
  OAI211_X1 U42415 ( .C1(n38204), .C2(n1764), .A(n38203), .B(n38572), .ZN(
        n38207) );
  NAND2_X1 U42416 ( .A1(n51394), .A2(n40972), .ZN(n38232) );
  NAND2_X1 U42417 ( .A1(n38552), .A2(n35175), .ZN(n38211) );
  NAND4_X1 U42418 ( .A1(n38211), .A2(n38210), .A3(n31355), .A4(n38221), .ZN(
        n38225) );
  NAND3_X1 U42419 ( .A1(n6734), .A2(n38212), .A3(n38213), .ZN(n38216) );
  NAND3_X1 U42420 ( .A1(n38214), .A2(n38213), .A3(n35175), .ZN(n38215) );
  NAND2_X1 U42421 ( .A1(n38557), .A2(n38550), .ZN(n38219) );
  NOR2_X1 U42422 ( .A1(n38221), .A2(n38226), .ZN(n38222) );
  NAND2_X1 U42423 ( .A1(n38222), .A2(n38553), .ZN(n38223) );
  NAND4_X1 U42425 ( .A1(n41375), .A2(n38885), .A3(n41380), .A4(n40967), .ZN(
        n38231) );
  AND2_X1 U42426 ( .A1(n40960), .A2(n40972), .ZN(n40953) );
  NAND2_X1 U42427 ( .A1(n40967), .A2(n40953), .ZN(n38896) );
  INV_X1 U42428 ( .A(n41374), .ZN(n38893) );
  NAND2_X1 U42429 ( .A1(n38893), .A2(n40960), .ZN(n40241) );
  INV_X1 U42430 ( .A(n40241), .ZN(n38887) );
  INV_X1 U42432 ( .A(n41380), .ZN(n40959) );
  NOR2_X1 U42433 ( .A1(n40967), .A2(n40972), .ZN(n38235) );
  NAND2_X1 U42434 ( .A1(n41380), .A2(n40972), .ZN(n38233) );
  OAI22_X1 U42435 ( .A1(n38233), .A2(n40241), .B1(n41378), .B2(n41380), .ZN(
        n38234) );
  AOI21_X1 U42436 ( .B1(n41373), .B2(n38235), .A(n38234), .ZN(n38236) );
  NAND2_X1 U42437 ( .A1(n39171), .A2(n38241), .ZN(n39168) );
  AOI21_X1 U42438 ( .B1(n39168), .B2(n38240), .A(n38239), .ZN(n38251) );
  AOI21_X1 U42439 ( .B1(n39176), .B2(n38241), .A(n7729), .ZN(n38244) );
  OAI211_X1 U42440 ( .C1(n39184), .C2(n38241), .A(n420), .B(n700), .ZN(n38242)
         );
  INV_X1 U42441 ( .A(n38242), .ZN(n38243) );
  OAI21_X1 U42442 ( .B1(n38244), .B2(n51496), .A(n38243), .ZN(n38249) );
  NAND2_X1 U42443 ( .A1(n38246), .A2(n38245), .ZN(n38674) );
  NAND2_X1 U42444 ( .A1(n38663), .A2(n39176), .ZN(n38247) );
  NAND4_X1 U42445 ( .A1(n38249), .A2(n38248), .A3(n38674), .A4(n38247), .ZN(
        n38250) );
  NAND3_X1 U42446 ( .A1(n38252), .A2(n38637), .A3(n38259), .ZN(n38253) );
  NAND3_X1 U42447 ( .A1(n38256), .A2(n38255), .A3(n38259), .ZN(n38268) );
  OAI21_X1 U42448 ( .B1(n38259), .B2(n2188), .A(n51360), .ZN(n38260) );
  NAND2_X1 U42449 ( .A1(n38265), .A2(n38264), .ZN(n38266) );
  NOR2_X1 U42451 ( .A1(n40874), .A2(n40868), .ZN(n40531) );
  MUX2_X1 U42452 ( .A(n38270), .B(n34529), .S(n38272), .Z(n38281) );
  OAI21_X1 U42453 ( .B1(n37629), .B2(n38272), .A(n38271), .ZN(n38274) );
  OAI21_X1 U42454 ( .B1(n38276), .B2(n38275), .A(n38274), .ZN(n38278) );
  NAND2_X1 U42455 ( .A1(n38278), .A2(n38277), .ZN(n38280) );
  OAI211_X1 U42456 ( .C1(n38282), .C2(n38281), .A(n38280), .B(n38279), .ZN(
        n38296) );
  AND2_X1 U42457 ( .A1(n38283), .A2(n2120), .ZN(n38287) );
  INV_X1 U42458 ( .A(n38288), .ZN(n38285) );
  AOI22_X1 U42459 ( .A1(n38287), .A2(n38286), .B1(n38285), .B2(n38284), .ZN(
        n38295) );
  OAI22_X1 U42460 ( .A1(n38291), .A2(n38290), .B1(n38289), .B2(n38288), .ZN(
        n38293) );
  NAND2_X1 U42461 ( .A1(n38293), .A2(n38292), .ZN(n38294) );
  NOR2_X1 U42462 ( .A1(n39221), .A2(n51736), .ZN(n39230) );
  NOR2_X1 U42463 ( .A1(n39246), .A2(n38701), .ZN(n38297) );
  NOR2_X1 U42464 ( .A1(n39230), .A2(n38297), .ZN(n38309) );
  OAI22_X1 U42465 ( .A1(n39233), .A2(n38706), .B1(n38298), .B2(n38303), .ZN(
        n38300) );
  NAND2_X1 U42466 ( .A1(n38300), .A2(n38299), .ZN(n38308) );
  NOR2_X1 U42467 ( .A1(n51063), .A2(n51507), .ZN(n38302) );
  NAND2_X1 U42468 ( .A1(n38303), .A2(n39243), .ZN(n38304) );
  NAND2_X1 U42469 ( .A1(n38305), .A2(n38304), .ZN(n38306) );
  NOR2_X1 U42470 ( .A1(n40531), .A2(n40876), .ZN(n38354) );
  OAI211_X1 U42472 ( .C1(n38730), .C2(n38314), .A(n39302), .B(n39300), .ZN(
        n38316) );
  NAND3_X1 U42473 ( .A1(n38720), .A2(n38732), .A3(n39300), .ZN(n38315) );
  MUX2_X1 U42474 ( .A(n7772), .B(n5593), .S(n38317), .Z(n38318) );
  NAND2_X1 U42475 ( .A1(n38318), .A2(n39288), .ZN(n38320) );
  AND2_X1 U42476 ( .A1(n8256), .A2(n40874), .ZN(n40535) );
  NAND2_X1 U42477 ( .A1(n40535), .A2(n39962), .ZN(n38353) );
  INV_X1 U42478 ( .A(n40874), .ZN(n40863) );
  NAND3_X1 U42479 ( .A1(n38323), .A2(n38338), .A3(n38330), .ZN(n38324) );
  INV_X1 U42480 ( .A(n38328), .ZN(n38333) );
  OAI22_X1 U42481 ( .A1(n6614), .A2(n38336), .B1(n38335), .B2(n38334), .ZN(
        n38344) );
  OAI22_X1 U42482 ( .A1(n35889), .A2(n38339), .B1(n38338), .B2(n38337), .ZN(
        n38343) );
  NOR2_X1 U42483 ( .A1(n38341), .A2(n38340), .ZN(n38342) );
  OAI21_X1 U42484 ( .B1(n40863), .B2(n39962), .A(n40862), .ZN(n38352) );
  INV_X1 U42485 ( .A(n40868), .ZN(n40856) );
  AND2_X1 U42486 ( .A1(n40856), .A2(n40869), .ZN(n40537) );
  INV_X1 U42487 ( .A(n40862), .ZN(n40533) );
  NAND2_X1 U42488 ( .A1(n40872), .A2(n40876), .ZN(n39969) );
  AND2_X1 U42489 ( .A1(n39969), .A2(n38355), .ZN(n38359) );
  NAND2_X1 U42490 ( .A1(n40874), .A2(n40868), .ZN(n39746) );
  NOR2_X1 U42491 ( .A1(n39746), .A2(n39962), .ZN(n40528) );
  NOR2_X1 U42492 ( .A1(n40528), .A2(n38356), .ZN(n38358) );
  NOR2_X1 U42493 ( .A1(n40874), .A2(n40862), .ZN(n39747) );
  NAND4_X2 U42494 ( .A1(n38359), .A2(n38360), .A3(n38358), .A4(n38357), .ZN(
        n44016) );
  XNOR2_X1 U42495 ( .A(n44016), .B(n44209), .ZN(n42870) );
  XNOR2_X1 U42496 ( .A(n44512), .B(n42870), .ZN(n42222) );
  AND2_X1 U42497 ( .A1(n41082), .A2(n41079), .ZN(n39704) );
  NAND2_X1 U42498 ( .A1(n39704), .A2(n41085), .ZN(n38867) );
  OAI211_X1 U42499 ( .C1(n38362), .C2(n39709), .A(n38867), .B(n38361), .ZN(
        n38367) );
  INV_X1 U42500 ( .A(n39707), .ZN(n39711) );
  NAND2_X1 U42501 ( .A1(n38364), .A2(n39146), .ZN(n38365) );
  OAI21_X1 U42502 ( .B1(n39713), .B2(n41079), .A(n38869), .ZN(n39702) );
  NAND2_X1 U42503 ( .A1(n39700), .A2(n39140), .ZN(n38366) );
  NAND2_X1 U42504 ( .A1(n40450), .A2(n40446), .ZN(n40445) );
  INV_X1 U42505 ( .A(n38368), .ZN(n38369) );
  NAND2_X1 U42506 ( .A1(n38369), .A2(n40447), .ZN(n40440) );
  OAI21_X1 U42507 ( .B1(n2854), .B2(n40445), .A(n40440), .ZN(n38371) );
  NOR2_X1 U42508 ( .A1(n40396), .A2(n39979), .ZN(n40401) );
  NOR2_X1 U42509 ( .A1(n38371), .A2(n40401), .ZN(n38378) );
  NAND2_X1 U42510 ( .A1(n39737), .A2(n40458), .ZN(n38372) );
  NAND2_X1 U42511 ( .A1(n40447), .A2(n40403), .ZN(n40437) );
  NAND2_X1 U42512 ( .A1(n40403), .A2(n40453), .ZN(n38374) );
  NOR2_X1 U42513 ( .A1(n40437), .A2(n38374), .ZN(n38377) );
  NAND2_X1 U42514 ( .A1(n40456), .A2(n40403), .ZN(n38375) );
  OAI22_X1 U42515 ( .A1(n40397), .A2(n38375), .B1(n38374), .B2(n40458), .ZN(
        n38376) );
  OR2_X1 U42516 ( .A1(n40397), .A2(n37345), .ZN(n40395) );
  NAND2_X1 U42517 ( .A1(n2848), .A2(n40403), .ZN(n40442) );
  NOR2_X1 U42518 ( .A1(n40395), .A2(n40442), .ZN(n39740) );
  XNOR2_X1 U42519 ( .A(n44006), .B(n51408), .ZN(n38399) );
  INV_X1 U42520 ( .A(n38782), .ZN(n38379) );
  NAND2_X1 U42521 ( .A1(n40125), .A2(n38379), .ZN(n40200) );
  NAND2_X1 U42522 ( .A1(n51233), .A2(n584), .ZN(n40201) );
  INV_X1 U42523 ( .A(n40119), .ZN(n40111) );
  NOR2_X1 U42524 ( .A1(n51325), .A2(n40120), .ZN(n38773) );
  NAND2_X1 U42525 ( .A1(n51325), .A2(n51352), .ZN(n40198) );
  XNOR2_X1 U42526 ( .A(n40120), .B(n51352), .ZN(n38381) );
  NAND4_X1 U42527 ( .A1(n40198), .A2(n38381), .A3(n40118), .A4(n40119), .ZN(
        n38382) );
  NAND2_X1 U42528 ( .A1(n38383), .A2(n38382), .ZN(n38387) );
  NAND2_X1 U42529 ( .A1(n40110), .A2(n38782), .ZN(n38784) );
  OAI21_X1 U42531 ( .B1(n507), .B2(n40120), .A(n40118), .ZN(n38385) );
  NOR2_X1 U42532 ( .A1(n40113), .A2(n40125), .ZN(n38384) );
  AOI22_X1 U42533 ( .A1(n39552), .A2(n38385), .B1(n38777), .B2(n38384), .ZN(
        n38386) );
  NOR2_X1 U42536 ( .A1(n40494), .A2(n41054), .ZN(n38392) );
  OR2_X1 U42537 ( .A1(n38389), .A2(n41065), .ZN(n40497) );
  NOR2_X1 U42538 ( .A1(n40513), .A2(n39129), .ZN(n38390) );
  AOI22_X1 U42539 ( .A1(n38392), .A2(n40497), .B1(n38391), .B2(n38390), .ZN(
        n38398) );
  NOR2_X1 U42540 ( .A1(n41064), .A2(n39129), .ZN(n38393) );
  OAI211_X1 U42541 ( .C1(n40499), .C2(n38393), .A(n41065), .B(n39604), .ZN(
        n38397) );
  OAI22_X1 U42542 ( .A1(n41064), .A2(n40512), .B1(n40493), .B2(n41047), .ZN(
        n38394) );
  NAND2_X1 U42543 ( .A1(n38394), .A2(n41055), .ZN(n38396) );
  OAI21_X1 U42544 ( .B1(n41052), .B2(n41063), .A(n41051), .ZN(n38395) );
  XNOR2_X1 U42547 ( .A(n45390), .B(n38399), .ZN(n40642) );
  AND2_X1 U42548 ( .A1(n660), .A2(n48273), .ZN(n44427) );
  NOR2_X1 U42549 ( .A1(n39929), .A2(n38401), .ZN(n38406) );
  INV_X1 U42551 ( .A(n40682), .ZN(n38402) );
  AOI211_X1 U42552 ( .C1(n38404), .C2(n40685), .A(n39673), .B(n40684), .ZN(
        n38405) );
  NAND2_X1 U42553 ( .A1(n40682), .A2(n40684), .ZN(n40679) );
  INV_X1 U42555 ( .A(n39680), .ZN(n39325) );
  OAI21_X1 U42556 ( .B1(n40693), .B2(n38406), .A(n39325), .ZN(n38407) );
  AND2_X1 U42557 ( .A1(n39674), .A2(n40672), .ZN(n39324) );
  INV_X1 U42558 ( .A(n39324), .ZN(n38414) );
  NAND2_X1 U42559 ( .A1(n40684), .A2(n39673), .ZN(n39927) );
  INV_X1 U42560 ( .A(n40690), .ZN(n38413) );
  INV_X1 U42561 ( .A(n38410), .ZN(n39321) );
  NAND2_X1 U42562 ( .A1(n6884), .A2(n38416), .ZN(n39670) );
  AND2_X1 U42563 ( .A1(n39103), .A2(n40003), .ZN(n40013) );
  NAND3_X1 U42564 ( .A1(n40013), .A2(n40002), .A3(n40015), .ZN(n38417) );
  AND3_X1 U42565 ( .A1(n38418), .A2(n39670), .A3(n38417), .ZN(n38435) );
  NAND2_X1 U42566 ( .A1(n38428), .A2(n51297), .ZN(n40001) );
  INV_X1 U42567 ( .A(n40001), .ZN(n38419) );
  NAND3_X1 U42568 ( .A1(n40013), .A2(n38424), .A3(n38419), .ZN(n38422) );
  INV_X1 U42569 ( .A(n39095), .ZN(n38420) );
  NAND3_X1 U42570 ( .A1(n39094), .A2(n39668), .A3(n38420), .ZN(n38421) );
  AND3_X1 U42571 ( .A1(n38423), .A2(n38422), .A3(n38421), .ZN(n38434) );
  NAND2_X1 U42572 ( .A1(n39101), .A2(n38424), .ZN(n39998) );
  INV_X1 U42573 ( .A(n39998), .ZN(n38425) );
  NAND2_X1 U42575 ( .A1(n40009), .A2(n38428), .ZN(n38431) );
  OAI21_X1 U42576 ( .B1(n39103), .B2(n39101), .A(n38429), .ZN(n38430) );
  NAND4_X1 U42577 ( .A1(n38431), .A2(n38430), .A3(n40003), .A4(n40014), .ZN(
        n38432) );
  AND2_X1 U42580 ( .A1(n39899), .A2(n51377), .ZN(n39914) );
  INV_X1 U42582 ( .A(n38438), .ZN(n38439) );
  NAND3_X1 U42583 ( .A1(n38440), .A2(n39565), .A3(n38439), .ZN(n38443) );
  NAND3_X1 U42584 ( .A1(n39915), .A2(n38441), .A3(n39565), .ZN(n38442) );
  AND3_X1 U42585 ( .A1(n38444), .A2(n38443), .A3(n38442), .ZN(n38463) );
  NAND2_X1 U42586 ( .A1(n39907), .A2(n38445), .ZN(n39790) );
  NAND3_X1 U42587 ( .A1(n38447), .A2(n38446), .A3(n39790), .ZN(n38462) );
  INV_X1 U42588 ( .A(n39785), .ZN(n39569) );
  NAND2_X1 U42589 ( .A1(n39565), .A2(n39908), .ZN(n38454) );
  INV_X1 U42590 ( .A(n39789), .ZN(n38451) );
  NAND2_X1 U42591 ( .A1(n39908), .A2(n51377), .ZN(n38450) );
  NAND3_X1 U42592 ( .A1(n38454), .A2(n38451), .A3(n38450), .ZN(n38452) );
  AND2_X1 U42593 ( .A1(n38452), .A2(n38453), .ZN(n38461) );
  NOR3_X1 U42594 ( .A1(n39785), .A2(n39565), .A3(n39912), .ZN(n38459) );
  NAND2_X1 U42595 ( .A1(n39906), .A2(n39899), .ZN(n39904) );
  INV_X1 U42596 ( .A(n39904), .ZN(n38458) );
  INV_X1 U42597 ( .A(n38454), .ZN(n38457) );
  INV_X1 U42598 ( .A(n38455), .ZN(n38456) );
  AOI22_X1 U42599 ( .A1(n38459), .A2(n38458), .B1(n38457), .B2(n38456), .ZN(
        n38460) );
  OAI22_X1 U42600 ( .A1(n38481), .A2(n36115), .B1(n38465), .B2(n38464), .ZN(
        n38470) );
  NOR2_X1 U42601 ( .A1(n38468), .A2(n38467), .ZN(n38469) );
  AOI21_X1 U42602 ( .B1(n38470), .B2(n38478), .A(n38469), .ZN(n38489) );
  AOI21_X1 U42603 ( .B1(n38473), .B2(n38472), .A(n38471), .ZN(n38474) );
  NAND2_X1 U42604 ( .A1(n38484), .A2(n38477), .ZN(n38482) );
  NAND2_X1 U42605 ( .A1(n38478), .A2(n1950), .ZN(n38479) );
  NAND4_X1 U42606 ( .A1(n38482), .A2(n38481), .A3(n38480), .A4(n38479), .ZN(
        n38488) );
  INV_X1 U42607 ( .A(n38482), .ZN(n38487) );
  NOR2_X1 U42608 ( .A1(n38484), .A2(n38483), .ZN(n38486) );
  INV_X1 U42609 ( .A(n41323), .ZN(n38511) );
  NAND2_X1 U42610 ( .A1(n38493), .A2(n38492), .ZN(n38498) );
  AOI21_X1 U42611 ( .B1(n38498), .B2(n38497), .A(n38496), .ZN(n38499) );
  NAND2_X1 U42612 ( .A1(n38502), .A2(n38501), .ZN(n38509) );
  OAI21_X1 U42613 ( .B1(n38505), .B2(n38504), .A(n38503), .ZN(n38507) );
  NAND2_X1 U42614 ( .A1(n38507), .A2(n38506), .ZN(n38508) );
  OAI22_X1 U42615 ( .A1(n38514), .A2(n37430), .B1(n38513), .B2(n38512), .ZN(
        n38516) );
  NOR2_X1 U42616 ( .A1(n37430), .A2(n38517), .ZN(n38519) );
  OAI21_X1 U42617 ( .B1(n38520), .B2(n38519), .A(n38518), .ZN(n38525) );
  NAND4_X1 U42618 ( .A1(n38526), .A2(n38525), .A3(n38524), .A4(n38523), .ZN(
        n38540) );
  OAI211_X1 U42619 ( .C1(n38535), .C2(n38534), .A(n38533), .B(n38532), .ZN(
        n38536) );
  OAI211_X1 U42620 ( .C1(n51363), .C2(n38538), .A(n38537), .B(n38536), .ZN(
        n38539) );
  NAND3_X1 U42621 ( .A1(n38544), .A2(n38543), .A3(n31355), .ZN(n38546) );
  OAI22_X1 U42622 ( .A1(n38555), .A2(n6734), .B1(n38553), .B2(n38552), .ZN(
        n38556) );
  OAI21_X1 U42623 ( .B1(n38558), .B2(n38557), .A(n38556), .ZN(n38559) );
  NOR2_X1 U42624 ( .A1(n41328), .A2(n41902), .ZN(n41318) );
  INV_X1 U42625 ( .A(n41318), .ZN(n38580) );
  OAI22_X1 U42626 ( .A1(n38567), .A2(n33062), .B1(n591), .B2(n1764), .ZN(
        n38563) );
  MUX2_X1 U42627 ( .A(n38564), .B(n38563), .S(n38562), .Z(n38579) );
  NOR2_X1 U42628 ( .A1(n38565), .A2(n33062), .ZN(n38568) );
  AOI22_X1 U42629 ( .A1(n38568), .A2(n38567), .B1(n38566), .B2(n6869), .ZN(
        n38578) );
  OAI22_X1 U42630 ( .A1(n38572), .A2(n38571), .B1(n38570), .B2(n38569), .ZN(
        n38574) );
  NAND2_X1 U42631 ( .A1(n38576), .A2(n591), .ZN(n38577) );
  NAND3_X1 U42632 ( .A1(n39814), .A2(n38580), .A3(n40730), .ZN(n38602) );
  NAND2_X1 U42633 ( .A1(n38582), .A2(n38581), .ZN(n38600) );
  AND2_X1 U42634 ( .A1(n38584), .A2(n38583), .ZN(n38597) );
  NAND2_X1 U42635 ( .A1(n38599), .A2(n38585), .ZN(n38586) );
  NOR2_X1 U42636 ( .A1(n51429), .A2(n38586), .ZN(n38588) );
  AOI22_X1 U42637 ( .A1(n38589), .A2(n38588), .B1(n38593), .B2(n38592), .ZN(
        n38595) );
  OAI211_X1 U42638 ( .C1(n38593), .C2(n38592), .A(n38591), .B(n38590), .ZN(
        n38594) );
  OAI211_X1 U42639 ( .C1(n38597), .C2(n38596), .A(n38595), .B(n38594), .ZN(
        n38598) );
  OAI211_X1 U42640 ( .C1(n40729), .C2(n40373), .A(n41326), .B(n40732), .ZN(
        n38601) );
  NOR2_X1 U42641 ( .A1(n41328), .A2(n41316), .ZN(n38606) );
  INV_X1 U42642 ( .A(n41324), .ZN(n38603) );
  NAND2_X1 U42643 ( .A1(n38603), .A2(n52214), .ZN(n39820) );
  NAND3_X1 U42644 ( .A1(n41902), .A2(n41319), .A3(n41332), .ZN(n40724) );
  NAND2_X1 U42645 ( .A1(n41320), .A2(n41328), .ZN(n38604) );
  AND3_X1 U42646 ( .A1(n39820), .A2(n40724), .A3(n38605), .ZN(n38609) );
  NAND2_X1 U42647 ( .A1(n38607), .A2(n38606), .ZN(n38608) );
  INV_X1 U42648 ( .A(n39839), .ZN(n38611) );
  INV_X1 U42649 ( .A(n41142), .ZN(n38614) );
  INV_X1 U42650 ( .A(n38612), .ZN(n41141) );
  AOI22_X1 U42651 ( .A1(n38614), .A2(n41141), .B1(n38613), .B2(n52083), .ZN(
        n38625) );
  INV_X1 U42652 ( .A(n40382), .ZN(n38619) );
  NAND2_X1 U42653 ( .A1(n38621), .A2(n682), .ZN(n38623) );
  XNOR2_X1 U42654 ( .A(n44198), .B(n38626), .ZN(n38752) );
  NAND3_X1 U42655 ( .A1(n38638), .A2(n38637), .A3(n35310), .ZN(n38639) );
  NAND2_X1 U42656 ( .A1(n38640), .A2(n38639), .ZN(n38642) );
  NAND2_X1 U42657 ( .A1(n38642), .A2(n38641), .ZN(n38643) );
  NAND2_X1 U42659 ( .A1(n39418), .A2(n38647), .ZN(n38648) );
  NAND2_X1 U42660 ( .A1(n38648), .A2(n39414), .ZN(n38657) );
  INV_X1 U42661 ( .A(n38649), .ZN(n38650) );
  AOI22_X1 U42662 ( .A1(n38938), .A2(n38650), .B1(n39422), .B2(n39426), .ZN(
        n38656) );
  INV_X1 U42663 ( .A(n39423), .ZN(n39201) );
  OAI21_X1 U42664 ( .B1(n38951), .B2(n39206), .A(n39201), .ZN(n38652) );
  OAI21_X1 U42666 ( .B1(n5151), .B2(n39410), .A(n39201), .ZN(n38653) );
  NAND3_X1 U42667 ( .A1(n38949), .A2(n39204), .A3(n38653), .ZN(n38654) );
  NAND2_X1 U42669 ( .A1(n38661), .A2(n38660), .ZN(n38683) );
  INV_X1 U42670 ( .A(n38662), .ZN(n38669) );
  INV_X1 U42671 ( .A(n38663), .ZN(n38675) );
  NAND2_X1 U42672 ( .A1(n700), .A2(n38664), .ZN(n39174) );
  NAND2_X1 U42673 ( .A1(n38664), .A2(n420), .ZN(n38665) );
  AOI21_X1 U42674 ( .B1(n38669), .B2(n39166), .A(n38668), .ZN(n38682) );
  AND2_X1 U42676 ( .A1(n38673), .A2(n38674), .ZN(n38681) );
  NAND4_X1 U42677 ( .A1(n38679), .A2(n419), .A3(n38678), .A4(n38677), .ZN(
        n38680) );
  NAND4_X2 U42678 ( .A1(n38682), .A2(n38680), .A3(n38683), .A4(n38681), .ZN(
        n41354) );
  NOR2_X1 U42679 ( .A1(n551), .A2(n39273), .ZN(n38685) );
  OAI21_X1 U42680 ( .B1(n39265), .B2(n38685), .A(n39259), .ZN(n38688) );
  NAND2_X1 U42681 ( .A1(n39016), .A2(n39262), .ZN(n38692) );
  INV_X1 U42682 ( .A(n39271), .ZN(n39013) );
  NAND3_X1 U42683 ( .A1(n38689), .A2(n39274), .A3(n551), .ZN(n38690) );
  MUX2_X1 U42686 ( .A(n38708), .B(n38698), .S(n39243), .Z(n38713) );
  OAI22_X1 U42687 ( .A1(n39227), .A2(n38702), .B1(n38701), .B2(n39221), .ZN(
        n38703) );
  NAND2_X1 U42688 ( .A1(n38703), .A2(n38704), .ZN(n38712) );
  NAND3_X1 U42689 ( .A1(n38706), .A2(n3874), .A3(n38704), .ZN(n38707) );
  NAND2_X1 U42690 ( .A1(n38710), .A2(n51736), .ZN(n38711) );
  INV_X1 U42691 ( .A(n41354), .ZN(n38740) );
  NAND2_X1 U42692 ( .A1(n8123), .A2(n52088), .ZN(n39889) );
  OAI211_X1 U42693 ( .C1(n6469), .C2(n41352), .A(n41345), .B(n39889), .ZN(
        n38714) );
  OAI21_X1 U42694 ( .B1(n41358), .B2(n40749), .A(n38714), .ZN(n38739) );
  NAND2_X1 U42695 ( .A1(n38715), .A2(n38716), .ZN(n38719) );
  INV_X1 U42696 ( .A(n38716), .ZN(n38717) );
  AOI21_X1 U42697 ( .B1(n38725), .B2(n38728), .A(n38724), .ZN(n38726) );
  OAI22_X1 U42698 ( .A1(n38734), .A2(n39300), .B1(n6748), .B2(n7772), .ZN(
        n38729) );
  AND2_X1 U42699 ( .A1(n38728), .A2(n38727), .ZN(n39298) );
  OAI21_X1 U42700 ( .B1(n38730), .B2(n38729), .A(n39298), .ZN(n38738) );
  INV_X1 U42701 ( .A(n39295), .ZN(n38737) );
  NAND3_X1 U42702 ( .A1(n39299), .A2(n7772), .A3(n38731), .ZN(n38733) );
  NAND2_X1 U42703 ( .A1(n39307), .A2(n38733), .ZN(n38736) );
  NAND2_X1 U42704 ( .A1(n38739), .A2(n41355), .ZN(n38751) );
  AND2_X1 U42705 ( .A1(n40740), .A2(n52087), .ZN(n41350) );
  NAND2_X1 U42706 ( .A1(n41350), .A2(n41348), .ZN(n40745) );
  XNOR2_X1 U42707 ( .A(n41348), .B(n41352), .ZN(n38743) );
  NAND2_X1 U42708 ( .A1(n41355), .A2(n41360), .ZN(n38742) );
  NOR2_X1 U42709 ( .A1(n38740), .A2(n52088), .ZN(n38741) );
  NAND4_X1 U42710 ( .A1(n38743), .A2(n38742), .A3(n6469), .A4(n38741), .ZN(
        n38744) );
  OAI211_X1 U42711 ( .C1(n38745), .C2(n40359), .A(n40745), .B(n38744), .ZN(
        n38750) );
  NOR2_X1 U42712 ( .A1(n41355), .A2(n52087), .ZN(n40737) );
  NAND2_X1 U42713 ( .A1(n52088), .A2(n41352), .ZN(n41343) );
  INV_X1 U42714 ( .A(n41343), .ZN(n38746) );
  NOR2_X1 U42715 ( .A1(n41355), .A2(n6469), .ZN(n41338) );
  NAND2_X1 U42716 ( .A1(n41354), .A2(n52087), .ZN(n39633) );
  INV_X1 U42717 ( .A(n39633), .ZN(n40360) );
  NAND2_X1 U42718 ( .A1(n41338), .A2(n40360), .ZN(n38749) );
  XNOR2_X1 U42719 ( .A(n38752), .B(n43909), .ZN(n45130) );
  XNOR2_X1 U42720 ( .A(n45130), .B(n38753), .ZN(n41254) );
  NAND3_X1 U42721 ( .A1(n43335), .A2(n39576), .A3(n39609), .ZN(n38758) );
  NOR2_X1 U42722 ( .A1(n43323), .A2(n39576), .ZN(n38756) );
  NAND4_X1 U42723 ( .A1(n39614), .A2(n38756), .A3(n43327), .A4(n38759), .ZN(
        n38757) );
  OAI21_X1 U42724 ( .B1(n40807), .B2(n38763), .A(n609), .ZN(n38767) );
  AND2_X1 U42725 ( .A1(n51357), .A2(n39576), .ZN(n40797) );
  NAND2_X1 U42726 ( .A1(n43323), .A2(n38764), .ZN(n40795) );
  INV_X1 U42727 ( .A(n40795), .ZN(n43326) );
  AOI22_X1 U42728 ( .A1(n43326), .A2(n38765), .B1(n40799), .B2(n43323), .ZN(
        n38766) );
  XNOR2_X1 U42729 ( .A(n42122), .B(n4482), .ZN(n43194) );
  INV_X1 U42730 ( .A(n38769), .ZN(n38770) );
  INV_X1 U42733 ( .A(n40194), .ZN(n38772) );
  NAND2_X1 U42734 ( .A1(n38772), .A2(n7239), .ZN(n40207) );
  OR2_X1 U42735 ( .A1(n40196), .A2(n40125), .ZN(n38775) );
  INV_X1 U42737 ( .A(n38773), .ZN(n38774) );
  NAND4_X1 U42738 ( .A1(n38775), .A2(n40194), .A3(n40192), .A4(n38774), .ZN(
        n38776) );
  AND2_X1 U42739 ( .A1(n38776), .A2(n40207), .ZN(n38791) );
  INV_X1 U42740 ( .A(n38777), .ZN(n38778) );
  OAI22_X1 U42741 ( .A1(n40192), .A2(n38778), .B1(n40204), .B2(n40111), .ZN(
        n38779) );
  AOI21_X1 U42742 ( .B1(n38781), .B2(n51325), .A(n39553), .ZN(n38788) );
  NOR2_X1 U42743 ( .A1(n38782), .A2(n584), .ZN(n38783) );
  NOR2_X1 U42744 ( .A1(n507), .A2(n38783), .ZN(n38787) );
  INV_X1 U42745 ( .A(n38784), .ZN(n40205) );
  NAND2_X1 U42746 ( .A1(n40205), .A2(n584), .ZN(n38786) );
  NAND2_X1 U42747 ( .A1(n40196), .A2(n40203), .ZN(n38785) );
  NAND4_X1 U42748 ( .A1(n38788), .A2(n38787), .A3(n38786), .A4(n38785), .ZN(
        n38789) );
  NAND4_X1 U42749 ( .A1(n40273), .A2(n40906), .A3(n40903), .A4(n2223), .ZN(
        n38793) );
  NAND3_X1 U42750 ( .A1(n38794), .A2(n40269), .A3(n38795), .ZN(n38798) );
  INV_X1 U42751 ( .A(n38795), .ZN(n38796) );
  NAND3_X1 U42752 ( .A1(n38796), .A2(n40906), .A3(n40903), .ZN(n38797) );
  OAI211_X1 U42753 ( .C1(n40906), .C2(n40900), .A(n38798), .B(n38797), .ZN(
        n38799) );
  NOR2_X1 U42754 ( .A1(n40273), .A2(n5072), .ZN(n40096) );
  OAI21_X1 U42755 ( .B1(n40910), .B2(n40903), .A(n40275), .ZN(n38803) );
  NOR2_X1 U42756 ( .A1(n2223), .A2(n40269), .ZN(n40904) );
  NAND2_X1 U42757 ( .A1(n40903), .A2(n40910), .ZN(n38800) );
  NAND2_X1 U42758 ( .A1(n38800), .A2(n40906), .ZN(n38802) );
  NAND4_X1 U42759 ( .A1(n38803), .A2(n40904), .A3(n38802), .A4(n38801), .ZN(
        n38804) );
  INV_X1 U42760 ( .A(n43635), .ZN(n43063) );
  XNOR2_X1 U42761 ( .A(n43194), .B(n51444), .ZN(n38864) );
  OR3_X1 U42762 ( .A1(n38805), .A2(n41792), .A3(n41796), .ZN(n38807) );
  AND2_X1 U42763 ( .A1(n43665), .A2(n40632), .ZN(n38809) );
  NAND3_X1 U42764 ( .A1(n38809), .A2(n41792), .A3(n41797), .ZN(n38806) );
  NAND4_X1 U42765 ( .A1(n38808), .A2(n51734), .A3(n38807), .A4(n38806), .ZN(
        n38811) );
  NAND2_X1 U42766 ( .A1(n51950), .A2(n41796), .ZN(n41801) );
  NAND4_X1 U42767 ( .A1(n38819), .A2(n51950), .A3(n40632), .A4(n41797), .ZN(
        n38813) );
  NAND3_X1 U42768 ( .A1(n38817), .A2(n43669), .A3(n51734), .ZN(n38818) );
  AND2_X1 U42769 ( .A1(n41793), .A2(n38818), .ZN(n38823) );
  INV_X1 U42770 ( .A(n38819), .ZN(n38821) );
  OAI211_X1 U42771 ( .C1(n41796), .C2(n43669), .A(n38821), .B(n38820), .ZN(
        n38822) );
  AND2_X1 U42773 ( .A1(n52095), .A2(n575), .ZN(n38828) );
  NAND3_X1 U42774 ( .A1(n39764), .A2(n38828), .A3(n39943), .ZN(n38825) );
  OAI21_X1 U42775 ( .B1(n39759), .B2(n39937), .A(n38825), .ZN(n38826) );
  INV_X1 U42777 ( .A(n38830), .ZN(n38833) );
  AND3_X1 U42779 ( .A1(n38835), .A2(n38836), .A3(n38834), .ZN(n38841) );
  NOR2_X1 U42780 ( .A1(n52095), .A2(n39754), .ZN(n38839) );
  NOR2_X1 U42781 ( .A1(n38838), .A2(n39943), .ZN(n39762) );
  XNOR2_X1 U42782 ( .A(n44189), .B(n45426), .ZN(n44325) );
  NAND3_X1 U42783 ( .A1(n39853), .A2(n38842), .A3(n40338), .ZN(n38846) );
  AND2_X1 U42784 ( .A1(n39857), .A2(n40342), .ZN(n40334) );
  NAND4_X1 U42785 ( .A1(n38843), .A2(n40329), .A3(n40341), .A4(n40330), .ZN(
        n38844) );
  AND2_X1 U42786 ( .A1(n39857), .A2(n40330), .ZN(n39850) );
  NAND3_X1 U42787 ( .A1(n39850), .A2(n39647), .A3(n40327), .ZN(n38847) );
  OAI21_X1 U42788 ( .B1(n38851), .B2(n40328), .A(n40329), .ZN(n38854) );
  INV_X1 U42789 ( .A(n40327), .ZN(n40343) );
  INV_X1 U42790 ( .A(n39850), .ZN(n38852) );
  NAND3_X1 U42791 ( .A1(n38852), .A2(n52101), .A3(n40338), .ZN(n38853) );
  NAND3_X1 U42792 ( .A1(n38854), .A2(n40343), .A3(n38853), .ZN(n38857) );
  NAND2_X1 U42793 ( .A1(n40328), .A2(n40340), .ZN(n39854) );
  OAI22_X1 U42794 ( .A1(n40337), .A2(n39647), .B1(n39854), .B2(n40330), .ZN(
        n38855) );
  NAND2_X1 U42795 ( .A1(n38855), .A2(n39862), .ZN(n38856) );
  XNOR2_X1 U42796 ( .A(n38860), .B(n38859), .ZN(n38861) );
  XNOR2_X1 U42797 ( .A(n51464), .B(n38861), .ZN(n38862) );
  XNOR2_X1 U42798 ( .A(n44325), .B(n38862), .ZN(n38863) );
  XNOR2_X1 U42799 ( .A(n38864), .B(n38863), .ZN(n38865) );
  XNOR2_X1 U42800 ( .A(n41254), .B(n38865), .ZN(n39093) );
  OAI21_X1 U42801 ( .B1(n41077), .B2(n38868), .A(n38875), .ZN(n38874) );
  NAND2_X1 U42802 ( .A1(n38869), .A2(n41085), .ZN(n39139) );
  INV_X1 U42803 ( .A(n39139), .ZN(n39143) );
  NAND3_X1 U42804 ( .A1(n39143), .A2(n38871), .A3(n41083), .ZN(n38873) );
  INV_X1 U42805 ( .A(n39145), .ZN(n38877) );
  NAND2_X1 U42806 ( .A1(n52108), .A2(n39712), .ZN(n39708) );
  AOI22_X1 U42807 ( .A1(n41087), .A2(n38875), .B1(n39143), .B2(n41077), .ZN(
        n38882) );
  OAI22_X1 U42808 ( .A1(n38877), .A2(n39140), .B1(n38876), .B2(n41083), .ZN(
        n38880) );
  AOI21_X1 U42809 ( .B1(n41085), .B2(n38878), .A(n41084), .ZN(n38879) );
  NAND2_X1 U42810 ( .A1(n38880), .A2(n38879), .ZN(n38881) );
  NOR2_X1 U42811 ( .A1(n41375), .A2(n40240), .ZN(n38899) );
  AND2_X1 U42812 ( .A1(n40960), .A2(n3775), .ZN(n38894) );
  NAND2_X1 U42813 ( .A1(n38894), .A2(n51853), .ZN(n38889) );
  NAND3_X1 U42814 ( .A1(n38887), .A2(n41380), .A3(n51853), .ZN(n38888) );
  OAI21_X1 U42815 ( .B1(n40917), .B2(n38889), .A(n38888), .ZN(n38892) );
  NAND4_X1 U42816 ( .A1(n41375), .A2(n40958), .A3(n676), .A4(n51394), .ZN(
        n38890) );
  OAI21_X1 U42817 ( .B1(n41372), .B2(n41374), .A(n38890), .ZN(n38891) );
  NOR2_X1 U42818 ( .A1(n38892), .A2(n38891), .ZN(n38904) );
  NAND3_X1 U42819 ( .A1(n41375), .A2(n40972), .A3(n40241), .ZN(n38897) );
  NAND3_X1 U42820 ( .A1(n38894), .A2(n40242), .A3(n51394), .ZN(n38895) );
  OAI211_X1 U42821 ( .C1(n38897), .C2(n40917), .A(n38896), .B(n38895), .ZN(
        n38898) );
  INV_X1 U42822 ( .A(n38898), .ZN(n38903) );
  INV_X1 U42823 ( .A(n40963), .ZN(n38901) );
  INV_X1 U42824 ( .A(n38899), .ZN(n38900) );
  AND2_X1 U42825 ( .A1(n40959), .A2(n40972), .ZN(n40966) );
  OAI211_X1 U42826 ( .C1(n38901), .C2(n51853), .A(n38900), .B(n40966), .ZN(
        n38902) );
  NAND2_X1 U42827 ( .A1(n41436), .A2(n41435), .ZN(n38906) );
  NAND4_X1 U42828 ( .A1(n38916), .A2(n40646), .A3(n40651), .A4(n38906), .ZN(
        n38908) );
  NAND3_X1 U42829 ( .A1(n41441), .A2(n41446), .A3(n5982), .ZN(n38907) );
  AND2_X1 U42830 ( .A1(n38908), .A2(n38907), .ZN(n38920) );
  INV_X1 U42831 ( .A(n40650), .ZN(n39766) );
  NOR2_X1 U42832 ( .A1(n39766), .A2(n40651), .ZN(n38911) );
  OAI22_X1 U42833 ( .A1(n41436), .A2(n41447), .B1(n38909), .B2(n7268), .ZN(
        n38910) );
  AOI21_X1 U42834 ( .B1(n40649), .B2(n38911), .A(n38910), .ZN(n38919) );
  INV_X1 U42835 ( .A(n38912), .ZN(n38914) );
  OAI21_X1 U42836 ( .B1(n39767), .B2(n41442), .A(n41436), .ZN(n38913) );
  OAI22_X1 U42837 ( .A1(n38914), .A2(n41434), .B1(n38913), .B2(n40651), .ZN(
        n38915) );
  OAI21_X1 U42838 ( .B1(n38916), .B2(n40646), .A(n38915), .ZN(n38918) );
  NOR2_X1 U42839 ( .A1(n40653), .A2(n41447), .ZN(n39776) );
  INV_X1 U42840 ( .A(n39776), .ZN(n38917) );
  NAND4_X2 U42841 ( .A1(n38920), .A2(n38919), .A3(n38918), .A4(n38917), .ZN(
        n45285) );
  XNOR2_X1 U42842 ( .A(n45285), .B(n3383), .ZN(n38936) );
  OAI21_X1 U42843 ( .B1(n38928), .B2(n41927), .A(n38921), .ZN(n38922) );
  NAND3_X1 U42844 ( .A1(n38924), .A2(n38923), .A3(n38922), .ZN(n38935) );
  NAND2_X1 U42845 ( .A1(n38926), .A2(n38925), .ZN(n38927) );
  NAND2_X1 U42846 ( .A1(n38927), .A2(n40250), .ZN(n38934) );
  NAND4_X1 U42847 ( .A1(n40251), .A2(n42202), .A3(n39543), .A4(n42205), .ZN(
        n38930) );
  NAND3_X1 U42848 ( .A1(n38928), .A2(n42202), .A3(n42205), .ZN(n38929) );
  AND2_X1 U42849 ( .A1(n38930), .A2(n38929), .ZN(n38933) );
  XNOR2_X1 U42850 ( .A(n38936), .B(n43170), .ZN(n42768) );
  XNOR2_X1 U42851 ( .A(n42768), .B(n52130), .ZN(n39091) );
  AOI22_X1 U42852 ( .A1(n38949), .A2(n39426), .B1(n38938), .B2(n38937), .ZN(
        n38939) );
  AND2_X1 U42853 ( .A1(n38941), .A2(n38940), .ZN(n39412) );
  OAI222_X1 U42854 ( .A1(n37907), .A2(n39207), .B1(n39411), .B2(n39429), .C1(
        n39422), .C2(n39430), .ZN(n38942) );
  NAND2_X1 U42855 ( .A1(n38949), .A2(n39414), .ZN(n38944) );
  NOR2_X1 U42856 ( .A1(n39417), .A2(n37900), .ZN(n39203) );
  NAND3_X1 U42857 ( .A1(n39203), .A2(n38946), .A3(n39207), .ZN(n39420) );
  INV_X1 U42859 ( .A(n38949), .ZN(n39424) );
  OAI21_X1 U42860 ( .B1(n38954), .B2(n38953), .A(n38952), .ZN(n38955) );
  NAND2_X1 U42861 ( .A1(n39198), .A2(n51322), .ZN(n38958) );
  AOI21_X1 U42862 ( .B1(n38959), .B2(n38958), .A(n39375), .ZN(n38970) );
  INV_X1 U42863 ( .A(n38960), .ZN(n38961) );
  NAND2_X1 U42864 ( .A1(n38961), .A2(n39381), .ZN(n38968) );
  XNOR2_X1 U42865 ( .A(n38963), .B(n39375), .ZN(n38964) );
  AOI22_X1 U42866 ( .A1(n39367), .A2(n38964), .B1(n38963), .B2(n38962), .ZN(
        n38967) );
  NAND3_X1 U42867 ( .A1(n39360), .A2(n39361), .A3(n39377), .ZN(n38965) );
  NAND4_X1 U42868 ( .A1(n38968), .A2(n38967), .A3(n38966), .A4(n38965), .ZN(
        n38969) );
  INV_X1 U42869 ( .A(n41693), .ZN(n41688) );
  NOR2_X1 U42870 ( .A1(n41702), .A2(n41688), .ZN(n39043) );
  INV_X1 U42871 ( .A(n38971), .ZN(n38976) );
  NAND2_X1 U42872 ( .A1(n2177), .A2(n473), .ZN(n38973) );
  AOI21_X1 U42873 ( .B1(n38976), .B2(n39486), .A(n38975), .ZN(n38990) );
  INV_X1 U42874 ( .A(n38977), .ZN(n38978) );
  OAI21_X1 U42875 ( .B1(n38979), .B2(n38978), .A(n39488), .ZN(n38989) );
  INV_X1 U42876 ( .A(n38980), .ZN(n38986) );
  INV_X1 U42877 ( .A(n38981), .ZN(n38985) );
  OAI21_X1 U42878 ( .B1(n38986), .B2(n38985), .A(n38984), .ZN(n38987) );
  NAND3_X1 U42879 ( .A1(n39400), .A2(n3735), .A3(n39395), .ZN(n38992) );
  AND3_X1 U42880 ( .A1(n38994), .A2(n38993), .A3(n38992), .ZN(n39006) );
  NAND2_X1 U42881 ( .A1(n39397), .A2(n38998), .ZN(n39001) );
  NAND3_X1 U42882 ( .A1(n39402), .A2(n39003), .A3(n38999), .ZN(n39000) );
  NAND3_X1 U42883 ( .A1(n39266), .A2(n39008), .A3(n39007), .ZN(n39010) );
  NAND4_X1 U42884 ( .A1(n39258), .A2(n39014), .A3(n39273), .A4(n39019), .ZN(
        n39009) );
  NAND3_X1 U42885 ( .A1(n39016), .A2(n39259), .A3(n39270), .ZN(n39018) );
  OAI211_X1 U42886 ( .C1(n39020), .C2(n39019), .A(n39018), .B(n39017), .ZN(
        n39021) );
  INV_X1 U42887 ( .A(n39021), .ZN(n39022) );
  MUX2_X1 U42888 ( .A(n39448), .B(n39032), .S(n39035), .Z(n39460) );
  NOR2_X1 U42889 ( .A1(n39445), .A2(n467), .ZN(n39029) );
  AOI21_X1 U42890 ( .B1(n39030), .B2(n39027), .A(n39029), .ZN(n39040) );
  NAND3_X1 U42891 ( .A1(n39033), .A2(n39032), .A3(n39031), .ZN(n39038) );
  OAI211_X1 U42892 ( .C1(n39036), .C2(n39035), .A(n39034), .B(n39450), .ZN(
        n39037) );
  AND2_X1 U42893 ( .A1(n39038), .A2(n39037), .ZN(n39039) );
  OAI21_X1 U42894 ( .B1(n41690), .B2(n41693), .A(n41697), .ZN(n39042) );
  INV_X1 U42895 ( .A(n41709), .ZN(n39877) );
  AND2_X1 U42896 ( .A1(n41693), .A2(n5475), .ZN(n41705) );
  INV_X1 U42897 ( .A(n41705), .ZN(n41170) );
  INV_X1 U42898 ( .A(n41689), .ZN(n39871) );
  NOR2_X1 U42900 ( .A1(n39043), .A2(n41166), .ZN(n39050) );
  INV_X1 U42901 ( .A(n41704), .ZN(n39870) );
  AND2_X1 U42902 ( .A1(n41690), .A2(n41621), .ZN(n39044) );
  MUX2_X1 U42903 ( .A(n39870), .B(n39044), .S(n41702), .Z(n39049) );
  NAND2_X1 U42904 ( .A1(n41690), .A2(n41691), .ZN(n39874) );
  INV_X1 U42905 ( .A(n39874), .ZN(n39045) );
  NAND3_X1 U42906 ( .A1(n41707), .A2(n41697), .A3(n39045), .ZN(n39047) );
  NAND3_X1 U42907 ( .A1(n41702), .A2(n41615), .A3(n41706), .ZN(n41711) );
  INV_X1 U42908 ( .A(n41699), .ZN(n39046) );
  AOI21_X1 U42909 ( .B1(n39050), .B2(n39049), .A(n39048), .ZN(n39051) );
  INV_X1 U42910 ( .A(n40295), .ZN(n39052) );
  OAI21_X1 U42911 ( .B1(n42061), .B2(n42441), .A(n39052), .ZN(n39056) );
  NAND2_X1 U42912 ( .A1(n39052), .A2(n42049), .ZN(n39055) );
  INV_X1 U42913 ( .A(n41482), .ZN(n39053) );
  NAND2_X1 U42914 ( .A1(n39053), .A2(n40295), .ZN(n39054) );
  XNOR2_X1 U42916 ( .A(n42441), .B(n679), .ZN(n39059) );
  NAND2_X1 U42917 ( .A1(n40295), .A2(n679), .ZN(n39058) );
  AND2_X1 U42918 ( .A1(n596), .A2(n480), .ZN(n42039) );
  AOI21_X1 U42919 ( .B1(n41481), .B2(n42049), .A(n42039), .ZN(n39057) );
  NAND4_X1 U42920 ( .A1(n39059), .A2(n39058), .A3(n39057), .A4(n42043), .ZN(
        n39060) );
  NAND2_X1 U42922 ( .A1(n40051), .A2(n42061), .ZN(n42041) );
  NAND2_X1 U42923 ( .A1(n40295), .A2(n42061), .ZN(n39062) );
  NAND2_X1 U42924 ( .A1(n39063), .A2(n41481), .ZN(n39066) );
  NOR2_X1 U42925 ( .A1(n39064), .A2(n42049), .ZN(n39065) );
  NOR2_X1 U42926 ( .A1(n42441), .A2(n41480), .ZN(n40292) );
  INV_X1 U42927 ( .A(n40292), .ZN(n41487) );
  OAI21_X1 U42929 ( .B1(n7488), .B2(n40836), .A(n39691), .ZN(n39070) );
  OAI21_X1 U42930 ( .B1(n51990), .B2(n51455), .A(n40839), .ZN(n39069) );
  NOR2_X1 U42931 ( .A1(n39070), .A2(n39069), .ZN(n39073) );
  INV_X1 U42932 ( .A(n39693), .ZN(n40826) );
  OAI21_X1 U42933 ( .B1(n39512), .B2(n40826), .A(n39071), .ZN(n39072) );
  AOI22_X1 U42934 ( .A1(n39074), .A2(n40840), .B1(n40835), .B2(n39513), .ZN(
        n39088) );
  NAND2_X1 U42935 ( .A1(n39512), .A2(n40815), .ZN(n40830) );
  OAI21_X1 U42938 ( .B1(n40838), .B2(n52151), .A(n40822), .ZN(n39076) );
  NAND3_X1 U42939 ( .A1(n39692), .A2(n40839), .A3(n39076), .ZN(n39081) );
  OR2_X1 U42940 ( .A1(n40818), .A2(n39077), .ZN(n39690) );
  INV_X1 U42941 ( .A(n39690), .ZN(n39079) );
  NAND2_X1 U42942 ( .A1(n40823), .A2(n52151), .ZN(n40816) );
  INV_X1 U42943 ( .A(n40816), .ZN(n39078) );
  INV_X1 U42946 ( .A(n39082), .ZN(n39087) );
  NAND3_X1 U42947 ( .A1(n39512), .A2(n40823), .A3(n40815), .ZN(n39083) );
  OAI21_X1 U42948 ( .B1(n39512), .B2(n40823), .A(n39083), .ZN(n39085) );
  INV_X1 U42949 ( .A(n39691), .ZN(n39084) );
  NAND2_X1 U42950 ( .A1(n39085), .A2(n39084), .ZN(n39086) );
  XNOR2_X1 U42951 ( .A(n42170), .B(n842), .ZN(n39090) );
  XNOR2_X1 U42952 ( .A(n43522), .B(n39090), .ZN(n43811) );
  XNOR2_X1 U42953 ( .A(n39091), .B(n43811), .ZN(n39092) );
  XNOR2_X1 U42954 ( .A(n39093), .B(n39092), .ZN(n39812) );
  AND2_X1 U42955 ( .A1(n40018), .A2(n39998), .ZN(n39109) );
  INV_X1 U42956 ( .A(n39094), .ZN(n39664) );
  OAI21_X1 U42957 ( .B1(n40003), .B2(n40015), .A(n39664), .ZN(n39096) );
  NAND2_X1 U42958 ( .A1(n39096), .A2(n39095), .ZN(n39108) );
  INV_X1 U42959 ( .A(n39101), .ZN(n39098) );
  NAND2_X1 U42960 ( .A1(n39101), .A2(n51297), .ZN(n39102) );
  OAI211_X1 U42961 ( .C1(n39098), .C2(n39103), .A(n40014), .B(n39102), .ZN(
        n39105) );
  INV_X1 U42962 ( .A(n39104), .ZN(n39997) );
  NAND2_X1 U42963 ( .A1(n39105), .A2(n39997), .ZN(n39106) );
  XNOR2_X1 U42964 ( .A(n44373), .B(n42327), .ZN(n39125) );
  OR2_X1 U42965 ( .A1(n52094), .A2(n39751), .ZN(n39940) );
  OAI211_X1 U42966 ( .C1(n2386), .C2(n39940), .A(n39942), .B(n39111), .ZN(
        n39110) );
  NAND2_X1 U42967 ( .A1(n39943), .A2(n52094), .ZN(n39954) );
  INV_X1 U42968 ( .A(n39954), .ZN(n39755) );
  AND2_X1 U42969 ( .A1(n39754), .A2(n575), .ZN(n39957) );
  INV_X1 U42970 ( .A(n39111), .ZN(n39951) );
  NAND3_X1 U42971 ( .A1(n39951), .A2(n39938), .A3(n39112), .ZN(n39113) );
  NAND2_X1 U42972 ( .A1(n40422), .A2(n41275), .ZN(n40429) );
  NAND2_X1 U42973 ( .A1(n40429), .A2(n41035), .ZN(n39116) );
  NOR2_X1 U42974 ( .A1(n52193), .A2(n40417), .ZN(n39726) );
  NAND2_X1 U42975 ( .A1(n39116), .A2(n39726), .ZN(n39124) );
  OR2_X1 U42976 ( .A1(n41276), .A2(n8291), .ZN(n39117) );
  NOR2_X1 U42977 ( .A1(n39117), .A2(n5324), .ZN(n39118) );
  INV_X1 U42978 ( .A(n41039), .ZN(n41280) );
  INV_X1 U42979 ( .A(n41287), .ZN(n41040) );
  INV_X1 U42980 ( .A(n39117), .ZN(n40428) );
  AOI22_X1 U42981 ( .A1(n39118), .A2(n41280), .B1(n41040), .B2(n40428), .ZN(
        n39123) );
  NAND2_X1 U42982 ( .A1(n41287), .A2(n41286), .ZN(n39120) );
  XNOR2_X1 U42983 ( .A(n40417), .B(n41275), .ZN(n39119) );
  AOI22_X1 U42984 ( .A1(n39120), .A2(n41280), .B1(n41040), .B2(n39119), .ZN(
        n39122) );
  NOR2_X1 U42985 ( .A1(n41039), .A2(n41276), .ZN(n39727) );
  NAND2_X1 U42986 ( .A1(n39121), .A2(n39727), .ZN(n41295) );
  INV_X1 U42987 ( .A(n40494), .ZN(n39127) );
  NAND2_X1 U42988 ( .A1(n51348), .A2(n39129), .ZN(n40511) );
  NAND2_X1 U42989 ( .A1(n41049), .A2(n40500), .ZN(n39126) );
  NAND2_X1 U42990 ( .A1(n6392), .A2(n41057), .ZN(n39603) );
  NOR2_X1 U42991 ( .A1(n39603), .A2(n40506), .ZN(n39128) );
  NOR2_X1 U42992 ( .A1(n41045), .A2(n39128), .ZN(n39136) );
  NAND3_X1 U42993 ( .A1(n40501), .A2(n39129), .A3(n41049), .ZN(n39135) );
  NAND2_X1 U42994 ( .A1(n41049), .A2(n41054), .ZN(n39130) );
  NAND2_X1 U42995 ( .A1(n39131), .A2(n39130), .ZN(n39133) );
  INV_X1 U42996 ( .A(n40513), .ZN(n39132) );
  NAND2_X1 U42997 ( .A1(n39133), .A2(n39132), .ZN(n39134) );
  NOR2_X1 U42998 ( .A1(n39712), .A2(n41082), .ZN(n39138) );
  NOR2_X1 U42999 ( .A1(n39139), .A2(n39138), .ZN(n41086) );
  OR2_X1 U43000 ( .A1(n39141), .A2(n39140), .ZN(n39142) );
  NAND2_X1 U43001 ( .A1(n41086), .A2(n39142), .ZN(n39153) );
  AOI21_X1 U43002 ( .B1(n39143), .B2(n39713), .A(n41087), .ZN(n39152) );
  NOR2_X1 U43003 ( .A1(n41085), .A2(n39144), .ZN(n41073) );
  NAND2_X1 U43004 ( .A1(n39145), .A2(n41073), .ZN(n39151) );
  NOR2_X1 U43006 ( .A1(n41085), .A2(n41082), .ZN(n39147) );
  AOI21_X1 U43007 ( .B1(n41084), .B2(n39147), .A(n8316), .ZN(n39148) );
  XNOR2_X2 U43009 ( .A(n43723), .B(n44501), .ZN(n43048) );
  XNOR2_X1 U43010 ( .A(n39154), .B(n43048), .ZN(n44975) );
  INV_X1 U43011 ( .A(n8759), .ZN(n40654) );
  NOR2_X1 U43012 ( .A1(n40654), .A2(n40655), .ZN(n39156) );
  INV_X1 U43013 ( .A(n5982), .ZN(n39155) );
  AOI22_X1 U43014 ( .A1(n39156), .A2(n40651), .B1(n39774), .B2(n39155), .ZN(
        n39165) );
  NAND3_X1 U43015 ( .A1(n40643), .A2(n39157), .A3(n40652), .ZN(n39159) );
  NOR2_X1 U43016 ( .A1(n7268), .A2(n41436), .ZN(n41450) );
  INV_X1 U43017 ( .A(n41450), .ZN(n39158) );
  AND2_X1 U43018 ( .A1(n39159), .A2(n39158), .ZN(n39164) );
  NOR2_X1 U43019 ( .A1(n40651), .A2(n41433), .ZN(n41451) );
  NAND2_X1 U43022 ( .A1(n41451), .A2(n39161), .ZN(n39163) );
  INV_X1 U43023 ( .A(n41430), .ZN(n39772) );
  NAND3_X1 U43024 ( .A1(n40653), .A2(n39772), .A3(n41435), .ZN(n39162) );
  NAND2_X1 U43025 ( .A1(n39170), .A2(n39169), .ZN(n39188) );
  INV_X1 U43026 ( .A(n39171), .ZN(n39177) );
  OAI211_X1 U43027 ( .C1(n39177), .C2(n39176), .A(n39175), .B(n39174), .ZN(
        n39178) );
  INV_X1 U43028 ( .A(n39178), .ZN(n39187) );
  INV_X1 U43029 ( .A(n39179), .ZN(n39180) );
  OAI22_X1 U43030 ( .A1(n39183), .A2(n39182), .B1(n420), .B2(n39180), .ZN(
        n39185) );
  NAND2_X1 U43031 ( .A1(n39185), .A2(n39184), .ZN(n39186) );
  NAND2_X1 U43032 ( .A1(n39189), .A2(n39380), .ZN(n39190) );
  AND2_X1 U43033 ( .A1(n39191), .A2(n39190), .ZN(n39199) );
  OAI21_X1 U43034 ( .B1(n39194), .B2(n39193), .A(n39192), .ZN(n39197) );
  NOR2_X1 U43035 ( .A1(n39194), .A2(n39387), .ZN(n39196) );
  NAND2_X1 U43036 ( .A1(n41238), .A2(n52198), .ZN(n40037) );
  NOR2_X1 U43037 ( .A1(n39203), .A2(n39202), .ZN(n39218) );
  NAND2_X1 U43038 ( .A1(n39205), .A2(n39204), .ZN(n39217) );
  INV_X1 U43039 ( .A(n39210), .ZN(n39212) );
  OAI21_X1 U43040 ( .B1(n39212), .B2(n39211), .A(n39430), .ZN(n39214) );
  NAND3_X1 U43041 ( .A1(n39214), .A2(n39213), .A3(n39422), .ZN(n39215) );
  AOI21_X1 U43043 ( .B1(n39227), .B2(n39219), .A(n51508), .ZN(n39220) );
  NOR2_X1 U43044 ( .A1(n39221), .A2(n39245), .ZN(n39222) );
  MUX2_X1 U43045 ( .A(n39223), .B(n39222), .S(n39240), .Z(n39229) );
  NAND3_X1 U43046 ( .A1(n39240), .A2(n39225), .A3(n51508), .ZN(n39226) );
  NOR2_X1 U43047 ( .A1(n39227), .A2(n39226), .ZN(n39228) );
  NOR2_X1 U43048 ( .A1(n39229), .A2(n39228), .ZN(n39256) );
  INV_X1 U43049 ( .A(n39234), .ZN(n39231) );
  NAND2_X1 U43050 ( .A1(n39231), .A2(n39230), .ZN(n39255) );
  AOI21_X1 U43051 ( .B1(n39236), .B2(n51507), .A(n51063), .ZN(n39237) );
  NAND2_X1 U43052 ( .A1(n39238), .A2(n39237), .ZN(n39253) );
  INV_X1 U43053 ( .A(n39239), .ZN(n39251) );
  INV_X1 U43054 ( .A(n39240), .ZN(n39250) );
  NAND2_X1 U43055 ( .A1(n39242), .A2(n51063), .ZN(n39244) );
  NAND2_X1 U43056 ( .A1(n39244), .A2(n39243), .ZN(n39249) );
  INV_X1 U43057 ( .A(n39245), .ZN(n39246) );
  NAND2_X1 U43060 ( .A1(n39285), .A2(n39258), .ZN(n39261) );
  NAND2_X1 U43061 ( .A1(n39259), .A2(n551), .ZN(n39260) );
  MUX2_X1 U43062 ( .A(n39261), .B(n39260), .S(n39266), .Z(n39279) );
  NOR2_X1 U43063 ( .A1(n39263), .A2(n39262), .ZN(n39267) );
  AOI22_X1 U43064 ( .A1(n39267), .A2(n39266), .B1(n39265), .B2(n39264), .ZN(
        n39278) );
  NAND4_X1 U43065 ( .A1(n39275), .A2(n39274), .A3(n39273), .A4(n39281), .ZN(
        n39276) );
  NAND4_X1 U43066 ( .A1(n39279), .A2(n39278), .A3(n39277), .A4(n39276), .ZN(
        n39287) );
  INV_X1 U43067 ( .A(n39280), .ZN(n39283) );
  NAND2_X1 U43069 ( .A1(n5593), .A2(n39289), .ZN(n39292) );
  AOI21_X1 U43070 ( .B1(n39292), .B2(n39291), .A(n39290), .ZN(n39296) );
  NAND2_X1 U43071 ( .A1(n39293), .A2(n8077), .ZN(n39294) );
  INV_X1 U43072 ( .A(n39298), .ZN(n39304) );
  NAND2_X1 U43073 ( .A1(n39300), .A2(n39299), .ZN(n39303) );
  OAI22_X1 U43074 ( .A1(n39304), .A2(n39303), .B1(n39302), .B2(n39301), .ZN(
        n39305) );
  INV_X1 U43075 ( .A(n39307), .ZN(n39310) );
  INV_X1 U43076 ( .A(n39308), .ZN(n39309) );
  INV_X1 U43078 ( .A(n39316), .ZN(n41679) );
  AND2_X1 U43079 ( .A1(n6335), .A2(n41685), .ZN(n41681) );
  AND2_X1 U43080 ( .A1(n39674), .A2(n39673), .ZN(n39320) );
  NOR2_X1 U43081 ( .A1(n40684), .A2(n40676), .ZN(n39319) );
  AOI22_X1 U43082 ( .A1(n39682), .A2(n39320), .B1(n40677), .B2(n39319), .ZN(
        n39328) );
  NAND2_X1 U43083 ( .A1(n39674), .A2(n40689), .ZN(n39676) );
  NAND3_X1 U43084 ( .A1(n39676), .A2(n39321), .A3(n40684), .ZN(n39323) );
  OAI21_X1 U43085 ( .B1(n39321), .B2(n40684), .A(n40675), .ZN(n39322) );
  AND2_X1 U43086 ( .A1(n39323), .A2(n39322), .ZN(n39327) );
  NAND2_X1 U43087 ( .A1(n39682), .A2(n40677), .ZN(n40696) );
  OAI21_X1 U43088 ( .B1(n39684), .B2(n39325), .A(n39324), .ZN(n39326) );
  XNOR2_X1 U43089 ( .A(n43363), .B(n45467), .ZN(n45361) );
  NAND2_X1 U43091 ( .A1(n39329), .A2(n43665), .ZN(n39333) );
  INV_X1 U43092 ( .A(n42104), .ZN(n39330) );
  AOI21_X1 U43093 ( .B1(n41794), .B2(n39330), .A(n41804), .ZN(n39332) );
  NOR2_X1 U43094 ( .A1(n41799), .A2(n43665), .ZN(n40640) );
  INV_X1 U43095 ( .A(n40640), .ZN(n39331) );
  NAND2_X1 U43096 ( .A1(n39335), .A2(n39348), .ZN(n39339) );
  NAND3_X1 U43097 ( .A1(n39337), .A2(n39336), .A3(n39339), .ZN(n39341) );
  NAND2_X1 U43098 ( .A1(n39343), .A2(n39342), .ZN(n39344) );
  NAND3_X1 U43100 ( .A1(n39349), .A2(n39348), .A3(n39347), .ZN(n39355) );
  NOR2_X1 U43101 ( .A1(n2089), .A2(n52054), .ZN(n39352) );
  OAI21_X1 U43102 ( .B1(n39353), .B2(n39352), .A(n39351), .ZN(n39354) );
  INV_X1 U43103 ( .A(n39358), .ZN(n39364) );
  NAND2_X1 U43104 ( .A1(n39359), .A2(n39381), .ZN(n39363) );
  AND2_X1 U43105 ( .A1(n39377), .A2(n39369), .ZN(n39368) );
  INV_X1 U43106 ( .A(n39360), .ZN(n39389) );
  OAI211_X1 U43107 ( .C1(n39364), .C2(n39390), .A(n39363), .B(n39362), .ZN(
        n39365) );
  INV_X1 U43108 ( .A(n39365), .ZN(n39392) );
  NAND2_X1 U43109 ( .A1(n39366), .A2(n39368), .ZN(n39372) );
  NAND3_X1 U43110 ( .A1(n39368), .A2(n39367), .A3(n39390), .ZN(n39371) );
  OAI21_X1 U43111 ( .B1(n39386), .B2(n39377), .A(n39369), .ZN(n39370) );
  NAND3_X1 U43112 ( .A1(n39379), .A2(n39378), .A3(n39377), .ZN(n39382) );
  AOI21_X1 U43114 ( .B1(n39401), .B2(n39400), .A(n39399), .ZN(n39403) );
  INV_X1 U43116 ( .A(n39406), .ZN(n39408) );
  NOR2_X1 U43117 ( .A1(n39408), .A2(n39407), .ZN(n39409) );
  NAND2_X1 U43118 ( .A1(n42006), .A2(n41581), .ZN(n41417) );
  OR2_X1 U43119 ( .A1(n42011), .A2(n41417), .ZN(n41502) );
  OAI21_X1 U43120 ( .B1(n39429), .B2(n39410), .A(n5151), .ZN(n39413) );
  NAND3_X1 U43121 ( .A1(n39413), .A2(n39412), .A3(n39411), .ZN(n39416) );
  OAI211_X1 U43122 ( .C1(n39418), .C2(n39417), .A(n39416), .B(n39415), .ZN(
        n39419) );
  INV_X1 U43123 ( .A(n39419), .ZN(n39436) );
  INV_X1 U43125 ( .A(n39422), .ZN(n39425) );
  AOI22_X1 U43126 ( .A1(n39426), .A2(n39425), .B1(n39424), .B2(n39423), .ZN(
        n39434) );
  AOI21_X1 U43127 ( .B1(n39430), .B2(n39429), .A(n39428), .ZN(n39431) );
  NOR2_X1 U43132 ( .A1(n39445), .A2(n39027), .ZN(n39446) );
  NOR2_X1 U43133 ( .A1(n39447), .A2(n39446), .ZN(n39458) );
  OAI22_X1 U43134 ( .A1(n39453), .A2(n39452), .B1(n39451), .B2(n39450), .ZN(
        n39455) );
  NAND2_X1 U43135 ( .A1(n39455), .A2(n39454), .ZN(n39456) );
  INV_X1 U43136 ( .A(n39460), .ZN(n39468) );
  OAI22_X1 U43137 ( .A1(n39463), .A2(n39462), .B1(n39461), .B2(n39027), .ZN(
        n39465) );
  NAND2_X1 U43138 ( .A1(n39465), .A2(n51389), .ZN(n39466) );
  OAI21_X1 U43139 ( .B1(n39468), .B2(n39467), .A(n39466), .ZN(n39469) );
  AOI21_X1 U43140 ( .B1(n39473), .B2(n39472), .A(n39471), .ZN(n39477) );
  NOR2_X1 U43141 ( .A1(n39475), .A2(n39474), .ZN(n39476) );
  OAI21_X1 U43142 ( .B1(n7159), .B2(n39479), .A(n39478), .ZN(n39482) );
  AOI22_X1 U43143 ( .A1(n39483), .A2(n39482), .B1(n39481), .B2(n1075), .ZN(
        n39490) );
  NAND3_X1 U43144 ( .A1(n39488), .A2(n39487), .A3(n39486), .ZN(n39489) );
  NAND2_X1 U43145 ( .A1(n42006), .A2(n4943), .ZN(n41576) );
  NAND3_X1 U43146 ( .A1(n41502), .A2(n41580), .A3(n41576), .ZN(n39498) );
  NAND2_X1 U43147 ( .A1(n41587), .A2(n41997), .ZN(n41503) );
  NAND2_X1 U43148 ( .A1(n41503), .A2(n41417), .ZN(n39492) );
  NAND2_X1 U43149 ( .A1(n41588), .A2(n42020), .ZN(n42007) );
  INV_X1 U43150 ( .A(n42007), .ZN(n41510) );
  NAND2_X1 U43151 ( .A1(n39492), .A2(n41510), .ZN(n39497) );
  INV_X1 U43152 ( .A(n42008), .ZN(n39493) );
  AND2_X1 U43153 ( .A1(n39494), .A2(n42000), .ZN(n39496) );
  NAND2_X1 U43154 ( .A1(n41588), .A2(n41587), .ZN(n41506) );
  NAND3_X1 U43155 ( .A1(n41504), .A2(n41506), .A3(n42020), .ZN(n39495) );
  XNOR2_X1 U43156 ( .A(n44374), .B(n45354), .ZN(n43816) );
  XNOR2_X1 U43157 ( .A(n45361), .B(n43816), .ZN(n43520) );
  XNOR2_X1 U43158 ( .A(n43520), .B(n44975), .ZN(n39591) );
  NAND2_X1 U43159 ( .A1(n40668), .A2(n40663), .ZN(n39504) );
  INV_X1 U43161 ( .A(n5060), .ZN(n40185) );
  INV_X1 U43162 ( .A(n39499), .ZN(n39500) );
  NAND2_X1 U43163 ( .A1(n39501), .A2(n39500), .ZN(n39503) );
  NAND3_X1 U43164 ( .A1(n5060), .A2(n41210), .A3(n40032), .ZN(n40030) );
  NAND4_X1 U43165 ( .A1(n39504), .A2(n39503), .A3(n40022), .A4(n40030), .ZN(
        n39510) );
  NAND2_X1 U43166 ( .A1(n40669), .A2(n40029), .ZN(n39508) );
  AND2_X1 U43167 ( .A1(n51052), .A2(n40029), .ZN(n41213) );
  AOI21_X1 U43168 ( .B1(n41213), .B2(n41207), .A(n41211), .ZN(n39507) );
  NAND2_X1 U43169 ( .A1(n39505), .A2(n51430), .ZN(n39506) );
  AOI22_X1 U43170 ( .A1(n39508), .A2(n41211), .B1(n39507), .B2(n39506), .ZN(
        n39509) );
  OAI21_X1 U43171 ( .B1(n40820), .B2(n51455), .A(n39511), .ZN(n39519) );
  OAI211_X1 U43172 ( .C1(n40822), .C2(n40816), .A(n39512), .B(n39689), .ZN(
        n39518) );
  AOI21_X1 U43173 ( .B1(n40820), .B2(n40831), .A(n39513), .ZN(n39517) );
  NAND2_X1 U43174 ( .A1(n40815), .A2(n52151), .ZN(n40824) );
  NAND2_X1 U43175 ( .A1(n39515), .A2(n39514), .ZN(n39516) );
  INV_X1 U43176 ( .A(n40535), .ZN(n39521) );
  NAND2_X1 U43177 ( .A1(n40862), .A2(n40868), .ZN(n39520) );
  AOI21_X1 U43178 ( .B1(n39521), .B2(n39520), .A(n40857), .ZN(n39523) );
  INV_X1 U43179 ( .A(n39969), .ZN(n39522) );
  NOR2_X1 U43180 ( .A1(n39962), .A2(n678), .ZN(n39971) );
  OAI21_X1 U43181 ( .B1(n40864), .B2(n40863), .A(n40862), .ZN(n39524) );
  OAI21_X1 U43182 ( .B1(n39971), .B2(n40540), .A(n39524), .ZN(n39526) );
  XNOR2_X1 U43183 ( .A(n43609), .B(n4065), .ZN(n44092) );
  XNOR2_X1 U43184 ( .A(n569), .B(n44092), .ZN(n39549) );
  NOR2_X1 U43185 ( .A1(n40778), .A2(n40774), .ZN(n39796) );
  INV_X1 U43186 ( .A(n39796), .ZN(n39528) );
  NAND2_X1 U43187 ( .A1(n39528), .A2(n39527), .ZN(n39530) );
  AND2_X1 U43188 ( .A1(n40768), .A2(n40785), .ZN(n40069) );
  INV_X1 U43189 ( .A(n39800), .ZN(n40784) );
  OAI211_X1 U43190 ( .C1(n40069), .C2(n40777), .A(n432), .B(n40784), .ZN(
        n39529) );
  NAND2_X1 U43191 ( .A1(n431), .A2(n40785), .ZN(n39795) );
  INV_X1 U43192 ( .A(n39795), .ZN(n39532) );
  AND2_X1 U43193 ( .A1(n40768), .A2(n40774), .ZN(n40583) );
  NAND2_X1 U43194 ( .A1(n426), .A2(n40778), .ZN(n40598) );
  INV_X1 U43195 ( .A(n40598), .ZN(n39531) );
  OAI21_X1 U43196 ( .B1(n39532), .B2(n40583), .A(n39531), .ZN(n39536) );
  INV_X1 U43197 ( .A(n40067), .ZN(n39534) );
  AND2_X1 U43198 ( .A1(n40778), .A2(n40774), .ZN(n39799) );
  INV_X1 U43199 ( .A(n39799), .ZN(n39533) );
  NAND3_X1 U43200 ( .A1(n39534), .A2(n426), .A3(n39533), .ZN(n39535) );
  XNOR2_X1 U43201 ( .A(n39538), .B(n39537), .ZN(n39539) );
  XNOR2_X1 U43202 ( .A(n43254), .B(n39539), .ZN(n39547) );
  NAND2_X1 U43203 ( .A1(n40250), .A2(n41927), .ZN(n41926) );
  NAND3_X1 U43204 ( .A1(n39542), .A2(n39541), .A3(n40249), .ZN(n39545) );
  OAI21_X1 U43205 ( .B1(n6580), .B2(n39543), .A(n41934), .ZN(n39544) );
  XNOR2_X1 U43206 ( .A(n39547), .B(n46137), .ZN(n39548) );
  XNOR2_X1 U43207 ( .A(n39549), .B(n39548), .ZN(n39589) );
  NAND2_X1 U43208 ( .A1(n39552), .A2(n40125), .ZN(n39558) );
  INV_X1 U43209 ( .A(n39553), .ZN(n39554) );
  NAND2_X1 U43210 ( .A1(n39555), .A2(n40192), .ZN(n39557) );
  OAI211_X1 U43211 ( .C1(n40203), .C2(n40119), .A(n40196), .B(n51352), .ZN(
        n39556) );
  INV_X1 U43212 ( .A(n39560), .ZN(n39561) );
  NAND2_X1 U43213 ( .A1(n39561), .A2(n39790), .ZN(n39574) );
  INV_X1 U43214 ( .A(n39562), .ZN(n39564) );
  NAND3_X1 U43215 ( .A1(n39906), .A2(n39565), .A3(n51377), .ZN(n39563) );
  AND2_X1 U43216 ( .A1(n39564), .A2(n39563), .ZN(n39573) );
  INV_X1 U43217 ( .A(n39566), .ZN(n39567) );
  OAI211_X1 U43218 ( .C1(n38448), .C2(n39782), .A(n39919), .B(n39567), .ZN(
        n39572) );
  NAND2_X1 U43219 ( .A1(n39907), .A2(n39912), .ZN(n39900) );
  NAND2_X1 U43220 ( .A1(n39908), .A2(n37356), .ZN(n39568) );
  NAND2_X1 U43221 ( .A1(n39900), .A2(n39568), .ZN(n39570) );
  NAND2_X1 U43222 ( .A1(n39570), .A2(n39569), .ZN(n39571) );
  NOR2_X1 U43223 ( .A1(n39575), .A2(n40807), .ZN(n40794) );
  NAND2_X1 U43224 ( .A1(n43328), .A2(n39613), .ZN(n39581) );
  NAND2_X1 U43225 ( .A1(n39578), .A2(n41010), .ZN(n39580) );
  AND2_X1 U43226 ( .A1(n40807), .A2(n43323), .ZN(n41011) );
  INV_X1 U43227 ( .A(n41011), .ZN(n39579) );
  NAND2_X1 U43228 ( .A1(n39582), .A2(n40896), .ZN(n39584) );
  INV_X1 U43229 ( .A(n40271), .ZN(n39583) );
  NAND2_X1 U43230 ( .A1(n39584), .A2(n39583), .ZN(n39588) );
  AND2_X1 U43231 ( .A1(n40903), .A2(n40269), .ZN(n40911) );
  AND2_X1 U43232 ( .A1(n2224), .A2(n40081), .ZN(n40090) );
  OAI21_X1 U43233 ( .B1(n40911), .B2(n40090), .A(n40273), .ZN(n39587) );
  NAND4_X1 U43234 ( .A1(n39585), .A2(n40900), .A3(n40274), .A4(n40909), .ZN(
        n39586) );
  XNOR2_X1 U43235 ( .A(n45357), .B(n41875), .ZN(n42764) );
  XNOR2_X1 U43236 ( .A(n44364), .B(n39589), .ZN(n39590) );
  INV_X1 U43237 ( .A(n39811), .ZN(n48264) );
  NAND2_X1 U43238 ( .A1(n48268), .A2(n48264), .ZN(n44425) );
  AND2_X1 U43239 ( .A1(n48268), .A2(n48273), .ZN(n48429) );
  OAI21_X1 U43240 ( .B1(n41256), .B2(n41123), .A(n41111), .ZN(n39592) );
  OAI21_X1 U43241 ( .B1(n41113), .B2(n41265), .A(n39592), .ZN(n39597) );
  INV_X1 U43242 ( .A(n39594), .ZN(n41736) );
  NAND4_X1 U43243 ( .A1(n41736), .A2(n41256), .A3(n41269), .A4(n41268), .ZN(
        n39595) );
  OAI211_X1 U43244 ( .C1(n41734), .C2(n39597), .A(n39596), .B(n39595), .ZN(
        n41117) );
  INV_X1 U43245 ( .A(n41115), .ZN(n41733) );
  NAND2_X1 U43246 ( .A1(n41112), .A2(n41265), .ZN(n41730) );
  NAND3_X1 U43247 ( .A1(n41733), .A2(n39598), .A3(n41730), .ZN(n40473) );
  INV_X1 U43248 ( .A(n41257), .ZN(n39599) );
  NAND2_X1 U43249 ( .A1(n40473), .A2(n41737), .ZN(n39600) );
  INV_X1 U43250 ( .A(n39601), .ZN(n39602) );
  NOR2_X1 U43251 ( .A1(n6392), .A2(n40502), .ZN(n41056) );
  NAND2_X1 U43252 ( .A1(n39602), .A2(n41056), .ZN(n39608) );
  NAND3_X1 U43253 ( .A1(n41045), .A2(n40502), .A3(n41066), .ZN(n39606) );
  NAND2_X1 U43254 ( .A1(n40499), .A2(n40501), .ZN(n39605) );
  XNOR2_X1 U43255 ( .A(n42590), .B(n43928), .ZN(n43657) );
  NAND2_X1 U43256 ( .A1(n51146), .A2(n40807), .ZN(n39610) );
  INV_X1 U43257 ( .A(n41010), .ZN(n41015) );
  OAI211_X1 U43258 ( .C1(n39610), .C2(n41015), .A(n40801), .B(n39609), .ZN(
        n39612) );
  AOI21_X1 U43259 ( .B1(n41010), .B2(n43323), .A(n39611), .ZN(n41007) );
  INV_X1 U43260 ( .A(n39614), .ZN(n39615) );
  INV_X1 U43261 ( .A(n39616), .ZN(n39617) );
  NAND2_X1 U43262 ( .A1(n39617), .A2(n41004), .ZN(n39618) );
  NOR2_X1 U43263 ( .A1(n41645), .A2(n41642), .ZN(n41640) );
  INV_X1 U43264 ( .A(n41640), .ZN(n41979) );
  NAND2_X1 U43265 ( .A1(n41103), .A2(n41646), .ZN(n40609) );
  NAND4_X1 U43266 ( .A1(n41979), .A2(n41986), .A3(n41977), .A4(n41650), .ZN(
        n39625) );
  AND2_X1 U43267 ( .A1(n41645), .A2(n41650), .ZN(n41984) );
  INV_X1 U43268 ( .A(n41984), .ZN(n39620) );
  AND2_X1 U43270 ( .A1(n6938), .A2(n41975), .ZN(n41093) );
  NAND2_X1 U43271 ( .A1(n41977), .A2(n41093), .ZN(n41099) );
  NAND2_X1 U43272 ( .A1(n41981), .A2(n41642), .ZN(n39621) );
  NAND4_X1 U43273 ( .A1(n41974), .A2(n39622), .A3(n41099), .A4(n39621), .ZN(
        n39624) );
  NOR2_X1 U43274 ( .A1(n41645), .A2(n6940), .ZN(n41095) );
  OR2_X1 U43275 ( .A1(n41642), .A2(n41646), .ZN(n40606) );
  NAND3_X1 U43276 ( .A1(n41095), .A2(n41647), .A3(n40606), .ZN(n39623) );
  XNOR2_X1 U43277 ( .A(n43657), .B(n43751), .ZN(n39661) );
  NOR2_X1 U43278 ( .A1(n41328), .A2(n41332), .ZN(n40371) );
  OAI22_X1 U43282 ( .A1(n40751), .A2(n39633), .B1(n41343), .B2(n39632), .ZN(
        n39883) );
  INV_X1 U43283 ( .A(n39883), .ZN(n39639) );
  OAI211_X1 U43284 ( .C1(n41353), .C2(n41356), .A(n41358), .B(n41339), .ZN(
        n39634) );
  NAND2_X1 U43285 ( .A1(n39634), .A2(n39884), .ZN(n39638) );
  INV_X1 U43286 ( .A(n41355), .ZN(n41349) );
  NAND4_X1 U43288 ( .A1(n41358), .A2(n41349), .A3(n41354), .A4(n41360), .ZN(
        n39636) );
  NAND4_X2 U43289 ( .A1(n39639), .A2(n39638), .A3(n39637), .A4(n39636), .ZN(
        n43655) );
  NAND3_X1 U43290 ( .A1(n39640), .A2(n39646), .A3(n40343), .ZN(n39641) );
  AND2_X1 U43291 ( .A1(n39642), .A2(n39641), .ZN(n39652) );
  INV_X1 U43292 ( .A(n39643), .ZN(n39645) );
  INV_X1 U43293 ( .A(n39644), .ZN(n40333) );
  NOR2_X1 U43294 ( .A1(n40327), .A2(n40338), .ZN(n39858) );
  NAND3_X1 U43295 ( .A1(n39645), .A2(n40333), .A3(n39858), .ZN(n39651) );
  OAI211_X1 U43296 ( .C1(n40335), .C2(n39857), .A(n40337), .B(n52101), .ZN(
        n39650) );
  NAND2_X1 U43297 ( .A1(n39647), .A2(n39646), .ZN(n39648) );
  NAND2_X1 U43298 ( .A1(n39648), .A2(n40337), .ZN(n39649) );
  NAND4_X2 U43299 ( .A1(n39652), .A2(n39651), .A3(n39650), .A4(n39649), .ZN(
        n45314) );
  NAND2_X1 U43300 ( .A1(n39654), .A2(n39653), .ZN(n39655) );
  INV_X1 U43301 ( .A(n40549), .ZN(n40318) );
  INV_X1 U43302 ( .A(n40573), .ZN(n40319) );
  NAND2_X1 U43303 ( .A1(n40559), .A2(n7848), .ZN(n39657) );
  XNOR2_X1 U43304 ( .A(n45314), .B(n43155), .ZN(n44347) );
  XNOR2_X1 U43305 ( .A(n43755), .B(n44347), .ZN(n39660) );
  NAND4_X1 U43306 ( .A1(n39663), .A2(n40013), .A3(n51297), .A4(n39662), .ZN(
        n39671) );
  NAND2_X1 U43307 ( .A1(n39664), .A2(n39997), .ZN(n39665) );
  OAI21_X1 U43308 ( .B1(n40685), .B2(n40684), .A(n39672), .ZN(n39679) );
  NOR2_X1 U43309 ( .A1(n39929), .A2(n39673), .ZN(n39678) );
  NAND2_X1 U43310 ( .A1(n39674), .A2(n51022), .ZN(n39675) );
  NAND2_X1 U43311 ( .A1(n39676), .A2(n39675), .ZN(n39677) );
  AOI22_X1 U43312 ( .A1(n39679), .A2(n39678), .B1(n39677), .B2(n40672), .ZN(
        n39688) );
  INV_X1 U43313 ( .A(n40693), .ZN(n39681) );
  AOI21_X1 U43314 ( .B1(n39682), .B2(n39681), .A(n39680), .ZN(n39926) );
  INV_X1 U43315 ( .A(n39926), .ZN(n39687) );
  NAND2_X1 U43316 ( .A1(n40674), .A2(n40690), .ZN(n39686) );
  OAI211_X1 U43317 ( .C1(n39684), .C2(n40672), .A(n40684), .B(n39683), .ZN(
        n39685) );
  NOR2_X1 U43318 ( .A1(n39690), .A2(n40836), .ZN(n39694) );
  AOI22_X1 U43319 ( .A1(n39694), .A2(n39693), .B1(n39692), .B2(n39691), .ZN(
        n39698) );
  XNOR2_X1 U43320 ( .A(n43014), .B(n45097), .ZN(n39699) );
  XNOR2_X1 U43321 ( .A(n39699), .B(n52171), .ZN(n45450) );
  NOR2_X1 U43322 ( .A1(n39702), .A2(n39701), .ZN(n39703) );
  INV_X1 U43323 ( .A(n41076), .ZN(n39717) );
  NAND2_X1 U43324 ( .A1(n39709), .A2(n39708), .ZN(n39710) );
  NAND2_X1 U43325 ( .A1(n39713), .A2(n39712), .ZN(n41074) );
  INV_X1 U43326 ( .A(n41074), .ZN(n39714) );
  XNOR2_X1 U43327 ( .A(n39719), .B(n39718), .ZN(n39722) );
  XNOR2_X1 U43328 ( .A(n39720), .B(n43537), .ZN(n39721) );
  XNOR2_X1 U43329 ( .A(n39722), .B(n39721), .ZN(n39723) );
  XNOR2_X1 U43330 ( .A(n44944), .B(n39723), .ZN(n39724) );
  XNOR2_X1 U43331 ( .A(n45450), .B(n39724), .ZN(n39725) );
  AND2_X1 U43332 ( .A1(n41276), .A2(n41275), .ZN(n41024) );
  NAND2_X1 U43333 ( .A1(n41024), .A2(n41039), .ZN(n41031) );
  INV_X1 U43334 ( .A(n39726), .ZN(n40430) );
  INV_X1 U43335 ( .A(n39727), .ZN(n39728) );
  NOR2_X1 U43336 ( .A1(n52192), .A2(n41292), .ZN(n41278) );
  INV_X1 U43337 ( .A(n41293), .ZN(n41034) );
  AOI21_X1 U43338 ( .B1(n40417), .B2(n5324), .A(n397), .ZN(n39733) );
  NAND2_X1 U43339 ( .A1(n40417), .A2(n41276), .ZN(n39731) );
  NAND2_X1 U43340 ( .A1(n39731), .A2(n40420), .ZN(n39732) );
  OR2_X1 U43341 ( .A1(n39738), .A2(n39737), .ZN(n40439) );
  NAND2_X1 U43342 ( .A1(n40396), .A2(n40404), .ZN(n39739) );
  AND2_X1 U43343 ( .A1(n39739), .A2(n40439), .ZN(n39743) );
  NAND2_X1 U43344 ( .A1(n39740), .A2(n40456), .ZN(n39742) );
  NAND2_X1 U43345 ( .A1(n39962), .A2(n40874), .ZN(n39744) );
  NOR2_X1 U43346 ( .A1(n40533), .A2(n39746), .ZN(n40861) );
  INV_X1 U43347 ( .A(n40857), .ZN(n40543) );
  NAND3_X1 U43348 ( .A1(n40859), .A2(n39747), .A3(n40868), .ZN(n39748) );
  NAND3_X1 U43349 ( .A1(n39937), .A2(n39942), .A3(n52094), .ZN(n39758) );
  NAND2_X1 U43350 ( .A1(n39955), .A2(n39751), .ZN(n39939) );
  INV_X1 U43351 ( .A(n39939), .ZN(n39753) );
  OAI21_X1 U43352 ( .B1(n39753), .B2(n39760), .A(n39957), .ZN(n39757) );
  NAND2_X1 U43353 ( .A1(n39755), .A2(n39754), .ZN(n39756) );
  OAI211_X1 U43354 ( .C1(n39759), .C2(n39758), .A(n39757), .B(n39756), .ZN(
        n39765) );
  NAND3_X1 U43355 ( .A1(n39762), .A2(n39938), .A3(n39761), .ZN(n39763) );
  XNOR2_X1 U43356 ( .A(n2206), .B(n42819), .ZN(n41159) );
  NOR2_X1 U43357 ( .A1(n39767), .A2(n40655), .ZN(n39769) );
  OAI21_X1 U43358 ( .B1(n40643), .B2(n39769), .A(n39768), .ZN(n39770) );
  MUX2_X1 U43359 ( .A(n39771), .B(n39770), .S(n40651), .Z(n39780) );
  AOI21_X1 U43360 ( .B1(n40652), .B2(n5982), .A(n39772), .ZN(n39778) );
  NAND2_X1 U43361 ( .A1(n41451), .A2(n39775), .ZN(n39777) );
  AOI21_X1 U43362 ( .B1(n39778), .B2(n39777), .A(n39776), .ZN(n39779) );
  INV_X1 U43363 ( .A(n39781), .ZN(n39784) );
  NOR2_X1 U43364 ( .A1(n39782), .A2(n39906), .ZN(n39783) );
  AOI21_X1 U43365 ( .B1(n39784), .B2(n39915), .A(n39783), .ZN(n39794) );
  OAI21_X1 U43366 ( .B1(n39919), .B2(n6645), .A(n39785), .ZN(n39786) );
  NAND2_X1 U43367 ( .A1(n39786), .A2(n39904), .ZN(n39793) );
  NAND2_X1 U43368 ( .A1(n39788), .A2(n39787), .ZN(n39792) );
  NOR2_X1 U43369 ( .A1(n39790), .A2(n39789), .ZN(n39905) );
  INV_X1 U43370 ( .A(n39905), .ZN(n39791) );
  XNOR2_X1 U43371 ( .A(n44559), .B(n46050), .ZN(n39808) );
  NAND2_X1 U43372 ( .A1(n40598), .A2(n681), .ZN(n39797) );
  NAND2_X1 U43374 ( .A1(n39800), .A2(n39799), .ZN(n40589) );
  NAND3_X1 U43375 ( .A1(n39802), .A2(n40783), .A3(n39801), .ZN(n39805) );
  INV_X1 U43376 ( .A(n40786), .ZN(n39803) );
  NAND3_X1 U43377 ( .A1(n40596), .A2(n39803), .A3(n40585), .ZN(n39804) );
  XNOR2_X1 U43378 ( .A(n43206), .B(n2117), .ZN(n39807) );
  XNOR2_X1 U43379 ( .A(n39808), .B(n39807), .ZN(n43012) );
  XNOR2_X1 U43380 ( .A(n41159), .B(n43012), .ZN(n39809) );
  XNOR2_X1 U43381 ( .A(n39810), .B(n39809), .ZN(n39813) );
  NAND3_X1 U43382 ( .A1(n48429), .A2(n44431), .A3(n48433), .ZN(n48426) );
  OAI21_X1 U43383 ( .B1(n44427), .B2(n44425), .A(n48426), .ZN(n45594) );
  INV_X1 U43384 ( .A(n39812), .ZN(n45589) );
  NAND2_X1 U43385 ( .A1(n48423), .A2(n45590), .ZN(n45588) );
  NOR2_X1 U43386 ( .A1(n39814), .A2(n40373), .ZN(n41895) );
  NOR2_X1 U43387 ( .A1(n2379), .A2(n41329), .ZN(n39815) );
  NOR2_X1 U43388 ( .A1(n41895), .A2(n39815), .ZN(n39829) );
  NAND3_X1 U43391 ( .A1(n39817), .A2(n41316), .A3(n39816), .ZN(n39819) );
  NAND2_X1 U43392 ( .A1(n39819), .A2(n39818), .ZN(n39826) );
  NAND2_X1 U43393 ( .A1(n39826), .A2(n39820), .ZN(n39824) );
  NAND2_X1 U43394 ( .A1(n674), .A2(n39821), .ZN(n39823) );
  NAND2_X1 U43395 ( .A1(n41902), .A2(n52215), .ZN(n40372) );
  NAND2_X1 U43396 ( .A1(n40371), .A2(n41331), .ZN(n40727) );
  INV_X1 U43397 ( .A(n40727), .ZN(n41894) );
  NAND3_X1 U43398 ( .A1(n41328), .A2(n52214), .A3(n41332), .ZN(n41898) );
  NOR2_X1 U43399 ( .A1(n41898), .A2(n41902), .ZN(n39825) );
  NOR2_X1 U43400 ( .A1(n41894), .A2(n39825), .ZN(n39828) );
  INV_X1 U43401 ( .A(n39826), .ZN(n41901) );
  NAND3_X1 U43402 ( .A1(n41901), .A2(n41329), .A3(n41900), .ZN(n39827) );
  NOR2_X1 U43404 ( .A1(n39843), .A2(n39830), .ZN(n39833) );
  OAI22_X1 U43405 ( .A1(n39842), .A2(n39839), .B1(n39831), .B2(n1931), .ZN(
        n39832) );
  NOR2_X1 U43406 ( .A1(n39833), .A2(n39832), .ZN(n39848) );
  OR2_X1 U43407 ( .A1(n40380), .A2(n40381), .ZN(n40378) );
  NAND3_X1 U43408 ( .A1(n40378), .A2(n40388), .A3(n40377), .ZN(n39847) );
  NAND2_X1 U43409 ( .A1(n1931), .A2(n39834), .ZN(n39838) );
  INV_X1 U43410 ( .A(n39835), .ZN(n39837) );
  NAND4_X1 U43411 ( .A1(n39838), .A2(n39837), .A3(n40385), .A4(n52083), .ZN(
        n39841) );
  NAND3_X1 U43412 ( .A1(n38611), .A2(n40382), .A3(n40377), .ZN(n39840) );
  AND2_X1 U43413 ( .A1(n39841), .A2(n39840), .ZN(n39846) );
  NAND3_X1 U43414 ( .A1(n40384), .A2(n39843), .A3(n39842), .ZN(n39844) );
  NAND2_X1 U43415 ( .A1(n39844), .A2(n40377), .ZN(n39845) );
  OAI21_X1 U43416 ( .B1(n39850), .B2(n40328), .A(n40343), .ZN(n39852) );
  NAND3_X1 U43417 ( .A1(n40333), .A2(n7117), .A3(n40327), .ZN(n39851) );
  AOI21_X1 U43418 ( .B1(n39852), .B2(n39851), .A(n52101), .ZN(n39869) );
  NAND3_X1 U43419 ( .A1(n40333), .A2(n40335), .A3(n52101), .ZN(n39861) );
  NAND2_X1 U43420 ( .A1(n39856), .A2(n39855), .ZN(n39860) );
  NAND3_X1 U43421 ( .A1(n39858), .A2(n7117), .A3(n39857), .ZN(n39859) );
  INV_X1 U43422 ( .A(n39862), .ZN(n39866) );
  NAND2_X1 U43423 ( .A1(n40328), .A2(n40330), .ZN(n39863) );
  INV_X1 U43424 ( .A(n40335), .ZN(n39864) );
  MUX2_X1 U43425 ( .A(n39866), .B(n39865), .S(n39864), .Z(n39867) );
  AOI22_X1 U43427 ( .A1(n39871), .A2(n41164), .B1(n41163), .B2(n39870), .ZN(
        n39881) );
  OAI211_X1 U43428 ( .C1(n41168), .C2(n41174), .A(n40353), .B(n39872), .ZN(
        n39880) );
  OAI21_X1 U43429 ( .B1(n2179), .B2(n41690), .A(n41609), .ZN(n39876) );
  NOR2_X1 U43430 ( .A1(n39874), .A2(n41703), .ZN(n39875) );
  AOI22_X1 U43431 ( .A1(n41702), .A2(n39876), .B1(n39875), .B2(n41707), .ZN(
        n39879) );
  INV_X1 U43432 ( .A(n41168), .ZN(n40355) );
  AND2_X1 U43433 ( .A1(n41706), .A2(n41691), .ZN(n41708) );
  OAI21_X1 U43434 ( .B1(n40355), .B2(n39877), .A(n41708), .ZN(n39878) );
  XNOR2_X1 U43436 ( .A(n44076), .B(n44960), .ZN(n43272) );
  NAND2_X1 U43437 ( .A1(n39883), .A2(n39882), .ZN(n39898) );
  AND2_X1 U43438 ( .A1(n41354), .A2(n41348), .ZN(n39886) );
  NOR2_X1 U43439 ( .A1(n41348), .A2(n41360), .ZN(n39885) );
  OAI21_X1 U43440 ( .B1(n39886), .B2(n39885), .A(n41355), .ZN(n39887) );
  NOR2_X1 U43441 ( .A1(n40744), .A2(n39888), .ZN(n39897) );
  INV_X1 U43442 ( .A(n39889), .ZN(n39890) );
  NAND3_X1 U43443 ( .A1(n39890), .A2(n6469), .A3(n41348), .ZN(n39894) );
  NAND3_X1 U43444 ( .A1(n41344), .A2(n39891), .A3(n41356), .ZN(n39893) );
  NAND2_X1 U43445 ( .A1(n39895), .A2(n41356), .ZN(n39896) );
  NOR2_X1 U43446 ( .A1(n39899), .A2(n51377), .ZN(n39901) );
  AOI21_X1 U43447 ( .B1(n39902), .B2(n39901), .A(n39900), .ZN(n39903) );
  OAI21_X1 U43448 ( .B1(n39905), .B2(n39904), .A(n39903), .ZN(n39924) );
  NOR2_X1 U43449 ( .A1(n39906), .A2(n39912), .ZN(n39911) );
  MUX2_X1 U43450 ( .A(n38448), .B(n39907), .S(n51377), .Z(n39909) );
  AOI22_X1 U43451 ( .A1(n39911), .A2(n39910), .B1(n39909), .B2(n39908), .ZN(
        n39923) );
  AND2_X1 U43452 ( .A1(n39912), .A2(n51377), .ZN(n39917) );
  NOR2_X1 U43453 ( .A1(n38448), .A2(n37356), .ZN(n39913) );
  AOI22_X1 U43454 ( .A1(n39915), .A2(n39914), .B1(n39917), .B2(n39913), .ZN(
        n39922) );
  NOR2_X1 U43455 ( .A1(n39916), .A2(n38448), .ZN(n39920) );
  AOI22_X1 U43456 ( .A1(n39920), .A2(n39919), .B1(n39918), .B2(n39917), .ZN(
        n39921) );
  NAND4_X1 U43457 ( .A1(n39924), .A2(n39923), .A3(n39922), .A4(n39921), .ZN(
        n44160) );
  OAI211_X1 U43458 ( .C1(n40685), .C2(n39929), .A(n40672), .B(n40689), .ZN(
        n39925) );
  NAND2_X1 U43459 ( .A1(n39926), .A2(n39925), .ZN(n39936) );
  NOR2_X1 U43460 ( .A1(n39927), .A2(n39929), .ZN(n40673) );
  NAND2_X1 U43461 ( .A1(n40673), .A2(n40683), .ZN(n39928) );
  AND2_X1 U43462 ( .A1(n39928), .A2(n40696), .ZN(n39935) );
  AND2_X1 U43463 ( .A1(n51022), .A2(n40676), .ZN(n40691) );
  AOI22_X1 U43465 ( .A1(n40691), .A2(n39930), .B1(n40693), .B2(n39929), .ZN(
        n39934) );
  OAI22_X1 U43466 ( .A1(n39931), .A2(n40676), .B1(n40692), .B2(n40689), .ZN(
        n39932) );
  NAND2_X1 U43467 ( .A1(n39932), .A2(n40677), .ZN(n39933) );
  OAI21_X1 U43468 ( .B1(n39940), .B2(n39955), .A(n39939), .ZN(n39941) );
  NAND2_X1 U43469 ( .A1(n39942), .A2(n575), .ZN(n39947) );
  NAND3_X1 U43470 ( .A1(n52073), .A2(n575), .A3(n39943), .ZN(n39946) );
  OAI21_X1 U43471 ( .B1(n39954), .B2(n39947), .A(n39946), .ZN(n39948) );
  INV_X1 U43472 ( .A(n39948), .ZN(n39960) );
  OAI21_X1 U43473 ( .B1(n684), .B2(n39950), .A(n39949), .ZN(n39952) );
  NAND2_X1 U43474 ( .A1(n39952), .A2(n39951), .ZN(n39959) );
  NAND2_X1 U43475 ( .A1(n39954), .A2(n39953), .ZN(n39956) );
  NAND2_X1 U43476 ( .A1(n39956), .A2(n39955), .ZN(n39958) );
  OAI211_X1 U43477 ( .C1(n40862), .C2(n40526), .A(n39962), .B(n40868), .ZN(
        n39963) );
  INV_X1 U43478 ( .A(n39963), .ZN(n39964) );
  NAND2_X1 U43479 ( .A1(n40876), .A2(n40874), .ZN(n39967) );
  MUX2_X1 U43480 ( .A(n39967), .B(n39966), .S(n40868), .Z(n39974) );
  AND2_X1 U43481 ( .A1(n6525), .A2(n40868), .ZN(n40541) );
  OAI21_X1 U43482 ( .B1(n40541), .B2(n40869), .A(n39968), .ZN(n39970) );
  AND2_X1 U43483 ( .A1(n39969), .A2(n39970), .ZN(n39973) );
  AOI22_X1 U43484 ( .A1(n39971), .A2(n40540), .B1(n40860), .B2(n40862), .ZN(
        n39972) );
  NAND4_X2 U43485 ( .A1(n39975), .A2(n39973), .A3(n39974), .A4(n39972), .ZN(
        n45484) );
  XNOR2_X1 U43486 ( .A(n45484), .B(n39976), .ZN(n39977) );
  XNOR2_X1 U43487 ( .A(n40979), .B(n39977), .ZN(n40021) );
  INV_X1 U43488 ( .A(n39978), .ZN(n40459) );
  INV_X1 U43489 ( .A(n39979), .ZN(n39980) );
  NAND2_X1 U43490 ( .A1(n39980), .A2(n40447), .ZN(n39981) );
  NAND3_X1 U43491 ( .A1(n40458), .A2(n40453), .A3(n40450), .ZN(n40454) );
  NOR2_X1 U43492 ( .A1(n40453), .A2(n40446), .ZN(n39985) );
  NAND2_X1 U43493 ( .A1(n39985), .A2(n40458), .ZN(n39982) );
  NAND2_X1 U43494 ( .A1(n40454), .A2(n39982), .ZN(n39983) );
  NOR2_X1 U43495 ( .A1(n40401), .A2(n39983), .ZN(n39993) );
  NAND3_X1 U43496 ( .A1(n40458), .A2(n40456), .A3(n40450), .ZN(n39984) );
  MUX2_X1 U43497 ( .A(n40395), .B(n39984), .S(n6851), .Z(n39992) );
  NAND2_X1 U43498 ( .A1(n2854), .A2(n40456), .ZN(n39989) );
  INV_X1 U43499 ( .A(n40458), .ZN(n39987) );
  INV_X1 U43500 ( .A(n39985), .ZN(n39986) );
  NAND3_X1 U43501 ( .A1(n39987), .A2(n39986), .A3(n40436), .ZN(n39988) );
  OAI211_X1 U43502 ( .C1(n39990), .C2(n39989), .A(n40404), .B(n39988), .ZN(
        n39991) );
  NAND2_X1 U43503 ( .A1(n40014), .A2(n51297), .ZN(n39996) );
  AND2_X1 U43504 ( .A1(n6861), .A2(n39996), .ZN(n39999) );
  MUX2_X1 U43505 ( .A(n39999), .B(n39998), .S(n39997), .Z(n40020) );
  OAI21_X1 U43506 ( .B1(n40015), .B2(n40001), .A(n40000), .ZN(n40007) );
  INV_X1 U43507 ( .A(n40002), .ZN(n40004) );
  AOI21_X1 U43508 ( .B1(n40005), .B2(n40004), .A(n40003), .ZN(n40006) );
  INV_X1 U43509 ( .A(n40008), .ZN(n40012) );
  INV_X1 U43510 ( .A(n40009), .ZN(n40010) );
  AOI22_X1 U43511 ( .A1(n40013), .A2(n40012), .B1(n40011), .B2(n40010), .ZN(
        n40019) );
  NAND3_X1 U43512 ( .A1(n40016), .A2(n40015), .A3(n40014), .ZN(n40017) );
  XNOR2_X1 U43513 ( .A(n45344), .B(n44398), .ZN(n40165) );
  OAI22_X1 U43514 ( .A1(n41212), .A2(n40023), .B1(n41200), .B2(n40028), .ZN(
        n40025) );
  NAND2_X1 U43515 ( .A1(n51430), .A2(n41202), .ZN(n40024) );
  MUX2_X1 U43516 ( .A(n40025), .B(n40024), .S(n685), .Z(n40027) );
  NAND2_X1 U43517 ( .A1(n40669), .A2(n5060), .ZN(n40026) );
  NAND2_X1 U43518 ( .A1(n40027), .A2(n40026), .ZN(n40036) );
  INV_X1 U43519 ( .A(n40028), .ZN(n40034) );
  OAI211_X1 U43520 ( .C1(n41207), .C2(n40034), .A(n40031), .B(n40030), .ZN(
        n40035) );
  INV_X1 U43521 ( .A(n41212), .ZN(n41193) );
  AOI21_X1 U43522 ( .B1(n40037), .B2(n40210), .A(n41245), .ZN(n40039) );
  INV_X1 U43524 ( .A(n40040), .ZN(n40038) );
  NAND2_X1 U43526 ( .A1(n40717), .A2(n41227), .ZN(n40041) );
  XNOR2_X1 U43527 ( .A(n44963), .B(n1341), .ZN(n40042) );
  XNOR2_X1 U43528 ( .A(n43079), .B(n40042), .ZN(n40080) );
  NOR3_X1 U43529 ( .A1(n40295), .A2(n41480), .A3(n42062), .ZN(n42443) );
  INV_X1 U43530 ( .A(n42443), .ZN(n42440) );
  NAND2_X1 U43531 ( .A1(n42062), .A2(n596), .ZN(n40045) );
  NAND2_X1 U43532 ( .A1(n42440), .A2(n40045), .ZN(n40044) );
  AND2_X1 U43533 ( .A1(n40049), .A2(n42062), .ZN(n40043) );
  AOI21_X1 U43534 ( .B1(n40044), .B2(n42441), .A(n40043), .ZN(n40057) );
  NAND3_X1 U43535 ( .A1(n42441), .A2(n42061), .A3(n480), .ZN(n40048) );
  INV_X1 U43536 ( .A(n40045), .ZN(n40046) );
  NAND2_X1 U43537 ( .A1(n40046), .A2(n679), .ZN(n40047) );
  MUX2_X1 U43538 ( .A(n40048), .B(n40047), .S(n40295), .Z(n40056) );
  OAI211_X1 U43539 ( .C1(n52128), .C2(n42052), .A(n40050), .B(n40293), .ZN(
        n40055) );
  INV_X1 U43540 ( .A(n40051), .ZN(n41485) );
  NAND2_X1 U43541 ( .A1(n41482), .A2(n480), .ZN(n40052) );
  OAI21_X1 U43542 ( .B1(n41485), .B2(n40052), .A(n40288), .ZN(n40053) );
  INV_X1 U43543 ( .A(n42053), .ZN(n40296) );
  NAND2_X1 U43544 ( .A1(n40053), .A2(n40296), .ZN(n40054) );
  NAND4_X2 U43545 ( .A1(n40057), .A2(n40056), .A3(n40055), .A4(n40054), .ZN(
        n44074) );
  INV_X1 U43546 ( .A(n40583), .ZN(n40058) );
  NOR2_X1 U43547 ( .A1(n40059), .A2(n40058), .ZN(n40068) );
  INV_X1 U43548 ( .A(n40774), .ZN(n40592) );
  NOR2_X1 U43549 ( .A1(n40592), .A2(n40768), .ZN(n40586) );
  NAND3_X1 U43550 ( .A1(n40062), .A2(n40061), .A3(n40060), .ZN(n40065) );
  INV_X1 U43551 ( .A(n40063), .ZN(n40064) );
  OAI21_X1 U43552 ( .B1(n40065), .B2(n40064), .A(n40785), .ZN(n40769) );
  INV_X1 U43553 ( .A(n40769), .ZN(n40066) );
  NAND2_X1 U43555 ( .A1(n40774), .A2(n40785), .ZN(n40072) );
  AOI22_X1 U43556 ( .A1(n40069), .A2(n432), .B1(n40072), .B2(n40778), .ZN(
        n40071) );
  NOR2_X1 U43557 ( .A1(n40768), .A2(n40785), .ZN(n40782) );
  AOI21_X1 U43558 ( .B1(n40782), .B2(n432), .A(n40777), .ZN(n40070) );
  OAI211_X1 U43559 ( .C1(n40768), .C2(n40072), .A(n40071), .B(n40070), .ZN(
        n40078) );
  MUX2_X1 U43560 ( .A(n40774), .B(n40777), .S(n40778), .Z(n40074) );
  AOI22_X1 U43561 ( .A1(n40074), .A2(n432), .B1(n40600), .B2(n40073), .ZN(
        n40077) );
  INV_X1 U43562 ( .A(n40589), .ZN(n40075) );
  NAND2_X1 U43563 ( .A1(n40075), .A2(n40591), .ZN(n40076) );
  XNOR2_X1 U43565 ( .A(n44074), .B(n51460), .ZN(n43884) );
  XNOR2_X1 U43566 ( .A(n40080), .B(n43884), .ZN(n42887) );
  NAND2_X1 U43567 ( .A1(n2616), .A2(n40081), .ZN(n40084) );
  INV_X1 U43568 ( .A(n40911), .ZN(n40082) );
  MUX2_X1 U43569 ( .A(n40084), .B(n40083), .S(n40082), .Z(n40103) );
  NAND2_X1 U43570 ( .A1(n40910), .A2(n40909), .ZN(n40905) );
  INV_X1 U43571 ( .A(n40905), .ZN(n40088) );
  NAND2_X1 U43572 ( .A1(n40900), .A2(n2223), .ZN(n40085) );
  NAND3_X1 U43574 ( .A1(n40089), .A2(n40906), .A3(n40088), .ZN(n40092) );
  NAND3_X1 U43575 ( .A1(n40090), .A2(n40900), .A3(n40903), .ZN(n40091) );
  AND2_X1 U43576 ( .A1(n40094), .A2(n2223), .ZN(n40095) );
  AOI22_X1 U43577 ( .A1(n40096), .A2(n40271), .B1(n5073), .B2(n40095), .ZN(
        n40101) );
  OAI21_X1 U43578 ( .B1(n40097), .B2(n40900), .A(n40271), .ZN(n40099) );
  INV_X1 U43579 ( .A(n40098), .ZN(n40895) );
  NAND2_X1 U43580 ( .A1(n40099), .A2(n40895), .ZN(n40100) );
  INV_X1 U43581 ( .A(n40104), .ZN(n40105) );
  XNOR2_X1 U43582 ( .A(n43074), .B(n40105), .ZN(n40106) );
  XNOR2_X1 U43583 ( .A(n40107), .B(n40106), .ZN(n40108) );
  XNOR2_X1 U43584 ( .A(n42316), .B(n40108), .ZN(n40132) );
  NAND3_X1 U43585 ( .A1(n40111), .A2(n40110), .A3(n584), .ZN(n40112) );
  AOI21_X1 U43586 ( .B1(n40112), .B2(n40125), .A(n40120), .ZN(n40131) );
  NAND2_X1 U43587 ( .A1(n40113), .A2(n40196), .ZN(n40116) );
  INV_X1 U43588 ( .A(n40114), .ZN(n40115) );
  NAND4_X1 U43589 ( .A1(n40116), .A2(n40115), .A3(n51325), .A4(n40195), .ZN(
        n40130) );
  NAND3_X1 U43590 ( .A1(n40119), .A2(n40118), .A3(n51352), .ZN(n40123) );
  MUX2_X1 U43591 ( .A(n40126), .B(n51233), .S(n507), .Z(n40128) );
  NAND2_X1 U43592 ( .A1(n40128), .A2(n40127), .ZN(n40129) );
  XNOR2_X1 U43593 ( .A(n40132), .B(n42500), .ZN(n40162) );
  OAI21_X1 U43594 ( .B1(n40133), .B2(n51455), .A(n40840), .ZN(n40145) );
  OAI21_X1 U43595 ( .B1(n40836), .B2(n40818), .A(n40839), .ZN(n40134) );
  NAND2_X1 U43596 ( .A1(n40134), .A2(n40831), .ZN(n40144) );
  NOR2_X1 U43597 ( .A1(n51455), .A2(n40828), .ZN(n40137) );
  NAND2_X1 U43598 ( .A1(n51990), .A2(n40823), .ZN(n40136) );
  NAND2_X1 U43599 ( .A1(n40823), .A2(n40828), .ZN(n40140) );
  OAI21_X1 U43600 ( .B1(n40822), .B2(n40818), .A(n40140), .ZN(n40142) );
  INV_X1 U43602 ( .A(n40148), .ZN(n40149) );
  NAND2_X1 U43605 ( .A1(n40556), .A2(n40565), .ZN(n40563) );
  NAND2_X1 U43606 ( .A1(n40556), .A2(n40558), .ZN(n40153) );
  INV_X1 U43607 ( .A(n40154), .ZN(n40576) );
  NOR2_X1 U43609 ( .A1(n40157), .A2(n40156), .ZN(n40158) );
  OAI21_X1 U43610 ( .B1(n40158), .B2(n40573), .A(n2597), .ZN(n40159) );
  XNOR2_X1 U43611 ( .A(n43106), .B(n45339), .ZN(n43069) );
  XNOR2_X1 U43612 ( .A(n40162), .B(n43069), .ZN(n40163) );
  XNOR2_X1 U43613 ( .A(n42887), .B(n40163), .ZN(n40164) );
  XNOR2_X1 U43614 ( .A(n40165), .B(n40164), .ZN(n40174) );
  AND2_X1 U43615 ( .A1(n48436), .A2(n48264), .ZN(n40168) );
  NAND2_X1 U43616 ( .A1(n45588), .A2(n40168), .ZN(n40180) );
  NAND2_X1 U43617 ( .A1(n48268), .A2(n660), .ZN(n40166) );
  OAI21_X1 U43618 ( .B1(n45590), .B2(n48259), .A(n40166), .ZN(n40167) );
  NAND3_X1 U43619 ( .A1(n40167), .A2(n48433), .A3(n48436), .ZN(n40171) );
  NAND2_X1 U43620 ( .A1(n48429), .A2(n40168), .ZN(n40170) );
  NAND2_X1 U43621 ( .A1(n48423), .A2(n44427), .ZN(n40169) );
  AND3_X1 U43622 ( .A1(n40171), .A2(n40170), .A3(n40169), .ZN(n40179) );
  INV_X1 U43623 ( .A(n45590), .ZN(n48260) );
  NAND2_X1 U43624 ( .A1(n48260), .A2(n48438), .ZN(n40173) );
  NAND2_X1 U43625 ( .A1(n48423), .A2(n48434), .ZN(n40172) );
  NAND2_X1 U43626 ( .A1(n40173), .A2(n40172), .ZN(n40178) );
  INV_X1 U43628 ( .A(n44427), .ZN(n48424) );
  NAND2_X1 U43629 ( .A1(n48424), .A2(n48438), .ZN(n40176) );
  INV_X1 U43630 ( .A(n40174), .ZN(n48269) );
  NAND2_X1 U43631 ( .A1(n40176), .A2(n40175), .ZN(n40177) );
  INV_X1 U43632 ( .A(n41213), .ZN(n40181) );
  NAND2_X1 U43633 ( .A1(n40181), .A2(n41210), .ZN(n40182) );
  INV_X1 U43635 ( .A(n40184), .ZN(n41215) );
  AND2_X1 U43636 ( .A1(n41215), .A2(n41207), .ZN(n40188) );
  OAI22_X1 U43637 ( .A1(n40186), .A2(n51430), .B1(n685), .B2(n51052), .ZN(
        n40187) );
  AND2_X1 U43638 ( .A1(n40188), .A2(n40187), .ZN(n40190) );
  AOI22_X1 U43639 ( .A1(n41196), .A2(n40662), .B1(n40664), .B2(n41207), .ZN(
        n40189) );
  OAI21_X2 U43640 ( .B1(n40191), .B2(n40190), .A(n40189), .ZN(n45306) );
  XNOR2_X1 U43641 ( .A(n45306), .B(n45097), .ZN(n44146) );
  XNOR2_X1 U43642 ( .A(n44146), .B(n43755), .ZN(n40209) );
  INV_X1 U43643 ( .A(n40192), .ZN(n40193) );
  INV_X1 U43644 ( .A(n40196), .ZN(n40197) );
  INV_X1 U43645 ( .A(n40198), .ZN(n40199) );
  NAND3_X1 U43646 ( .A1(n40200), .A2(n40199), .A3(n51233), .ZN(n40208) );
  INV_X1 U43647 ( .A(n40201), .ZN(n40202) );
  NAND4_X1 U43648 ( .A1(n40205), .A2(n40204), .A3(n40203), .A4(n40202), .ZN(
        n40206) );
  XNOR2_X1 U43649 ( .A(n40209), .B(n45303), .ZN(n42098) );
  INV_X1 U43650 ( .A(n41246), .ZN(n40213) );
  NAND2_X1 U43651 ( .A1(n3861), .A2(n3489), .ZN(n40708) );
  INV_X1 U43652 ( .A(n40708), .ZN(n40212) );
  NAND3_X1 U43653 ( .A1(n40213), .A2(n41234), .A3(n40212), .ZN(n40216) );
  INV_X1 U43654 ( .A(n41680), .ZN(n40215) );
  INV_X1 U43655 ( .A(n41684), .ZN(n40214) );
  NAND2_X1 U43656 ( .A1(n40215), .A2(n40214), .ZN(n41241) );
  INV_X1 U43658 ( .A(n52198), .ZN(n41237) );
  INV_X1 U43659 ( .A(n41681), .ZN(n41243) );
  NAND4_X1 U43660 ( .A1(n41227), .A2(n41234), .A3(n41683), .A4(n41673), .ZN(
        n40218) );
  OAI21_X1 U43661 ( .B1(n41237), .B2(n41243), .A(n40218), .ZN(n40219) );
  XNOR2_X1 U43662 ( .A(n40222), .B(n40221), .ZN(n40223) );
  XNOR2_X1 U43663 ( .A(n45314), .B(n40223), .ZN(n40224) );
  OR2_X1 U43664 ( .A1(n41544), .A2(n41554), .ZN(n40227) );
  NAND2_X1 U43665 ( .A1(n40936), .A2(n40989), .ZN(n40226) );
  INV_X1 U43666 ( .A(n41526), .ZN(n40225) );
  MUX2_X1 U43667 ( .A(n40227), .B(n40226), .S(n40225), .Z(n40237) );
  INV_X1 U43668 ( .A(n40228), .ZN(n40230) );
  NAND2_X1 U43669 ( .A1(n41553), .A2(n41394), .ZN(n40231) );
  NAND2_X1 U43670 ( .A1(n41554), .A2(n52120), .ZN(n41391) );
  NAND3_X1 U43671 ( .A1(n40230), .A2(n40229), .A3(n41391), .ZN(n40235) );
  INV_X1 U43672 ( .A(n41544), .ZN(n41543) );
  AND2_X1 U43673 ( .A1(n41554), .A2(n8754), .ZN(n40232) );
  NAND4_X1 U43674 ( .A1(n41543), .A2(n40232), .A3(n40231), .A4(n41394), .ZN(
        n40234) );
  NAND2_X1 U43675 ( .A1(n41539), .A2(n40986), .ZN(n41393) );
  INV_X1 U43676 ( .A(n41393), .ZN(n41525) );
  NAND2_X1 U43677 ( .A1(n41525), .A2(n41535), .ZN(n40233) );
  AND3_X1 U43678 ( .A1(n40235), .A2(n40234), .A3(n40233), .ZN(n40236) );
  NAND2_X2 U43679 ( .A1(n40236), .A2(n40237), .ZN(n45116) );
  XNOR2_X1 U43680 ( .A(n42098), .B(n40238), .ZN(n40286) );
  INV_X1 U43681 ( .A(n40921), .ZN(n41379) );
  NAND3_X1 U43682 ( .A1(n40924), .A2(n38901), .A3(n40239), .ZN(n42092) );
  NOR2_X1 U43683 ( .A1(n40967), .A2(n51853), .ZN(n40246) );
  NAND2_X1 U43684 ( .A1(n40241), .A2(n41380), .ZN(n40245) );
  INV_X1 U43685 ( .A(n40242), .ZN(n40244) );
  NAND2_X1 U43686 ( .A1(n41380), .A2(n3775), .ZN(n40243) );
  INV_X1 U43687 ( .A(n41944), .ZN(n40254) );
  NAND2_X1 U43688 ( .A1(n41934), .A2(n41940), .ZN(n40253) );
  NAND2_X1 U43689 ( .A1(n41942), .A2(n41931), .ZN(n41943) );
  INV_X1 U43690 ( .A(n41943), .ZN(n40252) );
  AOI21_X1 U43691 ( .B1(n40254), .B2(n40253), .A(n40252), .ZN(n40255) );
  XNOR2_X1 U43693 ( .A(n44042), .B(n44130), .ZN(n40283) );
  INV_X1 U43694 ( .A(n40257), .ZN(n42152) );
  INV_X1 U43696 ( .A(n40258), .ZN(n40264) );
  INV_X1 U43697 ( .A(n42156), .ZN(n41764) );
  NAND2_X1 U43698 ( .A1(n8332), .A2(n42136), .ZN(n42135) );
  NAND2_X1 U43699 ( .A1(n40264), .A2(n42135), .ZN(n40259) );
  NAND2_X1 U43700 ( .A1(n687), .A2(n51375), .ZN(n42146) );
  INV_X1 U43701 ( .A(n42146), .ZN(n40261) );
  INV_X1 U43702 ( .A(n42148), .ZN(n42749) );
  INV_X1 U43703 ( .A(n40262), .ZN(n40263) );
  OAI21_X1 U43704 ( .B1(n42157), .B2(n42145), .A(n40263), .ZN(n41762) );
  NAND2_X1 U43705 ( .A1(n42154), .A2(n41770), .ZN(n40882) );
  OAI21_X1 U43706 ( .B1(n42138), .B2(n42157), .A(n40882), .ZN(n41748) );
  NAND2_X1 U43707 ( .A1(n41762), .A2(n41748), .ZN(n40266) );
  NAND3_X1 U43708 ( .A1(n42158), .A2(n42145), .A3(n40264), .ZN(n40265) );
  NAND2_X1 U43709 ( .A1(n40268), .A2(n40267), .ZN(n40281) );
  NAND4_X2 U43712 ( .A1(n40281), .A2(n40279), .A3(n40280), .A4(n40278), .ZN(
        n45114) );
  XNOR2_X1 U43713 ( .A(n50987), .B(n45114), .ZN(n40282) );
  INV_X1 U43714 ( .A(n41159), .ZN(n40284) );
  XNOR2_X1 U43715 ( .A(n43148), .B(n40284), .ZN(n40285) );
  INV_X1 U43716 ( .A(n40288), .ZN(n40289) );
  AOI21_X1 U43717 ( .B1(n40290), .B2(n42049), .A(n40289), .ZN(n40301) );
  NAND2_X1 U43718 ( .A1(n42042), .A2(n596), .ZN(n40291) );
  NAND2_X1 U43719 ( .A1(n42443), .A2(n40291), .ZN(n40300) );
  OAI21_X1 U43720 ( .B1(n40294), .B2(n40293), .A(n40292), .ZN(n40299) );
  AOI22_X1 U43721 ( .A1(n40295), .A2(n480), .B1(n679), .B2(n42062), .ZN(n40297) );
  NAND4_X2 U43722 ( .A1(n40301), .A2(n40298), .A3(n40299), .A4(n40300), .ZN(
        n45358) );
  XNOR2_X1 U43723 ( .A(n46150), .B(n45358), .ZN(n40303) );
  XNOR2_X1 U43724 ( .A(n43609), .B(n45357), .ZN(n40302) );
  XNOR2_X1 U43725 ( .A(n40303), .B(n40302), .ZN(n40309) );
  XNOR2_X1 U43726 ( .A(n40305), .B(n40304), .ZN(n40306) );
  XNOR2_X1 U43727 ( .A(n43254), .B(n40306), .ZN(n40307) );
  XNOR2_X1 U43729 ( .A(n40309), .B(n40308), .ZN(n40326) );
  NAND2_X1 U43730 ( .A1(n40319), .A2(n40310), .ZN(n40313) );
  INV_X1 U43731 ( .A(n40311), .ZN(n40312) );
  NAND2_X1 U43732 ( .A1(n40313), .A2(n40312), .ZN(n40324) );
  NAND2_X1 U43733 ( .A1(n40317), .A2(n40316), .ZN(n40323) );
  NAND2_X1 U43734 ( .A1(n40318), .A2(n40565), .ZN(n40320) );
  MUX2_X1 U43735 ( .A(n40320), .B(n40319), .S(n52159), .Z(n40322) );
  XNOR2_X1 U43736 ( .A(n44182), .B(n4934), .ZN(n40325) );
  XNOR2_X1 U43737 ( .A(n40325), .B(n44373), .ZN(n41966) );
  XNOR2_X1 U43738 ( .A(n40326), .B(n41966), .ZN(n40394) );
  NAND3_X1 U43739 ( .A1(n40329), .A2(n40328), .A3(n40327), .ZN(n40332) );
  NAND3_X1 U43740 ( .A1(n52101), .A2(n40338), .A3(n40330), .ZN(n40331) );
  NAND3_X1 U43741 ( .A1(n40333), .A2(n40332), .A3(n40331), .ZN(n40347) );
  INV_X1 U43742 ( .A(n40337), .ZN(n40339) );
  OAI211_X1 U43743 ( .C1(n40341), .C2(n40340), .A(n40339), .B(n40338), .ZN(
        n40345) );
  NAND2_X1 U43744 ( .A1(n40343), .A2(n52101), .ZN(n40344) );
  INV_X1 U43745 ( .A(n41164), .ZN(n40348) );
  NAND2_X1 U43746 ( .A1(n41689), .A2(n40348), .ZN(n40351) );
  NAND3_X1 U43747 ( .A1(n41163), .A2(n41621), .A3(n41691), .ZN(n40350) );
  AND2_X1 U43748 ( .A1(n41702), .A2(n41692), .ZN(n41612) );
  NAND2_X1 U43749 ( .A1(n41612), .A2(n41695), .ZN(n40349) );
  INV_X1 U43750 ( .A(n41166), .ZN(n40352) );
  OAI21_X1 U43751 ( .B1(n41163), .B2(n40353), .A(n40352), .ZN(n40356) );
  AOI21_X1 U43752 ( .B1(n2179), .B2(n2867), .A(n41695), .ZN(n40354) );
  NAND2_X1 U43753 ( .A1(n40358), .A2(n41355), .ZN(n40752) );
  NAND3_X1 U43754 ( .A1(n40751), .A2(n41360), .A3(n39632), .ZN(n40363) );
  INV_X1 U43755 ( .A(n41353), .ZN(n40361) );
  OAI21_X1 U43756 ( .B1(n40361), .B2(n40360), .A(n40359), .ZN(n40362) );
  XNOR2_X1 U43757 ( .A(n46143), .B(n45467), .ZN(n43724) );
  XNOR2_X1 U43758 ( .A(n43724), .B(n45091), .ZN(n40393) );
  OR2_X1 U43759 ( .A1(n41902), .A2(n41317), .ZN(n40728) );
  INV_X1 U43760 ( .A(n40728), .ZN(n40365) );
  OAI21_X1 U43761 ( .B1(n40366), .B2(n40365), .A(n40727), .ZN(n40367) );
  NOR2_X1 U43762 ( .A1(n40730), .A2(n52215), .ZN(n40370) );
  INV_X1 U43763 ( .A(n40726), .ZN(n40369) );
  INV_X1 U43764 ( .A(n41320), .ZN(n40368) );
  AOI22_X1 U43765 ( .A1(n40371), .A2(n40370), .B1(n40369), .B2(n40368), .ZN(
        n40376) );
  INV_X1 U43766 ( .A(n40372), .ZN(n40374) );
  OAI21_X1 U43767 ( .B1(n41327), .B2(n40374), .A(n40373), .ZN(n40375) );
  AND2_X1 U43768 ( .A1(n40377), .A2(n682), .ZN(n40389) );
  NAND2_X1 U43769 ( .A1(n40378), .A2(n40389), .ZN(n40392) );
  AOI21_X1 U43770 ( .B1(n40381), .B2(n40380), .A(n40379), .ZN(n40391) );
  NAND2_X1 U43771 ( .A1(n40382), .A2(n41143), .ZN(n40383) );
  NAND3_X1 U43772 ( .A1(n40384), .A2(n40383), .A3(n41148), .ZN(n40387) );
  NAND3_X1 U43773 ( .A1(n41144), .A2(n40385), .A3(n41147), .ZN(n40386) );
  NAND3_X1 U43774 ( .A1(n40389), .A2(n677), .A3(n40388), .ZN(n40390) );
  XNOR2_X1 U43775 ( .A(n44098), .B(n40393), .ZN(n44378) );
  XNOR2_X1 U43776 ( .A(n40394), .B(n44378), .ZN(n40409) );
  OAI21_X1 U43777 ( .B1(n40436), .B2(n40403), .A(n40447), .ZN(n40398) );
  OAI22_X1 U43778 ( .A1(n40398), .A2(n40397), .B1(n6851), .B2(n40458), .ZN(
        n40399) );
  NOR2_X1 U43779 ( .A1(n40400), .A2(n40399), .ZN(n40407) );
  INV_X1 U43780 ( .A(n40401), .ZN(n40406) );
  INV_X1 U43781 ( .A(n40402), .ZN(n40444) );
  NOR2_X1 U43782 ( .A1(n40403), .A2(n40453), .ZN(n40460) );
  OAI21_X1 U43783 ( .B1(n40444), .B2(n40404), .A(n40460), .ZN(n40405) );
  INV_X1 U43784 ( .A(n43357), .ZN(n40408) );
  XNOR2_X1 U43785 ( .A(n44170), .B(n569), .ZN(n41408) );
  XNOR2_X2 U43786 ( .A(n40409), .B(n41408), .ZN(n46637) );
  INV_X1 U43787 ( .A(n41276), .ZN(n41285) );
  XNOR2_X1 U43788 ( .A(n52193), .B(n41292), .ZN(n40414) );
  INV_X1 U43789 ( .A(n40410), .ZN(n40411) );
  NAND3_X1 U43790 ( .A1(n40412), .A2(n40411), .A3(n41039), .ZN(n40413) );
  OAI211_X1 U43791 ( .C1(n40415), .C2(n40414), .A(n41028), .B(n40413), .ZN(
        n40416) );
  INV_X1 U43792 ( .A(n40416), .ZN(n40435) );
  INV_X1 U43793 ( .A(n40418), .ZN(n40419) );
  NAND2_X1 U43794 ( .A1(n40419), .A2(n41275), .ZN(n40426) );
  NAND4_X1 U43795 ( .A1(n40421), .A2(n41280), .A3(n41034), .A4(n41286), .ZN(
        n40425) );
  NAND3_X1 U43796 ( .A1(n40423), .A2(n41025), .A3(n41039), .ZN(n40424) );
  OR3_X1 U43797 ( .A1(n40429), .A2(n40428), .A3(n41039), .ZN(n40433) );
  NAND3_X1 U43798 ( .A1(n40431), .A2(n41276), .A3(n40430), .ZN(n40432) );
  AOI21_X1 U43799 ( .B1(n40437), .B2(n40436), .A(n40458), .ZN(n40438) );
  AND3_X1 U43800 ( .A1(n40441), .A2(n40440), .A3(n40439), .ZN(n40466) );
  INV_X1 U43801 ( .A(n40442), .ZN(n40443) );
  NAND3_X1 U43802 ( .A1(n40444), .A2(n40443), .A3(n40450), .ZN(n40452) );
  AND2_X1 U43803 ( .A1(n40445), .A2(n40453), .ZN(n40449) );
  OAI22_X1 U43804 ( .A1(n40447), .A2(n40456), .B1(n40446), .B2(n40450), .ZN(
        n40448) );
  OAI211_X1 U43805 ( .C1(n40450), .C2(n40458), .A(n40449), .B(n40448), .ZN(
        n40451) );
  AND2_X1 U43806 ( .A1(n40451), .A2(n40452), .ZN(n40465) );
  OR2_X1 U43807 ( .A1(n40458), .A2(n40453), .ZN(n40455) );
  OAI21_X1 U43808 ( .B1(n40459), .B2(n40455), .A(n40454), .ZN(n40457) );
  NAND2_X1 U43809 ( .A1(n40457), .A2(n40456), .ZN(n40464) );
  OAI211_X1 U43810 ( .C1(n40462), .C2(n40461), .A(n40460), .B(n40459), .ZN(
        n40463) );
  NAND2_X1 U43811 ( .A1(n40477), .A2(n41265), .ZN(n41121) );
  NAND2_X1 U43812 ( .A1(n40469), .A2(n41113), .ZN(n40472) );
  AND2_X1 U43813 ( .A1(n41113), .A2(n41256), .ZN(n41261) );
  NAND3_X1 U43814 ( .A1(n40482), .A2(n41124), .A3(n41261), .ZN(n40471) );
  OAI211_X1 U43815 ( .C1(n40473), .C2(n41121), .A(n40472), .B(n40471), .ZN(
        n40474) );
  INV_X1 U43816 ( .A(n40474), .ZN(n40492) );
  MUX2_X1 U43818 ( .A(n40486), .B(n40475), .S(n39593), .Z(n40491) );
  OAI21_X1 U43819 ( .B1(n41256), .B2(n41730), .A(n40476), .ZN(n40478) );
  NAND4_X1 U43820 ( .A1(n40478), .A2(n41263), .A3(n41110), .A4(n40477), .ZN(
        n40484) );
  AND2_X1 U43821 ( .A1(n41113), .A2(n41110), .ZN(n41120) );
  INV_X1 U43822 ( .A(n40479), .ZN(n40480) );
  NAND2_X1 U43823 ( .A1(n40480), .A2(n41735), .ZN(n40481) );
  NAND3_X1 U43824 ( .A1(n40482), .A2(n41120), .A3(n40481), .ZN(n40483) );
  AND2_X1 U43825 ( .A1(n40484), .A2(n40483), .ZN(n40490) );
  INV_X1 U43826 ( .A(n40485), .ZN(n40487) );
  NOR2_X1 U43827 ( .A1(n41256), .A2(n41112), .ZN(n41118) );
  INV_X1 U43828 ( .A(n41729), .ZN(n40488) );
  NAND4_X2 U43829 ( .A1(n40492), .A2(n40489), .A3(n40491), .A4(n40490), .ZN(
        n46058) );
  AOI22_X1 U43831 ( .A1(n40498), .A2(n40497), .B1(n40496), .B2(n41057), .ZN(
        n40519) );
  NAND4_X1 U43833 ( .A1(n40510), .A2(n40502), .A3(n41065), .A4(n41063), .ZN(
        n40503) );
  INV_X1 U43834 ( .A(n40506), .ZN(n40504) );
  NAND4_X1 U43835 ( .A1(n41052), .A2(n40504), .A3(n610), .A4(n41063), .ZN(
        n40507) );
  OAI22_X1 U43837 ( .A1(n40514), .A2(n40513), .B1(n40512), .B2(n40511), .ZN(
        n40515) );
  NAND2_X1 U43838 ( .A1(n40515), .A2(n41064), .ZN(n40518) );
  NAND2_X1 U43839 ( .A1(n41053), .A2(n41056), .ZN(n40517) );
  XNOR2_X1 U43840 ( .A(n40521), .B(n40520), .ZN(n40522) );
  XNOR2_X1 U43841 ( .A(n42170), .B(n40522), .ZN(n40523) );
  XNOR2_X1 U43842 ( .A(n44061), .B(n40523), .ZN(n40524) );
  NAND3_X1 U43843 ( .A1(n40541), .A2(n40525), .A3(n40529), .ZN(n40527) );
  NAND2_X1 U43844 ( .A1(n40874), .A2(n40526), .ZN(n40871) );
  AOI21_X1 U43845 ( .B1(n40527), .B2(n40871), .A(n40862), .ZN(n40539) );
  INV_X1 U43846 ( .A(n40529), .ZN(n40530) );
  NAND3_X1 U43847 ( .A1(n40531), .A2(n40530), .A3(n678), .ZN(n40532) );
  NOR2_X1 U43848 ( .A1(n40856), .A2(n40862), .ZN(n40536) );
  NAND3_X1 U43849 ( .A1(n40873), .A2(n40537), .A3(n40862), .ZN(n40538) );
  NAND2_X1 U43850 ( .A1(n40857), .A2(n40868), .ZN(n40547) );
  INV_X1 U43851 ( .A(n40873), .ZN(n40545) );
  INV_X1 U43852 ( .A(n40541), .ZN(n40542) );
  NAND4_X1 U43853 ( .A1(n40545), .A2(n40544), .A3(n40543), .A4(n40542), .ZN(
        n40546) );
  XNOR2_X1 U43854 ( .A(n43909), .B(n43781), .ZN(n40580) );
  OAI21_X1 U43855 ( .B1(n40549), .B2(n4950), .A(n40563), .ZN(n40551) );
  AOI21_X1 U43856 ( .B1(n40566), .B2(n40564), .A(n52159), .ZN(n40550) );
  INV_X1 U43857 ( .A(n40563), .ZN(n40553) );
  OAI21_X1 U43858 ( .B1(n40553), .B2(n4000), .A(n2597), .ZN(n40562) );
  OAI21_X1 U43859 ( .B1(n40564), .B2(n40565), .A(n4950), .ZN(n40557) );
  NAND4_X1 U43860 ( .A1(n40557), .A2(n4000), .A3(n40556), .A4(n40555), .ZN(
        n40561) );
  NAND2_X1 U43861 ( .A1(n40559), .A2(n40558), .ZN(n40560) );
  OAI211_X1 U43862 ( .C1(n40566), .C2(n40565), .A(n40564), .B(n40563), .ZN(
        n40577) );
  NAND2_X1 U43863 ( .A1(n7848), .A2(n40567), .ZN(n40569) );
  NAND3_X1 U43864 ( .A1(n40573), .A2(n52159), .A3(n40571), .ZN(n40574) );
  OAI211_X1 U43865 ( .C1(n40577), .C2(n40576), .A(n40575), .B(n40574), .ZN(
        n40578) );
  XNOR2_X1 U43866 ( .A(n40580), .B(n45432), .ZN(n40581) );
  NOR2_X1 U43867 ( .A1(n432), .A2(n40776), .ZN(n40582) );
  NAND2_X1 U43868 ( .A1(n40583), .A2(n40582), .ZN(n40772) );
  NOR3_X1 U43869 ( .A1(n40777), .A2(n6046), .A3(n40785), .ZN(n40584) );
  NOR2_X1 U43870 ( .A1(n40774), .A2(n40775), .ZN(n40587) );
  NAND4_X1 U43871 ( .A1(n40587), .A2(n426), .A3(n431), .A4(n40768), .ZN(n40588) );
  MUX2_X1 U43872 ( .A(n40784), .B(n40590), .S(n431), .Z(n40602) );
  NOR2_X1 U43873 ( .A1(n40591), .A2(n40768), .ZN(n40595) );
  NAND2_X1 U43874 ( .A1(n40592), .A2(n426), .ZN(n40593) );
  OAI21_X1 U43875 ( .B1(n40593), .B2(n432), .A(n681), .ZN(n40594) );
  AOI22_X1 U43876 ( .A1(n40600), .A2(n40595), .B1(n40594), .B2(n40783), .ZN(
        n40601) );
  INV_X1 U43877 ( .A(n40596), .ZN(n40597) );
  NAND3_X1 U43878 ( .A1(n40782), .A2(n6046), .A3(n40597), .ZN(n40599) );
  INV_X1 U43879 ( .A(n41104), .ZN(n40605) );
  NAND3_X1 U43880 ( .A1(n41977), .A2(n40608), .A3(n40605), .ZN(n40612) );
  INV_X1 U43881 ( .A(n40606), .ZN(n40607) );
  NAND4_X1 U43882 ( .A1(n40608), .A2(n40607), .A3(n41645), .A4(n41975), .ZN(
        n40611) );
  INV_X1 U43883 ( .A(n40609), .ZN(n40610) );
  AOI21_X1 U43884 ( .B1(n40612), .B2(n40611), .A(n40610), .ZN(n40613) );
  NOR2_X1 U43885 ( .A1(n40614), .A2(n40613), .ZN(n40629) );
  NAND3_X1 U43886 ( .A1(n41977), .A2(n40623), .A3(n41975), .ZN(n40620) );
  OR2_X1 U43887 ( .A1(n40615), .A2(n41642), .ZN(n40619) );
  AOI21_X1 U43888 ( .B1(n40617), .B2(n41642), .A(n41975), .ZN(n40616) );
  OAI211_X1 U43889 ( .C1(n40623), .C2(n40617), .A(n40616), .B(n41647), .ZN(
        n40618) );
  OAI211_X1 U43890 ( .C1(n40620), .C2(n41641), .A(n40619), .B(n40618), .ZN(
        n40621) );
  INV_X1 U43891 ( .A(n40621), .ZN(n40628) );
  NAND2_X1 U43892 ( .A1(n40622), .A2(n41977), .ZN(n40627) );
  INV_X1 U43893 ( .A(n40623), .ZN(n40624) );
  NOR2_X1 U43894 ( .A1(n41977), .A2(n40624), .ZN(n40625) );
  OAI21_X1 U43895 ( .B1(n41638), .B2(n40625), .A(n52080), .ZN(n40626) );
  XNOR2_X1 U43896 ( .A(n43197), .B(n43524), .ZN(n43173) );
  XNOR2_X1 U43897 ( .A(n44202), .B(n43173), .ZN(n40630) );
  INV_X1 U43899 ( .A(n46630), .ZN(n40950) );
  INV_X1 U43900 ( .A(n42870), .ZN(n40641) );
  AND2_X1 U43901 ( .A1(n40634), .A2(n42111), .ZN(n43672) );
  INV_X1 U43902 ( .A(n43672), .ZN(n40635) );
  OR2_X1 U43903 ( .A1(n40636), .A2(n41796), .ZN(n40638) );
  XNOR2_X1 U43904 ( .A(n40641), .B(n45393), .ZN(n43127) );
  XNOR2_X1 U43905 ( .A(n43127), .B(n40642), .ZN(n40766) );
  INV_X1 U43906 ( .A(n40643), .ZN(n41429) );
  NAND2_X1 U43907 ( .A1(n40645), .A2(n40644), .ZN(n40660) );
  NOR2_X1 U43908 ( .A1(n40647), .A2(n41436), .ZN(n40648) );
  AOI22_X1 U43909 ( .A1(n40649), .A2(n41433), .B1(n40648), .B2(n41451), .ZN(
        n40659) );
  OAI211_X1 U43910 ( .C1(n41450), .C2(n40651), .A(n40653), .B(n40650), .ZN(
        n40658) );
  NAND2_X1 U43911 ( .A1(n40653), .A2(n40652), .ZN(n40656) );
  NAND4_X1 U43912 ( .A1(n40656), .A2(n40655), .A3(n40654), .A4(n41436), .ZN(
        n40657) );
  NAND4_X2 U43913 ( .A1(n40660), .A2(n40659), .A3(n40658), .A4(n40657), .ZN(
        n44900) );
  MUX2_X1 U43914 ( .A(n41210), .B(n41202), .S(n41211), .Z(n40661) );
  AND2_X1 U43915 ( .A1(n685), .A2(n40665), .ZN(n40667) );
  INV_X1 U43916 ( .A(n41203), .ZN(n40666) );
  AOI21_X1 U43917 ( .B1(n41200), .B2(n40667), .A(n40666), .ZN(n40671) );
  NOR2_X1 U43918 ( .A1(n51430), .A2(n41207), .ZN(n41194) );
  OAI21_X1 U43919 ( .B1(n41194), .B2(n41212), .A(n40668), .ZN(n40670) );
  XNOR2_X2 U43920 ( .A(n44900), .B(n51406), .ZN(n45389) );
  NAND2_X1 U43922 ( .A1(n40677), .A2(n40676), .ZN(n40678) );
  NAND2_X1 U43923 ( .A1(n40682), .A2(n40685), .ZN(n40688) );
  NAND3_X1 U43924 ( .A1(n40685), .A2(n40684), .A3(n40683), .ZN(n40687) );
  MUX2_X1 U43925 ( .A(n40688), .B(n40687), .S(n51022), .Z(n40697) );
  NAND2_X1 U43926 ( .A1(n40690), .A2(n40689), .ZN(n40695) );
  NAND3_X1 U43927 ( .A1(n40693), .A2(n40692), .A3(n40691), .ZN(n40694) );
  NAND4_X1 U43928 ( .A1(n40697), .A2(n40696), .A3(n40695), .A4(n40694), .ZN(
        n40698) );
  NAND2_X1 U43929 ( .A1(n42018), .A2(n42020), .ZN(n42014) );
  NAND3_X1 U43930 ( .A1(n41997), .A2(n41581), .A3(n42018), .ZN(n41583) );
  NOR2_X1 U43931 ( .A1(n42018), .A2(n42020), .ZN(n41415) );
  NAND4_X1 U43932 ( .A1(n41415), .A2(n42011), .A3(n41587), .A4(n42006), .ZN(
        n40702) );
  NOR2_X1 U43933 ( .A1(n42018), .A2(n42010), .ZN(n41416) );
  NOR2_X1 U43934 ( .A1(n42006), .A2(n41997), .ZN(n41511) );
  NAND2_X1 U43935 ( .A1(n41416), .A2(n41511), .ZN(n40701) );
  AND2_X1 U43936 ( .A1(n40702), .A2(n40701), .ZN(n40706) );
  NAND2_X1 U43937 ( .A1(n41997), .A2(n42010), .ZN(n42019) );
  OR2_X1 U43938 ( .A1(n42018), .A2(n41587), .ZN(n41575) );
  OAI22_X1 U43939 ( .A1(n41588), .A2(n41576), .B1(n41575), .B2(n42006), .ZN(
        n40703) );
  NAND2_X1 U43940 ( .A1(n40703), .A2(n41997), .ZN(n40704) );
  NAND4_X2 U43941 ( .A1(n40704), .A2(n40705), .A3(n40707), .A4(n40706), .ZN(
        n44017) );
  NOR2_X1 U43942 ( .A1(n41685), .A2(n41679), .ZN(n41236) );
  NAND2_X1 U43943 ( .A1(n41246), .A2(n41236), .ZN(n40715) );
  NAND2_X1 U43944 ( .A1(n52198), .A2(n6335), .ZN(n40709) );
  NAND4_X1 U43948 ( .A1(n52198), .A2(n41245), .A3(n41685), .A4(n41670), .ZN(
        n40712) );
  NAND4_X1 U43949 ( .A1(n40715), .A2(n40714), .A3(n40713), .A4(n40712), .ZN(
        n40721) );
  OAI21_X1 U43951 ( .B1(n52198), .B2(n41685), .A(n41238), .ZN(n40718) );
  NAND3_X1 U43952 ( .A1(n41683), .A2(n40718), .A3(n41245), .ZN(n40719) );
  XNOR2_X1 U43953 ( .A(n40722), .B(n45389), .ZN(n44291) );
  AND3_X1 U43954 ( .A1(n40725), .A2(n40724), .A3(n40723), .ZN(n40735) );
  NAND2_X1 U43955 ( .A1(n40730), .A2(n52214), .ZN(n40731) );
  OAI22_X1 U43956 ( .A1(n41329), .A2(n41320), .B1(n40732), .B2(n40731), .ZN(
        n40733) );
  NAND2_X1 U43957 ( .A1(n40733), .A2(n41328), .ZN(n40734) );
  NAND2_X1 U43958 ( .A1(n40737), .A2(n40736), .ZN(n40739) );
  NOR2_X1 U43960 ( .A1(n41354), .A2(n41348), .ZN(n40742) );
  AND2_X1 U43961 ( .A1(n40740), .A2(n41352), .ZN(n40741) );
  AOI22_X1 U43962 ( .A1(n52049), .A2(n40742), .B1(n41345), .B2(n40741), .ZN(
        n40747) );
  NAND4_X1 U43963 ( .A1(n40748), .A2(n40747), .A3(n40746), .A4(n40745), .ZN(
        n40756) );
  INV_X1 U43964 ( .A(n39632), .ZN(n40754) );
  NAND2_X1 U43965 ( .A1(n40749), .A2(n41348), .ZN(n40750) );
  NOR2_X1 U43966 ( .A1(n40751), .A2(n40750), .ZN(n40753) );
  MUX2_X1 U43967 ( .A(n40754), .B(n40753), .S(n40752), .Z(n40755) );
  XNOR2_X1 U43969 ( .A(n41629), .B(n4800), .ZN(n43291) );
  XNOR2_X1 U43970 ( .A(n42067), .B(n43291), .ZN(n40763) );
  BUF_X2 U43971 ( .A(n40757), .Z(n44301) );
  XNOR2_X1 U43972 ( .A(n40759), .B(n40758), .ZN(n40760) );
  XNOR2_X1 U43973 ( .A(n43973), .B(n40760), .ZN(n40761) );
  XNOR2_X1 U43974 ( .A(n44301), .B(n40761), .ZN(n40762) );
  XNOR2_X1 U43975 ( .A(n40763), .B(n40762), .ZN(n40764) );
  XNOR2_X1 U43976 ( .A(n44291), .B(n40764), .ZN(n40765) );
  XNOR2_X1 U43977 ( .A(n45269), .B(n51681), .ZN(n45412) );
  NAND2_X1 U43978 ( .A1(n40769), .A2(n40778), .ZN(n40770) );
  NAND2_X1 U43979 ( .A1(n40771), .A2(n40770), .ZN(n40773) );
  NAND2_X1 U43980 ( .A1(n40773), .A2(n40772), .ZN(n40793) );
  AOI21_X1 U43981 ( .B1(n426), .B2(n40775), .A(n40774), .ZN(n40780) );
  NAND4_X1 U43982 ( .A1(n432), .A2(n40778), .A3(n40777), .A4(n40776), .ZN(
        n40779) );
  NAND3_X1 U43983 ( .A1(n40787), .A2(n40786), .A3(n40785), .ZN(n40788) );
  NAND3_X1 U43984 ( .A1(n40790), .A2(n40789), .A3(n40788), .ZN(n40791) );
  AOI21_X2 U43985 ( .B1(n40793), .B2(n426), .A(n40791), .ZN(n43236) );
  AOI22_X1 U43986 ( .A1(n40794), .A2(n609), .B1(n41010), .B2(n41009), .ZN(
        n40813) );
  NAND2_X1 U43987 ( .A1(n40795), .A2(n5911), .ZN(n40798) );
  NAND2_X1 U43988 ( .A1(n43323), .A2(n41004), .ZN(n40796) );
  NAND3_X1 U43989 ( .A1(n40798), .A2(n40797), .A3(n40796), .ZN(n40804) );
  NAND2_X1 U43990 ( .A1(n40800), .A2(n40799), .ZN(n40803) );
  AND2_X1 U43991 ( .A1(n51358), .A2(n43327), .ZN(n43330) );
  NAND2_X1 U43992 ( .A1(n43330), .A2(n40801), .ZN(n40802) );
  AND3_X1 U43993 ( .A1(n40804), .A2(n40803), .A3(n40802), .ZN(n40812) );
  AND2_X1 U43994 ( .A1(n43329), .A2(n41004), .ZN(n40805) );
  AOI22_X1 U43995 ( .A1(n43335), .A2(n43330), .B1(n40806), .B2(n40805), .ZN(
        n40810) );
  OAI22_X1 U43996 ( .A1(n43325), .A2(n43323), .B1(n40807), .B2(n41013), .ZN(
        n40808) );
  NAND2_X1 U43997 ( .A1(n40808), .A2(n43329), .ZN(n40809) );
  AND2_X1 U43998 ( .A1(n40809), .A2(n40810), .ZN(n40811) );
  NOR2_X1 U43999 ( .A1(n40816), .A2(n40815), .ZN(n40821) );
  NOR2_X1 U44000 ( .A1(n40818), .A2(n40817), .ZN(n40819) );
  AOI22_X1 U44001 ( .A1(n675), .A2(n40821), .B1(n40820), .B2(n40819), .ZN(
        n40844) );
  XNOR2_X1 U44002 ( .A(n40823), .B(n40822), .ZN(n40827) );
  INV_X1 U44003 ( .A(n40824), .ZN(n40825) );
  NAND3_X1 U44004 ( .A1(n40827), .A2(n40826), .A3(n40825), .ZN(n40843) );
  NAND3_X1 U44005 ( .A1(n7488), .A2(n40835), .A3(n40828), .ZN(n40834) );
  INV_X1 U44006 ( .A(n40831), .ZN(n40832) );
  NAND3_X1 U44007 ( .A1(n40834), .A2(n40833), .A3(n40832), .ZN(n40842) );
  NAND2_X1 U44008 ( .A1(n40836), .A2(n40835), .ZN(n40837) );
  OAI211_X1 U44009 ( .C1(n40840), .C2(n40839), .A(n51455), .B(n40837), .ZN(
        n40841) );
  XNOR2_X1 U44010 ( .A(n48843), .B(n4645), .ZN(n40845) );
  XNOR2_X1 U44011 ( .A(n42643), .B(n40845), .ZN(n40846) );
  XNOR2_X1 U44012 ( .A(n42729), .B(n40846), .ZN(n41310) );
  XNOR2_X1 U44013 ( .A(n41310), .B(n45412), .ZN(n40855) );
  XOR2_X1 U44014 ( .A(n42025), .B(n40847), .Z(n40848) );
  XNOR2_X1 U44015 ( .A(n40849), .B(n40848), .ZN(n40850) );
  XNOR2_X1 U44016 ( .A(n44879), .B(n40850), .ZN(n40851) );
  XNOR2_X1 U44017 ( .A(n40852), .B(n40851), .ZN(n40853) );
  XNOR2_X1 U44019 ( .A(n40853), .B(n43141), .ZN(n40854) );
  XNOR2_X1 U44020 ( .A(n40855), .B(n40854), .ZN(n40949) );
  AOI21_X1 U44021 ( .B1(n40857), .B2(n40856), .A(n678), .ZN(n40858) );
  OAI21_X1 U44022 ( .B1(n40859), .B2(n40858), .A(n40862), .ZN(n40880) );
  NAND2_X1 U44023 ( .A1(n40861), .A2(n40860), .ZN(n40867) );
  XNOR2_X1 U44024 ( .A(n40862), .B(n40863), .ZN(n40865) );
  NAND3_X1 U44025 ( .A1(n40865), .A2(n40864), .A3(n678), .ZN(n40866) );
  AND2_X1 U44026 ( .A1(n40868), .A2(n40869), .ZN(n40870) );
  AOI22_X1 U44027 ( .A1(n40873), .A2(n40872), .B1(n40871), .B2(n40870), .ZN(
        n40878) );
  NAND2_X1 U44028 ( .A1(n40876), .A2(n40875), .ZN(n40877) );
  XNOR2_X1 U44029 ( .A(n40881), .B(n46111), .ZN(n42035) );
  NAND2_X1 U44030 ( .A1(n42136), .A2(n42157), .ZN(n42155) );
  OAI211_X1 U44031 ( .C1(n42146), .C2(n52092), .A(n42131), .B(n42155), .ZN(
        n40884) );
  OAI21_X1 U44032 ( .B1(n42155), .B2(n41764), .A(n40882), .ZN(n40883) );
  NAND2_X1 U44033 ( .A1(n40884), .A2(n40883), .ZN(n40891) );
  AND2_X1 U44034 ( .A1(n52092), .A2(n42154), .ZN(n41773) );
  NOR2_X1 U44035 ( .A1(n42154), .A2(n51375), .ZN(n40885) );
  AOI22_X1 U44036 ( .A1(n41773), .A2(n42146), .B1(n40885), .B2(n42153), .ZN(
        n40890) );
  NOR2_X1 U44037 ( .A1(n52092), .A2(n42131), .ZN(n42151) );
  AOI22_X1 U44038 ( .A1(n42144), .A2(n41770), .B1(n40886), .B2(n42151), .ZN(
        n40889) );
  NAND2_X1 U44039 ( .A1(n40887), .A2(n42158), .ZN(n40888) );
  XNOR2_X1 U44041 ( .A(n42035), .B(n43143), .ZN(n40948) );
  NOR2_X1 U44042 ( .A1(n40906), .A2(n40892), .ZN(n40894) );
  AOI22_X1 U44043 ( .A1(n40895), .A2(n40894), .B1(n8708), .B2(n40911), .ZN(
        n40915) );
  NOR2_X1 U44044 ( .A1(n40905), .A2(n40906), .ZN(n40898) );
  AOI22_X1 U44045 ( .A1(n40898), .A2(n40903), .B1(n40897), .B2(n40896), .ZN(
        n40914) );
  INV_X1 U44046 ( .A(n40899), .ZN(n40902) );
  NAND3_X1 U44047 ( .A1(n40902), .A2(n40901), .A3(n40900), .ZN(n40908) );
  OR2_X1 U44048 ( .A1(n40904), .A2(n40903), .ZN(n40907) );
  NAND4_X1 U44049 ( .A1(n40908), .A2(n40907), .A3(n40906), .A4(n40905), .ZN(
        n40913) );
  OAI211_X1 U44050 ( .C1(n40911), .C2(n40910), .A(n2616), .B(n40909), .ZN(
        n40912) );
  INV_X1 U44051 ( .A(n40953), .ZN(n40955) );
  OAI22_X1 U44052 ( .A1(n40917), .A2(n40916), .B1(n38901), .B2(n40955), .ZN(
        n40920) );
  NAND2_X1 U44053 ( .A1(n40970), .A2(n51853), .ZN(n40918) );
  NOR2_X1 U44054 ( .A1(n40921), .A2(n40918), .ZN(n40919) );
  NOR2_X1 U44055 ( .A1(n40920), .A2(n40919), .ZN(n40930) );
  INV_X1 U44056 ( .A(n40965), .ZN(n40929) );
  AOI21_X1 U44057 ( .B1(n51394), .B2(n41374), .A(n41380), .ZN(n40923) );
  AND2_X1 U44058 ( .A1(n51853), .A2(n40972), .ZN(n41382) );
  INV_X1 U44059 ( .A(n41382), .ZN(n40922) );
  OR2_X1 U44060 ( .A1(n40923), .A2(n40922), .ZN(n40928) );
  OAI211_X1 U44061 ( .C1(n41375), .C2(n41380), .A(n40957), .B(n38901), .ZN(
        n40926) );
  AOI21_X1 U44062 ( .B1(n40959), .B2(n41378), .A(n40970), .ZN(n40925) );
  NAND3_X1 U44063 ( .A1(n40926), .A2(n40925), .A3(n40924), .ZN(n40927) );
  NOR2_X1 U44064 ( .A1(n52120), .A2(n40986), .ZN(n40931) );
  NOR2_X1 U44065 ( .A1(n40932), .A2(n40931), .ZN(n40934) );
  NOR2_X1 U44066 ( .A1(n41544), .A2(n41393), .ZN(n40933) );
  AOI22_X1 U44067 ( .A1(n41388), .A2(n40934), .B1(n40933), .B2(n41526), .ZN(
        n40947) );
  NAND2_X1 U44068 ( .A1(n40936), .A2(n40935), .ZN(n40946) );
  NAND2_X1 U44069 ( .A1(n41539), .A2(n41395), .ZN(n40988) );
  NOR2_X1 U44070 ( .A1(n41544), .A2(n40988), .ZN(n41531) );
  OAI21_X1 U44071 ( .B1(n41530), .B2(n40986), .A(n41393), .ZN(n40937) );
  OAI21_X1 U44072 ( .B1(n41531), .B2(n40937), .A(n41554), .ZN(n40945) );
  OAI21_X1 U44073 ( .B1(n41540), .B2(n40989), .A(n40941), .ZN(n40942) );
  NAND4_X2 U44074 ( .A1(n40947), .A2(n40945), .A3(n40946), .A4(n40944), .ZN(
        n46112) );
  XNOR2_X1 U44075 ( .A(n40948), .B(n42587), .ZN(n45063) );
  XNOR2_X1 U44076 ( .A(n40949), .B(n45063), .ZN(n40951) );
  NAND2_X1 U44078 ( .A1(n40950), .A2(n46631), .ZN(n44424) );
  INV_X1 U44079 ( .A(n46636), .ZN(n46627) );
  OR2_X1 U44080 ( .A1(n44652), .A2(n6741), .ZN(n44864) );
  INV_X1 U44081 ( .A(n44869), .ZN(n41132) );
  INV_X1 U44082 ( .A(n46631), .ZN(n44872) );
  OR2_X1 U44083 ( .A1(n44654), .A2(n46637), .ZN(n46641) );
  NAND2_X1 U44084 ( .A1(n46637), .A2(n46642), .ZN(n40952) );
  OR2_X1 U44085 ( .A1(n45757), .A2(n40952), .ZN(n44420) );
  OAI211_X1 U44086 ( .C1(n40955), .C2(n41372), .A(n41386), .B(n40954), .ZN(
        n40956) );
  INV_X1 U44087 ( .A(n40956), .ZN(n40978) );
  INV_X1 U44088 ( .A(n40957), .ZN(n40964) );
  NAND3_X1 U44089 ( .A1(n40958), .A2(n40970), .A3(n40967), .ZN(n40962) );
  NAND2_X1 U44091 ( .A1(n40966), .A2(n51853), .ZN(n40969) );
  MUX2_X1 U44092 ( .A(n40969), .B(n40968), .S(n38901), .Z(n40976) );
  INV_X1 U44093 ( .A(n40970), .ZN(n40971) );
  NAND2_X1 U44094 ( .A1(n40974), .A2(n51853), .ZN(n40975) );
  XNOR2_X2 U44096 ( .A(n45484), .B(n43318), .ZN(n46081) );
  XNOR2_X1 U44097 ( .A(n46081), .B(n40979), .ZN(n41002) );
  OR2_X1 U44098 ( .A1(n41544), .A2(n52120), .ZN(n40982) );
  OAI21_X1 U44099 ( .B1(n41524), .B2(n52120), .A(n41535), .ZN(n40980) );
  OAI22_X1 U44100 ( .A1(n40982), .A2(n40989), .B1(n41554), .B2(n40980), .ZN(
        n40985) );
  NOR2_X1 U44101 ( .A1(n40981), .A2(n41390), .ZN(n40984) );
  INV_X1 U44102 ( .A(n40982), .ZN(n40983) );
  OAI22_X1 U44103 ( .A1(n40985), .A2(n40984), .B1(n40983), .B2(n41394), .ZN(
        n40994) );
  AND3_X1 U44104 ( .A1(n41544), .A2(n41554), .A3(n40986), .ZN(n41533) );
  OAI21_X1 U44106 ( .B1(n40990), .B2(n40989), .A(n40988), .ZN(n40991) );
  NAND2_X1 U44107 ( .A1(n40991), .A2(n41540), .ZN(n40993) );
  NAND4_X1 U44108 ( .A1(n41544), .A2(n41524), .A3(n52120), .A4(n8754), .ZN(
        n40992) );
  XNOR2_X1 U44109 ( .A(n40996), .B(n40995), .ZN(n40997) );
  XNOR2_X1 U44110 ( .A(n43584), .B(n40997), .ZN(n41000) );
  INV_X1 U44111 ( .A(n44962), .ZN(n40999) );
  XNOR2_X1 U44112 ( .A(n41000), .B(n40999), .ZN(n41001) );
  XNOR2_X1 U44113 ( .A(n41002), .B(n41001), .ZN(n41023) );
  OAI21_X1 U44114 ( .B1(n51146), .B2(n41004), .A(n41003), .ZN(n43342) );
  OAI211_X1 U44115 ( .C1(n41007), .C2(n41006), .A(n43326), .B(n43342), .ZN(
        n41022) );
  NOR2_X1 U44116 ( .A1(n43323), .A2(n41013), .ZN(n43336) );
  OAI21_X1 U44117 ( .B1(n43336), .B2(n43327), .A(n43335), .ZN(n41012) );
  NAND2_X1 U44118 ( .A1(n41009), .A2(n41008), .ZN(n43339) );
  NAND2_X1 U44119 ( .A1(n41011), .A2(n41010), .ZN(n43338) );
  AND3_X1 U44120 ( .A1(n41012), .A2(n43339), .A3(n43338), .ZN(n41021) );
  INV_X1 U44121 ( .A(n43336), .ZN(n41016) );
  NAND3_X1 U44122 ( .A1(n43323), .A2(n41013), .A3(n43327), .ZN(n41014) );
  OAI21_X1 U44123 ( .B1(n41016), .B2(n41015), .A(n41014), .ZN(n41018) );
  NAND2_X1 U44124 ( .A1(n41018), .A2(n51357), .ZN(n41019) );
  XNOR2_X1 U44126 ( .A(n43890), .B(n45339), .ZN(n43098) );
  XNOR2_X1 U44127 ( .A(n43349), .B(n43098), .ZN(n45476) );
  XNOR2_X1 U44128 ( .A(n41023), .B(n45476), .ZN(n41130) );
  INV_X1 U44129 ( .A(n41024), .ZN(n41027) );
  NAND2_X1 U44130 ( .A1(n41025), .A2(n41276), .ZN(n41026) );
  NAND3_X1 U44131 ( .A1(n41028), .A2(n41027), .A3(n41026), .ZN(n41032) );
  NAND3_X1 U44132 ( .A1(n41034), .A2(n41276), .A3(n41291), .ZN(n41030) );
  NAND3_X1 U44133 ( .A1(n41032), .A2(n41031), .A3(n41030), .ZN(n41044) );
  OAI22_X1 U44134 ( .A1(n41274), .A2(n41035), .B1(n8613), .B2(n41034), .ZN(
        n41038) );
  OR2_X1 U44135 ( .A1(n41276), .A2(n41286), .ZN(n41036) );
  AOI21_X1 U44136 ( .B1(n8613), .B2(n41282), .A(n41036), .ZN(n41037) );
  NOR2_X1 U44137 ( .A1(n41039), .A2(n41286), .ZN(n41041) );
  AOI22_X1 U44138 ( .A1(n41041), .A2(n41040), .B1(n41278), .B2(n41039), .ZN(
        n41042) );
  XNOR2_X1 U44139 ( .A(n44164), .B(n43102), .ZN(n41072) );
  INV_X1 U44140 ( .A(n41051), .ZN(n41046) );
  NOR2_X1 U44141 ( .A1(n41047), .A2(n41065), .ZN(n41048) );
  AOI21_X1 U44142 ( .B1(n41050), .B2(n41049), .A(n41048), .ZN(n41070) );
  OAI21_X1 U44143 ( .B1(n41056), .B2(n41065), .A(n41054), .ZN(n41062) );
  INV_X1 U44144 ( .A(n41055), .ZN(n41061) );
  INV_X1 U44145 ( .A(n41056), .ZN(n41059) );
  NAND3_X1 U44146 ( .A1(n41059), .A2(n41058), .A3(n41057), .ZN(n41060) );
  NAND3_X1 U44147 ( .A1(n41062), .A2(n41061), .A3(n41060), .ZN(n41068) );
  OAI211_X1 U44148 ( .C1(n41066), .C2(n41065), .A(n41064), .B(n41063), .ZN(
        n41067) );
  INV_X1 U44149 ( .A(n44153), .ZN(n41071) );
  XNOR2_X1 U44150 ( .A(n41072), .B(n41071), .ZN(n41109) );
  NAND2_X1 U44151 ( .A1(n41074), .A2(n41073), .ZN(n41075) );
  NAND2_X1 U44152 ( .A1(n41076), .A2(n41075), .ZN(n41092) );
  INV_X1 U44153 ( .A(n41077), .ZN(n41078) );
  OAI21_X1 U44154 ( .B1(n8316), .B2(n41079), .A(n41085), .ZN(n41080) );
  OAI211_X1 U44155 ( .C1(n41088), .C2(n41085), .A(n41084), .B(n41083), .ZN(
        n41090) );
  OAI21_X1 U44156 ( .B1(n41088), .B2(n41087), .A(n41086), .ZN(n41089) );
  OAI21_X1 U44157 ( .B1(n41977), .B2(n41985), .A(n41093), .ZN(n41094) );
  INV_X1 U44158 ( .A(n41095), .ZN(n41097) );
  NOR2_X1 U44159 ( .A1(n41096), .A2(n41646), .ZN(n41649) );
  NAND2_X1 U44160 ( .A1(n41097), .A2(n41649), .ZN(n41100) );
  INV_X1 U44161 ( .A(n41101), .ZN(n41102) );
  NAND3_X1 U44162 ( .A1(n41102), .A2(n41645), .A3(n41647), .ZN(n41107) );
  INV_X1 U44163 ( .A(n41644), .ZN(n41105) );
  OAI21_X1 U44164 ( .B1(n41640), .B2(n41105), .A(n41978), .ZN(n41106) );
  XNOR2_X2 U44165 ( .A(n41956), .B(n44951), .ZN(n45068) );
  XNOR2_X1 U44166 ( .A(n41109), .B(n45068), .ZN(n43322) );
  OR2_X1 U44167 ( .A1(n41111), .A2(n41110), .ZN(n41262) );
  NAND3_X1 U44168 ( .A1(n41725), .A2(n41113), .A3(n41112), .ZN(n41114) );
  OAI21_X1 U44169 ( .B1(n41115), .B2(n41262), .A(n41114), .ZN(n41116) );
  INV_X1 U44171 ( .A(n41118), .ZN(n41119) );
  OAI21_X1 U44172 ( .B1(n41124), .B2(n41119), .A(n41262), .ZN(n41122) );
  AOI22_X1 U44173 ( .A1(n41736), .A2(n41122), .B1(n41121), .B2(n41120), .ZN(
        n41127) );
  NAND4_X1 U44174 ( .A1(n41728), .A2(n41124), .A3(n41123), .A4(n41735), .ZN(
        n41125) );
  XNOR2_X1 U44175 ( .A(n42979), .B(n43889), .ZN(n44079) );
  XNOR2_X1 U44176 ( .A(n42504), .B(n44079), .ZN(n41129) );
  XNOR2_X2 U44177 ( .A(n41130), .B(n8762), .ZN(n46635) );
  OAI211_X1 U44178 ( .C1(n44872), .C2(n46641), .A(n44420), .B(n47909), .ZN(
        n41131) );
  OAI21_X1 U44179 ( .B1(n44423), .B2(n45761), .A(n44868), .ZN(n41138) );
  NAND2_X1 U44180 ( .A1(n44652), .A2(n44873), .ZN(n41134) );
  NAND3_X1 U44181 ( .A1(n46635), .A2(n41134), .A3(n6741), .ZN(n41137) );
  NAND2_X1 U44182 ( .A1(n46631), .A2(n46637), .ZN(n44865) );
  INV_X1 U44183 ( .A(n44865), .ZN(n41136) );
  INV_X1 U44184 ( .A(n41134), .ZN(n41135) );
  AOI22_X1 U44185 ( .A1(n41138), .A2(n41137), .B1(n41136), .B2(n41135), .ZN(
        n41139) );
  INV_X1 U44186 ( .A(n44864), .ZN(n45760) );
  XNOR2_X1 U44187 ( .A(n46043), .B(n43014), .ZN(n42100) );
  OR2_X1 U44188 ( .A1(n41142), .A2(n41141), .ZN(n41154) );
  INV_X1 U44189 ( .A(n41146), .ZN(n41153) );
  XNOR2_X1 U44190 ( .A(n41156), .B(n41155), .ZN(n41157) );
  XNOR2_X1 U44191 ( .A(n51329), .B(n41157), .ZN(n41158) );
  XNOR2_X1 U44192 ( .A(n42100), .B(n41158), .ZN(n42430) );
  XNOR2_X1 U44193 ( .A(n41159), .B(n42430), .ZN(n41182) );
  XNOR2_X1 U44194 ( .A(n43655), .B(n51338), .ZN(n41160) );
  XNOR2_X1 U44195 ( .A(n41160), .B(n43657), .ZN(n41180) );
  INV_X1 U44196 ( .A(n4431), .ZN(n48775) );
  XNOR2_X1 U44197 ( .A(n41161), .B(n48775), .ZN(n41162) );
  XNOR2_X1 U44198 ( .A(n42938), .B(n41162), .ZN(n41178) );
  INV_X1 U44199 ( .A(n41163), .ZN(n41165) );
  NAND2_X1 U44200 ( .A1(n41165), .A2(n41164), .ZN(n41169) );
  NAND2_X1 U44201 ( .A1(n41166), .A2(n41692), .ZN(n41167) );
  NAND3_X1 U44202 ( .A1(n41169), .A2(n41168), .A3(n41167), .ZN(n41177) );
  NAND2_X1 U44203 ( .A1(n41692), .A2(n41706), .ZN(n41616) );
  OAI21_X1 U44204 ( .B1(n41170), .B2(n41616), .A(n41690), .ZN(n41173) );
  NAND2_X1 U44205 ( .A1(n41695), .A2(n2867), .ZN(n41171) );
  NAND4_X1 U44206 ( .A1(n41173), .A2(n41697), .A3(n41172), .A4(n41171), .ZN(
        n41176) );
  INV_X1 U44207 ( .A(n41174), .ZN(n41175) );
  XNOR2_X1 U44208 ( .A(n44937), .B(n4564), .ZN(n45100) );
  XNOR2_X1 U44209 ( .A(n41178), .B(n45100), .ZN(n41179) );
  XNOR2_X1 U44210 ( .A(n41180), .B(n41179), .ZN(n41181) );
  XNOR2_X1 U44211 ( .A(n41182), .B(n41181), .ZN(n41186) );
  XNOR2_X1 U44212 ( .A(n41183), .B(n4937), .ZN(n41184) );
  XNOR2_X1 U44213 ( .A(n516), .B(n41184), .ZN(n41185) );
  XNOR2_X1 U44214 ( .A(n43149), .B(n41185), .ZN(n43934) );
  XNOR2_X1 U44215 ( .A(n43168), .B(n43781), .ZN(n43392) );
  XNOR2_X1 U44216 ( .A(n41189), .B(n41188), .ZN(n41190) );
  XNOR2_X1 U44217 ( .A(n51464), .B(n41190), .ZN(n41191) );
  XNOR2_X1 U44218 ( .A(n43392), .B(n41191), .ZN(n42624) );
  XNOR2_X1 U44219 ( .A(n41192), .B(n42624), .ZN(n41253) );
  NAND3_X1 U44220 ( .A1(n41194), .A2(n41193), .A3(n51052), .ZN(n41199) );
  AND2_X1 U44221 ( .A1(n41212), .A2(n51052), .ZN(n41201) );
  NAND2_X1 U44222 ( .A1(n41201), .A2(n51430), .ZN(n41198) );
  INV_X1 U44223 ( .A(n41196), .ZN(n41197) );
  MUX2_X1 U44224 ( .A(n41199), .B(n41198), .S(n41197), .Z(n41222) );
  AND3_X1 U44225 ( .A1(n41204), .A2(n41205), .A3(n41203), .ZN(n41221) );
  OAI21_X1 U44226 ( .B1(n2408), .B2(n51052), .A(n41212), .ZN(n41218) );
  INV_X1 U44227 ( .A(n41209), .ZN(n41217) );
  OAI21_X1 U44228 ( .B1(n41212), .B2(n41211), .A(n41210), .ZN(n41214) );
  NOR2_X1 U44229 ( .A1(n41214), .A2(n41213), .ZN(n41216) );
  NAND4_X1 U44230 ( .A1(n41218), .A2(n41217), .A3(n41216), .A4(n41215), .ZN(
        n41219) );
  NAND4_X2 U44231 ( .A1(n41219), .A2(n41220), .A3(n41222), .A4(n41221), .ZN(
        n45293) );
  XOR2_X1 U44232 ( .A(n41567), .B(n41223), .Z(n41224) );
  XNOR2_X1 U44233 ( .A(n41225), .B(n41224), .ZN(n41226) );
  XNOR2_X1 U44234 ( .A(n43915), .B(n41226), .ZN(n41249) );
  NAND2_X1 U44235 ( .A1(n41229), .A2(n41228), .ZN(n41233) );
  INV_X1 U44236 ( .A(n41236), .ZN(n41230) );
  NAND2_X1 U44237 ( .A1(n41231), .A2(n41234), .ZN(n41232) );
  OAI22_X1 U44238 ( .A1(n41235), .A2(n39316), .B1(n41234), .B2(n41670), .ZN(
        n41240) );
  NAND3_X1 U44239 ( .A1(n41230), .A2(n41237), .A3(n41244), .ZN(n41239) );
  XNOR2_X1 U44240 ( .A(n41249), .B(n44923), .ZN(n41250) );
  XNOR2_X1 U44241 ( .A(n41251), .B(n41250), .ZN(n41252) );
  INV_X1 U44244 ( .A(n43218), .ZN(n41271) );
  OAI21_X1 U44246 ( .B1(n41258), .B2(n41734), .A(n41257), .ZN(n41631) );
  NOR2_X1 U44247 ( .A1(n41265), .A2(n41735), .ZN(n41259) );
  INV_X1 U44248 ( .A(n41728), .ZN(n41260) );
  NAND2_X1 U44249 ( .A1(n41261), .A2(n41260), .ZN(n41267) );
  NAND2_X1 U44250 ( .A1(n41731), .A2(n41263), .ZN(n41266) );
  NAND2_X1 U44251 ( .A1(n41269), .A2(n41268), .ZN(n41264) );
  NAND4_X1 U44252 ( .A1(n41267), .A2(n41266), .A3(n41265), .A4(n41264), .ZN(
        n41636) );
  OAI21_X1 U44253 ( .B1(n41631), .B2(n41632), .A(n41636), .ZN(n41270) );
  OAI21_X1 U44254 ( .B1(n41269), .B2(n41268), .A(n41729), .ZN(n41634) );
  NAND2_X1 U44255 ( .A1(n41270), .A2(n41634), .ZN(n45385) );
  XNOR2_X1 U44256 ( .A(n44288), .B(n45385), .ZN(n43831) );
  XNOR2_X1 U44257 ( .A(n41271), .B(n43831), .ZN(n41307) );
  XNOR2_X1 U44258 ( .A(n41629), .B(n41272), .ZN(n42663) );
  XNOR2_X1 U44259 ( .A(n2103), .B(n42663), .ZN(n41273) );
  XNOR2_X1 U44260 ( .A(n42222), .B(n41273), .ZN(n41306) );
  NOR2_X1 U44261 ( .A1(n41274), .A2(n8615), .ZN(n41279) );
  NAND2_X1 U44262 ( .A1(n52192), .A2(n41275), .ZN(n41281) );
  INV_X1 U44263 ( .A(n41281), .ZN(n41277) );
  AOI22_X1 U44264 ( .A1(n41279), .A2(n41278), .B1(n41277), .B2(n41276), .ZN(
        n41297) );
  XNOR2_X1 U44265 ( .A(n41281), .B(n8615), .ZN(n41290) );
  OAI21_X1 U44266 ( .B1(n52193), .B2(n41283), .A(n41282), .ZN(n41284) );
  INV_X1 U44267 ( .A(n41284), .ZN(n41289) );
  NAND3_X1 U44268 ( .A1(n41287), .A2(n41286), .A3(n41285), .ZN(n41288) );
  NAND3_X1 U44269 ( .A1(n41290), .A2(n41289), .A3(n41288), .ZN(n41296) );
  XNOR2_X1 U44270 ( .A(n44006), .B(n41298), .ZN(n43229) );
  XNOR2_X1 U44271 ( .A(n41300), .B(n41299), .ZN(n41301) );
  XNOR2_X1 U44272 ( .A(n43696), .B(n41301), .ZN(n41303) );
  XNOR2_X1 U44273 ( .A(n41303), .B(n41302), .ZN(n41304) );
  XNOR2_X1 U44274 ( .A(n43229), .B(n41304), .ZN(n41305) );
  XNOR2_X1 U44275 ( .A(n44525), .B(n45415), .ZN(n41309) );
  XNOR2_X1 U44276 ( .A(n43950), .B(n1354), .ZN(n41311) );
  XNOR2_X1 U44277 ( .A(n41311), .B(n2185), .ZN(n41312) );
  XNOR2_X1 U44278 ( .A(n2228), .B(n41312), .ZN(n45277) );
  XNOR2_X1 U44279 ( .A(n41314), .B(n41313), .ZN(n41315) );
  XNOR2_X1 U44280 ( .A(n51307), .B(n41315), .ZN(n41337) );
  NAND3_X1 U44281 ( .A1(n41318), .A2(n41317), .A3(n41316), .ZN(n41322) );
  OAI211_X1 U44282 ( .C1(n41320), .C2(n41332), .A(n41329), .B(n41319), .ZN(
        n41321) );
  OAI21_X1 U44283 ( .B1(n41333), .B2(n41332), .A(n41331), .ZN(n41334) );
  XNOR2_X1 U44284 ( .A(n44314), .B(n41337), .ZN(n41362) );
  INV_X1 U44285 ( .A(n41338), .ZN(n41341) );
  NAND4_X1 U44286 ( .A1(n41342), .A2(n41341), .A3(n38740), .A4(n41340), .ZN(
        n41361) );
  AND2_X1 U44287 ( .A1(n41355), .A2(n41352), .ZN(n41346) );
  AOI21_X1 U44288 ( .B1(n41349), .B2(n41352), .A(n41348), .ZN(n41351) );
  NAND2_X1 U44289 ( .A1(n41355), .A2(n41354), .ZN(n41357) );
  NAND2_X1 U44290 ( .A1(n41357), .A2(n52087), .ZN(n41359) );
  XNOR2_X1 U44291 ( .A(n44893), .B(n41362), .ZN(n41364) );
  XNOR2_X1 U44292 ( .A(n45279), .B(n43141), .ZN(n41363) );
  XNOR2_X1 U44293 ( .A(n41364), .B(n41363), .ZN(n41365) );
  XNOR2_X1 U44294 ( .A(n45467), .B(n41367), .ZN(n41368) );
  XNOR2_X1 U44295 ( .A(n41368), .B(n46143), .ZN(n42693) );
  XNOR2_X1 U44296 ( .A(n42693), .B(n43048), .ZN(n41371) );
  NAND3_X1 U44298 ( .A1(n41375), .A2(n3775), .A3(n41374), .ZN(n41376) );
  OAI211_X1 U44299 ( .C1(n41379), .C2(n41378), .A(n41377), .B(n41376), .ZN(
        n41381) );
  OAI21_X1 U44300 ( .B1(n41383), .B2(n41382), .A(n676), .ZN(n41384) );
  XNOR2_X1 U44301 ( .A(n41387), .B(n45355), .ZN(n41724) );
  OR2_X1 U44302 ( .A1(n41389), .A2(n41391), .ZN(n41398) );
  NAND2_X1 U44303 ( .A1(n41391), .A2(n41390), .ZN(n41392) );
  OAI211_X1 U44304 ( .C1(n41543), .C2(n41393), .A(n41392), .B(n8754), .ZN(
        n41397) );
  OAI211_X1 U44305 ( .C1(n41554), .C2(n52120), .A(n41544), .B(n7985), .ZN(
        n41396) );
  XNOR2_X1 U44306 ( .A(n4895), .B(n4923), .ZN(n41400) );
  XNOR2_X1 U44307 ( .A(n41401), .B(n41400), .ZN(n41402) );
  XNOR2_X1 U44308 ( .A(n41403), .B(n41402), .ZN(n41404) );
  XNOR2_X1 U44309 ( .A(n45089), .B(n41404), .ZN(n41405) );
  XNOR2_X1 U44310 ( .A(n41405), .B(n43363), .ZN(n41406) );
  XNOR2_X1 U44311 ( .A(n41724), .B(n41406), .ZN(n41407) );
  XNOR2_X2 U44312 ( .A(n41409), .B(n41408), .ZN(n46591) );
  INV_X1 U44313 ( .A(n46591), .ZN(n46709) );
  INV_X1 U44314 ( .A(n46596), .ZN(n41410) );
  INV_X1 U44315 ( .A(n46597), .ZN(n46572) );
  NAND2_X1 U44316 ( .A1(n46584), .A2(n46572), .ZN(n41469) );
  XNOR2_X1 U44317 ( .A(n43584), .B(n4733), .ZN(n41889) );
  NAND2_X1 U44318 ( .A1(n42007), .A2(n42006), .ZN(n41411) );
  NOR2_X1 U44319 ( .A1(n6236), .A2(n41997), .ZN(n42021) );
  AND2_X1 U44320 ( .A1(n41587), .A2(n41581), .ZN(n41577) );
  INV_X1 U44321 ( .A(n42014), .ZN(n41413) );
  NAND3_X1 U44322 ( .A1(n41414), .A2(n41413), .A3(n42010), .ZN(n41422) );
  NAND2_X1 U44323 ( .A1(n41416), .A2(n4943), .ZN(n41419) );
  INV_X1 U44324 ( .A(n41503), .ZN(n41418) );
  NAND4_X1 U44325 ( .A1(n41420), .A2(n41419), .A3(n41418), .A4(n41417), .ZN(
        n41421) );
  XOR2_X1 U44327 ( .A(n44963), .B(n51294), .Z(n41424) );
  XNOR2_X1 U44328 ( .A(n41889), .B(n41424), .ZN(n41425) );
  XNOR2_X1 U44329 ( .A(n41425), .B(n44478), .ZN(n41428) );
  XNOR2_X1 U44330 ( .A(n45067), .B(n41426), .ZN(n41427) );
  XNOR2_X1 U44331 ( .A(n43318), .B(n51461), .ZN(n43070) );
  XNOR2_X1 U44332 ( .A(n43070), .B(n41427), .ZN(n42680) );
  XNOR2_X1 U44333 ( .A(n42680), .B(n41428), .ZN(n41468) );
  AOI21_X1 U44334 ( .B1(n41430), .B2(n41440), .A(n41429), .ZN(n41431) );
  NOR2_X1 U44335 ( .A1(n41432), .A2(n41431), .ZN(n41456) );
  NOR2_X1 U44336 ( .A1(n41433), .A2(n41436), .ZN(n41439) );
  INV_X1 U44337 ( .A(n41434), .ZN(n41438) );
  NOR2_X1 U44338 ( .A1(n41442), .A2(n41435), .ZN(n41437) );
  AOI22_X1 U44339 ( .A1(n41439), .A2(n41438), .B1(n41437), .B2(n41436), .ZN(
        n41445) );
  INV_X1 U44340 ( .A(n41440), .ZN(n41443) );
  OAI21_X1 U44341 ( .B1(n41443), .B2(n41442), .A(n41441), .ZN(n41444) );
  AND2_X1 U44342 ( .A1(n41445), .A2(n41444), .ZN(n41455) );
  NOR2_X1 U44343 ( .A1(n41447), .A2(n41446), .ZN(n41449) );
  AOI22_X1 U44344 ( .A1(n41451), .A2(n41450), .B1(n41449), .B2(n41448), .ZN(
        n41454) );
  NAND2_X1 U44345 ( .A1(n41452), .A2(n2248), .ZN(n41453) );
  XNOR2_X1 U44346 ( .A(n42980), .B(n44164), .ZN(n41457) );
  XNOR2_X1 U44347 ( .A(n41457), .B(n43889), .ZN(n41458) );
  XNOR2_X1 U44348 ( .A(n4676), .B(n4237), .ZN(n41459) );
  XNOR2_X1 U44349 ( .A(n41460), .B(n41459), .ZN(n41461) );
  XNOR2_X1 U44350 ( .A(n41462), .B(n41461), .ZN(n41463) );
  XNOR2_X1 U44351 ( .A(n42500), .B(n41463), .ZN(n41464) );
  INV_X1 U44352 ( .A(Key[40]), .ZN(n48064) );
  XNOR2_X1 U44353 ( .A(n41465), .B(n42504), .ZN(n41466) );
  XNOR2_X1 U44354 ( .A(n41759), .B(n41466), .ZN(n41467) );
  AOI22_X1 U44355 ( .A1(n44845), .A2(n46707), .B1(n46584), .B2(n46574), .ZN(
        n41476) );
  INV_X1 U44356 ( .A(n46575), .ZN(n41475) );
  INV_X1 U44357 ( .A(n46580), .ZN(n41471) );
  INV_X1 U44358 ( .A(n41470), .ZN(n46595) );
  AOI22_X1 U44359 ( .A1(n41471), .A2(n46595), .B1(n46705), .B2(n405), .ZN(
        n41474) );
  AND2_X1 U44360 ( .A1(n46589), .A2(n46709), .ZN(n44704) );
  INV_X1 U44361 ( .A(n44704), .ZN(n41472) );
  OAI211_X1 U44362 ( .C1(n46584), .C2(n51396), .A(n46701), .B(n41472), .ZN(
        n41473) );
  OAI211_X1 U44363 ( .C1(n41476), .C2(n41475), .A(n41474), .B(n41473), .ZN(
        n41477) );
  XNOR2_X1 U44364 ( .A(n45116), .B(n41479), .ZN(n44050) );
  XNOR2_X1 U44365 ( .A(n52043), .B(n44050), .ZN(n41495) );
  NAND3_X1 U44366 ( .A1(n41482), .A2(n41481), .A3(n41480), .ZN(n41484) );
  OAI21_X1 U44367 ( .B1(n41485), .B2(n41484), .A(n41483), .ZN(n41486) );
  INV_X1 U44368 ( .A(n41486), .ZN(n41493) );
  NAND3_X1 U44370 ( .A1(n42048), .A2(n52128), .A3(n596), .ZN(n41490) );
  INV_X1 U44371 ( .A(n43206), .ZN(n41494) );
  XNOR2_X1 U44372 ( .A(n43655), .B(n43929), .ZN(n44038) );
  XNOR2_X1 U44373 ( .A(n44038), .B(n41495), .ZN(n41521) );
  XNOR2_X1 U44374 ( .A(n41497), .B(n41496), .ZN(n41498) );
  XNOR2_X1 U44375 ( .A(n41499), .B(n41498), .ZN(n41500) );
  XNOR2_X1 U44376 ( .A(n51338), .B(n41500), .ZN(n41501) );
  XNOR2_X1 U44377 ( .A(n41501), .B(n672), .ZN(n41519) );
  OAI21_X1 U44378 ( .B1(n41504), .B2(n41503), .A(n41502), .ZN(n41505) );
  INV_X1 U44379 ( .A(n41505), .ZN(n41517) );
  NAND2_X1 U44380 ( .A1(n41997), .A2(n4943), .ZN(n41507) );
  OR2_X1 U44381 ( .A1(n41507), .A2(n41506), .ZN(n41586) );
  AND2_X1 U44382 ( .A1(n41508), .A2(n41586), .ZN(n41516) );
  OAI21_X1 U44383 ( .B1(n42002), .B2(n41510), .A(n41509), .ZN(n41515) );
  NAND2_X1 U44384 ( .A1(n41513), .A2(n41512), .ZN(n41514) );
  XNOR2_X1 U44385 ( .A(n45099), .B(n52171), .ZN(n44565) );
  XNOR2_X1 U44386 ( .A(n44565), .B(n41519), .ZN(n41520) );
  XNOR2_X1 U44387 ( .A(n41520), .B(n41521), .ZN(n41523) );
  XNOR2_X1 U44388 ( .A(n42819), .B(n45303), .ZN(n43160) );
  XNOR2_X1 U44389 ( .A(n45454), .B(n43160), .ZN(n41522) );
  XNOR2_X1 U44390 ( .A(n43781), .B(n1326), .ZN(n41561) );
  OR2_X1 U44391 ( .A1(n41534), .A2(n41530), .ZN(n41528) );
  NAND2_X1 U44392 ( .A1(n41540), .A2(n41524), .ZN(n41545) );
  OAI211_X1 U44393 ( .C1(n41526), .C2(n41525), .A(n41534), .B(n41540), .ZN(
        n41527) );
  OAI21_X1 U44394 ( .B1(n41528), .B2(n41545), .A(n41527), .ZN(n41529) );
  INV_X1 U44395 ( .A(n41529), .ZN(n41560) );
  INV_X1 U44396 ( .A(n41530), .ZN(n41532) );
  AOI22_X1 U44397 ( .A1(n41533), .A2(n41532), .B1(n41531), .B2(n41554), .ZN(
        n41559) );
  NAND2_X1 U44398 ( .A1(n41539), .A2(n41535), .ZN(n41536) );
  NOR2_X1 U44399 ( .A1(n41540), .A2(n41536), .ZN(n41538) );
  AOI21_X1 U44400 ( .B1(n3559), .B2(n41538), .A(n41537), .ZN(n41550) );
  NOR2_X1 U44402 ( .A1(n41544), .A2(n41553), .ZN(n41547) );
  INV_X1 U44403 ( .A(n41545), .ZN(n41546) );
  NAND2_X1 U44404 ( .A1(n41547), .A2(n41546), .ZN(n41548) );
  INV_X1 U44406 ( .A(n41551), .ZN(n41552) );
  NOR2_X1 U44407 ( .A1(n41553), .A2(n41552), .ZN(n41555) );
  XNOR2_X1 U44408 ( .A(n41561), .B(n44547), .ZN(n43062) );
  XNOR2_X1 U44409 ( .A(n43909), .B(n44534), .ZN(n43802) );
  XNOR2_X1 U44410 ( .A(n41563), .B(n41562), .ZN(n41564) );
  XNOR2_X1 U44411 ( .A(n43915), .B(n41564), .ZN(n41565) );
  XNOR2_X1 U44412 ( .A(n43802), .B(n41565), .ZN(n41566) );
  XNOR2_X1 U44413 ( .A(n43062), .B(n41566), .ZN(n41571) );
  INV_X1 U44414 ( .A(n41567), .ZN(n41568) );
  XNOR2_X1 U44415 ( .A(n42284), .B(n41568), .ZN(n41569) );
  XNOR2_X1 U44416 ( .A(n44923), .B(n45285), .ZN(n44546) );
  XNOR2_X1 U44417 ( .A(n41570), .B(n44546), .ZN(n41823) );
  XNOR2_X1 U44418 ( .A(n41823), .B(n41571), .ZN(n41595) );
  NAND2_X1 U44419 ( .A1(n41587), .A2(n42020), .ZN(n42001) );
  INV_X1 U44420 ( .A(n42001), .ZN(n41572) );
  NAND4_X1 U44421 ( .A1(n41573), .A2(n41588), .A3(n41572), .A4(n42015), .ZN(
        n41574) );
  INV_X1 U44422 ( .A(n42000), .ZN(n41579) );
  INV_X1 U44423 ( .A(n41576), .ZN(n41578) );
  NOR2_X1 U44424 ( .A1(n41581), .A2(n42020), .ZN(n41582) );
  XNOR2_X1 U44425 ( .A(n52130), .B(n43197), .ZN(n41593) );
  XNOR2_X1 U44426 ( .A(n44056), .B(n41593), .ZN(n41594) );
  NOR2_X1 U44428 ( .A1(n46730), .A2(n51488), .ZN(n46737) );
  INV_X1 U44429 ( .A(n46737), .ZN(n45810) );
  XNOR2_X1 U44430 ( .A(n43973), .B(n42863), .ZN(n41596) );
  XNOR2_X1 U44431 ( .A(n41596), .B(n44301), .ZN(n43006) );
  XNOR2_X1 U44432 ( .A(n41597), .B(n2183), .ZN(n42069) );
  XNOR2_X1 U44433 ( .A(n42069), .B(n41598), .ZN(n41599) );
  XNOR2_X1 U44434 ( .A(n44016), .B(n41599), .ZN(n41600) );
  XNOR2_X1 U44435 ( .A(n44209), .B(n41600), .ZN(n41601) );
  XNOR2_X1 U44436 ( .A(n43229), .B(n41601), .ZN(n41602) );
  INV_X1 U44437 ( .A(n41603), .ZN(n41605) );
  OAI21_X1 U44438 ( .B1(n41606), .B2(n41605), .A(n41604), .ZN(n41608) );
  NAND2_X1 U44439 ( .A1(n41608), .A2(n41607), .ZN(n44300) );
  NOR2_X1 U44440 ( .A1(n41702), .A2(n2867), .ZN(n41687) );
  AOI22_X1 U44441 ( .A1(n41612), .A2(n41611), .B1(n41687), .B2(n41610), .ZN(
        n41628) );
  NAND2_X1 U44442 ( .A1(n41693), .A2(n41706), .ZN(n41620) );
  OAI22_X1 U44443 ( .A1(n41613), .A2(n41620), .B1(n41703), .B2(n41698), .ZN(
        n41614) );
  INV_X1 U44444 ( .A(n41614), .ZN(n41627) );
  NAND2_X1 U44445 ( .A1(n41618), .A2(n41697), .ZN(n41626) );
  NAND3_X1 U44446 ( .A1(n41688), .A2(n41706), .A3(n41691), .ZN(n41619) );
  NAND3_X1 U44447 ( .A1(n41695), .A2(n41621), .A3(n41706), .ZN(n41622) );
  NAND2_X1 U44448 ( .A1(n41702), .A2(n41622), .ZN(n41623) );
  NAND2_X1 U44449 ( .A1(n41624), .A2(n41623), .ZN(n41625) );
  XNOR2_X1 U44450 ( .A(n42869), .B(n41630), .ZN(n44516) );
  INV_X1 U44451 ( .A(n41631), .ZN(n41635) );
  INV_X1 U44452 ( .A(n41632), .ZN(n41633) );
  XNOR2_X1 U44453 ( .A(n44901), .B(n51408), .ZN(n41656) );
  NOR2_X1 U44454 ( .A1(n41647), .A2(n41646), .ZN(n41639) );
  AND2_X1 U44455 ( .A1(n41985), .A2(n41646), .ZN(n41637) );
  AOI22_X1 U44456 ( .A1(n41640), .A2(n41639), .B1(n41638), .B2(n41637), .ZN(
        n41654) );
  NOR2_X1 U44457 ( .A1(n41645), .A2(n41985), .ZN(n41651) );
  AND3_X1 U44458 ( .A1(n41647), .A2(n41975), .A3(n41646), .ZN(n41648) );
  AOI21_X1 U44459 ( .B1(n41651), .B2(n41649), .A(n41648), .ZN(n41653) );
  OAI21_X1 U44460 ( .B1(n41651), .B2(n41650), .A(n41986), .ZN(n41652) );
  INV_X1 U44461 ( .A(n44510), .ZN(n41655) );
  XNOR2_X1 U44462 ( .A(n42450), .B(n42339), .ZN(n46100) );
  XNOR2_X1 U44463 ( .A(n7101), .B(n46100), .ZN(n41657) );
  XNOR2_X1 U44464 ( .A(n46109), .B(n41657), .ZN(n41856) );
  INV_X1 U44465 ( .A(n41856), .ZN(n41658) );
  XNOR2_X1 U44466 ( .A(n41658), .B(n41659), .ZN(n41723) );
  XOR2_X1 U44467 ( .A(n46118), .B(n44320), .Z(n41722) );
  XNOR2_X1 U44468 ( .A(n51099), .B(n51100), .ZN(n41666) );
  XNOR2_X1 U44469 ( .A(n41661), .B(n41660), .ZN(n41662) );
  XNOR2_X1 U44470 ( .A(n41663), .B(n41662), .ZN(n41664) );
  XNOR2_X1 U44471 ( .A(n46128), .B(n41664), .ZN(n41665) );
  XNOR2_X1 U44472 ( .A(n41666), .B(n41665), .ZN(n41667) );
  XNOR2_X1 U44473 ( .A(n41667), .B(n43141), .ZN(n41720) );
  AND2_X1 U44474 ( .A1(n41680), .A2(n41670), .ZN(n41668) );
  NOR2_X1 U44475 ( .A1(n6335), .A2(n41670), .ZN(n41672) );
  NOR2_X1 U44476 ( .A1(n41673), .A2(n41672), .ZN(n41678) );
  NOR2_X1 U44477 ( .A1(n52198), .A2(n41679), .ZN(n41676) );
  XNOR2_X1 U44478 ( .A(n43619), .B(n45050), .ZN(n41686) );
  XNOR2_X1 U44479 ( .A(n43027), .B(n41686), .ZN(n43721) );
  NAND3_X1 U44480 ( .A1(n41689), .A2(n41688), .A3(n41687), .ZN(n41716) );
  NAND3_X1 U44481 ( .A1(n41693), .A2(n41692), .A3(n41691), .ZN(n41694) );
  OAI21_X1 U44482 ( .B1(n41699), .B2(n41698), .A(n41697), .ZN(n41700) );
  NAND4_X1 U44483 ( .A1(n41705), .A2(n41704), .A3(n2179), .A4(n41702), .ZN(
        n41714) );
  NAND2_X1 U44484 ( .A1(n41707), .A2(n41706), .ZN(n41712) );
  NAND2_X1 U44485 ( .A1(n41709), .A2(n41708), .ZN(n41710) );
  AND3_X1 U44486 ( .A1(n41712), .A2(n41711), .A3(n41710), .ZN(n41713) );
  XNOR2_X1 U44487 ( .A(n51101), .B(n46113), .ZN(n41718) );
  INV_X1 U44488 ( .A(n44879), .ZN(n41717) );
  XNOR2_X1 U44489 ( .A(n41718), .B(n41717), .ZN(n42352) );
  XNOR2_X1 U44490 ( .A(n43721), .B(n42352), .ZN(n41719) );
  XNOR2_X1 U44491 ( .A(n41719), .B(n41720), .ZN(n41721) );
  XNOR2_X1 U44493 ( .A(n41724), .B(n569), .ZN(n43258) );
  XNOR2_X1 U44494 ( .A(n44501), .B(n43943), .ZN(n43815) );
  AOI22_X1 U44495 ( .A1(n41729), .A2(n41728), .B1(n41727), .B2(n41726), .ZN(
        n41739) );
  INV_X1 U44496 ( .A(n41730), .ZN(n41732) );
  NAND3_X1 U44497 ( .A1(n41734), .A2(n41735), .A3(n39593), .ZN(n41738) );
  XNOR2_X1 U44498 ( .A(n43815), .B(n43725), .ZN(n41745) );
  XNOR2_X1 U44499 ( .A(n41740), .B(n2203), .ZN(n41741) );
  XNOR2_X1 U44500 ( .A(n41742), .B(n41741), .ZN(n41743) );
  XNOR2_X1 U44501 ( .A(n41745), .B(n41744), .ZN(n41746) );
  XNOR2_X1 U44502 ( .A(n43258), .B(n41746), .ZN(n41757) );
  NAND2_X1 U44503 ( .A1(n42149), .A2(n42136), .ZN(n42750) );
  NAND2_X1 U44504 ( .A1(n41748), .A2(n41747), .ZN(n41750) );
  OAI21_X1 U44505 ( .B1(n42144), .B2(n42145), .A(n51375), .ZN(n41749) );
  NAND2_X1 U44506 ( .A1(n41750), .A2(n41749), .ZN(n42753) );
  INV_X1 U44507 ( .A(n42753), .ZN(n41753) );
  OAI21_X1 U44508 ( .B1(n42154), .B2(n42157), .A(n41770), .ZN(n41752) );
  INV_X1 U44509 ( .A(n42155), .ZN(n41774) );
  OAI21_X1 U44510 ( .B1(n41752), .B2(n41774), .A(n41751), .ZN(n42751) );
  OAI211_X1 U44511 ( .C1(n42749), .C2(n42750), .A(n41753), .B(n42751), .ZN(
        n41754) );
  XNOR2_X1 U44512 ( .A(n41755), .B(n43819), .ZN(n44096) );
  XNOR2_X1 U44513 ( .A(n44096), .B(n41882), .ZN(n41756) );
  XNOR2_X1 U44515 ( .A(n42316), .B(n43584), .ZN(n43313) );
  XNOR2_X1 U44516 ( .A(n45490), .B(n43313), .ZN(n44479) );
  AND2_X1 U44517 ( .A1(n42154), .A2(n41764), .ZN(n41761) );
  AOI21_X1 U44518 ( .B1(n41761), .B2(n41760), .A(n42138), .ZN(n41769) );
  NAND2_X1 U44519 ( .A1(n41769), .A2(n41762), .ZN(n41768) );
  NOR2_X1 U44520 ( .A1(n687), .A2(n42154), .ZN(n41763) );
  OAI211_X1 U44521 ( .C1(n41763), .C2(n42153), .A(n52092), .B(n51375), .ZN(
        n41767) );
  AND2_X1 U44522 ( .A1(n41764), .A2(n41770), .ZN(n42139) );
  NAND2_X1 U44523 ( .A1(n42139), .A2(n687), .ZN(n41765) );
  NAND4_X1 U44524 ( .A1(n41768), .A2(n41767), .A3(n41766), .A4(n41765), .ZN(
        n41779) );
  INV_X1 U44525 ( .A(n41769), .ZN(n41777) );
  AND2_X1 U44526 ( .A1(n42154), .A2(n42157), .ZN(n41772) );
  AND2_X1 U44527 ( .A1(n41770), .A2(n42131), .ZN(n41771) );
  OAI21_X1 U44528 ( .B1(n41772), .B2(n52092), .A(n41771), .ZN(n41776) );
  NAND3_X1 U44529 ( .A1(n41774), .A2(n42138), .A3(n41773), .ZN(n41775) );
  OAI211_X1 U44530 ( .C1(n41777), .C2(n42142), .A(n41776), .B(n41775), .ZN(
        n41778) );
  XNOR2_X1 U44531 ( .A(n43496), .B(n4585), .ZN(n45076) );
  XNOR2_X1 U44532 ( .A(n42889), .B(Key[40]), .ZN(n41780) );
  XNOR2_X1 U44533 ( .A(n44954), .B(n41780), .ZN(n41781) );
  XNOR2_X1 U44534 ( .A(n41782), .B(n41781), .ZN(n41783) );
  XNOR2_X1 U44535 ( .A(n43102), .B(n41783), .ZN(n41784) );
  XNOR2_X1 U44536 ( .A(n45076), .B(n41784), .ZN(n41786) );
  XNOR2_X1 U44537 ( .A(n41956), .B(n44962), .ZN(n41785) );
  XNOR2_X1 U44538 ( .A(n41786), .B(n41785), .ZN(n41787) );
  INV_X1 U44539 ( .A(n41788), .ZN(n41790) );
  INV_X1 U44540 ( .A(n41794), .ZN(n41795) );
  NOR3_X1 U44541 ( .A1(n41797), .A2(n51684), .A3(n41796), .ZN(n41798) );
  NAND2_X1 U44542 ( .A1(n41799), .A2(n41798), .ZN(n41806) );
  NOR2_X1 U44543 ( .A1(n41801), .A2(n51684), .ZN(n41803) );
  OAI21_X1 U44544 ( .B1(n41804), .B2(n41803), .A(n41802), .ZN(n41805) );
  XNOR2_X1 U44545 ( .A(n43344), .B(n44963), .ZN(n41809) );
  XNOR2_X1 U44546 ( .A(n52103), .B(n41809), .ZN(n41810) );
  XNOR2_X1 U44547 ( .A(n41810), .B(n42504), .ZN(n44085) );
  NAND2_X1 U44548 ( .A1(n50965), .A2(n51344), .ZN(n46731) );
  AND2_X1 U44549 ( .A1(n41723), .A2(n46746), .ZN(n46739) );
  INV_X1 U44550 ( .A(n45804), .ZN(n44850) );
  NAND2_X1 U44551 ( .A1(n45186), .A2(n44850), .ZN(n45184) );
  INV_X1 U44552 ( .A(n45184), .ZN(n41811) );
  INV_X1 U44553 ( .A(n46731), .ZN(n45800) );
  AND2_X1 U44554 ( .A1(n46753), .A2(n51488), .ZN(n45799) );
  NAND2_X1 U44555 ( .A1(n45799), .A2(n46747), .ZN(n41812) );
  AND2_X1 U44556 ( .A1(n46746), .A2(n45190), .ZN(n41815) );
  NOR2_X1 U44557 ( .A1(n2092), .A2(n45188), .ZN(n41814) );
  AOI22_X1 U44558 ( .A1(n41815), .A2(n46737), .B1(n46743), .B2(n41814), .ZN(
        n41816) );
  INV_X1 U44559 ( .A(n47857), .ZN(n47879) );
  NAND2_X1 U44560 ( .A1(n47879), .A2(n51285), .ZN(n47876) );
  XNOR2_X1 U44561 ( .A(n43170), .B(n43781), .ZN(n41819) );
  BUF_X2 U44562 ( .A(n41820), .Z(n44542) );
  XNOR2_X1 U44563 ( .A(n44061), .B(n44542), .ZN(n41821) );
  XNOR2_X1 U44564 ( .A(n45426), .B(n75), .ZN(n41822) );
  XNOR2_X1 U44565 ( .A(n41822), .B(n45284), .ZN(n42129) );
  XNOR2_X1 U44566 ( .A(n42122), .B(n51444), .ZN(n42280) );
  INV_X1 U44569 ( .A(n45551), .ZN(n48206) );
  XNOR2_X1 U44570 ( .A(n43155), .B(n42938), .ZN(n41834) );
  XNOR2_X1 U44571 ( .A(n41825), .B(n4579), .ZN(n41826) );
  XNOR2_X1 U44572 ( .A(n41827), .B(n41826), .ZN(n41829) );
  XNOR2_X1 U44573 ( .A(n41829), .B(n41828), .ZN(n41830) );
  XNOR2_X1 U44574 ( .A(n41831), .B(n41830), .ZN(n41832) );
  XNOR2_X1 U44575 ( .A(n45114), .B(n41832), .ZN(n41833) );
  XNOR2_X1 U44576 ( .A(n41834), .B(n41833), .ZN(n41837) );
  XNOR2_X1 U44577 ( .A(n43014), .B(n41835), .ZN(n41836) );
  XNOR2_X1 U44578 ( .A(n41836), .B(n52171), .ZN(n45317) );
  XNOR2_X1 U44579 ( .A(n41837), .B(n45317), .ZN(n41838) );
  XNOR2_X1 U44580 ( .A(n42098), .B(n41838), .ZN(n41842) );
  XNOR2_X1 U44581 ( .A(n2206), .B(n43929), .ZN(n42377) );
  XNOR2_X1 U44582 ( .A(n44353), .B(n51329), .ZN(n41839) );
  XNOR2_X1 U44583 ( .A(n41839), .B(n51097), .ZN(n41840) );
  XNOR2_X1 U44584 ( .A(n42377), .B(n41840), .ZN(n41841) );
  XNOR2_X1 U44586 ( .A(n41844), .B(n41843), .ZN(n41845) );
  XNOR2_X1 U44587 ( .A(n42907), .B(n41845), .ZN(n41846) );
  XNOR2_X1 U44588 ( .A(n44301), .B(n41846), .ZN(n41847) );
  XNOR2_X1 U44589 ( .A(n42067), .B(n41847), .ZN(n41849) );
  XNOR2_X1 U44590 ( .A(n44006), .B(n44911), .ZN(n45394) );
  XNOR2_X1 U44591 ( .A(n45394), .B(n43291), .ZN(n41848) );
  XNOR2_X1 U44592 ( .A(n41848), .B(n41849), .ZN(n41855) );
  XNOR2_X1 U44593 ( .A(n41850), .B(n44900), .ZN(n41851) );
  XNOR2_X1 U44594 ( .A(n44016), .B(n41852), .ZN(n41853) );
  XNOR2_X1 U44595 ( .A(n43123), .B(n41853), .ZN(n44302) );
  XNOR2_X1 U44596 ( .A(n42218), .B(n44302), .ZN(n41854) );
  XNOR2_X1 U44597 ( .A(n41855), .B(n41854), .ZN(n41857) );
  INV_X1 U44599 ( .A(n48201), .ZN(n44996) );
  XNOR2_X1 U44600 ( .A(n41859), .B(n52096), .ZN(n44229) );
  XNOR2_X1 U44601 ( .A(n41860), .B(n44229), .ZN(n41863) );
  XNOR2_X1 U44602 ( .A(n44314), .B(n46113), .ZN(n41861) );
  XNOR2_X1 U44603 ( .A(n41861), .B(n44240), .ZN(n41862) );
  XNOR2_X1 U44604 ( .A(n44893), .B(n41862), .ZN(n45413) );
  XNOR2_X1 U44605 ( .A(n41863), .B(n45413), .ZN(n41871) );
  XNOR2_X1 U44606 ( .A(n44027), .B(n46128), .ZN(n44308) );
  XNOR2_X1 U44607 ( .A(n41865), .B(n41864), .ZN(n41866) );
  XNOR2_X1 U44608 ( .A(n42643), .B(n41866), .ZN(n41867) );
  INV_X1 U44609 ( .A(n42850), .ZN(n42923) );
  XNOR2_X1 U44610 ( .A(n41867), .B(n42923), .ZN(n41868) );
  XNOR2_X1 U44611 ( .A(n44308), .B(n41868), .ZN(n41869) );
  XNOR2_X1 U44612 ( .A(n44230), .B(n41869), .ZN(n41870) );
  NAND2_X1 U44613 ( .A1(n45539), .A2(n48210), .ZN(n41884) );
  XNOR2_X1 U44614 ( .A(n41873), .B(n41872), .ZN(n41874) );
  XNOR2_X1 U44615 ( .A(n43254), .B(n41874), .ZN(n41876) );
  XNOR2_X1 U44616 ( .A(n41876), .B(n43113), .ZN(n41877) );
  XNOR2_X1 U44617 ( .A(n41877), .B(n43048), .ZN(n41879) );
  XNOR2_X1 U44618 ( .A(n46150), .B(n41968), .ZN(n44372) );
  XNOR2_X1 U44619 ( .A(n43819), .B(n44372), .ZN(n41878) );
  XNOR2_X1 U44620 ( .A(n50967), .B(n43609), .ZN(n41880) );
  XNOR2_X1 U44621 ( .A(n41880), .B(n45355), .ZN(n44973) );
  XNOR2_X1 U44622 ( .A(n41966), .B(n44973), .ZN(n41881) );
  NOR2_X1 U44624 ( .A1(n48208), .A2(n45538), .ZN(n44270) );
  XNOR2_X1 U44625 ( .A(n41886), .B(n41885), .ZN(n41887) );
  XNOR2_X1 U44626 ( .A(n42980), .B(n41887), .ZN(n41888) );
  XNOR2_X1 U44627 ( .A(n41889), .B(n44964), .ZN(n41891) );
  XNOR2_X1 U44628 ( .A(n46081), .B(n44394), .ZN(n41890) );
  XNOR2_X1 U44629 ( .A(n41890), .B(n41891), .ZN(n41892) );
  XNOR2_X1 U44630 ( .A(n41892), .B(n41893), .ZN(n41907) );
  XNOR2_X1 U44631 ( .A(n41956), .B(n42500), .ZN(n45326) );
  XNOR2_X1 U44632 ( .A(n45326), .B(n42504), .ZN(n41906) );
  NOR2_X1 U44633 ( .A1(n41895), .A2(n41894), .ZN(n41896) );
  AND2_X1 U44634 ( .A1(n41897), .A2(n41896), .ZN(n41905) );
  INV_X1 U44635 ( .A(n41898), .ZN(n41899) );
  AOI21_X1 U44636 ( .B1(n41901), .B2(n41900), .A(n41899), .ZN(n41903) );
  MUX2_X1 U44637 ( .A(n41903), .B(n2379), .S(n41902), .Z(n41904) );
  NAND2_X1 U44638 ( .A1(n41905), .A2(n41904), .ZN(n44391) );
  XNOR2_X1 U44639 ( .A(n45490), .B(n44391), .ZN(n46082) );
  NAND2_X1 U44640 ( .A1(n44990), .A2(n52070), .ZN(n41909) );
  OAI211_X1 U44641 ( .C1(n45545), .C2(n48200), .A(n48205), .B(n41909), .ZN(
        n41910) );
  INV_X1 U44642 ( .A(n41910), .ZN(n41911) );
  NOR2_X1 U44643 ( .A1(n45540), .A2(n44992), .ZN(n48207) );
  INV_X1 U44645 ( .A(n44263), .ZN(n41921) );
  NAND3_X1 U44646 ( .A1(n48207), .A2(n52050), .A3(n41921), .ZN(n41917) );
  NAND2_X1 U44647 ( .A1(n44263), .A2(n44990), .ZN(n41914) );
  NAND2_X1 U44648 ( .A1(n45540), .A2(n48200), .ZN(n41913) );
  NAND3_X1 U44649 ( .A1(n41914), .A2(n41913), .A3(n48205), .ZN(n41915) );
  INV_X1 U44650 ( .A(n44992), .ZN(n44693) );
  NAND2_X1 U44652 ( .A1(n41915), .A2(n48214), .ZN(n41916) );
  AND2_X1 U44653 ( .A1(n45542), .A2(n52050), .ZN(n44269) );
  NAND2_X1 U44654 ( .A1(n48200), .A2(n48213), .ZN(n48204) );
  INV_X1 U44655 ( .A(n45539), .ZN(n41920) );
  NAND2_X1 U44656 ( .A1(n48205), .A2(n48200), .ZN(n41918) );
  NOR2_X1 U44657 ( .A1(n2119), .A2(n41918), .ZN(n41919) );
  INV_X1 U44658 ( .A(n45540), .ZN(n44696) );
  OAI21_X1 U44659 ( .B1(n44696), .B2(n52161), .A(n48208), .ZN(n41922) );
  AND2_X1 U44660 ( .A1(n41921), .A2(n44990), .ZN(n48221) );
  NAND2_X1 U44661 ( .A1(n41922), .A2(n48221), .ZN(n41923) );
  OR2_X1 U44662 ( .A1(n47876), .A2(n51470), .ZN(n47849) );
  XNOR2_X1 U44663 ( .A(n43496), .B(n42500), .ZN(n42289) );
  XNOR2_X1 U44664 ( .A(n42289), .B(n43313), .ZN(n43068) );
  NAND2_X1 U44665 ( .A1(n41929), .A2(n41928), .ZN(n41937) );
  OAI21_X1 U44666 ( .B1(n41931), .B2(n41930), .A(n42201), .ZN(n41936) );
  XNOR2_X1 U44668 ( .A(n41946), .B(n43596), .ZN(n41947) );
  XNOR2_X1 U44669 ( .A(n43068), .B(n41947), .ZN(n44969) );
  XNOR2_X1 U44670 ( .A(n41948), .B(n43764), .ZN(n41950) );
  XNOR2_X1 U44671 ( .A(n41950), .B(n41949), .ZN(n41951) );
  XNOR2_X1 U44672 ( .A(n45339), .B(n41951), .ZN(n41952) );
  XNOR2_X1 U44673 ( .A(n41952), .B(n44154), .ZN(n41953) );
  XNOR2_X1 U44674 ( .A(n41954), .B(n41953), .ZN(n41955) );
  XNOR2_X1 U44675 ( .A(n44969), .B(n41955), .ZN(n41959) );
  XNOR2_X1 U44676 ( .A(n42492), .B(n41956), .ZN(n44152) );
  XNOR2_X1 U44677 ( .A(n43349), .B(n44152), .ZN(n41957) );
  XNOR2_X1 U44678 ( .A(n44394), .B(n43889), .ZN(n44489) );
  XNOR2_X1 U44679 ( .A(n44489), .B(n41957), .ZN(n41958) );
  XNOR2_X1 U44680 ( .A(n41959), .B(n41958), .ZN(n42181) );
  XNOR2_X1 U44681 ( .A(n41961), .B(n41960), .ZN(n41962) );
  XNOR2_X1 U44682 ( .A(n43254), .B(n41962), .ZN(n41963) );
  XNOR2_X1 U44683 ( .A(n51398), .B(n44370), .ZN(n41964) );
  XNOR2_X1 U44684 ( .A(n41967), .B(n41966), .ZN(n41970) );
  XNOR2_X1 U44685 ( .A(n43724), .B(n41968), .ZN(n41969) );
  XNOR2_X1 U44686 ( .A(n41970), .B(n43936), .ZN(n41995) );
  INV_X1 U44687 ( .A(n41971), .ZN(n41972) );
  NAND2_X1 U44688 ( .A1(n41978), .A2(n41972), .ZN(n41973) );
  NAND2_X1 U44689 ( .A1(n41976), .A2(n41975), .ZN(n41990) );
  AND2_X1 U44690 ( .A1(n41980), .A2(n41979), .ZN(n41989) );
  OAI21_X1 U44691 ( .B1(n41984), .B2(n41983), .A(n41982), .ZN(n41988) );
  NAND2_X1 U44692 ( .A1(n41986), .A2(n41985), .ZN(n41987) );
  XNOR2_X1 U44693 ( .A(n46153), .B(n43609), .ZN(n43817) );
  XNOR2_X1 U44694 ( .A(n46150), .B(n41991), .ZN(n41993) );
  INV_X1 U44695 ( .A(n43048), .ZN(n41992) );
  XNOR2_X1 U44696 ( .A(n41993), .B(n41992), .ZN(n44185) );
  XNOR2_X1 U44697 ( .A(n44185), .B(n43817), .ZN(n41994) );
  XNOR2_X1 U44698 ( .A(n41995), .B(n41994), .ZN(n44825) );
  INV_X1 U44699 ( .A(n44825), .ZN(n44831) );
  XNOR2_X1 U44700 ( .A(n44027), .B(n41996), .ZN(n44521) );
  NAND2_X1 U44701 ( .A1(n41997), .A2(n42020), .ZN(n41998) );
  NAND2_X1 U44702 ( .A1(n41998), .A2(n42006), .ZN(n41999) );
  AOI21_X1 U44703 ( .B1(n42001), .B2(n42015), .A(n42010), .ZN(n42004) );
  NAND3_X1 U44704 ( .A1(n42005), .A2(n42004), .A3(n42003), .ZN(n42024) );
  INV_X1 U44705 ( .A(n42013), .ZN(n42009) );
  NAND4_X1 U44706 ( .A1(n42009), .A2(n42010), .A3(n42008), .A4(n42007), .ZN(
        n42017) );
  OAI211_X1 U44707 ( .C1(n42015), .C2(n42014), .A(n42013), .B(n42012), .ZN(
        n42016) );
  NAND2_X1 U44708 ( .A1(n42017), .A2(n42016), .ZN(n42023) );
  OAI211_X1 U44709 ( .C1(n42021), .C2(n42020), .A(n42019), .B(n42018), .ZN(
        n42022) );
  XNOR2_X1 U44710 ( .A(n44521), .B(n43856), .ZN(n42034) );
  XNOR2_X1 U44711 ( .A(n42025), .B(n42918), .ZN(n42027) );
  XNOR2_X1 U44712 ( .A(n42027), .B(n42026), .ZN(n42028) );
  XNOR2_X1 U44713 ( .A(n42029), .B(n42028), .ZN(n42030) );
  XNOR2_X1 U44714 ( .A(n43619), .B(n42030), .ZN(n42031) );
  XNOR2_X1 U44715 ( .A(n42031), .B(n2185), .ZN(n42032) );
  XNOR2_X1 U44716 ( .A(n43238), .B(n42032), .ZN(n42033) );
  XNOR2_X1 U44717 ( .A(n40814), .B(n43950), .ZN(n45416) );
  XNOR2_X1 U44718 ( .A(n42035), .B(n45416), .ZN(n42036) );
  XNOR2_X1 U44719 ( .A(n45279), .B(n44240), .ZN(n43569) );
  XNOR2_X1 U44720 ( .A(n44529), .B(n43569), .ZN(n42037) );
  NAND2_X1 U44721 ( .A1(n42039), .A2(n42441), .ZN(n42040) );
  AND2_X1 U44722 ( .A1(n42041), .A2(n42040), .ZN(n42437) );
  NAND2_X1 U44723 ( .A1(n42043), .A2(n42062), .ZN(n42046) );
  AND2_X1 U44724 ( .A1(n42046), .A2(n42045), .ZN(n42438) );
  AOI22_X1 U44725 ( .A1(n42047), .A2(n42438), .B1(n42443), .B2(n42441), .ZN(
        n42065) );
  NAND2_X1 U44726 ( .A1(n42051), .A2(n42050), .ZN(n42444) );
  OAI21_X1 U44727 ( .B1(n480), .B2(n42053), .A(n42052), .ZN(n42064) );
  OAI21_X1 U44728 ( .B1(n42056), .B2(n42055), .A(n42441), .ZN(n42060) );
  NAND2_X1 U44729 ( .A1(n42441), .A2(n42058), .ZN(n42059) );
  OAI211_X1 U44730 ( .C1(n42062), .C2(n42061), .A(n42060), .B(n42059), .ZN(
        n42063) );
  NAND2_X1 U44731 ( .A1(n42064), .A2(n42063), .ZN(n42445) );
  NAND4_X1 U44732 ( .A1(n42437), .A2(n42065), .A3(n42444), .A4(n42445), .ZN(
        n42066) );
  XNOR2_X1 U44733 ( .A(n42067), .B(n43833), .ZN(n46108) );
  XNOR2_X1 U44734 ( .A(n42869), .B(n42453), .ZN(n43707) );
  XNOR2_X1 U44735 ( .A(n46108), .B(n43707), .ZN(n42076) );
  XNOR2_X1 U44736 ( .A(n4624), .B(n4517), .ZN(n42068) );
  XNOR2_X1 U44737 ( .A(n44909), .B(n42068), .ZN(n42070) );
  XNOR2_X1 U44738 ( .A(n42070), .B(n42069), .ZN(n42071) );
  XNOR2_X1 U44739 ( .A(n43225), .B(n42071), .ZN(n42073) );
  XNOR2_X1 U44740 ( .A(n51406), .B(n44016), .ZN(n42072) );
  XNOR2_X1 U44741 ( .A(n42073), .B(n42072), .ZN(n42074) );
  XNOR2_X1 U44742 ( .A(n45252), .B(n42074), .ZN(n42075) );
  XNOR2_X1 U44743 ( .A(n42076), .B(n42075), .ZN(n42080) );
  XNOR2_X1 U44744 ( .A(n43219), .B(n44006), .ZN(n44913) );
  XNOR2_X1 U44745 ( .A(n44913), .B(n42570), .ZN(n42078) );
  XNOR2_X1 U44746 ( .A(n42078), .B(n45265), .ZN(n42079) );
  XNOR2_X1 U44747 ( .A(n42080), .B(n42079), .ZN(n42081) );
  NAND2_X1 U44748 ( .A1(n42180), .A2(n42081), .ZN(n44827) );
  INV_X1 U44749 ( .A(n44827), .ZN(n44281) );
  NOR2_X1 U44750 ( .A1(n45532), .A2(n44281), .ZN(n45522) );
  INV_X1 U44751 ( .A(n42180), .ZN(n44646) );
  INV_X1 U44752 ( .A(n42081), .ZN(n45828) );
  NAND2_X1 U44753 ( .A1(n45522), .A2(n45534), .ZN(n44814) );
  OR2_X1 U44755 ( .A1(n44822), .A2(n45827), .ZN(n45835) );
  NAND2_X1 U44756 ( .A1(n44814), .A2(n45835), .ZN(n42121) );
  XOR2_X1 U44757 ( .A(n42083), .B(n42082), .Z(n42085) );
  XNOR2_X1 U44758 ( .A(n42085), .B(n42084), .ZN(n42087) );
  INV_X1 U44759 ( .A(n42087), .ZN(n42093) );
  NAND2_X1 U44760 ( .A1(n42088), .A2(n42087), .ZN(n42091) );
  OAI211_X1 U44761 ( .C1(n42093), .C2(n42092), .A(n42091), .B(n42090), .ZN(
        n42094) );
  XNOR2_X1 U44762 ( .A(n42094), .B(n43380), .ZN(n42095) );
  XNOR2_X1 U44763 ( .A(n44353), .B(n44559), .ZN(n43925) );
  XNOR2_X1 U44764 ( .A(n42095), .B(n43925), .ZN(n42097) );
  XNOR2_X1 U44765 ( .A(n44561), .B(n4157), .ZN(n43754) );
  XNOR2_X1 U44766 ( .A(n44944), .B(n43754), .ZN(n42096) );
  XNOR2_X1 U44767 ( .A(n42097), .B(n42096), .ZN(n42099) );
  XNOR2_X1 U44768 ( .A(n42098), .B(n42099), .ZN(n42120) );
  XNOR2_X1 U44769 ( .A(n45099), .B(n42100), .ZN(n43658) );
  XNOR2_X1 U44770 ( .A(n45116), .B(n42101), .ZN(n44933) );
  XNOR2_X1 U44771 ( .A(n43155), .B(n42102), .ZN(n42117) );
  INV_X1 U44772 ( .A(n42103), .ZN(n42116) );
  INV_X1 U44773 ( .A(n42105), .ZN(n42107) );
  NAND4_X2 U44775 ( .A1(n42116), .A2(n42115), .A3(n42114), .A4(n42113), .ZN(
        n44134) );
  XNOR2_X1 U44776 ( .A(n44134), .B(n42117), .ZN(n46044) );
  XNOR2_X1 U44777 ( .A(n44933), .B(n46044), .ZN(n42118) );
  XNOR2_X1 U44778 ( .A(n43658), .B(n42118), .ZN(n42119) );
  INV_X1 U44779 ( .A(n42177), .ZN(n44813) );
  NAND2_X1 U44780 ( .A1(n42121), .A2(n44813), .ZN(n42189) );
  XNOR2_X1 U44781 ( .A(n42122), .B(n44547), .ZN(n42128) );
  XNOR2_X1 U44782 ( .A(n42123), .B(n1326), .ZN(n42124) );
  XNOR2_X1 U44783 ( .A(n42125), .B(n42124), .ZN(n42126) );
  XNOR2_X1 U44784 ( .A(n43781), .B(n42126), .ZN(n42127) );
  XNOR2_X1 U44785 ( .A(n42128), .B(n42127), .ZN(n42130) );
  XNOR2_X1 U44786 ( .A(n42129), .B(n42130), .ZN(n42168) );
  XNOR2_X1 U44787 ( .A(n44541), .B(n43915), .ZN(n43779) );
  AND2_X1 U44788 ( .A1(n42154), .A2(n42131), .ZN(n42134) );
  INV_X1 U44789 ( .A(n42132), .ZN(n42133) );
  OAI211_X1 U44790 ( .C1(n42135), .C2(n42145), .A(n42134), .B(n42133), .ZN(
        n42143) );
  NAND4_X1 U44791 ( .A1(n42139), .A2(n42138), .A3(n51375), .A4(n42136), .ZN(
        n42140) );
  INV_X1 U44792 ( .A(n42144), .ZN(n42147) );
  MUX2_X1 U44793 ( .A(n42147), .B(n42146), .S(n42145), .Z(n42165) );
  NOR2_X1 U44794 ( .A1(n42155), .A2(n42148), .ZN(n42150) );
  AOI22_X1 U44795 ( .A1(n42152), .A2(n42151), .B1(n42150), .B2(n42149), .ZN(
        n42164) );
  XNOR2_X1 U44796 ( .A(n42153), .B(n42154), .ZN(n42162) );
  NAND2_X1 U44797 ( .A1(n42155), .A2(n42154), .ZN(n42161) );
  AND2_X1 U44798 ( .A1(n42157), .A2(n52092), .ZN(n42160) );
  INV_X1 U44799 ( .A(n42158), .ZN(n42159) );
  NAND4_X1 U44800 ( .A1(n42162), .A2(n42161), .A3(n42160), .A4(n42159), .ZN(
        n42163) );
  XNOR2_X1 U44801 ( .A(n45421), .B(n43170), .ZN(n43059) );
  XNOR2_X1 U44803 ( .A(n46060), .B(n43779), .ZN(n42167) );
  XNOR2_X1 U44804 ( .A(n42168), .B(n42167), .ZN(n42174) );
  XNOR2_X1 U44805 ( .A(n42284), .B(n43635), .ZN(n42528) );
  XNOR2_X1 U44806 ( .A(n42528), .B(n44534), .ZN(n42169) );
  XNOR2_X1 U44807 ( .A(n42169), .B(n45122), .ZN(n45437) );
  XNOR2_X1 U44808 ( .A(n51464), .B(n44198), .ZN(n42530) );
  XNOR2_X1 U44809 ( .A(n42530), .B(n43168), .ZN(n44326) );
  XNOR2_X1 U44810 ( .A(n42170), .B(n4847), .ZN(n42171) );
  XNOR2_X1 U44811 ( .A(n42171), .B(n44542), .ZN(n44064) );
  XNOR2_X1 U44812 ( .A(n44064), .B(n44326), .ZN(n42172) );
  XNOR2_X1 U44813 ( .A(n45437), .B(n42172), .ZN(n42173) );
  OR2_X1 U44815 ( .A1(n42176), .A2(n45834), .ZN(n42178) );
  NOR2_X1 U44816 ( .A1(n42178), .A2(n45533), .ZN(n44832) );
  NOR2_X1 U44817 ( .A1(n42179), .A2(n44832), .ZN(n42188) );
  AND2_X1 U44818 ( .A1(n44640), .A2(n44825), .ZN(n44643) );
  AOI21_X1 U44819 ( .B1(n45819), .B2(n42176), .A(n44643), .ZN(n42184) );
  INV_X1 U44820 ( .A(n44280), .ZN(n44811) );
  NAND3_X1 U44821 ( .A1(n44811), .A2(n45524), .A3(n44831), .ZN(n42183) );
  INV_X1 U44822 ( .A(n44640), .ZN(n45829) );
  OR2_X1 U44823 ( .A1(n45829), .A2(n44828), .ZN(n42182) );
  OAI211_X1 U44824 ( .C1(n42184), .C2(n45834), .A(n42183), .B(n42182), .ZN(
        n42185) );
  INV_X1 U44825 ( .A(n42185), .ZN(n42187) );
  NAND2_X1 U44826 ( .A1(n42181), .A2(n44825), .ZN(n45830) );
  NOR2_X1 U44827 ( .A1(n45533), .A2(n45830), .ZN(n45530) );
  NAND2_X1 U44828 ( .A1(n45530), .A2(n44646), .ZN(n42186) );
  NAND4_X2 U44829 ( .A1(n42187), .A2(n42188), .A3(n42189), .A4(n42186), .ZN(
        n47831) );
  AND2_X1 U44830 ( .A1(n47842), .A2(n51285), .ZN(n42190) );
  MUX2_X1 U44831 ( .A(n47873), .B(n42190), .S(n47879), .Z(n42191) );
  NAND2_X1 U44832 ( .A1(n651), .A2(n47869), .ZN(n47874) );
  INV_X1 U44833 ( .A(n47874), .ZN(n47817) );
  NOR2_X1 U44834 ( .A1(n47879), .A2(n51469), .ZN(n47885) );
  NAND3_X1 U44835 ( .A1(n47885), .A2(n47842), .A3(n3798), .ZN(n42194) );
  NAND3_X1 U44836 ( .A1(n47831), .A2(n47873), .A3(n508), .ZN(n47834) );
  NAND2_X1 U44837 ( .A1(n47841), .A2(n42192), .ZN(n47880) );
  NOR2_X1 U44838 ( .A1(n47869), .A2(n47841), .ZN(n47850) );
  NAND2_X1 U44839 ( .A1(n47866), .A2(n47850), .ZN(n42196) );
  INV_X1 U44840 ( .A(n47880), .ZN(n42195) );
  NAND2_X1 U44841 ( .A1(n42195), .A2(n47855), .ZN(n47872) );
  NAND3_X1 U44842 ( .A1(n42198), .A2(n42197), .A3(n8769), .ZN(n42200) );
  INV_X1 U44843 ( .A(n4045), .ZN(n42199) );
  XNOR2_X1 U44844 ( .A(n42200), .B(n42199), .ZN(Plaintext[27]) );
  XNOR2_X1 U44845 ( .A(n44901), .B(n52058), .ZN(n42670) );
  NOR2_X1 U44846 ( .A1(n42202), .A2(n42201), .ZN(n42204) );
  AOI22_X1 U44847 ( .A1(n42206), .A2(n6578), .B1(n42204), .B2(n42203), .ZN(
        n42211) );
  NAND2_X1 U44848 ( .A1(n42208), .A2(n42207), .ZN(n42210) );
  MUX2_X1 U44849 ( .A(n42211), .B(n42210), .S(n42209), .Z(n42213) );
  NAND2_X1 U44850 ( .A1(n42213), .A2(n42212), .ZN(n44286) );
  XNOR2_X1 U44851 ( .A(n43216), .B(n44286), .ZN(n46102) );
  XNOR2_X1 U44852 ( .A(n43661), .B(n46102), .ZN(n42221) );
  XNOR2_X1 U44853 ( .A(n42215), .B(n42214), .ZN(n42216) );
  XNOR2_X1 U44854 ( .A(n42863), .B(n42216), .ZN(n42217) );
  XNOR2_X1 U44855 ( .A(n45263), .B(n42217), .ZN(n42219) );
  XNOR2_X1 U44856 ( .A(n42219), .B(n42218), .ZN(n42220) );
  XNOR2_X1 U44857 ( .A(n42221), .B(n42220), .ZN(n42223) );
  XNOR2_X1 U44858 ( .A(n51525), .B(n42223), .ZN(n45209) );
  XNOR2_X1 U44859 ( .A(n42850), .B(n51450), .ZN(n42224) );
  XNOR2_X1 U44860 ( .A(n51431), .B(n43623), .ZN(n42225) );
  XNOR2_X1 U44861 ( .A(n44879), .B(n42225), .ZN(n43301) );
  INV_X1 U44862 ( .A(n43301), .ZN(n42231) );
  XNOR2_X1 U44863 ( .A(n42227), .B(n42226), .ZN(n42228) );
  XNOR2_X1 U44864 ( .A(n43131), .B(n42228), .ZN(n42229) );
  XNOR2_X1 U44865 ( .A(n42229), .B(n46112), .ZN(n42230) );
  XNOR2_X1 U44866 ( .A(n42231), .B(n42230), .ZN(n42232) );
  XNOR2_X1 U44867 ( .A(n42414), .B(n42232), .ZN(n42238) );
  XNOR2_X1 U44868 ( .A(n42233), .B(n44027), .ZN(n42234) );
  XNOR2_X1 U44869 ( .A(n42234), .B(n51390), .ZN(n42853) );
  XNOR2_X1 U44870 ( .A(n51100), .B(n43244), .ZN(n42235) );
  XNOR2_X1 U44871 ( .A(n42853), .B(n42236), .ZN(n42237) );
  INV_X1 U44872 ( .A(n42271), .ZN(n44784) );
  XNOR2_X1 U44873 ( .A(n43209), .B(n45445), .ZN(n42239) );
  XNOR2_X1 U44874 ( .A(n42786), .B(n42239), .ZN(n42248) );
  XNOR2_X1 U44875 ( .A(n42240), .B(n3367), .ZN(n42242) );
  XNOR2_X1 U44876 ( .A(n42242), .B(n42241), .ZN(n42244) );
  XNOR2_X1 U44877 ( .A(n42244), .B(n42243), .ZN(n42245) );
  XNOR2_X1 U44878 ( .A(n45114), .B(n42245), .ZN(n42246) );
  XNOR2_X1 U44879 ( .A(n42246), .B(n43157), .ZN(n42247) );
  XNOR2_X1 U44882 ( .A(n43380), .B(n44044), .ZN(n42250) );
  XNOR2_X1 U44883 ( .A(n42250), .B(n43928), .ZN(n42251) );
  XNOR2_X1 U44884 ( .A(n45321), .B(n42251), .ZN(n43214) );
  XNOR2_X1 U44885 ( .A(n45306), .B(n4564), .ZN(n42253) );
  XNOR2_X1 U44886 ( .A(n45454), .B(n42253), .ZN(n42600) );
  INV_X1 U44887 ( .A(n42600), .ZN(n42254) );
  AND2_X1 U44888 ( .A1(n46243), .A2(n540), .ZN(n45215) );
  XNOR2_X1 U44889 ( .A(n45355), .B(n46138), .ZN(n42257) );
  XNOR2_X1 U44890 ( .A(n42329), .B(n4923), .ZN(n42255) );
  XNOR2_X1 U44891 ( .A(n50967), .B(n42255), .ZN(n42256) );
  XNOR2_X1 U44892 ( .A(n42257), .B(n42256), .ZN(n42260) );
  INV_X1 U44893 ( .A(n42258), .ZN(n42259) );
  XNOR2_X1 U44894 ( .A(n44374), .B(n42259), .ZN(n44184) );
  XNOR2_X1 U44895 ( .A(n42260), .B(n44184), .ZN(n42263) );
  XNOR2_X1 U44896 ( .A(n43254), .B(n42261), .ZN(n42262) );
  XNOR2_X1 U44897 ( .A(n43048), .B(n42262), .ZN(n42473) );
  XNOR2_X1 U44898 ( .A(n42264), .B(n42534), .ZN(n43604) );
  XNOR2_X1 U44899 ( .A(n44176), .B(n44182), .ZN(n42265) );
  XNOR2_X1 U44900 ( .A(n42265), .B(n51096), .ZN(n42269) );
  XNOR2_X1 U44901 ( .A(n42961), .B(n42266), .ZN(n42267) );
  XNOR2_X1 U44902 ( .A(n42267), .B(n43113), .ZN(n42268) );
  XNOR2_X1 U44903 ( .A(n43604), .B(n42872), .ZN(n42270) );
  OR2_X1 U44904 ( .A1(n45209), .A2(n49163), .ZN(n44783) );
  INV_X1 U44905 ( .A(n44783), .ZN(n49159) );
  AOI21_X1 U44906 ( .B1(n45215), .B2(n49161), .A(n49159), .ZN(n42310) );
  XNOR2_X1 U44907 ( .A(n46060), .B(n42272), .ZN(n42273) );
  XNOR2_X1 U44908 ( .A(n42273), .B(n43197), .ZN(n42953) );
  XNOR2_X1 U44909 ( .A(n42275), .B(n42274), .ZN(n42276) );
  XNOR2_X1 U44910 ( .A(n45293), .B(n42276), .ZN(n42277) );
  XNOR2_X1 U44911 ( .A(n42277), .B(n44547), .ZN(n42279) );
  XNOR2_X1 U44912 ( .A(n42278), .B(n46068), .ZN(n45429) );
  XNOR2_X1 U44913 ( .A(n45429), .B(n42279), .ZN(n42281) );
  XNOR2_X1 U44914 ( .A(n42281), .B(n42280), .ZN(n42282) );
  XNOR2_X1 U44915 ( .A(n42284), .B(n42283), .ZN(n42285) );
  XNOR2_X1 U44916 ( .A(n46058), .B(n42285), .ZN(n42286) );
  XNOR2_X1 U44917 ( .A(n42287), .B(n42286), .ZN(n43645) );
  AOI21_X1 U44918 ( .B1(n49159), .B2(n46252), .A(n46255), .ZN(n42304) );
  NAND2_X1 U44919 ( .A1(n49177), .A2(n539), .ZN(n49168) );
  NAND2_X1 U44921 ( .A1(n49163), .A2(n49161), .ZN(n46257) );
  NAND3_X1 U44922 ( .A1(n51376), .A2(n46244), .A3(n46257), .ZN(n42303) );
  XNOR2_X1 U44923 ( .A(n45490), .B(n42289), .ZN(n44081) );
  INV_X1 U44924 ( .A(n45068), .ZN(n42290) );
  XNOR2_X1 U44925 ( .A(n44081), .B(n42290), .ZN(n43763) );
  XNOR2_X1 U44926 ( .A(n43763), .B(n45344), .ZN(n42302) );
  XNOR2_X1 U44927 ( .A(n43079), .B(n43596), .ZN(n42491) );
  XNOR2_X1 U44928 ( .A(n44153), .B(n42291), .ZN(n44482) );
  XNOR2_X1 U44929 ( .A(n4823), .B(n4204), .ZN(n42292) );
  XNOR2_X1 U44930 ( .A(n42293), .B(n42292), .ZN(n42294) );
  XNOR2_X1 U44931 ( .A(n51460), .B(n42294), .ZN(n42295) );
  XNOR2_X1 U44932 ( .A(n44482), .B(n42295), .ZN(n42296) );
  XNOR2_X1 U44933 ( .A(n42491), .B(n42296), .ZN(n42300) );
  XNOR2_X1 U44934 ( .A(n42316), .B(n42980), .ZN(n45486) );
  XNOR2_X1 U44935 ( .A(n52125), .B(n42297), .ZN(n42298) );
  XNOR2_X1 U44936 ( .A(n45486), .B(n42298), .ZN(n42556) );
  INV_X1 U44937 ( .A(n42556), .ZN(n42299) );
  XNOR2_X1 U44938 ( .A(n42300), .B(n42299), .ZN(n42301) );
  XNOR2_X1 U44939 ( .A(n42302), .B(n42301), .ZN(n42305) );
  INV_X1 U44940 ( .A(n42305), .ZN(n46249) );
  NAND2_X1 U44941 ( .A1(n45649), .A2(n46249), .ZN(n49174) );
  NAND3_X1 U44942 ( .A1(n46249), .A2(n49163), .A3(n49170), .ZN(n42306) );
  OAI21_X1 U44943 ( .B1(n45648), .B2(n49174), .A(n42306), .ZN(n42307) );
  NAND2_X1 U44944 ( .A1(n42307), .A2(n540), .ZN(n42308) );
  INV_X1 U44945 ( .A(Key[160]), .ZN(n50546) );
  XNOR2_X1 U44946 ( .A(n4204), .B(n4835), .ZN(n42311) );
  XNOR2_X1 U44947 ( .A(n42311), .B(n49109), .ZN(n42312) );
  XNOR2_X1 U44948 ( .A(n42712), .B(n42312), .ZN(n42313) );
  XNOR2_X1 U44949 ( .A(n42314), .B(n42313), .ZN(n42315) );
  XNOR2_X1 U44950 ( .A(n42316), .B(n42315), .ZN(n42317) );
  XNOR2_X1 U44951 ( .A(n51494), .B(n42318), .ZN(n42320) );
  XNOR2_X1 U44952 ( .A(n52103), .B(n43890), .ZN(n42319) );
  XNOR2_X1 U44953 ( .A(n42319), .B(n42504), .ZN(n42985) );
  INV_X1 U44955 ( .A(n42980), .ZN(n42321) );
  XNOR2_X1 U44956 ( .A(n43889), .B(n42321), .ZN(n44395) );
  INV_X1 U44957 ( .A(n44395), .ZN(n42896) );
  XNOR2_X1 U44958 ( .A(n43102), .B(n42322), .ZN(n42323) );
  XNOR2_X1 U44959 ( .A(n42323), .B(n44153), .ZN(n44077) );
  XNOR2_X1 U44960 ( .A(n42896), .B(n44077), .ZN(n42324) );
  XNOR2_X1 U44961 ( .A(n43272), .B(n42324), .ZN(n42682) );
  XNOR2_X1 U44963 ( .A(n46138), .B(n43723), .ZN(n42326) );
  XNOR2_X1 U44964 ( .A(n42327), .B(n2203), .ZN(n42328) );
  XNOR2_X1 U44965 ( .A(n42329), .B(n42328), .ZN(n42330) );
  XNOR2_X1 U44966 ( .A(n42331), .B(n42330), .ZN(n42332) );
  XNOR2_X1 U44967 ( .A(n42961), .B(n42332), .ZN(n42333) );
  XNOR2_X1 U44968 ( .A(n42333), .B(n43113), .ZN(n42334) );
  XNOR2_X1 U44969 ( .A(n42335), .B(n42334), .ZN(n42336) );
  XNOR2_X1 U44970 ( .A(n42336), .B(n44096), .ZN(n42338) );
  XNOR2_X1 U44971 ( .A(n43354), .B(n45355), .ZN(n42470) );
  XNOR2_X1 U44972 ( .A(n44098), .B(n42470), .ZN(n42337) );
  XNOR2_X1 U44973 ( .A(n42534), .B(n43363), .ZN(n44503) );
  XNOR2_X1 U44974 ( .A(n42337), .B(n44503), .ZN(n42698) );
  OR2_X1 U44975 ( .A1(n46203), .A2(n52086), .ZN(n49270) );
  XNOR2_X1 U44976 ( .A(n52089), .B(n51408), .ZN(n44009) );
  XNOR2_X1 U44977 ( .A(n42863), .B(n42339), .ZN(n42340) );
  XNOR2_X1 U44978 ( .A(n42341), .B(n44009), .ZN(n42916) );
  XNOR2_X1 U44979 ( .A(n2183), .B(n4932), .ZN(n42858) );
  XNOR2_X1 U44980 ( .A(n42342), .B(n42858), .ZN(n42343) );
  XNOR2_X1 U44981 ( .A(n42344), .B(n42343), .ZN(n42345) );
  XNOR2_X1 U44982 ( .A(n43123), .B(n42345), .ZN(n42346) );
  XNOR2_X1 U44983 ( .A(n45393), .B(n42346), .ZN(n42347) );
  XNOR2_X1 U44984 ( .A(n44209), .B(n44911), .ZN(n42662) );
  XNOR2_X1 U44985 ( .A(n51509), .B(n42347), .ZN(n42348) );
  XNOR2_X1 U44986 ( .A(n43696), .B(n42349), .ZN(n42350) );
  XNOR2_X1 U44987 ( .A(n42353), .B(n42352), .ZN(n42361) );
  XNOR2_X1 U44988 ( .A(n43950), .B(n43623), .ZN(n42354) );
  XNOR2_X1 U44989 ( .A(n42354), .B(n43244), .ZN(n44032) );
  XNOR2_X1 U44990 ( .A(n42356), .B(n42355), .ZN(n42357) );
  XNOR2_X1 U44991 ( .A(n44314), .B(n42357), .ZN(n42358) );
  XNOR2_X1 U44992 ( .A(n44032), .B(n42359), .ZN(n42360) );
  XNOR2_X1 U44993 ( .A(n42361), .B(n42360), .ZN(n42364) );
  XNOR2_X1 U44994 ( .A(n44030), .B(n43131), .ZN(n42640) );
  XNOR2_X1 U44995 ( .A(n42640), .B(n43143), .ZN(n42362) );
  XNOR2_X1 U44996 ( .A(n44320), .B(n42362), .ZN(n42363) );
  NOR2_X1 U44997 ( .A1(n49270), .A2(n45667), .ZN(n42365) );
  AND2_X1 U44998 ( .A1(n49274), .A2(n46196), .ZN(n49261) );
  INV_X1 U44999 ( .A(n49261), .ZN(n46204) );
  XNOR2_X1 U45000 ( .A(n42367), .B(n42366), .ZN(n42368) );
  XNOR2_X1 U45001 ( .A(n42369), .B(n42368), .ZN(n42370) );
  XNOR2_X1 U45002 ( .A(n43155), .B(n42370), .ZN(n42371) );
  XNOR2_X1 U45003 ( .A(n42371), .B(n45116), .ZN(n42373) );
  XNOR2_X1 U45004 ( .A(n43157), .B(n44130), .ZN(n42372) );
  XNOR2_X1 U45005 ( .A(n42373), .B(n42372), .ZN(n42375) );
  INV_X1 U45006 ( .A(n43374), .ZN(n44133) );
  XNOR2_X1 U45007 ( .A(n44133), .B(n45114), .ZN(n42374) );
  XNOR2_X1 U45008 ( .A(n42590), .B(n4554), .ZN(n42376) );
  XNOR2_X1 U45009 ( .A(n42376), .B(n43928), .ZN(n44567) );
  XNOR2_X1 U45010 ( .A(n43209), .B(n43014), .ZN(n42791) );
  XNOR2_X1 U45011 ( .A(n44567), .B(n42791), .ZN(n44040) );
  XNOR2_X1 U45012 ( .A(n45454), .B(n42377), .ZN(n42378) );
  XNOR2_X1 U45013 ( .A(n45285), .B(n4755), .ZN(n42381) );
  XNOR2_X1 U45014 ( .A(n44923), .B(n42381), .ZN(n42382) );
  XNOR2_X1 U45015 ( .A(n42385), .B(n42384), .ZN(n42386) );
  XNOR2_X1 U45016 ( .A(n43170), .B(n3383), .ZN(n44342) );
  XNOR2_X1 U45017 ( .A(n42387), .B(n44342), .ZN(n42388) );
  XNOR2_X1 U45018 ( .A(n43635), .B(n44547), .ZN(n44066) );
  XNOR2_X1 U45019 ( .A(n42388), .B(n44066), .ZN(n42389) );
  XNOR2_X1 U45020 ( .A(n44055), .B(n42389), .ZN(n42392) );
  XNOR2_X1 U45021 ( .A(n44190), .B(n45293), .ZN(n42623) );
  XNOR2_X1 U45022 ( .A(n42623), .B(n52222), .ZN(n42390) );
  XNOR2_X1 U45023 ( .A(n44056), .B(n42390), .ZN(n42391) );
  OR2_X1 U45024 ( .A1(n49273), .A2(n51335), .ZN(n42394) );
  AND2_X1 U45025 ( .A1(n46203), .A2(n46201), .ZN(n45671) );
  INV_X1 U45026 ( .A(n46199), .ZN(n49262) );
  INV_X1 U45027 ( .A(n49263), .ZN(n49266) );
  NAND3_X1 U45028 ( .A1(n45671), .A2(n49262), .A3(n49275), .ZN(n42393) );
  OAI21_X1 U45029 ( .B1(n42394), .B2(n49267), .A(n42393), .ZN(n42397) );
  AND2_X1 U45030 ( .A1(n46196), .A2(n46201), .ZN(n44775) );
  OR2_X1 U45031 ( .A1(n44775), .A2(n46203), .ZN(n42395) );
  NOR2_X1 U45032 ( .A1(n45679), .A2(n42395), .ZN(n42396) );
  NAND3_X1 U45033 ( .A1(n666), .A2(n49263), .A3(n46196), .ZN(n42398) );
  NAND2_X1 U45034 ( .A1(n42398), .A2(n46201), .ZN(n42399) );
  NAND2_X1 U45035 ( .A1(n42399), .A2(n46203), .ZN(n42400) );
  NAND2_X1 U45036 ( .A1(n42401), .A2(n42400), .ZN(n42404) );
  AND2_X1 U45037 ( .A1(n49263), .A2(n666), .ZN(n45668) );
  INV_X1 U45038 ( .A(n45668), .ZN(n45680) );
  NAND2_X1 U45039 ( .A1(n49261), .A2(n49273), .ZN(n45665) );
  AOI21_X1 U45040 ( .B1(n49275), .B2(n45670), .A(n46201), .ZN(n42402) );
  OAI211_X1 U45041 ( .C1(n45680), .C2(n51335), .A(n45665), .B(n42402), .ZN(
        n42403) );
  MUX2_X1 U45042 ( .A(n45667), .B(n49261), .S(n46201), .Z(n42405) );
  AND2_X1 U45043 ( .A1(n49266), .A2(n666), .ZN(n49277) );
  OAI21_X1 U45044 ( .B1(n42405), .B2(n49278), .A(n49277), .ZN(n42406) );
  XNOR2_X1 U45045 ( .A(n43139), .B(n43623), .ZN(n42407) );
  XNOR2_X1 U45046 ( .A(n42407), .B(n51681), .ZN(n42584) );
  XNOR2_X1 U45047 ( .A(n42409), .B(n42408), .ZN(n42410) );
  XNOR2_X1 U45048 ( .A(n44314), .B(n42410), .ZN(n42411) );
  XNOR2_X1 U45049 ( .A(n42584), .B(n42412), .ZN(n42413) );
  XNOR2_X1 U45050 ( .A(n42414), .B(n42413), .ZN(n42418) );
  XNOR2_X1 U45051 ( .A(n45408), .B(n46113), .ZN(n42415) );
  XNOR2_X1 U45052 ( .A(n42415), .B(n46112), .ZN(n43962) );
  INV_X1 U45053 ( .A(n45269), .ZN(n42416) );
  XNOR2_X1 U45054 ( .A(n43962), .B(n42416), .ZN(n42417) );
  XNOR2_X1 U45055 ( .A(n42417), .B(n44320), .ZN(n44036) );
  XNOR2_X1 U45056 ( .A(n44036), .B(n42418), .ZN(n42508) );
  INV_X1 U45057 ( .A(n45305), .ZN(n44041) );
  XNOR2_X1 U45058 ( .A(n44041), .B(n44134), .ZN(n42422) );
  XNOR2_X1 U45059 ( .A(n42780), .B(n42419), .ZN(n42420) );
  XNOR2_X1 U45060 ( .A(n45314), .B(n42420), .ZN(n42421) );
  XNOR2_X1 U45061 ( .A(n42422), .B(n42421), .ZN(n42423) );
  XNOR2_X1 U45062 ( .A(n42423), .B(n42788), .ZN(n42426) );
  XNOR2_X1 U45063 ( .A(n43547), .B(n4565), .ZN(n42424) );
  XNOR2_X1 U45064 ( .A(n42424), .B(n44561), .ZN(n42425) );
  XNOR2_X1 U45065 ( .A(n42425), .B(n43929), .ZN(n42942) );
  XNOR2_X1 U45066 ( .A(n42426), .B(n42942), .ZN(n42432) );
  XNOR2_X1 U45067 ( .A(n43157), .B(n43380), .ZN(n42427) );
  XNOR2_X1 U45068 ( .A(n42786), .B(n42427), .ZN(n42428) );
  XNOR2_X1 U45069 ( .A(n516), .B(n42428), .ZN(n42429) );
  XNOR2_X1 U45070 ( .A(n42429), .B(n42430), .ZN(n42431) );
  AND2_X1 U45071 ( .A1(n42508), .A2(n46444), .ZN(n42512) );
  INV_X1 U45072 ( .A(n42433), .ZN(n42435) );
  XNOR2_X1 U45073 ( .A(n42435), .B(n42434), .ZN(n42436) );
  XNOR2_X1 U45074 ( .A(n43225), .B(n42436), .ZN(n42448) );
  INV_X1 U45075 ( .A(n42438), .ZN(n42439) );
  OAI21_X1 U45076 ( .B1(n42443), .B2(n42442), .A(n42441), .ZN(n42446) );
  XNOR2_X1 U45078 ( .A(n44288), .B(n44287), .ZN(n42746) );
  INV_X1 U45079 ( .A(n42746), .ZN(n42451) );
  XNOR2_X1 U45080 ( .A(n42456), .B(n42455), .ZN(n43843) );
  XNOR2_X1 U45081 ( .A(n42457), .B(n43843), .ZN(n48456) );
  XNOR2_X1 U45083 ( .A(n42458), .B(n44370), .ZN(n42459) );
  XNOR2_X1 U45084 ( .A(n42461), .B(n42460), .ZN(n42465) );
  XNOR2_X1 U45085 ( .A(n4895), .B(n4655), .ZN(n42462) );
  XNOR2_X1 U45086 ( .A(n42754), .B(n42462), .ZN(n42463) );
  XNOR2_X1 U45087 ( .A(n42463), .B(n45348), .ZN(n42464) );
  XNOR2_X1 U45088 ( .A(n42465), .B(n42464), .ZN(n42466) );
  XNOR2_X1 U45089 ( .A(n51323), .B(n42466), .ZN(n42467) );
  XNOR2_X1 U45090 ( .A(n45460), .B(n42467), .ZN(n42468) );
  XNOR2_X1 U45091 ( .A(n42469), .B(n42468), .ZN(n42472) );
  XNOR2_X1 U45092 ( .A(n42470), .B(n43819), .ZN(n42471) );
  XNOR2_X1 U45093 ( .A(n42472), .B(n42471), .ZN(n42474) );
  XNOR2_X1 U45094 ( .A(n42474), .B(n42473), .ZN(n42475) );
  INV_X1 U45095 ( .A(n44378), .ZN(n43828) );
  INV_X1 U45097 ( .A(n42476), .ZN(n42478) );
  XNOR2_X1 U45098 ( .A(n42478), .B(n42477), .ZN(n42479) );
  XNOR2_X1 U45099 ( .A(n44198), .B(n42479), .ZN(n42480) );
  XNOR2_X1 U45100 ( .A(n42480), .B(n45293), .ZN(n42481) );
  XNOR2_X1 U45101 ( .A(n44190), .B(n49887), .ZN(n43391) );
  XNOR2_X1 U45102 ( .A(n42481), .B(n43391), .ZN(n42484) );
  XNOR2_X1 U45103 ( .A(n45421), .B(n671), .ZN(n42482) );
  XNOR2_X1 U45104 ( .A(n45432), .B(n42482), .ZN(n42483) );
  XNOR2_X1 U45105 ( .A(n42484), .B(n42483), .ZN(n42485) );
  XNOR2_X1 U45106 ( .A(n42486), .B(n42485), .ZN(n42488) );
  XNOR2_X2 U45107 ( .A(n42488), .B(n42487), .ZN(n45614) );
  AOI21_X1 U45108 ( .B1(n46446), .B2(n45614), .A(n48459), .ZN(n42489) );
  INV_X1 U45109 ( .A(n45614), .ZN(n48451) );
  XNOR2_X1 U45111 ( .A(n42715), .B(n44074), .ZN(n45331) );
  XNOR2_X1 U45112 ( .A(n44160), .B(n4613), .ZN(n46090) );
  XNOR2_X1 U45113 ( .A(n45331), .B(n46090), .ZN(n42490) );
  XNOR2_X1 U45114 ( .A(n42491), .B(n42490), .ZN(n42495) );
  XNOR2_X1 U45115 ( .A(n43102), .B(n42492), .ZN(n42493) );
  XNOR2_X1 U45116 ( .A(n42493), .B(n44153), .ZN(n42494) );
  XNOR2_X1 U45117 ( .A(n42494), .B(n45068), .ZN(n44397) );
  XNOR2_X1 U45118 ( .A(n42495), .B(n44397), .ZN(n42507) );
  INV_X1 U45119 ( .A(n42496), .ZN(n42498) );
  XNOR2_X1 U45120 ( .A(n43766), .B(n43263), .ZN(n42497) );
  XNOR2_X1 U45121 ( .A(n42498), .B(n42497), .ZN(n42499) );
  XNOR2_X1 U45122 ( .A(n42500), .B(n42499), .ZN(n42502) );
  XNOR2_X1 U45123 ( .A(n42502), .B(n42501), .ZN(n42503) );
  XNOR2_X1 U45124 ( .A(n42503), .B(n42896), .ZN(n42505) );
  XNOR2_X1 U45125 ( .A(n42505), .B(n43892), .ZN(n42506) );
  AOI21_X1 U45126 ( .B1(n48449), .B2(n48457), .A(n46434), .ZN(n42511) );
  INV_X1 U45127 ( .A(n46441), .ZN(n42510) );
  INV_X1 U45128 ( .A(n42508), .ZN(n46412) );
  NOR2_X1 U45129 ( .A1(n7275), .A2(n51732), .ZN(n46411) );
  OAI21_X1 U45130 ( .B1(n42511), .B2(n42510), .A(n42509), .ZN(n42514) );
  INV_X1 U45131 ( .A(n48463), .ZN(n46415) );
  AND2_X1 U45132 ( .A1(n8569), .A2(n48459), .ZN(n48465) );
  INV_X1 U45133 ( .A(n48465), .ZN(n45207) );
  NAND2_X1 U45134 ( .A1(n45614), .A2(n46444), .ZN(n46435) );
  XNOR2_X1 U45137 ( .A(n44546), .B(n52222), .ZN(n42519) );
  INV_X1 U45138 ( .A(n44547), .ZN(n42517) );
  XNOR2_X1 U45139 ( .A(n45284), .B(n671), .ZN(n42525) );
  XNOR2_X1 U45140 ( .A(n42520), .B(n4847), .ZN(n42521) );
  XNOR2_X1 U45141 ( .A(n42522), .B(n42521), .ZN(n42523) );
  XNOR2_X1 U45142 ( .A(n44189), .B(n42523), .ZN(n42524) );
  XNOR2_X1 U45143 ( .A(n42525), .B(n42524), .ZN(n42526) );
  XNOR2_X1 U45144 ( .A(n52130), .B(n42526), .ZN(n42527) );
  INV_X1 U45145 ( .A(n46058), .ZN(n42949) );
  XNOR2_X1 U45146 ( .A(n42528), .B(n42949), .ZN(n43916) );
  XNOR2_X1 U45147 ( .A(n42529), .B(n42530), .ZN(n42531) );
  XNOR2_X1 U45148 ( .A(n42531), .B(n43916), .ZN(n42796) );
  XNOR2_X1 U45149 ( .A(n45467), .B(n44370), .ZN(n44177) );
  XNOR2_X1 U45150 ( .A(n43723), .B(n2203), .ZN(n42532) );
  XNOR2_X1 U45151 ( .A(n44177), .B(n42532), .ZN(n42762) );
  XNOR2_X1 U45153 ( .A(n43609), .B(n45355), .ZN(n42535) );
  INV_X1 U45155 ( .A(n4655), .ZN(n50077) );
  XNOR2_X1 U45156 ( .A(n42537), .B(n50077), .ZN(n42538) );
  XNOR2_X1 U45157 ( .A(n42539), .B(n42538), .ZN(n42540) );
  XNOR2_X1 U45158 ( .A(n42541), .B(n42540), .ZN(n42542) );
  XNOR2_X1 U45159 ( .A(n46137), .B(n42542), .ZN(n42543) );
  XNOR2_X1 U45160 ( .A(n42543), .B(n44182), .ZN(n42544) );
  XNOR2_X1 U45161 ( .A(n46138), .B(n45354), .ZN(n44086) );
  XNOR2_X1 U45162 ( .A(n42544), .B(n44086), .ZN(n42545) );
  XNOR2_X1 U45163 ( .A(n43360), .B(n42545), .ZN(n42546) );
  INV_X1 U45164 ( .A(n42605), .ZN(n45238) );
  AND2_X1 U45165 ( .A1(n46267), .A2(n45238), .ZN(n46360) );
  XNOR2_X1 U45166 ( .A(n45333), .B(n47679), .ZN(n42548) );
  XNOR2_X1 U45167 ( .A(n42549), .B(n42548), .ZN(n42550) );
  XNOR2_X1 U45168 ( .A(n42551), .B(n42550), .ZN(n42552) );
  XNOR2_X1 U45169 ( .A(n43106), .B(n42552), .ZN(n42553) );
  XNOR2_X1 U45170 ( .A(n42554), .B(n42553), .ZN(n42555) );
  XNOR2_X1 U45171 ( .A(n42556), .B(n42555), .ZN(n42557) );
  XNOR2_X1 U45172 ( .A(n42557), .B(n45476), .ZN(n42559) );
  XNOR2_X1 U45173 ( .A(n51494), .B(n44397), .ZN(n42558) );
  XNOR2_X2 U45174 ( .A(n42559), .B(n42558), .ZN(n46356) );
  XNOR2_X1 U45176 ( .A(n42563), .B(n42562), .ZN(n42564) );
  XNOR2_X1 U45177 ( .A(n43696), .B(n42564), .ZN(n42565) );
  XNOR2_X1 U45178 ( .A(n44296), .B(n42565), .ZN(n42566) );
  XNOR2_X1 U45179 ( .A(n42567), .B(n42566), .ZN(n42568) );
  XNOR2_X1 U45180 ( .A(n44901), .B(n45390), .ZN(n43700) );
  XNOR2_X1 U45181 ( .A(n43700), .B(n42568), .ZN(n42574) );
  INV_X1 U45182 ( .A(n44006), .ZN(n43832) );
  XNOR2_X1 U45183 ( .A(n43832), .B(n45263), .ZN(n42569) );
  XNOR2_X1 U45184 ( .A(n42569), .B(n45393), .ZN(n42906) );
  INV_X1 U45185 ( .A(n42906), .ZN(n42868) );
  XNOR2_X1 U45186 ( .A(n45389), .B(n42570), .ZN(n42571) );
  XNOR2_X1 U45187 ( .A(n42571), .B(n45252), .ZN(n42572) );
  XNOR2_X1 U45188 ( .A(n42868), .B(n42572), .ZN(n42573) );
  XNOR2_X1 U45189 ( .A(n51100), .B(n42575), .ZN(n43710) );
  XNOR2_X1 U45190 ( .A(n42576), .B(n43143), .ZN(n42577) );
  XNOR2_X1 U45191 ( .A(n42580), .B(n42579), .ZN(n42581) );
  XNOR2_X1 U45192 ( .A(n43950), .B(n42581), .ZN(n42582) );
  XNOR2_X1 U45193 ( .A(n42582), .B(n43244), .ZN(n42583) );
  XNOR2_X1 U45194 ( .A(n42584), .B(n42583), .ZN(n42585) );
  XNOR2_X1 U45195 ( .A(n46118), .B(n42587), .ZN(n42588) );
  XNOR2_X1 U45196 ( .A(n42589), .B(n42588), .ZN(n42604) );
  NAND3_X1 U45197 ( .A1(n46360), .A2(n46274), .A3(n46342), .ZN(n42603) );
  XNOR2_X1 U45198 ( .A(n43755), .B(n45303), .ZN(n45455) );
  XNOR2_X1 U45199 ( .A(n43148), .B(n45455), .ZN(n42599) );
  XNOR2_X1 U45200 ( .A(n43206), .B(n43380), .ZN(n44143) );
  XNOR2_X1 U45201 ( .A(n42791), .B(n44143), .ZN(n42597) );
  XNOR2_X1 U45202 ( .A(n42591), .B(n43746), .ZN(n42593) );
  XNOR2_X1 U45203 ( .A(n42593), .B(n42592), .ZN(n42594) );
  XNOR2_X1 U45204 ( .A(n45305), .B(n42594), .ZN(n42595) );
  XNOR2_X1 U45205 ( .A(n44944), .B(n42595), .ZN(n42596) );
  XNOR2_X1 U45206 ( .A(n42597), .B(n42596), .ZN(n42598) );
  NAND2_X1 U45209 ( .A1(n45697), .A2(n46276), .ZN(n46352) );
  AND2_X1 U45211 ( .A1(n42603), .A2(n45232), .ZN(n42612) );
  NAND2_X1 U45212 ( .A1(n46267), .A2(n46356), .ZN(n45689) );
  INV_X1 U45213 ( .A(n45689), .ZN(n42608) );
  INV_X1 U45214 ( .A(n42604), .ZN(n46359) );
  NOR3_X1 U45216 ( .A1(n45231), .A2(n46353), .A3(n46356), .ZN(n42607) );
  INV_X1 U45217 ( .A(n42606), .ZN(n46358) );
  AOI22_X1 U45218 ( .A1(n42608), .A2(n52187), .B1(n42607), .B2(n46346), .ZN(
        n42611) );
  NAND3_X1 U45219 ( .A1(n46344), .A2(n46353), .A3(n46276), .ZN(n44761) );
  NAND2_X1 U45220 ( .A1(n46358), .A2(n46267), .ZN(n45688) );
  NOR2_X1 U45221 ( .A1(n46357), .A2(n46274), .ZN(n42609) );
  OR2_X1 U45222 ( .A1(n46267), .A2(n46276), .ZN(n44766) );
  NAND4_X1 U45223 ( .A1(n45688), .A2(n42609), .A3(n46277), .A4(n44766), .ZN(
        n42610) );
  NAND4_X1 U45224 ( .A1(n42612), .A2(n42611), .A3(n44761), .A4(n42610), .ZN(
        n42617) );
  OR2_X1 U45225 ( .A1(n45688), .A2(n46356), .ZN(n46265) );
  INV_X1 U45226 ( .A(n46357), .ZN(n42613) );
  NAND3_X1 U45227 ( .A1(n44766), .A2(n42613), .A3(n46269), .ZN(n42615) );
  NAND3_X1 U45228 ( .A1(n46355), .A2(n46274), .A3(n46357), .ZN(n42614) );
  OAI211_X1 U45229 ( .C1(n46265), .C2(n46342), .A(n42615), .B(n42614), .ZN(
        n42616) );
  INV_X1 U45230 ( .A(n42810), .ZN(n46951) );
  NAND2_X1 U45231 ( .A1(n48975), .A2(n46951), .ZN(n48955) );
  INV_X1 U45232 ( .A(n48955), .ZN(n42618) );
  XNOR2_X1 U45233 ( .A(n42620), .B(n42619), .ZN(n42621) );
  XNOR2_X1 U45234 ( .A(n44189), .B(n42621), .ZN(n42622) );
  INV_X1 U45236 ( .A(n42684), .ZN(n49201) );
  XNOR2_X1 U45237 ( .A(n4564), .B(n4431), .ZN(n42629) );
  XNOR2_X1 U45238 ( .A(n4565), .B(n4587), .ZN(n42628) );
  XNOR2_X1 U45239 ( .A(n42629), .B(n42628), .ZN(n42631) );
  XNOR2_X1 U45240 ( .A(n42631), .B(n42630), .ZN(n42632) );
  XNOR2_X1 U45241 ( .A(n42633), .B(n42632), .ZN(n42634) );
  XNOR2_X1 U45242 ( .A(n43206), .B(n42634), .ZN(n42635) );
  XNOR2_X1 U45243 ( .A(n42822), .B(n42636), .ZN(n42637) );
  XNOR2_X1 U45244 ( .A(n42637), .B(n42788), .ZN(n42638) );
  XNOR2_X1 U45245 ( .A(n516), .B(n43149), .ZN(n44571) );
  XNOR2_X1 U45247 ( .A(n42640), .B(n51100), .ZN(n42641) );
  XNOR2_X1 U45248 ( .A(n2228), .B(n42641), .ZN(n42642) );
  XNOR2_X1 U45249 ( .A(n44318), .B(n42642), .ZN(n44532) );
  XNOR2_X1 U45250 ( .A(n42643), .B(n43954), .ZN(n42644) );
  XNOR2_X1 U45251 ( .A(n40814), .B(n42644), .ZN(n42645) );
  INV_X1 U45252 ( .A(n43303), .ZN(n42654) );
  XNOR2_X1 U45253 ( .A(n42646), .B(n49867), .ZN(n42648) );
  XNOR2_X1 U45254 ( .A(n42648), .B(n42647), .ZN(n42649) );
  XNOR2_X1 U45255 ( .A(n44314), .B(n42649), .ZN(n42651) );
  XNOR2_X1 U45256 ( .A(n42651), .B(n42650), .ZN(n42652) );
  XNOR2_X1 U45257 ( .A(n42652), .B(n51390), .ZN(n42653) );
  XNOR2_X1 U45258 ( .A(n42654), .B(n42653), .ZN(n42655) );
  INV_X1 U45259 ( .A(n42685), .ZN(n49198) );
  XNOR2_X1 U45260 ( .A(n42657), .B(n42656), .ZN(n42658) );
  XNOR2_X1 U45261 ( .A(n44904), .B(n42658), .ZN(n42660) );
  XNOR2_X1 U45262 ( .A(n44296), .B(n42660), .ZN(n42661) );
  XNOR2_X1 U45263 ( .A(n42661), .B(n51333), .ZN(n42665) );
  XNOR2_X1 U45264 ( .A(n51509), .B(n42663), .ZN(n42664) );
  XNOR2_X1 U45265 ( .A(n43219), .B(n42668), .ZN(n42669) );
  XNOR2_X1 U45266 ( .A(n42669), .B(n42863), .ZN(n42671) );
  XNOR2_X1 U45267 ( .A(n42670), .B(n42671), .ZN(n42672) );
  XNOR2_X1 U45268 ( .A(n43218), .B(n42672), .ZN(n44518) );
  XNOR2_X1 U45269 ( .A(n42673), .B(n44518), .ZN(n45966) );
  XNOR2_X1 U45270 ( .A(n42674), .B(n47679), .ZN(n42675) );
  XNOR2_X1 U45271 ( .A(n42676), .B(n42675), .ZN(n42677) );
  XNOR2_X1 U45272 ( .A(n43106), .B(n42677), .ZN(n42678) );
  XNOR2_X1 U45273 ( .A(n45325), .B(n42678), .ZN(n42679) );
  XNOR2_X1 U45274 ( .A(n44479), .B(n42679), .ZN(n42681) );
  XNOR2_X1 U45275 ( .A(n42681), .B(n42680), .ZN(n42683) );
  OAI21_X1 U45276 ( .B1(n46231), .B2(n45970), .A(n49216), .ZN(n49205) );
  XNOR2_X1 U45277 ( .A(n42686), .B(n4855), .ZN(n42687) );
  XNOR2_X1 U45278 ( .A(n42688), .B(n42687), .ZN(n42690) );
  XNOR2_X1 U45279 ( .A(n42690), .B(n42689), .ZN(n42691) );
  XNOR2_X1 U45280 ( .A(n43357), .B(n42691), .ZN(n42692) );
  XNOR2_X1 U45281 ( .A(n42693), .B(n42692), .ZN(n42695) );
  XNOR2_X1 U45282 ( .A(n44176), .B(n46137), .ZN(n42694) );
  XNOR2_X1 U45283 ( .A(n42694), .B(n43113), .ZN(n43044) );
  XNOR2_X1 U45284 ( .A(n42695), .B(n43044), .ZN(n42697) );
  XNOR2_X1 U45285 ( .A(n43937), .B(n42697), .ZN(n42699) );
  OAI21_X1 U45286 ( .B1(n49207), .B2(n44752), .A(n49199), .ZN(n42702) );
  NOR2_X1 U45287 ( .A1(n52105), .A2(n46232), .ZN(n42700) );
  INV_X1 U45288 ( .A(n45966), .ZN(n42703) );
  INV_X1 U45289 ( .A(n52106), .ZN(n42701) );
  NAND3_X1 U45290 ( .A1(n42701), .A2(n46226), .A3(n45970), .ZN(n46220) );
  OR2_X1 U45291 ( .A1(n49199), .A2(n45967), .ZN(n46210) );
  OAI21_X1 U45292 ( .B1(n46228), .B2(n49197), .A(n45970), .ZN(n42704) );
  NOR2_X1 U45293 ( .A1(n46210), .A2(n42704), .ZN(n42707) );
  NAND2_X1 U45294 ( .A1(n44752), .A2(n45966), .ZN(n46214) );
  INV_X1 U45295 ( .A(n46214), .ZN(n46227) );
  OAI21_X1 U45296 ( .B1(n46227), .B2(n52106), .A(n49209), .ZN(n42706) );
  INV_X1 U45297 ( .A(n46231), .ZN(n42705) );
  MUX2_X1 U45298 ( .A(n42707), .B(n42706), .S(n42705), .Z(n42708) );
  OR2_X2 U45299 ( .A1(n42709), .A2(n42708), .ZN(n47477) );
  INV_X1 U45300 ( .A(n44960), .ZN(n43094) );
  XNOR2_X1 U45301 ( .A(n43068), .B(n43094), .ZN(n42888) );
  XNOR2_X1 U45302 ( .A(n42711), .B(n42710), .ZN(n42713) );
  XNOR2_X1 U45303 ( .A(n42713), .B(n42712), .ZN(n42714) );
  XNOR2_X1 U45304 ( .A(n42715), .B(n42714), .ZN(n42716) );
  XNOR2_X1 U45305 ( .A(n42717), .B(n42716), .ZN(n42718) );
  XNOR2_X1 U45306 ( .A(n44156), .B(n4526), .ZN(n45328) );
  XNOR2_X1 U45307 ( .A(n42718), .B(n45328), .ZN(n42719) );
  XNOR2_X1 U45308 ( .A(n45067), .B(n43070), .ZN(n43995) );
  XNOR2_X1 U45309 ( .A(n42719), .B(n43995), .ZN(n42720) );
  XNOR2_X1 U45310 ( .A(n43139), .B(n43950), .ZN(n43716) );
  XNOR2_X1 U45311 ( .A(n42722), .B(n42721), .ZN(n42725) );
  INV_X1 U45312 ( .A(n42723), .ZN(n42724) );
  XNOR2_X1 U45313 ( .A(n42725), .B(n42724), .ZN(n42726) );
  XNOR2_X1 U45314 ( .A(n51101), .B(n42726), .ZN(n42727) );
  XNOR2_X1 U45315 ( .A(n43716), .B(n42727), .ZN(n42728) );
  XNOR2_X1 U45316 ( .A(n42729), .B(n43027), .ZN(n42731) );
  XNOR2_X1 U45317 ( .A(n42730), .B(n46112), .ZN(n43300) );
  XNOR2_X1 U45318 ( .A(n42731), .B(n43300), .ZN(n42732) );
  XNOR2_X1 U45319 ( .A(n42732), .B(n42733), .ZN(n42735) );
  XNOR2_X2 U45320 ( .A(n42734), .B(n42735), .ZN(n45661) );
  AND2_X1 U45321 ( .A1(n46498), .A2(n45661), .ZN(n42767) );
  INV_X1 U45322 ( .A(n43691), .ZN(n42736) );
  XNOR2_X1 U45323 ( .A(n43696), .B(n42736), .ZN(n42737) );
  XNOR2_X1 U45324 ( .A(n42863), .B(n42737), .ZN(n42738) );
  XNOR2_X1 U45325 ( .A(n43218), .B(n42738), .ZN(n43983) );
  XNOR2_X1 U45326 ( .A(n42739), .B(n45389), .ZN(n43297) );
  XNOR2_X1 U45327 ( .A(n44510), .B(n42740), .ZN(n45383) );
  XNOR2_X1 U45328 ( .A(n42742), .B(n42741), .ZN(n42743) );
  XNOR2_X1 U45329 ( .A(n43123), .B(n42743), .ZN(n42744) );
  XNOR2_X1 U45330 ( .A(n45383), .B(n42744), .ZN(n42745) );
  AOI21_X1 U45333 ( .B1(n42751), .B2(n42750), .A(n42749), .ZN(n42752) );
  OR2_X1 U45334 ( .A1(n42753), .A2(n42752), .ZN(n45365) );
  XNOR2_X1 U45335 ( .A(n43354), .B(n45365), .ZN(n42760) );
  XNOR2_X1 U45336 ( .A(n42755), .B(n42754), .ZN(n42756) );
  XNOR2_X1 U45337 ( .A(n42757), .B(n42756), .ZN(n42758) );
  XNOR2_X1 U45338 ( .A(n42760), .B(n42759), .ZN(n42761) );
  XNOR2_X1 U45339 ( .A(n42762), .B(n42761), .ZN(n42763) );
  XNOR2_X1 U45340 ( .A(n51420), .B(n42764), .ZN(n42765) );
  XNOR2_X1 U45341 ( .A(n43360), .B(n42765), .ZN(n42766) );
  OAI22_X1 U45342 ( .A1(n42767), .A2(n46380), .B1(n46493), .B2(n46487), .ZN(
        n42795) );
  XNOR2_X1 U45343 ( .A(n44535), .B(n46059), .ZN(n45298) );
  XOR2_X1 U45344 ( .A(n4325), .B(n42769), .Z(n42770) );
  XNOR2_X1 U45345 ( .A(n42771), .B(n42770), .ZN(n42772) );
  XNOR2_X1 U45346 ( .A(n42773), .B(n42772), .ZN(n42774) );
  XNOR2_X1 U45347 ( .A(n44190), .B(n42774), .ZN(n42775) );
  XNOR2_X1 U45348 ( .A(n45298), .B(n42775), .ZN(n42776) );
  XNOR2_X1 U45349 ( .A(n42777), .B(n44553), .ZN(n42797) );
  XNOR2_X1 U45350 ( .A(n44559), .B(n44562), .ZN(n42779) );
  INV_X1 U45351 ( .A(n44944), .ZN(n44131) );
  XNOR2_X1 U45352 ( .A(n42779), .B(n44131), .ZN(n42785) );
  XNOR2_X1 U45353 ( .A(n42781), .B(n42780), .ZN(n42782) );
  XNOR2_X1 U45354 ( .A(n43547), .B(n42782), .ZN(n42783) );
  XNOR2_X1 U45355 ( .A(n42783), .B(n43380), .ZN(n42784) );
  XNOR2_X1 U45356 ( .A(n42785), .B(n42784), .ZN(n42790) );
  XNOR2_X1 U45357 ( .A(n42786), .B(n44347), .ZN(n42787) );
  XNOR2_X1 U45358 ( .A(n42788), .B(n42787), .ZN(n42789) );
  XNOR2_X1 U45359 ( .A(n42789), .B(n42790), .ZN(n42793) );
  XNOR2_X1 U45360 ( .A(n42791), .B(n42938), .ZN(n43758) );
  XNOR2_X1 U45361 ( .A(n43758), .B(n43149), .ZN(n42792) );
  XNOR2_X2 U45362 ( .A(n42793), .B(n42792), .ZN(n46395) );
  INV_X1 U45363 ( .A(n46392), .ZN(n46385) );
  NAND2_X1 U45364 ( .A1(n46501), .A2(n46488), .ZN(n42794) );
  AOI22_X1 U45365 ( .A1(n42795), .A2(n46385), .B1(n46505), .B2(n42794), .ZN(
        n42803) );
  NAND2_X1 U45366 ( .A1(n46503), .A2(n45661), .ZN(n42798) );
  INV_X1 U45367 ( .A(n46498), .ZN(n45219) );
  NAND2_X1 U45368 ( .A1(n42798), .A2(n45219), .ZN(n42800) );
  INV_X1 U45370 ( .A(n46395), .ZN(n46491) );
  AND2_X1 U45373 ( .A1(n46488), .A2(n46491), .ZN(n46404) );
  NAND2_X1 U45374 ( .A1(n46404), .A2(n46501), .ZN(n45660) );
  INV_X1 U45375 ( .A(n46494), .ZN(n42801) );
  OR2_X1 U45376 ( .A1(n45660), .A2(n42801), .ZN(n42802) );
  INV_X1 U45377 ( .A(n48930), .ZN(n42804) );
  AND2_X1 U45378 ( .A1(n46951), .A2(n47477), .ZN(n47481) );
  NOR2_X1 U45379 ( .A1(n47477), .A2(n48973), .ZN(n48960) );
  NAND2_X1 U45380 ( .A1(n42805), .A2(n48960), .ZN(n48981) );
  NOR2_X1 U45381 ( .A1(n48974), .A2(n48935), .ZN(n47479) );
  NAND2_X1 U45382 ( .A1(n47479), .A2(n48976), .ZN(n47485) );
  INV_X1 U45383 ( .A(n48976), .ZN(n42808) );
  NAND3_X1 U45384 ( .A1(n42808), .A2(n48974), .A3(n48935), .ZN(n42809) );
  NOR2_X1 U45385 ( .A1(n48958), .A2(n48973), .ZN(n46957) );
  NAND2_X1 U45386 ( .A1(n46957), .A2(n51478), .ZN(n42812) );
  NAND2_X1 U45387 ( .A1(n42810), .A2(n47477), .ZN(n48950) );
  OR2_X1 U45388 ( .A1(n48950), .A2(n51478), .ZN(n42811) );
  MUX2_X1 U45389 ( .A(n42812), .B(n42811), .S(n51510), .Z(n42814) );
  NOR2_X1 U45390 ( .A1(n48950), .A2(n51510), .ZN(n48972) );
  NAND2_X1 U45391 ( .A1(n48935), .A2(n48957), .ZN(n48941) );
  INV_X1 U45392 ( .A(n48941), .ZN(n48951) );
  INV_X1 U45393 ( .A(n48952), .ZN(n47484) );
  AOI22_X1 U45394 ( .A1(n48972), .A2(n48951), .B1(n48974), .B2(n47484), .ZN(
        n42813) );
  INV_X1 U45395 ( .A(n4874), .ZN(n42815) );
  XNOR2_X1 U45396 ( .A(n45114), .B(n42816), .ZN(n42817) );
  XNOR2_X1 U45397 ( .A(n42817), .B(n51337), .ZN(n45451) );
  XNOR2_X1 U45398 ( .A(n45305), .B(n1224), .ZN(n42818) );
  XNOR2_X1 U45399 ( .A(n42818), .B(n45445), .ZN(n43872) );
  XNOR2_X1 U45400 ( .A(n43872), .B(n45451), .ZN(n42821) );
  INV_X1 U45401 ( .A(n4343), .ZN(n49817) );
  XNOR2_X1 U45402 ( .A(n45306), .B(n49817), .ZN(n42820) );
  XNOR2_X1 U45403 ( .A(n42820), .B(n42819), .ZN(n42943) );
  XNOR2_X1 U45404 ( .A(n42821), .B(n42943), .ZN(n42829) );
  XNOR2_X1 U45405 ( .A(n42822), .B(n43755), .ZN(n42941) );
  XNOR2_X1 U45406 ( .A(n42824), .B(n42823), .ZN(n42825) );
  XNOR2_X1 U45407 ( .A(n44130), .B(n42825), .ZN(n42826) );
  XNOR2_X1 U45408 ( .A(n42826), .B(n45116), .ZN(n42827) );
  XNOR2_X1 U45409 ( .A(n42941), .B(n42827), .ZN(n42828) );
  XNOR2_X1 U45410 ( .A(n42829), .B(n42828), .ZN(n42830) );
  XNOR2_X1 U45411 ( .A(n43658), .B(n45304), .ZN(n44949) );
  INV_X1 U45412 ( .A(n42883), .ZN(n49690) );
  XNOR2_X1 U45413 ( .A(n42831), .B(n4880), .ZN(n42832) );
  XNOR2_X1 U45414 ( .A(n42833), .B(n42832), .ZN(n42834) );
  XNOR2_X1 U45415 ( .A(n42835), .B(n42834), .ZN(n42836) );
  XNOR2_X1 U45416 ( .A(n43168), .B(n42836), .ZN(n42837) );
  XNOR2_X1 U45417 ( .A(n43522), .B(n42837), .ZN(n42840) );
  XNOR2_X1 U45418 ( .A(n51444), .B(n670), .ZN(n42839) );
  XNOR2_X1 U45419 ( .A(n42840), .B(n42839), .ZN(n42842) );
  INV_X1 U45420 ( .A(n42953), .ZN(n42841) );
  XNOR2_X1 U45421 ( .A(n42841), .B(n42842), .ZN(n42843) );
  XNOR2_X1 U45422 ( .A(n43642), .B(n42955), .ZN(n45136) );
  XNOR2_X1 U45423 ( .A(n44030), .B(n51099), .ZN(n43845) );
  XOR2_X1 U45424 ( .A(n42845), .B(n42844), .Z(n42847) );
  XNOR2_X1 U45425 ( .A(n42847), .B(n42846), .ZN(n42848) );
  XNOR2_X1 U45426 ( .A(n43139), .B(n42848), .ZN(n42849) );
  XNOR2_X1 U45427 ( .A(n43845), .B(n42849), .ZN(n42852) );
  XNOR2_X1 U45428 ( .A(n51431), .B(n44237), .ZN(n42851) );
  XNOR2_X1 U45429 ( .A(n42850), .B(n42851), .ZN(n43717) );
  XNOR2_X1 U45430 ( .A(n42852), .B(n43717), .ZN(n42854) );
  XNOR2_X1 U45431 ( .A(n42854), .B(n42853), .ZN(n42857) );
  XNOR2_X1 U45432 ( .A(n45416), .B(n43308), .ZN(n42855) );
  XNOR2_X1 U45433 ( .A(n44529), .B(n42855), .ZN(n42856) );
  INV_X1 U45434 ( .A(n49695), .ZN(n45921) );
  XNOR2_X1 U45435 ( .A(n43698), .B(n45389), .ZN(n42866) );
  XNOR2_X1 U45436 ( .A(n42859), .B(n42858), .ZN(n42860) );
  XNOR2_X1 U45437 ( .A(n42861), .B(n42860), .ZN(n42862) );
  XNOR2_X1 U45438 ( .A(n44904), .B(n42862), .ZN(n42864) );
  XNOR2_X1 U45439 ( .A(n42864), .B(n42863), .ZN(n42865) );
  XNOR2_X1 U45440 ( .A(n42866), .B(n42865), .ZN(n42867) );
  XNOR2_X1 U45441 ( .A(n42868), .B(n42867), .ZN(n42871) );
  XNOR2_X1 U45443 ( .A(n42870), .B(n43833), .ZN(n44903) );
  NAND2_X1 U45444 ( .A1(n45921), .A2(n49247), .ZN(n49686) );
  XNOR2_X1 U45445 ( .A(n46143), .B(n43609), .ZN(n42873) );
  XNOR2_X1 U45446 ( .A(n42873), .B(n45355), .ZN(n42874) );
  XNOR2_X1 U45447 ( .A(n42874), .B(n52085), .ZN(n43365) );
  XOR2_X1 U45448 ( .A(n45463), .B(n43739), .Z(n42875) );
  XNOR2_X1 U45449 ( .A(n42876), .B(n42875), .ZN(n42877) );
  XNOR2_X1 U45450 ( .A(n42877), .B(n43728), .ZN(n42878) );
  XNOR2_X1 U45451 ( .A(n50967), .B(n42878), .ZN(n42879) );
  INV_X1 U45452 ( .A(n42962), .ZN(n45468) );
  XNOR2_X1 U45453 ( .A(n42879), .B(n45468), .ZN(n42880) );
  XNOR2_X1 U45454 ( .A(n42880), .B(n43816), .ZN(n42881) );
  XNOR2_X1 U45455 ( .A(n43048), .B(n43725), .ZN(n43603) );
  XNOR2_X1 U45456 ( .A(n42881), .B(n43603), .ZN(n42882) );
  OR2_X1 U45457 ( .A1(n49686), .A2(n49231), .ZN(n42885) );
  AND2_X1 U45458 ( .A1(n49397), .A2(n51095), .ZN(n45913) );
  NAND2_X1 U45459 ( .A1(n45913), .A2(n43474), .ZN(n42884) );
  INV_X1 U45460 ( .A(n44743), .ZN(n45919) );
  MUX2_X1 U45461 ( .A(n45919), .B(n49254), .S(n49397), .Z(n42902) );
  XNOR2_X1 U45462 ( .A(n42888), .B(n42887), .ZN(n42901) );
  XNOR2_X1 U45463 ( .A(n52125), .B(n43890), .ZN(n45332) );
  XNOR2_X1 U45464 ( .A(n42889), .B(n49109), .ZN(n42890) );
  XNOR2_X1 U45465 ( .A(n42891), .B(n42890), .ZN(n42892) );
  XNOR2_X1 U45466 ( .A(n42893), .B(n42892), .ZN(n42894) );
  XNOR2_X1 U45467 ( .A(n43596), .B(n42894), .ZN(n42895) );
  XNOR2_X1 U45468 ( .A(n45332), .B(n42895), .ZN(n42897) );
  XNOR2_X1 U45469 ( .A(n42897), .B(n42896), .ZN(n42899) );
  XNOR2_X1 U45470 ( .A(n44153), .B(n43102), .ZN(n45487) );
  XOR2_X1 U45471 ( .A(n45487), .B(n44394), .Z(n42898) );
  XNOR2_X1 U45472 ( .A(n42899), .B(n42898), .ZN(n42900) );
  INV_X1 U45473 ( .A(n588), .ZN(n49230) );
  NOR2_X1 U45474 ( .A1(n49248), .A2(n49230), .ZN(n42904) );
  OAI21_X1 U45475 ( .B1(n43474), .B2(n49684), .A(n49686), .ZN(n42903) );
  OAI22_X1 U45476 ( .A1(n42904), .A2(n42903), .B1(n49242), .B2(n49696), .ZN(
        n42905) );
  XNOR2_X1 U45477 ( .A(n42907), .B(n43000), .ZN(n42912) );
  XNOR2_X1 U45478 ( .A(n42909), .B(n42908), .ZN(n42910) );
  XNOR2_X1 U45479 ( .A(n44017), .B(n42910), .ZN(n42911) );
  XNOR2_X1 U45480 ( .A(n42911), .B(n42912), .ZN(n42913) );
  XNOR2_X1 U45481 ( .A(n42913), .B(n43291), .ZN(n42914) );
  XNOR2_X1 U45482 ( .A(n44903), .B(n42914), .ZN(n42915) );
  XNOR2_X1 U45483 ( .A(n42906), .B(n42915), .ZN(n42917) );
  XNOR2_X1 U45484 ( .A(n46112), .B(n46113), .ZN(n44520) );
  XNOR2_X1 U45485 ( .A(n44520), .B(n44893), .ZN(n43859) );
  XNOR2_X1 U45486 ( .A(n42918), .B(n47802), .ZN(n42919) );
  XNOR2_X1 U45487 ( .A(n42920), .B(n42919), .ZN(n42921) );
  XNOR2_X1 U45488 ( .A(n46126), .B(n42921), .ZN(n42922) );
  XNOR2_X1 U45489 ( .A(n44237), .B(n42922), .ZN(n42924) );
  XNOR2_X1 U45490 ( .A(n42924), .B(n42923), .ZN(n42925) );
  XNOR2_X1 U45491 ( .A(n45269), .B(n42925), .ZN(n42926) );
  XNOR2_X1 U45492 ( .A(n43859), .B(n42926), .ZN(n42927) );
  XNOR2_X1 U45493 ( .A(n43575), .B(n42928), .ZN(n42932) );
  INV_X1 U45494 ( .A(n4649), .ZN(n47627) );
  XNOR2_X1 U45495 ( .A(n45408), .B(n47627), .ZN(n42930) );
  XNOR2_X1 U45496 ( .A(n42930), .B(n52096), .ZN(n42931) );
  XNOR2_X1 U45497 ( .A(n42932), .B(n42931), .ZN(n43250) );
  XNOR2_X1 U45498 ( .A(n4666), .B(n4793), .ZN(n42933) );
  XNOR2_X1 U45499 ( .A(n42934), .B(n42933), .ZN(n42935) );
  XNOR2_X1 U45500 ( .A(n42936), .B(n42935), .ZN(n42937) );
  XNOR2_X1 U45501 ( .A(n42938), .B(n42937), .ZN(n42939) );
  INV_X1 U45502 ( .A(n50987), .ZN(n42940) );
  XNOR2_X1 U45503 ( .A(n44130), .B(n42940), .ZN(n46052) );
  XNOR2_X1 U45504 ( .A(n45454), .B(n42943), .ZN(n42944) );
  XNOR2_X1 U45505 ( .A(n42945), .B(n42944), .ZN(n43464) );
  XNOR2_X1 U45506 ( .A(n42947), .B(n42946), .ZN(n42948) );
  XNOR2_X1 U45507 ( .A(n43781), .B(n42948), .ZN(n42950) );
  XNOR2_X1 U45508 ( .A(n42950), .B(n42949), .ZN(n42951) );
  XNOR2_X1 U45509 ( .A(n44056), .B(n42951), .ZN(n42952) );
  XNOR2_X1 U45510 ( .A(n42953), .B(n42952), .ZN(n42956) );
  INV_X1 U45511 ( .A(n45995), .ZN(n43460) );
  NAND2_X1 U45512 ( .A1(n42957), .A2(n49191), .ZN(n49188) );
  XNOR2_X1 U45513 ( .A(n42959), .B(n42958), .ZN(n42960) );
  XNOR2_X1 U45514 ( .A(n42961), .B(n42960), .ZN(n42963) );
  XNOR2_X1 U45515 ( .A(n42962), .B(n42963), .ZN(n42964) );
  XNOR2_X1 U45516 ( .A(n44170), .B(n42965), .ZN(n42967) );
  XNOR2_X1 U45517 ( .A(n51096), .B(n44182), .ZN(n42966) );
  XNOR2_X1 U45518 ( .A(n42966), .B(n51368), .ZN(n45363) );
  XNOR2_X1 U45519 ( .A(n42967), .B(n45363), .ZN(n42970) );
  XNOR2_X1 U45520 ( .A(n44979), .B(n52085), .ZN(n42968) );
  XNOR2_X1 U45521 ( .A(n43742), .B(n42968), .ZN(n46158) );
  INV_X1 U45522 ( .A(n46158), .ZN(n42969) );
  NAND2_X1 U45523 ( .A1(n49707), .A2(n49719), .ZN(n45989) );
  INV_X1 U45524 ( .A(n49725), .ZN(n43467) );
  AOI21_X1 U45525 ( .B1(n49188), .B2(n45989), .A(n43467), .ZN(n42988) );
  NAND2_X1 U45526 ( .A1(n43467), .A2(n49711), .ZN(n43470) );
  NAND3_X1 U45527 ( .A1(n43462), .A2(n49719), .A3(n43464), .ZN(n42972) );
  NOR2_X1 U45528 ( .A1(n43464), .A2(n49721), .ZN(n49184) );
  INV_X1 U45529 ( .A(n42971), .ZN(n49710) );
  XNOR2_X1 U45530 ( .A(n42973), .B(n4585), .ZN(n42974) );
  XNOR2_X1 U45531 ( .A(n42975), .B(n42974), .ZN(n42976) );
  XNOR2_X1 U45532 ( .A(n52125), .B(n42976), .ZN(n42977) );
  XNOR2_X1 U45533 ( .A(n42977), .B(n46079), .ZN(n42978) );
  XNOR2_X1 U45534 ( .A(n44960), .B(n42978), .ZN(n42984) );
  XNOR2_X1 U45535 ( .A(n42979), .B(n43079), .ZN(n42983) );
  XNOR2_X1 U45536 ( .A(n42980), .B(n44963), .ZN(n42981) );
  XNOR2_X1 U45537 ( .A(n42983), .B(n42982), .ZN(n43261) );
  XNOR2_X1 U45538 ( .A(n42984), .B(n43261), .ZN(n42987) );
  XNOR2_X1 U45539 ( .A(n42985), .B(n44479), .ZN(n42986) );
  XNOR2_X1 U45540 ( .A(n42987), .B(n42986), .ZN(n45909) );
  INV_X1 U45541 ( .A(n45909), .ZN(n49714) );
  OR2_X1 U45542 ( .A1(n43464), .A2(n45995), .ZN(n45999) );
  NAND2_X1 U45543 ( .A1(n51295), .A2(n42990), .ZN(n45907) );
  NOR2_X1 U45544 ( .A1(n45999), .A2(n45907), .ZN(n45994) );
  AND2_X1 U45545 ( .A1(n45909), .A2(n49719), .ZN(n49189) );
  AND2_X1 U45546 ( .A1(n49189), .A2(n42990), .ZN(n42989) );
  NOR2_X1 U45547 ( .A1(n45994), .A2(n42989), .ZN(n42994) );
  NAND2_X1 U45548 ( .A1(n49191), .A2(n42990), .ZN(n45897) );
  NAND3_X1 U45549 ( .A1(n45897), .A2(n45987), .A3(n45989), .ZN(n42991) );
  NAND2_X1 U45550 ( .A1(n42991), .A2(n45910), .ZN(n42993) );
  XNOR2_X1 U45551 ( .A(n45393), .B(n43698), .ZN(n43004) );
  XNOR2_X1 U45552 ( .A(n42996), .B(n42995), .ZN(n42997) );
  XNOR2_X1 U45553 ( .A(n42998), .B(n42997), .ZN(n42999) );
  XNOR2_X1 U45554 ( .A(n44017), .B(n42999), .ZN(n43001) );
  XNOR2_X1 U45555 ( .A(n51406), .B(n43001), .ZN(n43002) );
  XNOR2_X1 U45556 ( .A(n44207), .B(n43002), .ZN(n43003) );
  XNOR2_X1 U45557 ( .A(n43003), .B(n43004), .ZN(n43005) );
  XNOR2_X1 U45558 ( .A(n46108), .B(n43005), .ZN(n43007) );
  XNOR2_X1 U45559 ( .A(n43660), .B(n43006), .ZN(n44917) );
  XNOR2_X1 U45560 ( .A(n43007), .B(n44917), .ZN(n50293) );
  INV_X1 U45561 ( .A(n50293), .ZN(n49940) );
  XNOR2_X1 U45562 ( .A(n44561), .B(n44042), .ZN(n43008) );
  XNOR2_X1 U45563 ( .A(n44146), .B(n43008), .ZN(n43009) );
  XNOR2_X1 U45564 ( .A(n43009), .B(n43751), .ZN(n43213) );
  XNOR2_X1 U45565 ( .A(n43928), .B(n44134), .ZN(n43011) );
  XNOR2_X1 U45566 ( .A(n43155), .B(n4501), .ZN(n43010) );
  XNOR2_X1 U45567 ( .A(n43011), .B(n43010), .ZN(n43870) );
  XNOR2_X1 U45568 ( .A(n43012), .B(n43870), .ZN(n43013) );
  XNOR2_X1 U45569 ( .A(n43213), .B(n43013), .ZN(n43026) );
  XNOR2_X1 U45570 ( .A(n43014), .B(n4666), .ZN(n43015) );
  XNOR2_X1 U45571 ( .A(n52171), .B(n43015), .ZN(n43016) );
  XNOR2_X1 U45572 ( .A(n45099), .B(n43016), .ZN(n44149) );
  XNOR2_X1 U45573 ( .A(n50987), .B(n44046), .ZN(n43017) );
  XNOR2_X1 U45574 ( .A(n43017), .B(n44130), .ZN(n43759) );
  XNOR2_X1 U45575 ( .A(n43019), .B(n43018), .ZN(n43021) );
  XNOR2_X1 U45576 ( .A(n43021), .B(n43020), .ZN(n43022) );
  XNOR2_X1 U45577 ( .A(n43157), .B(n43022), .ZN(n43023) );
  XNOR2_X1 U45578 ( .A(n43759), .B(n43023), .ZN(n43024) );
  XNOR2_X1 U45579 ( .A(n44149), .B(n43024), .ZN(n43025) );
  NOR2_X1 U45580 ( .A1(n49940), .A2(n50294), .ZN(n49636) );
  XNOR2_X1 U45581 ( .A(n43028), .B(n45059), .ZN(n43960) );
  XNOR2_X1 U45582 ( .A(n43960), .B(n43029), .ZN(n43038) );
  XNOR2_X1 U45583 ( .A(n43954), .B(n47802), .ZN(n43243) );
  XNOR2_X1 U45584 ( .A(n43030), .B(n43849), .ZN(n43031) );
  XNOR2_X1 U45585 ( .A(n43032), .B(n43031), .ZN(n43033) );
  XNOR2_X1 U45586 ( .A(n43236), .B(n43033), .ZN(n43034) );
  XNOR2_X1 U45587 ( .A(n43243), .B(n43034), .ZN(n43035) );
  XNOR2_X1 U45588 ( .A(n44240), .B(n46112), .ZN(n44307) );
  XNOR2_X1 U45589 ( .A(n43035), .B(n44307), .ZN(n43036) );
  XNOR2_X1 U45590 ( .A(n51390), .B(n43143), .ZN(n46133) );
  XNOR2_X1 U45591 ( .A(n43036), .B(n46133), .ZN(n43037) );
  XNOR2_X1 U45592 ( .A(n43038), .B(n43037), .ZN(n43089) );
  XNOR2_X1 U45594 ( .A(n43943), .B(n4836), .ZN(n44971) );
  XNOR2_X1 U45595 ( .A(n51420), .B(n52085), .ZN(n43509) );
  XNOR2_X1 U45596 ( .A(n43509), .B(n43039), .ZN(n43047) );
  XNOR2_X1 U45597 ( .A(n43041), .B(n43040), .ZN(n43042) );
  XNOR2_X1 U45598 ( .A(n44979), .B(n43042), .ZN(n43043) );
  XNOR2_X1 U45599 ( .A(n43043), .B(n45468), .ZN(n43045) );
  XNOR2_X1 U45600 ( .A(n43045), .B(n43044), .ZN(n43046) );
  XNOR2_X1 U45601 ( .A(n43047), .B(n43046), .ZN(n43049) );
  AOI21_X1 U45602 ( .B1(n49636), .B2(n49946), .A(n50287), .ZN(n43088) );
  XNOR2_X1 U45603 ( .A(n43050), .B(n51409), .ZN(n43195) );
  XNOR2_X1 U45604 ( .A(n44189), .B(n46058), .ZN(n43051) );
  XNOR2_X1 U45605 ( .A(n43051), .B(n52222), .ZN(n43052) );
  XNOR2_X1 U45606 ( .A(n43195), .B(n43052), .ZN(n43067) );
  XNOR2_X1 U45607 ( .A(n43053), .B(n4931), .ZN(n43055) );
  XNOR2_X1 U45608 ( .A(n43055), .B(n43054), .ZN(n43056) );
  XNOR2_X1 U45609 ( .A(n43057), .B(n43056), .ZN(n43058) );
  XNOR2_X1 U45610 ( .A(n43168), .B(n43058), .ZN(n43060) );
  XNOR2_X1 U45611 ( .A(n43196), .B(n43060), .ZN(n43061) );
  XNOR2_X1 U45612 ( .A(n43062), .B(n43061), .ZN(n43065) );
  XNOR2_X1 U45613 ( .A(n52130), .B(n43064), .ZN(n44929) );
  XNOR2_X1 U45614 ( .A(n44929), .B(n43065), .ZN(n43066) );
  OAI21_X1 U45615 ( .B1(n51504), .B2(n51313), .A(n46035), .ZN(n43087) );
  XNOR2_X1 U45616 ( .A(n43069), .B(n43890), .ZN(n44392) );
  XNOR2_X1 U45617 ( .A(n43068), .B(n44392), .ZN(n43072) );
  XNOR2_X1 U45618 ( .A(n43070), .B(n44154), .ZN(n43071) );
  XNOR2_X1 U45619 ( .A(n43071), .B(n52135), .ZN(n44480) );
  XNOR2_X1 U45620 ( .A(n44480), .B(n43072), .ZN(n43085) );
  XNOR2_X1 U45621 ( .A(n43074), .B(n43073), .ZN(n43075) );
  XNOR2_X1 U45622 ( .A(n43076), .B(n43075), .ZN(n43077) );
  XNOR2_X1 U45623 ( .A(n44962), .B(n43077), .ZN(n43078) );
  XNOR2_X1 U45624 ( .A(n44391), .B(n43078), .ZN(n43081) );
  XNOR2_X1 U45625 ( .A(n43081), .B(n43080), .ZN(n43083) );
  XNOR2_X1 U45626 ( .A(n46079), .B(n46090), .ZN(n43082) );
  XNOR2_X1 U45627 ( .A(n43083), .B(n43082), .ZN(n43084) );
  AOI21_X1 U45629 ( .B1(n50299), .B2(n49946), .A(n51691), .ZN(n43086) );
  NAND2_X1 U45630 ( .A1(n49940), .A2(n43089), .ZN(n47307) );
  NAND2_X1 U45631 ( .A1(n50296), .A2(n51691), .ZN(n49945) );
  INV_X1 U45632 ( .A(n49945), .ZN(n49614) );
  INV_X1 U45633 ( .A(n46035), .ZN(n43090) );
  OAI211_X1 U45634 ( .C1(n47307), .C2(n49614), .A(n51504), .B(n43090), .ZN(
        n43093) );
  NOR2_X1 U45635 ( .A1(n49945), .A2(n51300), .ZN(n46033) );
  INV_X1 U45636 ( .A(n50294), .ZN(n49939) );
  INV_X1 U45638 ( .A(n50305), .ZN(n43091) );
  NAND2_X1 U45639 ( .A1(n49940), .A2(n49946), .ZN(n50297) );
  NAND3_X1 U45640 ( .A1(n50289), .A2(n49614), .A3(n50297), .ZN(n43092) );
  NOR2_X1 U45641 ( .A1(n51088), .A2(n49605), .ZN(n49573) );
  NOR2_X1 U45642 ( .A1(n49607), .A2(n49579), .ZN(n43188) );
  XNOR2_X1 U45643 ( .A(n43504), .B(n43094), .ZN(n43100) );
  XNOR2_X1 U45644 ( .A(n43096), .B(n43095), .ZN(n43097) );
  XNOR2_X1 U45645 ( .A(n43098), .B(n43097), .ZN(n43099) );
  XNOR2_X1 U45646 ( .A(n43100), .B(n43099), .ZN(n43101) );
  XNOR2_X1 U45647 ( .A(n44480), .B(n43101), .ZN(n43107) );
  XNOR2_X1 U45648 ( .A(n51294), .B(n43102), .ZN(n43103) );
  XNOR2_X1 U45649 ( .A(n43103), .B(n44153), .ZN(n43104) );
  XNOR2_X1 U45650 ( .A(n43320), .B(n44079), .ZN(n43996) );
  XNOR2_X1 U45651 ( .A(n43109), .B(n43108), .ZN(n43110) );
  XNOR2_X1 U45652 ( .A(n43112), .B(n51096), .ZN(n43115) );
  XNOR2_X1 U45653 ( .A(n46143), .B(n43113), .ZN(n43114) );
  INV_X1 U45654 ( .A(n4529), .ZN(n50759) );
  XNOR2_X1 U45655 ( .A(n46137), .B(n50759), .ZN(n43116) );
  XNOR2_X1 U45656 ( .A(n43116), .B(n45365), .ZN(n43117) );
  XNOR2_X1 U45657 ( .A(n43352), .B(n43117), .ZN(n43119) );
  XNOR2_X1 U45658 ( .A(n43119), .B(n43118), .ZN(n43259) );
  XNOR2_X1 U45659 ( .A(n43121), .B(n43120), .ZN(n43122) );
  XNOR2_X1 U45660 ( .A(n43123), .B(n43122), .ZN(n43124) );
  XNOR2_X1 U45661 ( .A(n44301), .B(n45385), .ZN(n43551) );
  XNOR2_X1 U45662 ( .A(n43125), .B(n43551), .ZN(n43126) );
  XNOR2_X1 U45663 ( .A(n44291), .B(n43126), .ZN(n43129) );
  XNOR2_X1 U45664 ( .A(n43218), .B(n43127), .ZN(n43128) );
  XNOR2_X1 U45665 ( .A(n43129), .B(n43128), .ZN(n43147) );
  XNOR2_X1 U45666 ( .A(n43131), .B(n43130), .ZN(n43567) );
  XNOR2_X1 U45667 ( .A(n52204), .B(n43567), .ZN(n43134) );
  XNOR2_X1 U45668 ( .A(n45415), .B(n43132), .ZN(n43133) );
  XNOR2_X1 U45669 ( .A(n43133), .B(n43134), .ZN(n43135) );
  XNOR2_X1 U45670 ( .A(n43135), .B(n44320), .ZN(n43146) );
  XNOR2_X1 U45671 ( .A(n43137), .B(n43136), .ZN(n43138) );
  XNOR2_X1 U45672 ( .A(n43139), .B(n43138), .ZN(n43140) );
  XNOR2_X1 U45673 ( .A(n44240), .B(n43140), .ZN(n43142) );
  XNOR2_X1 U45674 ( .A(n43142), .B(n43141), .ZN(n43144) );
  XNOR2_X1 U45675 ( .A(n43144), .B(n45418), .ZN(n43145) );
  XNOR2_X1 U45676 ( .A(n43146), .B(n43145), .ZN(n43184) );
  INV_X1 U45677 ( .A(n43184), .ZN(n49978) );
  XNOR2_X1 U45678 ( .A(n43929), .B(n45116), .ZN(n46054) );
  XNOR2_X1 U45679 ( .A(n43148), .B(n46054), .ZN(n43379) );
  XNOR2_X1 U45680 ( .A(n43151), .B(n43150), .ZN(n43152) );
  XNOR2_X1 U45681 ( .A(n43153), .B(n43152), .ZN(n43154) );
  XNOR2_X1 U45682 ( .A(n43155), .B(n43154), .ZN(n43156) );
  XNOR2_X1 U45683 ( .A(n44561), .B(n43156), .ZN(n43158) );
  XNOR2_X1 U45684 ( .A(n43157), .B(n44937), .ZN(n43536) );
  XNOR2_X1 U45685 ( .A(n43158), .B(n43536), .ZN(n43159) );
  BUF_X2 U45686 ( .A(n43181), .Z(n49627) );
  XNOR2_X1 U45687 ( .A(n4931), .B(n4880), .ZN(n43163) );
  XNOR2_X1 U45688 ( .A(n43164), .B(n43163), .ZN(n43165) );
  XNOR2_X1 U45689 ( .A(n43166), .B(n43165), .ZN(n43167) );
  XNOR2_X1 U45690 ( .A(n43168), .B(n43167), .ZN(n43169) );
  XNOR2_X1 U45691 ( .A(n51439), .B(n43169), .ZN(n43172) );
  XNOR2_X1 U45692 ( .A(n43170), .B(n44061), .ZN(n43171) );
  XNOR2_X1 U45693 ( .A(n43172), .B(n43171), .ZN(n43174) );
  XNOR2_X1 U45694 ( .A(n43174), .B(n43173), .ZN(n43177) );
  XNOR2_X1 U45695 ( .A(n44925), .B(n44923), .ZN(n43175) );
  XNOR2_X1 U45696 ( .A(n44338), .B(n43175), .ZN(n45133) );
  XNOR2_X1 U45697 ( .A(n43195), .B(n45133), .ZN(n43176) );
  XNOR2_X2 U45698 ( .A(n43177), .B(n43176), .ZN(n49629) );
  NAND2_X1 U45701 ( .A1(n49980), .A2(n49629), .ZN(n49988) );
  INV_X1 U45702 ( .A(n43180), .ZN(n49972) );
  OAI21_X1 U45703 ( .B1(n49982), .B2(n49972), .A(n47360), .ZN(n43183) );
  NOR2_X1 U45704 ( .A1(n47354), .A2(n49980), .ZN(n43182) );
  INV_X1 U45705 ( .A(n43181), .ZN(n49983) );
  OAI21_X1 U45706 ( .B1(n43183), .B2(n43182), .A(n49973), .ZN(n43187) );
  NAND2_X1 U45707 ( .A1(n47349), .A2(n47354), .ZN(n43455) );
  INV_X1 U45708 ( .A(n47349), .ZN(n43185) );
  OAI21_X1 U45709 ( .B1(n43185), .B2(n43184), .A(n49980), .ZN(n43186) );
  OAI21_X1 U45710 ( .B1(n49573), .B2(n43188), .A(n49606), .ZN(n43419) );
  NOR2_X1 U45711 ( .A1(n49580), .A2(n49569), .ZN(n49610) );
  OR2_X1 U45712 ( .A1(n49592), .A2(n49610), .ZN(n43408) );
  XNOR2_X1 U45713 ( .A(n43189), .B(n49887), .ZN(n43190) );
  XNOR2_X1 U45714 ( .A(n43191), .B(n43190), .ZN(n43192) );
  XNOR2_X1 U45715 ( .A(n44547), .B(n43192), .ZN(n43193) );
  XNOR2_X1 U45716 ( .A(n43196), .B(n43197), .ZN(n43638) );
  XNOR2_X1 U45718 ( .A(n4045), .B(n4940), .ZN(n43199) );
  XNOR2_X1 U45719 ( .A(n43200), .B(n43199), .ZN(n43201) );
  XNOR2_X1 U45720 ( .A(n43202), .B(n43201), .ZN(n43203) );
  XNOR2_X1 U45721 ( .A(n43204), .B(n43203), .ZN(n43205) );
  XNOR2_X1 U45722 ( .A(n43206), .B(n43205), .ZN(n43207) );
  XNOR2_X1 U45723 ( .A(n43207), .B(n44562), .ZN(n43208) );
  XNOR2_X1 U45724 ( .A(n43208), .B(n44944), .ZN(n43211) );
  XNOR2_X1 U45725 ( .A(n43209), .B(n51330), .ZN(n43210) );
  XNOR2_X1 U45726 ( .A(n43755), .B(n43210), .ZN(n46040) );
  XNOR2_X1 U45727 ( .A(n43211), .B(n46040), .ZN(n43212) );
  XNOR2_X1 U45728 ( .A(n43213), .B(n43212), .ZN(n43215) );
  XNOR2_X1 U45729 ( .A(n44207), .B(n43216), .ZN(n43217) );
  XNOR2_X1 U45730 ( .A(n43218), .B(n43217), .ZN(n43231) );
  XNOR2_X1 U45731 ( .A(n44510), .B(n43219), .ZN(n43227) );
  XNOR2_X1 U45732 ( .A(n43221), .B(n43220), .ZN(n43222) );
  XNOR2_X1 U45733 ( .A(n43223), .B(n43222), .ZN(n43224) );
  XNOR2_X1 U45734 ( .A(n43225), .B(n43224), .ZN(n43226) );
  XNOR2_X1 U45735 ( .A(n43227), .B(n43226), .ZN(n43228) );
  XNOR2_X1 U45736 ( .A(n43229), .B(n43228), .ZN(n43230) );
  XNOR2_X1 U45737 ( .A(n43231), .B(n43230), .ZN(n43232) );
  XNOR2_X1 U45738 ( .A(n51525), .B(n43232), .ZN(n43278) );
  INV_X1 U45739 ( .A(n43278), .ZN(n49672) );
  XNOR2_X1 U45740 ( .A(n43234), .B(n43233), .ZN(n43235) );
  XNOR2_X1 U45741 ( .A(n43623), .B(n43235), .ZN(n43237) );
  XNOR2_X1 U45742 ( .A(n43236), .B(n43237), .ZN(n43239) );
  XNOR2_X1 U45743 ( .A(n43238), .B(n43239), .ZN(n43242) );
  XNOR2_X1 U45744 ( .A(n51681), .B(n46113), .ZN(n43240) );
  XNOR2_X1 U45745 ( .A(n43241), .B(n43242), .ZN(n43248) );
  XNOR2_X1 U45746 ( .A(n45415), .B(n43243), .ZN(n43246) );
  XNOR2_X1 U45747 ( .A(n43244), .B(n43245), .ZN(n46116) );
  XNOR2_X1 U45748 ( .A(n43246), .B(n46116), .ZN(n43247) );
  XNOR2_X1 U45749 ( .A(n43248), .B(n43247), .ZN(n43249) );
  AND2_X1 U45750 ( .A1(n52211), .A2(n49672), .ZN(n50027) );
  XNOR2_X1 U45751 ( .A(n43252), .B(n43251), .ZN(n43253) );
  XNOR2_X1 U45752 ( .A(n43254), .B(n43253), .ZN(n43255) );
  XNOR2_X1 U45753 ( .A(n43255), .B(n46138), .ZN(n43256) );
  XNOR2_X1 U45754 ( .A(n43256), .B(n46153), .ZN(n43257) );
  XNOR2_X1 U45755 ( .A(n44480), .B(n43261), .ZN(n43275) );
  XNOR2_X1 U45756 ( .A(n43263), .B(n43262), .ZN(n43264) );
  XNOR2_X1 U45757 ( .A(n43265), .B(n43264), .ZN(n43266) );
  XNOR2_X1 U45758 ( .A(n43266), .B(n44070), .ZN(n43268) );
  XNOR2_X1 U45759 ( .A(n43268), .B(n43267), .ZN(n43269) );
  XNOR2_X1 U45760 ( .A(n43496), .B(n43269), .ZN(n43270) );
  XNOR2_X1 U45761 ( .A(n52103), .B(n43270), .ZN(n43271) );
  XNOR2_X1 U45762 ( .A(n43271), .B(n45325), .ZN(n43273) );
  XNOR2_X1 U45763 ( .A(n43272), .B(n43273), .ZN(n43274) );
  NOR2_X1 U45764 ( .A1(n49659), .A2(n46028), .ZN(n43276) );
  OAI21_X1 U45765 ( .B1(n49669), .B2(n43276), .A(n50027), .ZN(n43277) );
  AND3_X1 U45766 ( .A1(n49660), .A2(n43277), .A3(n46027), .ZN(n43287) );
  AND3_X1 U45767 ( .A1(n49657), .A2(n49667), .A3(n51733), .ZN(n45959) );
  INV_X1 U45768 ( .A(n45959), .ZN(n43279) );
  OAI21_X1 U45769 ( .B1(n46030), .B2(n49656), .A(n43279), .ZN(n43280) );
  NAND2_X1 U45770 ( .A1(n49651), .A2(n49667), .ZN(n49645) );
  NOR2_X1 U45771 ( .A1(n49647), .A2(n49645), .ZN(n43448) );
  OAI21_X1 U45772 ( .B1(n43280), .B2(n43448), .A(n46028), .ZN(n43286) );
  INV_X1 U45773 ( .A(n49654), .ZN(n43442) );
  NAND2_X1 U45774 ( .A1(n46028), .A2(n52212), .ZN(n43282) );
  NAND4_X1 U45776 ( .A1(n43442), .A2(n43281), .A3(n49659), .A4(n45957), .ZN(
        n43285) );
  INV_X1 U45777 ( .A(n46030), .ZN(n43284) );
  INV_X1 U45778 ( .A(n43282), .ZN(n43283) );
  XNOR2_X1 U45779 ( .A(n43289), .B(n43288), .ZN(n43290) );
  XNOR2_X1 U45780 ( .A(n44286), .B(n43290), .ZN(n43292) );
  XNOR2_X1 U45781 ( .A(n43292), .B(n43291), .ZN(n43296) );
  XNOR2_X1 U45782 ( .A(n44296), .B(n44904), .ZN(n43295) );
  XNOR2_X1 U45783 ( .A(n44510), .B(n43293), .ZN(n43294) );
  XNOR2_X1 U45784 ( .A(n43295), .B(n43294), .ZN(n43979) );
  XNOR2_X1 U45785 ( .A(n44512), .B(n45252), .ZN(n45045) );
  XNOR2_X1 U45786 ( .A(n42906), .B(n45045), .ZN(n43298) );
  XNOR2_X1 U45787 ( .A(n43299), .B(n43298), .ZN(n46290) );
  XNOR2_X1 U45788 ( .A(n43301), .B(n43300), .ZN(n43302) );
  XNOR2_X1 U45789 ( .A(n43303), .B(n43302), .ZN(n43312) );
  XNOR2_X1 U45790 ( .A(n43305), .B(n43304), .ZN(n43306) );
  XNOR2_X1 U45791 ( .A(n44314), .B(n43306), .ZN(n43307) );
  XNOR2_X1 U45792 ( .A(n44240), .B(n43307), .ZN(n43309) );
  XNOR2_X1 U45793 ( .A(n43309), .B(n43308), .ZN(n43310) );
  XNOR2_X1 U45794 ( .A(n43310), .B(n45418), .ZN(n43311) );
  XNOR2_X1 U45795 ( .A(n43313), .B(n44076), .ZN(n45070) );
  XNOR2_X1 U45796 ( .A(n43314), .B(n1341), .ZN(n43315) );
  XNOR2_X1 U45797 ( .A(n43316), .B(n43315), .ZN(n43317) );
  XNOR2_X1 U45798 ( .A(n51461), .B(n43317), .ZN(n43319) );
  AND2_X1 U45799 ( .A1(n7000), .A2(n43327), .ZN(n43324) );
  AOI22_X1 U45800 ( .A1(n43326), .A2(n43325), .B1(n2413), .B2(n43324), .ZN(
        n43333) );
  OAI21_X1 U45801 ( .B1(n43328), .B2(n43335), .A(n43327), .ZN(n43332) );
  NAND3_X1 U45802 ( .A1(n43336), .A2(n43330), .A3(n43329), .ZN(n43331) );
  NAND2_X1 U45804 ( .A1(n43346), .A2(n43342), .ZN(n43340) );
  NAND2_X1 U45805 ( .A1(n43336), .A2(n43335), .ZN(n43337) );
  AND3_X1 U45806 ( .A1(n43339), .A2(n43338), .A3(n43337), .ZN(n43341) );
  NAND3_X1 U45807 ( .A1(n43340), .A2(n43341), .A3(n45339), .ZN(n43347) );
  INV_X1 U45808 ( .A(n43341), .ZN(n43345) );
  OR2_X1 U45809 ( .A1(n43345), .A2(n43342), .ZN(n43343) );
  XNOR2_X1 U45810 ( .A(n43348), .B(n44395), .ZN(n43350) );
  INV_X1 U45813 ( .A(n49146), .ZN(n45944) );
  XNOR2_X1 U45814 ( .A(n43352), .B(n43819), .ZN(n43362) );
  XNOR2_X1 U45815 ( .A(n43354), .B(n43353), .ZN(n44171) );
  XNOR2_X1 U45816 ( .A(n43355), .B(n49790), .ZN(n43356) );
  XNOR2_X1 U45817 ( .A(n43357), .B(n43356), .ZN(n43358) );
  XNOR2_X1 U45818 ( .A(n44171), .B(n43358), .ZN(n43359) );
  XNOR2_X1 U45819 ( .A(n43360), .B(n43359), .ZN(n43361) );
  XNOR2_X1 U45820 ( .A(n43365), .B(n43364), .ZN(n45095) );
  NOR2_X1 U45821 ( .A1(n45936), .A2(n43401), .ZN(n49145) );
  AND2_X1 U45822 ( .A1(n49142), .A2(n45937), .ZN(n43398) );
  XNOR2_X1 U45823 ( .A(n45445), .B(n43368), .ZN(n44147) );
  XNOR2_X1 U45824 ( .A(n43370), .B(n43369), .ZN(n43372) );
  XNOR2_X1 U45825 ( .A(n43372), .B(n43371), .ZN(n43373) );
  XNOR2_X1 U45826 ( .A(n43374), .B(n43373), .ZN(n43375) );
  XNOR2_X1 U45827 ( .A(n45306), .B(n43375), .ZN(n43376) );
  XNOR2_X1 U45828 ( .A(n43377), .B(n43376), .ZN(n43378) );
  XNOR2_X1 U45829 ( .A(n43378), .B(n43379), .ZN(n43384) );
  XNOR2_X1 U45830 ( .A(n43380), .B(n2112), .ZN(n43381) );
  XNOR2_X1 U45831 ( .A(n43381), .B(n43928), .ZN(n43382) );
  XNOR2_X1 U45832 ( .A(n43382), .B(n45304), .ZN(n43383) );
  XNOR2_X1 U45833 ( .A(n45455), .B(n43383), .ZN(n45120) );
  XNOR2_X1 U45834 ( .A(n43385), .B(n274), .ZN(n43386) );
  XNOR2_X1 U45835 ( .A(n43387), .B(n43386), .ZN(n43388) );
  XNOR2_X1 U45836 ( .A(n45284), .B(n43388), .ZN(n43389) );
  XNOR2_X1 U45837 ( .A(n43389), .B(n46068), .ZN(n43390) );
  XNOR2_X1 U45838 ( .A(n43392), .B(n43391), .ZN(n43393) );
  XNOR2_X1 U45839 ( .A(n52130), .B(n670), .ZN(n43395) );
  XNOR2_X1 U45840 ( .A(n43534), .B(n43395), .ZN(n43396) );
  OAI21_X1 U45842 ( .B1(n49145), .B2(n43398), .A(n46292), .ZN(n43406) );
  INV_X1 U45843 ( .A(n49154), .ZN(n43421) );
  OR2_X1 U45844 ( .A1(n46288), .A2(n43421), .ZN(n44727) );
  OR2_X1 U45845 ( .A1(n44727), .A2(n44733), .ZN(n45939) );
  INV_X1 U45846 ( .A(n45939), .ZN(n43400) );
  AND2_X1 U45847 ( .A1(n43421), .A2(n46288), .ZN(n46281) );
  AND2_X1 U45848 ( .A1(n46281), .A2(n49138), .ZN(n43399) );
  NOR2_X1 U45849 ( .A1(n43400), .A2(n43399), .ZN(n43405) );
  OR2_X2 U45850 ( .A1(n46288), .A2(n49154), .ZN(n49150) );
  INV_X1 U45851 ( .A(n49150), .ZN(n46298) );
  INV_X1 U45852 ( .A(n49139), .ZN(n44731) );
  OAI21_X1 U45853 ( .B1(n43427), .B2(n46288), .A(n49150), .ZN(n44726) );
  NAND2_X1 U45854 ( .A1(n43402), .A2(n44726), .ZN(n43404) );
  AND2_X1 U45855 ( .A1(n7657), .A2(n44730), .ZN(n46297) );
  NAND3_X1 U45856 ( .A1(n46297), .A2(n49142), .A3(n51515), .ZN(n43403) );
  NAND4_X2 U45857 ( .A1(n43404), .A2(n43405), .A3(n43406), .A4(n43403), .ZN(
        n49599) );
  NAND4_X1 U45858 ( .A1(n43408), .A2(n49579), .A3(n49585), .A4(n43407), .ZN(
        n43414) );
  INV_X1 U45859 ( .A(n49608), .ZN(n49562) );
  AOI21_X1 U45860 ( .B1(n49562), .B2(n49580), .A(n49569), .ZN(n43412) );
  NOR2_X1 U45861 ( .A1(n49608), .A2(n49599), .ZN(n45719) );
  AND2_X1 U45862 ( .A1(n49608), .A2(n49598), .ZN(n43409) );
  OR2_X1 U45863 ( .A1(n45719), .A2(n43409), .ZN(n43411) );
  NAND2_X1 U45864 ( .A1(n49580), .A2(n49599), .ZN(n43410) );
  OAI211_X1 U45865 ( .C1(n43412), .C2(n49600), .A(n43411), .B(n43410), .ZN(
        n43413) );
  NAND2_X1 U45866 ( .A1(n49606), .A2(n49608), .ZN(n49603) );
  NOR2_X1 U45867 ( .A1(n49603), .A2(n51088), .ZN(n43415) );
  INV_X1 U45868 ( .A(n49603), .ZN(n49556) );
  NOR2_X1 U45869 ( .A1(n49580), .A2(n49599), .ZN(n45726) );
  AOI22_X1 U45870 ( .A1(n43416), .A2(n43415), .B1(n49556), .B2(n45726), .ZN(
        n43417) );
  INV_X1 U45871 ( .A(n4755), .ZN(n43420) );
  NAND3_X1 U45872 ( .A1(n45943), .A2(n46292), .A3(n49148), .ZN(n43423) );
  NAND2_X1 U45873 ( .A1(n49142), .A2(n43421), .ZN(n43422) );
  NAND2_X1 U45874 ( .A1(n51515), .A2(n49137), .ZN(n45949) );
  INV_X1 U45876 ( .A(n43428), .ZN(n43426) );
  OAI21_X1 U45877 ( .B1(n49150), .B2(n45937), .A(n49146), .ZN(n43425) );
  NAND2_X1 U45878 ( .A1(n43426), .A2(n43425), .ZN(n43431) );
  NAND2_X1 U45879 ( .A1(n43429), .A2(n43428), .ZN(n43430) );
  INV_X1 U45880 ( .A(n44727), .ZN(n45945) );
  INV_X1 U45881 ( .A(n49209), .ZN(n45969) );
  OR2_X1 U45882 ( .A1(n46231), .A2(n45969), .ZN(n43438) );
  NAND2_X1 U45883 ( .A1(n45967), .A2(n49208), .ZN(n44753) );
  INV_X1 U45884 ( .A(n44753), .ZN(n46223) );
  AOI21_X1 U45885 ( .B1(n49208), .B2(n46214), .A(n45967), .ZN(n43433) );
  INV_X1 U45886 ( .A(n46232), .ZN(n49225) );
  OAI211_X1 U45887 ( .C1(n46223), .C2(n43433), .A(n46226), .B(n49225), .ZN(
        n43437) );
  NAND2_X1 U45888 ( .A1(n46222), .A2(n45966), .ZN(n43434) );
  NAND3_X1 U45889 ( .A1(n49225), .A2(n43434), .A3(n46229), .ZN(n43436) );
  OR2_X1 U45890 ( .A1(n46214), .A2(n52106), .ZN(n43435) );
  NOR2_X1 U45892 ( .A1(n49197), .A2(n49207), .ZN(n46215) );
  NAND2_X1 U45893 ( .A1(n46223), .A2(n46215), .ZN(n49226) );
  NAND3_X1 U45894 ( .A1(n46229), .A2(n49208), .A3(n44752), .ZN(n49212) );
  NOR2_X1 U45895 ( .A1(n46222), .A2(n49198), .ZN(n49222) );
  INV_X1 U45898 ( .A(n49651), .ZN(n43443) );
  OR2_X1 U45899 ( .A1(n52212), .A2(n51733), .ZN(n43446) );
  AOI21_X1 U45900 ( .B1(n50020), .B2(n43446), .A(n50019), .ZN(n43447) );
  NAND2_X1 U45901 ( .A1(n43448), .A2(n49663), .ZN(n43450) );
  NAND3_X1 U45902 ( .A1(n49654), .A2(n50021), .A3(n49667), .ZN(n43449) );
  OAI211_X1 U45903 ( .C1(n49979), .C2(n49983), .A(n43452), .B(n49980), .ZN(
        n43453) );
  NAND2_X1 U45904 ( .A1(n43453), .A2(n47360), .ZN(n43459) );
  NAND2_X1 U45905 ( .A1(n49972), .A2(n49629), .ZN(n49984) );
  NAND4_X1 U45906 ( .A1(n47354), .A2(n49982), .A3(n7798), .A4(n49972), .ZN(
        n46013) );
  AOI21_X1 U45907 ( .B1(n46014), .B2(n46013), .A(n49978), .ZN(n43458) );
  NAND3_X1 U45908 ( .A1(n49990), .A2(n49972), .A3(n49982), .ZN(n43456) );
  MUX2_X1 U45909 ( .A(n49626), .B(n43456), .S(n47349), .Z(n43457) );
  INV_X1 U45910 ( .A(n45999), .ZN(n49713) );
  NAND2_X1 U45911 ( .A1(n49725), .A2(n52052), .ZN(n45896) );
  NAND3_X1 U45912 ( .A1(n49713), .A2(n45896), .A3(n45907), .ZN(n43461) );
  MUX2_X1 U45913 ( .A(n43461), .B(n43460), .S(n45909), .Z(n43473) );
  NAND2_X1 U45914 ( .A1(n49189), .A2(n49721), .ZN(n49190) );
  NAND2_X1 U45915 ( .A1(n45993), .A2(n49190), .ZN(n43463) );
  INV_X1 U45916 ( .A(n43464), .ZN(n45997) );
  NAND2_X1 U45917 ( .A1(n43463), .A2(n45997), .ZN(n43472) );
  INV_X1 U45918 ( .A(n45987), .ZN(n49726) );
  NAND3_X1 U45919 ( .A1(n49726), .A2(n52052), .A3(n49717), .ZN(n43469) );
  NAND2_X1 U45920 ( .A1(n43464), .A2(n45909), .ZN(n43465) );
  NAND2_X1 U45921 ( .A1(n43465), .A2(n45989), .ZN(n43466) );
  NAND2_X1 U45922 ( .A1(n43467), .A2(n43466), .ZN(n43468) );
  AND3_X1 U45923 ( .A1(n43470), .A2(n43469), .A3(n43468), .ZN(n43471) );
  OAI21_X1 U45924 ( .B1(n49534), .B2(n49514), .A(n43490), .ZN(n49480) );
  INV_X1 U45925 ( .A(n45024), .ZN(n43487) );
  INV_X1 U45927 ( .A(n49232), .ZN(n44745) );
  AND2_X1 U45928 ( .A1(n44745), .A2(n49251), .ZN(n49694) );
  NAND3_X1 U45929 ( .A1(n49694), .A2(n49690), .A3(n49235), .ZN(n43478) );
  INV_X1 U45932 ( .A(n49696), .ZN(n45914) );
  XNOR2_X1 U45933 ( .A(n588), .B(n51095), .ZN(n43480) );
  OAI21_X1 U45934 ( .B1(n49246), .B2(n45914), .A(n43480), .ZN(n43477) );
  NAND2_X1 U45935 ( .A1(n49231), .A2(n45922), .ZN(n49243) );
  OAI22_X1 U45936 ( .A1(n49243), .A2(n51095), .B1(n45919), .B2(n587), .ZN(
        n43475) );
  NAND2_X1 U45937 ( .A1(n43475), .A2(n49248), .ZN(n43476) );
  NAND2_X1 U45938 ( .A1(n42883), .A2(n43479), .ZN(n49688) );
  NOR2_X1 U45939 ( .A1(n49688), .A2(n49235), .ZN(n49252) );
  INV_X1 U45940 ( .A(n49252), .ZN(n43484) );
  INV_X1 U45942 ( .A(n43480), .ZN(n43481) );
  NAND3_X1 U45943 ( .A1(n51731), .A2(n43481), .A3(n49247), .ZN(n43483) );
  NAND3_X1 U45944 ( .A1(n49251), .A2(n49242), .A3(n49686), .ZN(n43482) );
  NAND3_X1 U45946 ( .A1(n49480), .A2(n43487), .A3(n49503), .ZN(n43489) );
  NAND2_X1 U45948 ( .A1(n51395), .A2(n49514), .ZN(n49512) );
  NAND4_X1 U45951 ( .A1(n49508), .A2(n49510), .A3(n49512), .A4(n45022), .ZN(
        n43488) );
  NAND2_X1 U45952 ( .A1(n49539), .A2(n49522), .ZN(n43491) );
  OR2_X1 U45953 ( .A1(n49522), .A2(n49503), .ZN(n49506) );
  NOR2_X1 U45954 ( .A1(n49534), .A2(n49539), .ZN(n49530) );
  NAND2_X1 U45955 ( .A1(n2193), .A2(n49511), .ZN(n49476) );
  INV_X1 U45956 ( .A(n49476), .ZN(n43492) );
  NAND2_X1 U45957 ( .A1(n49530), .A2(n43492), .ZN(n49543) );
  INV_X1 U45958 ( .A(n4213), .ZN(n43495) );
  XNOR2_X1 U45959 ( .A(n43496), .B(n44156), .ZN(n43498) );
  XNOR2_X1 U45960 ( .A(n52103), .B(n43498), .ZN(n46092) );
  XNOR2_X1 U45961 ( .A(n43890), .B(n51294), .ZN(n43503) );
  XNOR2_X1 U45962 ( .A(n43500), .B(n43499), .ZN(n43501) );
  XNOR2_X1 U45963 ( .A(n45339), .B(n43501), .ZN(n43502) );
  XNOR2_X1 U45964 ( .A(n43503), .B(n43502), .ZN(n43505) );
  XNOR2_X1 U45965 ( .A(n43505), .B(n43504), .ZN(n43506) );
  XNOR2_X1 U45966 ( .A(n43584), .B(n51460), .ZN(n43507) );
  XNOR2_X1 U45967 ( .A(n43507), .B(n44074), .ZN(n43508) );
  XNOR2_X1 U45968 ( .A(n43508), .B(n45325), .ZN(n43774) );
  XNOR2_X1 U45969 ( .A(n51096), .B(n46153), .ZN(n43614) );
  XNOR2_X1 U45970 ( .A(n43509), .B(n43614), .ZN(n43519) );
  XNOR2_X1 U45971 ( .A(n44501), .B(n45089), .ZN(n43515) );
  XNOR2_X1 U45972 ( .A(n46144), .B(n43510), .ZN(n43511) );
  XNOR2_X1 U45973 ( .A(n43512), .B(n43511), .ZN(n43513) );
  XNOR2_X1 U45974 ( .A(n46150), .B(n43513), .ZN(n43514) );
  XNOR2_X1 U45975 ( .A(n43515), .B(n43514), .ZN(n43517) );
  XNOR2_X1 U45976 ( .A(n43516), .B(n45365), .ZN(n43946) );
  XNOR2_X1 U45977 ( .A(n43517), .B(n43946), .ZN(n43518) );
  INV_X1 U45978 ( .A(n46062), .ZN(n43521) );
  XNOR2_X1 U45979 ( .A(n46059), .B(n43521), .ZN(n43911) );
  INV_X1 U45980 ( .A(n43911), .ZN(n43523) );
  XNOR2_X1 U45981 ( .A(n43523), .B(n43522), .ZN(n43526) );
  XNOR2_X1 U45982 ( .A(n43642), .B(n52222), .ZN(n43525) );
  XNOR2_X1 U45983 ( .A(n44330), .B(n47244), .ZN(n43527) );
  XNOR2_X1 U45984 ( .A(n43528), .B(n43527), .ZN(n43529) );
  XNOR2_X1 U45985 ( .A(n43530), .B(n43529), .ZN(n43531) );
  XNOR2_X1 U45986 ( .A(n51464), .B(n43531), .ZN(n43532) );
  XNOR2_X1 U45987 ( .A(n43532), .B(n44923), .ZN(n43533) );
  XNOR2_X1 U45988 ( .A(n44061), .B(n44534), .ZN(n46073) );
  XNOR2_X1 U45990 ( .A(n44565), .B(n43657), .ZN(n43546) );
  XNOR2_X1 U45991 ( .A(n43929), .B(n43536), .ZN(n43544) );
  XNOR2_X1 U45992 ( .A(n43538), .B(n43537), .ZN(n43540) );
  XNOR2_X1 U45993 ( .A(n43540), .B(n43539), .ZN(n43541) );
  XNOR2_X1 U45994 ( .A(n46050), .B(n43541), .ZN(n43542) );
  XNOR2_X1 U45995 ( .A(n43751), .B(n43542), .ZN(n43543) );
  XNOR2_X1 U45996 ( .A(n43544), .B(n43543), .ZN(n43545) );
  XNOR2_X1 U45997 ( .A(n43546), .B(n43545), .ZN(n43550) );
  XNOR2_X1 U45998 ( .A(n46049), .B(n44130), .ZN(n43548) );
  XNOR2_X1 U45999 ( .A(n43548), .B(n44944), .ZN(n45449) );
  XNOR2_X1 U46000 ( .A(n51503), .B(n45449), .ZN(n43549) );
  NAND2_X1 U46002 ( .A1(n50314), .A2(n52224), .ZN(n43581) );
  INV_X1 U46003 ( .A(n43581), .ZN(n50006) );
  XOR2_X1 U46004 ( .A(n43553), .B(n43552), .Z(n43554) );
  XNOR2_X1 U46005 ( .A(n44300), .B(n43554), .ZN(n43555) );
  XNOR2_X1 U46006 ( .A(n45393), .B(n43555), .ZN(n43556) );
  XNOR2_X1 U46007 ( .A(n43557), .B(n43556), .ZN(n43559) );
  XNOR2_X1 U46008 ( .A(n43558), .B(n43559), .ZN(n43562) );
  XNOR2_X1 U46009 ( .A(n51448), .B(n44288), .ZN(n43976) );
  INV_X1 U46010 ( .A(n43976), .ZN(n43561) );
  XNOR2_X1 U46011 ( .A(n43698), .B(n43560), .ZN(n43830) );
  XNOR2_X1 U46012 ( .A(n43564), .B(n43563), .ZN(n43565) );
  XNOR2_X1 U46013 ( .A(n46113), .B(n43565), .ZN(n43566) );
  XNOR2_X1 U46014 ( .A(n43566), .B(n43567), .ZN(n43568) );
  XNOR2_X1 U46015 ( .A(n43568), .B(n46131), .ZN(n43570) );
  XNOR2_X1 U46016 ( .A(n43570), .B(n43569), .ZN(n43574) );
  XNOR2_X1 U46017 ( .A(n46128), .B(n43571), .ZN(n43572) );
  XNOR2_X1 U46018 ( .A(n608), .B(n43572), .ZN(n43846) );
  XNOR2_X1 U46019 ( .A(n43846), .B(n43717), .ZN(n43573) );
  XNOR2_X1 U46021 ( .A(n43575), .B(n43856), .ZN(n45281) );
  XNOR2_X1 U46022 ( .A(n45281), .B(n45059), .ZN(n43629) );
  NAND3_X1 U46023 ( .A1(n49994), .A2(n50006), .A3(n50322), .ZN(n46010) );
  INV_X1 U46024 ( .A(n50317), .ZN(n43577) );
  OR2_X1 U46025 ( .A1(n49995), .A2(n43581), .ZN(n50332) );
  NAND2_X1 U46026 ( .A1(n46008), .A2(n50325), .ZN(n50331) );
  INV_X1 U46027 ( .A(n50314), .ZN(n50321) );
  AND2_X1 U46029 ( .A1(n50314), .A2(n43577), .ZN(n49996) );
  NAND4_X1 U46030 ( .A1(n47369), .A2(n49996), .A3(n47368), .A4(n50322), .ZN(
        n43579) );
  OR2_X1 U46031 ( .A1(n43581), .A2(n51526), .ZN(n50013) );
  NAND2_X1 U46032 ( .A1(n50013), .A2(n49993), .ZN(n43582) );
  INV_X1 U46033 ( .A(n50325), .ZN(n50015) );
  NAND4_X1 U46034 ( .A1(n43582), .A2(n50015), .A3(n1812), .A4(n50322), .ZN(
        n43583) );
  XNOR2_X1 U46035 ( .A(n45327), .B(n43584), .ZN(n43595) );
  XNOR2_X1 U46036 ( .A(n4823), .B(n4733), .ZN(n43585) );
  XNOR2_X1 U46037 ( .A(n43586), .B(n43585), .ZN(n43587) );
  XNOR2_X1 U46038 ( .A(n43588), .B(n43587), .ZN(n43590) );
  XNOR2_X1 U46039 ( .A(n43590), .B(n43589), .ZN(n43591) );
  XNOR2_X1 U46040 ( .A(n43592), .B(n43591), .ZN(n43593) );
  XNOR2_X1 U46041 ( .A(n45484), .B(n43593), .ZN(n43594) );
  XNOR2_X1 U46042 ( .A(n43595), .B(n43594), .ZN(n43600) );
  XNOR2_X1 U46044 ( .A(n43596), .B(n44074), .ZN(n43597) );
  XNOR2_X1 U46045 ( .A(n43598), .B(n43597), .ZN(n43599) );
  XNOR2_X1 U46046 ( .A(n43600), .B(n43599), .ZN(n43601) );
  XNOR2_X1 U46047 ( .A(n43763), .B(n43601), .ZN(n43602) );
  XNOR2_X1 U46048 ( .A(n43604), .B(n43603), .ZN(n43617) );
  XNOR2_X1 U46049 ( .A(n43605), .B(n49790), .ZN(n43606) );
  XNOR2_X1 U46050 ( .A(n43607), .B(n43606), .ZN(n43608) );
  XNOR2_X1 U46051 ( .A(n45354), .B(n43608), .ZN(n43611) );
  XNOR2_X1 U46052 ( .A(n43609), .B(n45358), .ZN(n43610) );
  XNOR2_X1 U46053 ( .A(n43611), .B(n43610), .ZN(n43613) );
  INV_X1 U46054 ( .A(n45365), .ZN(n43734) );
  XNOR2_X1 U46055 ( .A(n43734), .B(n44373), .ZN(n43612) );
  XNOR2_X1 U46056 ( .A(n43613), .B(n43612), .ZN(n43615) );
  XNOR2_X1 U46057 ( .A(n43615), .B(n43614), .ZN(n43616) );
  INV_X1 U46059 ( .A(n45165), .ZN(n43631) );
  XNOR2_X1 U46060 ( .A(n51450), .B(n608), .ZN(n43618) );
  XNOR2_X1 U46061 ( .A(n43859), .B(n43618), .ZN(n43628) );
  XNOR2_X1 U46062 ( .A(n45274), .B(n43710), .ZN(n43626) );
  XNOR2_X1 U46063 ( .A(n43621), .B(n43620), .ZN(n43622) );
  XNOR2_X1 U46064 ( .A(n43623), .B(n4781), .ZN(n45057) );
  XNOR2_X1 U46065 ( .A(n43624), .B(n45057), .ZN(n43625) );
  XNOR2_X1 U46066 ( .A(n43626), .B(n43625), .ZN(n43627) );
  XNOR2_X1 U46067 ( .A(n43628), .B(n43627), .ZN(n43630) );
  NAND2_X1 U46068 ( .A1(n43631), .A2(n47162), .ZN(n46995) );
  XNOR2_X1 U46069 ( .A(n4035), .B(n4752), .ZN(n43632) );
  XNOR2_X1 U46070 ( .A(n43633), .B(n43632), .ZN(n43634) );
  XNOR2_X1 U46071 ( .A(n43635), .B(n43634), .ZN(n43636) );
  XNOR2_X1 U46072 ( .A(n44534), .B(n43636), .ZN(n43637) );
  XNOR2_X1 U46073 ( .A(n2196), .B(n44327), .ZN(n45287) );
  XNOR2_X1 U46074 ( .A(n43637), .B(n45287), .ZN(n43639) );
  XNOR2_X1 U46075 ( .A(n44535), .B(n43640), .ZN(n45434) );
  XNOR2_X1 U46076 ( .A(n42170), .B(n45426), .ZN(n43641) );
  XNOR2_X1 U46077 ( .A(n45434), .B(n43641), .ZN(n43643) );
  XNOR2_X1 U46078 ( .A(n43642), .B(n43643), .ZN(n43644) );
  XNOR2_X1 U46079 ( .A(n44043), .B(n43647), .ZN(n43648) );
  XNOR2_X1 U46080 ( .A(n43649), .B(n43648), .ZN(n43650) );
  XNOR2_X1 U46081 ( .A(n43920), .B(n43650), .ZN(n43651) );
  XNOR2_X1 U46082 ( .A(n45305), .B(n43651), .ZN(n43652) );
  XNOR2_X1 U46083 ( .A(n43652), .B(n51097), .ZN(n43653) );
  XNOR2_X1 U46084 ( .A(n51503), .B(n43653), .ZN(n43659) );
  XNOR2_X1 U46085 ( .A(n45097), .B(n43654), .ZN(n43656) );
  XNOR2_X1 U46086 ( .A(n43655), .B(n43656), .ZN(n44932) );
  XNOR2_X1 U46087 ( .A(n43657), .B(n44562), .ZN(n45320) );
  INV_X1 U46088 ( .A(n45159), .ZN(n46994) );
  XNOR2_X1 U46089 ( .A(n43661), .B(n43660), .ZN(n43681) );
  XNOR2_X1 U46090 ( .A(n44006), .B(n51371), .ZN(n43664) );
  INV_X1 U46091 ( .A(n43662), .ZN(n43663) );
  XNOR2_X1 U46092 ( .A(n44510), .B(n43663), .ZN(n45262) );
  XNOR2_X1 U46093 ( .A(n43664), .B(n45262), .ZN(n43679) );
  OAI21_X1 U46094 ( .B1(n43667), .B2(n43666), .A(n43665), .ZN(n43668) );
  AND3_X1 U46095 ( .A1(n43670), .A2(n43669), .A3(n43668), .ZN(n43673) );
  XNOR2_X1 U46096 ( .A(n43675), .B(n43674), .ZN(n43676) );
  XNOR2_X1 U46097 ( .A(n45041), .B(n43676), .ZN(n43677) );
  XNOR2_X1 U46098 ( .A(n45258), .B(n43677), .ZN(n43678) );
  XNOR2_X1 U46099 ( .A(n43679), .B(n43678), .ZN(n43680) );
  XNOR2_X1 U46100 ( .A(n43681), .B(n43680), .ZN(n43682) );
  NAND2_X2 U46101 ( .A1(n8655), .A2(n388), .ZN(n47159) );
  NAND4_X1 U46102 ( .A1(n46995), .A2(n46994), .A3(n47159), .A4(n43683), .ZN(
        n43690) );
  OAI211_X1 U46103 ( .C1(n46999), .C2(n47151), .A(n47153), .B(n47162), .ZN(
        n43684) );
  OAI21_X1 U46104 ( .B1(n47159), .B2(n45164), .A(n43684), .ZN(n43685) );
  AND2_X1 U46105 ( .A1(n47152), .A2(n663), .ZN(n47003) );
  NAND3_X1 U46106 ( .A1(n47150), .A2(n2751), .A3(n46999), .ZN(n43686) );
  NAND2_X1 U46107 ( .A1(n46999), .A2(n389), .ZN(n44471) );
  NAND2_X1 U46108 ( .A1(n45157), .A2(n45159), .ZN(n43689) );
  AND2_X1 U46109 ( .A1(n44471), .A2(n47153), .ZN(n45153) );
  NAND2_X1 U46110 ( .A1(n45156), .A2(n46998), .ZN(n44473) );
  NAND2_X1 U46111 ( .A1(n45156), .A2(n663), .ZN(n46894) );
  XNOR2_X1 U46113 ( .A(n43692), .B(n43691), .ZN(n43693) );
  XNOR2_X1 U46114 ( .A(n43694), .B(n43693), .ZN(n43695) );
  XNOR2_X1 U46115 ( .A(n43696), .B(n43695), .ZN(n43697) );
  XNOR2_X1 U46116 ( .A(n44301), .B(n43697), .ZN(n43699) );
  XNOR2_X1 U46117 ( .A(n43699), .B(n43698), .ZN(n43701) );
  XNOR2_X1 U46118 ( .A(n43701), .B(n43700), .ZN(n43706) );
  XNOR2_X1 U46119 ( .A(n44216), .B(n45262), .ZN(n43704) );
  XNOR2_X1 U46120 ( .A(n44017), .B(n43702), .ZN(n44905) );
  XNOR2_X1 U46121 ( .A(n44905), .B(n43703), .ZN(n43978) );
  XNOR2_X1 U46122 ( .A(n43704), .B(n43978), .ZN(n43705) );
  XNOR2_X1 U46123 ( .A(n43706), .B(n43705), .ZN(n43709) );
  XNOR2_X1 U46124 ( .A(n45394), .B(n45393), .ZN(n43708) );
  XNOR2_X1 U46125 ( .A(n43708), .B(n43707), .ZN(n45047) );
  XNOR2_X1 U46126 ( .A(n44525), .B(n43710), .ZN(n43711) );
  XNOR2_X1 U46127 ( .A(n43962), .B(n43711), .ZN(n43720) );
  XNOR2_X1 U46128 ( .A(n43713), .B(n43712), .ZN(n43714) );
  XNOR2_X1 U46129 ( .A(n51681), .B(n43714), .ZN(n43715) );
  XNOR2_X1 U46130 ( .A(n43716), .B(n43715), .ZN(n43718) );
  XNOR2_X1 U46131 ( .A(n43718), .B(n43717), .ZN(n43719) );
  XNOR2_X1 U46132 ( .A(n43720), .B(n43719), .ZN(n43722) );
  INV_X1 U46133 ( .A(n46971), .ZN(n46969) );
  XNOR2_X1 U46134 ( .A(n45460), .B(n43723), .ZN(n44099) );
  XNOR2_X1 U46135 ( .A(n44099), .B(n52123), .ZN(n43947) );
  INV_X1 U46136 ( .A(n43947), .ZN(n43726) );
  XNOR2_X1 U46137 ( .A(n43725), .B(n43724), .ZN(n44983) );
  XNOR2_X1 U46138 ( .A(n43726), .B(n44983), .ZN(n43738) );
  XNOR2_X1 U46139 ( .A(n43728), .B(n43727), .ZN(n43729) );
  XNOR2_X1 U46140 ( .A(n43730), .B(n43729), .ZN(n43731) );
  XNOR2_X1 U46141 ( .A(n45354), .B(n43731), .ZN(n43733) );
  XNOR2_X1 U46142 ( .A(n46150), .B(n51398), .ZN(n43732) );
  XNOR2_X1 U46143 ( .A(n43733), .B(n43732), .ZN(n43736) );
  XNOR2_X1 U46144 ( .A(n44374), .B(n43734), .ZN(n43735) );
  XNOR2_X1 U46145 ( .A(n43736), .B(n43735), .ZN(n43737) );
  XNOR2_X1 U46146 ( .A(n43738), .B(n43737), .ZN(n43743) );
  XNOR2_X1 U46147 ( .A(n52084), .B(n43739), .ZN(n43741) );
  XNOR2_X1 U46148 ( .A(n43742), .B(n43741), .ZN(n45473) );
  BUF_X2 U46149 ( .A(n46978), .Z(n50367) );
  XNOR2_X1 U46150 ( .A(n43745), .B(n43744), .ZN(n43747) );
  XNOR2_X1 U46151 ( .A(n43747), .B(n43746), .ZN(n43748) );
  XNOR2_X1 U46152 ( .A(n51330), .B(n43748), .ZN(n43749) );
  XNOR2_X1 U46153 ( .A(n51097), .B(n43749), .ZN(n43750) );
  XNOR2_X1 U46154 ( .A(n43750), .B(n45303), .ZN(n43753) );
  XNOR2_X1 U46155 ( .A(n44134), .B(n44562), .ZN(n45447) );
  XNOR2_X1 U46156 ( .A(n45447), .B(n43751), .ZN(n43752) );
  XNOR2_X1 U46157 ( .A(n43753), .B(n43752), .ZN(n43762) );
  XNOR2_X1 U46158 ( .A(n43755), .B(n43754), .ZN(n43756) );
  XNOR2_X1 U46159 ( .A(n516), .B(n43756), .ZN(n43760) );
  XNOR2_X1 U46160 ( .A(n43758), .B(n43759), .ZN(n43932) );
  NOR2_X1 U46161 ( .A1(n47139), .A2(n50364), .ZN(n43777) );
  NAND2_X1 U46162 ( .A1(n50364), .A2(n50367), .ZN(n50365) );
  XNOR2_X1 U46163 ( .A(n43764), .B(n4654), .ZN(n43765) );
  XNOR2_X1 U46164 ( .A(n43766), .B(n43765), .ZN(n43767) );
  XNOR2_X1 U46165 ( .A(n43768), .B(n43767), .ZN(n43770) );
  XNOR2_X1 U46166 ( .A(n43770), .B(n43769), .ZN(n43771) );
  XNOR2_X1 U46167 ( .A(n45327), .B(n43771), .ZN(n43772) );
  XNOR2_X1 U46168 ( .A(n43772), .B(n44154), .ZN(n43773) );
  XNOR2_X1 U46169 ( .A(n43774), .B(n43773), .ZN(n43775) );
  OAI21_X1 U46170 ( .B1(n50365), .B2(n667), .A(n43798), .ZN(n43776) );
  NOR2_X1 U46171 ( .A1(n43777), .A2(n43776), .ZN(n43778) );
  OAI21_X1 U46172 ( .B1(n46977), .B2(n50367), .A(n43778), .ZN(n43801) );
  INV_X1 U46173 ( .A(n46978), .ZN(n46989) );
  NAND2_X1 U46174 ( .A1(n46989), .A2(n50364), .ZN(n46982) );
  XNOR2_X1 U46175 ( .A(n44547), .B(n45421), .ZN(n43904) );
  XNOR2_X1 U46176 ( .A(n43904), .B(n43779), .ZN(n43780) );
  XNOR2_X1 U46177 ( .A(n43916), .B(n43780), .ZN(n43793) );
  INV_X1 U46178 ( .A(n43781), .ZN(n43782) );
  XNOR2_X1 U46179 ( .A(n43782), .B(n51464), .ZN(n44548) );
  XOR2_X1 U46180 ( .A(n4706), .B(n842), .Z(n43783) );
  XNOR2_X1 U46181 ( .A(n43784), .B(n43783), .ZN(n43785) );
  XNOR2_X1 U46182 ( .A(n43786), .B(n43785), .ZN(n43787) );
  XNOR2_X1 U46183 ( .A(n671), .B(n43787), .ZN(n43788) );
  XNOR2_X1 U46184 ( .A(n44548), .B(n43788), .ZN(n43791) );
  XNOR2_X1 U46185 ( .A(n44061), .B(n46068), .ZN(n43789) );
  XNOR2_X1 U46186 ( .A(n43789), .B(n45434), .ZN(n43790) );
  XNOR2_X1 U46187 ( .A(n43791), .B(n43790), .ZN(n43792) );
  XNOR2_X1 U46188 ( .A(n43793), .B(n43792), .ZN(n43794) );
  XNOR2_X1 U46189 ( .A(n45439), .B(n43794), .ZN(n43795) );
  NOR2_X1 U46190 ( .A1(n46982), .A2(n50366), .ZN(n43796) );
  INV_X1 U46191 ( .A(n43795), .ZN(n50368) );
  AOI22_X1 U46192 ( .A1(n43796), .A2(n50363), .B1(n50368), .B2(n43798), .ZN(
        n43800) );
  AND2_X1 U46193 ( .A1(n46984), .A2(n50370), .ZN(n47143) );
  NAND2_X1 U46194 ( .A1(n47139), .A2(n50368), .ZN(n47142) );
  XNOR2_X1 U46196 ( .A(n43196), .B(n43802), .ZN(n43809) );
  XNOR2_X1 U46197 ( .A(n43803), .B(n47244), .ZN(n43804) );
  XNOR2_X1 U46198 ( .A(n43805), .B(n43804), .ZN(n43806) );
  XNOR2_X1 U46199 ( .A(n44327), .B(n43806), .ZN(n43807) );
  XNOR2_X1 U46200 ( .A(n43807), .B(n45432), .ZN(n43808) );
  XNOR2_X1 U46201 ( .A(n43809), .B(n43808), .ZN(n43810) );
  XNOR2_X1 U46202 ( .A(n45133), .B(n43810), .ZN(n43814) );
  XNOR2_X1 U46203 ( .A(n43812), .B(n43811), .ZN(n43813) );
  XNOR2_X1 U46205 ( .A(n43816), .B(n43815), .ZN(n43818) );
  XNOR2_X1 U46206 ( .A(n43818), .B(n43817), .ZN(n43827) );
  XNOR2_X1 U46207 ( .A(n43821), .B(n43820), .ZN(n43822) );
  XNOR2_X1 U46208 ( .A(n45358), .B(n43822), .ZN(n43823) );
  XNOR2_X1 U46209 ( .A(n45089), .B(n43823), .ZN(n43824) );
  XNOR2_X1 U46210 ( .A(n43825), .B(n43824), .ZN(n43826) );
  XNOR2_X1 U46211 ( .A(n43827), .B(n43826), .ZN(n43829) );
  INV_X1 U46212 ( .A(n50350), .ZN(n47030) );
  INV_X1 U46213 ( .A(n50349), .ZN(n47293) );
  XNOR2_X1 U46214 ( .A(n43831), .B(n43830), .ZN(n43842) );
  XNOR2_X1 U46215 ( .A(n44300), .B(n43832), .ZN(n43834) );
  XNOR2_X1 U46216 ( .A(n43834), .B(n51333), .ZN(n43840) );
  XNOR2_X1 U46217 ( .A(n43836), .B(n43835), .ZN(n43837) );
  XNOR2_X1 U46218 ( .A(n43973), .B(n43837), .ZN(n43838) );
  XNOR2_X1 U46219 ( .A(n45258), .B(n43838), .ZN(n43839) );
  XNOR2_X1 U46220 ( .A(n43840), .B(n43839), .ZN(n43841) );
  XNOR2_X1 U46221 ( .A(n43841), .B(n43842), .ZN(n43844) );
  XNOR2_X1 U46222 ( .A(n43845), .B(n45274), .ZN(n44321) );
  XNOR2_X1 U46225 ( .A(n43849), .B(n43848), .ZN(n43851) );
  XNOR2_X1 U46226 ( .A(n43851), .B(n43850), .ZN(n43853) );
  XNOR2_X1 U46227 ( .A(n43853), .B(n43852), .ZN(n43854) );
  XNOR2_X1 U46228 ( .A(n51431), .B(n43854), .ZN(n43855) );
  XNOR2_X1 U46229 ( .A(n43855), .B(n51681), .ZN(n43857) );
  XNOR2_X1 U46230 ( .A(n43857), .B(n51390), .ZN(n43858) );
  XNOR2_X1 U46231 ( .A(n43859), .B(n43858), .ZN(n43860) );
  AND2_X1 U46233 ( .A1(n47278), .A2(n51386), .ZN(n50347) );
  XNOR2_X1 U46234 ( .A(n43863), .B(n43862), .ZN(n43864) );
  XNOR2_X1 U46235 ( .A(n45105), .B(n43864), .ZN(n43865) );
  XNOR2_X1 U46236 ( .A(n43866), .B(n43865), .ZN(n43867) );
  XNOR2_X1 U46237 ( .A(n44937), .B(n43867), .ZN(n43868) );
  XNOR2_X1 U46238 ( .A(n43868), .B(n43920), .ZN(n43869) );
  XNOR2_X1 U46239 ( .A(n43869), .B(n2206), .ZN(n43871) );
  XNOR2_X1 U46240 ( .A(n43871), .B(n43870), .ZN(n43874) );
  XNOR2_X1 U46241 ( .A(n43872), .B(n44038), .ZN(n43873) );
  XNOR2_X1 U46242 ( .A(n43873), .B(n43874), .ZN(n43877) );
  XNOR2_X1 U46243 ( .A(n45116), .B(n52171), .ZN(n43875) );
  XNOR2_X1 U46244 ( .A(n43875), .B(n44131), .ZN(n43876) );
  XNOR2_X1 U46245 ( .A(n43148), .B(n43876), .ZN(n44361) );
  INV_X1 U46246 ( .A(n50344), .ZN(n50348) );
  XOR2_X1 U46247 ( .A(n43879), .B(n43878), .Z(n43880) );
  XNOR2_X1 U46248 ( .A(n43881), .B(n43880), .ZN(n43882) );
  XNOR2_X1 U46249 ( .A(n44963), .B(n43882), .ZN(n43883) );
  XNOR2_X1 U46250 ( .A(n43883), .B(n44391), .ZN(n43886) );
  XNOR2_X1 U46251 ( .A(n43884), .B(n46090), .ZN(n43885) );
  XNOR2_X1 U46252 ( .A(n43886), .B(n43885), .ZN(n43888) );
  XNOR2_X1 U46253 ( .A(n43887), .B(n43888), .ZN(n43895) );
  XNOR2_X1 U46254 ( .A(n45325), .B(n43889), .ZN(n43891) );
  XNOR2_X1 U46255 ( .A(n43890), .B(n44962), .ZN(n43992) );
  XNOR2_X1 U46256 ( .A(n43891), .B(n43992), .ZN(n43893) );
  XNOR2_X1 U46257 ( .A(n43893), .B(n43892), .ZN(n43894) );
  NAND3_X1 U46258 ( .A1(n50347), .A2(n50348), .A3(n47271), .ZN(n47023) );
  NOR2_X1 U46259 ( .A1(n47030), .A2(n51026), .ZN(n47031) );
  XNOR2_X1 U46260 ( .A(n51386), .B(n50344), .ZN(n43896) );
  NAND2_X1 U46261 ( .A1(n43896), .A2(n505), .ZN(n43897) );
  OAI21_X1 U46262 ( .B1(n50347), .B2(n47031), .A(n43897), .ZN(n43899) );
  OR2_X1 U46263 ( .A1(n50352), .A2(n51725), .ZN(n43898) );
  OAI21_X1 U46264 ( .B1(n50348), .B2(n51386), .A(n47271), .ZN(n43901) );
  INV_X1 U46266 ( .A(n47291), .ZN(n43900) );
  OR2_X1 U46267 ( .A1(n505), .A2(n51025), .ZN(n47270) );
  NAND3_X1 U46268 ( .A1(n43901), .A2(n43900), .A3(n47270), .ZN(n43902) );
  OR2_X1 U46270 ( .A1(n50620), .A2(n50578), .ZN(n50591) );
  XNOR2_X1 U46271 ( .A(n44548), .B(n44327), .ZN(n43905) );
  XNOR2_X1 U46272 ( .A(n43905), .B(n43904), .ZN(n44188) );
  XNOR2_X1 U46273 ( .A(n43907), .B(n43906), .ZN(n43908) );
  XNOR2_X1 U46274 ( .A(n43909), .B(n43908), .ZN(n43910) );
  XNOR2_X1 U46275 ( .A(n44542), .B(n43910), .ZN(n43912) );
  XNOR2_X1 U46276 ( .A(n43912), .B(n43911), .ZN(n43913) );
  XNOR2_X1 U46277 ( .A(n44188), .B(n43913), .ZN(n43919) );
  XNOR2_X1 U46278 ( .A(n51439), .B(n43915), .ZN(n46074) );
  XNOR2_X1 U46279 ( .A(n43916), .B(n46074), .ZN(n43917) );
  XNOR2_X1 U46280 ( .A(n44553), .B(n43917), .ZN(n43918) );
  INV_X1 U46282 ( .A(n50265), .ZN(n44583) );
  XNOR2_X1 U46283 ( .A(n44134), .B(n43920), .ZN(n43924) );
  XNOR2_X1 U46284 ( .A(n4637), .B(n4885), .ZN(n43921) );
  XNOR2_X1 U46285 ( .A(n43921), .B(n4045), .ZN(n43923) );
  XNOR2_X1 U46286 ( .A(n43926), .B(n43925), .ZN(n43931) );
  XNOR2_X1 U46287 ( .A(n43928), .B(n43927), .ZN(n44945) );
  XNOR2_X1 U46288 ( .A(n44945), .B(n43929), .ZN(n43930) );
  XNOR2_X1 U46289 ( .A(n43931), .B(n43930), .ZN(n43933) );
  XNOR2_X1 U46290 ( .A(n43932), .B(n43933), .ZN(n43935) );
  INV_X1 U46291 ( .A(n50276), .ZN(n43966) );
  XNOR2_X1 U46292 ( .A(n43939), .B(n43938), .ZN(n43940) );
  XNOR2_X1 U46293 ( .A(n43941), .B(n43940), .ZN(n43942) );
  XNOR2_X1 U46294 ( .A(n45358), .B(n43942), .ZN(n43944) );
  XNOR2_X1 U46295 ( .A(n43944), .B(n43943), .ZN(n43945) );
  XNOR2_X1 U46296 ( .A(n43946), .B(n43945), .ZN(n43948) );
  AND2_X1 U46297 ( .A1(n44583), .A2(n50280), .ZN(n50252) );
  INV_X1 U46298 ( .A(n47058), .ZN(n50270) );
  XNOR2_X1 U46299 ( .A(n51681), .B(n44027), .ZN(n43949) );
  XNOR2_X1 U46300 ( .A(n43949), .B(n45274), .ZN(n43958) );
  XNOR2_X1 U46301 ( .A(n43950), .B(n46111), .ZN(n43956) );
  XNOR2_X1 U46302 ( .A(n43952), .B(n43951), .ZN(n43953) );
  XNOR2_X1 U46303 ( .A(n43954), .B(n43953), .ZN(n43955) );
  XNOR2_X1 U46304 ( .A(n43956), .B(n43955), .ZN(n43957) );
  XNOR2_X1 U46305 ( .A(n43958), .B(n43957), .ZN(n43959) );
  XNOR2_X1 U46306 ( .A(n43960), .B(n43959), .ZN(n43964) );
  INV_X1 U46307 ( .A(n51307), .ZN(n43961) );
  XNOR2_X1 U46308 ( .A(n608), .B(n43961), .ZN(n45049) );
  XNOR2_X1 U46309 ( .A(n43962), .B(n45049), .ZN(n43963) );
  NAND2_X1 U46310 ( .A1(n50281), .A2(n44001), .ZN(n43965) );
  XNOR2_X1 U46311 ( .A(n47737), .B(n4641), .ZN(n43967) );
  XNOR2_X1 U46312 ( .A(n43968), .B(n43967), .ZN(n43969) );
  XNOR2_X1 U46313 ( .A(n43970), .B(n43969), .ZN(n43971) );
  XNOR2_X1 U46314 ( .A(n44016), .B(n43971), .ZN(n43972) );
  XNOR2_X1 U46315 ( .A(n43972), .B(n44216), .ZN(n43975) );
  XNOR2_X1 U46316 ( .A(n43973), .B(n45258), .ZN(n43974) );
  XNOR2_X1 U46317 ( .A(n43975), .B(n43974), .ZN(n43977) );
  XNOR2_X1 U46318 ( .A(n43977), .B(n43976), .ZN(n43981) );
  XNOR2_X1 U46319 ( .A(n43979), .B(n43978), .ZN(n43980) );
  XNOR2_X1 U46320 ( .A(n43981), .B(n43980), .ZN(n43982) );
  NAND2_X1 U46321 ( .A1(n47044), .A2(n47341), .ZN(n47334) );
  NAND2_X1 U46322 ( .A1(n43984), .A2(n47334), .ZN(n44117) );
  XNOR2_X1 U46323 ( .A(n43068), .B(n45325), .ZN(n44168) );
  XNOR2_X1 U46324 ( .A(n43985), .B(n48814), .ZN(n43987) );
  XNOR2_X1 U46325 ( .A(n43987), .B(n43986), .ZN(n43989) );
  XNOR2_X1 U46326 ( .A(n43989), .B(n43988), .ZN(n43990) );
  XNOR2_X1 U46327 ( .A(n44156), .B(n43990), .ZN(n43991) );
  XNOR2_X1 U46328 ( .A(n43992), .B(n43991), .ZN(n43993) );
  XNOR2_X1 U46329 ( .A(n43993), .B(n45068), .ZN(n43994) );
  XNOR2_X1 U46330 ( .A(n44168), .B(n43994), .ZN(n43998) );
  XNOR2_X1 U46331 ( .A(n43995), .B(n43996), .ZN(n43997) );
  XNOR2_X1 U46332 ( .A(n43998), .B(n43997), .ZN(n44118) );
  NAND2_X1 U46333 ( .A1(n44117), .A2(n44118), .ZN(n44004) );
  INV_X1 U46334 ( .A(n47334), .ZN(n50255) );
  NAND2_X1 U46335 ( .A1(n50281), .A2(n50255), .ZN(n47340) );
  NAND2_X1 U46336 ( .A1(n47335), .A2(n50252), .ZN(n43999) );
  AND2_X1 U46337 ( .A1(n47340), .A2(n43999), .ZN(n44116) );
  NOR3_X1 U46338 ( .A1(n47058), .A2(n51410), .A3(n47341), .ZN(n44000) );
  NOR2_X1 U46339 ( .A1(n47058), .A2(n50254), .ZN(n44586) );
  OAI21_X1 U46340 ( .B1(n44000), .B2(n44586), .A(n47046), .ZN(n44115) );
  AND2_X1 U46341 ( .A1(n5237), .A2(n50254), .ZN(n50278) );
  NAND2_X1 U46342 ( .A1(n50276), .A2(n50278), .ZN(n47062) );
  NAND4_X1 U46343 ( .A1(n44116), .A2(n50277), .A3(n44115), .A4(n47062), .ZN(
        n44003) );
  OR2_X1 U46344 ( .A1(n50261), .A2(n47333), .ZN(n47061) );
  NAND3_X1 U46345 ( .A1(n50262), .A2(n50251), .A3(n50253), .ZN(n44002) );
  NAND3_X1 U46346 ( .A1(n47061), .A2(n44002), .A3(n47064), .ZN(n44121) );
  AOI21_X2 U46347 ( .B1(n44004), .B2(n44003), .A(n44121), .ZN(n50618) );
  NOR2_X1 U46348 ( .A1(n50618), .A2(n50638), .ZN(n44124) );
  INV_X1 U46349 ( .A(n44124), .ZN(n44005) );
  OAI21_X1 U46350 ( .B1(n50610), .B2(n50591), .A(n44005), .ZN(n44114) );
  XNOR2_X1 U46351 ( .A(n44006), .B(n44301), .ZN(n44007) );
  XNOR2_X1 U46352 ( .A(n44009), .B(n44008), .ZN(n44021) );
  XNOR2_X1 U46353 ( .A(n44010), .B(n47737), .ZN(n44011) );
  XNOR2_X1 U46354 ( .A(n44012), .B(n44011), .ZN(n44013) );
  XNOR2_X1 U46355 ( .A(n45041), .B(n44013), .ZN(n44014) );
  XNOR2_X1 U46356 ( .A(n44216), .B(n44014), .ZN(n44019) );
  XNOR2_X1 U46357 ( .A(n44016), .B(n44015), .ZN(n44018) );
  XNOR2_X1 U46358 ( .A(n44018), .B(n44017), .ZN(n44514) );
  XNOR2_X1 U46359 ( .A(n44019), .B(n44514), .ZN(n44020) );
  XNOR2_X1 U46360 ( .A(n44021), .B(n44020), .ZN(n44023) );
  XNOR2_X1 U46362 ( .A(n44025), .B(n44024), .ZN(n44026) );
  XNOR2_X1 U46363 ( .A(n44027), .B(n44026), .ZN(n44028) );
  XNOR2_X1 U46364 ( .A(n44240), .B(n44028), .ZN(n44029) );
  XNOR2_X1 U46365 ( .A(n44893), .B(n44029), .ZN(n44035) );
  INV_X1 U46366 ( .A(n4826), .ZN(n48657) );
  XNOR2_X1 U46367 ( .A(n44030), .B(n48657), .ZN(n44877) );
  XNOR2_X1 U46368 ( .A(n44877), .B(n608), .ZN(n44033) );
  XNOR2_X1 U46369 ( .A(n44033), .B(n44032), .ZN(n44034) );
  XNOR2_X1 U46370 ( .A(n44035), .B(n44034), .ZN(n44037) );
  AND2_X1 U46371 ( .A1(n46810), .A2(n46828), .ZN(n47075) );
  XNOR2_X1 U46372 ( .A(n46050), .B(n45114), .ZN(n44940) );
  XNOR2_X1 U46373 ( .A(n52043), .B(n44940), .ZN(n44039) );
  XNOR2_X1 U46374 ( .A(n44041), .B(n51337), .ZN(n44049) );
  XNOR2_X1 U46375 ( .A(n44044), .B(n44043), .ZN(n44045) );
  XNOR2_X1 U46376 ( .A(n44046), .B(n44045), .ZN(n44047) );
  XNOR2_X1 U46377 ( .A(n44134), .B(n44047), .ZN(n44048) );
  XNOR2_X1 U46378 ( .A(n44049), .B(n44048), .ZN(n44051) );
  XNOR2_X1 U46379 ( .A(n44051), .B(n44050), .ZN(n44053) );
  XNOR2_X1 U46380 ( .A(n44353), .B(n50987), .ZN(n44052) );
  XNOR2_X1 U46381 ( .A(n44052), .B(n51097), .ZN(n44568) );
  XNOR2_X1 U46382 ( .A(n44053), .B(n44568), .ZN(n44054) );
  XNOR2_X1 U46383 ( .A(n44057), .B(n4639), .ZN(n44058) );
  XNOR2_X1 U46384 ( .A(n44059), .B(n44058), .ZN(n44060) );
  XNOR2_X1 U46385 ( .A(n45421), .B(n44060), .ZN(n44062) );
  XNOR2_X1 U46386 ( .A(n44061), .B(n44062), .ZN(n44063) );
  XNOR2_X1 U46387 ( .A(n44064), .B(n44063), .ZN(n44068) );
  XNOR2_X1 U46388 ( .A(n671), .B(n46058), .ZN(n44065) );
  XNOR2_X1 U46389 ( .A(n44066), .B(n44065), .ZN(n44067) );
  AND2_X1 U46390 ( .A1(n47076), .A2(n46828), .ZN(n46775) );
  XNOR2_X1 U46391 ( .A(n44070), .B(n44069), .ZN(n44071) );
  XNOR2_X1 U46392 ( .A(n44072), .B(n44071), .ZN(n44073) );
  XNOR2_X1 U46393 ( .A(n44074), .B(n44073), .ZN(n44075) );
  XNOR2_X1 U46394 ( .A(n44076), .B(n44075), .ZN(n44078) );
  XNOR2_X1 U46395 ( .A(n44078), .B(n44077), .ZN(n44083) );
  XNOR2_X1 U46396 ( .A(n46079), .B(n44079), .ZN(n44080) );
  XNOR2_X1 U46397 ( .A(n44081), .B(n44080), .ZN(n44082) );
  XNOR2_X1 U46398 ( .A(n44083), .B(n44082), .ZN(n44084) );
  XNOR2_X1 U46399 ( .A(n44086), .B(n44372), .ZN(n44095) );
  XOR2_X1 U46400 ( .A(n4869), .B(n4836), .Z(n44087) );
  XNOR2_X1 U46401 ( .A(n44088), .B(n44087), .ZN(n44089) );
  XNOR2_X1 U46402 ( .A(n44090), .B(n44089), .ZN(n44091) );
  XNOR2_X1 U46403 ( .A(n44979), .B(n44091), .ZN(n44093) );
  XNOR2_X1 U46404 ( .A(n44093), .B(n44092), .ZN(n44094) );
  XNOR2_X1 U46405 ( .A(n44095), .B(n44094), .ZN(n44097) );
  XNOR2_X1 U46406 ( .A(n44097), .B(n44096), .ZN(n44102) );
  XNOR2_X1 U46407 ( .A(n44098), .B(n44099), .ZN(n44100) );
  XNOR2_X1 U46408 ( .A(n44100), .B(n44503), .ZN(n44101) );
  XNOR2_X1 U46409 ( .A(n44102), .B(n44101), .ZN(n46774) );
  AND2_X1 U46410 ( .A1(n46774), .A2(n46816), .ZN(n46832) );
  AOI22_X1 U46411 ( .A1(n47075), .A2(n46822), .B1(n46775), .B2(n46832), .ZN(
        n44106) );
  INV_X1 U46412 ( .A(n46832), .ZN(n44103) );
  OR2_X1 U46413 ( .A1(n44103), .A2(n46772), .ZN(n46766) );
  INV_X1 U46414 ( .A(n46774), .ZN(n45179) );
  AND2_X1 U46415 ( .A1(n45179), .A2(n46816), .ZN(n46823) );
  NAND3_X1 U46416 ( .A1(n47069), .A2(n400), .A3(n46822), .ZN(n44104) );
  AND4_X1 U46417 ( .A1(n44106), .A2(n46766), .A3(n44105), .A4(n44104), .ZN(
        n44112) );
  INV_X1 U46418 ( .A(n46772), .ZN(n44110) );
  NAND2_X1 U46419 ( .A1(n47069), .A2(n44458), .ZN(n46831) );
  AND2_X1 U46420 ( .A1(n45176), .A2(n51292), .ZN(n44108) );
  MUX2_X1 U46421 ( .A(n51419), .B(n51456), .S(n46774), .Z(n44107) );
  AOI22_X1 U46422 ( .A1(n44110), .A2(n46831), .B1(n44108), .B2(n44107), .ZN(
        n44111) );
  NAND3_X1 U46423 ( .A1(n44458), .A2(n46824), .A3(n400), .ZN(n46778) );
  AOI21_X1 U46424 ( .B1(n44114), .B2(n50630), .A(n50575), .ZN(n44125) );
  INV_X1 U46425 ( .A(n50620), .ZN(n50598) );
  NOR2_X1 U46426 ( .A1(n50598), .A2(n52226), .ZN(n50588) );
  NAND3_X1 U46427 ( .A1(n44116), .A2(n44115), .A3(n47062), .ZN(n44120) );
  INV_X1 U46428 ( .A(n44117), .ZN(n44119) );
  MUX2_X1 U46429 ( .A(n44120), .B(n44119), .S(n44118), .Z(n44122) );
  NAND2_X1 U46430 ( .A1(n50620), .A2(n51029), .ZN(n47217) );
  INV_X1 U46433 ( .A(n50618), .ZN(n50644) );
  NAND3_X1 U46434 ( .A1(n50644), .A2(n50609), .A3(n52226), .ZN(n50593) );
  NAND2_X1 U46435 ( .A1(n50642), .A2(n52081), .ZN(n47221) );
  NAND2_X1 U46436 ( .A1(n52082), .A2(n50578), .ZN(n50579) );
  NAND2_X1 U46437 ( .A1(n47221), .A2(n50579), .ZN(n44127) );
  INV_X1 U46438 ( .A(n50575), .ZN(n44126) );
  NAND4_X1 U46439 ( .A1(n44128), .A2(n50641), .A3(n44127), .A4(n44126), .ZN(
        n44129) );
  XNOR2_X1 U46440 ( .A(n44559), .B(n44130), .ZN(n44132) );
  XNOR2_X1 U46441 ( .A(n44132), .B(n44131), .ZN(n44142) );
  XNOR2_X1 U46442 ( .A(n44133), .B(n44134), .ZN(n44140) );
  INV_X1 U46443 ( .A(n44135), .ZN(n44137) );
  XNOR2_X1 U46444 ( .A(n44137), .B(n44136), .ZN(n44138) );
  XNOR2_X1 U46445 ( .A(n45114), .B(n44138), .ZN(n44139) );
  XNOR2_X1 U46446 ( .A(n44140), .B(n44139), .ZN(n44141) );
  XNOR2_X1 U46447 ( .A(n44142), .B(n44141), .ZN(n44145) );
  XNOR2_X1 U46448 ( .A(n607), .B(n44143), .ZN(n44144) );
  XNOR2_X1 U46449 ( .A(n44144), .B(n45303), .ZN(n44359) );
  XNOR2_X1 U46450 ( .A(n44359), .B(n44145), .ZN(n44151) );
  INV_X1 U46451 ( .A(n44146), .ZN(n44148) );
  XNOR2_X1 U46452 ( .A(n44148), .B(n44147), .ZN(n46041) );
  XNOR2_X1 U46453 ( .A(n46041), .B(n44149), .ZN(n44150) );
  XNOR2_X1 U46454 ( .A(n44151), .B(n44150), .ZN(n44206) );
  INV_X1 U46455 ( .A(n44206), .ZN(n46474) );
  XNOR2_X1 U46456 ( .A(n44152), .B(n46081), .ZN(n44159) );
  XNOR2_X1 U46457 ( .A(n44153), .B(n44154), .ZN(n44158) );
  XNOR2_X1 U46458 ( .A(n44156), .B(n44155), .ZN(n44157) );
  XNOR2_X1 U46459 ( .A(n44158), .B(n44157), .ZN(n45078) );
  XNOR2_X1 U46460 ( .A(n44159), .B(n45078), .ZN(n44167) );
  XNOR2_X1 U46461 ( .A(n44160), .B(n51461), .ZN(n45489) );
  XNOR2_X1 U46462 ( .A(n44162), .B(n44161), .ZN(n44163) );
  XNOR2_X1 U46463 ( .A(n44164), .B(n44163), .ZN(n44165) );
  XNOR2_X1 U46464 ( .A(n45489), .B(n44165), .ZN(n44166) );
  INV_X1 U46465 ( .A(n46313), .ZN(n44246) );
  XNOR2_X1 U46466 ( .A(n46138), .B(n50967), .ZN(n44169) );
  XNOR2_X1 U46467 ( .A(n44170), .B(n44169), .ZN(n45093) );
  XNOR2_X1 U46468 ( .A(n45358), .B(n46137), .ZN(n44362) );
  XNOR2_X1 U46469 ( .A(n44171), .B(n44362), .ZN(n44180) );
  XNOR2_X1 U46470 ( .A(n44172), .B(n4895), .ZN(n44174) );
  XNOR2_X1 U46471 ( .A(n44174), .B(n44173), .ZN(n44175) );
  XNOR2_X1 U46472 ( .A(n44176), .B(n44175), .ZN(n44178) );
  XNOR2_X1 U46473 ( .A(n44178), .B(n44177), .ZN(n44179) );
  XNOR2_X1 U46474 ( .A(n44180), .B(n44179), .ZN(n44181) );
  XNOR2_X1 U46475 ( .A(n45093), .B(n44181), .ZN(n44187) );
  XNOR2_X1 U46476 ( .A(n44182), .B(n44373), .ZN(n44183) );
  XNOR2_X1 U46477 ( .A(n44184), .B(n44183), .ZN(n46142) );
  XNOR2_X1 U46478 ( .A(n46142), .B(n44185), .ZN(n44186) );
  XNOR2_X1 U46479 ( .A(n44188), .B(n45437), .ZN(n44205) );
  XNOR2_X1 U46480 ( .A(n44189), .B(n44190), .ZN(n44200) );
  INV_X1 U46481 ( .A(n44191), .ZN(n44192) );
  XNOR2_X1 U46482 ( .A(n44192), .B(n4639), .ZN(n44194) );
  XNOR2_X1 U46483 ( .A(n44194), .B(n44193), .ZN(n44195) );
  XNOR2_X1 U46484 ( .A(n44196), .B(n44195), .ZN(n44197) );
  XNOR2_X1 U46485 ( .A(n44198), .B(n44197), .ZN(n44199) );
  XNOR2_X1 U46486 ( .A(n44200), .B(n44199), .ZN(n44201) );
  XNOR2_X1 U46487 ( .A(n45429), .B(n44201), .ZN(n44203) );
  XNOR2_X1 U46488 ( .A(n44203), .B(n44202), .ZN(n44204) );
  XNOR2_X1 U46492 ( .A(n44207), .B(n44299), .ZN(n44214) );
  INV_X1 U46493 ( .A(n44208), .ZN(n44210) );
  XNOR2_X1 U46494 ( .A(n44209), .B(n44210), .ZN(n44211) );
  XNOR2_X1 U46495 ( .A(n51448), .B(n44211), .ZN(n44213) );
  XNOR2_X1 U46496 ( .A(n44213), .B(n44214), .ZN(n44215) );
  XNOR2_X1 U46497 ( .A(n44215), .B(n45376), .ZN(n44228) );
  XNOR2_X1 U46498 ( .A(n44216), .B(n44286), .ZN(n44219) );
  XNOR2_X1 U46499 ( .A(n7101), .B(n47737), .ZN(n44218) );
  XNOR2_X1 U46500 ( .A(n44219), .B(n44218), .ZN(n45378) );
  INV_X1 U46501 ( .A(n44220), .ZN(n44222) );
  XNOR2_X1 U46502 ( .A(n44222), .B(n44221), .ZN(n44223) );
  XNOR2_X1 U46503 ( .A(n44900), .B(n44224), .ZN(n44225) );
  XNOR2_X1 U46504 ( .A(n44288), .B(n44225), .ZN(n44226) );
  XNOR2_X1 U46505 ( .A(n45378), .B(n44226), .ZN(n44227) );
  XNOR2_X1 U46507 ( .A(n44230), .B(n44229), .ZN(n44231) );
  XNOR2_X1 U46508 ( .A(n44318), .B(n44231), .ZN(n44245) );
  XNOR2_X1 U46509 ( .A(n45403), .B(n4668), .ZN(n44232) );
  XNOR2_X1 U46510 ( .A(n44233), .B(n44232), .ZN(n44235) );
  XNOR2_X1 U46511 ( .A(n44235), .B(n44234), .ZN(n44236) );
  XNOR2_X1 U46512 ( .A(n46128), .B(n44236), .ZN(n44239) );
  XNOR2_X1 U46513 ( .A(n45408), .B(n44237), .ZN(n44238) );
  XNOR2_X1 U46514 ( .A(n44239), .B(n44238), .ZN(n44242) );
  XNOR2_X1 U46515 ( .A(n44242), .B(n44241), .ZN(n44243) );
  XNOR2_X1 U46516 ( .A(n44529), .B(n44243), .ZN(n44244) );
  OR2_X1 U46518 ( .A1(n46322), .A2(n52066), .ZN(n48196) );
  AOI22_X1 U46519 ( .A1(n44246), .A2(n46478), .B1(n48512), .B2(n48196), .ZN(
        n44253) );
  INV_X1 U46520 ( .A(n46322), .ZN(n46475) );
  INV_X1 U46522 ( .A(n48521), .ZN(n44252) );
  OR2_X1 U46523 ( .A1(n46474), .A2(n52202), .ZN(n44249) );
  INV_X1 U46524 ( .A(n44249), .ZN(n44248) );
  NAND3_X1 U46527 ( .A1(n44248), .A2(n48510), .A3(n48498), .ZN(n44251) );
  NOR2_X1 U46528 ( .A1(n48196), .A2(n44249), .ZN(n46315) );
  INV_X1 U46529 ( .A(n46315), .ZN(n44250) );
  OAI211_X1 U46530 ( .C1(n44253), .C2(n44252), .A(n44251), .B(n44250), .ZN(
        n44254) );
  INV_X1 U46531 ( .A(n45559), .ZN(n45562) );
  AND2_X1 U46532 ( .A1(n48505), .A2(n45562), .ZN(n45558) );
  NAND2_X1 U46533 ( .A1(n45558), .A2(n46471), .ZN(n48189) );
  NOR2_X1 U46534 ( .A1(n48521), .A2(n46474), .ZN(n44257) );
  MUX2_X1 U46535 ( .A(n46322), .B(n52066), .S(n46471), .Z(n44256) );
  AND2_X1 U46536 ( .A1(n48505), .A2(n52203), .ZN(n48508) );
  INV_X1 U46537 ( .A(n48508), .ZN(n44255) );
  OAI22_X1 U46538 ( .A1(n48189), .A2(n44257), .B1(n44256), .B2(n44255), .ZN(
        n44258) );
  INV_X1 U46539 ( .A(n44258), .ZN(n44260) );
  MUX2_X1 U46540 ( .A(n46318), .B(n48521), .S(n48512), .Z(n45557) );
  NAND3_X1 U46541 ( .A1(n45557), .A2(n48510), .A3(n46474), .ZN(n44259) );
  NAND2_X1 U46542 ( .A1(n48207), .A2(n48221), .ZN(n44261) );
  NAND2_X1 U46543 ( .A1(n44262), .A2(n48205), .ZN(n44274) );
  INV_X1 U46545 ( .A(n44998), .ZN(n44266) );
  NOR2_X1 U46546 ( .A1(n48210), .A2(n48200), .ZN(n44265) );
  AND2_X1 U46547 ( .A1(n44263), .A2(n52050), .ZN(n44264) );
  AOI22_X1 U46548 ( .A1(n44266), .A2(n44265), .B1(n44264), .B2(n48214), .ZN(
        n44273) );
  AND2_X1 U46549 ( .A1(n52161), .A2(n48210), .ZN(n45544) );
  NAND2_X1 U46550 ( .A1(n48205), .A2(n44693), .ZN(n45541) );
  INV_X1 U46551 ( .A(n45541), .ZN(n44268) );
  NAND2_X1 U46552 ( .A1(n45540), .A2(n44992), .ZN(n48218) );
  OAI21_X1 U46553 ( .B1(n45538), .B2(n45547), .A(n48218), .ZN(n44267) );
  AOI21_X1 U46554 ( .B1(n45544), .B2(n44268), .A(n44267), .ZN(n44272) );
  OAI21_X1 U46555 ( .B1(n44270), .B2(n45545), .A(n44269), .ZN(n44271) );
  AND2_X1 U46556 ( .A1(n48051), .A2(n48084), .ZN(n48021) );
  NAND2_X1 U46557 ( .A1(n45524), .A2(n45818), .ZN(n44275) );
  OAI21_X1 U46558 ( .B1(n45533), .B2(n45827), .A(n44275), .ZN(n44276) );
  NAND2_X1 U46559 ( .A1(n44276), .A2(n44828), .ZN(n44285) );
  OR2_X1 U46560 ( .A1(n45524), .A2(n42176), .ZN(n44279) );
  NAND2_X1 U46561 ( .A1(n44831), .A2(n44640), .ZN(n44277) );
  NAND2_X1 U46562 ( .A1(n45834), .A2(n44277), .ZN(n44641) );
  INV_X1 U46563 ( .A(n44641), .ZN(n44278) );
  AOI22_X1 U46564 ( .A1(n44279), .A2(n44278), .B1(n45523), .B2(n45829), .ZN(
        n44284) );
  NAND2_X1 U46565 ( .A1(n45524), .A2(n44281), .ZN(n44282) );
  INV_X1 U46566 ( .A(n45532), .ZN(n44283) );
  XNOR2_X1 U46568 ( .A(n44287), .B(n44286), .ZN(n44289) );
  XNOR2_X1 U46569 ( .A(n44288), .B(n44289), .ZN(n44290) );
  XNOR2_X1 U46570 ( .A(n44291), .B(n44290), .ZN(n44306) );
  INV_X1 U46571 ( .A(n44292), .ZN(n44294) );
  XNOR2_X1 U46572 ( .A(n44294), .B(n44293), .ZN(n44295) );
  XNOR2_X1 U46573 ( .A(n44911), .B(n44295), .ZN(n44297) );
  XNOR2_X1 U46574 ( .A(n44296), .B(n44297), .ZN(n44298) );
  XNOR2_X1 U46575 ( .A(n44299), .B(n44298), .ZN(n44304) );
  XNOR2_X1 U46576 ( .A(n44301), .B(n44300), .ZN(n46103) );
  XNOR2_X1 U46577 ( .A(n46103), .B(n44302), .ZN(n44303) );
  XNOR2_X1 U46578 ( .A(n44304), .B(n44303), .ZN(n44305) );
  XNOR2_X1 U46579 ( .A(n44306), .B(n44305), .ZN(n44409) );
  INV_X1 U46580 ( .A(n44409), .ZN(n44673) );
  XNOR2_X1 U46581 ( .A(n44307), .B(n44308), .ZN(n44317) );
  XOR2_X1 U46582 ( .A(n4535), .B(n4668), .Z(n44309) );
  XNOR2_X1 U46583 ( .A(n44310), .B(n44309), .ZN(n44312) );
  XNOR2_X1 U46584 ( .A(n44312), .B(n44311), .ZN(n44313) );
  XNOR2_X1 U46585 ( .A(n44314), .B(n44313), .ZN(n44315) );
  XNOR2_X1 U46586 ( .A(n44317), .B(n44316), .ZN(n44319) );
  XNOR2_X1 U46587 ( .A(n44318), .B(n44319), .ZN(n44323) );
  XNOR2_X1 U46588 ( .A(n44321), .B(n44320), .ZN(n44322) );
  INV_X1 U46589 ( .A(n48251), .ZN(n44380) );
  XNOR2_X1 U46590 ( .A(n46068), .B(n44542), .ZN(n44324) );
  XNOR2_X1 U46591 ( .A(n44327), .B(n45293), .ZN(n44337) );
  INV_X1 U46592 ( .A(n44328), .ZN(n44334) );
  XNOR2_X1 U46593 ( .A(n44330), .B(n44329), .ZN(n44331) );
  XNOR2_X1 U46594 ( .A(n44332), .B(n44331), .ZN(n44333) );
  XNOR2_X1 U46595 ( .A(n44334), .B(n44333), .ZN(n44335) );
  XNOR2_X1 U46596 ( .A(n45285), .B(n44335), .ZN(n44336) );
  XNOR2_X1 U46597 ( .A(n44337), .B(n44336), .ZN(n44339) );
  XNOR2_X1 U46598 ( .A(n44338), .B(n44339), .ZN(n44340) );
  XNOR2_X1 U46599 ( .A(n44341), .B(n44340), .ZN(n44346) );
  XNOR2_X1 U46600 ( .A(n670), .B(n44342), .ZN(n44343) );
  XNOR2_X1 U46601 ( .A(n44344), .B(n44343), .ZN(n44345) );
  XNOR2_X1 U46602 ( .A(n45097), .B(n45445), .ZN(n44348) );
  XNOR2_X1 U46603 ( .A(n44348), .B(n44347), .ZN(n44357) );
  XNOR2_X1 U46604 ( .A(n44350), .B(n44349), .ZN(n44351) );
  XNOR2_X1 U46605 ( .A(n51330), .B(n44351), .ZN(n44355) );
  INV_X1 U46606 ( .A(n44353), .ZN(n44354) );
  XNOR2_X1 U46607 ( .A(n44355), .B(n44354), .ZN(n44356) );
  XNOR2_X1 U46608 ( .A(n44357), .B(n44356), .ZN(n44358) );
  XNOR2_X1 U46609 ( .A(n44359), .B(n44358), .ZN(n44360) );
  INV_X1 U46610 ( .A(n48485), .ZN(n44402) );
  XNOR2_X1 U46611 ( .A(n45355), .B(n44501), .ZN(n44363) );
  XNOR2_X1 U46612 ( .A(n44363), .B(n44362), .ZN(n44365) );
  XNOR2_X1 U46613 ( .A(n44364), .B(n44365), .ZN(n44377) );
  XNOR2_X1 U46614 ( .A(n44366), .B(n44493), .ZN(n44368) );
  XNOR2_X1 U46615 ( .A(n44368), .B(n44367), .ZN(n44369) );
  XNOR2_X1 U46616 ( .A(n44370), .B(n44369), .ZN(n44371) );
  XNOR2_X1 U46617 ( .A(n44372), .B(n44371), .ZN(n44375) );
  XNOR2_X1 U46618 ( .A(n44374), .B(n44373), .ZN(n45462) );
  XNOR2_X1 U46619 ( .A(n44375), .B(n45462), .ZN(n44376) );
  XNOR2_X1 U46620 ( .A(n44376), .B(n44377), .ZN(n44379) );
  NAND3_X1 U46621 ( .A1(n44380), .A2(n44402), .A3(n48487), .ZN(n44383) );
  INV_X1 U46622 ( .A(n48479), .ZN(n48246) );
  NOR2_X1 U46623 ( .A1(n46458), .A2(n48246), .ZN(n48253) );
  INV_X1 U46624 ( .A(n48253), .ZN(n44382) );
  NAND2_X1 U46625 ( .A1(n48246), .A2(n44673), .ZN(n44410) );
  AND2_X1 U46626 ( .A1(n44410), .A2(n48248), .ZN(n46456) );
  NAND2_X1 U46627 ( .A1(n46456), .A2(n44681), .ZN(n44381) );
  NAND3_X1 U46628 ( .A1(n44383), .A2(n44382), .A3(n44381), .ZN(n44408) );
  INV_X1 U46629 ( .A(n48474), .ZN(n45600) );
  OR2_X1 U46630 ( .A1(n48487), .A2(n44409), .ZN(n44400) );
  NAND2_X1 U46631 ( .A1(n48487), .A2(n44409), .ZN(n44384) );
  NAND4_X1 U46632 ( .A1(n45600), .A2(n44400), .A3(n48479), .A4(n44384), .ZN(
        n44404) );
  INV_X1 U46633 ( .A(n44385), .ZN(n44388) );
  XNOR2_X1 U46634 ( .A(n44386), .B(n47679), .ZN(n44387) );
  XNOR2_X1 U46635 ( .A(n44388), .B(n44387), .ZN(n44389) );
  XNOR2_X1 U46636 ( .A(n51460), .B(n44389), .ZN(n44390) );
  XNOR2_X1 U46637 ( .A(n44391), .B(n44390), .ZN(n44393) );
  XNOR2_X1 U46638 ( .A(n44393), .B(n44392), .ZN(n44396) );
  XNOR2_X1 U46639 ( .A(n44395), .B(n44394), .ZN(n44967) );
  XNOR2_X1 U46640 ( .A(n44396), .B(n44967), .ZN(n44399) );
  INV_X1 U46641 ( .A(n44400), .ZN(n44401) );
  NAND2_X1 U46642 ( .A1(n44402), .A2(n44401), .ZN(n44403) );
  NAND3_X1 U46643 ( .A1(n44404), .A2(n48478), .A3(n44403), .ZN(n44407) );
  NAND3_X1 U46644 ( .A1(n48251), .A2(n45600), .A3(n48475), .ZN(n44405) );
  NAND2_X1 U46645 ( .A1(n44405), .A2(n48482), .ZN(n44406) );
  OAI21_X1 U46646 ( .B1(n44408), .B2(n44407), .A(n44406), .ZN(n44416) );
  AND2_X1 U46647 ( .A1(n48487), .A2(n48491), .ZN(n45598) );
  AND2_X1 U46648 ( .A1(n44410), .A2(n48482), .ZN(n48493) );
  AND3_X1 U46649 ( .A1(n45598), .A2(n48493), .A3(n48247), .ZN(n44412) );
  AND2_X1 U46650 ( .A1(n48474), .A2(n48248), .ZN(n44411) );
  AND2_X1 U46651 ( .A1(n48493), .A2(n44411), .ZN(n44679) );
  NOR2_X1 U46652 ( .A1(n44412), .A2(n44679), .ZN(n44415) );
  OAI21_X1 U46653 ( .B1(n45598), .B2(n46456), .A(n48478), .ZN(n44413) );
  NAND2_X1 U46654 ( .A1(n44413), .A2(n48244), .ZN(n44414) );
  INV_X1 U46656 ( .A(n48083), .ZN(n48041) );
  NOR2_X1 U46657 ( .A1(n48041), .A2(n51092), .ZN(n48081) );
  OR2_X1 U46658 ( .A1(n44652), .A2(n46642), .ZN(n46623) );
  NOR2_X1 U46659 ( .A1(n46632), .A2(n46623), .ZN(n46626) );
  OAI21_X1 U46660 ( .B1(n44423), .B2(n46633), .A(n46628), .ZN(n44417) );
  AND2_X1 U46661 ( .A1(n52153), .A2(n47909), .ZN(n44418) );
  AND2_X1 U46662 ( .A1(n47907), .A2(n44418), .ZN(n44866) );
  NAND4_X1 U46663 ( .A1(n44864), .A2(n44868), .A3(n45761), .A4(n46633), .ZN(
        n44419) );
  NAND2_X1 U46664 ( .A1(n48084), .A2(n48074), .ZN(n48053) );
  NOR2_X1 U46665 ( .A1(n48260), .A2(n48267), .ZN(n44670) );
  OR3_X1 U46666 ( .A1(n44670), .A2(n48267), .A3(n48264), .ZN(n44434) );
  OAI21_X1 U46667 ( .B1(n44431), .B2(n48436), .A(n44425), .ZN(n44428) );
  NAND2_X1 U46668 ( .A1(n48432), .A2(n44427), .ZN(n48263) );
  NAND2_X1 U46670 ( .A1(n48263), .A2(n48261), .ZN(n44426) );
  AOI21_X1 U46671 ( .B1(n44428), .B2(n44427), .A(n44426), .ZN(n44433) );
  NAND2_X1 U46672 ( .A1(n48438), .A2(n48436), .ZN(n48274) );
  OAI21_X1 U46673 ( .B1(n48264), .B2(n48273), .A(n48434), .ZN(n44429) );
  OR2_X1 U46674 ( .A1(n48274), .A2(n44429), .ZN(n44432) );
  NAND4_X1 U46675 ( .A1(n48021), .A2(n48081), .A3(n48053), .A4(n44442), .ZN(
        n44438) );
  NOR2_X1 U46676 ( .A1(n48084), .A2(n48051), .ZN(n48067) );
  OR2_X1 U46677 ( .A1(n48074), .A2(n48077), .ZN(n48032) );
  NOR2_X1 U46678 ( .A1(n48032), .A2(n52127), .ZN(n44435) );
  AND2_X1 U46679 ( .A1(n51092), .A2(n48074), .ZN(n48002) );
  AOI22_X1 U46680 ( .A1(n48067), .A2(n44435), .B1(n48021), .B2(n48002), .ZN(
        n44437) );
  NOR2_X1 U46681 ( .A1(n51343), .A2(n48077), .ZN(n48009) );
  INV_X1 U46682 ( .A(n48084), .ZN(n48039) );
  AND2_X1 U46683 ( .A1(n48009), .A2(n48039), .ZN(n44441) );
  NAND3_X1 U46684 ( .A1(n48039), .A2(n48077), .A3(n48074), .ZN(n44439) );
  NAND2_X1 U46685 ( .A1(n48069), .A2(n44439), .ZN(n44440) );
  OAI21_X1 U46686 ( .B1(n44441), .B2(n48069), .A(n44440), .ZN(n44448) );
  INV_X1 U46687 ( .A(n44442), .ZN(n48066) );
  NOR2_X1 U46688 ( .A1(n48051), .A2(n48041), .ZN(n48019) );
  NAND2_X1 U46689 ( .A1(n51092), .A2(n48039), .ZN(n48042) );
  NAND3_X1 U46690 ( .A1(n48066), .A2(n48019), .A3(n48042), .ZN(n44447) );
  AND2_X1 U46691 ( .A1(n48051), .A2(n48077), .ZN(n44443) );
  NAND3_X1 U46692 ( .A1(n48054), .A2(n44443), .A3(n48041), .ZN(n44445) );
  AND2_X1 U46693 ( .A1(n48083), .A2(n48074), .ZN(n48007) );
  AOI22_X1 U46694 ( .A1(n48007), .A2(n44443), .B1(n48002), .B2(n52127), .ZN(
        n44444) );
  INV_X1 U46695 ( .A(n4754), .ZN(n44450) );
  XNOR2_X1 U46696 ( .A(n44451), .B(n44450), .ZN(Plaintext[37]) );
  NAND2_X1 U46697 ( .A1(n47069), .A2(n7046), .ZN(n44453) );
  NOR2_X1 U46698 ( .A1(n51292), .A2(n46774), .ZN(n44459) );
  NAND2_X1 U46699 ( .A1(n44458), .A2(n44459), .ZN(n47073) );
  OAI21_X1 U46700 ( .B1(n44453), .B2(n47073), .A(n44452), .ZN(n44457) );
  OR2_X1 U46701 ( .A1(n46816), .A2(n46830), .ZN(n47080) );
  INV_X1 U46702 ( .A(n47080), .ZN(n45177) );
  NAND2_X1 U46703 ( .A1(n45177), .A2(n7046), .ZN(n44455) );
  NAND3_X1 U46704 ( .A1(n46822), .A2(n46823), .A3(n51304), .ZN(n44454) );
  NAND2_X1 U46705 ( .A1(n46772), .A2(n400), .ZN(n44461) );
  INV_X1 U46706 ( .A(n44459), .ZN(n44460) );
  OR2_X1 U46707 ( .A1(n44460), .A2(n46772), .ZN(n46782) );
  MUX2_X1 U46708 ( .A(n44461), .B(n46782), .S(n46781), .Z(n44466) );
  INV_X1 U46709 ( .A(n46775), .ZN(n44462) );
  INV_X1 U46710 ( .A(n47069), .ZN(n45172) );
  MUX2_X1 U46711 ( .A(n44464), .B(n44463), .S(n45179), .Z(n44465) );
  NAND2_X1 U46712 ( .A1(n45165), .A2(n389), .ZN(n46997) );
  OAI22_X1 U46713 ( .A1(n44473), .A2(n46997), .B1(n47152), .B2(n47153), .ZN(
        n44469) );
  INV_X1 U46714 ( .A(n44469), .ZN(n44477) );
  OR2_X1 U46715 ( .A1(n47160), .A2(n46888), .ZN(n44476) );
  INV_X1 U46716 ( .A(n47154), .ZN(n47149) );
  OR2_X1 U46717 ( .A1(n44473), .A2(n44472), .ZN(n44474) );
  NAND4_X2 U46718 ( .A1(n44475), .A2(n44476), .A3(n44477), .A4(n44474), .ZN(
        n50716) );
  XNOR2_X1 U46719 ( .A(n44479), .B(n44478), .ZN(n44481) );
  XNOR2_X1 U46720 ( .A(n44483), .B(n4526), .ZN(n44484) );
  XNOR2_X1 U46721 ( .A(n44485), .B(n44484), .ZN(n44486) );
  XNOR2_X1 U46722 ( .A(n45327), .B(n44486), .ZN(n44487) );
  XNOR2_X1 U46723 ( .A(n44951), .B(n44487), .ZN(n44488) );
  XNOR2_X1 U46724 ( .A(n44490), .B(n44489), .ZN(n44491) );
  XNOR2_X1 U46725 ( .A(n44979), .B(n51398), .ZN(n44500) );
  XNOR2_X1 U46726 ( .A(n44493), .B(n4065), .ZN(n44494) );
  XNOR2_X1 U46727 ( .A(n44495), .B(n44494), .ZN(n44496) );
  XNOR2_X1 U46728 ( .A(n44497), .B(n44496), .ZN(n44498) );
  XNOR2_X1 U46729 ( .A(n50967), .B(n44498), .ZN(n44499) );
  XNOR2_X1 U46730 ( .A(n44500), .B(n44499), .ZN(n44502) );
  XNOR2_X1 U46731 ( .A(n44501), .B(n45365), .ZN(n46140) );
  XNOR2_X1 U46732 ( .A(n44502), .B(n46140), .ZN(n44504) );
  XNOR2_X1 U46733 ( .A(n44506), .B(n4932), .ZN(n44507) );
  XNOR2_X1 U46734 ( .A(n44508), .B(n44507), .ZN(n44509) );
  XNOR2_X1 U46735 ( .A(n44510), .B(n44509), .ZN(n44511) );
  XNOR2_X1 U46736 ( .A(n44511), .B(n44900), .ZN(n44513) );
  XNOR2_X1 U46737 ( .A(n44512), .B(n44513), .ZN(n44515) );
  XNOR2_X1 U46738 ( .A(n44515), .B(n44514), .ZN(n44517) );
  XNOR2_X1 U46739 ( .A(n44516), .B(n44517), .ZN(n44519) );
  XNOR2_X1 U46740 ( .A(n44520), .B(n44521), .ZN(n44528) );
  XNOR2_X1 U46741 ( .A(n44523), .B(n44522), .ZN(n44524) );
  XNOR2_X1 U46742 ( .A(n2185), .B(n44524), .ZN(n44526) );
  XNOR2_X1 U46743 ( .A(n44525), .B(n44526), .ZN(n44527) );
  XNOR2_X1 U46744 ( .A(n44528), .B(n44527), .ZN(n44531) );
  INV_X1 U46745 ( .A(n44529), .ZN(n44530) );
  XNOR2_X1 U46746 ( .A(n44530), .B(n44531), .ZN(n44533) );
  XNOR2_X1 U46747 ( .A(n44535), .B(n44534), .ZN(n44536) );
  XNOR2_X1 U46748 ( .A(n44537), .B(n4847), .ZN(n44538) );
  XNOR2_X1 U46749 ( .A(n44539), .B(n44538), .ZN(n44540) );
  XNOR2_X1 U46750 ( .A(n44541), .B(n44540), .ZN(n44543) );
  XNOR2_X1 U46751 ( .A(n44542), .B(n44543), .ZN(n44544) );
  XNOR2_X1 U46752 ( .A(n44545), .B(n44544), .ZN(n44551) );
  XNOR2_X1 U46753 ( .A(n670), .B(n44546), .ZN(n44550) );
  XNOR2_X1 U46754 ( .A(n46058), .B(n44547), .ZN(n44549) );
  XNOR2_X1 U46755 ( .A(n44548), .B(n44549), .ZN(n44927) );
  XOR2_X1 U46756 ( .A(n4638), .B(n2117), .Z(n44554) );
  XNOR2_X1 U46757 ( .A(n44555), .B(n44554), .ZN(n44556) );
  XNOR2_X1 U46758 ( .A(n44557), .B(n44556), .ZN(n44558) );
  XNOR2_X1 U46759 ( .A(n45114), .B(n44558), .ZN(n44560) );
  XNOR2_X1 U46760 ( .A(n44560), .B(n44559), .ZN(n44564) );
  XNOR2_X1 U46761 ( .A(n44561), .B(n44562), .ZN(n44563) );
  XNOR2_X1 U46762 ( .A(n44564), .B(n44563), .ZN(n44566) );
  XNOR2_X1 U46763 ( .A(n44565), .B(n44566), .ZN(n44570) );
  XNOR2_X1 U46764 ( .A(n44567), .B(n44568), .ZN(n44569) );
  XNOR2_X1 U46765 ( .A(n44569), .B(n44570), .ZN(n44572) );
  NAND2_X1 U46766 ( .A1(n47111), .A2(n2159), .ZN(n44574) );
  NAND2_X1 U46767 ( .A1(n44574), .A2(n44573), .ZN(n44575) );
  AND2_X1 U46768 ( .A1(n46872), .A2(n47096), .ZN(n47112) );
  INV_X1 U46769 ( .A(n47088), .ZN(n47093) );
  NAND2_X1 U46771 ( .A1(n47104), .A2(n44576), .ZN(n44577) );
  AND2_X1 U46772 ( .A1(n46877), .A2(n44577), .ZN(n44579) );
  AND2_X1 U46773 ( .A1(n51410), .A2(n50280), .ZN(n47339) );
  INV_X1 U46774 ( .A(n47339), .ZN(n44581) );
  NAND2_X1 U46775 ( .A1(n44581), .A2(n50266), .ZN(n44585) );
  INV_X1 U46776 ( .A(n50259), .ZN(n44582) );
  INV_X1 U46777 ( .A(n44585), .ZN(n44587) );
  NAND3_X1 U46778 ( .A1(n44587), .A2(n44586), .A3(n50277), .ZN(n44593) );
  NAND2_X1 U46779 ( .A1(n50262), .A2(n50255), .ZN(n44588) );
  NAND2_X1 U46780 ( .A1(n44589), .A2(n44588), .ZN(n44590) );
  OR2_X1 U46781 ( .A1(n47333), .A2(n44001), .ZN(n47042) );
  NAND2_X1 U46782 ( .A1(n50276), .A2(n47044), .ZN(n44591) );
  NAND2_X1 U46783 ( .A1(n47042), .A2(n44591), .ZN(n44592) );
  NAND2_X1 U46784 ( .A1(n52126), .A2(n50679), .ZN(n44632) );
  INV_X1 U46785 ( .A(n44632), .ZN(n50667) );
  INV_X1 U46786 ( .A(n46984), .ZN(n46803) );
  NAND2_X1 U46787 ( .A1(n43798), .A2(n50367), .ZN(n46805) );
  OAI21_X1 U46788 ( .B1(n47139), .B2(n46803), .A(n46805), .ZN(n50362) );
  NAND2_X1 U46789 ( .A1(n50362), .A2(n3607), .ZN(n44598) );
  INV_X1 U46790 ( .A(n50364), .ZN(n44595) );
  INV_X1 U46791 ( .A(n50372), .ZN(n44594) );
  INV_X1 U46792 ( .A(n50363), .ZN(n46983) );
  NAND3_X1 U46793 ( .A1(n44594), .A2(n46983), .A3(n50370), .ZN(n44597) );
  AND2_X1 U46794 ( .A1(n46971), .A2(n50370), .ZN(n46975) );
  NAND3_X1 U46795 ( .A1(n44598), .A2(n44597), .A3(n44596), .ZN(n44606) );
  NOR2_X1 U46796 ( .A1(n47139), .A2(n51421), .ZN(n47145) );
  OR2_X1 U46797 ( .A1(n50364), .A2(n667), .ZN(n44601) );
  NOR2_X1 U46798 ( .A1(n50361), .A2(n44601), .ZN(n44599) );
  OAI21_X1 U46799 ( .B1(n47145), .B2(n44599), .A(n50368), .ZN(n44600) );
  AND2_X1 U46800 ( .A1(n50364), .A2(n50368), .ZN(n47144) );
  NAND3_X1 U46801 ( .A1(n47144), .A2(n3607), .A3(n51421), .ZN(n46797) );
  NOR2_X1 U46802 ( .A1(n50364), .A2(n50366), .ZN(n47137) );
  AND2_X1 U46803 ( .A1(n47137), .A2(n51421), .ZN(n44604) );
  INV_X1 U46804 ( .A(n44601), .ZN(n44602) );
  OAI211_X1 U46805 ( .C1(n44602), .C2(n50368), .A(n43798), .B(n50363), .ZN(
        n44603) );
  OAI22_X1 U46806 ( .A1(n46800), .A2(n46971), .B1(n44604), .B2(n44603), .ZN(
        n44605) );
  OAI21_X1 U46807 ( .B1(n50710), .B2(n50667), .A(n50681), .ZN(n44623) );
  NAND2_X1 U46808 ( .A1(n47026), .A2(n50343), .ZN(n50337) );
  OR2_X1 U46809 ( .A1(n44607), .A2(n50337), .ZN(n47282) );
  NAND2_X1 U46810 ( .A1(n51725), .A2(n47030), .ZN(n50342) );
  NAND2_X1 U46811 ( .A1(n47294), .A2(n47030), .ZN(n47273) );
  INV_X1 U46812 ( .A(n47273), .ZN(n44611) );
  AND2_X1 U46813 ( .A1(n47288), .A2(n505), .ZN(n47290) );
  NAND2_X1 U46814 ( .A1(n47271), .A2(n50344), .ZN(n44609) );
  NOR2_X1 U46815 ( .A1(n47290), .A2(n44609), .ZN(n44610) );
  INV_X1 U46816 ( .A(n50347), .ZN(n47028) );
  AOI22_X1 U46817 ( .A1(n44611), .A2(n44610), .B1(n49961), .B2(n47028), .ZN(
        n44620) );
  AND2_X1 U46818 ( .A1(n555), .A2(n51386), .ZN(n47289) );
  NAND2_X1 U46819 ( .A1(n50352), .A2(n47289), .ZN(n44612) );
  NAND2_X1 U46820 ( .A1(n44613), .A2(n44612), .ZN(n44618) );
  OR2_X1 U46821 ( .A1(n50337), .A2(n47030), .ZN(n44616) );
  NOR3_X1 U46822 ( .A1(n47271), .A2(n50344), .A3(n51026), .ZN(n44615) );
  NAND2_X1 U46823 ( .A1(n50335), .A2(n47030), .ZN(n44614) );
  AOI21_X1 U46824 ( .B1(n50689), .B2(n50680), .A(n51367), .ZN(n44622) );
  INV_X1 U46825 ( .A(n50681), .ZN(n50731) );
  OAI21_X1 U46826 ( .B1(n50692), .B2(n50721), .A(n50731), .ZN(n44621) );
  NAND2_X1 U46828 ( .A1(n50700), .A2(n50721), .ZN(n44625) );
  NAND2_X1 U46829 ( .A1(n50700), .A2(n50680), .ZN(n44624) );
  NAND3_X1 U46830 ( .A1(n50718), .A2(n44625), .A3(n44624), .ZN(n44627) );
  NOR2_X1 U46831 ( .A1(n50721), .A2(n50727), .ZN(n50723) );
  INV_X1 U46832 ( .A(n50679), .ZN(n50704) );
  NAND2_X1 U46833 ( .A1(n50723), .A2(n50704), .ZN(n44626) );
  NOR2_X1 U46834 ( .A1(n50727), .A2(n52126), .ZN(n50676) );
  NAND2_X1 U46835 ( .A1(n50676), .A2(n50679), .ZN(n44629) );
  AND2_X1 U46836 ( .A1(n50716), .A2(n50679), .ZN(n50726) );
  OAI21_X1 U46837 ( .B1(n50726), .B2(n50705), .A(n50727), .ZN(n44628) );
  NAND4_X1 U46838 ( .A1(n44630), .A2(n44629), .A3(n50721), .A4(n44628), .ZN(
        n44635) );
  NAND2_X1 U46839 ( .A1(n50727), .A2(n50680), .ZN(n44631) );
  NOR2_X1 U46840 ( .A1(n44632), .A2(n44631), .ZN(n44633) );
  NOR2_X1 U46841 ( .A1(n50731), .A2(n50721), .ZN(n50707) );
  NAND2_X1 U46842 ( .A1(n50716), .A2(n50708), .ZN(n50650) );
  INV_X1 U46843 ( .A(n50650), .ZN(n50655) );
  AOI22_X1 U46844 ( .A1(n44633), .A2(n50707), .B1(n50655), .B2(n51367), .ZN(
        n44634) );
  INV_X1 U46845 ( .A(n4838), .ZN(n44638) );
  AOI21_X1 U46846 ( .B1(n45820), .B2(n45819), .A(n44640), .ZN(n44642) );
  NAND3_X1 U46847 ( .A1(n45524), .A2(n45827), .A3(n44831), .ZN(n45525) );
  NAND2_X1 U46849 ( .A1(n45836), .A2(n45827), .ZN(n44815) );
  NOR2_X1 U46850 ( .A1(n45524), .A2(n44643), .ZN(n44644) );
  AOI21_X1 U46851 ( .B1(n44815), .B2(n44644), .A(n45820), .ZN(n44645) );
  NOR2_X1 U46852 ( .A1(n45533), .A2(n44827), .ZN(n45531) );
  INV_X1 U46853 ( .A(n45531), .ZN(n44650) );
  NOR2_X1 U46854 ( .A1(n44822), .A2(n44646), .ZN(n45520) );
  INV_X1 U46855 ( .A(n45520), .ZN(n44649) );
  NOR2_X1 U46856 ( .A1(n45532), .A2(n44826), .ZN(n44823) );
  NAND2_X1 U46857 ( .A1(n44823), .A2(n45521), .ZN(n44648) );
  INV_X1 U46858 ( .A(n45830), .ZN(n44817) );
  NAND4_X1 U46860 ( .A1(n44817), .A2(n45819), .A3(n45534), .A4(n44827), .ZN(
        n44647) );
  NAND4_X1 U46861 ( .A1(n44650), .A2(n44649), .A3(n44648), .A4(n44647), .ZN(
        n47891) );
  NAND2_X1 U46862 ( .A1(n45757), .A2(n47909), .ZN(n44651) );
  NAND3_X1 U46864 ( .A1(n44651), .A2(n46631), .A3(n45756), .ZN(n47913) );
  XNOR2_X1 U46865 ( .A(n46627), .B(n6741), .ZN(n44653) );
  NAND3_X1 U46866 ( .A1(n44868), .A2(n5325), .A3(n44653), .ZN(n47914) );
  NAND2_X1 U46867 ( .A1(n46628), .A2(n44654), .ZN(n47912) );
  OR2_X1 U46868 ( .A1(n46632), .A2(n46642), .ZN(n47911) );
  NAND2_X1 U46869 ( .A1(n47991), .A2(n47937), .ZN(n47925) );
  NAND3_X1 U46872 ( .A1(n48260), .A2(n48438), .A3(n2346), .ZN(n44657) );
  OAI21_X1 U46873 ( .B1(n44658), .B2(n48438), .A(n44657), .ZN(n44663) );
  OR2_X1 U46874 ( .A1(n48434), .A2(n48264), .ZN(n44666) );
  NAND3_X1 U46875 ( .A1(n44659), .A2(n44666), .A3(n48436), .ZN(n44662) );
  NAND2_X1 U46876 ( .A1(n48434), .A2(n48259), .ZN(n44660) );
  NOR2_X1 U46877 ( .A1(n52178), .A2(n44660), .ZN(n44661) );
  AOI21_X1 U46878 ( .B1(n44663), .B2(n44662), .A(n44661), .ZN(n44672) );
  AOI21_X1 U46879 ( .B1(n48423), .B2(n48437), .A(n48433), .ZN(n44664) );
  INV_X1 U46880 ( .A(n44666), .ZN(n44667) );
  AOI21_X1 U46881 ( .B1(n44667), .B2(n48438), .A(n48269), .ZN(n44668) );
  NAND2_X2 U46882 ( .A1(n44672), .A2(n44671), .ZN(n47945) );
  AOI21_X1 U46883 ( .B1(n48251), .B2(n51301), .A(n48479), .ZN(n44676) );
  NAND2_X1 U46884 ( .A1(n48478), .A2(n48248), .ZN(n44682) );
  NAND3_X1 U46885 ( .A1(n44674), .A2(n48251), .A3(n45600), .ZN(n44675) );
  OAI21_X1 U46886 ( .B1(n44676), .B2(n44682), .A(n44675), .ZN(n44677) );
  INV_X1 U46887 ( .A(n44677), .ZN(n44690) );
  NAND2_X1 U46888 ( .A1(n44679), .A2(n44678), .ZN(n44689) );
  OAI21_X1 U46889 ( .B1(n48487), .B2(n48478), .A(n48246), .ZN(n44680) );
  OR2_X1 U46890 ( .A1(n48474), .A2(n44682), .ZN(n45601) );
  AND2_X1 U46891 ( .A1(n44683), .A2(n45601), .ZN(n44688) );
  NOR2_X1 U46892 ( .A1(n48247), .A2(n48248), .ZN(n44684) );
  AND2_X1 U46893 ( .A1(n48251), .A2(n44684), .ZN(n45604) );
  OR2_X1 U46894 ( .A1(n44409), .A2(n48248), .ZN(n48477) );
  NOR2_X1 U46895 ( .A1(n44685), .A2(n48477), .ZN(n44686) );
  OAI21_X1 U46896 ( .B1(n45604), .B2(n44686), .A(n48478), .ZN(n44687) );
  OR2_X1 U46898 ( .A1(n45539), .A2(n44691), .ZN(n44700) );
  XNOR2_X1 U46899 ( .A(n52070), .B(n45538), .ZN(n44692) );
  NAND4_X1 U46900 ( .A1(n44692), .A2(n44992), .A3(n52050), .A4(n48200), .ZN(
        n44698) );
  NAND2_X1 U46901 ( .A1(n45538), .A2(n48200), .ZN(n44695) );
  NAND2_X1 U46902 ( .A1(n48205), .A2(n44992), .ZN(n45552) );
  OAI21_X1 U46903 ( .B1(n44693), .B2(n48213), .A(n45552), .ZN(n44694) );
  NAND4_X1 U46904 ( .A1(n44998), .A2(n44696), .A3(n44695), .A4(n44694), .ZN(
        n44697) );
  NAND2_X1 U46905 ( .A1(n47936), .A2(n47945), .ZN(n47965) );
  NAND2_X1 U46906 ( .A1(n47965), .A2(n51805), .ZN(n44710) );
  INV_X1 U46907 ( .A(n46705), .ZN(n46586) );
  INV_X1 U46908 ( .A(n46708), .ZN(n46583) );
  NAND2_X1 U46909 ( .A1(n46583), .A2(n46591), .ZN(n44701) );
  NOR2_X1 U46910 ( .A1(n46587), .A2(n44701), .ZN(n44702) );
  INV_X1 U46911 ( .A(n46587), .ZN(n46699) );
  NAND3_X1 U46912 ( .A1(n44704), .A2(n46714), .A3(n45790), .ZN(n44846) );
  OAI21_X1 U46913 ( .B1(n45788), .B2(n46586), .A(n44846), .ZN(n44705) );
  XNOR2_X1 U46914 ( .A(n44706), .B(n46714), .ZN(n44707) );
  NOR2_X1 U46915 ( .A1(n46580), .A2(n46587), .ZN(n46573) );
  NAND2_X1 U46916 ( .A1(n46573), .A2(n46584), .ZN(n44708) );
  NAND3_X1 U46917 ( .A1(n44710), .A2(n47988), .A3(n47966), .ZN(n44712) );
  NOR2_X1 U46918 ( .A1(n52056), .A2(n47937), .ZN(n47926) );
  NAND3_X1 U46919 ( .A1(n567), .A2(n47926), .A3(n47945), .ZN(n44711) );
  INV_X1 U46920 ( .A(n47965), .ZN(n47995) );
  AND2_X1 U46921 ( .A1(n52056), .A2(n47936), .ZN(n47974) );
  AOI22_X1 U46922 ( .A1(n567), .A2(n47995), .B1(n47974), .B2(n47941), .ZN(
        n44720) );
  NOR2_X1 U46923 ( .A1(n47989), .A2(n47936), .ZN(n47944) );
  NAND2_X1 U46924 ( .A1(n47991), .A2(n47944), .ZN(n44713) );
  NAND2_X1 U46925 ( .A1(n44713), .A2(n47990), .ZN(n44715) );
  OR2_X1 U46926 ( .A1(n47966), .A2(n52057), .ZN(n47950) );
  OAI21_X1 U46927 ( .B1(n47950), .B2(n52162), .A(n47945), .ZN(n44714) );
  NAND2_X1 U46928 ( .A1(n44715), .A2(n44714), .ZN(n44718) );
  NOR2_X1 U46929 ( .A1(n567), .A2(n47937), .ZN(n47943) );
  OAI211_X1 U46931 ( .C1(n47990), .C2(n52057), .A(n47943), .B(n44716), .ZN(
        n44717) );
  INV_X1 U46933 ( .A(n75), .ZN(n44722) );
  XNOR2_X1 U46934 ( .A(n44723), .B(n44722), .ZN(Plaintext[30]) );
  NAND2_X1 U46935 ( .A1(n44730), .A2(n46287), .ZN(n44734) );
  NOR2_X1 U46936 ( .A1(n44734), .A2(n49146), .ZN(n44724) );
  INV_X1 U46937 ( .A(n44725), .ZN(n44739) );
  AND2_X1 U46938 ( .A1(n44726), .A2(n46282), .ZN(n44729) );
  NAND2_X1 U46939 ( .A1(n49139), .A2(n43421), .ZN(n46302) );
  AND2_X1 U46942 ( .A1(n49137), .A2(n49146), .ZN(n46291) );
  AOI22_X1 U46943 ( .A1(n44729), .A2(n46302), .B1(n44728), .B2(n46291), .ZN(
        n44738) );
  INV_X1 U46944 ( .A(n44730), .ZN(n46280) );
  MUX2_X1 U46945 ( .A(n44731), .B(n46280), .S(n46287), .Z(n44732) );
  OAI21_X1 U46946 ( .B1(n44732), .B2(n45944), .A(n46292), .ZN(n44737) );
  AOI21_X1 U46947 ( .B1(n44734), .B2(n44733), .A(n49149), .ZN(n44735) );
  OAI21_X1 U46948 ( .B1(n49145), .B2(n44735), .A(n46288), .ZN(n44736) );
  INV_X1 U46949 ( .A(n49119), .ZN(n49054) );
  NOR2_X1 U46950 ( .A1(n49696), .A2(n49232), .ZN(n49237) );
  AOI21_X1 U46951 ( .B1(n49248), .B2(n49237), .A(n49252), .ZN(n49703) );
  NAND2_X1 U46952 ( .A1(n45914), .A2(n51095), .ZN(n49395) );
  OAI21_X1 U46953 ( .B1(n49242), .B2(n49689), .A(n51095), .ZN(n44740) );
  OAI21_X1 U46954 ( .B1(n656), .B2(n44740), .A(n49251), .ZN(n44741) );
  NAND3_X1 U46955 ( .A1(n45914), .A2(n656), .A3(n44743), .ZN(n49256) );
  OAI211_X1 U46956 ( .C1(n49395), .C2(n49683), .A(n44741), .B(n49256), .ZN(
        n44742) );
  NAND2_X1 U46957 ( .A1(n49397), .A2(n49231), .ZN(n45918) );
  NAND2_X1 U46958 ( .A1(n44743), .A2(n588), .ZN(n44744) );
  OAI22_X1 U46959 ( .A1(n45918), .A2(n44744), .B1(n49683), .B2(n49686), .ZN(
        n44748) );
  NAND3_X1 U46960 ( .A1(n587), .A2(n49231), .A3(n49247), .ZN(n44746) );
  OAI22_X1 U46961 ( .A1(n49233), .A2(n44746), .B1(n49688), .B2(n44745), .ZN(
        n44747) );
  NAND2_X1 U46962 ( .A1(n49054), .A2(n49127), .ZN(n49085) );
  NAND2_X1 U46963 ( .A1(n49208), .A2(n49198), .ZN(n44750) );
  NAND3_X1 U46964 ( .A1(n46226), .A2(n46214), .A3(n44750), .ZN(n44751) );
  MUX2_X1 U46965 ( .A(n44751), .B(n49207), .S(n45967), .Z(n44759) );
  OAI22_X1 U46966 ( .A1(n49203), .A2(n44753), .B1(n52105), .B2(n44752), .ZN(
        n44754) );
  NAND2_X1 U46967 ( .A1(n44754), .A2(n49197), .ZN(n44758) );
  NAND3_X1 U46968 ( .A1(n46229), .A2(n49208), .A3(n45970), .ZN(n44757) );
  NAND2_X1 U46969 ( .A1(n49216), .A2(n49207), .ZN(n45968) );
  INV_X1 U46970 ( .A(n46226), .ZN(n44755) );
  NAND3_X1 U46971 ( .A1(n45968), .A2(n44755), .A3(n45969), .ZN(n44756) );
  NOR2_X1 U46973 ( .A1(n45686), .A2(n45231), .ZN(n45245) );
  AND2_X1 U46975 ( .A1(n44761), .A2(n44760), .ZN(n44771) );
  NAND2_X1 U46976 ( .A1(n45232), .A2(n46353), .ZN(n44763) );
  OAI22_X1 U46977 ( .A1(n46277), .A2(n52187), .B1(n46358), .B2(n46342), .ZN(
        n44762) );
  NAND3_X1 U46978 ( .A1(n44763), .A2(n46274), .A3(n44762), .ZN(n44770) );
  INV_X1 U46979 ( .A(n46277), .ZN(n44764) );
  AOI22_X1 U46980 ( .A1(n45245), .A2(n44764), .B1(n46355), .B2(n46342), .ZN(
        n44769) );
  NAND2_X1 U46981 ( .A1(n45697), .A2(n46354), .ZN(n45229) );
  OAI21_X1 U46982 ( .B1(n46359), .B2(n46345), .A(n45229), .ZN(n44767) );
  NAND3_X1 U46983 ( .A1(n44767), .A2(n46269), .A3(n44766), .ZN(n44768) );
  NAND4_X2 U46984 ( .A1(n44769), .A2(n44771), .A3(n44770), .A4(n44768), .ZN(
        n49117) );
  INV_X1 U46985 ( .A(n49117), .ZN(n44772) );
  NOR2_X1 U46986 ( .A1(n49267), .A2(n49272), .ZN(n45927) );
  AND3_X1 U46987 ( .A1(n51335), .A2(n49277), .A3(n49278), .ZN(n44773) );
  NOR2_X1 U46988 ( .A1(n45927), .A2(n44773), .ZN(n44782) );
  AND2_X1 U46989 ( .A1(n49266), .A2(n52086), .ZN(n45675) );
  NAND3_X1 U46990 ( .A1(n45675), .A2(n49265), .A3(n46203), .ZN(n44774) );
  NAND2_X1 U46991 ( .A1(n45665), .A2(n44774), .ZN(n44777) );
  XNOR2_X1 U46994 ( .A(n49274), .B(n49272), .ZN(n44778) );
  NAND3_X1 U46995 ( .A1(n44779), .A2(n46203), .A3(n44778), .ZN(n44781) );
  NAND2_X1 U46996 ( .A1(n46255), .A2(n49161), .ZN(n46250) );
  AND2_X1 U46997 ( .A1(n46250), .A2(n44783), .ZN(n44788) );
  NOR2_X1 U46998 ( .A1(n46243), .A2(n540), .ZN(n46256) );
  OAI21_X1 U46999 ( .B1(n49168), .B2(n44784), .A(n49162), .ZN(n44785) );
  OAI21_X1 U47000 ( .B1(n44788), .B2(n46256), .A(n44785), .ZN(n44791) );
  AND2_X1 U47001 ( .A1(n45649), .A2(n49162), .ZN(n49171) );
  NAND3_X1 U47002 ( .A1(n46258), .A2(n49171), .A3(n49170), .ZN(n44790) );
  AOI21_X1 U47003 ( .B1(n46244), .B2(n46249), .A(n664), .ZN(n44787) );
  AND2_X1 U47004 ( .A1(n539), .A2(n46255), .ZN(n49165) );
  OAI21_X1 U47005 ( .B1(n44788), .B2(n44787), .A(n49165), .ZN(n44789) );
  NAND2_X1 U47007 ( .A1(n44798), .A2(n49112), .ZN(n49104) );
  INV_X1 U47008 ( .A(n49104), .ZN(n44793) );
  INV_X1 U47009 ( .A(n49128), .ZN(n44792) );
  NAND4_X1 U47011 ( .A1(n44793), .A2(n49127), .A3(n44792), .A4(n49107), .ZN(
        n44796) );
  INV_X1 U47012 ( .A(n49126), .ZN(n44800) );
  OR2_X1 U47013 ( .A1(n49117), .A2(n49070), .ZN(n49100) );
  NOR2_X1 U47014 ( .A1(n49112), .A2(n49117), .ZN(n49068) );
  AOI21_X1 U47015 ( .B1(n49083), .B2(n49100), .A(n49068), .ZN(n44794) );
  NAND2_X1 U47016 ( .A1(n49119), .A2(n49126), .ZN(n49103) );
  NAND2_X1 U47017 ( .A1(n49103), .A2(n49127), .ZN(n49072) );
  NAND3_X1 U47018 ( .A1(n44794), .A2(n49072), .A3(n49107), .ZN(n44795) );
  INV_X1 U47019 ( .A(n44798), .ZN(n49094) );
  NAND2_X1 U47020 ( .A1(n49094), .A2(n49119), .ZN(n44799) );
  NAND2_X1 U47021 ( .A1(n49089), .A2(n49066), .ZN(n49124) );
  AND2_X1 U47022 ( .A1(n49119), .A2(n44772), .ZN(n49080) );
  NAND3_X1 U47023 ( .A1(n49065), .A2(n44800), .A3(n49080), .ZN(n44805) );
  NOR2_X1 U47024 ( .A1(n49119), .A2(n1501), .ZN(n44801) );
  NAND3_X1 U47025 ( .A1(n44801), .A2(n49126), .A3(n49112), .ZN(n44803) );
  NAND2_X1 U47026 ( .A1(n44808), .A2(n44807), .ZN(n44810) );
  INV_X1 U47027 ( .A(n4865), .ZN(n44809) );
  XNOR2_X1 U47028 ( .A(n44810), .B(n44809), .ZN(Plaintext[97]) );
  INV_X1 U47029 ( .A(n45533), .ZN(n45817) );
  NAND3_X1 U47030 ( .A1(n44811), .A2(n45817), .A3(n45523), .ZN(n45825) );
  NAND3_X1 U47031 ( .A1(n44817), .A2(n45524), .A3(n45828), .ZN(n44812) );
  AND2_X1 U47032 ( .A1(n44812), .A2(n45825), .ZN(n44821) );
  OR2_X1 U47033 ( .A1(n44814), .A2(n44813), .ZN(n44820) );
  AND2_X1 U47034 ( .A1(n44828), .A2(n44831), .ZN(n45821) );
  NAND2_X1 U47035 ( .A1(n44816), .A2(n45821), .ZN(n44819) );
  OAI211_X1 U47036 ( .C1(n45531), .C2(n45836), .A(n44817), .B(n113), .ZN(
        n44818) );
  INV_X1 U47037 ( .A(n44826), .ZN(n45816) );
  MUX2_X1 U47039 ( .A(n44827), .B(n44826), .S(n44825), .Z(n44829) );
  NAND2_X1 U47040 ( .A1(n44829), .A2(n44828), .ZN(n44830) );
  AOI22_X1 U47041 ( .A1(n44832), .A2(n44831), .B1(n44830), .B2(n45521), .ZN(
        n44833) );
  NOR2_X1 U47042 ( .A1(n46574), .A2(n51396), .ZN(n44837) );
  NAND2_X1 U47043 ( .A1(n46589), .A2(n46591), .ZN(n46713) );
  INV_X1 U47044 ( .A(n46713), .ZN(n44838) );
  OAI211_X1 U47045 ( .C1(n405), .C2(n46580), .A(n44840), .B(n44839), .ZN(
        n44841) );
  INV_X1 U47046 ( .A(n46584), .ZN(n44842) );
  INV_X1 U47047 ( .A(n46707), .ZN(n44843) );
  NAND3_X1 U47048 ( .A1(n44845), .A2(n46587), .A3(n46575), .ZN(n44847) );
  AND2_X1 U47049 ( .A1(n44847), .A2(n44846), .ZN(n44848) );
  NAND2_X1 U47050 ( .A1(n45877), .A2(n47786), .ZN(n47781) );
  OR2_X1 U47051 ( .A1(n46730), .A2(n51344), .ZN(n45802) );
  NAND3_X1 U47052 ( .A1(n45802), .A2(n2092), .A3(n46747), .ZN(n44851) );
  NAND2_X1 U47053 ( .A1(n44851), .A2(n44850), .ZN(n44855) );
  NAND2_X1 U47054 ( .A1(n46755), .A2(n51488), .ZN(n45801) );
  INV_X1 U47056 ( .A(n45190), .ZN(n44852) );
  NAND2_X1 U47057 ( .A1(n44853), .A2(n44852), .ZN(n44854) );
  NAND2_X1 U47059 ( .A1(n46738), .A2(n45188), .ZN(n44856) );
  AND2_X1 U47060 ( .A1(n44857), .A2(n44856), .ZN(n44862) );
  XNOR2_X1 U47061 ( .A(n51344), .B(n46730), .ZN(n44858) );
  NAND2_X1 U47062 ( .A1(n44858), .A2(n51488), .ZN(n46561) );
  INV_X1 U47063 ( .A(n46747), .ZN(n46560) );
  NAND4_X1 U47064 ( .A1(n46561), .A2(n46753), .A3(n46740), .A4(n46560), .ZN(
        n44861) );
  AND2_X1 U47065 ( .A1(n46755), .A2(n41723), .ZN(n44859) );
  OAI21_X1 U47066 ( .B1(n46739), .B2(n44859), .A(n46743), .ZN(n44860) );
  AND2_X1 U47067 ( .A1(n44864), .A2(n44654), .ZN(n46629) );
  NAND3_X1 U47068 ( .A1(n44866), .A2(n46629), .A3(n44865), .ZN(n44876) );
  AOI22_X1 U47069 ( .A1(n44867), .A2(n46623), .B1(n46635), .B2(n44873), .ZN(
        n44875) );
  INV_X1 U47070 ( .A(n44868), .ZN(n44870) );
  AND2_X1 U47071 ( .A1(n46628), .A2(n6741), .ZN(n44871) );
  OAI211_X1 U47072 ( .C1(n46635), .C2(n44873), .A(n44872), .B(n46632), .ZN(
        n44874) );
  NAND2_X1 U47073 ( .A1(n47763), .A2(n47745), .ZN(n45008) );
  XNOR2_X1 U47074 ( .A(n44878), .B(n44877), .ZN(n44883) );
  XNOR2_X1 U47075 ( .A(n44879), .B(n46112), .ZN(n44881) );
  XNOR2_X1 U47076 ( .A(n44881), .B(n44880), .ZN(n44882) );
  XNOR2_X1 U47077 ( .A(n44883), .B(n44882), .ZN(n44884) );
  XNOR2_X1 U47078 ( .A(n45281), .B(n44884), .ZN(n44898) );
  XNOR2_X1 U47079 ( .A(n46122), .B(n44885), .ZN(n44886) );
  XNOR2_X1 U47080 ( .A(n44887), .B(n44886), .ZN(n44888) );
  XNOR2_X1 U47081 ( .A(n44889), .B(n44888), .ZN(n44890) );
  XNOR2_X1 U47082 ( .A(n51101), .B(n44890), .ZN(n44892) );
  XNOR2_X1 U47083 ( .A(n44892), .B(n51681), .ZN(n44894) );
  XNOR2_X1 U47084 ( .A(n44893), .B(n44894), .ZN(n44896) );
  XNOR2_X1 U47085 ( .A(n44896), .B(n44895), .ZN(n44897) );
  XNOR2_X1 U47086 ( .A(n51371), .B(n44900), .ZN(n44902) );
  XNOR2_X1 U47087 ( .A(n44901), .B(n44902), .ZN(n45043) );
  XNOR2_X1 U47088 ( .A(n44903), .B(n45043), .ZN(n44916) );
  XNOR2_X1 U47089 ( .A(n44905), .B(n44904), .ZN(n46104) );
  XNOR2_X1 U47090 ( .A(n44907), .B(n44906), .ZN(n44908) );
  XNOR2_X1 U47091 ( .A(n44909), .B(n44908), .ZN(n44910) );
  XNOR2_X1 U47092 ( .A(n44911), .B(n44910), .ZN(n44912) );
  XNOR2_X1 U47093 ( .A(n44913), .B(n44912), .ZN(n44914) );
  XNOR2_X1 U47094 ( .A(n46104), .B(n44914), .ZN(n44915) );
  XNOR2_X1 U47095 ( .A(n44916), .B(n44915), .ZN(n44918) );
  INV_X1 U47096 ( .A(n4880), .ZN(n50056) );
  XNOR2_X1 U47097 ( .A(n44919), .B(n50056), .ZN(n44920) );
  XNOR2_X1 U47098 ( .A(n44921), .B(n44920), .ZN(n44922) );
  XNOR2_X1 U47099 ( .A(n45426), .B(n44922), .ZN(n44924) );
  XNOR2_X1 U47100 ( .A(n44924), .B(n44923), .ZN(n44926) );
  XNOR2_X1 U47101 ( .A(n670), .B(n44926), .ZN(n44928) );
  XNOR2_X1 U47102 ( .A(n44928), .B(n44927), .ZN(n44930) );
  XNOR2_X1 U47103 ( .A(n44933), .B(n44932), .ZN(n44943) );
  XNOR2_X1 U47104 ( .A(n44935), .B(n2608), .ZN(n44936) );
  XNOR2_X1 U47105 ( .A(n44937), .B(n44936), .ZN(n44939) );
  XNOR2_X1 U47106 ( .A(n44939), .B(n50987), .ZN(n44941) );
  XNOR2_X1 U47107 ( .A(n44941), .B(n44940), .ZN(n44942) );
  XNOR2_X1 U47108 ( .A(n44943), .B(n44942), .ZN(n44948) );
  XNOR2_X1 U47109 ( .A(n44945), .B(n44944), .ZN(n44946) );
  XNOR2_X1 U47110 ( .A(n45321), .B(n44946), .ZN(n44947) );
  XNOR2_X1 U47111 ( .A(n44947), .B(n44948), .ZN(n44950) );
  AND2_X1 U47112 ( .A1(n46901), .A2(n46614), .ZN(n46920) );
  XNOR2_X1 U47113 ( .A(n51294), .B(n44951), .ZN(n44959) );
  XNOR2_X1 U47114 ( .A(n44952), .B(n4676), .ZN(n44953) );
  XNOR2_X1 U47115 ( .A(n44954), .B(n44953), .ZN(n44955) );
  XNOR2_X1 U47116 ( .A(n44956), .B(n44955), .ZN(n44957) );
  XNOR2_X1 U47117 ( .A(n45484), .B(n44957), .ZN(n44958) );
  XNOR2_X1 U47118 ( .A(n44959), .B(n44958), .ZN(n44961) );
  XOR2_X1 U47119 ( .A(n44963), .B(n44962), .Z(n44965) );
  XNOR2_X1 U47120 ( .A(n44965), .B(n44964), .ZN(n44966) );
  XNOR2_X1 U47121 ( .A(n44968), .B(n44967), .ZN(n44970) );
  XNOR2_X1 U47123 ( .A(n569), .B(n44971), .ZN(n44974) );
  XNOR2_X1 U47124 ( .A(n44977), .B(n44976), .ZN(n44978) );
  XNOR2_X1 U47125 ( .A(n44979), .B(n44978), .ZN(n44981) );
  INV_X1 U47126 ( .A(n45089), .ZN(n44980) );
  XNOR2_X1 U47127 ( .A(n44981), .B(n44980), .ZN(n44982) );
  XNOR2_X1 U47128 ( .A(n44982), .B(n51368), .ZN(n44984) );
  INV_X1 U47129 ( .A(n44985), .ZN(n46905) );
  INV_X1 U47130 ( .A(n46692), .ZN(n44986) );
  NAND3_X1 U47131 ( .A1(n46905), .A2(n46693), .A3(n45848), .ZN(n44987) );
  NAND2_X1 U47132 ( .A1(n46905), .A2(n51359), .ZN(n45031) );
  NAND2_X1 U47133 ( .A1(n44987), .A2(n45031), .ZN(n44988) );
  OAI21_X1 U47134 ( .B1(n46901), .B2(n45848), .A(n46913), .ZN(n44989) );
  INV_X1 U47135 ( .A(n48208), .ZN(n44995) );
  NAND2_X1 U47136 ( .A1(n44990), .A2(n48205), .ZN(n44991) );
  AOI21_X1 U47137 ( .B1(n52161), .B2(n45538), .A(n44991), .ZN(n44994) );
  OR2_X1 U47138 ( .A1(n45542), .A2(n44992), .ZN(n44993) );
  AOI22_X1 U47139 ( .A1(n44995), .A2(n48210), .B1(n44994), .B2(n44993), .ZN(
        n45006) );
  INV_X1 U47140 ( .A(n48210), .ZN(n45549) );
  INV_X1 U47141 ( .A(n45547), .ZN(n48216) );
  OAI211_X1 U47142 ( .C1(n45549), .C2(n48216), .A(n45539), .B(n2119), .ZN(
        n45001) );
  INV_X1 U47143 ( .A(n45552), .ZN(n48220) );
  NAND2_X1 U47144 ( .A1(n44996), .A2(n48200), .ZN(n44997) );
  NAND2_X1 U47145 ( .A1(n45002), .A2(n45545), .ZN(n48212) );
  INV_X1 U47146 ( .A(n45554), .ZN(n45003) );
  NAND2_X1 U47147 ( .A1(n45003), .A2(n48207), .ZN(n45004) );
  AND2_X1 U47148 ( .A1(n47745), .A2(n47777), .ZN(n47755) );
  OAI211_X1 U47149 ( .C1(n47781), .C2(n45008), .A(n47785), .B(n45007), .ZN(
        n45010) );
  INV_X1 U47150 ( .A(n47744), .ZN(n47730) );
  NOR2_X1 U47151 ( .A1(n45010), .A2(n45009), .ZN(n45019) );
  NAND2_X1 U47152 ( .A1(n47797), .A2(n51468), .ZN(n47766) );
  OAI211_X1 U47153 ( .C1(n47777), .C2(n47766), .A(n45011), .B(n45877), .ZN(
        n45014) );
  NAND3_X1 U47154 ( .A1(n47711), .A2(n47790), .A3(n47745), .ZN(n45012) );
  AOI21_X1 U47155 ( .B1(n45012), .B2(n52149), .A(n47786), .ZN(n45013) );
  NAND2_X1 U47156 ( .A1(n45014), .A2(n45013), .ZN(n45018) );
  XNOR2_X1 U47157 ( .A(n47763), .B(n51467), .ZN(n47760) );
  NOR2_X1 U47158 ( .A1(n47745), .A2(n47777), .ZN(n47716) );
  NAND4_X1 U47159 ( .A1(n47760), .A2(n47716), .A3(n47786), .A4(n47782), .ZN(
        n45017) );
  OR2_X1 U47160 ( .A1(n47771), .A2(n47786), .ZN(n47710) );
  OAI21_X1 U47161 ( .B1(n47710), .B2(n47711), .A(n47742), .ZN(n45015) );
  INV_X1 U47162 ( .A(n45015), .ZN(n45016) );
  INV_X1 U47163 ( .A(n4429), .ZN(n45020) );
  NAND2_X1 U47164 ( .A1(n49521), .A2(n49511), .ZN(n49538) );
  NAND2_X1 U47165 ( .A1(n49534), .A2(n49539), .ZN(n49494) );
  NAND2_X1 U47166 ( .A1(n49510), .A2(n49511), .ZN(n49495) );
  NAND2_X1 U47167 ( .A1(n49495), .A2(n51395), .ZN(n45025) );
  OR2_X1 U47168 ( .A1(n49534), .A2(n43490), .ZN(n49479) );
  AOI21_X1 U47169 ( .B1(n49479), .B2(n49529), .A(n49512), .ZN(n45026) );
  INV_X1 U47170 ( .A(n4721), .ZN(n45027) );
  INV_X1 U47171 ( .A(n46913), .ZN(n45845) );
  AND2_X1 U47172 ( .A1(n45848), .A2(n46904), .ZN(n46902) );
  INV_X1 U47173 ( .A(n46902), .ZN(n46616) );
  NAND3_X1 U47174 ( .A1(n45845), .A2(n46919), .A3(n46616), .ZN(n46910) );
  NAND3_X1 U47175 ( .A1(n46694), .A2(n46692), .A3(n46901), .ZN(n45030) );
  NAND3_X1 U47176 ( .A1(n46920), .A2(n46689), .A3(n46606), .ZN(n45029) );
  NAND3_X1 U47177 ( .A1(n46919), .A2(n46913), .A3(n46606), .ZN(n45028) );
  INV_X1 U47178 ( .A(n46912), .ZN(n46613) );
  NOR2_X1 U47179 ( .A1(n46613), .A2(n45848), .ZN(n45032) );
  OAI21_X1 U47180 ( .B1(n46915), .B2(n45032), .A(n46689), .ZN(n45036) );
  MUX2_X1 U47181 ( .A(n659), .B(n52169), .S(n46903), .Z(n45034) );
  OAI21_X1 U47182 ( .B1(n45034), .B2(n51399), .A(n46607), .ZN(n45035) );
  INV_X1 U47183 ( .A(n45192), .ZN(n50929) );
  XNOR2_X1 U47184 ( .A(n45044), .B(n45043), .ZN(n45046) );
  XNOR2_X1 U47185 ( .A(n45046), .B(n45045), .ZN(n45048) );
  XNOR2_X1 U47186 ( .A(n45048), .B(n45047), .ZN(n45138) );
  XNOR2_X1 U47188 ( .A(n45051), .B(n2604), .ZN(n45053) );
  XOR2_X1 U47189 ( .A(n45053), .B(n45052), .Z(n45054) );
  XNOR2_X1 U47190 ( .A(n45055), .B(n45054), .ZN(n45056) );
  XNOR2_X1 U47191 ( .A(n51101), .B(n45056), .ZN(n45058) );
  XNOR2_X1 U47192 ( .A(n45058), .B(n45057), .ZN(n45060) );
  XNOR2_X1 U47193 ( .A(n45060), .B(n45059), .ZN(n45061) );
  XNOR2_X1 U47194 ( .A(n45062), .B(n45061), .ZN(n45064) );
  XNOR2_X1 U47195 ( .A(n45064), .B(n45063), .ZN(n45065) );
  INV_X1 U47196 ( .A(n45065), .ZN(n45772) );
  INV_X1 U47197 ( .A(n46859), .ZN(n45066) );
  XNOR2_X1 U47199 ( .A(n45067), .B(n45068), .ZN(n45069) );
  XNOR2_X1 U47200 ( .A(n45070), .B(n45069), .ZN(n45080) );
  XOR2_X1 U47201 ( .A(n45072), .B(n45071), .Z(n45073) );
  XNOR2_X1 U47202 ( .A(n51294), .B(n45073), .ZN(n45075) );
  XNOR2_X1 U47203 ( .A(n45076), .B(n45075), .ZN(n45077) );
  XNOR2_X1 U47204 ( .A(n45078), .B(n45077), .ZN(n45079) );
  XNOR2_X1 U47205 ( .A(n45080), .B(n45079), .ZN(n45081) );
  XNOR2_X1 U47206 ( .A(n45083), .B(n45082), .ZN(n45084) );
  XNOR2_X1 U47207 ( .A(n45085), .B(n45084), .ZN(n45086) );
  XNOR2_X1 U47208 ( .A(n45087), .B(n45086), .ZN(n45088) );
  XNOR2_X1 U47209 ( .A(n45089), .B(n45088), .ZN(n45090) );
  XNOR2_X1 U47210 ( .A(n52123), .B(n45092), .ZN(n45094) );
  XNOR2_X1 U47211 ( .A(n45094), .B(n45093), .ZN(n45096) );
  XNOR2_X1 U47212 ( .A(n45095), .B(n45096), .ZN(n46649) );
  INV_X1 U47213 ( .A(n46649), .ZN(n47127) );
  NAND2_X1 U47214 ( .A1(n46842), .A2(n47127), .ZN(n46845) );
  XNOR2_X1 U47215 ( .A(n45305), .B(n45097), .ZN(n45098) );
  XNOR2_X1 U47216 ( .A(n45099), .B(n45098), .ZN(n45103) );
  XNOR2_X1 U47217 ( .A(n52043), .B(n45100), .ZN(n45102) );
  XNOR2_X1 U47218 ( .A(n45102), .B(n45103), .ZN(n45119) );
  XNOR2_X1 U47219 ( .A(n45105), .B(n45104), .ZN(n45110) );
  XNOR2_X1 U47220 ( .A(n45106), .B(n4793), .ZN(n45108) );
  XNOR2_X1 U47221 ( .A(n45108), .B(n45107), .ZN(n45109) );
  XNOR2_X1 U47222 ( .A(n45110), .B(n45109), .ZN(n45112) );
  XNOR2_X1 U47223 ( .A(n45112), .B(n45111), .ZN(n45113) );
  XNOR2_X1 U47224 ( .A(n45114), .B(n45113), .ZN(n45115) );
  XNOR2_X1 U47225 ( .A(n45116), .B(n45115), .ZN(n45117) );
  XNOR2_X1 U47226 ( .A(n45117), .B(n46052), .ZN(n45118) );
  XNOR2_X1 U47227 ( .A(n45119), .B(n45118), .ZN(n45121) );
  XNOR2_X1 U47228 ( .A(n45120), .B(n45121), .ZN(n46844) );
  INV_X1 U47229 ( .A(n47121), .ZN(n45139) );
  XNOR2_X1 U47230 ( .A(n45123), .B(n50586), .ZN(n45124) );
  XNOR2_X1 U47231 ( .A(n45125), .B(n45124), .ZN(n45126) );
  XNOR2_X1 U47232 ( .A(n45426), .B(n45126), .ZN(n45128) );
  XNOR2_X1 U47233 ( .A(n671), .B(n45128), .ZN(n45129) );
  XNOR2_X1 U47234 ( .A(n45130), .B(n45129), .ZN(n45131) );
  XNOR2_X1 U47235 ( .A(n45131), .B(n45132), .ZN(n45134) );
  XNOR2_X1 U47236 ( .A(n45134), .B(n45133), .ZN(n45135) );
  INV_X1 U47237 ( .A(n45771), .ZN(n47126) );
  NAND3_X1 U47238 ( .A1(n45139), .A2(n46840), .A3(n47126), .ZN(n46857) );
  NOR2_X1 U47239 ( .A1(n47127), .A2(n47122), .ZN(n45137) );
  INV_X1 U47240 ( .A(n46648), .ZN(n45773) );
  AND2_X1 U47241 ( .A1(n46860), .A2(n47127), .ZN(n46839) );
  NAND2_X1 U47242 ( .A1(n46839), .A2(n47118), .ZN(n45140) );
  NAND2_X1 U47243 ( .A1(n50929), .A2(n50950), .ZN(n45170) );
  NOR2_X1 U47244 ( .A1(n47095), .A2(n47088), .ZN(n47086) );
  INV_X1 U47245 ( .A(n47086), .ZN(n45142) );
  INV_X1 U47246 ( .A(n45143), .ZN(n45152) );
  INV_X1 U47247 ( .A(n47104), .ZN(n45144) );
  NAND2_X1 U47248 ( .A1(n47110), .A2(n46872), .ZN(n46725) );
  NAND2_X1 U47249 ( .A1(n45146), .A2(n47111), .ZN(n45150) );
  INV_X1 U47250 ( .A(n47098), .ZN(n45147) );
  NOR2_X1 U47251 ( .A1(n45147), .A2(n47109), .ZN(n46871) );
  INV_X1 U47252 ( .A(n47109), .ZN(n46875) );
  OR2_X1 U47253 ( .A1(n47096), .A2(n46869), .ZN(n46873) );
  OAI22_X1 U47254 ( .A1(n46875), .A2(n46873), .B1(n47108), .B2(n47111), .ZN(
        n45148) );
  OAI21_X1 U47255 ( .B1(n46871), .B2(n45148), .A(n46872), .ZN(n45149) );
  NAND2_X1 U47257 ( .A1(n47153), .A2(n47151), .ZN(n45161) );
  NOR2_X1 U47258 ( .A1(n45156), .A2(n45159), .ZN(n47156) );
  AOI21_X1 U47259 ( .B1(n45157), .B2(n2751), .A(n47156), .ZN(n47010) );
  INV_X1 U47260 ( .A(n45158), .ZN(n45163) );
  NAND2_X1 U47261 ( .A1(n46998), .A2(n46999), .ZN(n45160) );
  NAND2_X1 U47262 ( .A1(n45160), .A2(n45159), .ZN(n45162) );
  INV_X1 U47263 ( .A(n45161), .ZN(n47006) );
  AOI22_X1 U47264 ( .A1(n45163), .A2(n45162), .B1(n47006), .B2(n47154), .ZN(
        n45168) );
  NOR2_X1 U47265 ( .A1(n45164), .A2(n46888), .ZN(n47164) );
  AND2_X1 U47266 ( .A1(n45165), .A2(n47000), .ZN(n45166) );
  OAI21_X1 U47267 ( .B1(n47164), .B2(n45166), .A(n47162), .ZN(n45167) );
  BUF_X2 U47268 ( .A(n45194), .Z(n50955) );
  OR2_X1 U47269 ( .A1(n51298), .A2(n45194), .ZN(n47399) );
  NOR2_X1 U47270 ( .A1(n45170), .A2(n47399), .ZN(n50917) );
  OR2_X1 U47271 ( .A1(n47074), .A2(n51404), .ZN(n46817) );
  NAND3_X1 U47272 ( .A1(n46817), .A2(n47076), .A3(n45179), .ZN(n45171) );
  INV_X1 U47273 ( .A(n47075), .ZN(n46811) );
  NAND3_X1 U47274 ( .A1(n45171), .A2(n46811), .A3(n46812), .ZN(n45175) );
  AOI22_X1 U47275 ( .A1(n45172), .A2(n46824), .B1(n399), .B2(n51456), .ZN(
        n45174) );
  INV_X1 U47276 ( .A(n45176), .ZN(n45178) );
  NAND3_X1 U47277 ( .A1(n45178), .A2(n7046), .A3(n45177), .ZN(n45180) );
  MUX2_X1 U47278 ( .A(n46813), .B(n45180), .S(n45179), .Z(n45181) );
  NAND2_X1 U47279 ( .A1(n46747), .A2(n46554), .ZN(n45183) );
  AND2_X1 U47280 ( .A1(n46755), .A2(n50965), .ZN(n46749) );
  NAND2_X1 U47282 ( .A1(n45186), .A2(n51488), .ZN(n45187) );
  NAND3_X1 U47283 ( .A1(n45189), .A2(n45188), .A3(n45187), .ZN(n45809) );
  NAND3_X1 U47284 ( .A1(n46738), .A2(n46744), .A3(n45190), .ZN(n46733) );
  NAND2_X1 U47285 ( .A1(n50950), .A2(n50906), .ZN(n47228) );
  NAND2_X1 U47286 ( .A1(n50955), .A2(n51299), .ZN(n45193) );
  NAND2_X1 U47287 ( .A1(n47228), .A2(n45193), .ZN(n47392) );
  INV_X1 U47288 ( .A(n45194), .ZN(n50928) );
  OAI21_X1 U47289 ( .B1(n50928), .B2(n50929), .A(n47236), .ZN(n45195) );
  AOI22_X1 U47290 ( .A1(n50917), .A2(n50901), .B1(n47392), .B2(n45195), .ZN(
        n45200) );
  INV_X1 U47292 ( .A(n47396), .ZN(n45196) );
  NAND2_X1 U47293 ( .A1(n50909), .A2(n45196), .ZN(n45199) );
  INV_X1 U47294 ( .A(n50949), .ZN(n47230) );
  AND2_X1 U47295 ( .A1(n50913), .A2(n51299), .ZN(n50959) );
  NAND3_X1 U47296 ( .A1(n47230), .A2(n50959), .A3(n50929), .ZN(n45198) );
  NAND2_X1 U47297 ( .A1(n51299), .A2(n5365), .ZN(n50946) );
  INV_X1 U47298 ( .A(n50946), .ZN(n45197) );
  NAND2_X1 U47299 ( .A1(n45197), .A2(n50949), .ZN(n50910) );
  NAND3_X1 U47300 ( .A1(n45200), .A2(n45199), .A3(n8767), .ZN(n45202) );
  INV_X1 U47301 ( .A(Key[190]), .ZN(n45201) );
  XNOR2_X1 U47302 ( .A(n45202), .B(n45201), .ZN(Plaintext[190]) );
  MUX2_X1 U47304 ( .A(n48457), .B(n48450), .S(n48463), .Z(n45204) );
  NAND2_X1 U47305 ( .A1(n51732), .A2(n48459), .ZN(n45203) );
  NAND2_X1 U47306 ( .A1(n8585), .A2(n48455), .ZN(n45205) );
  MUX2_X1 U47307 ( .A(n46412), .B(n48455), .S(n7275), .Z(n45208) );
  AOI21_X1 U47308 ( .B1(n48449), .B2(n46441), .A(n46434), .ZN(n45206) );
  NOR2_X1 U47309 ( .A1(n46258), .A2(n45215), .ZN(n45210) );
  INV_X1 U47310 ( .A(n45649), .ZN(n45212) );
  OR2_X1 U47311 ( .A1(n46255), .A2(n540), .ZN(n49158) );
  OR2_X1 U47312 ( .A1(n46244), .A2(n46255), .ZN(n49157) );
  OAI21_X1 U47313 ( .B1(n45212), .B2(n49158), .A(n49157), .ZN(n45647) );
  OAI21_X1 U47314 ( .B1(n49159), .B2(n539), .A(n45647), .ZN(n45213) );
  NAND2_X1 U47315 ( .A1(n49178), .A2(n45216), .ZN(n45217) );
  AND2_X1 U47316 ( .A1(n45649), .A2(n49170), .ZN(n46239) );
  NAND3_X1 U47317 ( .A1(n46239), .A2(n49165), .A3(n46249), .ZN(n49181) );
  NAND2_X1 U47318 ( .A1(n46505), .A2(n45661), .ZN(n45218) );
  AOI21_X1 U47319 ( .B1(n51426), .B2(n46491), .A(n46488), .ZN(n45220) );
  NAND2_X1 U47320 ( .A1(n45221), .A2(n46501), .ZN(n45226) );
  NAND3_X1 U47321 ( .A1(n46502), .A2(n46487), .A3(n46385), .ZN(n45225) );
  AND2_X1 U47322 ( .A1(n8207), .A2(n52136), .ZN(n46483) );
  INV_X1 U47323 ( .A(n46483), .ZN(n45222) );
  NAND3_X1 U47324 ( .A1(n45222), .A2(n46503), .A3(n46494), .ZN(n45224) );
  NAND2_X1 U47325 ( .A1(n46488), .A2(n51426), .ZN(n45223) );
  NAND4_X1 U47326 ( .A1(n45226), .A2(n45225), .A3(n45224), .A4(n45223), .ZN(
        n45227) );
  NOR2_X1 U47327 ( .A1(n46267), .A2(n46359), .ZN(n45230) );
  AOI21_X1 U47328 ( .B1(n45230), .B2(n45229), .A(n45238), .ZN(n45695) );
  NAND2_X1 U47329 ( .A1(n46344), .A2(n46357), .ZN(n45696) );
  NAND2_X1 U47330 ( .A1(n45695), .A2(n45696), .ZN(n45236) );
  INV_X1 U47331 ( .A(n45231), .ZN(n46343) );
  NAND2_X1 U47332 ( .A1(n46355), .A2(n46343), .ZN(n45234) );
  NAND2_X1 U47333 ( .A1(n46344), .A2(n45237), .ZN(n45233) );
  NAND4_X1 U47334 ( .A1(n45234), .A2(n45233), .A3(n45238), .A4(n45232), .ZN(
        n45235) );
  AND2_X1 U47335 ( .A1(n45237), .A2(n45238), .ZN(n45239) );
  AOI21_X1 U47336 ( .B1(n45239), .B2(n46359), .A(n46356), .ZN(n45241) );
  OAI21_X1 U47337 ( .B1(n45688), .B2(n45241), .A(n45240), .ZN(n45244) );
  NOR2_X1 U47338 ( .A1(n45697), .A2(n46359), .ZN(n46273) );
  NAND4_X1 U47339 ( .A1(n46273), .A2(n46354), .A3(n46353), .A4(n46267), .ZN(
        n45242) );
  NOR2_X1 U47340 ( .A1(n45244), .A2(n45243), .ZN(n45248) );
  INV_X1 U47341 ( .A(n45245), .ZN(n45246) );
  NAND3_X1 U47342 ( .A1(n45246), .A2(n46350), .A3(n46356), .ZN(n45247) );
  XNOR2_X1 U47343 ( .A(n51408), .B(n45250), .ZN(n45251) );
  XNOR2_X1 U47344 ( .A(n45252), .B(n45251), .ZN(n45261) );
  XNOR2_X1 U47345 ( .A(n45254), .B(n45253), .ZN(n45255) );
  XNOR2_X1 U47346 ( .A(n45256), .B(n45255), .ZN(n45257) );
  XNOR2_X1 U47347 ( .A(n45258), .B(n45257), .ZN(n45259) );
  XNOR2_X1 U47348 ( .A(n45259), .B(n45390), .ZN(n45260) );
  XNOR2_X1 U47349 ( .A(n45261), .B(n45260), .ZN(n45267) );
  XNOR2_X1 U47350 ( .A(n45263), .B(n45262), .ZN(n45264) );
  XNOR2_X1 U47351 ( .A(n45265), .B(n45264), .ZN(n45266) );
  XNOR2_X1 U47352 ( .A(n45266), .B(n45267), .ZN(n45268) );
  XNOR2_X1 U47353 ( .A(n45268), .B(n51525), .ZN(n45370) );
  XNOR2_X1 U47354 ( .A(n45271), .B(n45270), .ZN(n45272) );
  XNOR2_X1 U47355 ( .A(n46113), .B(n45272), .ZN(n45273) );
  XNOR2_X1 U47356 ( .A(n45274), .B(n45273), .ZN(n45275) );
  XNOR2_X1 U47357 ( .A(n45275), .B(n45276), .ZN(n45278) );
  XNOR2_X1 U47358 ( .A(n45278), .B(n45277), .ZN(n45283) );
  XNOR2_X1 U47359 ( .A(n45281), .B(n45280), .ZN(n45282) );
  XNOR2_X1 U47360 ( .A(n45284), .B(n45285), .ZN(n45286) );
  XNOR2_X1 U47361 ( .A(n45287), .B(n45286), .ZN(n45296) );
  XNOR2_X1 U47362 ( .A(n45288), .B(n4931), .ZN(n45290) );
  XNOR2_X1 U47363 ( .A(n45290), .B(n45289), .ZN(n45291) );
  XNOR2_X1 U47364 ( .A(n51465), .B(n45291), .ZN(n45294) );
  XNOR2_X1 U47365 ( .A(n45293), .B(n45294), .ZN(n45295) );
  XNOR2_X1 U47366 ( .A(n45296), .B(n45295), .ZN(n45297) );
  XNOR2_X1 U47367 ( .A(n45437), .B(n45297), .ZN(n45302) );
  XNOR2_X1 U47368 ( .A(n45300), .B(n45299), .ZN(n45301) );
  INV_X1 U47369 ( .A(n45628), .ZN(n45631) );
  XNOR2_X1 U47370 ( .A(n45305), .B(n45306), .ZN(n45316) );
  INV_X1 U47371 ( .A(n45307), .ZN(n45309) );
  XOR2_X1 U47372 ( .A(n4739), .B(n4565), .Z(n45308) );
  XNOR2_X1 U47373 ( .A(n45309), .B(n45308), .ZN(n45312) );
  INV_X1 U47374 ( .A(n45310), .ZN(n45311) );
  XNOR2_X1 U47375 ( .A(n45312), .B(n45311), .ZN(n45313) );
  XNOR2_X1 U47376 ( .A(n45314), .B(n45313), .ZN(n45315) );
  XNOR2_X1 U47377 ( .A(n45316), .B(n45315), .ZN(n45318) );
  XNOR2_X1 U47378 ( .A(n45318), .B(n45317), .ZN(n45319) );
  XNOR2_X1 U47379 ( .A(n51503), .B(n45320), .ZN(n45322) );
  INV_X1 U47380 ( .A(n48535), .ZN(n45324) );
  NAND2_X1 U47382 ( .A1(n48227), .A2(n48239), .ZN(n48238) );
  OR2_X1 U47383 ( .A1(n48524), .A2(n46464), .ZN(n45636) );
  OAI22_X1 U47384 ( .A1(n48548), .A2(n45324), .B1(n48238), .B2(n45636), .ZN(
        n45346) );
  XNOR2_X1 U47385 ( .A(n45326), .B(n45325), .ZN(n45330) );
  XNOR2_X1 U47386 ( .A(n45327), .B(n45328), .ZN(n45329) );
  XNOR2_X1 U47387 ( .A(n45330), .B(n45329), .ZN(n45477) );
  XNOR2_X1 U47388 ( .A(n45332), .B(n45331), .ZN(n45342) );
  XNOR2_X1 U47389 ( .A(n45333), .B(n49109), .ZN(n45334) );
  XNOR2_X1 U47390 ( .A(n45335), .B(n45334), .ZN(n45337) );
  XNOR2_X1 U47391 ( .A(n45337), .B(n45336), .ZN(n45338) );
  XNOR2_X1 U47392 ( .A(n45339), .B(n45338), .ZN(n45340) );
  XNOR2_X1 U47393 ( .A(n45486), .B(n45340), .ZN(n45341) );
  XNOR2_X1 U47394 ( .A(n45342), .B(n45341), .ZN(n45343) );
  XNOR2_X1 U47395 ( .A(n45477), .B(n45343), .ZN(n45345) );
  NAND2_X1 U47396 ( .A1(n45346), .A2(n52059), .ZN(n45375) );
  INV_X1 U47397 ( .A(n45347), .ZN(n45352) );
  XNOR2_X1 U47398 ( .A(n45348), .B(n4818), .ZN(n45349) );
  XNOR2_X1 U47399 ( .A(n45350), .B(n45349), .ZN(n45351) );
  XNOR2_X1 U47400 ( .A(n45352), .B(n45351), .ZN(n45353) );
  XNOR2_X1 U47401 ( .A(n45354), .B(n45353), .ZN(n45356) );
  XNOR2_X1 U47402 ( .A(n45356), .B(n45355), .ZN(n45360) );
  XNOR2_X1 U47403 ( .A(n45358), .B(n45357), .ZN(n45359) );
  XNOR2_X1 U47404 ( .A(n45360), .B(n45359), .ZN(n45362) );
  XNOR2_X1 U47405 ( .A(n45366), .B(n45365), .ZN(n45367) );
  XNOR2_X1 U47406 ( .A(n45368), .B(n45367), .ZN(n45474) );
  XNOR2_X2 U47407 ( .A(n45369), .B(n45474), .ZN(n48546) );
  NOR2_X1 U47408 ( .A1(n48531), .A2(n48546), .ZN(n48536) );
  INV_X1 U47409 ( .A(n45370), .ZN(n48534) );
  AND2_X1 U47410 ( .A1(n48551), .A2(n48536), .ZN(n45630) );
  INV_X1 U47411 ( .A(n45636), .ZN(n48528) );
  NAND3_X1 U47412 ( .A1(n45630), .A2(n48528), .A3(n48534), .ZN(n45374) );
  NAND2_X1 U47413 ( .A1(n45631), .A2(n48546), .ZN(n46369) );
  OAI211_X1 U47414 ( .C1(n48535), .C2(n52059), .A(n46369), .B(n48526), .ZN(
        n45371) );
  NAND3_X1 U47415 ( .A1(n48535), .A2(n48227), .A3(n48547), .ZN(n48554) );
  INV_X1 U47416 ( .A(n48546), .ZN(n45372) );
  NOR2_X1 U47417 ( .A1(n48531), .A2(n2207), .ZN(n48233) );
  AOI22_X1 U47418 ( .A1(n48540), .A2(n48524), .B1(n48233), .B2(n48237), .ZN(
        n45373) );
  INV_X1 U47419 ( .A(n45376), .ZN(n45377) );
  XNOR2_X1 U47420 ( .A(n45377), .B(n45378), .ZN(n45398) );
  XNOR2_X1 U47421 ( .A(n45380), .B(n45379), .ZN(n45381) );
  XNOR2_X1 U47422 ( .A(n45382), .B(n45381), .ZN(n45384) );
  XNOR2_X1 U47423 ( .A(n45383), .B(n45384), .ZN(n45388) );
  XNOR2_X1 U47424 ( .A(n51408), .B(n45385), .ZN(n45387) );
  XNOR2_X1 U47425 ( .A(n45388), .B(n45387), .ZN(n45392) );
  XNOR2_X1 U47426 ( .A(n45390), .B(n45389), .ZN(n45391) );
  XNOR2_X1 U47427 ( .A(n45392), .B(n45391), .ZN(n45396) );
  XNOR2_X1 U47428 ( .A(n45393), .B(n4121), .ZN(n45395) );
  XNOR2_X1 U47429 ( .A(n51101), .B(n51099), .ZN(n45410) );
  XNOR2_X1 U47430 ( .A(n45402), .B(n45401), .ZN(n45404) );
  XNOR2_X1 U47431 ( .A(n45404), .B(n45403), .ZN(n45405) );
  XNOR2_X1 U47432 ( .A(n45406), .B(n45405), .ZN(n45407) );
  XNOR2_X1 U47433 ( .A(n45408), .B(n45407), .ZN(n45409) );
  XNOR2_X1 U47434 ( .A(n45410), .B(n45409), .ZN(n45411) );
  XNOR2_X1 U47435 ( .A(n45412), .B(n45411), .ZN(n45414) );
  XNOR2_X1 U47436 ( .A(n45414), .B(n45413), .ZN(n45420) );
  XNOR2_X1 U47437 ( .A(n45415), .B(n45416), .ZN(n45417) );
  XNOR2_X1 U47438 ( .A(n45418), .B(n45417), .ZN(n45419) );
  INV_X1 U47439 ( .A(n45422), .ZN(n45423) );
  XNOR2_X1 U47440 ( .A(n45424), .B(n45423), .ZN(n45425) );
  XNOR2_X1 U47441 ( .A(n45426), .B(n45425), .ZN(n45427) );
  XNOR2_X1 U47442 ( .A(n45428), .B(n45427), .ZN(n45431) );
  INV_X1 U47443 ( .A(n45429), .ZN(n45430) );
  XNOR2_X1 U47444 ( .A(n45430), .B(n45431), .ZN(n45436) );
  INV_X1 U47445 ( .A(n45432), .ZN(n45433) );
  XNOR2_X1 U47446 ( .A(n45434), .B(n45433), .ZN(n45435) );
  XNOR2_X1 U47447 ( .A(n45436), .B(n45435), .ZN(n45440) );
  INV_X1 U47448 ( .A(n45437), .ZN(n45438) );
  BUF_X2 U47449 ( .A(n45497), .Z(n48417) );
  INV_X1 U47450 ( .A(n45441), .ZN(n45443) );
  XNOR2_X1 U47451 ( .A(n45443), .B(n45442), .ZN(n45444) );
  XNOR2_X1 U47452 ( .A(n45445), .B(n45444), .ZN(n45446) );
  XNOR2_X1 U47453 ( .A(n45447), .B(n45446), .ZN(n45448) );
  XNOR2_X1 U47454 ( .A(n45448), .B(n45449), .ZN(n45453) );
  XNOR2_X1 U47455 ( .A(n45451), .B(n45450), .ZN(n45452) );
  XNOR2_X1 U47456 ( .A(n45453), .B(n45452), .ZN(n45457) );
  XNOR2_X1 U47457 ( .A(n45455), .B(n45454), .ZN(n45456) );
  NAND2_X1 U47459 ( .A1(n48417), .A2(n51068), .ZN(n45574) );
  INV_X1 U47460 ( .A(n45574), .ZN(n45579) );
  INV_X1 U47461 ( .A(n46336), .ZN(n48180) );
  AND2_X1 U47462 ( .A1(n45579), .A2(n48410), .ZN(n45458) );
  NOR2_X1 U47463 ( .A1(n46518), .A2(n45458), .ZN(n45500) );
  XNOR2_X1 U47464 ( .A(n45460), .B(n50967), .ZN(n45461) );
  XNOR2_X1 U47465 ( .A(n45462), .B(n45461), .ZN(n45471) );
  XNOR2_X1 U47466 ( .A(n45463), .B(n4529), .ZN(n45464) );
  XNOR2_X1 U47467 ( .A(n45465), .B(n45464), .ZN(n45466) );
  XNOR2_X1 U47468 ( .A(n45467), .B(n45466), .ZN(n45469) );
  XNOR2_X1 U47469 ( .A(n45469), .B(n45468), .ZN(n45470) );
  XNOR2_X1 U47470 ( .A(n45471), .B(n45470), .ZN(n45472) );
  XNOR2_X1 U47471 ( .A(n45473), .B(n45472), .ZN(n45475) );
  XNOR2_X1 U47472 ( .A(n45475), .B(n45474), .ZN(n48413) );
  INV_X1 U47473 ( .A(n45478), .ZN(n45482) );
  XNOR2_X1 U47474 ( .A(n45480), .B(n45479), .ZN(n45481) );
  XNOR2_X1 U47475 ( .A(n45482), .B(n45481), .ZN(n45483) );
  XNOR2_X1 U47476 ( .A(n45484), .B(n45483), .ZN(n45485) );
  XNOR2_X1 U47477 ( .A(n45486), .B(n45485), .ZN(n45488) );
  XNOR2_X1 U47478 ( .A(n45488), .B(n45487), .ZN(n45493) );
  INV_X1 U47479 ( .A(n45489), .ZN(n45491) );
  XNOR2_X1 U47480 ( .A(n45490), .B(n45491), .ZN(n45492) );
  XNOR2_X1 U47481 ( .A(n45493), .B(n45492), .ZN(n45494) );
  XNOR2_X2 U47482 ( .A(n45495), .B(n45494), .ZN(n48416) );
  OAI21_X1 U47483 ( .B1(n46336), .B2(n51068), .A(n46337), .ZN(n45496) );
  NAND2_X1 U47484 ( .A1(n1752), .A2(n45496), .ZN(n45498) );
  INV_X1 U47485 ( .A(n48403), .ZN(n45575) );
  INV_X1 U47486 ( .A(n45497), .ZN(n46522) );
  NAND2_X1 U47487 ( .A1(n46522), .A2(n46511), .ZN(n45503) );
  INV_X1 U47488 ( .A(n45503), .ZN(n48414) );
  NAND3_X1 U47489 ( .A1(n45575), .A2(n48165), .A3(n48414), .ZN(n45584) );
  NAND4_X1 U47490 ( .A1(n45500), .A2(n45499), .A3(n45498), .A4(n45584), .ZN(
        n45507) );
  NOR3_X1 U47491 ( .A1(n48416), .A2(n2742), .A3(n46511), .ZN(n45501) );
  NAND3_X1 U47492 ( .A1(n45501), .A2(n48166), .A3(n48165), .ZN(n48182) );
  NOR2_X1 U47493 ( .A1(n48403), .A2(n668), .ZN(n46517) );
  NAND2_X1 U47495 ( .A1(n46517), .A2(n46521), .ZN(n45505) );
  NAND2_X1 U47496 ( .A1(n506), .A2(n48404), .ZN(n45502) );
  NOR2_X1 U47497 ( .A1(n45503), .A2(n45502), .ZN(n46514) );
  INV_X1 U47498 ( .A(n46514), .ZN(n45504) );
  OAI211_X1 U47499 ( .C1(n48182), .C2(n48417), .A(n45505), .B(n45504), .ZN(
        n45506) );
  NAND2_X1 U47501 ( .A1(n2034), .A2(n51328), .ZN(n48830) );
  OAI22_X1 U47503 ( .A1(n48819), .A2(n45510), .B1(n45509), .B2(n45743), .ZN(
        n45515) );
  AND2_X1 U47504 ( .A1(n52434), .A2(n48792), .ZN(n48804) );
  NAND3_X1 U47505 ( .A1(n48829), .A2(n48804), .A3(n45752), .ZN(n45513) );
  NAND2_X1 U47506 ( .A1(n51328), .A2(n48792), .ZN(n48793) );
  OAI21_X1 U47507 ( .B1(n45752), .B2(n48808), .A(n48793), .ZN(n45511) );
  OAI21_X1 U47508 ( .B1(n45513), .B2(n48834), .A(n45512), .ZN(n45514) );
  OAI21_X1 U47509 ( .B1(n48817), .B2(n48796), .A(n48833), .ZN(n45517) );
  NOR2_X1 U47510 ( .A1(n52091), .A2(n2034), .ZN(n48824) );
  INV_X1 U47511 ( .A(n4451), .ZN(n45519) );
  NAND2_X1 U47512 ( .A1(n45520), .A2(n45521), .ZN(n45526) );
  NOR2_X1 U47513 ( .A1(n45830), .A2(n45819), .ZN(n45527) );
  MUX2_X1 U47514 ( .A(n45527), .B(n45836), .S(n45834), .Z(n45528) );
  NOR2_X1 U47515 ( .A1(n45529), .A2(n45528), .ZN(n45537) );
  OR2_X1 U47516 ( .A1(n45531), .A2(n45530), .ZN(n45826) );
  NOR2_X1 U47517 ( .A1(n45533), .A2(n45532), .ZN(n45535) );
  OAI21_X1 U47518 ( .B1(n45826), .B2(n45535), .A(n45534), .ZN(n45536) );
  AOI22_X1 U47519 ( .A1(n45545), .A2(n45540), .B1(n45539), .B2(n45538), .ZN(
        n45556) );
  NOR2_X1 U47520 ( .A1(n45541), .A2(n48200), .ZN(n45543) );
  INV_X1 U47521 ( .A(n45545), .ZN(n45548) );
  NAND2_X1 U47522 ( .A1(n48206), .A2(n52050), .ZN(n45546) );
  OAI211_X1 U47523 ( .C1(n45548), .C2(n48200), .A(n45547), .B(n45546), .ZN(
        n45550) );
  NAND2_X1 U47524 ( .A1(n52161), .A2(n52070), .ZN(n48219) );
  OR2_X1 U47525 ( .A1(n3911), .A2(n8061), .ZN(n46539) );
  NAND2_X1 U47526 ( .A1(n45557), .A2(n48510), .ZN(n45573) );
  NAND2_X1 U47527 ( .A1(n48498), .A2(n46474), .ZN(n48192) );
  AND3_X1 U47528 ( .A1(n48192), .A2(n45558), .A3(n46318), .ZN(n45565) );
  NAND2_X1 U47529 ( .A1(n52203), .A2(n46474), .ZN(n48518) );
  OR2_X1 U47530 ( .A1(n48518), .A2(n46322), .ZN(n45561) );
  AOI21_X1 U47531 ( .B1(n45561), .B2(n46471), .A(n48522), .ZN(n45564) );
  NAND3_X1 U47532 ( .A1(n7110), .A2(n51451), .A3(n48517), .ZN(n48519) );
  NOR2_X1 U47533 ( .A1(n48505), .A2(n46471), .ZN(n45566) );
  AND2_X1 U47534 ( .A1(n45566), .A2(n46318), .ZN(n48188) );
  AOI21_X1 U47535 ( .B1(n51451), .B2(n46322), .A(n46474), .ZN(n45567) );
  NAND2_X1 U47536 ( .A1(n48188), .A2(n45567), .ZN(n46317) );
  NOR2_X1 U47537 ( .A1(n46318), .A2(n48505), .ZN(n48500) );
  NAND2_X1 U47538 ( .A1(n48500), .A2(n48512), .ZN(n45568) );
  NOR2_X1 U47539 ( .A1(n46318), .A2(n46478), .ZN(n45570) );
  OAI21_X1 U47540 ( .B1(n48498), .B2(n46471), .A(n48505), .ZN(n45569) );
  OAI211_X1 U47541 ( .C1(n45570), .C2(n45569), .A(n48517), .B(n52203), .ZN(
        n45571) );
  OAI21_X1 U47542 ( .B1(n48417), .B2(n48404), .A(n48179), .ZN(n45576) );
  OAI22_X1 U47543 ( .A1(n46336), .A2(n48417), .B1(n668), .B2(n51068), .ZN(
        n45577) );
  AND2_X1 U47544 ( .A1(n506), .A2(n48416), .ZN(n48174) );
  NAND2_X1 U47545 ( .A1(n45577), .A2(n48174), .ZN(n45583) );
  NAND2_X1 U47546 ( .A1(n48410), .A2(n45578), .ZN(n45580) );
  NAND2_X1 U47547 ( .A1(n45580), .A2(n45579), .ZN(n45582) );
  NAND4_X1 U47548 ( .A1(n45584), .A2(n45583), .A3(n45582), .A4(n45581), .ZN(
        n45585) );
  AND2_X1 U47549 ( .A1(n48112), .A2(n46542), .ZN(n48125) );
  NAND4_X1 U47550 ( .A1(n45587), .A2(n45588), .A3(n48263), .A4(n48436), .ZN(
        n45593) );
  NAND3_X1 U47551 ( .A1(n45589), .A2(n48259), .A3(n48273), .ZN(n45591) );
  AOI21_X1 U47552 ( .B1(n48267), .B2(n45591), .A(n45590), .ZN(n45592) );
  OR2_X1 U47553 ( .A1(n48261), .A2(n48437), .ZN(n45596) );
  NAND2_X1 U47555 ( .A1(n48125), .A2(n8689), .ZN(n48093) );
  AND2_X1 U47556 ( .A1(n48248), .A2(n45597), .ZN(n48480) );
  AOI22_X1 U47557 ( .A1(n45598), .A2(n48493), .B1(n48480), .B2(n48246), .ZN(
        n45599) );
  OR2_X1 U47558 ( .A1(n45599), .A2(n48247), .ZN(n45608) );
  NAND2_X1 U47559 ( .A1(n45602), .A2(n45601), .ZN(n45603) );
  NAND2_X1 U47560 ( .A1(n45603), .A2(n48491), .ZN(n45607) );
  OAI21_X1 U47561 ( .B1(n45604), .B2(n48482), .A(n48488), .ZN(n45605) );
  OAI21_X1 U47562 ( .B1(n48125), .B2(n48110), .A(n48156), .ZN(n45610) );
  AND2_X1 U47563 ( .A1(n48159), .A2(n48140), .ZN(n46535) );
  NAND3_X1 U47564 ( .A1(n8061), .A2(n48100), .A3(n48155), .ZN(n45609) );
  INV_X1 U47565 ( .A(n48159), .ZN(n48117) );
  AND2_X1 U47566 ( .A1(n48117), .A2(n48140), .ZN(n48154) );
  OR2_X1 U47567 ( .A1(n48155), .A2(n48156), .ZN(n48128) );
  INV_X1 U47568 ( .A(n4869), .ZN(n45612) );
  NAND2_X1 U47569 ( .A1(n48455), .A2(n45614), .ZN(n45613) );
  AND2_X1 U47570 ( .A1(n45613), .A2(n46435), .ZN(n45619) );
  XNOR2_X1 U47571 ( .A(n45614), .B(n51732), .ZN(n45615) );
  NAND2_X1 U47572 ( .A1(n46415), .A2(n45615), .ZN(n45620) );
  NAND2_X1 U47573 ( .A1(n48450), .A2(n46444), .ZN(n45616) );
  NAND2_X1 U47574 ( .A1(n45616), .A2(n7275), .ZN(n45617) );
  OAI211_X1 U47575 ( .C1(n45619), .C2(n45618), .A(n45620), .B(n45617), .ZN(
        n45627) );
  INV_X1 U47576 ( .A(n45620), .ZN(n45622) );
  NAND3_X1 U47577 ( .A1(n45622), .A2(n7275), .A3(n45621), .ZN(n45626) );
  OR2_X1 U47578 ( .A1(n46435), .A2(n48456), .ZN(n46433) );
  NAND2_X1 U47579 ( .A1(n48448), .A2(n46412), .ZN(n45623) );
  NAND2_X1 U47580 ( .A1(n46433), .A2(n45623), .ZN(n45624) );
  NAND2_X1 U47581 ( .A1(n45624), .A2(n7275), .ZN(n45625) );
  INV_X1 U47582 ( .A(n46464), .ZN(n48552) );
  OAI21_X1 U47583 ( .B1(n48552), .B2(n48227), .A(n48539), .ZN(n45629) );
  NAND2_X1 U47584 ( .A1(n48531), .A2(n2207), .ZN(n46374) );
  AND2_X1 U47585 ( .A1(n48546), .A2(n2207), .ZN(n48527) );
  NAND3_X1 U47586 ( .A1(n45635), .A2(n48551), .A3(n48237), .ZN(n45633) );
  NOR2_X1 U47587 ( .A1(n45631), .A2(n46464), .ZN(n48234) );
  NAND2_X1 U47588 ( .A1(n48234), .A2(n48526), .ZN(n45632) );
  AND2_X1 U47589 ( .A1(n45633), .A2(n45632), .ZN(n45638) );
  OR2_X1 U47590 ( .A1(n48548), .A2(n48539), .ZN(n48543) );
  NAND3_X1 U47591 ( .A1(n48535), .A2(n48540), .A3(n48551), .ZN(n45634) );
  OR2_X1 U47592 ( .A1(n48549), .A2(n45636), .ZN(n45637) );
  NAND2_X1 U47594 ( .A1(n49167), .A2(n45648), .ZN(n45640) );
  NAND2_X1 U47595 ( .A1(n664), .A2(n540), .ZN(n49169) );
  OAI21_X1 U47596 ( .B1(n49169), .B2(n49177), .A(n49170), .ZN(n45646) );
  INV_X1 U47597 ( .A(n46243), .ZN(n45642) );
  NAND3_X1 U47598 ( .A1(n45642), .A2(n46255), .A3(n540), .ZN(n45644) );
  NAND3_X1 U47599 ( .A1(n49177), .A2(n46252), .A3(n44784), .ZN(n45643) );
  NAND4_X1 U47601 ( .A1(n45650), .A2(n46252), .A3(n46249), .A4(n45649), .ZN(
        n45652) );
  NAND3_X1 U47602 ( .A1(n46239), .A2(n46249), .A3(n49168), .ZN(n45651) );
  OR2_X1 U47603 ( .A1(n45653), .A2(n49162), .ZN(n45655) );
  NAND4_X1 U47604 ( .A1(n49159), .A2(n49162), .A3(n49161), .A4(n49177), .ZN(
        n45654) );
  OAI211_X1 U47605 ( .C1(n45656), .C2(n49162), .A(n45655), .B(n45654), .ZN(
        n45657) );
  INV_X1 U47606 ( .A(n46505), .ZN(n46189) );
  OAI22_X1 U47607 ( .A1(n46396), .A2(n993), .B1(n46501), .B2(n45659), .ZN(
        n45658) );
  NAND2_X1 U47608 ( .A1(n45659), .A2(n46491), .ZN(n46484) );
  NAND2_X1 U47609 ( .A1(n46488), .A2(n46493), .ZN(n46397) );
  NAND2_X1 U47610 ( .A1(n46395), .A2(n46487), .ZN(n46497) );
  OR2_X1 U47611 ( .A1(n46397), .A2(n46497), .ZN(n46190) );
  NOR2_X1 U47612 ( .A1(n46395), .A2(n45661), .ZN(n45662) );
  OR2_X1 U47613 ( .A1(n46488), .A2(n45662), .ZN(n45663) );
  OAI211_X1 U47614 ( .C1(n46490), .C2(n46386), .A(n46502), .B(n45663), .ZN(
        n45664) );
  INV_X1 U47615 ( .A(n49267), .ZN(n45681) );
  INV_X1 U47616 ( .A(n51335), .ZN(n45930) );
  INV_X1 U47617 ( .A(n49265), .ZN(n45669) );
  AOI22_X1 U47618 ( .A1(n45669), .A2(n45668), .B1(n51335), .B2(n49273), .ZN(
        n45673) );
  NAND3_X1 U47619 ( .A1(n45671), .A2(n49277), .A3(n45670), .ZN(n45672) );
  AND2_X1 U47620 ( .A1(n45673), .A2(n45672), .ZN(n45685) );
  AND2_X1 U47621 ( .A1(n52079), .A2(n52086), .ZN(n45678) );
  OAI21_X1 U47622 ( .B1(n52079), .B2(n52086), .A(n46203), .ZN(n45674) );
  INV_X1 U47623 ( .A(n45674), .ZN(n45677) );
  NAND2_X1 U47624 ( .A1(n45675), .A2(n49272), .ZN(n45676) );
  OAI211_X1 U47625 ( .C1(n45678), .C2(n46199), .A(n45677), .B(n45676), .ZN(
        n45684) );
  OAI21_X1 U47626 ( .B1(n45680), .B2(n49261), .A(n45679), .ZN(n45682) );
  NAND2_X1 U47627 ( .A1(n45682), .A2(n45681), .ZN(n45683) );
  INV_X1 U47628 ( .A(n45686), .ZN(n45687) );
  NOR2_X1 U47629 ( .A1(n45688), .A2(n46342), .ZN(n45690) );
  NAND2_X1 U47630 ( .A1(n45697), .A2(n46359), .ZN(n46266) );
  NAND2_X1 U47631 ( .A1(n46274), .A2(n45693), .ZN(n45694) );
  NOR2_X1 U47632 ( .A1(n46274), .A2(n45697), .ZN(n45698) );
  AND2_X1 U47634 ( .A1(n48912), .A2(n48888), .ZN(n48879) );
  NAND2_X1 U47635 ( .A1(n48879), .A2(n51689), .ZN(n48877) );
  NOR2_X1 U47636 ( .A1(n48919), .A2(n51688), .ZN(n48882) );
  INV_X1 U47637 ( .A(n48887), .ZN(n45703) );
  NOR2_X1 U47638 ( .A1(n48905), .A2(n48912), .ZN(n48910) );
  AND2_X1 U47639 ( .A1(n48908), .A2(n48919), .ZN(n48852) );
  OAI211_X1 U47641 ( .C1(n48918), .C2(n5081), .A(n45700), .B(n48886), .ZN(
        n45701) );
  AOI22_X1 U47642 ( .A1(n45703), .A2(n48910), .B1(n48852), .B2(n45701), .ZN(
        n45706) );
  NOR2_X1 U47643 ( .A1(n48853), .A2(n48905), .ZN(n45702) );
  NAND2_X1 U47645 ( .A1(n48847), .A2(n48875), .ZN(n48893) );
  INV_X1 U47646 ( .A(n4824), .ZN(n45708) );
  NAND2_X1 U47647 ( .A1(n52434), .A2(n2034), .ZN(n45746) );
  NOR2_X1 U47648 ( .A1(n48834), .A2(n52434), .ZN(n48798) );
  NAND2_X1 U47649 ( .A1(n45711), .A2(n48808), .ZN(n48836) );
  NOR2_X1 U47650 ( .A1(n45752), .A2(n48836), .ZN(n45712) );
  AND2_X1 U47651 ( .A1(n45711), .A2(n45739), .ZN(n48816) );
  NAND2_X1 U47652 ( .A1(n52090), .A2(n45739), .ZN(n45713) );
  NAND2_X1 U47653 ( .A1(n48816), .A2(n48792), .ZN(n45714) );
  AOI21_X1 U47654 ( .B1(n48817), .B2(n45743), .A(n45714), .ZN(n45715) );
  NOR2_X1 U47655 ( .A1(n45747), .A2(n45715), .ZN(n45716) );
  INV_X1 U47656 ( .A(n4536), .ZN(n45717) );
  XNOR2_X1 U47657 ( .A(n45718), .B(n45717), .ZN(Plaintext[72]) );
  NAND3_X1 U47658 ( .A1(n49564), .A2(n6985), .A3(n51088), .ZN(n45720) );
  AND2_X1 U47659 ( .A1(n49608), .A2(n49599), .ZN(n49586) );
  NAND2_X1 U47660 ( .A1(n49586), .A2(n49579), .ZN(n45723) );
  NOR2_X1 U47661 ( .A1(n49579), .A2(n49599), .ZN(n49609) );
  NAND3_X1 U47662 ( .A1(n49609), .A2(n51088), .A3(n49608), .ZN(n45722) );
  OAI211_X1 U47663 ( .C1(n49592), .C2(n49574), .A(n45723), .B(n45722), .ZN(
        n45724) );
  INV_X1 U47664 ( .A(n49599), .ZN(n49583) );
  NAND2_X1 U47665 ( .A1(n49583), .A2(n49579), .ZN(n49604) );
  INV_X1 U47666 ( .A(n49604), .ZN(n45725) );
  AND2_X1 U47667 ( .A1(n49580), .A2(n49598), .ZN(n49584) );
  NAND3_X1 U47668 ( .A1(n45725), .A2(n49562), .A3(n49584), .ZN(n45733) );
  INV_X1 U47669 ( .A(n49585), .ZN(n45727) );
  AND2_X1 U47670 ( .A1(n49569), .A2(n49579), .ZN(n49551) );
  NAND3_X1 U47671 ( .A1(n45727), .A2(n49551), .A3(n45726), .ZN(n45731) );
  AND2_X1 U47672 ( .A1(n49579), .A2(n49599), .ZN(n49593) );
  NAND3_X1 U47673 ( .A1(n49593), .A2(n49580), .A3(n49569), .ZN(n45730) );
  NAND2_X1 U47674 ( .A1(n49586), .A2(n49598), .ZN(n45729) );
  AND2_X1 U47675 ( .A1(n49608), .A2(n49569), .ZN(n49595) );
  AND4_X1 U47676 ( .A1(n45731), .A2(n45730), .A3(n45729), .A4(n45728), .ZN(
        n45732) );
  INV_X1 U47677 ( .A(n45736), .ZN(n45737) );
  OR2_X1 U47678 ( .A1(n48821), .A2(n45752), .ZN(n45742) );
  OR2_X1 U47679 ( .A1(n48828), .A2(n48808), .ZN(n45740) );
  NOR2_X1 U47680 ( .A1(n52434), .A2(n48792), .ZN(n45745) );
  NOR2_X1 U47681 ( .A1(n2034), .A2(n2033), .ZN(n45750) );
  NAND2_X1 U47682 ( .A1(n2034), .A2(n2033), .ZN(n45748) );
  OAI211_X1 U47683 ( .C1(n45750), .C2(n52091), .A(n52434), .B(n45748), .ZN(
        n45751) );
  NAND2_X1 U47684 ( .A1(n48834), .A2(n45752), .ZN(n45753) );
  INV_X1 U47685 ( .A(n4923), .ZN(n45755) );
  OAI22_X1 U47687 ( .A1(n45758), .A2(n46631), .B1(n45757), .B2(n46623), .ZN(
        n45759) );
  AND2_X1 U47688 ( .A1(n47909), .A2(n46637), .ZN(n46622) );
  OAI21_X1 U47689 ( .B1(n45762), .B2(n46635), .A(n45761), .ZN(n45768) );
  NAND2_X1 U47690 ( .A1(n47907), .A2(n52153), .ZN(n45764) );
  OAI21_X1 U47691 ( .B1(n46630), .B2(n6741), .A(n46637), .ZN(n45765) );
  NAND2_X1 U47692 ( .A1(n45766), .A2(n46627), .ZN(n45767) );
  INV_X1 U47693 ( .A(n47689), .ZN(n45857) );
  NOR2_X1 U47695 ( .A1(n47123), .A2(n46676), .ZN(n45774) );
  OAI21_X1 U47696 ( .B1(n45775), .B2(n45774), .A(n47129), .ZN(n45784) );
  INV_X1 U47697 ( .A(n47123), .ZN(n46847) );
  AND2_X1 U47698 ( .A1(n52053), .A2(n47127), .ZN(n45776) );
  AOI22_X1 U47699 ( .A1(n46847), .A2(n46854), .B1(n46860), .B2(n45776), .ZN(
        n45779) );
  AND2_X1 U47700 ( .A1(n51425), .A2(n3892), .ZN(n47124) );
  NAND2_X1 U47701 ( .A1(n47124), .A2(n47121), .ZN(n45778) );
  INV_X1 U47702 ( .A(n46845), .ZN(n46660) );
  NAND3_X1 U47703 ( .A1(n46660), .A2(n46840), .A3(n46859), .ZN(n45777) );
  AND2_X1 U47704 ( .A1(n46844), .A2(n47126), .ZN(n47119) );
  OAI211_X1 U47705 ( .C1(n51425), .C2(n47128), .A(n47119), .B(n46859), .ZN(
        n45780) );
  NOR2_X1 U47706 ( .A1(n45782), .A2(n45781), .ZN(n45783) );
  AND2_X2 U47707 ( .A1(n45784), .A2(n45783), .ZN(n47655) );
  OR2_X1 U47708 ( .A1(n46707), .A2(n46591), .ZN(n46585) );
  INV_X1 U47709 ( .A(n46585), .ZN(n45787) );
  NAND2_X1 U47710 ( .A1(n46589), .A2(n46708), .ZN(n45785) );
  OAI21_X1 U47711 ( .B1(n46713), .B2(n46701), .A(n45785), .ZN(n45786) );
  AOI21_X1 U47712 ( .B1(n45787), .B2(n46584), .A(n45786), .ZN(n45798) );
  OR2_X1 U47713 ( .A1(n46580), .A2(n46714), .ZN(n46702) );
  OAI21_X1 U47714 ( .B1(n45788), .B2(n46574), .A(n46702), .ZN(n45789) );
  NOR2_X1 U47715 ( .A1(n46583), .A2(n45790), .ZN(n45792) );
  INV_X1 U47716 ( .A(n46701), .ZN(n45791) );
  OAI21_X1 U47717 ( .B1(n44845), .B2(n45792), .A(n45791), .ZN(n45797) );
  NAND2_X1 U47718 ( .A1(n46591), .A2(n405), .ZN(n45794) );
  AOI21_X1 U47719 ( .B1(n46701), .B2(n45794), .A(n51396), .ZN(n45795) );
  NAND2_X1 U47720 ( .A1(n46705), .A2(n45795), .ZN(n45796) );
  AOI21_X1 U47721 ( .B1(n45857), .B2(n47655), .A(n47686), .ZN(n45843) );
  MUX2_X1 U47722 ( .A(n46730), .B(n51488), .S(n46747), .Z(n45805) );
  MUX2_X1 U47723 ( .A(n45806), .B(n45805), .S(n46740), .Z(n45815) );
  NAND2_X1 U47724 ( .A1(n46739), .A2(n46730), .ZN(n45808) );
  NAND3_X1 U47725 ( .A1(n46743), .A2(n46744), .A3(n51344), .ZN(n45807) );
  OAI211_X1 U47726 ( .C1(n46561), .C2(n45809), .A(n45808), .B(n45807), .ZN(
        n45813) );
  MUX2_X1 U47727 ( .A(n46747), .B(n46756), .S(n51344), .Z(n45811) );
  NOR2_X1 U47728 ( .A1(n45811), .A2(n45810), .ZN(n45812) );
  NOR2_X1 U47729 ( .A1(n45813), .A2(n45812), .ZN(n45814) );
  NAND2_X2 U47730 ( .A1(n45814), .A2(n45815), .ZN(n47688) );
  INV_X1 U47731 ( .A(n47688), .ZN(n45886) );
  NAND2_X1 U47732 ( .A1(n45817), .A2(n45816), .ZN(n45824) );
  OAI22_X1 U47733 ( .A1(n44280), .A2(n45819), .B1(n45818), .B2(n45829), .ZN(
        n45822) );
  NAND2_X1 U47734 ( .A1(n45822), .A2(n45821), .ZN(n45823) );
  AND3_X1 U47735 ( .A1(n45825), .A2(n45824), .A3(n45823), .ZN(n45841) );
  INV_X1 U47736 ( .A(n45826), .ZN(n45840) );
  AOI21_X1 U47737 ( .B1(n45829), .B2(n45828), .A(n45827), .ZN(n45831) );
  OR2_X1 U47738 ( .A1(n45831), .A2(n45830), .ZN(n45832) );
  AND2_X1 U47739 ( .A1(n45833), .A2(n45832), .ZN(n45839) );
  NAND2_X1 U47740 ( .A1(n45835), .A2(n45834), .ZN(n45837) );
  NAND2_X1 U47741 ( .A1(n45837), .A2(n45836), .ZN(n45838) );
  NAND2_X1 U47743 ( .A1(n45886), .A2(n47687), .ZN(n47629) );
  INV_X1 U47744 ( .A(n45859), .ZN(n47684) );
  AND2_X1 U47745 ( .A1(n47689), .A2(n47655), .ZN(n45860) );
  INV_X1 U47746 ( .A(n45860), .ZN(n45890) );
  NAND3_X1 U47747 ( .A1(n47684), .A2(n45890), .A3(n47687), .ZN(n45842) );
  NAND2_X1 U47750 ( .A1(n46607), .A2(n46904), .ZN(n45847) );
  NAND2_X1 U47751 ( .A1(n46912), .A2(n46903), .ZN(n45851) );
  INV_X1 U47752 ( .A(n46919), .ZN(n45850) );
  NAND2_X1 U47753 ( .A1(n45852), .A2(n46609), .ZN(n45854) );
  NAND2_X1 U47754 ( .A1(n46919), .A2(n46614), .ZN(n45853) );
  INV_X1 U47755 ( .A(n47651), .ZN(n47675) );
  NAND2_X1 U47756 ( .A1(n45856), .A2(n47675), .ZN(n45865) );
  NOR2_X1 U47757 ( .A1(n47655), .A2(n47689), .ZN(n47685) );
  INV_X1 U47758 ( .A(n47655), .ZN(n47673) );
  INV_X1 U47759 ( .A(n47686), .ZN(n47650) );
  AOI22_X1 U47761 ( .A1(n47685), .A2(n47698), .B1(n47699), .B2(n45857), .ZN(
        n45858) );
  AND2_X1 U47763 ( .A1(n47687), .A2(n47651), .ZN(n47702) );
  NAND2_X1 U47764 ( .A1(n47665), .A2(n47702), .ZN(n47697) );
  NOR2_X1 U47765 ( .A1(n47687), .A2(n47651), .ZN(n47691) );
  NAND3_X1 U47766 ( .A1(n45860), .A2(n47691), .A3(n47688), .ZN(n45862) );
  NAND2_X1 U47767 ( .A1(n47702), .A2(n47688), .ZN(n45861) );
  NAND3_X1 U47768 ( .A1(n47673), .A2(n47687), .A3(n47686), .ZN(n47645) );
  AND4_X1 U47769 ( .A1(n47697), .A2(n45862), .A3(n45861), .A4(n47645), .ZN(
        n45863) );
  NOR3_X1 U47772 ( .A1(n47790), .A2(n51467), .A3(n47786), .ZN(n45868) );
  INV_X1 U47773 ( .A(n51468), .ZN(n45876) );
  NAND2_X1 U47774 ( .A1(n45876), .A2(n47745), .ZN(n47761) );
  NOR2_X1 U47775 ( .A1(n47761), .A2(n47777), .ZN(n45870) );
  NAND2_X1 U47776 ( .A1(n47778), .A2(n47721), .ZN(n47752) );
  NOR2_X1 U47777 ( .A1(n51467), .A2(n47721), .ZN(n45873) );
  NAND4_X1 U47778 ( .A1(n45877), .A2(n47790), .A3(n45873), .A4(n47786), .ZN(
        n45874) );
  OAI211_X1 U47779 ( .C1(n47762), .C2(n47752), .A(n47785), .B(n45874), .ZN(
        n45875) );
  INV_X1 U47780 ( .A(n45875), .ZN(n45881) );
  NAND3_X1 U47782 ( .A1(n644), .A2(n47716), .A3(n51467), .ZN(n45880) );
  INV_X1 U47784 ( .A(n45883), .ZN(n45884) );
  INV_X1 U47786 ( .A(n47702), .ZN(n47664) );
  NAND2_X1 U47787 ( .A1(n47698), .A2(n47655), .ZN(n47668) );
  NOR2_X1 U47788 ( .A1(n45886), .A2(n47655), .ZN(n47683) );
  AND2_X1 U47789 ( .A1(n47689), .A2(n47686), .ZN(n47694) );
  INV_X1 U47792 ( .A(n47642), .ZN(n47667) );
  INV_X1 U47793 ( .A(n47685), .ZN(n45887) );
  AOI22_X1 U47794 ( .A1(n47665), .A2(n47651), .B1(n47702), .B2(n47650), .ZN(
        n45892) );
  INV_X1 U47795 ( .A(n47629), .ZN(n45889) );
  AND2_X1 U47796 ( .A1(n47689), .A2(n47651), .ZN(n47656) );
  INV_X1 U47797 ( .A(n47656), .ZN(n45888) );
  OAI211_X1 U47798 ( .C1(n45892), .C2(n47688), .A(n45891), .B(n47697), .ZN(
        n45893) );
  NOR2_X1 U47799 ( .A1(n45894), .A2(n45893), .ZN(n45895) );
  XNOR2_X1 U47800 ( .A(n45895), .B(n4723), .ZN(Plaintext[14]) );
  INV_X1 U47801 ( .A(n45896), .ZN(n45899) );
  INV_X1 U47802 ( .A(n49191), .ZN(n45901) );
  OR2_X1 U47803 ( .A1(n45907), .A2(n49707), .ZN(n45900) );
  NAND2_X1 U47804 ( .A1(n45901), .A2(n45900), .ZN(n45902) );
  NAND2_X1 U47805 ( .A1(n45902), .A2(n46001), .ZN(n45905) );
  AOI21_X1 U47806 ( .B1(n49726), .B2(n51094), .A(n52052), .ZN(n45904) );
  INV_X1 U47807 ( .A(n45907), .ZN(n45908) );
  NAND2_X1 U47808 ( .A1(n46001), .A2(n49189), .ZN(n45988) );
  MUX2_X1 U47809 ( .A(n45911), .B(n45988), .S(n45999), .Z(n45912) );
  NAND2_X1 U47810 ( .A1(n49235), .A2(n49397), .ZN(n45917) );
  NAND2_X1 U47811 ( .A1(n45914), .A2(n45913), .ZN(n45916) );
  NOR2_X1 U47812 ( .A1(n49686), .A2(n587), .ZN(n49394) );
  NAND2_X1 U47813 ( .A1(n49394), .A2(n49690), .ZN(n45915) );
  OAI211_X1 U47814 ( .C1(n45917), .C2(n49691), .A(n45916), .B(n45915), .ZN(
        n45926) );
  OAI211_X1 U47815 ( .C1(n45919), .C2(n45918), .A(n588), .B(n49686), .ZN(
        n45920) );
  NAND2_X1 U47816 ( .A1(n49242), .A2(n45920), .ZN(n45925) );
  AND2_X1 U47817 ( .A1(n588), .A2(n45921), .ZN(n45923) );
  OAI211_X1 U47818 ( .C1(n49251), .C2(n45923), .A(n656), .B(n49235), .ZN(
        n45924) );
  NAND2_X1 U47819 ( .A1(n45925), .A2(n45924), .ZN(n49400) );
  NOR2_X1 U47820 ( .A1(n49457), .A2(n49465), .ZN(n49462) );
  AND2_X1 U47821 ( .A1(n45929), .A2(n45928), .ZN(n45934) );
  NOR2_X1 U47822 ( .A1(n666), .A2(n49274), .ZN(n45932) );
  XNOR2_X1 U47823 ( .A(n46203), .B(n52086), .ZN(n45931) );
  OAI211_X1 U47824 ( .C1(n49273), .C2(n45932), .A(n45931), .B(n45930), .ZN(
        n45933) );
  NAND3_X1 U47825 ( .A1(n46281), .A2(n45944), .A3(n45937), .ZN(n45938) );
  NAND2_X1 U47826 ( .A1(n45939), .A2(n45938), .ZN(n45940) );
  NAND2_X1 U47828 ( .A1(n45942), .A2(n49142), .ZN(n45948) );
  NAND3_X1 U47829 ( .A1(n45945), .A2(n46299), .A3(n45944), .ZN(n45946) );
  AND3_X1 U47830 ( .A1(n45948), .A2(n45947), .A3(n45946), .ZN(n45955) );
  NAND3_X1 U47831 ( .A1(n49138), .A2(n45949), .A3(n49146), .ZN(n45951) );
  AOI21_X1 U47832 ( .B1(n49148), .B2(n46288), .A(n51515), .ZN(n45950) );
  OR2_X1 U47833 ( .A1(n45951), .A2(n45950), .ZN(n45954) );
  NAND3_X1 U47834 ( .A1(n49151), .A2(n46292), .A3(n49146), .ZN(n45952) );
  AND2_X1 U47835 ( .A1(n46286), .A2(n45952), .ZN(n45953) );
  AND2_X1 U47837 ( .A1(n52107), .A2(n49443), .ZN(n45976) );
  INV_X1 U47838 ( .A(n45976), .ZN(n45977) );
  OR2_X1 U47839 ( .A1(n49654), .A2(n45957), .ZN(n49677) );
  NAND2_X1 U47840 ( .A1(n45961), .A2(n49657), .ZN(n45965) );
  AOI22_X1 U47841 ( .A1(n49669), .A2(n49657), .B1(n45962), .B2(n49656), .ZN(
        n45964) );
  AOI21_X1 U47842 ( .B1(n49671), .B2(n45962), .A(n49667), .ZN(n45963) );
  INV_X1 U47843 ( .A(n46229), .ZN(n49215) );
  NOR2_X1 U47844 ( .A1(n45967), .A2(n49208), .ZN(n46233) );
  NAND4_X1 U47845 ( .A1(n49215), .A2(n45969), .A3(n46233), .A4(n45968), .ZN(
        n45973) );
  INV_X1 U47846 ( .A(n45970), .ZN(n49213) );
  NAND3_X1 U47847 ( .A1(n46223), .A2(n49213), .A3(n46215), .ZN(n45972) );
  OR2_X1 U47848 ( .A1(n52105), .A2(n49201), .ZN(n45971) );
  OAI21_X1 U47849 ( .B1(n49462), .B2(n45977), .A(n47202), .ZN(n49456) );
  NOR2_X1 U47850 ( .A1(n47195), .A2(n51453), .ZN(n47203) );
  OAI21_X1 U47851 ( .B1(n49442), .B2(n51315), .A(n47203), .ZN(n45978) );
  NAND2_X1 U47852 ( .A1(n49456), .A2(n45978), .ZN(n45985) );
  NOR2_X1 U47853 ( .A1(n49450), .A2(n51315), .ZN(n45979) );
  AOI22_X1 U47854 ( .A1(n49434), .A2(n45979), .B1(n47192), .B2(n49418), .ZN(
        n45984) );
  INV_X1 U47855 ( .A(n49434), .ZN(n45980) );
  OR2_X1 U47856 ( .A1(n47195), .A2(n49442), .ZN(n49460) );
  NAND3_X1 U47857 ( .A1(n45980), .A2(n49460), .A3(n2857), .ZN(n45982) );
  NOR2_X1 U47858 ( .A1(n49443), .A2(n51091), .ZN(n49390) );
  NAND2_X1 U47859 ( .A1(n49390), .A2(n49393), .ZN(n45981) );
  AND2_X1 U47860 ( .A1(n49390), .A2(n49407), .ZN(n47199) );
  OAI21_X1 U47861 ( .B1(n47199), .B2(n49423), .A(n47195), .ZN(n45983) );
  INV_X1 U47862 ( .A(n4287), .ZN(n45986) );
  INV_X1 U47863 ( .A(n45989), .ZN(n45991) );
  NOR2_X1 U47864 ( .A1(n49714), .A2(n49721), .ZN(n45990) );
  AOI22_X1 U47865 ( .A1(n49191), .A2(n49725), .B1(n45991), .B2(n45990), .ZN(
        n45992) );
  INV_X1 U47866 ( .A(n45994), .ZN(n46004) );
  INV_X1 U47867 ( .A(n49722), .ZN(n46000) );
  NAND2_X1 U47868 ( .A1(n51295), .A2(n49707), .ZN(n45996) );
  NAND4_X1 U47869 ( .A1(n45997), .A2(n49719), .A3(n49714), .A4(n45996), .ZN(
        n45998) );
  OAI21_X1 U47870 ( .B1(n46000), .B2(n45999), .A(n45998), .ZN(n46002) );
  NAND2_X1 U47871 ( .A1(n46002), .A2(n46001), .ZN(n46003) );
  NAND2_X1 U47872 ( .A1(n49996), .A2(n50315), .ZN(n46005) );
  OR2_X1 U47873 ( .A1(n50001), .A2(n50325), .ZN(n50330) );
  INV_X1 U47874 ( .A(n50330), .ZN(n46006) );
  INV_X1 U47875 ( .A(n50322), .ZN(n46009) );
  OAI21_X1 U47876 ( .B1(n46009), .B2(n46008), .A(n52124), .ZN(n46011) );
  NAND2_X1 U47877 ( .A1(n49932), .A2(n49923), .ZN(n49909) );
  INV_X1 U47878 ( .A(n49973), .ZN(n46015) );
  OAI211_X1 U47879 ( .C1(n49987), .C2(n46015), .A(n46014), .B(n46013), .ZN(
        n46024) );
  NAND2_X1 U47880 ( .A1(n49979), .A2(n47349), .ZN(n46016) );
  NAND3_X1 U47881 ( .A1(n47350), .A2(n47360), .A3(n46016), .ZN(n46023) );
  INV_X1 U47882 ( .A(n49989), .ZN(n46018) );
  OR2_X1 U47883 ( .A1(n49988), .A2(n47354), .ZN(n46017) );
  OAI211_X1 U47884 ( .C1(n46018), .C2(n49979), .A(n46017), .B(n49990), .ZN(
        n46022) );
  NAND3_X1 U47885 ( .A1(n51093), .A2(n49978), .A3(n7798), .ZN(n46020) );
  AOI21_X1 U47886 ( .B1(n49984), .B2(n46020), .A(n49979), .ZN(n46021) );
  OAI22_X1 U47887 ( .A1(n46024), .A2(n46023), .B1(n46022), .B2(n46021), .ZN(
        n46026) );
  AND2_X1 U47888 ( .A1(n49626), .A2(n47352), .ZN(n46025) );
  NAND2_X1 U47889 ( .A1(n46026), .A2(n46025), .ZN(n49889) );
  OR2_X1 U47890 ( .A1(n49654), .A2(n52212), .ZN(n46032) );
  INV_X1 U47891 ( .A(n50027), .ZN(n49661) );
  OAI211_X1 U47892 ( .C1(n49673), .C2(n49667), .A(n49661), .B(n46030), .ZN(
        n46031) );
  AND2_X1 U47893 ( .A1(n51691), .A2(n50287), .ZN(n50308) );
  AND2_X1 U47894 ( .A1(n50309), .A2(n50308), .ZN(n49643) );
  OAI21_X1 U47895 ( .B1(n49643), .B2(n46033), .A(n50294), .ZN(n46039) );
  NAND2_X1 U47896 ( .A1(n50294), .A2(n49635), .ZN(n49637) );
  INV_X1 U47897 ( .A(n49637), .ZN(n50288) );
  OAI21_X1 U47898 ( .B1(n46035), .B2(n50296), .A(n28), .ZN(n46036) );
  NAND2_X1 U47899 ( .A1(n46036), .A2(n50292), .ZN(n46038) );
  INV_X1 U47900 ( .A(n50307), .ZN(n49616) );
  OAI211_X1 U47901 ( .C1(n28), .C2(n50294), .A(n49616), .B(n49953), .ZN(n46037) );
  INV_X1 U47902 ( .A(n49899), .ZN(n47423) );
  NOR2_X1 U47903 ( .A1(n49923), .A2(n49889), .ZN(n49934) );
  XNOR2_X1 U47904 ( .A(n46041), .B(n46040), .ZN(n46047) );
  XNOR2_X1 U47905 ( .A(n52171), .B(n51097), .ZN(n46045) );
  XNOR2_X1 U47906 ( .A(n46045), .B(n46044), .ZN(n46046) );
  XNOR2_X1 U47907 ( .A(n46047), .B(n46046), .ZN(n46057) );
  XNOR2_X1 U47908 ( .A(n46049), .B(n46048), .ZN(n46051) );
  XNOR2_X1 U47909 ( .A(n46051), .B(n46050), .ZN(n46053) );
  XNOR2_X1 U47910 ( .A(n46053), .B(n46052), .ZN(n46055) );
  XNOR2_X1 U47911 ( .A(n46055), .B(n46054), .ZN(n46056) );
  XNOR2_X1 U47912 ( .A(n46058), .B(n46059), .ZN(n46061) );
  XNOR2_X1 U47913 ( .A(n46061), .B(n43196), .ZN(n46072) );
  XNOR2_X1 U47914 ( .A(n46062), .B(n4490), .ZN(n46063) );
  XNOR2_X1 U47915 ( .A(n46064), .B(n46063), .ZN(n46066) );
  XNOR2_X1 U47916 ( .A(n46066), .B(n46065), .ZN(n46067) );
  XNOR2_X1 U47917 ( .A(n46068), .B(n46067), .ZN(n46070) );
  XNOR2_X1 U47918 ( .A(n51409), .B(n46070), .ZN(n46071) );
  XNOR2_X1 U47919 ( .A(n46071), .B(n46072), .ZN(n46076) );
  XNOR2_X1 U47920 ( .A(n46074), .B(n46073), .ZN(n46075) );
  XNOR2_X1 U47921 ( .A(n46075), .B(n46076), .ZN(n46078) );
  AND2_X1 U47922 ( .A1(n50386), .A2(n2199), .ZN(n47322) );
  INV_X1 U47923 ( .A(n47322), .ZN(n46161) );
  INV_X1 U47924 ( .A(n46079), .ZN(n46080) );
  XNOR2_X1 U47925 ( .A(n46080), .B(n46081), .ZN(n46083) );
  XNOR2_X1 U47926 ( .A(n46083), .B(n46082), .ZN(n46094) );
  XNOR2_X1 U47927 ( .A(n46084), .B(n4204), .ZN(n46085) );
  XNOR2_X1 U47928 ( .A(n46086), .B(n46085), .ZN(n46087) );
  XNOR2_X1 U47929 ( .A(n51461), .B(n46087), .ZN(n46089) );
  XNOR2_X1 U47930 ( .A(n46090), .B(n46089), .ZN(n46091) );
  XNOR2_X1 U47931 ( .A(n46092), .B(n46091), .ZN(n46093) );
  XNOR2_X1 U47932 ( .A(n46094), .B(n46093), .ZN(n46096) );
  INV_X1 U47933 ( .A(n47013), .ZN(n50377) );
  XNOR2_X1 U47934 ( .A(n46098), .B(n46097), .ZN(n46099) );
  XNOR2_X1 U47935 ( .A(n46100), .B(n46099), .ZN(n46101) );
  XNOR2_X1 U47936 ( .A(n46102), .B(n46101), .ZN(n46106) );
  XNOR2_X1 U47937 ( .A(n46104), .B(n46103), .ZN(n46105) );
  XNOR2_X1 U47938 ( .A(n46106), .B(n46105), .ZN(n46107) );
  XNOR2_X1 U47939 ( .A(n46108), .B(n46109), .ZN(n46110) );
  XNOR2_X1 U47940 ( .A(n46112), .B(n46111), .ZN(n46115) );
  XNOR2_X1 U47941 ( .A(n46115), .B(n46114), .ZN(n46117) );
  XNOR2_X1 U47942 ( .A(n46117), .B(n46116), .ZN(n46119) );
  XNOR2_X1 U47943 ( .A(n46118), .B(n46119), .ZN(n46136) );
  XNOR2_X1 U47944 ( .A(n51100), .B(n46120), .ZN(n46130) );
  XNOR2_X1 U47945 ( .A(n46122), .B(n49937), .ZN(n46123) );
  XNOR2_X1 U47946 ( .A(n46124), .B(n46123), .ZN(n46125) );
  XNOR2_X1 U47947 ( .A(n46126), .B(n46125), .ZN(n46127) );
  XNOR2_X1 U47948 ( .A(n46128), .B(n46127), .ZN(n46129) );
  XNOR2_X1 U47949 ( .A(n46130), .B(n46129), .ZN(n46132) );
  XNOR2_X1 U47950 ( .A(n46132), .B(n46131), .ZN(n46134) );
  XNOR2_X1 U47951 ( .A(n46134), .B(n46133), .ZN(n46135) );
  XNOR2_X1 U47952 ( .A(n46137), .B(n46138), .ZN(n46139) );
  XNOR2_X1 U47953 ( .A(n46140), .B(n46139), .ZN(n46141) );
  XNOR2_X1 U47954 ( .A(n46142), .B(n46141), .ZN(n46156) );
  XNOR2_X1 U47955 ( .A(n46144), .B(n50759), .ZN(n46145) );
  XNOR2_X1 U47956 ( .A(n46146), .B(n46145), .ZN(n46147) );
  XNOR2_X1 U47957 ( .A(n46148), .B(n46147), .ZN(n46149) );
  XNOR2_X1 U47958 ( .A(n46150), .B(n46149), .ZN(n46151) );
  XNOR2_X1 U47959 ( .A(n46152), .B(n46151), .ZN(n46154) );
  XNOR2_X1 U47960 ( .A(n46154), .B(n51368), .ZN(n46155) );
  XNOR2_X1 U47961 ( .A(n46156), .B(n46155), .ZN(n46157) );
  INV_X1 U47963 ( .A(n2198), .ZN(n50033) );
  AND2_X1 U47964 ( .A1(n51058), .A2(n423), .ZN(n46167) );
  NAND2_X1 U47965 ( .A1(n49731), .A2(n51058), .ZN(n49736) );
  OAI211_X1 U47966 ( .C1(n47012), .C2(n46167), .A(n47322), .B(n49736), .ZN(
        n46159) );
  OAI211_X1 U47967 ( .C1(n46161), .C2(n50377), .A(n46160), .B(n46159), .ZN(
        n46162) );
  INV_X1 U47968 ( .A(n46162), .ZN(n46172) );
  INV_X1 U47969 ( .A(n49731), .ZN(n46163) );
  NAND2_X1 U47970 ( .A1(n46163), .A2(n423), .ZN(n49740) );
  INV_X1 U47971 ( .A(n50374), .ZN(n49743) );
  NAND4_X1 U47972 ( .A1(n50389), .A2(n49743), .A3(n50033), .A4(n47309), .ZN(
        n46166) );
  NAND2_X1 U47973 ( .A1(n50387), .A2(n51058), .ZN(n50044) );
  INV_X1 U47974 ( .A(n50375), .ZN(n47018) );
  OR2_X1 U47975 ( .A1(n49731), .A2(n51058), .ZN(n46164) );
  NAND4_X1 U47976 ( .A1(n50044), .A2(n47018), .A3(n50377), .A4(n46164), .ZN(
        n46165) );
  AND2_X1 U47977 ( .A1(n46165), .A2(n46166), .ZN(n46171) );
  NAND2_X1 U47978 ( .A1(n49738), .A2(n423), .ZN(n47326) );
  INV_X1 U47979 ( .A(n46167), .ZN(n47321) );
  AND2_X1 U47980 ( .A1(n49740), .A2(n50386), .ZN(n47310) );
  INV_X1 U47981 ( .A(n49742), .ZN(n46168) );
  OAI211_X1 U47982 ( .C1(n47310), .C2(n49743), .A(n47019), .B(n46168), .ZN(
        n46169) );
  INV_X1 U47983 ( .A(n49928), .ZN(n49917) );
  NOR2_X1 U47984 ( .A1(n7345), .A2(n49899), .ZN(n46176) );
  OR3_X1 U47985 ( .A1(n49923), .A2(n47420), .A3(n49892), .ZN(n47430) );
  OAI211_X1 U47986 ( .C1(n49929), .C2(n47426), .A(n46177), .B(n47430), .ZN(
        n46178) );
  INV_X1 U47987 ( .A(n46178), .ZN(n46182) );
  NAND2_X1 U47988 ( .A1(n49889), .A2(n46173), .ZN(n49878) );
  INV_X1 U47989 ( .A(n49878), .ZN(n49925) );
  NAND2_X1 U47990 ( .A1(n49923), .A2(n49899), .ZN(n49907) );
  NAND3_X1 U47991 ( .A1(n49925), .A2(n49907), .A3(n49916), .ZN(n46181) );
  INV_X1 U47992 ( .A(n49907), .ZN(n49891) );
  NAND4_X1 U47993 ( .A1(n49891), .A2(n46179), .A3(n49933), .A4(n49889), .ZN(
        n46180) );
  INV_X1 U47995 ( .A(n4782), .ZN(n46184) );
  NAND2_X1 U47997 ( .A1(n46186), .A2(n46404), .ZN(n46195) );
  OR2_X1 U47998 ( .A1(n46501), .A2(n46484), .ZN(n46187) );
  OAI211_X1 U47999 ( .C1(n46397), .C2(n46189), .A(n46188), .B(n46187), .ZN(
        n46192) );
  NAND2_X1 U48000 ( .A1(n46398), .A2(n46190), .ZN(n46191) );
  NOR2_X1 U48001 ( .A1(n46192), .A2(n46191), .ZN(n46194) );
  INV_X1 U48002 ( .A(n46503), .ZN(n46193) );
  NOR2_X1 U48003 ( .A1(n46392), .A2(n46386), .ZN(n46486) );
  NOR2_X1 U48004 ( .A1(n49267), .A2(n46196), .ZN(n46198) );
  NAND3_X1 U48005 ( .A1(n49275), .A2(n46201), .A3(n46199), .ZN(n46200) );
  NAND2_X1 U48006 ( .A1(n49265), .A2(n46201), .ZN(n46202) );
  NAND4_X1 U48007 ( .A1(n46204), .A2(n49273), .A3(n46203), .A4(n46202), .ZN(
        n46208) );
  INV_X1 U48008 ( .A(n49273), .ZN(n46206) );
  NAND2_X1 U48009 ( .A1(n49265), .A2(n49263), .ZN(n46205) );
  NAND3_X1 U48010 ( .A1(n46206), .A2(n49278), .A3(n46205), .ZN(n46207) );
  NOR2_X1 U48011 ( .A1(n46231), .A2(n49198), .ZN(n49218) );
  NAND2_X1 U48012 ( .A1(n49213), .A2(n46229), .ZN(n46209) );
  INV_X1 U48014 ( .A(n46210), .ZN(n46211) );
  NAND2_X1 U48016 ( .A1(n46232), .A2(n49199), .ZN(n46213) );
  OAI211_X1 U48017 ( .C1(n49199), .C2(n46214), .A(n46213), .B(n49216), .ZN(
        n46216) );
  NAND2_X1 U48018 ( .A1(n46216), .A2(n46215), .ZN(n46219) );
  INV_X1 U48019 ( .A(n49203), .ZN(n46217) );
  INV_X1 U48020 ( .A(n49197), .ZN(n49200) );
  NAND3_X1 U48021 ( .A1(n46217), .A2(n49200), .A3(n46223), .ZN(n46218) );
  OR2_X1 U48022 ( .A1(n46226), .A2(n52106), .ZN(n46225) );
  NAND2_X1 U48023 ( .A1(n46223), .A2(n46226), .ZN(n46224) );
  MUX2_X1 U48024 ( .A(n46225), .B(n46224), .S(n46232), .Z(n46236) );
  NAND2_X1 U48025 ( .A1(n46227), .A2(n46226), .ZN(n49223) );
  NAND2_X1 U48026 ( .A1(n46229), .A2(n46228), .ZN(n46230) );
  OAI211_X1 U48027 ( .C1(n46232), .C2(n46231), .A(n49223), .B(n46230), .ZN(
        n46234) );
  NAND2_X1 U48028 ( .A1(n46234), .A2(n46233), .ZN(n46235) );
  NAND2_X1 U48029 ( .A1(n46236), .A2(n46235), .ZN(n46237) );
  NAND3_X1 U48030 ( .A1(n46239), .A2(n49178), .A3(n49162), .ZN(n46242) );
  NAND2_X1 U48031 ( .A1(n49158), .A2(n49161), .ZN(n49175) );
  NOR2_X1 U48032 ( .A1(n49162), .A2(n49163), .ZN(n46240) );
  NAND2_X1 U48033 ( .A1(n49175), .A2(n46240), .ZN(n46241) );
  AND2_X1 U48034 ( .A1(n46242), .A2(n46241), .ZN(n46263) );
  AND2_X1 U48035 ( .A1(n46243), .A2(n46249), .ZN(n46247) );
  INV_X1 U48036 ( .A(n46244), .ZN(n46246) );
  AOI22_X1 U48037 ( .A1(n46248), .A2(n46247), .B1(n46246), .B2(n539), .ZN(
        n46262) );
  AOI21_X1 U48038 ( .B1(n49159), .B2(n49170), .A(n46249), .ZN(n46254) );
  INV_X1 U48039 ( .A(n46250), .ZN(n46251) );
  OAI21_X1 U48040 ( .B1(n46252), .B2(n49163), .A(n46251), .ZN(n46253) );
  OAI211_X1 U48041 ( .C1(n46256), .C2(n46255), .A(n46254), .B(n46253), .ZN(
        n46261) );
  NOR2_X1 U48042 ( .A1(n46257), .A2(n49162), .ZN(n46259) );
  OAI21_X1 U48043 ( .B1(n49171), .B2(n46259), .A(n46258), .ZN(n46260) );
  OR2_X1 U48044 ( .A1(n46342), .A2(n46353), .ZN(n46264) );
  NAND3_X1 U48045 ( .A1(n46266), .A2(n46354), .A3(n46356), .ZN(n46272) );
  NAND2_X1 U48046 ( .A1(n46267), .A2(n46353), .ZN(n46268) );
  OAI211_X1 U48047 ( .C1(n46344), .C2(n46356), .A(n46342), .B(n46268), .ZN(
        n46271) );
  NAND2_X1 U48048 ( .A1(n46345), .A2(n46269), .ZN(n46270) );
  OAI21_X1 U48049 ( .B1(n46277), .B2(n46276), .A(n46275), .ZN(n46278) );
  NOR2_X1 U48050 ( .A1(n653), .A2(n49020), .ZN(n49004) );
  NAND2_X1 U48051 ( .A1(n46298), .A2(n46280), .ZN(n46285) );
  NAND2_X1 U48052 ( .A1(n49151), .A2(n46281), .ZN(n46284) );
  NAND3_X1 U48053 ( .A1(n46289), .A2(n46299), .A3(n49146), .ZN(n46294) );
  NAND3_X1 U48054 ( .A1(n46292), .A2(n46291), .A3(n46290), .ZN(n46293) );
  NAND2_X1 U48055 ( .A1(n46294), .A2(n46293), .ZN(n46295) );
  NOR2_X1 U48056 ( .A1(n46296), .A2(n46295), .ZN(n46305) );
  NAND2_X1 U48057 ( .A1(n46297), .A2(n51515), .ZN(n46301) );
  NAND2_X1 U48058 ( .A1(n46299), .A2(n46298), .ZN(n46300) );
  OAI211_X1 U48059 ( .C1(n7657), .C2(n46302), .A(n46301), .B(n46300), .ZN(
        n46303) );
  NAND2_X1 U48060 ( .A1(n46303), .A2(n49142), .ZN(n46304) );
  AOI22_X1 U48061 ( .A1(n49008), .A2(n49004), .B1(n48988), .B2(n48984), .ZN(
        n46308) );
  NAND2_X1 U48062 ( .A1(n46934), .A2(n49020), .ZN(n49042) );
  NAND2_X1 U48063 ( .A1(n49037), .A2(n49019), .ZN(n49024) );
  OAI21_X1 U48064 ( .B1(n52179), .B2(n49021), .A(n49024), .ZN(n46306) );
  NAND3_X1 U48065 ( .A1(n49042), .A2(n51321), .A3(n46306), .ZN(n46307) );
  OAI211_X1 U48066 ( .C1(n48989), .C2(n49019), .A(n46308), .B(n46307), .ZN(
        n46311) );
  NOR2_X1 U48067 ( .A1(n49047), .A2(n49020), .ZN(n49002) );
  OAI21_X1 U48068 ( .B1(n6389), .B2(n51310), .A(n52179), .ZN(n46309) );
  NAND2_X1 U48069 ( .A1(n46309), .A2(n49029), .ZN(n46310) );
  NAND2_X1 U48071 ( .A1(n46312), .A2(n46474), .ZN(n46314) );
  NAND3_X1 U48072 ( .A1(n46314), .A2(n45562), .A3(n46313), .ZN(n46316) );
  AND2_X1 U48074 ( .A1(n46471), .A2(n46318), .ZN(n48499) );
  INV_X1 U48075 ( .A(n48498), .ZN(n48513) );
  NOR2_X1 U48076 ( .A1(n46322), .A2(n48517), .ZN(n46319) );
  OR2_X1 U48077 ( .A1(n48512), .A2(n46319), .ZN(n46320) );
  OAI211_X1 U48078 ( .C1(n48499), .C2(n48513), .A(n48505), .B(n46320), .ZN(
        n46329) );
  OR2_X1 U48079 ( .A1(n52066), .A2(n46471), .ZN(n46321) );
  NOR2_X1 U48080 ( .A1(n48518), .A2(n46321), .ZN(n48523) );
  INV_X1 U48081 ( .A(n48523), .ZN(n46328) );
  NAND2_X1 U48082 ( .A1(n48498), .A2(n45562), .ZN(n46326) );
  NAND2_X1 U48083 ( .A1(n46322), .A2(n46474), .ZN(n46324) );
  NAND2_X1 U48084 ( .A1(n46324), .A2(n52066), .ZN(n46325) );
  NAND3_X1 U48085 ( .A1(n46326), .A2(n48510), .A3(n46325), .ZN(n46327) );
  NAND2_X1 U48087 ( .A1(n48416), .A2(n51068), .ZN(n46332) );
  XNOR2_X1 U48088 ( .A(n48410), .B(n46332), .ZN(n46334) );
  NAND2_X1 U48089 ( .A1(n48416), .A2(n48417), .ZN(n48405) );
  AND2_X1 U48090 ( .A1(n2742), .A2(n48405), .ZN(n46333) );
  NAND2_X1 U48091 ( .A1(n46335), .A2(n48421), .ZN(n46341) );
  NAND2_X1 U48092 ( .A1(n46336), .A2(n46511), .ZN(n48171) );
  NAND2_X1 U48093 ( .A1(n48171), .A2(n46337), .ZN(n46338) );
  NAND2_X1 U48094 ( .A1(n48404), .A2(n48417), .ZN(n48402) );
  NAND3_X1 U48095 ( .A1(n46338), .A2(n48416), .A3(n48402), .ZN(n46340) );
  NAND2_X1 U48096 ( .A1(n46346), .A2(n44765), .ZN(n46347) );
  OAI211_X1 U48097 ( .C1(n46355), .C2(n46354), .A(n46353), .B(n46352), .ZN(
        n46363) );
  AOI21_X1 U48098 ( .B1(n46358), .B2(n46357), .A(n46356), .ZN(n46362) );
  NAND2_X1 U48099 ( .A1(n46360), .A2(n46359), .ZN(n46361) );
  NAND3_X1 U48100 ( .A1(n46363), .A2(n46362), .A3(n46361), .ZN(n46364) );
  INV_X2 U48101 ( .A(n47442), .ZN(n48722) );
  INV_X1 U48102 ( .A(n48550), .ZN(n46367) );
  OAI211_X1 U48103 ( .C1(n48535), .C2(n46367), .A(n52059), .B(n48238), .ZN(
        n46368) );
  AND2_X1 U48104 ( .A1(n48543), .A2(n46368), .ZN(n46379) );
  NOR2_X1 U48105 ( .A1(n48233), .A2(n46369), .ZN(n46372) );
  OR2_X1 U48106 ( .A1(n46464), .A2(n2207), .ZN(n48229) );
  AOI22_X1 U48107 ( .A1(n48552), .A2(n48227), .B1(n48229), .B2(n48531), .ZN(
        n46371) );
  NOR2_X1 U48108 ( .A1(n48550), .A2(n48531), .ZN(n46370) );
  AOI22_X1 U48109 ( .A1(n46372), .A2(n46371), .B1(n46370), .B2(n48526), .ZN(
        n48556) );
  INV_X1 U48110 ( .A(n48526), .ZN(n46373) );
  NAND3_X1 U48111 ( .A1(n46373), .A2(n48552), .A3(n48536), .ZN(n46378) );
  INV_X1 U48112 ( .A(n46374), .ZN(n46376) );
  NOR2_X1 U48114 ( .A1(n48722), .A2(n48769), .ZN(n48766) );
  NAND2_X1 U48115 ( .A1(n48745), .A2(n48766), .ZN(n47441) );
  INV_X1 U48117 ( .A(n48749), .ZN(n46421) );
  NAND2_X1 U48118 ( .A1(n46380), .A2(n46395), .ZN(n46383) );
  AOI21_X1 U48119 ( .B1(n46489), .B2(n46491), .A(n8207), .ZN(n46382) );
  NAND2_X1 U48120 ( .A1(n52136), .A2(n46488), .ZN(n46381) );
  OAI211_X1 U48121 ( .C1(n46488), .C2(n46383), .A(n46382), .B(n46381), .ZN(
        n46384) );
  NAND2_X1 U48122 ( .A1(n46384), .A2(n46505), .ZN(n46390) );
  NAND3_X1 U48123 ( .A1(n46385), .A2(n46492), .A3(n46403), .ZN(n46389) );
  NAND3_X1 U48124 ( .A1(n46387), .A2(n46386), .A3(n46503), .ZN(n46388) );
  AND3_X1 U48125 ( .A1(n46390), .A2(n46389), .A3(n46388), .ZN(n46402) );
  OAI21_X1 U48126 ( .B1(n46394), .B2(n46393), .A(n46494), .ZN(n46401) );
  NAND4_X1 U48127 ( .A1(n46398), .A2(n46493), .A3(n46403), .A4(n46397), .ZN(
        n46399) );
  NAND4_X1 U48128 ( .A1(n46402), .A2(n46401), .A3(n46400), .A4(n46399), .ZN(
        n46410) );
  INV_X1 U48129 ( .A(n46484), .ZN(n46500) );
  INV_X1 U48130 ( .A(n46403), .ZN(n46405) );
  OAI21_X1 U48131 ( .B1(n46405), .B2(n46483), .A(n46404), .ZN(n46406) );
  INV_X1 U48132 ( .A(n46406), .ZN(n46408) );
  MUX2_X1 U48133 ( .A(n46500), .B(n46408), .S(n46407), .Z(n46409) );
  NAND2_X1 U48134 ( .A1(n46441), .A2(n46412), .ZN(n48464) );
  AOI21_X1 U48135 ( .B1(n48451), .B2(n7275), .A(n46444), .ZN(n46413) );
  OR2_X1 U48136 ( .A1(n46413), .A2(n48450), .ZN(n46416) );
  AND2_X1 U48137 ( .A1(n46448), .A2(n48455), .ZN(n46414) );
  AOI22_X1 U48138 ( .A1(n46416), .A2(n46415), .B1(n46414), .B2(n8585), .ZN(
        n46419) );
  OAI21_X1 U48139 ( .B1(n46448), .B2(n48449), .A(n48463), .ZN(n46417) );
  AND3_X2 U48140 ( .A1(n46420), .A2(n46419), .A3(n46418), .ZN(n48734) );
  AOI21_X1 U48142 ( .B1(n47441), .B2(n48786), .A(n46422), .ZN(n46430) );
  NOR3_X1 U48143 ( .A1(n48730), .A2(n48722), .A3(n48751), .ZN(n46425) );
  AND3_X1 U48144 ( .A1(n48722), .A2(n48734), .A3(n48751), .ZN(n46424) );
  NAND3_X1 U48145 ( .A1(n48778), .A2(n52067), .A3(n48722), .ZN(n46423) );
  OAI21_X1 U48146 ( .B1(n46425), .B2(n46424), .A(n46423), .ZN(n46428) );
  NAND2_X1 U48147 ( .A1(n48722), .A2(n48729), .ZN(n46426) );
  OR2_X1 U48148 ( .A1(n46426), .A2(n48730), .ZN(n48720) );
  NAND3_X1 U48149 ( .A1(n48750), .A2(n52067), .A3(n48729), .ZN(n46427) );
  XNOR2_X1 U48150 ( .A(n46431), .B(n4744), .ZN(Plaintext[71]) );
  NAND2_X1 U48151 ( .A1(n48451), .A2(n48449), .ZN(n46432) );
  AOI21_X1 U48152 ( .B1(n46433), .B2(n46432), .A(n46434), .ZN(n46440) );
  AOI21_X1 U48153 ( .B1(n48450), .B2(n46446), .A(n883), .ZN(n46439) );
  INV_X1 U48154 ( .A(n46434), .ZN(n46436) );
  OAI211_X1 U48155 ( .C1(n46440), .C2(n51732), .A(n46439), .B(n46438), .ZN(
        n46454) );
  NAND2_X1 U48156 ( .A1(n48455), .A2(n46441), .ZN(n46442) );
  MUX2_X1 U48157 ( .A(n46443), .B(n46442), .S(n48448), .Z(n46453) );
  NOR2_X1 U48158 ( .A1(n7275), .A2(n46444), .ZN(n46445) );
  OAI211_X1 U48159 ( .C1(n46449), .C2(n46448), .A(n7275), .B(n46447), .ZN(
        n46450) );
  NAND2_X1 U48160 ( .A1(n46450), .A2(n48457), .ZN(n46451) );
  OAI21_X1 U48161 ( .B1(n48485), .B2(n44409), .A(n48474), .ZN(n46455) );
  OAI211_X1 U48162 ( .C1(n48254), .C2(n46456), .A(n48478), .B(n46455), .ZN(
        n46461) );
  XNOR2_X1 U48163 ( .A(n48485), .B(n48487), .ZN(n46459) );
  NAND2_X1 U48164 ( .A1(n604), .A2(n48247), .ZN(n46457) );
  NAND4_X1 U48165 ( .A1(n46459), .A2(n48493), .A3(n46458), .A4(n46457), .ZN(
        n46460) );
  NOR2_X1 U48166 ( .A1(n48659), .A2(n48674), .ZN(n48669) );
  NAND3_X1 U48168 ( .A1(n48236), .A2(n48237), .A3(n48547), .ZN(n46469) );
  NAND3_X1 U48169 ( .A1(n48230), .A2(n48547), .A3(n48526), .ZN(n46467) );
  NAND2_X1 U48170 ( .A1(n48531), .A2(n48552), .ZN(n46465) );
  OAI21_X1 U48171 ( .B1(n48526), .B2(n46465), .A(n48524), .ZN(n46466) );
  NAND2_X1 U48172 ( .A1(n46467), .A2(n46466), .ZN(n46468) );
  NAND2_X1 U48174 ( .A1(n48669), .A2(n48703), .ZN(n47404) );
  NAND2_X1 U48175 ( .A1(n48517), .A2(n46471), .ZN(n46472) );
  NOR2_X1 U48176 ( .A1(n48196), .A2(n46472), .ZN(n46473) );
  AOI22_X1 U48177 ( .A1(n46473), .A2(n48508), .B1(n45562), .B2(n48510), .ZN(
        n46482) );
  NAND3_X1 U48178 ( .A1(n48498), .A2(n48522), .A3(n46474), .ZN(n46477) );
  OAI21_X1 U48179 ( .B1(n48521), .B2(n48505), .A(n48517), .ZN(n46476) );
  NAND2_X1 U48180 ( .A1(n48518), .A2(n48505), .ZN(n46479) );
  NAND2_X1 U48181 ( .A1(n48507), .A2(n46479), .ZN(n46480) );
  NOR2_X1 U48182 ( .A1(n46484), .A2(n46483), .ZN(n46485) );
  OAI21_X1 U48183 ( .B1(n46486), .B2(n46485), .A(n46505), .ZN(n46509) );
  OAI22_X1 U48184 ( .A1(n46490), .A2(n46489), .B1(n46488), .B2(n46487), .ZN(
        n46496) );
  AOI21_X1 U48185 ( .B1(n46492), .B2(n991), .A(n51426), .ZN(n46495) );
  AOI22_X1 U48186 ( .A1(n46496), .A2(n46495), .B1(n46494), .B2(n46493), .ZN(
        n46508) );
  NOR2_X1 U48187 ( .A1(n51426), .A2(n46497), .ZN(n46499) );
  INV_X1 U48188 ( .A(n46501), .ZN(n46504) );
  OAI211_X1 U48189 ( .C1(n46505), .C2(n46504), .A(n46503), .B(n46502), .ZN(
        n46506) );
  NOR2_X1 U48192 ( .A1(n46511), .A2(n668), .ZN(n46512) );
  MUX2_X1 U48193 ( .A(n2742), .B(n46512), .S(n48417), .Z(n46513) );
  OAI21_X1 U48194 ( .B1(n46513), .B2(n48414), .A(n48412), .ZN(n46516) );
  NOR2_X1 U48196 ( .A1(n46518), .A2(n46517), .ZN(n46526) );
  AND2_X1 U48197 ( .A1(n48166), .A2(n51068), .ZN(n46520) );
  NAND2_X1 U48198 ( .A1(n48179), .A2(n46522), .ZN(n46523) );
  MUX2_X1 U48199 ( .A(n46524), .B(n46523), .S(n48410), .Z(n46525) );
  AND2_X1 U48200 ( .A1(n48702), .A2(n48674), .ZN(n48696) );
  INV_X1 U48201 ( .A(n48697), .ZN(n48664) );
  OR2_X1 U48202 ( .A1(n48664), .A2(n48674), .ZN(n47247) );
  OAI211_X1 U48203 ( .C1(n48696), .C2(n48698), .A(n47247), .B(n48687), .ZN(
        n46529) );
  NAND2_X1 U48204 ( .A1(n51658), .A2(n48702), .ZN(n48688) );
  NAND2_X1 U48205 ( .A1(n48697), .A2(n48674), .ZN(n48682) );
  INV_X1 U48206 ( .A(n48659), .ZN(n47410) );
  NAND2_X1 U48207 ( .A1(n51659), .A2(n48674), .ZN(n46532) );
  AND4_X1 U48208 ( .A1(n48702), .A2(n47410), .A3(n46532), .A4(n48664), .ZN(
        n46533) );
  XNOR2_X1 U48209 ( .A(n46534), .B(n4737), .ZN(Plaintext[64]) );
  NOR2_X1 U48210 ( .A1(n48159), .A2(n48112), .ZN(n48135) );
  INV_X1 U48211 ( .A(n48160), .ZN(n46536) );
  NAND2_X1 U48212 ( .A1(n46536), .A2(n46535), .ZN(n46537) );
  OAI211_X1 U48213 ( .C1(n46540), .C2(n46539), .A(n46538), .B(n46537), .ZN(
        n46541) );
  INV_X1 U48214 ( .A(n46541), .ZN(n46551) );
  AND2_X1 U48215 ( .A1(n48159), .A2(n48156), .ZN(n48097) );
  NOR2_X1 U48216 ( .A1(n48140), .A2(n48100), .ZN(n48130) );
  NAND3_X1 U48218 ( .A1(n48097), .A2(n48130), .A3(n48136), .ZN(n46544) );
  NAND3_X1 U48219 ( .A1(n48136), .A2(n48112), .A3(n48140), .ZN(n48094) );
  NAND3_X1 U48220 ( .A1(n48112), .A2(n46547), .A3(n48155), .ZN(n46543) );
  AND3_X1 U48221 ( .A1(n48094), .A2(n46544), .A3(n46543), .ZN(n46550) );
  AND3_X1 U48222 ( .A1(n48140), .A2(n48100), .A3(n48155), .ZN(n46546) );
  AOI22_X1 U48225 ( .A1(n46546), .A2(n48095), .B1(n48141), .B2(n48136), .ZN(
        n46549) );
  OAI211_X1 U48226 ( .C1(n48100), .C2(n48136), .A(n48153), .B(n48154), .ZN(
        n46548) );
  INV_X1 U48227 ( .A(n46552), .ZN(n46553) );
  AOI22_X1 U48228 ( .A1(n46744), .A2(n46743), .B1(n51344), .B2(n44850), .ZN(
        n46559) );
  INV_X1 U48229 ( .A(n46739), .ZN(n46557) );
  NAND2_X1 U48230 ( .A1(n46557), .A2(n46738), .ZN(n46558) );
  MUX2_X1 U48231 ( .A(n46559), .B(n46558), .S(n46740), .Z(n46563) );
  NAND2_X1 U48232 ( .A1(n46561), .A2(n46560), .ZN(n46562) );
  NAND2_X1 U48233 ( .A1(n47103), .A2(n47108), .ZN(n47105) );
  OAI21_X1 U48234 ( .B1(n47104), .B2(n47087), .A(n47106), .ZN(n46566) );
  NAND2_X1 U48235 ( .A1(n46570), .A2(n47109), .ZN(n46571) );
  INV_X1 U48237 ( .A(n47608), .ZN(n47616) );
  AND2_X1 U48238 ( .A1(n46572), .A2(n46591), .ZN(n46581) );
  AOI22_X1 U48239 ( .A1(n46581), .A2(n46714), .B1(n51396), .B2(n46587), .ZN(
        n46578) );
  NAND2_X1 U48240 ( .A1(n46586), .A2(n46573), .ZN(n46577) );
  INV_X1 U48241 ( .A(n46574), .ZN(n46592) );
  NAND4_X1 U48242 ( .A1(n46699), .A2(n46592), .A3(n46710), .A4(n46575), .ZN(
        n46576) );
  OAI211_X1 U48243 ( .C1(n46578), .C2(n46586), .A(n46577), .B(n46576), .ZN(
        n46579) );
  INV_X1 U48244 ( .A(n46579), .ZN(n46602) );
  INV_X1 U48245 ( .A(n46581), .ZN(n46582) );
  NAND2_X1 U48246 ( .A1(n46587), .A2(n46595), .ZN(n46588) );
  OAI211_X1 U48247 ( .C1(n46591), .C2(n46589), .A(n46588), .B(n46710), .ZN(
        n46590) );
  INV_X1 U48248 ( .A(n46590), .ZN(n46594) );
  NOR2_X1 U48249 ( .A1(n46708), .A2(n46591), .ZN(n46715) );
  NAND2_X1 U48250 ( .A1(n46592), .A2(n46715), .ZN(n46593) );
  OAI211_X1 U48251 ( .C1(n46596), .C2(n46595), .A(n46594), .B(n46593), .ZN(
        n46601) );
  OAI211_X1 U48252 ( .C1(n46705), .C2(n46703), .A(n46714), .B(n46715), .ZN(
        n46599) );
  NOR2_X1 U48253 ( .A1(n46703), .A2(n51317), .ZN(n46598) );
  OR2_X1 U48254 ( .A1(n46599), .A2(n46598), .ZN(n46600) );
  AOI22_X1 U48255 ( .A1(n46607), .A2(n46603), .B1(n46903), .B2(n46901), .ZN(
        n46605) );
  AND2_X1 U48256 ( .A1(n46918), .A2(n46908), .ZN(n46685) );
  AND3_X1 U48257 ( .A1(n46607), .A2(n51399), .A3(n52169), .ZN(n46608) );
  NOR2_X1 U48258 ( .A1(n46608), .A2(n46915), .ZN(n46620) );
  NAND3_X1 U48259 ( .A1(n46609), .A2(n46689), .A3(n46905), .ZN(n46610) );
  INV_X1 U48260 ( .A(n46611), .ZN(n46619) );
  INV_X1 U48261 ( .A(n46920), .ZN(n46612) );
  NAND2_X1 U48262 ( .A1(n46614), .A2(n46904), .ZN(n46615) );
  NAND4_X1 U48263 ( .A1(n46617), .A2(n51399), .A3(n46616), .A4(n46615), .ZN(
        n46618) );
  NAND3_X1 U48266 ( .A1(n46623), .A2(n52154), .A3(n46622), .ZN(n46624) );
  NAND3_X1 U48267 ( .A1(n46629), .A2(n46628), .A3(n46627), .ZN(n46645) );
  OAI22_X1 U48268 ( .A1(n46633), .A2(n46632), .B1(n46631), .B2(n46630), .ZN(
        n46634) );
  INV_X1 U48269 ( .A(n46634), .ZN(n46644) );
  AOI21_X1 U48270 ( .B1(n44654), .B2(n46637), .A(n46635), .ZN(n46640) );
  NOR2_X1 U48271 ( .A1(n52154), .A2(n46642), .ZN(n46638) );
  OAI21_X1 U48272 ( .B1(n46638), .B2(n46637), .A(n5325), .ZN(n46639) );
  OAI211_X1 U48273 ( .C1(n46642), .C2(n46641), .A(n46640), .B(n46639), .ZN(
        n46643) );
  INV_X1 U48275 ( .A(n47586), .ZN(n47589) );
  AND2_X1 U48276 ( .A1(n47592), .A2(n47589), .ZN(n46669) );
  NAND2_X1 U48277 ( .A1(n47118), .A2(n51425), .ZN(n46651) );
  INV_X1 U48278 ( .A(n46840), .ZN(n46846) );
  NAND2_X1 U48279 ( .A1(n46650), .A2(n46863), .ZN(n47134) );
  NOR2_X1 U48280 ( .A1(n46860), .A2(n46842), .ZN(n46681) );
  INV_X1 U48281 ( .A(n46681), .ZN(n46657) );
  OAI211_X1 U48282 ( .C1(n47128), .C2(n46842), .A(n46654), .B(n47127), .ZN(
        n46652) );
  AND2_X1 U48283 ( .A1(n47121), .A2(n46652), .ZN(n46656) );
  NAND2_X1 U48284 ( .A1(n46840), .A2(n46676), .ZN(n46653) );
  OAI21_X1 U48285 ( .B1(n47123), .B2(n46654), .A(n46653), .ZN(n46655) );
  AOI21_X1 U48286 ( .B1(n46657), .B2(n46656), .A(n46655), .ZN(n46663) );
  INV_X1 U48287 ( .A(n47129), .ZN(n46659) );
  NAND2_X1 U48288 ( .A1(n46854), .A2(n46860), .ZN(n46658) );
  OAI21_X1 U48289 ( .B1(n46659), .B2(n47118), .A(n46658), .ZN(n46661) );
  NAND2_X1 U48290 ( .A1(n46661), .A2(n46660), .ZN(n46662) );
  OR2_X1 U48291 ( .A1(n46668), .A2(n2163), .ZN(n47587) );
  INV_X1 U48292 ( .A(n47587), .ZN(n46664) );
  NAND4_X1 U48294 ( .A1(n46669), .A2(n46664), .A3(n8448), .A4(n47617), .ZN(
        n46667) );
  NAND2_X1 U48295 ( .A1(n46668), .A2(n47599), .ZN(n47468) );
  INV_X1 U48296 ( .A(n47468), .ZN(n46665) );
  NAND2_X1 U48297 ( .A1(n46665), .A2(n47462), .ZN(n46666) );
  OAI211_X1 U48298 ( .C1(n47616), .C2(n47622), .A(n46667), .B(n46666), .ZN(
        n46674) );
  AND2_X1 U48300 ( .A1(n47596), .A2(n2163), .ZN(n47266) );
  NAND2_X1 U48301 ( .A1(n46669), .A2(n47266), .ZN(n46672) );
  OR2_X1 U48302 ( .A1(n51401), .A2(n46668), .ZN(n47614) );
  NAND2_X1 U48303 ( .A1(n47589), .A2(n47618), .ZN(n46670) );
  NAND3_X1 U48304 ( .A1(n1187), .A2(n47614), .A3(n46670), .ZN(n46671) );
  NAND3_X1 U48305 ( .A1(n47615), .A2(n46672), .A3(n46671), .ZN(n46673) );
  NOR2_X1 U48306 ( .A1(n46674), .A2(n46673), .ZN(n46675) );
  XNOR2_X1 U48307 ( .A(n46675), .B(n4835), .ZN(Plaintext[10]) );
  NAND2_X1 U48308 ( .A1(n46863), .A2(n3892), .ZN(n46678) );
  OAI211_X1 U48309 ( .C1(n46852), .C2(n46678), .A(n2469), .B(n46677), .ZN(
        n46684) );
  INV_X1 U48310 ( .A(n46863), .ZN(n46679) );
  OAI211_X1 U48311 ( .C1(n47124), .C2(n46845), .A(n46679), .B(n52053), .ZN(
        n46682) );
  OAI21_X1 U48312 ( .B1(n46903), .B2(n51359), .A(n46685), .ZN(n46688) );
  OAI21_X1 U48313 ( .B1(n46905), .B2(n51399), .A(n46921), .ZN(n46687) );
  MUX2_X1 U48314 ( .A(n46688), .B(n46687), .S(n46913), .Z(n46698) );
  NOR2_X1 U48315 ( .A1(n46902), .A2(n46901), .ZN(n46916) );
  INV_X1 U48316 ( .A(n46689), .ZN(n46690) );
  OAI211_X1 U48317 ( .C1(n46916), .C2(n51399), .A(n46905), .B(n46690), .ZN(
        n46697) );
  NAND3_X1 U48318 ( .A1(n46919), .A2(n46693), .A3(n46904), .ZN(n46696) );
  NAND3_X1 U48319 ( .A1(n46694), .A2(n46693), .A3(n46692), .ZN(n46695) );
  NAND2_X1 U48321 ( .A1(n46702), .A2(n46701), .ZN(n46704) );
  AOI22_X1 U48322 ( .A1(n46706), .A2(n46705), .B1(n46704), .B2(n46703), .ZN(
        n46718) );
  OAI21_X1 U48323 ( .B1(n46710), .B2(n46709), .A(n46707), .ZN(n46712) );
  AOI21_X1 U48324 ( .B1(n46710), .B2(n46709), .A(n51396), .ZN(n46711) );
  OAI211_X1 U48325 ( .C1(n46714), .C2(n46713), .A(n46712), .B(n46711), .ZN(
        n46717) );
  NAND2_X1 U48326 ( .A1(n46871), .A2(n47104), .ZN(n46729) );
  NAND2_X1 U48327 ( .A1(n47095), .A2(n46719), .ZN(n46720) );
  NAND2_X1 U48328 ( .A1(n47089), .A2(n51341), .ZN(n46723) );
  OR2_X1 U48329 ( .A1(n47088), .A2(n46721), .ZN(n46722) );
  AND3_X1 U48330 ( .A1(n46724), .A2(n46723), .A3(n46722), .ZN(n46728) );
  OAI211_X1 U48331 ( .C1(n51341), .C2(n669), .A(n46725), .B(n47109), .ZN(
        n46726) );
  NOR2_X1 U48333 ( .A1(n47505), .A2(n47527), .ZN(n46780) );
  OR2_X1 U48334 ( .A1(n46731), .A2(n46730), .ZN(n46734) );
  OAI211_X1 U48335 ( .C1(n46735), .C2(n46734), .A(n46733), .B(n46732), .ZN(
        n46736) );
  INV_X1 U48336 ( .A(n46736), .ZN(n46764) );
  NAND2_X1 U48337 ( .A1(n46739), .A2(n46737), .ZN(n46742) );
  NAND2_X1 U48338 ( .A1(n46739), .A2(n46738), .ZN(n46741) );
  MUX2_X1 U48339 ( .A(n46742), .B(n46741), .S(n46740), .Z(n46763) );
  NAND2_X1 U48340 ( .A1(n46753), .A2(n46746), .ZN(n46748) );
  AOI21_X1 U48341 ( .B1(n46748), .B2(n46747), .A(n44850), .ZN(n46750) );
  OAI21_X1 U48342 ( .B1(n46751), .B2(n46750), .A(n46749), .ZN(n46762) );
  MUX2_X1 U48343 ( .A(n50965), .B(n46756), .S(n46753), .Z(n46760) );
  NAND2_X1 U48344 ( .A1(n46756), .A2(n46755), .ZN(n46752) );
  OAI21_X1 U48345 ( .B1(n46753), .B2(n46756), .A(n46752), .ZN(n46754) );
  OAI21_X1 U48346 ( .B1(n46756), .B2(n46755), .A(n50965), .ZN(n46757) );
  INV_X1 U48347 ( .A(n46814), .ZN(n46768) );
  NOR2_X1 U48348 ( .A1(n47073), .A2(n46770), .ZN(n46783) );
  OAI21_X1 U48349 ( .B1(n47073), .B2(n46772), .A(n46784), .ZN(n46773) );
  NOR2_X1 U48350 ( .A1(n46783), .A2(n46773), .ZN(n46779) );
  OR2_X1 U48351 ( .A1(n7046), .A2(n46774), .ZN(n47070) );
  INV_X1 U48352 ( .A(n47070), .ZN(n46776) );
  OAI21_X1 U48353 ( .B1(n46776), .B2(n400), .A(n46775), .ZN(n46777) );
  AND2_X1 U48354 ( .A1(n46778), .A2(n46777), .ZN(n46785) );
  NOR2_X1 U48355 ( .A1(n51346), .A2(n47573), .ZN(n47514) );
  AND2_X1 U48356 ( .A1(n47563), .A2(n51302), .ZN(n46793) );
  INV_X1 U48357 ( .A(n46783), .ZN(n46786) );
  NAND3_X1 U48358 ( .A1(n46786), .A2(n46785), .A3(n46784), .ZN(n46787) );
  OAI21_X1 U48359 ( .B1(n52044), .B2(n47554), .A(n414), .ZN(n46789) );
  OAI21_X1 U48360 ( .B1(n51290), .B2(n47574), .A(n46789), .ZN(n46790) );
  AND2_X1 U48361 ( .A1(n47570), .A2(n47571), .ZN(n47502) );
  NAND3_X1 U48363 ( .A1(n47505), .A2(n51346), .A3(n47542), .ZN(n46792) );
  OAI211_X1 U48364 ( .C1(n52045), .C2(n51302), .A(n47542), .B(n51289), .ZN(
        n46791) );
  AND3_X1 U48365 ( .A1(n51346), .A2(n46793), .A3(n47573), .ZN(n47580) );
  NOR2_X1 U48366 ( .A1(n47539), .A2(n51346), .ZN(n46794) );
  MUX2_X1 U48367 ( .A(n47580), .B(n46794), .S(n51286), .Z(n46795) );
  INV_X1 U48368 ( .A(n46800), .ZN(n46801) );
  NAND2_X1 U48369 ( .A1(n46801), .A2(n46977), .ZN(n46809) );
  NAND2_X1 U48370 ( .A1(n46803), .A2(n46802), .ZN(n46804) );
  OAI211_X1 U48371 ( .C1(n50367), .C2(n50361), .A(n46804), .B(n46975), .ZN(
        n46808) );
  INV_X1 U48372 ( .A(n46805), .ZN(n47141) );
  NAND2_X1 U48373 ( .A1(n46806), .A2(n47141), .ZN(n46807) );
  AND3_X1 U48375 ( .A1(n46814), .A2(n46815), .A3(n46813), .ZN(n46837) );
  OR2_X1 U48376 ( .A1(n51292), .A2(n7046), .ZN(n46820) );
  INV_X1 U48377 ( .A(n46817), .ZN(n46818) );
  NAND3_X1 U48378 ( .A1(n46818), .A2(n46822), .A3(n47069), .ZN(n46819) );
  OAI21_X1 U48379 ( .B1(n47071), .B2(n46820), .A(n46819), .ZN(n46821) );
  INV_X1 U48380 ( .A(n46821), .ZN(n46836) );
  NAND2_X1 U48381 ( .A1(n46822), .A2(n47074), .ZN(n46827) );
  NAND2_X1 U48382 ( .A1(n46824), .A2(n46823), .ZN(n46826) );
  INV_X1 U48383 ( .A(n400), .ZN(n46825) );
  NAND3_X1 U48384 ( .A1(n46827), .A2(n46826), .A3(n46825), .ZN(n46829) );
  NAND2_X1 U48385 ( .A1(n46829), .A2(n51304), .ZN(n46835) );
  OAI22_X1 U48386 ( .A1(n46831), .A2(n51419), .B1(n47075), .B2(n51456), .ZN(
        n46833) );
  NAND2_X1 U48387 ( .A1(n46833), .A2(n46832), .ZN(n46834) );
  NAND4_X2 U48388 ( .A1(n46837), .A2(n46836), .A3(n46835), .A4(n46834), .ZN(
        n50837) );
  NAND2_X1 U48389 ( .A1(n46839), .A2(n46838), .ZN(n46843) );
  NAND2_X1 U48390 ( .A1(n47123), .A2(n47122), .ZN(n46841) );
  NAND3_X1 U48391 ( .A1(n46841), .A2(n46840), .A3(n47118), .ZN(n47131) );
  MUX2_X1 U48392 ( .A(n46843), .B(n47131), .S(n46842), .Z(n46868) );
  OR2_X1 U48393 ( .A1(n46845), .A2(n46844), .ZN(n46851) );
  NAND3_X1 U48394 ( .A1(n46847), .A2(n46859), .A3(n46846), .ZN(n46850) );
  OAI21_X1 U48395 ( .B1(n46859), .B2(n47127), .A(n47126), .ZN(n46848) );
  NAND2_X1 U48396 ( .A1(n46848), .A2(n47129), .ZN(n46849) );
  OAI211_X1 U48397 ( .C1(n46852), .C2(n46851), .A(n46850), .B(n46849), .ZN(
        n46853) );
  INV_X1 U48398 ( .A(n46853), .ZN(n46867) );
  NAND2_X1 U48399 ( .A1(n46854), .A2(n47129), .ZN(n46856) );
  NAND3_X1 U48400 ( .A1(n47124), .A2(n52053), .A3(n47126), .ZN(n46855) );
  NAND3_X1 U48401 ( .A1(n46857), .A2(n46856), .A3(n46855), .ZN(n46858) );
  NAND2_X1 U48402 ( .A1(n46858), .A2(n47127), .ZN(n46866) );
  NAND2_X1 U48403 ( .A1(n47124), .A2(n46859), .ZN(n46862) );
  NAND2_X1 U48404 ( .A1(n46860), .A2(n47128), .ZN(n46861) );
  NAND2_X1 U48405 ( .A1(n46864), .A2(n46863), .ZN(n46865) );
  NAND4_X2 U48406 ( .A1(n46867), .A2(n46868), .A3(n46866), .A4(n46865), .ZN(
        n50850) );
  NAND2_X1 U48407 ( .A1(n50848), .A2(n50850), .ZN(n50873) );
  NOR2_X1 U48408 ( .A1(n46872), .A2(n51341), .ZN(n46870) );
  NOR2_X1 U48409 ( .A1(n46871), .A2(n46870), .ZN(n46887) );
  MUX2_X1 U48410 ( .A(n2159), .B(n47088), .S(n46872), .Z(n46874) );
  NAND2_X1 U48411 ( .A1(n46874), .A2(n46873), .ZN(n46876) );
  NAND2_X1 U48412 ( .A1(n46876), .A2(n46875), .ZN(n46886) );
  NAND2_X1 U48413 ( .A1(n46879), .A2(n7919), .ZN(n46885) );
  AND2_X1 U48414 ( .A1(n47087), .A2(n2159), .ZN(n46883) );
  AND2_X1 U48415 ( .A1(n47111), .A2(n47096), .ZN(n46882) );
  NOR2_X1 U48417 ( .A1(n51312), .A2(n50850), .ZN(n50853) );
  AND2_X1 U48418 ( .A1(n50837), .A2(n50826), .ZN(n50829) );
  AOI21_X1 U48419 ( .B1(n46994), .B2(n389), .A(n43683), .ZN(n46898) );
  OAI22_X1 U48420 ( .A1(n47154), .A2(n46889), .B1(n46888), .B2(n47153), .ZN(
        n46897) );
  INV_X1 U48421 ( .A(n46890), .ZN(n46892) );
  INV_X1 U48422 ( .A(n47150), .ZN(n46891) );
  NOR2_X1 U48423 ( .A1(n43683), .A2(n46999), .ZN(n46893) );
  OAI211_X1 U48424 ( .C1(n46894), .C2(n46893), .A(n2751), .B(n47154), .ZN(
        n46895) );
  NAND2_X1 U48425 ( .A1(n46900), .A2(n51513), .ZN(n46909) );
  NAND2_X1 U48426 ( .A1(n46902), .A2(n46901), .ZN(n46907) );
  NAND3_X1 U48427 ( .A1(n46905), .A2(n46904), .A3(n46903), .ZN(n46906) );
  NAND4_X1 U48428 ( .A1(n46909), .A2(n46908), .A3(n46907), .A4(n46906), .ZN(
        n46911) );
  AND2_X1 U48429 ( .A1(n46911), .A2(n46910), .ZN(n46926) );
  AOI21_X1 U48431 ( .B1(n46917), .B2(n46916), .A(n46915), .ZN(n46924) );
  OAI21_X1 U48432 ( .B1(n46922), .B2(n46921), .A(n46920), .ZN(n46923) );
  AND2_X1 U48433 ( .A1(n50865), .A2(n50826), .ZN(n50872) );
  INV_X1 U48434 ( .A(n50854), .ZN(n50863) );
  INV_X1 U48435 ( .A(n50864), .ZN(n46927) );
  INV_X1 U48436 ( .A(n50837), .ZN(n50890) );
  OR2_X1 U48437 ( .A1(n50865), .A2(n601), .ZN(n50861) );
  AOI21_X1 U48438 ( .B1(n50861), .B2(n50890), .A(n50894), .ZN(n46929) );
  OAI21_X1 U48439 ( .B1(n50851), .B2(n50831), .A(n46929), .ZN(n46931) );
  NOR2_X1 U48440 ( .A1(n50850), .A2(n50826), .ZN(n50883) );
  AND2_X1 U48441 ( .A1(n601), .A2(n52098), .ZN(n50888) );
  OAI21_X1 U48442 ( .B1(n50851), .B2(n50883), .A(n50888), .ZN(n46930) );
  INV_X1 U48443 ( .A(n4890), .ZN(n46932) );
  AND2_X1 U48444 ( .A1(n49021), .A2(n49037), .ZN(n49006) );
  AND2_X1 U48445 ( .A1(n49004), .A2(n49006), .ZN(n48987) );
  NAND2_X1 U48446 ( .A1(n49019), .A2(n49020), .ZN(n46933) );
  NAND2_X1 U48447 ( .A1(n49003), .A2(n51397), .ZN(n48994) );
  NAND2_X1 U48448 ( .A1(n46935), .A2(n6389), .ZN(n46940) );
  NAND2_X1 U48449 ( .A1(n49007), .A2(n51397), .ZN(n49025) );
  AND2_X1 U48451 ( .A1(n46279), .A2(n49021), .ZN(n49040) );
  NAND2_X1 U48452 ( .A1(n52179), .A2(n49037), .ZN(n49017) );
  INV_X1 U48453 ( .A(n49008), .ZN(n49044) );
  AND2_X1 U48454 ( .A1(n51397), .A2(n49020), .ZN(n49046) );
  OAI211_X1 U48455 ( .C1(n49040), .C2(n49017), .A(n49044), .B(n49046), .ZN(
        n46938) );
  NAND4_X1 U48456 ( .A1(n46941), .A2(n46940), .A3(n46939), .A4(n46938), .ZN(
        n46943) );
  INV_X1 U48457 ( .A(n4884), .ZN(n46942) );
  XNOR2_X1 U48458 ( .A(n46943), .B(n46942), .ZN(Plaintext[95]) );
  OAI21_X1 U48459 ( .B1(n48975), .B2(n48944), .A(n48958), .ZN(n48937) );
  INV_X1 U48460 ( .A(n48937), .ZN(n46944) );
  NAND2_X1 U48461 ( .A1(n46944), .A2(n48972), .ZN(n46949) );
  INV_X1 U48462 ( .A(n48934), .ZN(n46948) );
  NAND3_X1 U48463 ( .A1(n48954), .A2(n46951), .A3(n48931), .ZN(n46947) );
  NAND2_X1 U48464 ( .A1(n48973), .A2(n51478), .ZN(n48932) );
  INV_X1 U48465 ( .A(n48932), .ZN(n46945) );
  NAND4_X1 U48466 ( .A1(n46949), .A2(n46948), .A3(n46947), .A4(n46946), .ZN(
        n46962) );
  NAND2_X1 U48468 ( .A1(n51511), .A2(n48957), .ZN(n46956) );
  NAND2_X1 U48469 ( .A1(n48973), .A2(n48935), .ZN(n46953) );
  NAND2_X1 U48470 ( .A1(n48935), .A2(n47477), .ZN(n48928) );
  INV_X1 U48471 ( .A(n48928), .ZN(n46958) );
  NAND2_X1 U48472 ( .A1(n46958), .A2(n51511), .ZN(n47482) );
  NAND4_X1 U48473 ( .A1(n46960), .A2(n46959), .A3(n47482), .A4(n48981), .ZN(
        n46961) );
  NAND2_X1 U48474 ( .A1(n50007), .A2(n49996), .ZN(n46963) );
  MUX2_X1 U48475 ( .A(n46963), .B(n2489), .S(n50015), .Z(n46966) );
  OR2_X1 U48476 ( .A1(n50325), .A2(n50315), .ZN(n46964) );
  OAI211_X1 U48477 ( .C1(n50329), .C2(n50010), .A(n46964), .B(n47368), .ZN(
        n46965) );
  AND2_X1 U48478 ( .A1(n50321), .A2(n50325), .ZN(n46967) );
  NOR2_X1 U48479 ( .A1(n50330), .A2(n52224), .ZN(n46968) );
  OAI211_X1 U48480 ( .C1(n51421), .C2(n46971), .A(n46970), .B(n50370), .ZN(
        n46972) );
  AOI22_X1 U48481 ( .A1(n47141), .A2(n46973), .B1(n46972), .B2(n47137), .ZN(
        n46993) );
  NOR2_X1 U48482 ( .A1(n47135), .A2(n50364), .ZN(n46976) );
  NOR2_X1 U48483 ( .A1(n50372), .A2(n51421), .ZN(n46974) );
  AOI22_X1 U48484 ( .A1(n46977), .A2(n46976), .B1(n46975), .B2(n46974), .ZN(
        n46992) );
  AOI21_X1 U48485 ( .B1(n47144), .B2(n46979), .A(n43798), .ZN(n46981) );
  NAND2_X1 U48486 ( .A1(n50361), .A2(n46984), .ZN(n46980) );
  OAI21_X1 U48487 ( .B1(n46983), .B2(n46982), .A(n50370), .ZN(n46986) );
  NAND3_X1 U48488 ( .A1(n46984), .A2(n667), .A3(n50363), .ZN(n46985) );
  NAND2_X1 U48489 ( .A1(n46986), .A2(n46985), .ZN(n46987) );
  NAND3_X1 U48491 ( .A1(n47143), .A2(n47139), .A3(n51421), .ZN(n46990) );
  NAND3_X1 U48492 ( .A1(n46995), .A2(n46994), .A3(n47159), .ZN(n47009) );
  OAI211_X1 U48493 ( .C1(n47159), .C2(n46998), .A(n47150), .B(n47161), .ZN(
        n47008) );
  NAND2_X1 U48494 ( .A1(n46997), .A2(n47154), .ZN(n47005) );
  NAND2_X1 U48495 ( .A1(n47159), .A2(n46998), .ZN(n47002) );
  NAND2_X1 U48496 ( .A1(n47000), .A2(n46999), .ZN(n47001) );
  AOI22_X1 U48497 ( .A1(n47006), .A2(n47005), .B1(n47004), .B2(n47003), .ZN(
        n47007) );
  AND4_X2 U48498 ( .A1(n47010), .A2(n47009), .A3(n47008), .A4(n47007), .ZN(
        n50550) );
  NAND2_X1 U48499 ( .A1(n47019), .A2(n51058), .ZN(n50039) );
  AOI21_X1 U48500 ( .B1(n47310), .B2(n2199), .A(n49742), .ZN(n47011) );
  NOR2_X1 U48501 ( .A1(n50375), .A2(n49731), .ZN(n50385) );
  NOR2_X1 U48502 ( .A1(n47013), .A2(n51058), .ZN(n49730) );
  AND2_X1 U48503 ( .A1(n49743), .A2(n47013), .ZN(n50035) );
  NAND3_X1 U48504 ( .A1(n50035), .A2(n423), .A3(n2199), .ZN(n47014) );
  INV_X1 U48505 ( .A(n49740), .ZN(n47016) );
  NAND2_X1 U48506 ( .A1(n47016), .A2(n49742), .ZN(n47314) );
  NAND2_X1 U48507 ( .A1(n50378), .A2(n49738), .ZN(n47017) );
  AND2_X1 U48508 ( .A1(n47314), .A2(n47017), .ZN(n47020) );
  NAND3_X1 U48509 ( .A1(n47019), .A2(n47018), .A3(n49743), .ZN(n49744) );
  NAND2_X1 U48510 ( .A1(n50550), .A2(n50533), .ZN(n50563) );
  OR2_X1 U48511 ( .A1(n47273), .A2(n51725), .ZN(n47277) );
  NAND2_X1 U48512 ( .A1(n50337), .A2(n50348), .ZN(n47021) );
  NOR2_X1 U48513 ( .A1(n47277), .A2(n47021), .ZN(n47025) );
  NAND2_X1 U48514 ( .A1(n47275), .A2(n47289), .ZN(n47022) );
  OAI211_X1 U48515 ( .C1(n51025), .C2(n47023), .A(n47022), .B(n47282), .ZN(
        n47024) );
  NOR2_X1 U48516 ( .A1(n47025), .A2(n47024), .ZN(n47038) );
  INV_X1 U48517 ( .A(n50351), .ZN(n47027) );
  NAND2_X1 U48518 ( .A1(n47027), .A2(n49961), .ZN(n49969) );
  NAND2_X1 U48519 ( .A1(n47028), .A2(n50349), .ZN(n47029) );
  AOI21_X1 U48520 ( .B1(n49969), .B2(n47029), .A(n51725), .ZN(n47036) );
  OAI211_X1 U48521 ( .C1(n49961), .C2(n47030), .A(n51725), .B(n51386), .ZN(
        n47034) );
  OAI211_X1 U48522 ( .C1(n50352), .C2(n50349), .A(n51725), .B(n50351), .ZN(
        n47033) );
  NAND3_X1 U48523 ( .A1(n44608), .A2(n51725), .A3(n47031), .ZN(n47032) );
  NAND3_X1 U48524 ( .A1(n47034), .A2(n47033), .A3(n47032), .ZN(n47035) );
  NOR2_X1 U48525 ( .A1(n47036), .A2(n47035), .ZN(n47037) );
  INV_X1 U48528 ( .A(n47042), .ZN(n47043) );
  NAND2_X1 U48529 ( .A1(n47043), .A2(n50280), .ZN(n47048) );
  NAND2_X1 U48530 ( .A1(n47058), .A2(n44001), .ZN(n47045) );
  NAND2_X1 U48532 ( .A1(n50269), .A2(n47058), .ZN(n47047) );
  INV_X1 U48534 ( .A(n50526), .ZN(n47049) );
  OR2_X1 U48535 ( .A1(n50521), .A2(n50520), .ZN(n50527) );
  NAND4_X1 U48536 ( .A1(n47049), .A2(n50564), .A3(n50542), .A4(n50527), .ZN(
        n47050) );
  AND2_X1 U48537 ( .A1(n47050), .A2(n50494), .ZN(n47054) );
  INV_X1 U48538 ( .A(n50552), .ZN(n50508) );
  OAI21_X1 U48539 ( .B1(n50564), .B2(n50533), .A(n50508), .ZN(n50525) );
  NAND3_X1 U48540 ( .A1(n50541), .A2(n50525), .A3(n50521), .ZN(n47053) );
  AND2_X1 U48541 ( .A1(n50564), .A2(n50552), .ZN(n50534) );
  NOR2_X1 U48542 ( .A1(n50555), .A2(n50533), .ZN(n47051) );
  AND2_X1 U48543 ( .A1(n50520), .A2(n50552), .ZN(n50490) );
  NAND4_X1 U48544 ( .A1(n47055), .A2(n47054), .A3(n47053), .A4(n47052), .ZN(
        n47057) );
  INV_X1 U48545 ( .A(n4482), .ZN(n47056) );
  XNOR2_X1 U48546 ( .A(n47057), .B(n47056), .ZN(Plaintext[156]) );
  NOR2_X1 U48547 ( .A1(n47335), .A2(n51372), .ZN(n47059) );
  AND2_X1 U48548 ( .A1(n50277), .A2(n50280), .ZN(n50275) );
  OAI21_X1 U48549 ( .B1(n47065), .B2(n47059), .A(n50275), .ZN(n47063) );
  NAND2_X1 U48550 ( .A1(n47335), .A2(n50281), .ZN(n47060) );
  NAND2_X1 U48551 ( .A1(n47065), .A2(n50251), .ZN(n47066) );
  MUX2_X1 U48552 ( .A(n47334), .B(n50279), .S(n47333), .Z(n50260) );
  NAND3_X1 U48553 ( .A1(n50260), .A2(n50259), .A3(n50276), .ZN(n47348) );
  NAND2_X1 U48554 ( .A1(n47069), .A2(n51419), .ZN(n47072) );
  OAI22_X1 U48555 ( .A1(n47073), .A2(n47072), .B1(n47071), .B2(n47070), .ZN(
        n47083) );
  XNOR2_X1 U48556 ( .A(n47074), .B(n7046), .ZN(n47077) );
  OAI21_X1 U48557 ( .B1(n47077), .B2(n47076), .A(n47075), .ZN(n47081) );
  NAND3_X1 U48558 ( .A1(n51419), .A2(n400), .A3(n661), .ZN(n47079) );
  NAND3_X1 U48559 ( .A1(n47081), .A2(n47080), .A3(n47079), .ZN(n47082) );
  NAND2_X1 U48560 ( .A1(n47086), .A2(n47104), .ZN(n47092) );
  NAND3_X1 U48561 ( .A1(n47089), .A2(n47106), .A3(n47088), .ZN(n47091) );
  NAND3_X1 U48562 ( .A1(n47094), .A2(n47093), .A3(n7332), .ZN(n47102) );
  INV_X1 U48563 ( .A(n47095), .ZN(n47097) );
  NAND3_X1 U48564 ( .A1(n47097), .A2(n47098), .A3(n47096), .ZN(n47100) );
  NAND2_X1 U48565 ( .A1(n47098), .A2(n7332), .ZN(n47099) );
  INV_X1 U48566 ( .A(n47103), .ZN(n47107) );
  OAI211_X1 U48567 ( .C1(n47107), .C2(n47106), .A(n47105), .B(n47104), .ZN(
        n47116) );
  NOR2_X1 U48568 ( .A1(n47111), .A2(n47110), .ZN(n47113) );
  OAI21_X1 U48569 ( .B1(n47114), .B2(n47113), .A(n47112), .ZN(n47115) );
  NAND2_X1 U48570 ( .A1(n50786), .A2(n2095), .ZN(n50815) );
  NAND3_X1 U48571 ( .A1(n47119), .A2(n47127), .A3(n47118), .ZN(n47120) );
  OAI21_X1 U48572 ( .B1(n47123), .B2(n52053), .A(n47121), .ZN(n47125) );
  NAND2_X1 U48573 ( .A1(n47125), .A2(n47124), .ZN(n47132) );
  NAND4_X1 U48574 ( .A1(n47129), .A2(n47128), .A3(n47127), .A4(n47126), .ZN(
        n47130) );
  OAI22_X1 U48575 ( .A1(n47136), .A2(n50361), .B1(n47135), .B2(n50363), .ZN(
        n47138) );
  INV_X1 U48576 ( .A(n47139), .ZN(n50371) );
  AND2_X1 U48577 ( .A1(n43798), .A2(n50366), .ZN(n47140) );
  AOI22_X1 U48578 ( .A1(n47142), .A2(n47141), .B1(n50371), .B2(n47140), .ZN(
        n47148) );
  NAND2_X1 U48579 ( .A1(n47143), .A2(n667), .ZN(n47147) );
  OR2_X1 U48580 ( .A1(n51730), .A2(n50808), .ZN(n50811) );
  AND2_X1 U48581 ( .A1(n47151), .A2(n47152), .ZN(n47158) );
  OR2_X1 U48582 ( .A1(n47154), .A2(n47153), .ZN(n47155) );
  AOI21_X1 U48583 ( .B1(n47158), .B2(n47157), .A(n47156), .ZN(n47166) );
  OAI211_X1 U48584 ( .C1(n47164), .C2(n43683), .A(n47163), .B(n47162), .ZN(
        n47165) );
  NOR2_X1 U48585 ( .A1(n50779), .A2(n50809), .ZN(n47167) );
  NAND2_X1 U48587 ( .A1(n51296), .A2(n50772), .ZN(n50783) );
  INV_X1 U48588 ( .A(n50783), .ZN(n50762) );
  OAI21_X1 U48589 ( .B1(n47167), .B2(n50804), .A(n50762), .ZN(n47171) );
  NOR2_X1 U48590 ( .A1(n51296), .A2(n51730), .ZN(n50764) );
  NAND3_X1 U48591 ( .A1(n50764), .A2(n52076), .A3(n2095), .ZN(n47170) );
  NOR2_X1 U48592 ( .A1(n50771), .A2(n50772), .ZN(n50797) );
  NAND3_X1 U48593 ( .A1(n50798), .A2(n52076), .A3(n50797), .ZN(n47169) );
  NAND2_X1 U48594 ( .A1(n50751), .A2(n51296), .ZN(n50761) );
  NAND3_X1 U48595 ( .A1(n50761), .A2(n51354), .A3(n51730), .ZN(n47168) );
  AND4_X1 U48596 ( .A1(n47171), .A2(n47170), .A3(n47169), .A4(n47168), .ZN(
        n47176) );
  AND2_X1 U48597 ( .A1(n50773), .A2(n50772), .ZN(n50752) );
  OR2_X1 U48598 ( .A1(n50752), .A2(n50781), .ZN(n47172) );
  OAI21_X1 U48599 ( .B1(n47172), .B2(n50797), .A(n50751), .ZN(n47173) );
  OR2_X1 U48600 ( .A1(n51354), .A2(n51730), .ZN(n47183) );
  NAND4_X1 U48601 ( .A1(n47174), .A2(n47173), .A3(n50808), .A4(n47183), .ZN(
        n47175) );
  OAI211_X1 U48602 ( .C1(n50815), .C2(n50811), .A(n47176), .B(n47175), .ZN(
        n47178) );
  INV_X1 U48603 ( .A(n4325), .ZN(n47177) );
  XNOR2_X1 U48604 ( .A(n47178), .B(n47177), .ZN(Plaintext[174]) );
  AOI21_X1 U48605 ( .B1(n47179), .B2(n50781), .A(n51353), .ZN(n47181) );
  OR2_X1 U48606 ( .A1(n50751), .A2(n50787), .ZN(n50747) );
  NAND2_X1 U48607 ( .A1(n50798), .A2(n51296), .ZN(n47180) );
  NAND4_X1 U48608 ( .A1(n47182), .A2(n47181), .A3(n50747), .A4(n47180), .ZN(
        n47186) );
  AND2_X1 U48609 ( .A1(n2095), .A2(n50809), .ZN(n47184) );
  OAI211_X1 U48610 ( .C1(n50798), .C2(n51730), .A(n47184), .B(n47183), .ZN(
        n47185) );
  OAI211_X1 U48611 ( .C1(n50783), .C2(n51730), .A(n47186), .B(n47185), .ZN(
        n47190) );
  NAND4_X1 U48612 ( .A1(n50798), .A2(n50781), .A3(n51354), .A4(n50808), .ZN(
        n50739) );
  AND2_X1 U48613 ( .A1(n51354), .A2(n50809), .ZN(n47187) );
  OAI21_X1 U48614 ( .B1(n50773), .B2(n50739), .A(n47188), .ZN(n47189) );
  NOR2_X1 U48615 ( .A1(n47190), .A2(n47189), .ZN(n47191) );
  XNOR2_X1 U48616 ( .A(n47191), .B(n4627), .ZN(Plaintext[179]) );
  NOR2_X1 U48618 ( .A1(n49443), .A2(n52107), .ZN(n49409) );
  AND2_X1 U48619 ( .A1(n49452), .A2(n51315), .ZN(n47200) );
  OAI211_X1 U48620 ( .C1(n49461), .C2(n51516), .A(n47196), .B(n47200), .ZN(
        n47198) );
  INV_X1 U48621 ( .A(n47200), .ZN(n49417) );
  NAND2_X1 U48622 ( .A1(n49445), .A2(n51315), .ZN(n49403) );
  AND2_X1 U48623 ( .A1(n49461), .A2(n49403), .ZN(n49441) );
  AND2_X1 U48624 ( .A1(n49443), .A2(n49465), .ZN(n49458) );
  OR2_X1 U48625 ( .A1(n47203), .A2(n49458), .ZN(n49440) );
  NAND2_X1 U48626 ( .A1(n49445), .A2(n52107), .ZN(n49424) );
  INV_X1 U48627 ( .A(n2231), .ZN(n47205) );
  NAND2_X1 U48628 ( .A1(n47206), .A2(n47586), .ZN(n47610) );
  XNOR2_X1 U48629 ( .A(n47618), .B(n8448), .ZN(n47207) );
  NOR2_X1 U48630 ( .A1(n47617), .A2(n47620), .ZN(n47595) );
  NAND2_X1 U48631 ( .A1(n47257), .A2(n47595), .ZN(n47208) );
  OAI211_X1 U48632 ( .C1(n47610), .C2(n47616), .A(n47209), .B(n47208), .ZN(
        n47215) );
  NAND2_X1 U48634 ( .A1(n8448), .A2(n47586), .ZN(n47256) );
  NAND3_X1 U48635 ( .A1(n47210), .A2(n47256), .A3(n47618), .ZN(n47211) );
  NAND3_X1 U48636 ( .A1(n47463), .A2(n47266), .A3(n47617), .ZN(n47606) );
  INV_X1 U48637 ( .A(n47618), .ZN(n47461) );
  NAND2_X1 U48638 ( .A1(n47461), .A2(n52158), .ZN(n47212) );
  NOR2_X1 U48639 ( .A1(n47215), .A2(n47214), .ZN(n47216) );
  XNOR2_X1 U48640 ( .A(n47216), .B(n842), .ZN(Plaintext[6]) );
  NOR2_X1 U48641 ( .A1(n47217), .A2(n50611), .ZN(n47218) );
  NOR2_X1 U48642 ( .A1(n52225), .A2(n51029), .ZN(n50634) );
  OAI21_X1 U48643 ( .B1(n47218), .B2(n50634), .A(n50642), .ZN(n47219) );
  NAND2_X1 U48644 ( .A1(n47219), .A2(n50633), .ZN(n47225) );
  NOR2_X1 U48645 ( .A1(n50618), .A2(n50630), .ZN(n50573) );
  INV_X1 U48646 ( .A(n50631), .ZN(n47220) );
  OR3_X1 U48647 ( .A1(n50573), .A2(n47220), .A3(n50578), .ZN(n47224) );
  NAND2_X1 U48648 ( .A1(n50624), .A2(n47221), .ZN(n47222) );
  NAND2_X1 U48649 ( .A1(n47222), .A2(n50599), .ZN(n47223) );
  NAND4_X1 U48650 ( .A1(n47225), .A2(n47224), .A3(n47223), .A4(n50622), .ZN(
        n47227) );
  INV_X1 U48651 ( .A(n4800), .ZN(n47226) );
  XNOR2_X1 U48652 ( .A(n47227), .B(n47226), .ZN(Plaintext[164]) );
  NOR2_X1 U48653 ( .A1(n50929), .A2(n51299), .ZN(n50903) );
  NAND2_X1 U48654 ( .A1(n47391), .A2(n47228), .ZN(n47229) );
  OAI211_X1 U48655 ( .C1(n50903), .C2(n50913), .A(n47230), .B(n47229), .ZN(
        n47233) );
  NAND2_X1 U48656 ( .A1(n50913), .A2(n50955), .ZN(n47231) );
  AOI21_X1 U48657 ( .B1(n47231), .B2(n50958), .A(n50950), .ZN(n47232) );
  OR2_X1 U48658 ( .A1(n47233), .A2(n47232), .ZN(n47243) );
  NOR2_X1 U48659 ( .A1(n47236), .A2(n50906), .ZN(n50957) );
  NAND2_X1 U48660 ( .A1(n50957), .A2(n51298), .ZN(n50920) );
  OR2_X1 U48661 ( .A1(n50920), .A2(n5365), .ZN(n47242) );
  AND2_X1 U48662 ( .A1(n50958), .A2(n50950), .ZN(n50925) );
  AOI22_X1 U48663 ( .A1(n50903), .A2(n47391), .B1(n50925), .B2(n50928), .ZN(
        n47241) );
  OR2_X1 U48664 ( .A1(n50950), .A2(n50955), .ZN(n47234) );
  INV_X1 U48666 ( .A(n47236), .ZN(n50937) );
  AND3_X1 U48667 ( .A1(n50951), .A2(n5365), .A3(n50906), .ZN(n50947) );
  NAND2_X1 U48668 ( .A1(n50937), .A2(n50947), .ZN(n47238) );
  NAND3_X1 U48669 ( .A1(n50959), .A2(n50958), .A3(n50906), .ZN(n47237) );
  NAND2_X1 U48670 ( .A1(n47238), .A2(n47237), .ZN(n47239) );
  NOR2_X1 U48671 ( .A1(n50938), .A2(n47239), .ZN(n47240) );
  INV_X1 U48672 ( .A(n48702), .ZN(n48667) );
  AOI21_X1 U48673 ( .B1(n48667), .B2(n48687), .A(n48697), .ZN(n47246) );
  NOR2_X1 U48674 ( .A1(n48659), .A2(n52157), .ZN(n48707) );
  NAND2_X1 U48675 ( .A1(n48667), .A2(n48707), .ZN(n47245) );
  NAND2_X1 U48676 ( .A1(n52004), .A2(n48714), .ZN(n48711) );
  INV_X1 U48677 ( .A(n48711), .ZN(n47249) );
  AOI21_X1 U48679 ( .B1(n51291), .B2(n48659), .A(n47247), .ZN(n47248) );
  NAND2_X1 U48680 ( .A1(n47249), .A2(n47248), .ZN(n47254) );
  INV_X1 U48681 ( .A(n48688), .ZN(n47250) );
  NAND2_X1 U48682 ( .A1(n48659), .A2(n48697), .ZN(n48713) );
  INV_X1 U48683 ( .A(n48713), .ZN(n48675) );
  NAND3_X1 U48684 ( .A1(n47250), .A2(n52157), .A3(n48675), .ZN(n47253) );
  NOR2_X1 U48685 ( .A1(n48701), .A2(n51659), .ZN(n47413) );
  INV_X1 U48686 ( .A(n47413), .ZN(n47252) );
  NAND2_X1 U48687 ( .A1(n48659), .A2(n52157), .ZN(n48704) );
  NAND3_X1 U48688 ( .A1(n48687), .A2(n47407), .A3(n48704), .ZN(n47251) );
  NAND4_X1 U48689 ( .A1(n47254), .A2(n47253), .A3(n47252), .A4(n47251), .ZN(
        n47255) );
  OR3_X1 U48690 ( .A1(n47256), .A2(n47592), .A3(n47468), .ZN(n47264) );
  NOR2_X1 U48691 ( .A1(n8450), .A2(n2163), .ZN(n47259) );
  NOR2_X1 U48692 ( .A1(n47586), .A2(n2163), .ZN(n47258) );
  AOI22_X1 U48693 ( .A1(n47259), .A2(n8449), .B1(n47620), .B2(n47258), .ZN(
        n47262) );
  INV_X1 U48694 ( .A(n47619), .ZN(n47260) );
  NAND3_X1 U48695 ( .A1(n47260), .A2(n47617), .A3(n47468), .ZN(n47261) );
  NAND4_X1 U48696 ( .A1(n47264), .A2(n47263), .A3(n47262), .A4(n47261), .ZN(
        n47267) );
  XNOR2_X1 U48697 ( .A(n47269), .B(n47268), .ZN(Plaintext[7]) );
  NAND2_X1 U48698 ( .A1(n51025), .A2(n47271), .ZN(n50346) );
  NOR2_X1 U48699 ( .A1(n50346), .A2(n52062), .ZN(n47272) );
  AND2_X1 U48700 ( .A1(n47273), .A2(n47272), .ZN(n47274) );
  AOI22_X1 U48701 ( .A1(n47276), .A2(n47275), .B1(n47274), .B2(n47282), .ZN(
        n47299) );
  INV_X1 U48702 ( .A(n49961), .ZN(n49963) );
  NOR2_X1 U48703 ( .A1(n47277), .A2(n49963), .ZN(n47284) );
  NOR2_X1 U48704 ( .A1(n51725), .A2(n555), .ZN(n47279) );
  INV_X1 U48705 ( .A(n47279), .ZN(n47281) );
  NAND3_X1 U48706 ( .A1(n50352), .A2(n47279), .A3(n47278), .ZN(n47280) );
  OAI21_X1 U48707 ( .B1(n47282), .B2(n47281), .A(n47280), .ZN(n47283) );
  NOR2_X1 U48708 ( .A1(n47284), .A2(n47283), .ZN(n47298) );
  INV_X1 U48709 ( .A(n50342), .ZN(n49965) );
  NAND2_X1 U48710 ( .A1(n49965), .A2(n47294), .ZN(n47287) );
  INV_X1 U48711 ( .A(n47289), .ZN(n47285) );
  NAND3_X1 U48712 ( .A1(n50351), .A2(n51725), .A3(n47285), .ZN(n47286) );
  AOI22_X1 U48713 ( .A1(n47290), .A2(n47289), .B1(n51725), .B2(n47288), .ZN(
        n47292) );
  NAND3_X1 U48714 ( .A1(n50337), .A2(n47294), .A3(n47291), .ZN(n50341) );
  OAI211_X1 U48715 ( .C1(n47294), .C2(n47293), .A(n47292), .B(n50341), .ZN(
        n47295) );
  NAND2_X1 U48716 ( .A1(n47295), .A2(n50348), .ZN(n47296) );
  INV_X1 U48718 ( .A(n49639), .ZN(n49954) );
  NAND2_X1 U48719 ( .A1(n49954), .A2(n50307), .ZN(n47301) );
  OR2_X1 U48720 ( .A1(n49638), .A2(n49956), .ZN(n47300) );
  OR2_X1 U48723 ( .A1(n49637), .A2(n51300), .ZN(n47302) );
  NAND2_X1 U48724 ( .A1(n50299), .A2(n51691), .ZN(n47304) );
  NAND2_X1 U48725 ( .A1(n49956), .A2(n28), .ZN(n47306) );
  OAI211_X1 U48726 ( .C1(n51504), .C2(n50296), .A(n47307), .B(n47306), .ZN(
        n47308) );
  AND2_X1 U48727 ( .A1(n50233), .A2(n50189), .ZN(n50178) );
  AOI22_X1 U48728 ( .A1(n47310), .A2(n47309), .B1(n2199), .B2(n50378), .ZN(
        n47312) );
  INV_X1 U48729 ( .A(n49730), .ZN(n47311) );
  OR2_X1 U48730 ( .A1(n47312), .A2(n47311), .ZN(n47332) );
  NAND2_X1 U48731 ( .A1(n50035), .A2(n423), .ZN(n47313) );
  AND2_X1 U48732 ( .A1(n47314), .A2(n47313), .ZN(n47331) );
  INV_X1 U48733 ( .A(n49738), .ZN(n47315) );
  NAND2_X1 U48734 ( .A1(n49739), .A2(n47322), .ZN(n47319) );
  NAND2_X1 U48735 ( .A1(n2199), .A2(n51058), .ZN(n50379) );
  OAI21_X1 U48736 ( .B1(n50379), .B2(n47316), .A(n50377), .ZN(n47317) );
  INV_X1 U48737 ( .A(n47317), .ZN(n47318) );
  NAND3_X1 U48738 ( .A1(n47320), .A2(n47319), .A3(n47318), .ZN(n47325) );
  NAND3_X1 U48739 ( .A1(n47322), .A2(n49731), .A3(n47321), .ZN(n47323) );
  NAND2_X1 U48740 ( .A1(n47323), .A2(n50390), .ZN(n47324) );
  NAND2_X1 U48741 ( .A1(n47325), .A2(n47324), .ZN(n47330) );
  OAI21_X1 U48742 ( .B1(n47327), .B2(n50375), .A(n47326), .ZN(n47328) );
  NAND2_X1 U48743 ( .A1(n47328), .A2(n50390), .ZN(n47329) );
  OAI211_X1 U48744 ( .C1(n47335), .C2(n50259), .A(n658), .B(n47334), .ZN(
        n47338) );
  NAND2_X1 U48745 ( .A1(n50281), .A2(n50266), .ZN(n47337) );
  NAND3_X1 U48746 ( .A1(n50281), .A2(n47341), .A3(n50259), .ZN(n47336) );
  AND3_X1 U48747 ( .A1(n47338), .A2(n47337), .A3(n47336), .ZN(n47347) );
  NAND3_X1 U48748 ( .A1(n47340), .A2(n47339), .A3(n50277), .ZN(n47346) );
  OR2_X1 U48749 ( .A1(n50281), .A2(n50280), .ZN(n47343) );
  NAND2_X1 U48750 ( .A1(n47344), .A2(n50277), .ZN(n47345) );
  XNOR2_X1 U48751 ( .A(n51480), .B(n50192), .ZN(n47378) );
  NAND2_X1 U48752 ( .A1(n49618), .A2(n47352), .ZN(n47353) );
  NAND2_X1 U48753 ( .A1(n47353), .A2(n49973), .ZN(n47364) );
  NAND2_X1 U48754 ( .A1(n47355), .A2(n47354), .ZN(n47357) );
  OAI21_X1 U48755 ( .B1(n47357), .B2(n47356), .A(n49626), .ZN(n47358) );
  INV_X1 U48756 ( .A(n47358), .ZN(n47363) );
  NAND2_X1 U48757 ( .A1(n49629), .A2(n51326), .ZN(n47359) );
  AND3_X1 U48758 ( .A1(n47360), .A2(n49627), .A3(n47359), .ZN(n49625) );
  NAND2_X1 U48759 ( .A1(n49625), .A2(n47361), .ZN(n47362) );
  OAI21_X1 U48760 ( .B1(n50314), .B2(n50325), .A(n50329), .ZN(n47367) );
  OAI211_X1 U48761 ( .C1(n50329), .C2(n1812), .A(n50015), .B(n47368), .ZN(
        n47366) );
  MUX2_X1 U48762 ( .A(n47367), .B(n47366), .S(n52124), .Z(n47377) );
  NAND2_X1 U48763 ( .A1(n50320), .A2(n47369), .ZN(n50003) );
  NAND3_X1 U48764 ( .A1(n50325), .A2(n50008), .A3(n1812), .ZN(n47370) );
  NAND2_X1 U48765 ( .A1(n50003), .A2(n47370), .ZN(n47375) );
  NAND3_X1 U48766 ( .A1(n47371), .A2(n50006), .A3(n50010), .ZN(n47373) );
  NAND2_X1 U48767 ( .A1(n50325), .A2(n50314), .ZN(n47372) );
  NAND2_X1 U48768 ( .A1(n47373), .A2(n47372), .ZN(n47374) );
  NAND2_X1 U48769 ( .A1(n47378), .A2(n50227), .ZN(n47380) );
  NOR2_X1 U48770 ( .A1(n602), .A2(n50235), .ZN(n50161) );
  OAI21_X1 U48771 ( .B1(n50161), .B2(n50222), .A(n50227), .ZN(n47379) );
  AOI22_X1 U48772 ( .A1(n50178), .A2(n47380), .B1(n47379), .B2(n5799), .ZN(
        n47387) );
  INV_X1 U48773 ( .A(n47382), .ZN(n50209) );
  NAND2_X1 U48774 ( .A1(n50209), .A2(n50234), .ZN(n50198) );
  NAND3_X1 U48775 ( .A1(n50189), .A2(n50196), .A3(n50235), .ZN(n50180) );
  NOR2_X1 U48776 ( .A1(n47382), .A2(n50235), .ZN(n50210) );
  AOI22_X1 U48777 ( .A1(n50210), .A2(n602), .B1(n50233), .B2(n50235), .ZN(
        n47383) );
  NOR2_X1 U48778 ( .A1(n50189), .A2(n50192), .ZN(n50205) );
  NAND2_X1 U48779 ( .A1(n50205), .A2(n50233), .ZN(n50230) );
  NAND2_X1 U48780 ( .A1(n50235), .A2(n50196), .ZN(n50236) );
  OAI22_X1 U48781 ( .A1(n47383), .A2(n50234), .B1(n50230), .B2(n50236), .ZN(
        n47384) );
  NOR2_X1 U48782 ( .A1(n47385), .A2(n47384), .ZN(n47386) );
  INV_X1 U48783 ( .A(n4651), .ZN(n47388) );
  NOR2_X1 U48786 ( .A1(n5365), .A2(n50950), .ZN(n47390) );
  NAND2_X1 U48787 ( .A1(n47392), .A2(n47391), .ZN(n47393) );
  NAND3_X1 U48788 ( .A1(n47395), .A2(n47394), .A3(n47393), .ZN(n47400) );
  OAI211_X1 U48790 ( .C1(n50935), .C2(n47399), .A(n50933), .B(n47398), .ZN(
        n50945) );
  NOR2_X1 U48791 ( .A1(n47400), .A2(n50945), .ZN(n47402) );
  XNOR2_X1 U48792 ( .A(n47402), .B(n47401), .ZN(Plaintext[188]) );
  NAND2_X1 U48793 ( .A1(n48659), .A2(n48703), .ZN(n48708) );
  NOR2_X1 U48795 ( .A1(n48708), .A2(n48685), .ZN(n47406) );
  NOR2_X1 U48796 ( .A1(n47404), .A2(n47407), .ZN(n47405) );
  MUX2_X1 U48797 ( .A(n47406), .B(n47405), .S(n48667), .Z(n47418) );
  INV_X1 U48798 ( .A(n48687), .ZN(n47408) );
  AOI22_X1 U48799 ( .A1(n47408), .A2(n48685), .B1(n51291), .B2(n47407), .ZN(
        n47409) );
  NAND2_X1 U48800 ( .A1(n48702), .A2(n52157), .ZN(n48709) );
  OR2_X1 U48801 ( .A1(n48711), .A2(n48713), .ZN(n48677) );
  NAND3_X1 U48802 ( .A1(n48696), .A2(n47410), .A3(n48703), .ZN(n48663) );
  OAI211_X1 U48803 ( .C1(n47409), .C2(n48709), .A(n48677), .B(n48663), .ZN(
        n47417) );
  NOR2_X1 U48804 ( .A1(n47410), .A2(n48702), .ZN(n48666) );
  OAI21_X1 U48805 ( .B1(n51659), .B2(n48703), .A(n52157), .ZN(n47411) );
  OAI211_X1 U48806 ( .C1(n52157), .C2(n48685), .A(n48666), .B(n47411), .ZN(
        n47415) );
  NOR2_X1 U48807 ( .A1(n48682), .A2(n48659), .ZN(n47412) );
  NOR2_X1 U48808 ( .A1(n47413), .A2(n47412), .ZN(n47414) );
  OAI211_X1 U48809 ( .C1(n48682), .C2(n48688), .A(n47415), .B(n47414), .ZN(
        n47416) );
  NOR3_X1 U48810 ( .A1(n47418), .A2(n47417), .A3(n47416), .ZN(n47419) );
  XNOR2_X1 U48811 ( .A(n47419), .B(n4691), .ZN(Plaintext[61]) );
  NAND2_X1 U48812 ( .A1(n49909), .A2(n49889), .ZN(n49900) );
  NAND3_X1 U48813 ( .A1(n47423), .A2(n49923), .A3(n49894), .ZN(n49926) );
  INV_X1 U48814 ( .A(n49923), .ZN(n47424) );
  NAND2_X1 U48816 ( .A1(n49933), .A2(n652), .ZN(n49901) );
  NAND2_X1 U48817 ( .A1(n49901), .A2(n47420), .ZN(n47421) );
  NAND2_X1 U48818 ( .A1(n49903), .A2(n47421), .ZN(n47422) );
  OAI21_X1 U48819 ( .B1(n49900), .B2(n49926), .A(n47422), .ZN(n47433) );
  NOR2_X1 U48820 ( .A1(n47423), .A2(n49923), .ZN(n49930) );
  OAI21_X1 U48821 ( .B1(n49917), .B2(n47425), .A(n49930), .ZN(n47431) );
  NAND2_X1 U48822 ( .A1(n49892), .A2(n49894), .ZN(n49882) );
  NAND4_X1 U48823 ( .A1(n47425), .A2(n49928), .A3(n47424), .A4(n49882), .ZN(
        n47429) );
  AND2_X1 U48824 ( .A1(n49889), .A2(n49932), .ZN(n49919) );
  INV_X1 U48825 ( .A(n49919), .ZN(n49908) );
  NOR2_X1 U48828 ( .A1(n47433), .A2(n47432), .ZN(n47434) );
  XNOR2_X1 U48829 ( .A(n47434), .B(n4605), .ZN(Plaintext[135]) );
  INV_X1 U48830 ( .A(n48734), .ZN(n48762) );
  NAND2_X1 U48831 ( .A1(n47435), .A2(n48751), .ZN(n47449) );
  NAND2_X1 U48832 ( .A1(n48726), .A2(n47449), .ZN(n47436) );
  NAND2_X1 U48833 ( .A1(n47436), .A2(n48769), .ZN(n47439) );
  NAND3_X1 U48834 ( .A1(n48778), .A2(n52067), .A3(n48759), .ZN(n48763) );
  NAND4_X1 U48835 ( .A1(n47439), .A2(n47438), .A3(n48763), .A4(n47437), .ZN(
        n48773) );
  NAND2_X1 U48836 ( .A1(n47442), .A2(n48747), .ZN(n48780) );
  NAND4_X1 U48837 ( .A1(n48780), .A2(n48730), .A3(n48751), .A4(n48729), .ZN(
        n47440) );
  NAND2_X1 U48838 ( .A1(n47441), .A2(n47440), .ZN(n48777) );
  NAND2_X1 U48839 ( .A1(n48773), .A2(n48777), .ZN(n47458) );
  INV_X1 U48840 ( .A(n48745), .ZN(n47444) );
  NAND2_X1 U48841 ( .A1(n47442), .A2(n48751), .ZN(n48779) );
  NAND4_X1 U48842 ( .A1(n48779), .A2(n48729), .A3(n48778), .A4(n48762), .ZN(
        n47443) );
  NAND3_X1 U48843 ( .A1(n48747), .A2(n48722), .A3(n995), .ZN(n48764) );
  OAI211_X1 U48844 ( .C1(n48778), .C2(n47444), .A(n47443), .B(n48764), .ZN(
        n47448) );
  NOR2_X1 U48846 ( .A1(n48747), .A2(n48729), .ZN(n47445) );
  NAND4_X1 U48847 ( .A1(n47452), .A2(n48730), .A3(n47445), .A4(n48762), .ZN(
        n47446) );
  AND2_X1 U48850 ( .A1(n48778), .A2(n48759), .ZN(n48744) );
  INV_X1 U48852 ( .A(n48780), .ZN(n48770) );
  INV_X1 U48853 ( .A(n47449), .ZN(n47450) );
  NAND3_X1 U48854 ( .A1(n48770), .A2(n48769), .A3(n47450), .ZN(n47451) );
  AND2_X1 U48855 ( .A1(n48736), .A2(n47451), .ZN(n47456) );
  INV_X1 U48856 ( .A(n48760), .ZN(n47453) );
  OAI22_X1 U48857 ( .A1(n47453), .A2(n48730), .B1(n47452), .B2(n48769), .ZN(
        n47454) );
  NAND3_X1 U48858 ( .A1(n47454), .A2(n48734), .A3(n52067), .ZN(n47455) );
  INV_X1 U48859 ( .A(n47622), .ZN(n47466) );
  NAND3_X1 U48860 ( .A1(n47616), .A2(n47461), .A3(n8448), .ZN(n47465) );
  OR2_X1 U48861 ( .A1(n47462), .A2(n47618), .ZN(n47605) );
  NAND4_X1 U48862 ( .A1(n47466), .A2(n47465), .A3(n47605), .A4(n47464), .ZN(
        n47473) );
  MUX2_X1 U48863 ( .A(n47587), .B(n47468), .S(n51400), .Z(n47467) );
  NOR2_X1 U48864 ( .A1(n47467), .A2(n52158), .ZN(n47472) );
  INV_X1 U48865 ( .A(n2163), .ZN(n47613) );
  NOR2_X1 U48866 ( .A1(n47468), .A2(n8450), .ZN(n47469) );
  NOR3_X1 U48867 ( .A1(n47473), .A2(n47472), .A3(n47471), .ZN(n47474) );
  XNOR2_X1 U48868 ( .A(n47474), .B(n4647), .ZN(Plaintext[8]) );
  OAI211_X1 U48869 ( .C1(n51510), .C2(n48935), .A(n48955), .B(n48974), .ZN(
        n47475) );
  AOI21_X1 U48870 ( .B1(n51511), .B2(n47477), .A(n47476), .ZN(n47478) );
  AOI21_X1 U48871 ( .B1(n47479), .B2(n47476), .A(n47478), .ZN(n47480) );
  NAND2_X1 U48872 ( .A1(n47481), .A2(n48957), .ZN(n48943) );
  INV_X1 U48873 ( .A(n48950), .ZN(n48968) );
  AND3_X1 U48874 ( .A1(n48943), .A2(n47483), .A3(n47482), .ZN(n47486) );
  OR2_X1 U48875 ( .A1(n47528), .A2(n51303), .ZN(n47558) );
  OR2_X1 U48876 ( .A1(n47558), .A2(n47557), .ZN(n47550) );
  AND2_X1 U48877 ( .A1(n47573), .A2(n47570), .ZN(n47538) );
  AND2_X1 U48878 ( .A1(n47570), .A2(n52045), .ZN(n47501) );
  NAND3_X1 U48879 ( .A1(n47501), .A2(n47539), .A3(n47579), .ZN(n47489) );
  OAI21_X1 U48880 ( .B1(n47574), .B2(n414), .A(n51303), .ZN(n47487) );
  NAND2_X1 U48881 ( .A1(n47519), .A2(n47487), .ZN(n47488) );
  AND4_X1 U48882 ( .A1(n47489), .A2(n47490), .A3(n47550), .A4(n47488), .ZN(
        n47497) );
  NAND4_X1 U48883 ( .A1(n47541), .A2(n47542), .A3(n47574), .A4(n47570), .ZN(
        n47492) );
  NAND2_X1 U48884 ( .A1(n47541), .A2(n47502), .ZN(n47491) );
  AND2_X1 U48885 ( .A1(n52045), .A2(n51289), .ZN(n47511) );
  NAND2_X1 U48886 ( .A1(n47511), .A2(n47573), .ZN(n47530) );
  AND3_X1 U48887 ( .A1(n47492), .A2(n47491), .A3(n47530), .ZN(n47496) );
  NAND2_X1 U48888 ( .A1(n47571), .A2(n51289), .ZN(n47518) );
  OAI21_X1 U48889 ( .B1(n47539), .B2(n47570), .A(n47518), .ZN(n47493) );
  NOR2_X1 U48890 ( .A1(n51287), .A2(n52044), .ZN(n47556) );
  NAND3_X1 U48891 ( .A1(n47493), .A2(n47542), .A3(n47556), .ZN(n47495) );
  INV_X1 U48892 ( .A(n4926), .ZN(n47498) );
  AND2_X1 U48893 ( .A1(n47541), .A2(n47542), .ZN(n47546) );
  AOI22_X1 U48894 ( .A1(n47546), .A2(n51303), .B1(n47501), .B2(n47499), .ZN(
        n47508) );
  NAND2_X1 U48895 ( .A1(n47573), .A2(n51287), .ZN(n47500) );
  INV_X1 U48896 ( .A(n47501), .ZN(n47504) );
  INV_X1 U48897 ( .A(n47502), .ZN(n47503) );
  NAND3_X1 U48898 ( .A1(n47504), .A2(n47503), .A3(n47541), .ZN(n47507) );
  INV_X1 U48899 ( .A(n4517), .ZN(n47509) );
  XNOR2_X1 U48900 ( .A(n47510), .B(n47509), .ZN(Plaintext[2]) );
  INV_X1 U48901 ( .A(n47511), .ZN(n47513) );
  OR2_X1 U48902 ( .A1(n47573), .A2(n51289), .ZN(n47512) );
  NAND4_X1 U48903 ( .A1(n47513), .A2(n414), .A3(n51346), .A4(n47512), .ZN(
        n47517) );
  INV_X1 U48904 ( .A(n47558), .ZN(n47515) );
  NAND3_X1 U48905 ( .A1(n47515), .A2(n47514), .A3(n47572), .ZN(n47516) );
  OAI211_X1 U48906 ( .C1(n47542), .C2(n47518), .A(n47517), .B(n47516), .ZN(
        n47526) );
  NAND2_X1 U48907 ( .A1(n47519), .A2(n51289), .ZN(n47525) );
  NAND2_X1 U48908 ( .A1(n47526), .A2(n47525), .ZN(n47524) );
  OAI211_X1 U48909 ( .C1(n51286), .C2(n47527), .A(n4564), .B(n47530), .ZN(
        n47520) );
  NOR2_X1 U48910 ( .A1(n47521), .A2(n47520), .ZN(n47523) );
  AND2_X1 U48911 ( .A1(n52045), .A2(n47527), .ZN(n47545) );
  NAND2_X1 U48912 ( .A1(n47534), .A2(n47545), .ZN(n47522) );
  NAND3_X1 U48913 ( .A1(n47524), .A2(n47523), .A3(n47522), .ZN(n47537) );
  NAND3_X1 U48914 ( .A1(n47526), .A2(n47533), .A3(n47525), .ZN(n47536) );
  INV_X1 U48915 ( .A(n47527), .ZN(n47575) );
  OAI211_X1 U48919 ( .C1(n47534), .C2(n47575), .A(n47533), .B(n47532), .ZN(
        n47535) );
  NAND2_X1 U48920 ( .A1(n47538), .A2(n52045), .ZN(n47540) );
  OAI211_X1 U48921 ( .C1(n47542), .C2(n47541), .A(n47540), .B(n47539), .ZN(
        n47544) );
  NAND2_X1 U48922 ( .A1(n47544), .A2(n47543), .ZN(n47551) );
  NAND4_X1 U48923 ( .A1(n47551), .A2(n47550), .A3(n47549), .A4(n47548), .ZN(
        n47553) );
  INV_X1 U48924 ( .A(n4237), .ZN(n47552) );
  XNOR2_X1 U48925 ( .A(n47553), .B(n47552), .ZN(Plaintext[4]) );
  NAND2_X1 U48926 ( .A1(n47573), .A2(n51289), .ZN(n47555) );
  NOR2_X1 U48927 ( .A1(n47556), .A2(n47555), .ZN(n47561) );
  INV_X1 U48928 ( .A(n51290), .ZN(n47560) );
  NOR2_X1 U48929 ( .A1(n47558), .A2(n52044), .ZN(n47559) );
  AOI22_X1 U48930 ( .A1(n51346), .A2(n47561), .B1(n47560), .B2(n47559), .ZN(
        n47583) );
  OAI21_X1 U48931 ( .B1(n47579), .B2(n47573), .A(n52044), .ZN(n47564) );
  NAND2_X1 U48932 ( .A1(n47574), .A2(n47570), .ZN(n47565) );
  NAND3_X1 U48933 ( .A1(n47564), .A2(n47575), .A3(n47565), .ZN(n47568) );
  INV_X1 U48934 ( .A(n47565), .ZN(n47566) );
  NAND3_X1 U48935 ( .A1(n47566), .A2(n47573), .A3(n47579), .ZN(n47567) );
  OAI21_X1 U48936 ( .B1(n47573), .B2(n47574), .A(n47572), .ZN(n47569) );
  NAND3_X1 U48937 ( .A1(n47569), .A2(n47570), .A3(n47579), .ZN(n47578) );
  NAND3_X1 U48938 ( .A1(n47572), .A2(n47571), .A3(n47570), .ZN(n47577) );
  NAND3_X1 U48939 ( .A1(n47575), .A2(n47574), .A3(n47573), .ZN(n47576) );
  AND3_X1 U48940 ( .A1(n47578), .A2(n47577), .A3(n47576), .ZN(n47582) );
  NAND2_X1 U48941 ( .A1(n47580), .A2(n47579), .ZN(n47581) );
  INV_X1 U48942 ( .A(n4535), .ZN(n47584) );
  NOR2_X1 U48943 ( .A1(n46668), .A2(n47586), .ZN(n47607) );
  AOI21_X1 U48944 ( .B1(n47588), .B2(n47587), .A(n47607), .ZN(n47594) );
  OAI21_X1 U48945 ( .B1(n47619), .B2(n47591), .A(n47590), .ZN(n47593) );
  XNOR2_X1 U48946 ( .A(n51401), .B(n2163), .ZN(n47598) );
  OAI211_X1 U48947 ( .C1(n2163), .C2(n47617), .A(n47598), .B(n51340), .ZN(
        n47600) );
  NOR2_X1 U48948 ( .A1(n47603), .A2(n47602), .ZN(n47604) );
  XNOR2_X1 U48949 ( .A(n47604), .B(n4312), .ZN(Plaintext[9]) );
  AND2_X1 U48950 ( .A1(n47606), .A2(n47605), .ZN(n47626) );
  NAND2_X1 U48951 ( .A1(n47608), .A2(n47607), .ZN(n47609) );
  OAI211_X1 U48952 ( .C1(n46668), .C2(n47619), .A(n47610), .B(n47609), .ZN(
        n47612) );
  INV_X1 U48953 ( .A(n47612), .ZN(n47625) );
  AOI21_X1 U48954 ( .B1(n47619), .B2(n47618), .A(n47617), .ZN(n47621) );
  OAI21_X1 U48955 ( .B1(n47622), .B2(n47621), .A(n1187), .ZN(n47623) );
  NAND2_X1 U48956 ( .A1(n47675), .A2(n47689), .ZN(n47628) );
  OR2_X1 U48957 ( .A1(n47629), .A2(n47628), .ZN(n47644) );
  OR2_X1 U48958 ( .A1(n47655), .A2(n47686), .ZN(n47700) );
  AND2_X1 U48959 ( .A1(n47689), .A2(n47688), .ZN(n47630) );
  OAI21_X1 U48960 ( .B1(n47700), .B2(n47630), .A(n47702), .ZN(n47633) );
  OAI21_X1 U48961 ( .B1(n47656), .B2(n47687), .A(n47699), .ZN(n47632) );
  NAND4_X1 U48962 ( .A1(n47685), .A2(n47688), .A3(n47651), .A4(n47686), .ZN(
        n47631) );
  NAND4_X1 U48963 ( .A1(n47644), .A2(n47633), .A3(n47632), .A4(n47631), .ZN(
        n47639) );
  AOI21_X1 U48964 ( .B1(n47665), .B2(n47655), .A(n47694), .ZN(n47637) );
  NOR2_X1 U48965 ( .A1(n47650), .A2(n47687), .ZN(n47634) );
  NAND4_X1 U48966 ( .A1(n47673), .A2(n47675), .A3(n47634), .A4(n47689), .ZN(
        n47636) );
  NAND3_X1 U48967 ( .A1(n47656), .A2(n47698), .A3(n47674), .ZN(n47635) );
  OAI211_X1 U48968 ( .C1(n47637), .C2(n47688), .A(n47636), .B(n47635), .ZN(
        n47638) );
  INV_X1 U48970 ( .A(n4578), .ZN(n47640) );
  XNOR2_X1 U48971 ( .A(n47641), .B(n47640), .ZN(Plaintext[12]) );
  NAND3_X1 U48972 ( .A1(n47642), .A2(n47694), .A3(n47688), .ZN(n47643) );
  AND3_X1 U48973 ( .A1(n47645), .A2(n47644), .A3(n47643), .ZN(n47661) );
  AND2_X1 U48974 ( .A1(n47688), .A2(n47655), .ZN(n47695) );
  NAND3_X1 U48975 ( .A1(n47667), .A2(n47695), .A3(n47665), .ZN(n47649) );
  NAND2_X1 U48976 ( .A1(n47688), .A2(n47686), .ZN(n47646) );
  NAND2_X1 U48977 ( .A1(n47646), .A2(n47651), .ZN(n47647) );
  NAND2_X1 U48978 ( .A1(n47685), .A2(n47647), .ZN(n47648) );
  AND2_X1 U48979 ( .A1(n47649), .A2(n47648), .ZN(n47660) );
  AND2_X1 U48980 ( .A1(n47675), .A2(n47687), .ZN(n47671) );
  OR2_X1 U48981 ( .A1(n47689), .A2(n47650), .ZN(n47669) );
  NAND2_X1 U48982 ( .A1(n47665), .A2(n47698), .ZN(n47653) );
  OAI21_X1 U48983 ( .B1(n47651), .B2(n47686), .A(n47688), .ZN(n47652) );
  NOR3_X1 U48984 ( .A1(n47655), .A2(n47688), .A3(n47687), .ZN(n47657) );
  AOI22_X1 U48985 ( .A1(n47683), .A2(n47691), .B1(n47657), .B2(n47656), .ZN(
        n47658) );
  NAND4_X1 U48986 ( .A1(n47661), .A2(n47660), .A3(n47659), .A4(n47658), .ZN(
        n47663) );
  INV_X1 U48987 ( .A(n4908), .ZN(n47662) );
  XNOR2_X1 U48988 ( .A(n47663), .B(n47662), .ZN(Plaintext[13]) );
  INV_X1 U48989 ( .A(n47691), .ZN(n47666) );
  INV_X1 U48990 ( .A(n47668), .ZN(n47672) );
  INV_X1 U48991 ( .A(n47669), .ZN(n47670) );
  OAI211_X1 U48992 ( .C1(n47674), .C2(n47694), .A(n47684), .B(n47673), .ZN(
        n47677) );
  OR2_X1 U48993 ( .A1(n47689), .A2(n47675), .ZN(n47681) );
  INV_X1 U48994 ( .A(n47681), .ZN(n47676) );
  INV_X1 U48995 ( .A(n47679), .ZN(n47680) );
  NAND2_X1 U48996 ( .A1(n47681), .A2(n47686), .ZN(n47682) );
  OAI211_X1 U48997 ( .C1(n47684), .C2(n47691), .A(n47683), .B(n47682), .ZN(
        n47707) );
  OAI211_X1 U48998 ( .C1(n47698), .C2(n47686), .A(n47685), .B(n47687), .ZN(
        n47693) );
  AND2_X1 U48999 ( .A1(n47688), .A2(n47687), .ZN(n47690) );
  OAI21_X1 U49000 ( .B1(n47691), .B2(n47690), .A(n47689), .ZN(n47692) );
  AND2_X1 U49001 ( .A1(n47693), .A2(n47692), .ZN(n47706) );
  NAND2_X1 U49002 ( .A1(n47695), .A2(n47694), .ZN(n47696) );
  AND2_X1 U49003 ( .A1(n47697), .A2(n47696), .ZN(n47705) );
  NAND2_X1 U49005 ( .A1(n47701), .A2(n47700), .ZN(n47703) );
  NAND2_X1 U49006 ( .A1(n47703), .A2(n47702), .ZN(n47704) );
  INV_X1 U49010 ( .A(n47710), .ZN(n47715) );
  NAND3_X1 U49011 ( .A1(n47712), .A2(n47797), .A3(n47711), .ZN(n47714) );
  AND2_X1 U49012 ( .A1(n47745), .A2(n47721), .ZN(n47789) );
  INV_X1 U49013 ( .A(n47779), .ZN(n47713) );
  INV_X1 U49014 ( .A(n47716), .ZN(n47718) );
  NAND2_X1 U49015 ( .A1(n47790), .A2(n51468), .ZN(n47764) );
  NOR2_X1 U49016 ( .A1(n47745), .A2(n47721), .ZN(n47717) );
  OAI22_X1 U49017 ( .A1(n47718), .A2(n47780), .B1(n47764), .B2(n47717), .ZN(
        n47720) );
  AOI21_X1 U49018 ( .B1(n47781), .B2(n47797), .A(n47752), .ZN(n47719) );
  NOR2_X1 U49019 ( .A1(n47720), .A2(n47719), .ZN(n47724) );
  NAND2_X1 U49020 ( .A1(n45877), .A2(n47745), .ZN(n47731) );
  NOR2_X1 U49021 ( .A1(n47731), .A2(n47777), .ZN(n47788) );
  NAND2_X1 U49022 ( .A1(n47788), .A2(n47721), .ZN(n47723) );
  INV_X1 U49025 ( .A(n4542), .ZN(n47725) );
  OR2_X1 U49027 ( .A1(n47792), .A2(n45877), .ZN(n47796) );
  OAI21_X1 U49028 ( .B1(n47755), .B2(n47752), .A(n47796), .ZN(n47727) );
  NAND2_X1 U49029 ( .A1(n47727), .A2(n47762), .ZN(n47736) );
  OAI21_X1 U49030 ( .B1(n47752), .B2(n47745), .A(n52118), .ZN(n47729) );
  AND2_X1 U49031 ( .A1(n47728), .A2(n51468), .ZN(n47791) );
  OAI21_X1 U49032 ( .B1(n47729), .B2(n47791), .A(n52149), .ZN(n47735) );
  NAND2_X1 U49033 ( .A1(n47730), .A2(n47791), .ZN(n47734) );
  NAND2_X1 U49034 ( .A1(n645), .A2(n47731), .ZN(n47732) );
  NAND4_X1 U49035 ( .A1(n47736), .A2(n47735), .A3(n47734), .A4(n47733), .ZN(
        n47739) );
  INV_X1 U49036 ( .A(n47737), .ZN(n47738) );
  XNOR2_X1 U49037 ( .A(n47739), .B(n47738), .ZN(Plaintext[20]) );
  MUX2_X1 U49038 ( .A(n47786), .B(n47740), .S(n47763), .Z(n47772) );
  INV_X1 U49039 ( .A(n47772), .ZN(n47750) );
  NAND2_X1 U49040 ( .A1(n47743), .A2(n45877), .ZN(n47741) );
  INV_X1 U49042 ( .A(n47798), .ZN(n47749) );
  AND2_X1 U49043 ( .A1(n52149), .A2(n4628), .ZN(n47748) );
  NOR2_X1 U49044 ( .A1(n47744), .A2(n51468), .ZN(n47746) );
  OAI21_X1 U49045 ( .B1(n47747), .B2(n47746), .A(n47745), .ZN(n47757) );
  NAND4_X1 U49046 ( .A1(n47757), .A2(n47749), .A3(n47748), .A4(n47750), .ZN(
        n47776) );
  NAND2_X1 U49047 ( .A1(n47771), .A2(n52118), .ZN(n47751) );
  OAI211_X1 U49048 ( .C1(n645), .C2(n47752), .A(n4628), .B(n47751), .ZN(n47753) );
  NOR2_X1 U49049 ( .A1(n47753), .A2(n47798), .ZN(n47759) );
  INV_X1 U49050 ( .A(n47754), .ZN(n47758) );
  NAND4_X1 U49051 ( .A1(n47759), .A2(n47758), .A3(n47757), .A4(n47756), .ZN(
        n47775) );
  AOI22_X1 U49052 ( .A1(n47762), .A2(n47761), .B1(n47760), .B2(n47797), .ZN(
        n47769) );
  AOI21_X1 U49053 ( .B1(n52118), .B2(n47763), .A(n4628), .ZN(n47765) );
  OAI211_X1 U49054 ( .C1(n47766), .C2(n47786), .A(n47765), .B(n47764), .ZN(
        n47767) );
  INV_X1 U49055 ( .A(n47767), .ZN(n47768) );
  OAI21_X1 U49056 ( .B1(n47769), .B2(n45877), .A(n47768), .ZN(n47774) );
  INV_X1 U49057 ( .A(n4628), .ZN(n47770) );
  NAND4_X1 U49058 ( .A1(n47772), .A2(n52149), .A3(n52118), .A4(n47770), .ZN(
        n47773) );
  NAND4_X1 U49059 ( .A1(n47776), .A2(n47775), .A3(n47774), .A4(n47773), .ZN(
        Plaintext[22]) );
  NAND2_X1 U49060 ( .A1(n51468), .A2(n47777), .ZN(n47793) );
  NOR2_X1 U49061 ( .A1(n47784), .A2(n47783), .ZN(n47801) );
  OAI21_X1 U49062 ( .B1(n47788), .B2(n47787), .A(n47786), .ZN(n47800) );
  OAI21_X1 U49063 ( .B1(n651), .B2(n51285), .A(n47880), .ZN(n47840) );
  AOI21_X1 U49064 ( .B1(n47840), .B2(n51469), .A(n47803), .ZN(n47805) );
  NOR2_X1 U49065 ( .A1(n47875), .A2(n47841), .ZN(n47807) );
  NAND2_X1 U49066 ( .A1(n47842), .A2(n508), .ZN(n47827) );
  NAND2_X1 U49067 ( .A1(n47827), .A2(n51285), .ZN(n47806) );
  AOI22_X1 U49068 ( .A1(n47807), .A2(n47806), .B1(n47824), .B2(n47855), .ZN(
        n47811) );
  NAND2_X1 U49069 ( .A1(n47831), .A2(n47841), .ZN(n47839) );
  NOR2_X1 U49070 ( .A1(n47839), .A2(n3798), .ZN(n47886) );
  NAND2_X1 U49071 ( .A1(n51469), .A2(n47841), .ZN(n47828) );
  AOI22_X1 U49072 ( .A1(n47842), .A2(n47828), .B1(n47883), .B2(n508), .ZN(
        n47809) );
  OAI21_X1 U49073 ( .B1(n47883), .B2(n508), .A(n47880), .ZN(n47808) );
  AOI22_X1 U49074 ( .A1(n47886), .A2(n47885), .B1(n47809), .B2(n47808), .ZN(
        n47810) );
  INV_X1 U49075 ( .A(n4659), .ZN(n47812) );
  XNOR2_X1 U49076 ( .A(n47813), .B(n47812), .ZN(Plaintext[24]) );
  NAND2_X1 U49077 ( .A1(n51285), .A2(n47857), .ZN(n47882) );
  NOR2_X1 U49079 ( .A1(n47882), .A2(n47814), .ZN(n47865) );
  NOR2_X1 U49082 ( .A1(n47865), .A2(n47816), .ZN(n47823) );
  INV_X1 U49083 ( .A(n51469), .ZN(n47881) );
  INV_X1 U49084 ( .A(n47839), .ZN(n47867) );
  NAND3_X1 U49085 ( .A1(n3386), .A2(n47881), .A3(n47867), .ZN(n47821) );
  XNOR2_X1 U49086 ( .A(n47883), .B(n51285), .ZN(n47819) );
  NOR3_X1 U49087 ( .A1(n508), .A2(n51470), .A3(n47873), .ZN(n47818) );
  NAND4_X1 U49089 ( .A1(n47823), .A2(n47822), .A3(n47821), .A4(n47820), .ZN(
        n47836) );
  AND2_X1 U49093 ( .A1(n508), .A2(n47831), .ZN(n47870) );
  NAND3_X1 U49094 ( .A1(n47870), .A2(n47881), .A3(n51285), .ZN(n47832) );
  OR2_X1 U49095 ( .A1(n47836), .A2(n47835), .ZN(n47838) );
  INV_X1 U49096 ( .A(n4836), .ZN(n47837) );
  XNOR2_X1 U49097 ( .A(n47838), .B(n47837), .ZN(Plaintext[25]) );
  AOI21_X1 U49098 ( .B1(n47839), .B2(n508), .A(n47881), .ZN(n47846) );
  OAI21_X1 U49099 ( .B1(n47866), .B2(n47855), .A(n47840), .ZN(n47845) );
  NAND2_X1 U49100 ( .A1(n47842), .A2(n47841), .ZN(n47851) );
  INV_X1 U49101 ( .A(n47851), .ZN(n47854) );
  NAND2_X1 U49102 ( .A1(n47882), .A2(n47875), .ZN(n47843) );
  AOI21_X1 U49103 ( .B1(n47854), .B2(n47843), .A(n47885), .ZN(n47844) );
  OAI211_X1 U49104 ( .C1(n47846), .C2(n47858), .A(n47845), .B(n47844), .ZN(
        n47848) );
  INV_X1 U49105 ( .A(n4353), .ZN(n47847) );
  XNOR2_X1 U49106 ( .A(n47848), .B(n47847), .ZN(Plaintext[26]) );
  OR2_X1 U49107 ( .A1(n47849), .A2(n651), .ZN(n47863) );
  INV_X1 U49108 ( .A(n47850), .ZN(n47852) );
  AOI21_X1 U49109 ( .B1(n47852), .B2(n47851), .A(n47855), .ZN(n47853) );
  OAI21_X1 U49110 ( .B1(n47866), .B2(n47854), .A(n47853), .ZN(n47862) );
  INV_X1 U49111 ( .A(n47865), .ZN(n47861) );
  INV_X1 U49112 ( .A(n47875), .ZN(n47859) );
  NAND2_X1 U49113 ( .A1(n47855), .A2(n47880), .ZN(n47856) );
  OAI211_X1 U49114 ( .C1(n47859), .C2(n47858), .A(n508), .B(n47856), .ZN(
        n47860) );
  INV_X1 U49115 ( .A(n4502), .ZN(n47864) );
  OAI211_X1 U49116 ( .C1(n47870), .C2(n51469), .A(n51285), .B(n47873), .ZN(
        n47871) );
  NAND2_X1 U49117 ( .A1(n47872), .A2(n47871), .ZN(n47878) );
  OAI22_X1 U49118 ( .A1(n47876), .A2(n47875), .B1(n47874), .B2(n47873), .ZN(
        n47877) );
  NOR2_X1 U49119 ( .A1(n47878), .A2(n47877), .ZN(n47889) );
  OAI22_X1 U49120 ( .A1(n47882), .A2(n47881), .B1(n47880), .B2(n47879), .ZN(
        n47884) );
  NAND2_X1 U49121 ( .A1(n47884), .A2(n47883), .ZN(n47888) );
  OAI21_X1 U49122 ( .B1(n47886), .B2(n3386), .A(n47885), .ZN(n47887) );
  INV_X1 U49123 ( .A(n4720), .ZN(n47890) );
  NOR2_X1 U49124 ( .A1(n47966), .A2(n47989), .ZN(n47957) );
  AOI21_X1 U49125 ( .B1(n47962), .B2(n47891), .A(n47989), .ZN(n47894) );
  NAND2_X1 U49126 ( .A1(n47892), .A2(n47962), .ZN(n47893) );
  NAND2_X1 U49127 ( .A1(n47894), .A2(n47893), .ZN(n47895) );
  OAI21_X1 U49128 ( .B1(n47957), .B2(n47936), .A(n47895), .ZN(n47897) );
  NAND2_X1 U49129 ( .A1(n47928), .A2(n47996), .ZN(n47896) );
  MUX2_X1 U49130 ( .A(n47897), .B(n47896), .S(n51805), .Z(n47923) );
  OAI21_X1 U49131 ( .B1(n47945), .B2(n47935), .A(n47980), .ZN(n47898) );
  NAND3_X1 U49133 ( .A1(n47899), .A2(n567), .A3(n47944), .ZN(n47902) );
  NAND2_X1 U49134 ( .A1(n47966), .A2(n52057), .ZN(n47900) );
  AND3_X1 U49135 ( .A1(n47903), .A2(n47902), .A3(n47901), .ZN(n47922) );
  NAND2_X1 U49137 ( .A1(n51805), .A2(n47936), .ZN(n47984) );
  NOR2_X1 U49138 ( .A1(n47984), .A2(n47989), .ZN(n47906) );
  NOR2_X1 U49139 ( .A1(n47991), .A2(n47965), .ZN(n47905) );
  AOI22_X1 U49142 ( .A1(n47960), .A2(n47906), .B1(n47905), .B2(n47961), .ZN(
        n47921) );
  NAND2_X1 U49143 ( .A1(n47908), .A2(n47907), .ZN(n47910) );
  NAND2_X1 U49144 ( .A1(n47910), .A2(n47909), .ZN(n47916) );
  AND2_X1 U49145 ( .A1(n47912), .A2(n47911), .ZN(n47915) );
  NAND4_X1 U49146 ( .A1(n47916), .A2(n47915), .A3(n47914), .A4(n47913), .ZN(
        n47917) );
  NAND4_X1 U49147 ( .A1(n47991), .A2(n47988), .A3(n47936), .A4(n47917), .ZN(
        n47918) );
  NAND2_X1 U49148 ( .A1(n47918), .A2(n47941), .ZN(n47919) );
  NAND2_X1 U49149 ( .A1(n47919), .A2(n47990), .ZN(n47920) );
  INV_X1 U49150 ( .A(n2203), .ZN(n47924) );
  NOR2_X1 U49151 ( .A1(n47925), .A2(n51805), .ZN(n47949) );
  OAI21_X1 U49152 ( .B1(n47949), .B2(n47990), .A(n47989), .ZN(n47934) );
  OAI21_X1 U49153 ( .B1(n648), .B2(n47986), .A(n51805), .ZN(n47931) );
  NAND2_X1 U49154 ( .A1(n47935), .A2(n47966), .ZN(n47973) );
  OAI21_X1 U49155 ( .B1(n648), .B2(n47973), .A(n47986), .ZN(n47930) );
  NAND2_X1 U49156 ( .A1(n47931), .A2(n47930), .ZN(n47932) );
  AND2_X1 U49157 ( .A1(n47935), .A2(n52057), .ZN(n47940) );
  XNOR2_X1 U49158 ( .A(n47937), .B(n47936), .ZN(n47938) );
  OAI211_X1 U49160 ( .C1(n47990), .C2(n47941), .A(n47940), .B(n47939), .ZN(
        n47942) );
  NOR2_X1 U49162 ( .A1(n47945), .A2(n47944), .ZN(n47946) );
  AOI21_X1 U49163 ( .B1(n47979), .B2(n47946), .A(n52057), .ZN(n47953) );
  NAND2_X1 U49164 ( .A1(n47990), .A2(n47988), .ZN(n47947) );
  NAND2_X1 U49165 ( .A1(n47947), .A2(n47962), .ZN(n47948) );
  NAND2_X1 U49166 ( .A1(n47949), .A2(n47948), .ZN(n47952) );
  NOR2_X1 U49167 ( .A1(n47950), .A2(n47990), .ZN(n47976) );
  NAND2_X1 U49168 ( .A1(n47996), .A2(n47976), .ZN(n47951) );
  INV_X1 U49170 ( .A(n4896), .ZN(n47955) );
  XNOR2_X1 U49171 ( .A(n47956), .B(n47955), .ZN(Plaintext[33]) );
  AND2_X1 U49172 ( .A1(n47957), .A2(n47974), .ZN(n47959) );
  INV_X1 U49173 ( .A(n47980), .ZN(n47958) );
  AOI22_X1 U49174 ( .A1(n47960), .A2(n47959), .B1(n648), .B2(n47958), .ZN(
        n47970) );
  NAND2_X1 U49175 ( .A1(n47979), .A2(n47961), .ZN(n47964) );
  INV_X1 U49176 ( .A(n47981), .ZN(n47963) );
  NAND2_X1 U49177 ( .A1(n47964), .A2(n47963), .ZN(n47969) );
  OR2_X1 U49178 ( .A1(n47965), .A2(n47988), .ZN(n47968) );
  AND2_X1 U49179 ( .A1(n47990), .A2(n47966), .ZN(n47985) );
  OAI211_X1 U49180 ( .C1(n47988), .C2(n52056), .A(n648), .B(n47985), .ZN(
        n47967) );
  NAND4_X1 U49181 ( .A1(n47970), .A2(n47969), .A3(n47968), .A4(n47967), .ZN(
        n47972) );
  INV_X1 U49182 ( .A(n4317), .ZN(n47971) );
  XNOR2_X1 U49183 ( .A(n47972), .B(n47971), .ZN(Plaintext[34]) );
  INV_X1 U49184 ( .A(n47973), .ZN(n47975) );
  NAND3_X1 U49185 ( .A1(n47975), .A2(n567), .A3(n47974), .ZN(n47978) );
  INV_X1 U49186 ( .A(n47976), .ZN(n47977) );
  INV_X1 U49187 ( .A(n47979), .ZN(n47983) );
  NAND2_X1 U49188 ( .A1(n47981), .A2(n47980), .ZN(n47982) );
  OAI211_X1 U49189 ( .C1(n47985), .C2(n47984), .A(n47983), .B(n47982), .ZN(
        n47998) );
  OAI21_X1 U49190 ( .B1(n47988), .B2(n47987), .A(n47986), .ZN(n47994) );
  AND3_X1 U49191 ( .A1(n47990), .A2(n47989), .A3(n52057), .ZN(n47992) );
  NAND2_X1 U49192 ( .A1(n47996), .A2(n47995), .ZN(n47997) );
  INV_X1 U49193 ( .A(n4837), .ZN(n48000) );
  XNOR2_X1 U49194 ( .A(n48001), .B(n48000), .ZN(Plaintext[35]) );
  INV_X1 U49195 ( .A(n48002), .ZN(n48003) );
  NAND3_X1 U49196 ( .A1(n48005), .A2(n48004), .A3(n48068), .ZN(n48006) );
  NAND2_X1 U49197 ( .A1(n48006), .A2(n650), .ZN(n48017) );
  NAND2_X1 U49198 ( .A1(n48007), .A2(n48051), .ZN(n48008) );
  NAND2_X1 U49199 ( .A1(n48008), .A2(n48084), .ZN(n48012) );
  NAND2_X1 U49200 ( .A1(n51343), .A2(n48077), .ZN(n48010) );
  AOI21_X1 U49201 ( .B1(n48074), .B2(n48010), .A(n48009), .ZN(n48011) );
  NAND2_X1 U49202 ( .A1(n48012), .A2(n48011), .ZN(n48016) );
  OR2_X1 U49203 ( .A1(n48084), .A2(n48083), .ZN(n48070) );
  INV_X1 U49204 ( .A(n48070), .ZN(n48014) );
  XNOR2_X1 U49205 ( .A(n48051), .B(n51343), .ZN(n48013) );
  NAND2_X1 U49206 ( .A1(n48014), .A2(n48013), .ZN(n48015) );
  INV_X1 U49207 ( .A(n4454), .ZN(n48018) );
  AND2_X1 U49208 ( .A1(n48039), .A2(n48019), .ZN(n48076) );
  AOI21_X1 U49209 ( .B1(n48072), .B2(n48067), .A(n48076), .ZN(n48027) );
  AND2_X1 U49210 ( .A1(n48051), .A2(n48074), .ZN(n48078) );
  OAI21_X1 U49211 ( .B1(n6355), .B2(n48078), .A(n48020), .ZN(n48026) );
  INV_X1 U49212 ( .A(n48021), .ZN(n48022) );
  NAND3_X1 U49213 ( .A1(n48022), .A2(n48059), .A3(n51343), .ZN(n48025) );
  NOR3_X1 U49214 ( .A1(n48084), .A2(n48051), .A3(n48077), .ZN(n48023) );
  OAI21_X1 U49215 ( .B1(n48023), .B2(n52127), .A(n48074), .ZN(n48024) );
  NAND4_X1 U49216 ( .A1(n48027), .A2(n48026), .A3(n48025), .A4(n48024), .ZN(
        n48029) );
  INV_X1 U49217 ( .A(n3336), .ZN(n48028) );
  XNOR2_X1 U49218 ( .A(n48029), .B(n48028), .ZN(Plaintext[38]) );
  NOR2_X1 U49219 ( .A1(n48082), .A2(n48084), .ZN(n48075) );
  NOR2_X1 U49220 ( .A1(n48039), .A2(n48085), .ZN(n48031) );
  INV_X1 U49221 ( .A(n48069), .ZN(n48030) );
  OAI22_X1 U49222 ( .A1(n48075), .A2(n48031), .B1(n48030), .B2(n52127), .ZN(
        n48048) );
  NAND3_X1 U49223 ( .A1(n48032), .A2(n52127), .A3(n48084), .ZN(n48035) );
  NAND2_X1 U49224 ( .A1(n48051), .A2(n51343), .ZN(n48034) );
  OAI22_X1 U49225 ( .A1(n48035), .A2(n48078), .B1(n48084), .B2(n48034), .ZN(
        n48036) );
  INV_X1 U49226 ( .A(n48036), .ZN(n48047) );
  INV_X1 U49227 ( .A(n48059), .ZN(n48056) );
  OAI21_X1 U49228 ( .B1(n52127), .B2(n48074), .A(n48082), .ZN(n48037) );
  INV_X1 U49229 ( .A(n48037), .ZN(n48040) );
  NAND4_X1 U49230 ( .A1(n48056), .A2(n48040), .A3(n48039), .A4(n48038), .ZN(
        n48046) );
  INV_X1 U49231 ( .A(n48042), .ZN(n48043) );
  NAND3_X1 U49232 ( .A1(n48044), .A2(n48043), .A3(n650), .ZN(n48045) );
  NAND4_X1 U49233 ( .A1(n48048), .A2(n48047), .A3(n48046), .A4(n48045), .ZN(
        n48050) );
  INV_X1 U49234 ( .A(n4937), .ZN(n48049) );
  XNOR2_X1 U49235 ( .A(n48050), .B(n48049), .ZN(Plaintext[39]) );
  NAND3_X1 U49236 ( .A1(n48053), .A2(n48081), .A3(n48051), .ZN(n48052) );
  NAND3_X1 U49237 ( .A1(n48076), .A2(n51092), .A3(n48066), .ZN(n48062) );
  NAND2_X1 U49238 ( .A1(n48054), .A2(n48053), .ZN(n48055) );
  NAND2_X1 U49239 ( .A1(n48056), .A2(n48055), .ZN(n48061) );
  NAND2_X1 U49240 ( .A1(n48084), .A2(n51092), .ZN(n48058) );
  NAND2_X1 U49241 ( .A1(n48059), .A2(n48058), .ZN(n48079) );
  NAND2_X1 U49242 ( .A1(n48079), .A2(n48078), .ZN(n48060) );
  NAND4_X1 U49243 ( .A1(n48063), .A2(n48062), .A3(n48061), .A4(n48060), .ZN(
        n48065) );
  XNOR2_X1 U49244 ( .A(n48065), .B(n48064), .ZN(Plaintext[40]) );
  AND2_X1 U49245 ( .A1(n48067), .A2(n48066), .ZN(n48073) );
  AOI21_X1 U49246 ( .B1(n48073), .B2(n48072), .A(n48071), .ZN(n48090) );
  OAI21_X1 U49247 ( .B1(n48076), .B2(n48075), .A(n48074), .ZN(n48089) );
  NAND2_X1 U49248 ( .A1(n48084), .A2(n48077), .ZN(n48080) );
  OAI211_X1 U49249 ( .C1(n48081), .C2(n48080), .A(n48079), .B(n48078), .ZN(
        n48088) );
  MUX2_X1 U49250 ( .A(n48086), .B(n48085), .S(n48084), .Z(n48087) );
  INV_X1 U49251 ( .A(n4537), .ZN(n48091) );
  INV_X1 U49252 ( .A(n48095), .ZN(n48099) );
  INV_X1 U49253 ( .A(n48127), .ZN(n48098) );
  NAND2_X1 U49254 ( .A1(n48160), .A2(n48155), .ZN(n48096) );
  AOI22_X1 U49255 ( .A1(n48099), .A2(n48098), .B1(n48097), .B2(n48096), .ZN(
        n48107) );
  NAND2_X1 U49256 ( .A1(n48152), .A2(n48112), .ZN(n48106) );
  INV_X1 U49257 ( .A(n48158), .ZN(n48104) );
  NAND2_X1 U49258 ( .A1(n48157), .A2(n3911), .ZN(n48101) );
  NAND2_X1 U49259 ( .A1(n48101), .A2(n48100), .ZN(n48134) );
  NAND4_X1 U49260 ( .A1(n48104), .A2(n48103), .A3(n48134), .A4(n48102), .ZN(
        n48105) );
  INV_X1 U49261 ( .A(n274), .ZN(n48108) );
  AOI21_X1 U49262 ( .B1(n48141), .B2(n48115), .A(n48135), .ZN(n48121) );
  AND2_X1 U49263 ( .A1(n48110), .A2(n8689), .ZN(n48111) );
  OAI21_X1 U49264 ( .B1(n48152), .B2(n48111), .A(n48117), .ZN(n48120) );
  NAND2_X1 U49265 ( .A1(n48155), .A2(n48156), .ZN(n48113) );
  OAI22_X1 U49266 ( .A1(n48160), .A2(n48113), .B1(n48116), .B2(n48112), .ZN(
        n48114) );
  INV_X1 U49267 ( .A(n48114), .ZN(n48119) );
  NAND4_X1 U49268 ( .A1(n48121), .A2(n48120), .A3(n48119), .A4(n48118), .ZN(
        n48123) );
  XNOR2_X1 U49269 ( .A(n48123), .B(n48122), .ZN(Plaintext[44]) );
  MUX2_X1 U49270 ( .A(n48127), .B(n48126), .S(n48159), .Z(n48150) );
  INV_X1 U49271 ( .A(n48128), .ZN(n48133) );
  NOR2_X1 U49272 ( .A1(n48157), .A2(n3911), .ZN(n48129) );
  OAI211_X1 U49273 ( .C1(n48157), .C2(n48140), .A(n48136), .B(n48156), .ZN(
        n48131) );
  OAI21_X1 U49274 ( .B1(n48131), .B2(n48130), .A(n4501), .ZN(n48132) );
  AOI21_X1 U49275 ( .B1(n48133), .B2(n48139), .A(n48132), .ZN(n48138) );
  NAND2_X1 U49276 ( .A1(n48134), .A2(n48152), .ZN(n48144) );
  OAI21_X1 U49277 ( .B1(n48135), .B2(n48151), .A(n8306), .ZN(n48145) );
  OR2_X1 U49278 ( .A1(n48145), .A2(n48136), .ZN(n48137) );
  NAND4_X1 U49279 ( .A1(n48150), .A2(n48138), .A3(n48144), .A4(n48137), .ZN(
        n48149) );
  AOI21_X1 U49280 ( .B1(n48156), .B2(n48140), .A(n48155), .ZN(n48143) );
  INV_X1 U49281 ( .A(n48141), .ZN(n48142) );
  INV_X1 U49282 ( .A(n48144), .ZN(n48147) );
  AOI21_X1 U49283 ( .B1(n48145), .B2(n48155), .A(n4501), .ZN(n48146) );
  OAI21_X1 U49284 ( .B1(n48155), .B2(n48154), .A(n48153), .ZN(n48163) );
  INV_X1 U49285 ( .A(n4048), .ZN(n48164) );
  NAND2_X1 U49286 ( .A1(n48165), .A2(n2742), .ZN(n48177) );
  NAND2_X1 U49287 ( .A1(n48166), .A2(n48174), .ZN(n48167) );
  INV_X1 U49288 ( .A(n48169), .ZN(n48170) );
  INV_X1 U49289 ( .A(n48412), .ZN(n48173) );
  INV_X1 U49290 ( .A(n48402), .ZN(n48172) );
  AOI22_X1 U49291 ( .A1(n48173), .A2(n48414), .B1(n48172), .B2(n48171), .ZN(
        n48176) );
  INV_X1 U49292 ( .A(n48174), .ZN(n48175) );
  INV_X1 U49293 ( .A(n48177), .ZN(n48178) );
  INV_X1 U49294 ( .A(n48405), .ZN(n48409) );
  NAND3_X1 U49295 ( .A1(n48414), .A2(n48180), .A3(n48179), .ZN(n48181) );
  NAND3_X1 U49296 ( .A1(n48183), .A2(n48182), .A3(n48181), .ZN(n48184) );
  NOR2_X1 U49297 ( .A1(n48185), .A2(n48184), .ZN(n48186) );
  INV_X1 U49298 ( .A(n48510), .ZN(n48191) );
  INV_X1 U49299 ( .A(n48188), .ZN(n48190) );
  OAI211_X1 U49300 ( .C1(n51451), .C2(n48191), .A(n48190), .B(n48189), .ZN(
        n48194) );
  INV_X1 U49301 ( .A(n48192), .ZN(n48193) );
  NAND2_X1 U49302 ( .A1(n48194), .A2(n48193), .ZN(n48199) );
  XNOR2_X1 U49303 ( .A(n48505), .B(n48517), .ZN(n48195) );
  NAND2_X1 U49304 ( .A1(n48195), .A2(n45562), .ZN(n48197) );
  INV_X1 U49305 ( .A(n48196), .ZN(n48501) );
  AOI22_X1 U49306 ( .A1(n48197), .A2(n48501), .B1(n48522), .B2(n52202), .ZN(
        n48198) );
  INV_X1 U49307 ( .A(n48381), .ZN(n48392) );
  INV_X1 U49308 ( .A(n48369), .ZN(n48276) );
  NAND3_X1 U49309 ( .A1(n52050), .A2(n52070), .A3(n48200), .ZN(n48203) );
  MUX2_X1 U49310 ( .A(n48210), .B(n48209), .S(n48208), .Z(n48226) );
  AND2_X1 U49311 ( .A1(n48212), .A2(n48211), .ZN(n48225) );
  NAND2_X1 U49312 ( .A1(n48214), .A2(n48213), .ZN(n48215) );
  NAND2_X1 U49313 ( .A1(n48215), .A2(n48218), .ZN(n48217) );
  NAND2_X1 U49314 ( .A1(n48217), .A2(n48216), .ZN(n48224) );
  INV_X1 U49315 ( .A(n48218), .ZN(n48222) );
  OAI211_X1 U49316 ( .C1(n48222), .C2(n48221), .A(n48220), .B(n48219), .ZN(
        n48223) );
  OAI21_X1 U49317 ( .B1(n48227), .B2(n48524), .A(n48546), .ZN(n48228) );
  OAI211_X1 U49318 ( .C1(n48534), .C2(n48229), .A(n48550), .B(n48228), .ZN(
        n48231) );
  NAND2_X1 U49319 ( .A1(n48232), .A2(n48547), .ZN(n48243) );
  NAND3_X1 U49321 ( .A1(n48236), .A2(n52060), .A3(n48234), .ZN(n48241) );
  AND2_X1 U49322 ( .A1(n48238), .A2(n48237), .ZN(n48530) );
  OAI21_X1 U49323 ( .B1(n48239), .B2(n48540), .A(n48530), .ZN(n48240) );
  AND2_X1 U49325 ( .A1(n48247), .A2(n44409), .ZN(n48492) );
  NAND3_X1 U49326 ( .A1(n48492), .A2(n48246), .A3(n51301), .ZN(n48250) );
  AND2_X1 U49327 ( .A1(n48250), .A2(n48249), .ZN(n48310) );
  NAND4_X1 U49328 ( .A1(n48311), .A2(n48310), .A3(n48478), .A4(n48309), .ZN(
        n48257) );
  OAI211_X1 U49329 ( .C1(n48253), .C2(n48488), .A(n48252), .B(n48251), .ZN(
        n48314) );
  NAND2_X1 U49330 ( .A1(n48314), .A2(n48482), .ZN(n48256) );
  AND2_X1 U49331 ( .A1(n48480), .A2(n48479), .ZN(n48255) );
  OR2_X1 U49332 ( .A1(n48255), .A2(n48254), .ZN(n48308) );
  NOR2_X1 U49333 ( .A1(n48341), .A2(n52172), .ZN(n48361) );
  OAI21_X1 U49334 ( .B1(n48259), .B2(n48430), .A(n48269), .ZN(n48258) );
  INV_X1 U49336 ( .A(n48261), .ZN(n48262) );
  AOI21_X1 U49337 ( .B1(n48263), .B2(n48436), .A(n48262), .ZN(n48265) );
  NAND2_X1 U49338 ( .A1(n48267), .A2(n48436), .ZN(n48271) );
  OAI211_X1 U49339 ( .C1(n48269), .C2(n660), .A(n48268), .B(n48433), .ZN(
        n48270) );
  NAND3_X1 U49340 ( .A1(n48271), .A2(n48270), .A3(n48424), .ZN(n48272) );
  OAI21_X1 U49341 ( .B1(n48274), .B2(n48273), .A(n48272), .ZN(n48275) );
  OAI211_X1 U49342 ( .C1(n48276), .C2(n48361), .A(n48353), .B(n4035), .ZN(
        n48280) );
  OAI21_X1 U49343 ( .B1(n48369), .B2(n51072), .A(n6986), .ZN(n48278) );
  NOR2_X1 U49344 ( .A1(n52172), .A2(n51072), .ZN(n48340) );
  INV_X1 U49345 ( .A(n48340), .ZN(n48277) );
  AND2_X1 U49346 ( .A1(n51318), .A2(n51072), .ZN(n48359) );
  INV_X1 U49347 ( .A(n48359), .ZN(n48328) );
  NAND3_X1 U49348 ( .A1(n51356), .A2(n48277), .A3(n48328), .ZN(n48290) );
  NAND4_X1 U49349 ( .A1(n48278), .A2(n48290), .A3(n4035), .A4(n48380), .ZN(
        n48279) );
  NAND2_X1 U49350 ( .A1(n48280), .A2(n48279), .ZN(n48283) );
  AND2_X1 U49351 ( .A1(n51728), .A2(n48353), .ZN(n48329) );
  AND2_X1 U49352 ( .A1(n48381), .A2(n51072), .ZN(n48345) );
  INV_X1 U49353 ( .A(n48345), .ZN(n48306) );
  OAI22_X1 U49354 ( .A1(n48329), .A2(n48306), .B1(n48395), .B2(n48332), .ZN(
        n48286) );
  NAND3_X1 U49355 ( .A1(n51087), .A2(n48353), .A3(n48359), .ZN(n48304) );
  OAI21_X1 U49356 ( .B1(n48360), .B2(n48281), .A(n48304), .ZN(n48285) );
  NOR2_X1 U49357 ( .A1(n48286), .A2(n48285), .ZN(n48282) );
  NAND2_X1 U49358 ( .A1(n48283), .A2(n48282), .ZN(n48295) );
  INV_X1 U49359 ( .A(n4035), .ZN(n48284) );
  OAI21_X1 U49360 ( .B1(n48286), .B2(n48285), .A(n48284), .ZN(n48294) );
  INV_X1 U49361 ( .A(n48341), .ZN(n48287) );
  AOI21_X1 U49362 ( .B1(n48303), .B2(n48287), .A(n4035), .ZN(n48292) );
  NAND2_X1 U49363 ( .A1(n48369), .A2(n6986), .ZN(n48289) );
  NAND2_X1 U49364 ( .A1(n51072), .A2(n6986), .ZN(n48288) );
  NAND4_X1 U49365 ( .A1(n48290), .A2(n48380), .A3(n48289), .A4(n48288), .ZN(
        n48291) );
  OAI211_X1 U49366 ( .C1(n48369), .C2(n48380), .A(n48292), .B(n48291), .ZN(
        n48293) );
  NAND3_X1 U49367 ( .A1(n48295), .A2(n48294), .A3(n48293), .ZN(Plaintext[48])
         );
  NAND2_X1 U49368 ( .A1(n51728), .A2(n48381), .ZN(n48298) );
  NOR2_X1 U49369 ( .A1(n48381), .A2(n51072), .ZN(n48302) );
  NAND3_X1 U49370 ( .A1(n48302), .A2(n6986), .A3(n48380), .ZN(n48297) );
  AOI21_X1 U49371 ( .B1(n48298), .B2(n48297), .A(n48296), .ZN(n48301) );
  NAND2_X1 U49372 ( .A1(n48345), .A2(n51728), .ZN(n48347) );
  NOR2_X1 U49373 ( .A1(n48301), .A2(n48300), .ZN(n48323) );
  NAND2_X1 U49374 ( .A1(n48353), .A2(n48382), .ZN(n48388) );
  OR2_X1 U49375 ( .A1(n48388), .A2(n48366), .ZN(n48372) );
  NOR2_X1 U49376 ( .A1(n48302), .A2(n51728), .ZN(n48378) );
  OAI211_X1 U49377 ( .C1(n48392), .C2(n51087), .A(n48378), .B(n48303), .ZN(
        n48305) );
  AND3_X1 U49378 ( .A1(n48372), .A2(n48305), .A3(n48304), .ZN(n48322) );
  INV_X1 U49379 ( .A(n48307), .ZN(n48321) );
  NOR2_X1 U49380 ( .A1(n51356), .A2(n51728), .ZN(n48350) );
  NAND2_X1 U49381 ( .A1(n48381), .A2(n48382), .ZN(n48344) );
  INV_X1 U49382 ( .A(n48308), .ZN(n48317) );
  NAND2_X1 U49383 ( .A1(n48310), .A2(n48309), .ZN(n48313) );
  INV_X1 U49384 ( .A(n48311), .ZN(n48312) );
  OAI21_X1 U49385 ( .B1(n48313), .B2(n48312), .A(n48478), .ZN(n48316) );
  OR2_X1 U49386 ( .A1(n48314), .A2(n48478), .ZN(n48315) );
  NAND4_X1 U49387 ( .A1(n51072), .A2(n48317), .A3(n48316), .A4(n48315), .ZN(
        n48326) );
  NOR2_X1 U49388 ( .A1(n48381), .A2(n48326), .ZN(n48318) );
  AOI22_X1 U49389 ( .A1(n48350), .A2(n48319), .B1(n48351), .B2(n48318), .ZN(
        n48320) );
  NAND4_X1 U49390 ( .A1(n48323), .A2(n48322), .A3(n48321), .A4(n48320), .ZN(
        n48325) );
  INV_X1 U49391 ( .A(n4916), .ZN(n48324) );
  XNOR2_X1 U49392 ( .A(n48325), .B(n48324), .ZN(Plaintext[49]) );
  INV_X1 U49393 ( .A(n48326), .ZN(n48327) );
  NOR2_X1 U49394 ( .A1(n51356), .A2(n48340), .ZN(n48331) );
  OAI21_X1 U49395 ( .B1(n48353), .B2(n48381), .A(n48328), .ZN(n48330) );
  AOI22_X1 U49396 ( .A1(n48331), .A2(n48330), .B1(n48329), .B2(n48359), .ZN(
        n48336) );
  NAND2_X1 U49397 ( .A1(n48366), .A2(n48382), .ZN(n48334) );
  AOI21_X1 U49398 ( .B1(n48332), .B2(n51072), .A(n48353), .ZN(n48333) );
  OAI21_X1 U49399 ( .B1(n48369), .B2(n48334), .A(n48333), .ZN(n48335) );
  OAI211_X1 U49400 ( .C1(n48369), .C2(n48337), .A(n48336), .B(n48335), .ZN(
        n48339) );
  INV_X1 U49401 ( .A(n42668), .ZN(n48338) );
  XNOR2_X1 U49402 ( .A(n48339), .B(n48338), .ZN(Plaintext[50]) );
  NAND4_X1 U49403 ( .A1(n51356), .A2(n6986), .A3(n48353), .A4(n48340), .ZN(
        n48343) );
  INV_X1 U49404 ( .A(n48344), .ZN(n48349) );
  NAND3_X1 U49405 ( .A1(n48345), .A2(n52172), .A3(n48353), .ZN(n48346) );
  NAND2_X1 U49406 ( .A1(n48347), .A2(n48346), .ZN(n48348) );
  AOI21_X1 U49407 ( .B1(n48350), .B2(n48349), .A(n48348), .ZN(n48357) );
  INV_X1 U49408 ( .A(n48351), .ZN(n48352) );
  NAND4_X1 U49409 ( .A1(n48352), .A2(n48353), .A3(n51072), .A4(n48395), .ZN(
        n48356) );
  INV_X1 U49410 ( .A(n48395), .ZN(n48354) );
  NOR2_X1 U49411 ( .A1(n8103), .A2(n48382), .ZN(n48396) );
  INV_X1 U49412 ( .A(n4637), .ZN(n48358) );
  AND2_X1 U49413 ( .A1(n48359), .A2(n48381), .ZN(n48363) );
  INV_X1 U49414 ( .A(n48360), .ZN(n48362) );
  NAND2_X1 U49415 ( .A1(n48366), .A2(n51072), .ZN(n48367) );
  NAND3_X1 U49416 ( .A1(n48395), .A2(n48368), .A3(n48367), .ZN(n48371) );
  NAND2_X1 U49417 ( .A1(n48369), .A2(n51728), .ZN(n48370) );
  INV_X1 U49418 ( .A(n4827), .ZN(n48374) );
  XNOR2_X1 U49419 ( .A(n48375), .B(n48374), .ZN(Plaintext[52]) );
  INV_X1 U49420 ( .A(n48376), .ZN(n48379) );
  INV_X1 U49421 ( .A(n48388), .ZN(n48377) );
  AOI22_X1 U49422 ( .A1(n48379), .A2(n48378), .B1(n48377), .B2(n51356), .ZN(
        n48399) );
  OR2_X1 U49423 ( .A1(n48381), .A2(n51318), .ZN(n48386) );
  AOI21_X1 U49424 ( .B1(n51356), .B2(n52172), .A(n6986), .ZN(n48390) );
  INV_X1 U49425 ( .A(n48386), .ZN(n48387) );
  NAND2_X1 U49426 ( .A1(n48392), .A2(n51728), .ZN(n48393) );
  NAND3_X1 U49427 ( .A1(n48395), .A2(n48394), .A3(n48393), .ZN(n48397) );
  NAND2_X1 U49428 ( .A1(n48397), .A2(n48396), .ZN(n48398) );
  INV_X1 U49429 ( .A(n4781), .ZN(n48400) );
  XNOR2_X1 U49430 ( .A(n48401), .B(n48400), .ZN(Plaintext[53]) );
  NOR2_X1 U49431 ( .A1(n48405), .A2(n506), .ZN(n48406) );
  NOR3_X1 U49432 ( .A1(n48408), .A2(n48407), .A3(n48406), .ZN(n48422) );
  NOR3_X1 U49433 ( .A1(n48411), .A2(n48410), .A3(n48409), .ZN(n48419) );
  NAND3_X1 U49434 ( .A1(n48414), .A2(n506), .A3(n48412), .ZN(n48415) );
  OAI21_X1 U49435 ( .B1(n48417), .B2(n48416), .A(n48415), .ZN(n48418) );
  NOR2_X1 U49436 ( .A1(n48419), .A2(n48418), .ZN(n48420) );
  INV_X1 U49438 ( .A(n48438), .ZN(n48427) );
  NAND2_X1 U49439 ( .A1(n48424), .A2(n48423), .ZN(n48425) );
  OAI211_X1 U49440 ( .C1(n52178), .C2(n48427), .A(n48426), .B(n48425), .ZN(
        n48428) );
  INV_X1 U49441 ( .A(n48428), .ZN(n48447) );
  OR2_X1 U49442 ( .A1(n48430), .A2(n48429), .ZN(n48431) );
  NAND2_X1 U49443 ( .A1(n48432), .A2(n48434), .ZN(n48441) );
  NAND2_X1 U49444 ( .A1(n48434), .A2(n48433), .ZN(n48435) );
  NAND4_X1 U49445 ( .A1(n48438), .A2(n48437), .A3(n48436), .A4(n48435), .ZN(
        n48439) );
  OAI21_X1 U49446 ( .B1(n48441), .B2(n52178), .A(n48439), .ZN(n48442) );
  INV_X1 U49447 ( .A(n48442), .ZN(n48445) );
  NAND2_X1 U49448 ( .A1(n48443), .A2(n660), .ZN(n48444) );
  NAND2_X1 U49449 ( .A1(n51350), .A2(n48567), .ZN(n48587) );
  INV_X1 U49450 ( .A(n48587), .ZN(n48497) );
  INV_X1 U49451 ( .A(n48448), .ZN(n48468) );
  NAND3_X1 U49452 ( .A1(n48450), .A2(n48449), .A3(n7275), .ZN(n48453) );
  INV_X1 U49453 ( .A(n48455), .ZN(n48460) );
  OAI21_X1 U49454 ( .B1(n48460), .B2(n48459), .A(n48458), .ZN(n48467) );
  NOR2_X1 U49455 ( .A1(n51732), .A2(n48461), .ZN(n48466) );
  OR2_X1 U49456 ( .A1(n48469), .A2(n48468), .ZN(n48471) );
  OAI21_X1 U49457 ( .B1(n48474), .B2(n48479), .A(n48473), .ZN(n48476) );
  NAND3_X1 U49458 ( .A1(n48476), .A2(n48478), .A3(n48475), .ZN(n48496) );
  OAI21_X1 U49459 ( .B1(n48479), .B2(n48478), .A(n48477), .ZN(n48486) );
  INV_X1 U49460 ( .A(n48480), .ZN(n48484) );
  NAND2_X1 U49461 ( .A1(n48482), .A2(n51301), .ZN(n48483) );
  OAI211_X1 U49462 ( .C1(n48486), .C2(n48485), .A(n48484), .B(n48483), .ZN(
        n48490) );
  NAND2_X1 U49463 ( .A1(n48490), .A2(n48489), .ZN(n48495) );
  NAND3_X1 U49464 ( .A1(n48493), .A2(n48492), .A3(n48491), .ZN(n48494) );
  NOR2_X1 U49466 ( .A1(n48652), .A2(n48647), .ZN(n48605) );
  NAND2_X1 U49467 ( .A1(n48497), .A2(n48605), .ZN(n48562) );
  NAND3_X1 U49468 ( .A1(n48499), .A2(n48505), .A3(n48498), .ZN(n48504) );
  NAND2_X1 U49469 ( .A1(n48500), .A2(n52202), .ZN(n48503) );
  NAND2_X1 U49470 ( .A1(n48501), .A2(n48508), .ZN(n48502) );
  NAND3_X1 U49471 ( .A1(n48504), .A2(n48503), .A3(n48502), .ZN(n48516) );
  NAND2_X1 U49472 ( .A1(n48505), .A2(n48517), .ZN(n48506) );
  NOR2_X1 U49473 ( .A1(n48521), .A2(n48506), .ZN(n48509) );
  OAI21_X1 U49474 ( .B1(n48509), .B2(n48508), .A(n48507), .ZN(n48515) );
  AOI22_X1 U49475 ( .A1(n48513), .A2(n48512), .B1(n51451), .B2(n48510), .ZN(
        n48514) );
  NAND2_X1 U49476 ( .A1(n48519), .A2(n48518), .ZN(n48520) );
  OAI211_X1 U49477 ( .C1(n48523), .C2(n48522), .A(n48521), .B(n48520), .ZN(
        n48564) );
  NAND2_X1 U49478 ( .A1(n48546), .A2(n48524), .ZN(n48525) );
  OR2_X1 U49479 ( .A1(n48526), .A2(n48525), .ZN(n48533) );
  INV_X1 U49480 ( .A(n48527), .ZN(n48529) );
  AOI21_X1 U49481 ( .B1(n48530), .B2(n48529), .A(n48528), .ZN(n48532) );
  MUX2_X1 U49482 ( .A(n48533), .B(n48532), .S(n52059), .Z(n48560) );
  NAND2_X1 U49483 ( .A1(n48535), .A2(n48534), .ZN(n48537) );
  INV_X1 U49484 ( .A(n48536), .ZN(n48542) );
  AOI21_X1 U49485 ( .B1(n48538), .B2(n48537), .A(n48542), .ZN(n48545) );
  NAND3_X1 U49486 ( .A1(n48540), .A2(n48551), .A3(n48539), .ZN(n48541) );
  OAI21_X1 U49487 ( .B1(n48543), .B2(n48542), .A(n48541), .ZN(n48544) );
  NOR2_X1 U49488 ( .A1(n48545), .A2(n48544), .ZN(n48559) );
  NAND2_X1 U49489 ( .A1(n48553), .A2(n48552), .ZN(n48558) );
  INV_X1 U49490 ( .A(n48554), .ZN(n48555) );
  NAND2_X1 U49491 ( .A1(n48556), .A2(n48555), .ZN(n48557) );
  NAND2_X1 U49492 ( .A1(n48652), .A2(n52042), .ZN(n48600) );
  NAND4_X1 U49494 ( .A1(n48562), .A2(n48561), .A3(n48633), .A4(n48618), .ZN(
        n48563) );
  NAND2_X1 U49495 ( .A1(n48604), .A2(n48647), .ZN(n48616) );
  INV_X1 U49496 ( .A(n48633), .ZN(n48646) );
  OAI21_X1 U49497 ( .B1(n48616), .B2(n48587), .A(n48646), .ZN(n48579) );
  NAND2_X1 U49498 ( .A1(n48563), .A2(n48579), .ZN(n48573) );
  NAND3_X1 U49499 ( .A1(n48565), .A2(n48564), .A3(n48652), .ZN(n48566) );
  AND3_X1 U49500 ( .A1(n48581), .A2(n48633), .A3(n48566), .ZN(n48642) );
  INV_X1 U49501 ( .A(n48606), .ZN(n48638) );
  NOR2_X1 U49502 ( .A1(n48639), .A2(n48638), .ZN(n48568) );
  OAI21_X1 U49503 ( .B1(n48642), .B2(n48568), .A(n48647), .ZN(n48572) );
  NOR2_X1 U49504 ( .A1(n48606), .A2(n48633), .ZN(n48622) );
  NAND3_X1 U49505 ( .A1(n48649), .A2(n51382), .A3(n48622), .ZN(n48571) );
  AOI22_X1 U49506 ( .A1(n48583), .A2(n51350), .B1(n51382), .B2(n48647), .ZN(
        n48569) );
  OR2_X1 U49507 ( .A1(n48569), .A2(n48640), .ZN(n48570) );
  NAND4_X1 U49508 ( .A1(n48573), .A2(n48572), .A3(n48571), .A4(n48570), .ZN(
        n48575) );
  INV_X1 U49509 ( .A(n2947), .ZN(n48574) );
  XNOR2_X1 U49510 ( .A(n48575), .B(n48574), .ZN(Plaintext[54]) );
  NAND3_X1 U49511 ( .A1(n48604), .A2(n48640), .A3(n51382), .ZN(n48588) );
  OR2_X1 U49512 ( .A1(n51350), .A2(n52042), .ZN(n48641) );
  AND2_X1 U49513 ( .A1(n51382), .A2(n48606), .ZN(n48648) );
  OR2_X1 U49514 ( .A1(n48604), .A2(n52042), .ZN(n48612) );
  NAND2_X1 U49515 ( .A1(n6788), .A2(n48567), .ZN(n48615) );
  NAND3_X1 U49516 ( .A1(n48638), .A2(n51382), .A3(n48652), .ZN(n48580) );
  OAI22_X1 U49517 ( .A1(n48612), .A2(n48615), .B1(n48604), .B2(n48580), .ZN(
        n48577) );
  NAND2_X1 U49518 ( .A1(n48618), .A2(n48633), .ZN(n48576) );
  NAND2_X1 U49519 ( .A1(n48633), .A2(n51350), .ZN(n48589) );
  NAND2_X1 U49520 ( .A1(n48580), .A2(n48589), .ZN(n48582) );
  NAND4_X1 U49521 ( .A1(n48582), .A2(n48604), .A3(n48641), .A4(n48581), .ZN(
        n48584) );
  OR2_X1 U49522 ( .A1(n48587), .A2(n48640), .ZN(n48609) );
  INV_X1 U49523 ( .A(n4855), .ZN(n48585) );
  XNOR2_X1 U49524 ( .A(n48586), .B(n48585), .ZN(Plaintext[55]) );
  NOR2_X1 U49525 ( .A1(n48639), .A2(n48647), .ZN(n48593) );
  OR2_X1 U49526 ( .A1(n48646), .A2(n48587), .ZN(n48627) );
  NAND3_X1 U49527 ( .A1(n48613), .A2(n48649), .A3(n48627), .ZN(n48596) );
  AND2_X1 U49528 ( .A1(n48588), .A2(n48646), .ZN(n48592) );
  NAND2_X1 U49529 ( .A1(n48641), .A2(n51382), .ZN(n48591) );
  NAND2_X1 U49530 ( .A1(n48604), .A2(n48567), .ZN(n48621) );
  NAND2_X1 U49531 ( .A1(n48621), .A2(n48589), .ZN(n48590) );
  AOI22_X1 U49532 ( .A1(n48592), .A2(n48591), .B1(n48590), .B2(n48624), .ZN(
        n48595) );
  OR2_X1 U49533 ( .A1(n48593), .A2(n48618), .ZN(n48594) );
  NAND3_X1 U49534 ( .A1(n48596), .A2(n48595), .A3(n48594), .ZN(n48599) );
  INV_X1 U49535 ( .A(n48597), .ZN(n48598) );
  XNOR2_X1 U49536 ( .A(n48599), .B(n48598), .ZN(Plaintext[56]) );
  INV_X1 U49537 ( .A(n48600), .ZN(n48607) );
  AND2_X1 U49538 ( .A1(n48640), .A2(n51350), .ZN(n48632) );
  NAND2_X1 U49539 ( .A1(n48632), .A2(n51382), .ZN(n48602) );
  OAI211_X1 U49540 ( .C1(n48615), .C2(n48604), .A(n48603), .B(n48602), .ZN(
        n48611) );
  NAND3_X1 U49542 ( .A1(n51331), .A2(n48605), .A3(n48604), .ZN(n48610) );
  NAND3_X1 U49543 ( .A1(n48649), .A2(n48607), .A3(n51350), .ZN(n48608) );
  INV_X1 U49544 ( .A(n48648), .ZN(n48617) );
  INV_X1 U49545 ( .A(n48615), .ZN(n48625) );
  OAI21_X1 U49546 ( .B1(n48621), .B2(n48622), .A(n48620), .ZN(n48636) );
  INV_X1 U49547 ( .A(n48636), .ZN(n48628) );
  INV_X1 U49548 ( .A(n48622), .ZN(n48623) );
  OAI21_X1 U49549 ( .B1(n48625), .B2(n48624), .A(n48623), .ZN(n48626) );
  NAND4_X1 U49550 ( .A1(n48629), .A2(n48628), .A3(n48627), .A4(n48626), .ZN(
        n48631) );
  INV_X1 U49551 ( .A(n4654), .ZN(n48630) );
  XNOR2_X1 U49552 ( .A(n48631), .B(n48630), .ZN(Plaintext[58]) );
  OAI21_X1 U49553 ( .B1(n52042), .B2(n48633), .A(n48632), .ZN(n48635) );
  NAND2_X1 U49554 ( .A1(n48636), .A2(n48635), .ZN(n48656) );
  OAI21_X1 U49555 ( .B1(n48649), .B2(n48638), .A(n51331), .ZN(n48644) );
  OAI21_X1 U49556 ( .B1(n48641), .B2(n48640), .A(n48639), .ZN(n48643) );
  AOI21_X1 U49557 ( .B1(n48644), .B2(n48643), .A(n48642), .ZN(n48655) );
  NAND3_X1 U49558 ( .A1(n48649), .A2(n48646), .A3(n48567), .ZN(n48651) );
  NAND3_X1 U49559 ( .A1(n48649), .A2(n48648), .A3(n48647), .ZN(n48650) );
  NAND2_X1 U49560 ( .A1(n48651), .A2(n48650), .ZN(n48653) );
  NAND2_X1 U49561 ( .A1(n48653), .A2(n48652), .ZN(n48654) );
  NAND3_X1 U49562 ( .A1(n48656), .A2(n48655), .A3(n48654), .ZN(n48658) );
  XNOR2_X1 U49563 ( .A(n48658), .B(n48657), .ZN(Plaintext[59]) );
  NAND3_X1 U49564 ( .A1(n48702), .A2(n48714), .A3(n48659), .ZN(n48712) );
  NAND2_X1 U49565 ( .A1(n48708), .A2(n51659), .ZN(n48661) );
  NAND2_X1 U49566 ( .A1(n48661), .A2(n52157), .ZN(n48662) );
  NAND3_X1 U49567 ( .A1(n48663), .A2(n48712), .A3(n48662), .ZN(n48665) );
  NAND2_X1 U49568 ( .A1(n48665), .A2(n48664), .ZN(n48679) );
  NAND2_X1 U49569 ( .A1(n48666), .A2(n48685), .ZN(n48672) );
  NAND2_X1 U49570 ( .A1(n48713), .A2(n48703), .ZN(n48668) );
  OAI211_X1 U49571 ( .C1(n48669), .C2(n48703), .A(n48668), .B(n48667), .ZN(
        n48671) );
  NAND3_X1 U49572 ( .A1(n48682), .A2(n48714), .A3(n48703), .ZN(n48670) );
  AND3_X1 U49573 ( .A1(n48671), .A2(n48672), .A3(n48670), .ZN(n48678) );
  NAND3_X1 U49574 ( .A1(n48675), .A2(n48695), .A3(n48674), .ZN(n48676) );
  INV_X1 U49578 ( .A(n48682), .ZN(n48683) );
  AOI21_X1 U49579 ( .B1(n48684), .B2(n48713), .A(n48683), .ZN(n48692) );
  INV_X1 U49580 ( .A(n48708), .ZN(n48686) );
  OAI21_X1 U49581 ( .B1(n48686), .B2(n48696), .A(n48685), .ZN(n48691) );
  NOR2_X1 U49582 ( .A1(n48687), .A2(n48697), .ZN(n48689) );
  AOI21_X1 U49583 ( .B1(n48689), .B2(n48688), .A(n48707), .ZN(n48690) );
  OAI211_X1 U49584 ( .C1(n48692), .C2(n48711), .A(n48691), .B(n48690), .ZN(
        n48694) );
  NAND2_X1 U49587 ( .A1(n48702), .A2(n48703), .ZN(n48700) );
  AOI21_X1 U49588 ( .B1(n48701), .B2(n51659), .A(n48697), .ZN(n48699) );
  OAI21_X1 U49589 ( .B1(n48707), .B2(n48700), .A(n48699), .ZN(n48706) );
  OAI22_X1 U49590 ( .A1(n48704), .A2(n48703), .B1(n48702), .B2(n48701), .ZN(
        n48705) );
  NOR2_X1 U49591 ( .A1(n48706), .A2(n48705), .ZN(n48717) );
  INV_X1 U49592 ( .A(n48707), .ZN(n48710) );
  OAI22_X1 U49593 ( .A1(n48711), .A2(n48710), .B1(n48709), .B2(n48708), .ZN(
        n48716) );
  OAI21_X1 U49594 ( .B1(n48714), .B2(n48713), .A(n48712), .ZN(n48715) );
  NOR3_X1 U49595 ( .A1(n48717), .A2(n48716), .A3(n48715), .ZN(n48718) );
  INV_X1 U49596 ( .A(n4645), .ZN(n48719) );
  AND2_X1 U49597 ( .A1(n48721), .A2(n48720), .ZN(n48724) );
  OAI21_X1 U49598 ( .B1(n48750), .B2(n48722), .A(n52067), .ZN(n48723) );
  AOI21_X1 U49599 ( .B1(n48724), .B2(n48723), .A(n48759), .ZN(n48743) );
  OR2_X1 U49600 ( .A1(n48730), .A2(n48729), .ZN(n48725) );
  NOR2_X1 U49601 ( .A1(n48779), .A2(n48725), .ZN(n48728) );
  NOR2_X1 U49602 ( .A1(n48745), .A2(n48726), .ZN(n48727) );
  NOR2_X1 U49603 ( .A1(n48728), .A2(n48727), .ZN(n48737) );
  NAND2_X1 U49604 ( .A1(n48780), .A2(n48729), .ZN(n48733) );
  NAND2_X1 U49605 ( .A1(n52067), .A2(n48730), .ZN(n48731) );
  NAND2_X1 U49606 ( .A1(n48731), .A2(n48734), .ZN(n48732) );
  OAI211_X1 U49607 ( .C1(n48734), .C2(n48744), .A(n48733), .B(n48732), .ZN(
        n48735) );
  NAND4_X1 U49608 ( .A1(n48737), .A2(n4490), .A3(n48735), .A4(n48736), .ZN(
        n48742) );
  INV_X1 U49609 ( .A(n4490), .ZN(n48738) );
  NAND2_X1 U49610 ( .A1(n48743), .A2(n48738), .ZN(n48741) );
  NAND3_X1 U49611 ( .A1(n48737), .A2(n48736), .A3(n48735), .ZN(n48739) );
  NAND2_X1 U49612 ( .A1(n48739), .A2(n48738), .ZN(n48740) );
  OAI211_X1 U49613 ( .C1(n48743), .C2(n48742), .A(n48741), .B(n48740), .ZN(
        Plaintext[66]) );
  NAND2_X1 U49614 ( .A1(n48750), .A2(n48747), .ZN(n48785) );
  AOI21_X1 U49616 ( .B1(n48785), .B2(n52051), .A(n52223), .ZN(n48756) );
  AOI21_X1 U49617 ( .B1(n48768), .B2(n48747), .A(n48760), .ZN(n48755) );
  INV_X1 U49618 ( .A(n48779), .ZN(n48748) );
  OAI21_X1 U49619 ( .B1(n48750), .B2(n48749), .A(n48748), .ZN(n48754) );
  INV_X1 U49620 ( .A(n48766), .ZN(n48752) );
  NAND3_X1 U49621 ( .A1(n48752), .A2(n994), .A3(n48751), .ZN(n48753) );
  INV_X1 U49623 ( .A(n4558), .ZN(n48757) );
  AND2_X1 U49625 ( .A1(n48759), .A2(n48760), .ZN(n48783) );
  OAI211_X1 U49626 ( .C1(n48768), .C2(n48762), .A(n48783), .B(n52067), .ZN(
        n48774) );
  INV_X1 U49627 ( .A(n48763), .ZN(n48767) );
  INV_X1 U49628 ( .A(n48764), .ZN(n48765) );
  AOI21_X1 U49629 ( .B1(n48767), .B2(n48766), .A(n48765), .ZN(n48772) );
  NAND3_X1 U49630 ( .A1(n48770), .A2(n48769), .A3(n48768), .ZN(n48771) );
  NAND4_X1 U49631 ( .A1(n48774), .A2(n48773), .A3(n48772), .A4(n48771), .ZN(
        n48776) );
  XNOR2_X1 U49632 ( .A(n48776), .B(n48775), .ZN(Plaintext[69]) );
  INV_X1 U49633 ( .A(n48777), .ZN(n48788) );
  NAND2_X1 U49634 ( .A1(n48780), .A2(n48779), .ZN(n48781) );
  AOI22_X1 U49635 ( .A1(n48784), .A2(n48783), .B1(n48782), .B2(n48781), .ZN(
        n48787) );
  NAND4_X1 U49636 ( .A1(n48788), .A2(n48787), .A3(n48786), .A4(n48785), .ZN(
        n48790) );
  INV_X1 U49637 ( .A(n4845), .ZN(n48789) );
  XNOR2_X1 U49638 ( .A(n48790), .B(n48789), .ZN(Plaintext[70]) );
  OAI21_X1 U49639 ( .B1(n48817), .B2(n48792), .A(n48791), .ZN(n48795) );
  INV_X1 U49640 ( .A(n48819), .ZN(n48838) );
  NAND2_X1 U49641 ( .A1(n48793), .A2(n48830), .ZN(n48794) );
  AOI22_X1 U49642 ( .A1(n48796), .A2(n48795), .B1(n48838), .B2(n48794), .ZN(
        n48802) );
  INV_X1 U49643 ( .A(n48806), .ZN(n48797) );
  OAI21_X1 U49644 ( .B1(n48798), .B2(n48816), .A(n48797), .ZN(n48801) );
  INV_X1 U49645 ( .A(n4650), .ZN(n48803) );
  NAND3_X1 U49646 ( .A1(n48838), .A2(n48805), .A3(n48804), .ZN(n48813) );
  NAND2_X1 U49647 ( .A1(n48806), .A2(n52434), .ZN(n48807) );
  OAI211_X1 U49648 ( .C1(n48819), .C2(n48816), .A(n48831), .B(n48807), .ZN(
        n48811) );
  INV_X1 U49649 ( .A(n48823), .ZN(n48809) );
  NAND3_X1 U49650 ( .A1(n48817), .A2(n48809), .A3(n45743), .ZN(n48810) );
  INV_X1 U49651 ( .A(n48814), .ZN(n48815) );
  NAND3_X1 U49652 ( .A1(n48817), .A2(n52434), .A3(n48816), .ZN(n48818) );
  NAND2_X1 U49653 ( .A1(n48820), .A2(n48819), .ZN(n48842) );
  AOI21_X1 U49654 ( .B1(n48824), .B2(n48823), .A(n48834), .ZN(n48825) );
  OAI21_X1 U49655 ( .B1(n48827), .B2(n48826), .A(n48825), .ZN(n48841) );
  NOR2_X1 U49656 ( .A1(n48829), .A2(n48828), .ZN(n48835) );
  NAND2_X1 U49657 ( .A1(n48831), .A2(n48830), .ZN(n48832) );
  AOI22_X1 U49658 ( .A1(n48835), .A2(n48834), .B1(n48833), .B2(n48832), .ZN(
        n48840) );
  NOR2_X1 U49659 ( .A1(n48836), .A2(n51328), .ZN(n48837) );
  NAND2_X1 U49660 ( .A1(n48838), .A2(n48837), .ZN(n48839) );
  NAND4_X1 U49661 ( .A1(n48842), .A2(n48841), .A3(n48840), .A4(n48839), .ZN(
        n48845) );
  INV_X1 U49662 ( .A(n48843), .ZN(n48844) );
  XNOR2_X1 U49663 ( .A(n48845), .B(n48844), .ZN(Plaintext[77]) );
  NOR2_X1 U49664 ( .A1(n48853), .A2(n51688), .ZN(n48854) );
  OAI21_X1 U49665 ( .B1(n48854), .B2(n48888), .A(n48846), .ZN(n48849) );
  INV_X1 U49666 ( .A(n48912), .ZN(n48900) );
  MUX2_X1 U49667 ( .A(n48849), .B(n48848), .S(n48900), .Z(n48858) );
  NAND2_X1 U49668 ( .A1(n48918), .A2(n48886), .ZN(n48851) );
  INV_X1 U49669 ( .A(n48919), .ZN(n48862) );
  NAND2_X1 U49670 ( .A1(n5078), .A2(n48912), .ZN(n48906) );
  NOR2_X1 U49671 ( .A1(n3631), .A2(n48906), .ZN(n48850) );
  AND2_X1 U49672 ( .A1(n48919), .A2(n48853), .ZN(n48874) );
  INV_X1 U49673 ( .A(n48908), .ZN(n48899) );
  NOR2_X1 U49674 ( .A1(n48899), .A2(n48905), .ZN(n48855) );
  AOI22_X1 U49675 ( .A1(n48874), .A2(n48855), .B1(n48854), .B2(n48898), .ZN(
        n48856) );
  INV_X1 U49676 ( .A(n1336), .ZN(n48859) );
  AOI21_X1 U49677 ( .B1(n51689), .B2(n48886), .A(n48899), .ZN(n48861) );
  OAI21_X1 U49678 ( .B1(n48920), .B2(n48874), .A(n5081), .ZN(n48860) );
  OAI21_X1 U49679 ( .B1(n48861), .B2(n48862), .A(n48860), .ZN(n48869) );
  NAND3_X1 U49680 ( .A1(n48913), .A2(n48862), .A3(n48905), .ZN(n48864) );
  NAND2_X1 U49681 ( .A1(n48905), .A2(n51689), .ZN(n48863) );
  OAI22_X1 U49682 ( .A1(n48875), .A2(n48864), .B1(n48920), .B2(n48863), .ZN(
        n48865) );
  INV_X1 U49683 ( .A(n48865), .ZN(n48868) );
  INV_X1 U49684 ( .A(n48918), .ZN(n48866) );
  OAI21_X1 U49685 ( .B1(n48915), .B2(n48898), .A(n48866), .ZN(n48867) );
  NAND3_X1 U49686 ( .A1(n48869), .A2(n48868), .A3(n48867), .ZN(n48871) );
  INV_X1 U49687 ( .A(n4939), .ZN(n48870) );
  XNOR2_X1 U49688 ( .A(n48871), .B(n48870), .ZN(Plaintext[80]) );
  AND2_X1 U49689 ( .A1(n48919), .A2(n51689), .ZN(n48872) );
  INV_X1 U49690 ( .A(n48886), .ZN(n48881) );
  NAND3_X1 U49691 ( .A1(n48875), .A2(n5081), .A3(n48874), .ZN(n48876) );
  OAI21_X1 U49692 ( .B1(n48908), .B2(n48906), .A(n48877), .ZN(n48878) );
  INV_X1 U49693 ( .A(n48878), .ZN(n48884) );
  NOR2_X1 U49694 ( .A1(n48879), .A2(n48919), .ZN(n48880) );
  OAI211_X1 U49695 ( .C1(n48882), .C2(n48888), .A(n48881), .B(n48908), .ZN(
        n48883) );
  OR3_X1 U49696 ( .A1(n48887), .A2(n48905), .A3(n48886), .ZN(n48895) );
  INV_X1 U49698 ( .A(n48911), .ZN(n48891) );
  AOI22_X1 U49699 ( .A1(n48916), .A2(n48889), .B1(n48891), .B2(n48915), .ZN(
        n48894) );
  NAND2_X1 U49700 ( .A1(n48918), .A2(n3782), .ZN(n48890) );
  OAI211_X1 U49701 ( .C1(n48898), .C2(n48900), .A(n48891), .B(n48890), .ZN(
        n48892) );
  NAND4_X1 U49702 ( .A1(n48895), .A2(n48894), .A3(n48893), .A4(n48892), .ZN(
        n48897) );
  INV_X1 U49703 ( .A(n4026), .ZN(n48896) );
  XNOR2_X1 U49704 ( .A(n48897), .B(n48896), .ZN(Plaintext[82]) );
  NAND2_X1 U49705 ( .A1(n48899), .A2(n48898), .ZN(n48903) );
  INV_X1 U49706 ( .A(n48906), .ZN(n48907) );
  NOR2_X1 U49707 ( .A1(n48900), .A2(n48919), .ZN(n48901) );
  AOI22_X1 U49708 ( .A1(n48905), .A2(n48907), .B1(n48901), .B2(n48908), .ZN(
        n48902) );
  MUX2_X1 U49709 ( .A(n48903), .B(n48902), .S(n51688), .Z(n48924) );
  NOR3_X1 U49710 ( .A1(n48906), .A2(n48905), .A3(n51688), .ZN(n48909) );
  AOI22_X1 U49711 ( .A1(n48909), .A2(n48908), .B1(n48911), .B2(n48907), .ZN(
        n48923) );
  INV_X1 U49712 ( .A(n48910), .ZN(n48917) );
  OAI21_X1 U49713 ( .B1(n48913), .B2(n48912), .A(n48911), .ZN(n48914) );
  OAI211_X1 U49714 ( .C1(n48917), .C2(n48916), .A(n48915), .B(n48914), .ZN(
        n48922) );
  NAND3_X1 U49715 ( .A1(n48920), .A2(n48919), .A3(n48918), .ZN(n48921) );
  NAND4_X1 U49716 ( .A1(n48924), .A2(n48923), .A3(n48922), .A4(n48921), .ZN(
        n48926) );
  INV_X1 U49717 ( .A(n4653), .ZN(n48925) );
  XNOR2_X1 U49718 ( .A(n48926), .B(n48925), .ZN(Plaintext[83]) );
  MUX2_X1 U49719 ( .A(n48929), .B(n48928), .S(n48927), .Z(n48940) );
  OAI22_X1 U49720 ( .A1(n48932), .A2(n48931), .B1(n51510), .B2(n48930), .ZN(
        n48933) );
  NOR2_X1 U49721 ( .A1(n48934), .A2(n48933), .ZN(n48939) );
  NAND2_X1 U49722 ( .A1(n48952), .A2(n48935), .ZN(n48936) );
  NAND3_X1 U49723 ( .A1(n48937), .A2(n48973), .A3(n48936), .ZN(n48938) );
  NOR2_X1 U49724 ( .A1(n48955), .A2(n48941), .ZN(n48946) );
  NAND2_X1 U49725 ( .A1(n48943), .A2(n48942), .ZN(n48945) );
  MUX2_X1 U49726 ( .A(n48946), .B(n48945), .S(n51478), .Z(n48947) );
  NOR2_X1 U49727 ( .A1(n48948), .A2(n48947), .ZN(n48949) );
  XNOR2_X1 U49728 ( .A(n48949), .B(n4752), .ZN(Plaintext[84]) );
  NOR2_X1 U49729 ( .A1(n48951), .A2(n48950), .ZN(n48953) );
  OAI22_X1 U49730 ( .A1(n48972), .A2(n48953), .B1(n51510), .B2(n48952), .ZN(
        n48964) );
  INV_X1 U49731 ( .A(n48954), .ZN(n48967) );
  NAND2_X1 U49732 ( .A1(n48955), .A2(n48967), .ZN(n48956) );
  NAND2_X1 U49733 ( .A1(n48956), .A2(n48970), .ZN(n48963) );
  NAND2_X1 U49734 ( .A1(n48958), .A2(n48957), .ZN(n48959) );
  OAI21_X1 U49735 ( .B1(n48960), .B2(n48959), .A(n46954), .ZN(n48961) );
  NAND2_X1 U49736 ( .A1(n48961), .A2(n47476), .ZN(n48962) );
  NAND3_X1 U49737 ( .A1(n48964), .A2(n48963), .A3(n48962), .ZN(n48966) );
  INV_X1 U49738 ( .A(n4208), .ZN(n48965) );
  XNOR2_X1 U49739 ( .A(n48966), .B(n48965), .ZN(Plaintext[86]) );
  NAND2_X1 U49740 ( .A1(n48968), .A2(n48967), .ZN(n48969) );
  OAI211_X1 U49741 ( .C1(n48970), .C2(n51511), .A(n48969), .B(n48971), .ZN(
        n48980) );
  AOI21_X1 U49742 ( .B1(n51511), .B2(n48974), .A(n48973), .ZN(n48977) );
  NAND2_X1 U49743 ( .A1(n48977), .A2(n48976), .ZN(n48978) );
  NAND4_X1 U49744 ( .A1(n48981), .A2(n48980), .A3(n48979), .A4(n48978), .ZN(
        n48983) );
  INV_X1 U49745 ( .A(n4823), .ZN(n48982) );
  XNOR2_X1 U49746 ( .A(n48983), .B(n48982), .ZN(Plaintext[88]) );
  NOR2_X1 U49747 ( .A1(n49020), .A2(n49021), .ZN(n49030) );
  NAND2_X1 U49748 ( .A1(n49030), .A2(n51310), .ZN(n48985) );
  OAI22_X1 U49749 ( .A1(n48985), .A2(n49017), .B1(n48984), .B2(n51321), .ZN(
        n48986) );
  AOI21_X1 U49750 ( .B1(n51310), .B2(n48987), .A(n48986), .ZN(n48998) );
  OAI22_X1 U49751 ( .A1(n48988), .A2(n49019), .B1(n6389), .B2(n51321), .ZN(
        n48991) );
  INV_X1 U49752 ( .A(n48992), .ZN(n48997) );
  NAND4_X1 U49753 ( .A1(n49016), .A2(n49029), .A3(n49008), .A4(n49021), .ZN(
        n48993) );
  OAI22_X1 U49754 ( .A1(n49006), .A2(n52179), .B1(n49029), .B2(n49019), .ZN(
        n48995) );
  NAND4_X1 U49755 ( .A1(n48995), .A2(n49007), .A3(n48994), .A4(n51321), .ZN(
        n48996) );
  INV_X1 U49756 ( .A(n4818), .ZN(n48999) );
  AND2_X1 U49757 ( .A1(n51310), .A2(n51397), .ZN(n49001) );
  OAI21_X1 U49758 ( .B1(n49006), .B2(n49029), .A(n51321), .ZN(n49000) );
  OAI21_X1 U49759 ( .B1(n49002), .B2(n49001), .A(n49000), .ZN(n49013) );
  AND2_X1 U49760 ( .A1(n52179), .A2(n49021), .ZN(n49005) );
  AOI22_X1 U49761 ( .A1(n49046), .A2(n49005), .B1(n49004), .B2(n49003), .ZN(
        n49012) );
  NAND3_X1 U49762 ( .A1(n49006), .A2(n51321), .A3(n52179), .ZN(n49010) );
  NAND3_X1 U49763 ( .A1(n49008), .A2(n49007), .A3(n49021), .ZN(n49009) );
  AND2_X1 U49764 ( .A1(n49010), .A2(n49009), .ZN(n49011) );
  NAND4_X1 U49765 ( .A1(n49013), .A2(n49012), .A3(n49011), .A4(n49031), .ZN(
        n49015) );
  INV_X1 U49766 ( .A(n4624), .ZN(n49014) );
  XNOR2_X1 U49767 ( .A(n49015), .B(n49014), .ZN(Plaintext[92]) );
  NOR2_X1 U49768 ( .A1(n51397), .A2(n49021), .ZN(n49043) );
  NOR2_X1 U49769 ( .A1(n49017), .A2(n653), .ZN(n49018) );
  NAND3_X1 U49770 ( .A1(n51321), .A2(n49019), .A3(n51397), .ZN(n49023) );
  AOI21_X1 U49771 ( .B1(n49021), .B2(n49020), .A(n52179), .ZN(n49022) );
  OAI211_X1 U49772 ( .C1(n49024), .C2(n51321), .A(n49023), .B(n49022), .ZN(
        n49027) );
  OAI21_X1 U49773 ( .B1(n49025), .B2(n51321), .A(n52179), .ZN(n49026) );
  AND2_X1 U49774 ( .A1(n49029), .A2(n51310), .ZN(n49038) );
  NAND2_X1 U49775 ( .A1(n49034), .A2(n51321), .ZN(n49035) );
  AND2_X1 U49776 ( .A1(n49036), .A2(n49035), .ZN(n49051) );
  NAND3_X1 U49777 ( .A1(n49039), .A2(n49038), .A3(n49037), .ZN(n49050) );
  INV_X1 U49778 ( .A(n49040), .ZN(n49041) );
  OR2_X1 U49779 ( .A1(n49042), .A2(n49041), .ZN(n49049) );
  INV_X1 U49780 ( .A(n49043), .ZN(n49045) );
  OAI211_X1 U49781 ( .C1(n52179), .C2(n49046), .A(n49045), .B(n49044), .ZN(
        n49048) );
  NAND4_X1 U49782 ( .A1(n49051), .A2(n49050), .A3(n49049), .A4(n49048), .ZN(
        n49053) );
  INV_X1 U49783 ( .A(n4275), .ZN(n49052) );
  XNOR2_X1 U49784 ( .A(n49053), .B(n49052), .ZN(Plaintext[94]) );
  OR2_X1 U49785 ( .A1(n49065), .A2(n49054), .ZN(n49073) );
  INV_X1 U49786 ( .A(n49073), .ZN(n49056) );
  INV_X1 U49787 ( .A(n49103), .ZN(n49055) );
  AOI22_X1 U49788 ( .A1(n49056), .A2(n49067), .B1(n49081), .B2(n49055), .ZN(
        n49062) );
  INV_X1 U49789 ( .A(n49101), .ZN(n49092) );
  AND2_X1 U49790 ( .A1(n49112), .A2(n49117), .ZN(n49071) );
  NAND2_X1 U49791 ( .A1(n49101), .A2(n49071), .ZN(n49125) );
  NOR2_X1 U49792 ( .A1(n49125), .A2(n49128), .ZN(n49058) );
  NAND2_X1 U49793 ( .A1(n49115), .A2(n49117), .ZN(n49059) );
  NAND3_X1 U49794 ( .A1(n49072), .A2(n49100), .A3(n49059), .ZN(n49060) );
  INV_X1 U49795 ( .A(n4597), .ZN(n49063) );
  AOI22_X1 U49797 ( .A1(n49067), .A2(n49092), .B1(n49066), .B2(n49065), .ZN(
        n49077) );
  OR2_X1 U49798 ( .A1(n49119), .A2(n49112), .ZN(n49093) );
  INV_X1 U49800 ( .A(n49118), .ZN(n49076) );
  OR2_X1 U49801 ( .A1(n49068), .A2(n49127), .ZN(n49069) );
  OAI211_X1 U49802 ( .C1(n49072), .C2(n49071), .A(n49070), .B(n49069), .ZN(
        n49075) );
  NAND3_X1 U49803 ( .A1(n49073), .A2(n49117), .A3(n49103), .ZN(n49074) );
  NAND4_X1 U49804 ( .A1(n49077), .A2(n49076), .A3(n49075), .A4(n49074), .ZN(
        n49079) );
  INV_X1 U49805 ( .A(n2903), .ZN(n49078) );
  XNOR2_X1 U49806 ( .A(n49079), .B(n49078), .ZN(Plaintext[98]) );
  INV_X1 U49807 ( .A(n51320), .ZN(n49084) );
  OAI22_X1 U49808 ( .A1(n49085), .A2(n49084), .B1(n49083), .B2(n49082), .ZN(
        n49086) );
  AOI21_X1 U49809 ( .B1(n49088), .B2(n49087), .A(n49086), .ZN(n49097) );
  INV_X1 U49810 ( .A(n49100), .ZN(n49090) );
  OAI21_X1 U49811 ( .B1(n49118), .B2(n49091), .A(n49090), .ZN(n49108) );
  NAND2_X1 U49812 ( .A1(n49092), .A2(n49122), .ZN(n49131) );
  INV_X1 U49813 ( .A(n49093), .ZN(n49095) );
  NAND2_X1 U49814 ( .A1(n49095), .A2(n49094), .ZN(n49096) );
  NAND4_X1 U49815 ( .A1(n49097), .A2(n49108), .A3(n49131), .A4(n49096), .ZN(
        n49099) );
  INV_X1 U49816 ( .A(n4554), .ZN(n49098) );
  XNOR2_X1 U49817 ( .A(n49099), .B(n49098), .ZN(Plaintext[99]) );
  NAND3_X1 U49818 ( .A1(n49101), .A2(n49127), .A3(n49100), .ZN(n49102) );
  OAI22_X1 U49819 ( .A1(n49104), .A2(n49128), .B1(n44772), .B2(n49103), .ZN(
        n49105) );
  OAI211_X1 U49820 ( .C1(n49108), .C2(n49107), .A(n8768), .B(n49106), .ZN(
        n49111) );
  INV_X1 U49821 ( .A(n49109), .ZN(n49110) );
  XNOR2_X1 U49822 ( .A(n49111), .B(n49110), .ZN(Plaintext[100]) );
  OAI21_X1 U49823 ( .B1(n49114), .B2(n51320), .A(n49112), .ZN(n49116) );
  NAND2_X1 U49824 ( .A1(n49116), .A2(n49115), .ZN(n49120) );
  AOI22_X1 U49825 ( .A1(n49120), .A2(n49119), .B1(n49117), .B2(n49118), .ZN(
        n49134) );
  NAND2_X1 U49826 ( .A1(n49123), .A2(n49122), .ZN(n49133) );
  NAND2_X1 U49827 ( .A1(n49125), .A2(n49124), .ZN(n49130) );
  NAND3_X1 U49828 ( .A1(n49128), .A2(n49127), .A3(n49126), .ZN(n49129) );
  NAND2_X1 U49829 ( .A1(n49130), .A2(n49129), .ZN(n49132) );
  NAND4_X1 U49830 ( .A1(n49134), .A2(n49133), .A3(n49132), .A4(n49131), .ZN(
        n49136) );
  INV_X1 U49831 ( .A(n1313), .ZN(n49135) );
  XNOR2_X1 U49832 ( .A(n49136), .B(n49135), .ZN(Plaintext[101]) );
  NAND2_X1 U49833 ( .A1(n49138), .A2(n49137), .ZN(n49140) );
  NAND3_X1 U49834 ( .A1(n49141), .A2(n49140), .A3(n49139), .ZN(n49144) );
  OAI21_X1 U49835 ( .B1(n49148), .B2(n49147), .A(n49146), .ZN(n49153) );
  AND2_X1 U49836 ( .A1(n49150), .A2(n49149), .ZN(n49152) );
  AOI22_X1 U49837 ( .A1(n51515), .A2(n49153), .B1(n49152), .B2(n49151), .ZN(
        n49155) );
  OAI21_X1 U49839 ( .B1(n49159), .B2(n49158), .A(n49157), .ZN(n49160) );
  INV_X1 U49840 ( .A(n49160), .ZN(n49180) );
  NOR3_X1 U49841 ( .A1(n49162), .A2(n49163), .A3(n49161), .ZN(n49166) );
  NOR2_X1 U49842 ( .A1(n49170), .A2(n49163), .ZN(n49164) );
  NAND2_X1 U49843 ( .A1(n49169), .A2(n49168), .ZN(n49172) );
  NAND3_X1 U49844 ( .A1(n49172), .A2(n49171), .A3(n49170), .ZN(n49173) );
  NOR2_X1 U49845 ( .A1(n49175), .A2(n49174), .ZN(n49176) );
  INV_X1 U49847 ( .A(n49342), .ZN(n49229) );
  NAND3_X1 U49848 ( .A1(n49721), .A2(n49707), .A3(n49719), .ZN(n49182) );
  AND2_X1 U49849 ( .A1(n49182), .A2(n49714), .ZN(n49187) );
  NAND2_X1 U49850 ( .A1(n49710), .A2(n51295), .ZN(n49183) );
  OR2_X1 U49851 ( .A1(n49184), .A2(n49183), .ZN(n49186) );
  NAND2_X1 U49852 ( .A1(n49191), .A2(n52052), .ZN(n49185) );
  NAND4_X1 U49853 ( .A1(n49188), .A2(n49187), .A3(n49186), .A4(n49185), .ZN(
        n49196) );
  OAI211_X1 U49854 ( .C1(n49189), .C2(n49725), .A(n49713), .B(n49717), .ZN(
        n49194) );
  NAND2_X1 U49855 ( .A1(n49190), .A2(n49725), .ZN(n49192) );
  NAND2_X1 U49856 ( .A1(n49192), .A2(n49191), .ZN(n49193) );
  NOR2_X1 U49857 ( .A1(n49198), .A2(n49197), .ZN(n49202) );
  AOI22_X1 U49858 ( .A1(n49202), .A2(n49201), .B1(n49200), .B2(n49199), .ZN(
        n49204) );
  OR2_X1 U49861 ( .A1(n49208), .A2(n49207), .ZN(n49214) );
  INV_X1 U49862 ( .A(n49214), .ZN(n49210) );
  NAND2_X1 U49863 ( .A1(n49210), .A2(n49209), .ZN(n49211) );
  NAND2_X1 U49864 ( .A1(n49212), .A2(n49211), .ZN(n49220) );
  AOI21_X1 U49865 ( .B1(n49215), .B2(n49214), .A(n49213), .ZN(n49217) );
  INV_X1 U49866 ( .A(n49222), .ZN(n49224) );
  OAI211_X1 U49867 ( .C1(n49226), .C2(n49225), .A(n49224), .B(n49223), .ZN(
        n49227) );
  INV_X1 U49868 ( .A(n49227), .ZN(n49228) );
  OAI21_X1 U49869 ( .B1(n49229), .B2(n49376), .A(n49285), .ZN(n49284) );
  NAND2_X1 U49870 ( .A1(n49230), .A2(n49232), .ZN(n49240) );
  INV_X1 U49872 ( .A(n49243), .ZN(n49236) );
  NAND2_X1 U49873 ( .A1(n49236), .A2(n49235), .ZN(n49238) );
  OAI21_X1 U49874 ( .B1(n51095), .B2(n49242), .A(n49241), .ZN(n49245) );
  AOI21_X1 U49875 ( .B1(n49397), .B2(n49254), .A(n49243), .ZN(n49244) );
  NAND2_X1 U49876 ( .A1(n49245), .A2(n49244), .ZN(n49259) );
  NAND2_X1 U49878 ( .A1(n49248), .A2(n49247), .ZN(n49249) );
  NAND2_X1 U49879 ( .A1(n49250), .A2(n49249), .ZN(n49253) );
  OAI21_X1 U49880 ( .B1(n49253), .B2(n49252), .A(n49251), .ZN(n49258) );
  AND2_X1 U49881 ( .A1(n49255), .A2(n49256), .ZN(n49257) );
  AOI22_X1 U49882 ( .A1(n49262), .A2(n49277), .B1(n49261), .B2(n49275), .ZN(
        n49271) );
  OR2_X1 U49883 ( .A1(n49263), .A2(n52086), .ZN(n49264) );
  OAI211_X1 U49884 ( .C1(n49278), .C2(n49275), .A(n49265), .B(n49264), .ZN(
        n49269) );
  OR2_X1 U49885 ( .A1(n49267), .A2(n49266), .ZN(n49268) );
  OAI211_X1 U49886 ( .C1(n49271), .C2(n49270), .A(n49269), .B(n49268), .ZN(
        n49281) );
  AOI22_X1 U49887 ( .A1(n49275), .A2(n49274), .B1(n49273), .B2(n49272), .ZN(
        n49279) );
  AND2_X1 U49888 ( .A1(n49367), .A2(n523), .ZN(n49364) );
  INV_X1 U49889 ( .A(n49370), .ZN(n49378) );
  OR2_X1 U49890 ( .A1(n51729), .A2(n49366), .ZN(n49282) );
  AOI22_X1 U49891 ( .A1(n49284), .A2(n49364), .B1(n49378), .B2(n49283), .ZN(
        n49292) );
  OR2_X1 U49892 ( .A1(n49375), .A2(n522), .ZN(n49313) );
  INV_X1 U49893 ( .A(n49313), .ZN(n49332) );
  OAI211_X1 U49894 ( .C1(n49332), .C2(n49366), .A(n49376), .B(n49344), .ZN(
        n49291) );
  NAND2_X1 U49895 ( .A1(n49342), .A2(n49370), .ZN(n49286) );
  AOI21_X1 U49896 ( .B1(n49286), .B2(n49347), .A(n523), .ZN(n49287) );
  NAND2_X1 U49897 ( .A1(n49288), .A2(n49287), .ZN(n49290) );
  OR2_X1 U49898 ( .A1(n49313), .A2(n49380), .ZN(n49289) );
  INV_X1 U49899 ( .A(n4665), .ZN(n49293) );
  INV_X1 U49900 ( .A(n49366), .ZN(n49302) );
  NAND2_X1 U49901 ( .A1(n49302), .A2(n49347), .ZN(n49382) );
  OAI21_X1 U49902 ( .B1(n49382), .B2(n49313), .A(n49344), .ZN(n49294) );
  INV_X1 U49903 ( .A(n522), .ZN(n49377) );
  NAND2_X1 U49904 ( .A1(n8021), .A2(n49366), .ZN(n49296) );
  NAND2_X1 U49905 ( .A1(n8021), .A2(n51729), .ZN(n49295) );
  NAND4_X1 U49906 ( .A1(n49350), .A2(n49367), .A3(n49296), .A4(n49295), .ZN(
        n49300) );
  NAND4_X1 U49907 ( .A1(n49349), .A2(n49302), .A3(n49370), .A4(n49376), .ZN(
        n49299) );
  NAND2_X1 U49908 ( .A1(n49370), .A2(n49366), .ZN(n49372) );
  INV_X1 U49909 ( .A(n49372), .ZN(n49297) );
  OR2_X1 U49910 ( .A1(n522), .A2(n49376), .ZN(n49312) );
  NAND3_X1 U49911 ( .A1(n49297), .A2(n49367), .A3(n49312), .ZN(n49298) );
  NAND4_X1 U49912 ( .A1(n49301), .A2(n49300), .A3(n49299), .A4(n49298), .ZN(
        n49309) );
  OR2_X1 U49913 ( .A1(n49367), .A2(n49371), .ZN(n49319) );
  NOR2_X1 U49914 ( .A1(n49302), .A2(n49367), .ZN(n49351) );
  OAI21_X1 U49915 ( .B1(n49347), .B2(n49312), .A(n51729), .ZN(n49304) );
  AOI21_X1 U49916 ( .B1(n523), .B2(n49376), .A(n49370), .ZN(n49303) );
  OAI211_X1 U49917 ( .C1(n49351), .C2(n51729), .A(n49304), .B(n49303), .ZN(
        n49307) );
  AOI22_X1 U49918 ( .A1(n49305), .A2(n49347), .B1(n49342), .B2(n49376), .ZN(
        n49306) );
  OAI211_X1 U49919 ( .C1(n49372), .C2(n49319), .A(n49307), .B(n49306), .ZN(
        n49308) );
  INV_X1 U49920 ( .A(n4895), .ZN(n49310) );
  XNOR2_X1 U49921 ( .A(n49311), .B(n49310), .ZN(Plaintext[103]) );
  INV_X1 U49922 ( .A(n49380), .ZN(n49316) );
  INV_X1 U49923 ( .A(n49312), .ZN(n49315) );
  NAND2_X1 U49924 ( .A1(n49313), .A2(n49344), .ZN(n49314) );
  AOI22_X1 U49925 ( .A1(n49316), .A2(n49315), .B1(n49350), .B2(n49314), .ZN(
        n49321) );
  OAI21_X1 U49926 ( .B1(n49371), .B2(n49366), .A(n49367), .ZN(n49317) );
  NAND2_X1 U49927 ( .A1(n49350), .A2(n49317), .ZN(n49318) );
  AND2_X1 U49928 ( .A1(n49318), .A2(n49319), .ZN(n49320) );
  OAI211_X1 U49929 ( .C1(n49322), .C2(n523), .A(n49321), .B(n49320), .ZN(
        n49325) );
  INV_X1 U49930 ( .A(n49323), .ZN(n49324) );
  XNOR2_X1 U49931 ( .A(n49325), .B(n49324), .ZN(Plaintext[104]) );
  NAND2_X1 U49932 ( .A1(n49366), .A2(n49365), .ZN(n49358) );
  INV_X1 U49933 ( .A(n49358), .ZN(n49326) );
  NAND3_X1 U49934 ( .A1(n49326), .A2(n49371), .A3(n49347), .ZN(n49328) );
  AND2_X1 U49935 ( .A1(n49365), .A2(n51729), .ZN(n49346) );
  NAND3_X1 U49936 ( .A1(n49347), .A2(n49378), .A3(n49346), .ZN(n49327) );
  AND3_X1 U49937 ( .A1(n49329), .A2(n49328), .A3(n49327), .ZN(n49339) );
  NAND3_X1 U49938 ( .A1(n49349), .A2(n49347), .A3(n49350), .ZN(n49331) );
  NAND3_X1 U49939 ( .A1(n49350), .A2(n523), .A3(n49366), .ZN(n49330) );
  AND2_X1 U49940 ( .A1(n49331), .A2(n49330), .ZN(n49338) );
  INV_X1 U49941 ( .A(n49363), .ZN(n49334) );
  NOR2_X1 U49942 ( .A1(n49332), .A2(n49365), .ZN(n49333) );
  OAI211_X1 U49943 ( .C1(n49364), .C2(n49366), .A(n49334), .B(n49333), .ZN(
        n49337) );
  NAND2_X1 U49944 ( .A1(n49382), .A2(n49378), .ZN(n49335) );
  NAND3_X1 U49945 ( .A1(n49335), .A2(n49376), .A3(n8021), .ZN(n49336) );
  NAND4_X1 U49946 ( .A1(n49339), .A2(n49338), .A3(n49337), .A4(n49336), .ZN(
        n49341) );
  INV_X1 U49947 ( .A(n4868), .ZN(n49340) );
  XNOR2_X1 U49948 ( .A(n49341), .B(n49340), .ZN(Plaintext[105]) );
  NAND2_X1 U49949 ( .A1(n49342), .A2(n49367), .ZN(n49343) );
  AND2_X1 U49951 ( .A1(n49370), .A2(n51729), .ZN(n49359) );
  INV_X1 U49952 ( .A(n49349), .ZN(n49345) );
  OAI211_X1 U49953 ( .C1(n49365), .C2(n49359), .A(n49345), .B(n49382), .ZN(
        n49354) );
  INV_X1 U49954 ( .A(n49346), .ZN(n49348) );
  NAND4_X1 U49955 ( .A1(n49348), .A2(n49347), .A3(n49370), .A4(n8021), .ZN(
        n49353) );
  NAND3_X1 U49956 ( .A1(n49351), .A2(n49350), .A3(n49349), .ZN(n49352) );
  NAND4_X1 U49957 ( .A1(n51309), .A2(n49354), .A3(n49353), .A4(n49352), .ZN(
        n49357) );
  INV_X1 U49958 ( .A(n4585), .ZN(n49356) );
  XNOR2_X1 U49959 ( .A(n49357), .B(n49356), .ZN(Plaintext[106]) );
  NAND3_X1 U49960 ( .A1(n49360), .A2(n49359), .A3(n49358), .ZN(n49386) );
  OAI21_X1 U49961 ( .B1(n49366), .B2(n49376), .A(n49370), .ZN(n49361) );
  INV_X1 U49962 ( .A(n49361), .ZN(n49362) );
  AOI22_X1 U49963 ( .A1(n49365), .A2(n49364), .B1(n49363), .B2(n49362), .ZN(
        n49385) );
  XNOR2_X1 U49964 ( .A(n51729), .B(n49366), .ZN(n49368) );
  OAI21_X1 U49965 ( .B1(n49368), .B2(n523), .A(n49367), .ZN(n49374) );
  OAI21_X1 U49966 ( .B1(n49371), .B2(n49370), .A(n523), .ZN(n49373) );
  NAND4_X1 U49967 ( .A1(n49374), .A2(n49376), .A3(n49373), .A4(n49372), .ZN(
        n49384) );
  OAI21_X1 U49968 ( .B1(n49377), .B2(n49376), .A(n51729), .ZN(n49379) );
  NOR2_X1 U49969 ( .A1(n49379), .A2(n49378), .ZN(n49381) );
  NAND3_X1 U49970 ( .A1(n49382), .A2(n49381), .A3(n49380), .ZN(n49383) );
  NOR2_X1 U49971 ( .A1(n49445), .A2(n49442), .ZN(n49448) );
  AND2_X1 U49972 ( .A1(n51091), .A2(n49443), .ZN(n49389) );
  NOR2_X1 U49973 ( .A1(n49445), .A2(n49389), .ZN(n49392) );
  AOI22_X1 U49974 ( .A1(n49448), .A2(n49393), .B1(n49392), .B2(n49391), .ZN(
        n49413) );
  INV_X1 U49975 ( .A(n49394), .ZN(n49399) );
  INV_X1 U49976 ( .A(n49395), .ZN(n49396) );
  NOR2_X1 U49977 ( .A1(n49396), .A2(n49699), .ZN(n49398) );
  MUX2_X1 U49978 ( .A(n49399), .B(n49398), .S(n49397), .Z(n49402) );
  NAND2_X1 U49980 ( .A1(n49402), .A2(n52072), .ZN(n49406) );
  INV_X1 U49981 ( .A(n49403), .ZN(n49405) );
  AND2_X1 U49982 ( .A1(n52107), .A2(n49442), .ZN(n49436) );
  AOI22_X1 U49983 ( .A1(n49418), .A2(n52107), .B1(n49436), .B2(n49450), .ZN(
        n49404) );
  OAI211_X1 U49984 ( .C1(n49407), .C2(n49406), .A(n49405), .B(n49404), .ZN(
        n49412) );
  INV_X1 U49985 ( .A(n49452), .ZN(n49408) );
  AOI22_X1 U49986 ( .A1(n49408), .A2(n51316), .B1(n49459), .B2(n49458), .ZN(
        n49411) );
  NAND2_X1 U49987 ( .A1(n49409), .A2(n49462), .ZN(n49410) );
  NAND4_X1 U49988 ( .A1(n49413), .A2(n49412), .A3(n49411), .A4(n49410), .ZN(
        n49416) );
  INV_X1 U49989 ( .A(n49414), .ZN(n49415) );
  XNOR2_X1 U49990 ( .A(n49416), .B(n49415), .ZN(Plaintext[108]) );
  NAND2_X1 U49991 ( .A1(n49417), .A2(n49443), .ZN(n49428) );
  NAND2_X1 U49992 ( .A1(n51316), .A2(n49465), .ZN(n49419) );
  OAI22_X1 U49993 ( .A1(n49424), .A2(n49420), .B1(n49460), .B2(n49419), .ZN(
        n49421) );
  INV_X1 U49994 ( .A(n49421), .ZN(n49427) );
  INV_X1 U49995 ( .A(n49457), .ZN(n49449) );
  INV_X1 U49996 ( .A(n49458), .ZN(n49422) );
  NAND4_X1 U49997 ( .A1(n49428), .A2(n49427), .A3(n49426), .A4(n49425), .ZN(
        n49431) );
  INV_X1 U49998 ( .A(n49429), .ZN(n49430) );
  XNOR2_X1 U49999 ( .A(n49431), .B(n49430), .ZN(Plaintext[110]) );
  NAND2_X1 U50000 ( .A1(n49449), .A2(n49432), .ZN(n49433) );
  NAND3_X1 U50001 ( .A1(n49434), .A2(n49442), .A3(n49465), .ZN(n49439) );
  XNOR2_X1 U50002 ( .A(n49442), .B(n49465), .ZN(n49435) );
  NAND4_X1 U50004 ( .A1(n49445), .A2(n49436), .A3(n49450), .A4(n51315), .ZN(
        n49437) );
  NAND2_X1 U50005 ( .A1(n49443), .A2(n2858), .ZN(n49444) );
  NOR2_X1 U50006 ( .A1(n49445), .A2(n49444), .ZN(n49446) );
  AOI22_X1 U50007 ( .A1(n49448), .A2(n52107), .B1(n49446), .B2(n51316), .ZN(
        n49454) );
  NOR2_X1 U50008 ( .A1(n49452), .A2(n49451), .ZN(n49466) );
  INV_X1 U50009 ( .A(n49466), .ZN(n49453) );
  INV_X1 U50010 ( .A(n4316), .ZN(n49455) );
  INV_X1 U50011 ( .A(n49456), .ZN(n49470) );
  AOI22_X1 U50012 ( .A1(n49461), .A2(n49459), .B1(n49458), .B2(n51316), .ZN(
        n49469) );
  NAND2_X1 U50013 ( .A1(n49461), .A2(n49460), .ZN(n49464) );
  INV_X1 U50014 ( .A(n49462), .ZN(n49463) );
  NAND2_X1 U50015 ( .A1(n49464), .A2(n49463), .ZN(n49468) );
  NAND2_X1 U50016 ( .A1(n49466), .A2(n49465), .ZN(n49467) );
  NAND4_X1 U50017 ( .A1(n49470), .A2(n49469), .A3(n49468), .A4(n49467), .ZN(
        n49472) );
  INV_X1 U50018 ( .A(n4803), .ZN(n49471) );
  XNOR2_X1 U50019 ( .A(n49472), .B(n49471), .ZN(Plaintext[112]) );
  XNOR2_X1 U50020 ( .A(n49521), .B(n49534), .ZN(n49475) );
  NOR2_X1 U50021 ( .A1(n49534), .A2(n49521), .ZN(n49490) );
  NAND2_X1 U50022 ( .A1(n49490), .A2(n43490), .ZN(n49474) );
  NAND2_X1 U50023 ( .A1(n49510), .A2(n43490), .ZN(n49536) );
  NAND2_X1 U50024 ( .A1(n49514), .A2(n49503), .ZN(n49526) );
  AND3_X1 U50025 ( .A1(n49511), .A2(n49536), .A3(n49526), .ZN(n49473) );
  OAI211_X1 U50026 ( .C1(n49475), .C2(n2193), .A(n49474), .B(n49473), .ZN(
        n49484) );
  NAND3_X1 U50027 ( .A1(n49491), .A2(n2193), .A3(n49539), .ZN(n49478) );
  NAND4_X1 U50028 ( .A1(n49529), .A2(n49534), .A3(n49476), .A4(n49503), .ZN(
        n49477) );
  AND2_X1 U50029 ( .A1(n49478), .A2(n49477), .ZN(n49482) );
  NAND3_X1 U50030 ( .A1(n49480), .A2(n49479), .A3(n49503), .ZN(n49481) );
  NAND4_X1 U50031 ( .A1(n49484), .A2(n49483), .A3(n49482), .A4(n49481), .ZN(
        n49486) );
  INV_X1 U50032 ( .A(n3383), .ZN(n49485) );
  XNOR2_X1 U50033 ( .A(n49486), .B(n49485), .ZN(Plaintext[114]) );
  OR2_X1 U50034 ( .A1(n49534), .A2(n49522), .ZN(n49528) );
  INV_X1 U50035 ( .A(n49528), .ZN(n49489) );
  INV_X1 U50036 ( .A(n49487), .ZN(n49488) );
  NAND3_X1 U50037 ( .A1(n49489), .A2(n43490), .A3(n49488), .ZN(n49501) );
  INV_X1 U50038 ( .A(n49490), .ZN(n49500) );
  AND2_X1 U50039 ( .A1(n2193), .A2(n49503), .ZN(n49540) );
  NAND2_X1 U50040 ( .A1(n49493), .A2(n49540), .ZN(n49499) );
  NAND2_X1 U50041 ( .A1(n49494), .A2(n49512), .ZN(n49497) );
  INV_X1 U50042 ( .A(n49495), .ZN(n49496) );
  NAND2_X1 U50043 ( .A1(n49497), .A2(n49496), .ZN(n49498) );
  INV_X1 U50044 ( .A(n4817), .ZN(n49502) );
  OR2_X1 U50045 ( .A1(n2193), .A2(n49521), .ZN(n49537) );
  INV_X1 U50046 ( .A(n49537), .ZN(n49507) );
  AND2_X1 U50047 ( .A1(n49522), .A2(n49503), .ZN(n49504) );
  NAND4_X1 U50048 ( .A1(n49539), .A2(n49504), .A3(n49521), .A4(n2192), .ZN(
        n49505) );
  OAI21_X1 U50049 ( .B1(n49507), .B2(n49506), .A(n49505), .ZN(n49509) );
  NAND2_X1 U50050 ( .A1(n49509), .A2(n49508), .ZN(n49518) );
  INV_X1 U50051 ( .A(n49512), .ZN(n49531) );
  NAND2_X1 U50052 ( .A1(n43490), .A2(n2193), .ZN(n49524) );
  NAND3_X1 U50053 ( .A1(n49531), .A2(n49522), .A3(n49524), .ZN(n49516) );
  OAI211_X1 U50054 ( .C1(n49539), .C2(n51395), .A(n49534), .B(n49514), .ZN(
        n49515) );
  NAND4_X1 U50055 ( .A1(n49518), .A2(n49517), .A3(n49516), .A4(n49515), .ZN(
        n49520) );
  INV_X1 U50056 ( .A(n4204), .ZN(n49519) );
  XNOR2_X1 U50057 ( .A(n49520), .B(n49519), .ZN(Plaintext[118]) );
  OR2_X1 U50058 ( .A1(n49522), .A2(n49521), .ZN(n49523) );
  NOR2_X1 U50059 ( .A1(n49524), .A2(n49523), .ZN(n49525) );
  OR3_X1 U50060 ( .A1(n49534), .A2(n49510), .A3(n49526), .ZN(n49547) );
  NAND3_X1 U50061 ( .A1(n49528), .A2(n49510), .A3(n49539), .ZN(n49533) );
  NAND4_X1 U50063 ( .A1(n49537), .A2(n49536), .A3(n51395), .A4(n49534), .ZN(
        n49544) );
  INV_X1 U50064 ( .A(n49538), .ZN(n49541) );
  NAND3_X1 U50065 ( .A1(n49541), .A2(n49540), .A3(n49539), .ZN(n49542) );
  INV_X1 U50066 ( .A(n4879), .ZN(n49549) );
  NOR2_X1 U50067 ( .A1(n49580), .A2(n49608), .ZN(n49601) );
  INV_X1 U50068 ( .A(n49601), .ZN(n49552) );
  OAI211_X1 U50069 ( .C1(n49552), .C2(n49551), .A(n49583), .B(n49605), .ZN(
        n49553) );
  INV_X1 U50070 ( .A(n49606), .ZN(n49563) );
  NAND2_X1 U50071 ( .A1(n49553), .A2(n49563), .ZN(n49560) );
  NAND2_X1 U50072 ( .A1(n49573), .A2(n49599), .ZN(n49559) );
  INV_X1 U50073 ( .A(n49586), .ZN(n49568) );
  NAND3_X1 U50074 ( .A1(n49568), .A2(n49554), .A3(n51088), .ZN(n49558) );
  INV_X1 U50075 ( .A(n49607), .ZN(n49555) );
  OAI21_X1 U50076 ( .B1(n49556), .B2(n49593), .A(n49555), .ZN(n49557) );
  NAND4_X1 U50077 ( .A1(n49560), .A2(n49559), .A3(n49558), .A4(n49557), .ZN(
        n49561) );
  XNOR2_X1 U50078 ( .A(n49561), .B(n6926), .ZN(Plaintext[122]) );
  OAI211_X1 U50079 ( .C1(n49563), .C2(n49599), .A(n49584), .B(n49585), .ZN(
        n49567) );
  NAND2_X1 U50080 ( .A1(n49595), .A2(n49574), .ZN(n49566) );
  NAND2_X1 U50081 ( .A1(n49564), .A2(n49600), .ZN(n49565) );
  AND4_X1 U50082 ( .A1(n49567), .A2(n49602), .A3(n49566), .A4(n49565), .ZN(
        n49576) );
  OAI211_X1 U50083 ( .C1(n6985), .C2(n49580), .A(n49568), .B(n49598), .ZN(
        n49572) );
  NAND2_X1 U50084 ( .A1(n49580), .A2(n49606), .ZN(n49570) );
  OAI21_X1 U50085 ( .B1(n49604), .B2(n49570), .A(n49569), .ZN(n49571) );
  NAND2_X1 U50086 ( .A1(n49572), .A2(n49571), .ZN(n49575) );
  XNOR2_X1 U50087 ( .A(n49578), .B(n49577), .ZN(Plaintext[123]) );
  AND2_X1 U50088 ( .A1(n49580), .A2(n49579), .ZN(n49582) );
  AOI21_X1 U50089 ( .B1(n49583), .B2(n49580), .A(n49598), .ZN(n49581) );
  OAI21_X1 U50090 ( .B1(n49585), .B2(n49582), .A(n49581), .ZN(n49590) );
  NAND4_X1 U50091 ( .A1(n49584), .A2(n49600), .A3(n49583), .A4(n49608), .ZN(
        n49589) );
  NAND2_X1 U50092 ( .A1(n49593), .A2(n49585), .ZN(n49588) );
  NAND2_X1 U50093 ( .A1(n49586), .A2(n49606), .ZN(n49587) );
  XNOR2_X1 U50094 ( .A(n49591), .B(n4518), .ZN(Plaintext[124]) );
  INV_X1 U50095 ( .A(n49593), .ZN(n49594) );
  AOI21_X1 U50096 ( .B1(n647), .B2(n49595), .A(n49594), .ZN(n49596) );
  NAND3_X1 U50097 ( .A1(n49610), .A2(n49609), .A3(n49608), .ZN(n49611) );
  INV_X1 U50098 ( .A(n3481), .ZN(n49612) );
  OR2_X1 U50099 ( .A1(n50305), .A2(n49946), .ZN(n49955) );
  OAI21_X1 U50100 ( .B1(n49954), .B2(n49637), .A(n49613), .ZN(n49615) );
  NOR2_X1 U50101 ( .A1(n50297), .A2(n28), .ZN(n49948) );
  MUX2_X1 U50102 ( .A(n50297), .B(n49638), .S(n50287), .Z(n49617) );
  AOI21_X1 U50103 ( .B1(n28), .B2(n49617), .A(n49616), .ZN(n49752) );
  INV_X1 U50104 ( .A(n49618), .ZN(n49619) );
  NAND2_X1 U50105 ( .A1(n49619), .A2(n49627), .ZN(n49634) );
  NOR2_X1 U50106 ( .A1(n49978), .A2(n49980), .ZN(n49620) );
  AOI21_X1 U50107 ( .B1(n49620), .B2(n49627), .A(n49629), .ZN(n49621) );
  OAI21_X1 U50108 ( .B1(n49987), .B2(n49627), .A(n49621), .ZN(n49622) );
  NAND2_X1 U50109 ( .A1(n49622), .A2(n49990), .ZN(n49633) );
  NAND4_X1 U50110 ( .A1(n49626), .A2(n49625), .A3(n49624), .A4(n49623), .ZN(
        n49632) );
  NAND2_X1 U50111 ( .A1(n49980), .A2(n49627), .ZN(n49628) );
  OAI21_X1 U50112 ( .B1(n49979), .B2(n49628), .A(n49987), .ZN(n49630) );
  NAND2_X1 U50113 ( .A1(n49630), .A2(n49629), .ZN(n49631) );
  NOR2_X1 U50114 ( .A1(n49704), .A2(n49853), .ZN(n49644) );
  NAND2_X1 U50115 ( .A1(n49636), .A2(n51504), .ZN(n49942) );
  OR2_X1 U50116 ( .A1(n49638), .A2(n49637), .ZN(n50303) );
  OR2_X1 U50117 ( .A1(n49639), .A2(n49956), .ZN(n49640) );
  NAND3_X1 U50118 ( .A1(n49641), .A2(n50287), .A3(n49640), .ZN(n49642) );
  NAND2_X1 U50119 ( .A1(n49643), .A2(n49939), .ZN(n49762) );
  AND2_X1 U50120 ( .A1(n49810), .A2(n49762), .ZN(n49706) );
  INV_X1 U50121 ( .A(n49823), .ZN(n49848) );
  INV_X1 U50122 ( .A(n49645), .ZN(n49649) );
  NAND2_X1 U50123 ( .A1(n49647), .A2(n49646), .ZN(n49648) );
  NAND2_X1 U50124 ( .A1(n49652), .A2(n49651), .ZN(n49653) );
  OR2_X1 U50125 ( .A1(n49654), .A2(n49653), .ZN(n50022) );
  INV_X1 U50126 ( .A(n49671), .ZN(n50028) );
  NAND3_X1 U50127 ( .A1(n50022), .A2(n49655), .A3(n50028), .ZN(n49682) );
  NAND4_X1 U50128 ( .A1(n49660), .A2(n49677), .A3(n49659), .A4(n49658), .ZN(
        n49680) );
  NAND2_X1 U50129 ( .A1(n49669), .A2(n49661), .ZN(n49665) );
  NAND3_X1 U50130 ( .A1(n50027), .A2(n49663), .A3(n51733), .ZN(n49664) );
  NAND2_X1 U50131 ( .A1(n49646), .A2(n49667), .ZN(n49668) );
  NAND2_X1 U50132 ( .A1(n49671), .A2(n52212), .ZN(n49675) );
  NAND2_X1 U50133 ( .A1(n49673), .A2(n49672), .ZN(n49674) );
  NAND4_X1 U50134 ( .A1(n49677), .A2(n49676), .A3(n49675), .A4(n49674), .ZN(
        n49678) );
  OAI21_X1 U50135 ( .B1(n49680), .B2(n49679), .A(n49678), .ZN(n49681) );
  INV_X1 U50136 ( .A(n49683), .ZN(n49687) );
  NOR2_X1 U50137 ( .A1(n49684), .A2(n51095), .ZN(n49685) );
  AOI22_X1 U50138 ( .A1(n49687), .A2(n49686), .B1(n49248), .B2(n49685), .ZN(
        n49702) );
  OAI21_X1 U50139 ( .B1(n49690), .B2(n49689), .A(n49688), .ZN(n49693) );
  AOI22_X1 U50140 ( .A1(n49694), .A2(n49693), .B1(n656), .B2(n49692), .ZN(
        n49701) );
  NOR2_X1 U50141 ( .A1(n49696), .A2(n51095), .ZN(n49698) );
  OAI21_X1 U50142 ( .B1(n49699), .B2(n49698), .A(n51731), .ZN(n49700) );
  OR2_X1 U50144 ( .A1(n49850), .A2(n49871), .ZN(n49774) );
  NOR2_X1 U50145 ( .A1(n49848), .A2(n49774), .ZN(n49751) );
  NOR2_X1 U50146 ( .A1(n49710), .A2(n49707), .ZN(n49709) );
  OAI21_X1 U50147 ( .B1(n49709), .B2(n49725), .A(n49708), .ZN(n49716) );
  NOR2_X1 U50148 ( .A1(n49725), .A2(n49710), .ZN(n49712) );
  AOI22_X1 U50149 ( .A1(n49721), .A2(n49713), .B1(n49712), .B2(n49711), .ZN(
        n49715) );
  MUX2_X1 U50150 ( .A(n49716), .B(n49715), .S(n49714), .Z(n49771) );
  OR2_X1 U50151 ( .A1(n49718), .A2(n49717), .ZN(n49728) );
  OR2_X1 U50152 ( .A1(n51295), .A2(n49719), .ZN(n49724) );
  NAND2_X1 U50153 ( .A1(n49722), .A2(n49721), .ZN(n49723) );
  NAND4_X1 U50154 ( .A1(n49726), .A2(n49725), .A3(n49724), .A4(n49723), .ZN(
        n49727) );
  AND2_X1 U50155 ( .A1(n49728), .A2(n49727), .ZN(n49770) );
  OR2_X1 U50156 ( .A1(n49841), .A2(n49782), .ZN(n49856) );
  NAND3_X1 U50157 ( .A1(n49850), .A2(n49871), .A3(n49853), .ZN(n49779) );
  NAND2_X1 U50158 ( .A1(n50377), .A2(n2198), .ZN(n49735) );
  NAND2_X1 U50159 ( .A1(n2198), .A2(n50034), .ZN(n49729) );
  OAI211_X1 U50160 ( .C1(n49732), .C2(n49731), .A(n49730), .B(n49729), .ZN(
        n49733) );
  OAI211_X1 U50161 ( .C1(n49736), .C2(n49735), .A(n49734), .B(n49733), .ZN(
        n49737) );
  INV_X1 U50162 ( .A(n49737), .ZN(n49748) );
  OAI211_X1 U50165 ( .C1(n50378), .C2(n49743), .A(n49742), .B(n50387), .ZN(
        n49745) );
  NAND3_X1 U50166 ( .A1(n49820), .A2(n49863), .A3(n49853), .ZN(n49749) );
  OAI21_X1 U50167 ( .B1(n49856), .B2(n49779), .A(n49749), .ZN(n49750) );
  NOR2_X1 U50168 ( .A1(n49751), .A2(n49750), .ZN(n49759) );
  NAND2_X1 U50169 ( .A1(n49829), .A2(n49841), .ZN(n49758) );
  INV_X1 U50170 ( .A(n49819), .ZN(n49796) );
  NAND4_X1 U50171 ( .A1(n49793), .A2(n49796), .A3(n49862), .A4(n49841), .ZN(
        n49757) );
  NAND2_X1 U50172 ( .A1(n49766), .A2(n49854), .ZN(n49826) );
  INV_X1 U50173 ( .A(n49826), .ZN(n49825) );
  NAND2_X1 U50174 ( .A1(n49850), .A2(n49782), .ZN(n49777) );
  INV_X1 U50175 ( .A(n49752), .ZN(n49764) );
  NAND2_X1 U50176 ( .A1(n49762), .A2(n49764), .ZN(n49808) );
  OR2_X1 U50177 ( .A1(n49808), .A2(n49809), .ZN(n49805) );
  INV_X1 U50178 ( .A(n49810), .ZN(n49753) );
  NAND2_X1 U50180 ( .A1(n49862), .A2(n49863), .ZN(n49851) );
  NAND2_X1 U50181 ( .A1(n51314), .A2(n49851), .ZN(n49755) );
  NAND2_X1 U50182 ( .A1(n49862), .A2(n49871), .ZN(n49754) );
  OAI211_X1 U50183 ( .C1(n49825), .C2(n49777), .A(n49755), .B(n49754), .ZN(
        n49756) );
  NAND4_X1 U50184 ( .A1(n49759), .A2(n49758), .A3(n49757), .A4(n49756), .ZN(
        n49761) );
  INV_X1 U50185 ( .A(n4705), .ZN(n49760) );
  XNOR2_X1 U50186 ( .A(n49761), .B(n49760), .ZN(Plaintext[126]) );
  INV_X1 U50187 ( .A(n49762), .ZN(n49763) );
  NOR2_X1 U50188 ( .A1(n49763), .A2(n49809), .ZN(n49765) );
  NAND4_X1 U50189 ( .A1(n49765), .A2(n49854), .A3(n49764), .A4(n49810), .ZN(
        n49767) );
  INV_X1 U50190 ( .A(n49766), .ZN(n49839) );
  NAND2_X1 U50191 ( .A1(n49767), .A2(n49839), .ZN(n49768) );
  NAND3_X1 U50192 ( .A1(n49768), .A2(n49853), .A3(n49826), .ZN(n49803) );
  NAND3_X1 U50193 ( .A1(n49823), .A2(n49839), .A3(n49862), .ZN(n49769) );
  MUX2_X1 U50194 ( .A(n49803), .B(n49769), .S(n49819), .Z(n49789) );
  INV_X1 U50195 ( .A(n49853), .ZN(n49811) );
  AND2_X1 U50196 ( .A1(n49811), .A2(n49863), .ZN(n49836) );
  INV_X1 U50198 ( .A(n49850), .ZN(n49837) );
  NAND4_X1 U50199 ( .A1(n49841), .A2(n49837), .A3(n49871), .A4(n49784), .ZN(
        n49773) );
  NAND4_X1 U50200 ( .A1(n49841), .A2(n49782), .A3(n49837), .A4(n49863), .ZN(
        n49772) );
  OAI211_X1 U50201 ( .C1(n49775), .C2(n49774), .A(n49773), .B(n49772), .ZN(
        n49776) );
  INV_X1 U50202 ( .A(n49776), .ZN(n49788) );
  OAI21_X1 U50203 ( .B1(n49777), .B2(n49863), .A(n49841), .ZN(n49781) );
  NOR2_X1 U50204 ( .A1(n49871), .A2(n49811), .ZN(n49847) );
  NAND3_X1 U50205 ( .A1(n49837), .A2(n49847), .A3(n49862), .ZN(n49778) );
  NAND3_X1 U50206 ( .A1(n49779), .A2(n49778), .A3(n49820), .ZN(n49780) );
  NAND2_X1 U50207 ( .A1(n49781), .A2(n49780), .ZN(n49787) );
  INV_X1 U50208 ( .A(n49836), .ZN(n49783) );
  NAND2_X1 U50209 ( .A1(n49782), .A2(n49839), .ZN(n49794) );
  OAI21_X1 U50210 ( .B1(n49783), .B2(n49794), .A(n51314), .ZN(n49785) );
  NAND3_X1 U50211 ( .A1(n49785), .A2(n49850), .A3(n49842), .ZN(n49786) );
  NAND4_X1 U50212 ( .A1(n49789), .A2(n49788), .A3(n49787), .A4(n49786), .ZN(
        n49792) );
  INV_X1 U50213 ( .A(n49790), .ZN(n49791) );
  XNOR2_X1 U50214 ( .A(n49792), .B(n49791), .ZN(Plaintext[127]) );
  NOR2_X1 U50215 ( .A1(n49841), .A2(n49839), .ZN(n49843) );
  OAI21_X1 U50216 ( .B1(n49844), .B2(n49843), .A(n49816), .ZN(n49800) );
  NOR2_X1 U50217 ( .A1(n51314), .A2(n49839), .ZN(n49824) );
  AND2_X1 U50218 ( .A1(n49823), .A2(n49862), .ZN(n49797) );
  NAND2_X1 U50219 ( .A1(n49850), .A2(n49871), .ZN(n49822) );
  NAND2_X1 U50220 ( .A1(n51314), .A2(n49822), .ZN(n49795) );
  AOI22_X1 U50221 ( .A1(n49797), .A2(n49796), .B1(n49795), .B2(n49784), .ZN(
        n49799) );
  NAND2_X1 U50222 ( .A1(n49829), .A2(n49871), .ZN(n49798) );
  OAI211_X1 U50223 ( .C1(n49800), .C2(n49824), .A(n49799), .B(n49798), .ZN(
        n49802) );
  INV_X1 U50224 ( .A(n3276), .ZN(n49801) );
  XNOR2_X1 U50225 ( .A(n49802), .B(n49801), .ZN(Plaintext[128]) );
  OAI21_X1 U50226 ( .B1(n49841), .B2(n49871), .A(n49811), .ZN(n49804) );
  INV_X1 U50227 ( .A(n49805), .ZN(n49806) );
  NAND4_X1 U50228 ( .A1(n49806), .A2(n49811), .A3(n49782), .A4(n49810), .ZN(
        n49807) );
  INV_X1 U50229 ( .A(n49808), .ZN(n49813) );
  INV_X1 U50230 ( .A(n49809), .ZN(n49812) );
  NAND4_X1 U50231 ( .A1(n49813), .A2(n49812), .A3(n49811), .A4(n49810), .ZN(
        n49814) );
  NAND3_X1 U50232 ( .A1(n49837), .A2(n49862), .A3(n49814), .ZN(n49815) );
  XNOR2_X1 U50233 ( .A(n49818), .B(n49817), .ZN(Plaintext[129]) );
  OAI21_X1 U50234 ( .B1(n49823), .B2(n49822), .A(n49821), .ZN(n49861) );
  NOR2_X1 U50235 ( .A1(n49861), .A2(n49824), .ZN(n49833) );
  OAI21_X1 U50236 ( .B1(n49784), .B2(n49825), .A(n49848), .ZN(n49832) );
  INV_X1 U50237 ( .A(n49856), .ZN(n49827) );
  NAND3_X1 U50238 ( .A1(n49827), .A2(n49826), .A3(n49850), .ZN(n49831) );
  NAND3_X1 U50239 ( .A1(n49829), .A2(n49847), .A3(n49828), .ZN(n49830) );
  NAND4_X1 U50240 ( .A1(n49833), .A2(n49832), .A3(n49831), .A4(n49830), .ZN(
        n49835) );
  INV_X1 U50241 ( .A(n4733), .ZN(n49834) );
  XNOR2_X1 U50242 ( .A(n49835), .B(n49834), .ZN(Plaintext[130]) );
  AND2_X1 U50243 ( .A1(n49836), .A2(n49862), .ZN(n49868) );
  NOR2_X1 U50244 ( .A1(n51314), .A2(n49837), .ZN(n49872) );
  MUX2_X1 U50245 ( .A(n49868), .B(n49872), .S(n49839), .Z(n49840) );
  INV_X1 U50246 ( .A(n49840), .ZN(n49859) );
  NAND2_X1 U50247 ( .A1(n49842), .A2(n49841), .ZN(n49846) );
  INV_X1 U50248 ( .A(n49843), .ZN(n49845) );
  INV_X1 U50249 ( .A(n49847), .ZN(n49849) );
  OAI21_X1 U50250 ( .B1(n49850), .B2(n49849), .A(n49848), .ZN(n49864) );
  INV_X1 U50251 ( .A(n49851), .ZN(n49852) );
  AOI21_X1 U50252 ( .B1(n49864), .B2(n49852), .A(n49867), .ZN(n49858) );
  AND2_X1 U50253 ( .A1(n49854), .A2(n49853), .ZN(n49855) );
  NAND2_X1 U50254 ( .A1(n49856), .A2(n49855), .ZN(n49860) );
  NAND2_X1 U50255 ( .A1(n49861), .A2(n49860), .ZN(n49857) );
  NAND3_X1 U50256 ( .A1(n49861), .A2(n49867), .A3(n49860), .ZN(n49866) );
  NAND4_X1 U50257 ( .A1(n49864), .A2(n49867), .A3(n49863), .A4(n49862), .ZN(
        n49865) );
  AND2_X1 U50258 ( .A1(n49866), .A2(n49865), .ZN(n49875) );
  INV_X1 U50259 ( .A(n49868), .ZN(n49869) );
  AOI21_X1 U50260 ( .B1(n49869), .B2(n49871), .A(n1354), .ZN(n49870) );
  OAI21_X1 U50261 ( .B1(n49872), .B2(n49871), .A(n49870), .ZN(n49873) );
  NAND4_X1 U50262 ( .A1(n49876), .A2(n49875), .A3(n49874), .A4(n49873), .ZN(
        Plaintext[131]) );
  MUX2_X1 U50263 ( .A(n49877), .B(n49907), .S(n49894), .Z(n49886) );
  AOI21_X1 U50264 ( .B1(n49919), .B2(n49899), .A(n49894), .ZN(n49879) );
  OAI22_X1 U50265 ( .A1(n49880), .A2(n49879), .B1(n49923), .B2(n49905), .ZN(
        n49881) );
  OAI21_X1 U50266 ( .B1(n49903), .B2(n49916), .A(n49881), .ZN(n49885) );
  OAI21_X1 U50267 ( .B1(n49882), .B2(n47420), .A(n49923), .ZN(n49883) );
  OAI211_X1 U50268 ( .C1(n49892), .C2(n49925), .A(n49883), .B(n49899), .ZN(
        n49884) );
  OAI211_X1 U50269 ( .C1(n49886), .C2(n49889), .A(n49885), .B(n49884), .ZN(
        n49888) );
  XNOR2_X1 U50270 ( .A(n49888), .B(n49887), .ZN(Plaintext[132]) );
  AND2_X1 U50271 ( .A1(n49923), .A2(n49889), .ZN(n49906) );
  AND2_X1 U50272 ( .A1(n49916), .A2(n49894), .ZN(n49902) );
  OAI21_X1 U50273 ( .B1(n49919), .B2(n49902), .A(n49891), .ZN(n49897) );
  OR2_X1 U50274 ( .A1(n652), .A2(n49916), .ZN(n49927) );
  NAND2_X1 U50275 ( .A1(n49899), .A2(n49892), .ZN(n49893) );
  NAND3_X1 U50276 ( .A1(n49927), .A2(n49894), .A3(n49893), .ZN(n49895) );
  NAND2_X1 U50277 ( .A1(n49934), .A2(n49895), .ZN(n49896) );
  INV_X1 U50278 ( .A(n4932), .ZN(n49898) );
  NAND2_X1 U50279 ( .A1(n49899), .A2(n49933), .ZN(n49915) );
  OR2_X1 U50280 ( .A1(n49900), .A2(n49915), .ZN(n49913) );
  NOR2_X1 U50281 ( .A1(n49901), .A2(n47420), .ZN(n49904) );
  AOI22_X1 U50282 ( .A1(n49904), .A2(n49903), .B1(n49902), .B2(n49932), .ZN(
        n49912) );
  NAND2_X1 U50283 ( .A1(n49906), .A2(n49905), .ZN(n49918) );
  NAND3_X1 U50284 ( .A1(n49909), .A2(n49908), .A3(n49907), .ZN(n49910) );
  NAND2_X1 U50285 ( .A1(n49910), .A2(n49928), .ZN(n49911) );
  NAND4_X1 U50286 ( .A1(n49913), .A2(n49912), .A3(n49918), .A4(n49911), .ZN(
        n49914) );
  XNOR2_X1 U50287 ( .A(n49914), .B(n6311), .ZN(Plaintext[136]) );
  NAND2_X1 U50290 ( .A1(n49918), .A2(n49917), .ZN(n49920) );
  NAND3_X1 U50291 ( .A1(n49929), .A2(n49928), .A3(n49927), .ZN(n49931) );
  NAND2_X1 U50292 ( .A1(n49931), .A2(n49930), .ZN(n49936) );
  NAND3_X1 U50293 ( .A1(n49934), .A2(n49933), .A3(n49932), .ZN(n49935) );
  INV_X1 U50294 ( .A(n49937), .ZN(n49938) );
  AOI22_X1 U50295 ( .A1(n50307), .A2(n49940), .B1(n49939), .B2(n50296), .ZN(
        n49941) );
  NAND2_X1 U50296 ( .A1(n49942), .A2(n49941), .ZN(n49944) );
  NAND3_X1 U50297 ( .A1(n49944), .A2(n28), .A3(n50309), .ZN(n49951) );
  OAI21_X1 U50298 ( .B1(n49946), .B2(n49945), .A(n50303), .ZN(n49947) );
  INV_X1 U50299 ( .A(n49947), .ZN(n49950) );
  NAND2_X1 U50300 ( .A1(n49948), .A2(n50307), .ZN(n49949) );
  NAND3_X1 U50301 ( .A1(n49951), .A2(n49950), .A3(n49949), .ZN(n49960) );
  NAND2_X1 U50302 ( .A1(n50287), .A2(n51300), .ZN(n49952) );
  OR2_X1 U50303 ( .A1(n49956), .A2(n49952), .ZN(n50304) );
  OAI21_X1 U50304 ( .B1(n49953), .B2(n7724), .A(n50304), .ZN(n49958) );
  AOI21_X1 U50305 ( .B1(n49956), .B2(n49955), .A(n49954), .ZN(n49957) );
  MUX2_X1 U50306 ( .A(n49958), .B(n49957), .S(n51691), .Z(n49959) );
  INV_X1 U50308 ( .A(n50337), .ZN(n49964) );
  OAI21_X1 U50309 ( .B1(n49964), .B2(n49963), .A(n49962), .ZN(n49966) );
  AOI21_X1 U50310 ( .B1(n50349), .B2(n52062), .A(n51725), .ZN(n49968) );
  NAND2_X1 U50311 ( .A1(n50144), .A2(n50115), .ZN(n50082) );
  NAND2_X1 U50312 ( .A1(n49989), .A2(n51326), .ZN(n49975) );
  NAND2_X1 U50313 ( .A1(n49979), .A2(n49983), .ZN(n49981) );
  OAI211_X1 U50314 ( .C1(n49983), .C2(n49982), .A(n49981), .B(n49980), .ZN(
        n49985) );
  NAND2_X1 U50315 ( .A1(n49985), .A2(n49984), .ZN(n49986) );
  OAI211_X1 U50316 ( .C1(n49990), .C2(n49989), .A(n49988), .B(n49987), .ZN(
        n49991) );
  OR2_X1 U50317 ( .A1(n50082), .A2(n51645), .ZN(n50102) );
  NAND2_X1 U50318 ( .A1(n50331), .A2(n50322), .ZN(n49992) );
  NAND3_X1 U50319 ( .A1(n49992), .A2(n52124), .A3(n50325), .ZN(n50000) );
  NAND3_X1 U50320 ( .A1(n49994), .A2(n49993), .A3(n50322), .ZN(n49999) );
  NOR2_X1 U50321 ( .A1(n49995), .A2(n50315), .ZN(n49997) );
  OAI21_X1 U50322 ( .B1(n49997), .B2(n50325), .A(n49996), .ZN(n49998) );
  AND3_X1 U50323 ( .A1(n50000), .A2(n49999), .A3(n49998), .ZN(n50018) );
  OR2_X1 U50324 ( .A1(n50322), .A2(n50001), .ZN(n50002) );
  NAND2_X1 U50325 ( .A1(n50003), .A2(n50002), .ZN(n50005) );
  NAND2_X1 U50326 ( .A1(n50005), .A2(n43577), .ZN(n50017) );
  NAND2_X1 U50327 ( .A1(n50007), .A2(n50006), .ZN(n50011) );
  NOR2_X1 U50328 ( .A1(n50316), .A2(n50008), .ZN(n50324) );
  INV_X1 U50329 ( .A(n50316), .ZN(n50012) );
  NAND2_X1 U50330 ( .A1(n50012), .A2(n50322), .ZN(n50014) );
  NAND4_X1 U50331 ( .A1(n50328), .A2(n50014), .A3(n1812), .A4(n50013), .ZN(
        n50016) );
  OR2_X1 U50332 ( .A1(n50020), .A2(n50019), .ZN(n50024) );
  INV_X1 U50333 ( .A(n50021), .ZN(n50023) );
  OAI21_X1 U50334 ( .B1(n50024), .B2(n50023), .A(n50022), .ZN(n50026) );
  NOR2_X1 U50335 ( .A1(n50026), .A2(n50025), .ZN(n50032) );
  NOR2_X1 U50336 ( .A1(n50030), .A2(n50029), .ZN(n50031) );
  NAND2_X1 U50337 ( .A1(n50378), .A2(n51058), .ZN(n50037) );
  NAND2_X1 U50338 ( .A1(n50033), .A2(n50377), .ZN(n50380) );
  INV_X1 U50339 ( .A(n50380), .ZN(n50036) );
  AOI22_X1 U50340 ( .A1(n50037), .A2(n50036), .B1(n50035), .B2(n50034), .ZN(
        n50038) );
  NAND2_X1 U50342 ( .A1(n50378), .A2(n50377), .ZN(n50040) );
  NAND2_X1 U50343 ( .A1(n50040), .A2(n2199), .ZN(n50043) );
  NAND2_X1 U50344 ( .A1(n50386), .A2(n50390), .ZN(n50041) );
  OR2_X1 U50345 ( .A1(n50378), .A2(n50041), .ZN(n50042) );
  OAI211_X1 U50346 ( .C1(n50044), .C2(n50375), .A(n50043), .B(n50042), .ZN(
        n50045) );
  AND2_X1 U50347 ( .A1(n51644), .A2(n562), .ZN(n50148) );
  NAND2_X1 U50348 ( .A1(n50148), .A2(n50145), .ZN(n50047) );
  INV_X1 U50349 ( .A(n50048), .ZN(n50055) );
  OR2_X1 U50350 ( .A1(n52055), .A2(n51727), .ZN(n50059) );
  NOR2_X1 U50351 ( .A1(n50079), .A2(n50059), .ZN(n50066) );
  NAND3_X1 U50353 ( .A1(n4203), .A2(n8603), .A3(n562), .ZN(n50138) );
  OAI21_X1 U50354 ( .B1(n50068), .B2(n51442), .A(n50138), .ZN(n50049) );
  OAI21_X1 U50355 ( .B1(n50066), .B2(n50049), .A(n51644), .ZN(n50054) );
  NAND2_X1 U50356 ( .A1(n50143), .A2(n50097), .ZN(n50087) );
  OAI21_X1 U50357 ( .B1(n50064), .B2(n50097), .A(n50087), .ZN(n50051) );
  NOR2_X1 U50358 ( .A1(n50088), .A2(n51442), .ZN(n50050) );
  OAI21_X1 U50359 ( .B1(n50051), .B2(n50050), .A(n52055), .ZN(n50053) );
  NOR2_X1 U50360 ( .A1(n50062), .A2(n50128), .ZN(n50135) );
  NAND2_X1 U50361 ( .A1(n50135), .A2(n50113), .ZN(n50052) );
  NAND4_X1 U50362 ( .A1(n50055), .A2(n50054), .A3(n50053), .A4(n50052), .ZN(
        n50057) );
  XNOR2_X1 U50363 ( .A(n50057), .B(n50056), .ZN(Plaintext[138]) );
  NAND2_X1 U50364 ( .A1(n50082), .A2(n50097), .ZN(n50058) );
  NAND2_X1 U50365 ( .A1(n50058), .A2(n50114), .ZN(n50061) );
  AND2_X1 U50366 ( .A1(n50145), .A2(n51442), .ZN(n50120) );
  NAND2_X1 U50367 ( .A1(n50113), .A2(n562), .ZN(n50060) );
  INV_X1 U50368 ( .A(n50059), .ZN(n50136) );
  OR2_X1 U50369 ( .A1(n50145), .A2(n50144), .ZN(n50129) );
  NOR2_X1 U50370 ( .A1(n50129), .A2(n50062), .ZN(n50134) );
  NOR2_X1 U50371 ( .A1(n50134), .A2(n50063), .ZN(n50075) );
  NAND2_X1 U50372 ( .A1(n4203), .A2(n51442), .ZN(n50065) );
  NOR3_X1 U50373 ( .A1(n50065), .A2(n50064), .A3(n50088), .ZN(n50067) );
  NOR2_X1 U50374 ( .A1(n50067), .A2(n50066), .ZN(n50074) );
  NAND2_X1 U50375 ( .A1(n50068), .A2(n51442), .ZN(n50072) );
  NOR2_X1 U50376 ( .A1(n50098), .A2(n4203), .ZN(n50071) );
  OAI211_X1 U50377 ( .C1(n50101), .C2(n50143), .A(n50097), .B(n50145), .ZN(
        n50070) );
  NAND4_X1 U50378 ( .A1(n50072), .A2(n50071), .A3(n50070), .A4(n50069), .ZN(
        n50073) );
  NAND4_X1 U50379 ( .A1(n50076), .A2(n50075), .A3(n50074), .A4(n50073), .ZN(
        n50078) );
  XNOR2_X1 U50380 ( .A(n50078), .B(n50077), .ZN(Plaintext[139]) );
  NOR2_X1 U50381 ( .A1(n50113), .A2(n50101), .ZN(n50081) );
  AND2_X1 U50382 ( .A1(n52055), .A2(n51645), .ZN(n50086) );
  INV_X1 U50383 ( .A(n50079), .ZN(n50080) );
  AOI21_X1 U50384 ( .B1(n50081), .B2(n50086), .A(n50080), .ZN(n50094) );
  INV_X1 U50385 ( .A(n50082), .ZN(n50085) );
  NAND2_X1 U50386 ( .A1(n50083), .A2(n50097), .ZN(n50084) );
  NAND2_X1 U50387 ( .A1(n50085), .A2(n50084), .ZN(n50093) );
  OAI21_X1 U50390 ( .B1(n50148), .B2(n50086), .A(n52078), .ZN(n50092) );
  NAND2_X1 U50391 ( .A1(n50129), .A2(n50087), .ZN(n50090) );
  INV_X1 U50392 ( .A(n50088), .ZN(n50089) );
  NAND2_X1 U50393 ( .A1(n50090), .A2(n50089), .ZN(n50091) );
  NAND4_X1 U50394 ( .A1(n50094), .A2(n50093), .A3(n50092), .A4(n50091), .ZN(
        n50096) );
  INV_X1 U50395 ( .A(n4568), .ZN(n50095) );
  XNOR2_X1 U50396 ( .A(n50096), .B(n50095), .ZN(Plaintext[140]) );
  NAND3_X1 U50397 ( .A1(n4203), .A2(n50114), .A3(n50101), .ZN(n50116) );
  NOR2_X1 U50398 ( .A1(n50145), .A2(n562), .ZN(n50111) );
  AND2_X1 U50399 ( .A1(n51442), .A2(n52055), .ZN(n50141) );
  NAND2_X1 U50400 ( .A1(n50111), .A2(n50141), .ZN(n50099) );
  INV_X1 U50401 ( .A(n50100), .ZN(n50106) );
  AND2_X1 U50402 ( .A1(n50101), .A2(n50143), .ZN(n50131) );
  AOI22_X1 U50403 ( .A1(n50120), .A2(n50131), .B1(n52078), .B2(n50148), .ZN(
        n50105) );
  NOR2_X1 U50404 ( .A1(n50145), .A2(n50101), .ZN(n50140) );
  AOI22_X1 U50405 ( .A1(n50140), .A2(n50143), .B1(n50148), .B2(n4203), .ZN(
        n50104) );
  INV_X1 U50406 ( .A(n50102), .ZN(n50121) );
  OAI21_X1 U50407 ( .B1(n50120), .B2(n50143), .A(n50121), .ZN(n50103) );
  INV_X1 U50409 ( .A(n4793), .ZN(n50107) );
  NAND2_X1 U50411 ( .A1(n4203), .A2(n51644), .ZN(n50110) );
  OAI21_X1 U50412 ( .B1(n50111), .B2(n50110), .A(n50128), .ZN(n50112) );
  OAI21_X1 U50413 ( .B1(n51442), .B2(n50113), .A(n50112), .ZN(n50124) );
  AOI22_X1 U50414 ( .A1(n50129), .A2(n562), .B1(n50114), .B2(n50145), .ZN(
        n50119) );
  NAND2_X1 U50415 ( .A1(n52078), .A2(n50116), .ZN(n50118) );
  NAND2_X1 U50416 ( .A1(n50119), .A2(n50118), .ZN(n50123) );
  NAND3_X1 U50417 ( .A1(n50121), .A2(n50120), .A3(n50143), .ZN(n50122) );
  NAND3_X1 U50418 ( .A1(n50124), .A2(n50123), .A3(n50122), .ZN(n50126) );
  INV_X1 U50419 ( .A(n4486), .ZN(n50125) );
  XNOR2_X1 U50420 ( .A(n50126), .B(n50125), .ZN(Plaintext[142]) );
  NAND2_X1 U50421 ( .A1(n51442), .A2(n51645), .ZN(n50130) );
  AOI21_X1 U50422 ( .B1(n50131), .B2(n50130), .A(n50129), .ZN(n50132) );
  OAI21_X1 U50423 ( .B1(n50134), .B2(n50133), .A(n50132), .ZN(n50153) );
  INV_X1 U50424 ( .A(n50142), .ZN(n50137) );
  AOI21_X1 U50425 ( .B1(n50137), .B2(n50136), .A(n50135), .ZN(n50152) );
  INV_X1 U50426 ( .A(n50138), .ZN(n50139) );
  AOI21_X1 U50427 ( .B1(n50141), .B2(n50140), .A(n50139), .ZN(n50151) );
  NAND2_X1 U50428 ( .A1(n50142), .A2(n52077), .ZN(n50147) );
  NAND3_X1 U50429 ( .A1(n50145), .A2(n52055), .A3(n50143), .ZN(n50146) );
  NAND2_X1 U50430 ( .A1(n50147), .A2(n50146), .ZN(n50149) );
  NAND2_X1 U50431 ( .A1(n50149), .A2(n50148), .ZN(n50150) );
  NAND4_X1 U50432 ( .A1(n50153), .A2(n50152), .A3(n50151), .A4(n50150), .ZN(
        n50155) );
  INV_X1 U50433 ( .A(n4286), .ZN(n50154) );
  XNOR2_X1 U50434 ( .A(n50155), .B(n50154), .ZN(Plaintext[143]) );
  NAND4_X1 U50435 ( .A1(n50178), .A2(n50226), .A3(n51480), .A4(n50196), .ZN(
        n50156) );
  AND2_X1 U50436 ( .A1(n50157), .A2(n50156), .ZN(n50172) );
  NOR2_X1 U50437 ( .A1(n50198), .A2(n50222), .ZN(n50214) );
  NOR2_X1 U50438 ( .A1(n51480), .A2(n50192), .ZN(n50199) );
  NAND2_X1 U50439 ( .A1(n50226), .A2(n50196), .ZN(n50213) );
  NOR2_X1 U50440 ( .A1(n50235), .A2(n50196), .ZN(n50188) );
  NOR2_X1 U50441 ( .A1(n50192), .A2(n50222), .ZN(n50158) );
  AOI21_X1 U50442 ( .B1(n50198), .B2(n50158), .A(n50187), .ZN(n50164) );
  NAND3_X1 U50443 ( .A1(n7201), .A2(n51480), .A3(n50233), .ZN(n50160) );
  NAND2_X1 U50444 ( .A1(n51480), .A2(n602), .ZN(n50159) );
  AND2_X1 U50445 ( .A1(n50160), .A2(n50159), .ZN(n50163) );
  NAND3_X1 U50446 ( .A1(n50161), .A2(n50233), .A3(n50192), .ZN(n50162) );
  NAND4_X1 U50447 ( .A1(n50165), .A2(n50164), .A3(n50163), .A4(n50162), .ZN(
        n50170) );
  NAND2_X1 U50448 ( .A1(n5799), .A2(n50222), .ZN(n50166) );
  AND2_X1 U50449 ( .A1(n50168), .A2(n50167), .ZN(n50169) );
  INV_X1 U50450 ( .A(n4897), .ZN(n50173) );
  INV_X1 U50451 ( .A(n50213), .ZN(n50176) );
  AND2_X1 U50452 ( .A1(n50234), .A2(n50189), .ZN(n50175) );
  NOR2_X1 U50453 ( .A1(n50233), .A2(n602), .ZN(n50231) );
  AOI21_X1 U50454 ( .B1(n50176), .B2(n50175), .A(n50231), .ZN(n50184) );
  INV_X1 U50455 ( .A(n50199), .ZN(n50177) );
  OAI211_X1 U50456 ( .C1(n50187), .C2(n50232), .A(n50177), .B(n50209), .ZN(
        n50183) );
  INV_X1 U50457 ( .A(n50224), .ZN(n50179) );
  NAND2_X1 U50458 ( .A1(n50179), .A2(n50178), .ZN(n50182) );
  NAND3_X1 U50460 ( .A1(n50232), .A2(n50208), .A3(n50180), .ZN(n50181) );
  NAND4_X1 U50461 ( .A1(n50184), .A2(n50183), .A3(n50182), .A4(n50181), .ZN(
        n50186) );
  INV_X1 U50462 ( .A(n3014), .ZN(n50185) );
  XNOR2_X1 U50463 ( .A(n50186), .B(n50185), .ZN(Plaintext[146]) );
  AND2_X1 U50464 ( .A1(n50196), .A2(n50234), .ZN(n50204) );
  OAI21_X1 U50465 ( .B1(n50188), .B2(n50204), .A(n50226), .ZN(n50195) );
  AND2_X1 U50466 ( .A1(n50189), .A2(n50192), .ZN(n50239) );
  NAND3_X1 U50467 ( .A1(n50191), .A2(n51480), .A3(n50239), .ZN(n50194) );
  NAND4_X1 U50468 ( .A1(n50209), .A2(n52099), .A3(n50222), .A4(n50192), .ZN(
        n50193) );
  NOR2_X1 U50469 ( .A1(n50233), .A2(n50196), .ZN(n50215) );
  OAI211_X1 U50470 ( .C1(n50215), .C2(n50235), .A(n50232), .B(n50222), .ZN(
        n50201) );
  INV_X1 U50471 ( .A(n50208), .ZN(n50197) );
  NAND3_X1 U50472 ( .A1(n50199), .A2(n50198), .A3(n50197), .ZN(n50200) );
  INV_X1 U50473 ( .A(n4739), .ZN(n50203) );
  INV_X1 U50474 ( .A(n50204), .ZN(n50207) );
  NAND2_X1 U50475 ( .A1(n50205), .A2(n50204), .ZN(n50206) );
  OAI21_X1 U50476 ( .B1(n50207), .B2(n50210), .A(n50206), .ZN(n50223) );
  INV_X1 U50477 ( .A(n50223), .ZN(n50219) );
  OAI22_X1 U50479 ( .A1(n50211), .A2(n50210), .B1(n50209), .B2(n50236), .ZN(
        n50212) );
  INV_X1 U50480 ( .A(n50212), .ZN(n50218) );
  NAND2_X1 U50481 ( .A1(n50214), .A2(n50213), .ZN(n50217) );
  NAND4_X1 U50482 ( .A1(n50232), .A2(n50222), .A3(n50215), .A4(n50235), .ZN(
        n50216) );
  INV_X1 U50484 ( .A(n4676), .ZN(n50220) );
  NOR2_X1 U50486 ( .A1(n50233), .A2(n50222), .ZN(n50225) );
  INV_X1 U50487 ( .A(n50242), .ZN(n50250) );
  NAND2_X1 U50488 ( .A1(n50227), .A2(n50226), .ZN(n50228) );
  NAND3_X1 U50489 ( .A1(n50228), .A2(n50233), .A3(n50234), .ZN(n50229) );
  AND2_X1 U50490 ( .A1(n50230), .A2(n50229), .ZN(n50244) );
  NAND2_X1 U50491 ( .A1(n50232), .A2(n50231), .ZN(n50240) );
  NAND3_X1 U50492 ( .A1(n52099), .A2(n602), .A3(n50233), .ZN(n50238) );
  NAND2_X1 U50493 ( .A1(n50235), .A2(n50234), .ZN(n50237) );
  NAND4_X1 U50494 ( .A1(n50239), .A2(n50238), .A3(n50237), .A4(n50236), .ZN(
        n50241) );
  NAND4_X1 U50495 ( .A1(n50244), .A2(n4618), .A3(n50240), .A4(n50241), .ZN(
        n50249) );
  INV_X1 U50496 ( .A(n4618), .ZN(n50245) );
  NAND2_X1 U50497 ( .A1(n50243), .A2(n50245), .ZN(n50248) );
  INV_X1 U50498 ( .A(n50244), .ZN(n50246) );
  NAND2_X1 U50499 ( .A1(n50246), .A2(n50245), .ZN(n50247) );
  OAI211_X1 U50500 ( .C1(n50250), .C2(n50249), .A(n50248), .B(n50247), .ZN(
        Plaintext[149]) );
  NAND3_X1 U50501 ( .A1(n658), .A2(n50251), .A3(n50253), .ZN(n50258) );
  NAND3_X1 U50502 ( .A1(n50253), .A2(n50252), .A3(n51372), .ZN(n50257) );
  AND2_X1 U50503 ( .A1(n6132), .A2(n50254), .ZN(n50264) );
  NAND3_X1 U50504 ( .A1(n50276), .A2(n50255), .A3(n50264), .ZN(n50256) );
  NAND2_X1 U50505 ( .A1(n50260), .A2(n50259), .ZN(n50273) );
  OAI21_X1 U50506 ( .B1(n50261), .B2(n50280), .A(n50277), .ZN(n50263) );
  NAND2_X1 U50507 ( .A1(n50263), .A2(n50262), .ZN(n50268) );
  NAND3_X1 U50508 ( .A1(n50266), .A2(n51410), .A3(n50264), .ZN(n50267) );
  NAND3_X1 U50509 ( .A1(n50281), .A2(n50278), .A3(n50277), .ZN(n50284) );
  NAND3_X1 U50510 ( .A1(n50281), .A2(n50280), .A3(n50279), .ZN(n50282) );
  AND2_X1 U50511 ( .A1(n51691), .A2(n50297), .ZN(n50290) );
  NAND2_X1 U50512 ( .A1(n50291), .A2(n50290), .ZN(n50313) );
  NAND2_X1 U50513 ( .A1(n51313), .A2(n50292), .ZN(n50295) );
  NAND4_X1 U50514 ( .A1(n50297), .A2(n50296), .A3(n50295), .A4(n50294), .ZN(
        n50302) );
  MUX2_X1 U50515 ( .A(n50302), .B(n50301), .S(n51691), .Z(n50312) );
  OAI211_X1 U50516 ( .C1(n7724), .C2(n50305), .A(n50304), .B(n50303), .ZN(
        n50306) );
  INV_X1 U50517 ( .A(n50306), .ZN(n50311) );
  NAND3_X1 U50518 ( .A1(n50309), .A2(n50308), .A3(n50307), .ZN(n50310) );
  AOI21_X1 U50519 ( .B1(n50315), .B2(n50314), .A(n6172), .ZN(n50318) );
  NAND2_X1 U50520 ( .A1(n50320), .A2(n50319), .ZN(n50327) );
  NOR2_X1 U50521 ( .A1(n50321), .A2(n50322), .ZN(n50323) );
  NOR2_X1 U50522 ( .A1(n50324), .A2(n50323), .ZN(n50326) );
  MUX2_X1 U50523 ( .A(n50327), .B(n50326), .S(n50325), .Z(n50407) );
  OAI21_X1 U50524 ( .B1(n50330), .B2(n50329), .A(n50328), .ZN(n50334) );
  NAND2_X1 U50525 ( .A1(n50332), .A2(n50331), .ZN(n50333) );
  NOR2_X1 U50526 ( .A1(n50334), .A2(n50333), .ZN(n50406) );
  NAND2_X1 U50527 ( .A1(n50335), .A2(n555), .ZN(n50336) );
  MUX2_X1 U50528 ( .A(n50340), .B(n51026), .S(n51725), .Z(n50356) );
  OAI21_X1 U50529 ( .B1(n51386), .B2(n50342), .A(n50341), .ZN(n50345) );
  NAND2_X1 U50530 ( .A1(n50345), .A2(n50344), .ZN(n50355) );
  OAI211_X1 U50531 ( .C1(n50349), .C2(n50348), .A(n50347), .B(n50346), .ZN(
        n50354) );
  NAND3_X1 U50532 ( .A1(n50352), .A2(n50351), .A3(n555), .ZN(n50353) );
  NAND2_X1 U50533 ( .A1(n50486), .A2(n50452), .ZN(n50357) );
  INV_X1 U50534 ( .A(n50452), .ZN(n50459) );
  NAND2_X1 U50536 ( .A1(n50470), .A2(n50482), .ZN(n50358) );
  NAND3_X1 U50537 ( .A1(n50368), .A2(n50367), .A3(n667), .ZN(n50369) );
  OAI21_X1 U50539 ( .B1(n50436), .B2(n50401), .A(n50373), .ZN(n50396) );
  AOI21_X1 U50540 ( .B1(n2198), .B2(n50390), .A(n51058), .ZN(n50376) );
  AOI21_X1 U50541 ( .B1(n50376), .B2(n50375), .A(n50378), .ZN(n50395) );
  NAND3_X1 U50542 ( .A1(n50378), .A2(n50386), .A3(n50377), .ZN(n50381) );
  NAND3_X1 U50543 ( .A1(n50381), .A2(n50380), .A3(n50379), .ZN(n50394) );
  NOR3_X1 U50544 ( .A1(n2198), .A2(n50386), .A3(n423), .ZN(n50384) );
  NOR2_X1 U50545 ( .A1(n50385), .A2(n50384), .ZN(n50392) );
  NAND2_X1 U50546 ( .A1(n50387), .A2(n50386), .ZN(n50388) );
  NAND2_X1 U50547 ( .A1(n50389), .A2(n50388), .ZN(n50391) );
  MUX2_X1 U50548 ( .A(n50392), .B(n50391), .S(n50390), .Z(n50393) );
  NOR2_X1 U50549 ( .A1(n50433), .A2(n50465), .ZN(n50457) );
  INV_X1 U50550 ( .A(n50457), .ZN(n50397) );
  OAI21_X1 U50551 ( .B1(n50397), .B2(n50483), .A(n50486), .ZN(n50399) );
  NAND2_X1 U50552 ( .A1(n50483), .A2(n50452), .ZN(n50412) );
  NOR2_X1 U50553 ( .A1(n50485), .A2(n50452), .ZN(n50408) );
  NAND3_X1 U50554 ( .A1(n50436), .A2(n7114), .A3(n50408), .ZN(n50398) );
  INV_X1 U50555 ( .A(n50433), .ZN(n50479) );
  NAND4_X1 U50556 ( .A1(n7114), .A2(n50479), .A3(n50482), .A4(n50483), .ZN(
        n50410) );
  INV_X1 U50557 ( .A(n4296), .ZN(n50400) );
  INV_X1 U50558 ( .A(n50401), .ZN(n50405) );
  NAND2_X1 U50559 ( .A1(n50433), .A2(n50485), .ZN(n50468) );
  NOR2_X1 U50560 ( .A1(n50436), .A2(n50468), .ZN(n50404) );
  OAI21_X1 U50561 ( .B1(n50465), .B2(n50483), .A(n50433), .ZN(n50453) );
  NAND2_X1 U50562 ( .A1(n7139), .A2(n50459), .ZN(n50402) );
  NOR2_X1 U50563 ( .A1(n50453), .A2(n50402), .ZN(n50403) );
  AOI22_X1 U50564 ( .A1(n50405), .A2(n50404), .B1(n50455), .B2(n50403), .ZN(
        n50423) );
  AND3_X1 U50565 ( .A1(n50407), .A2(n50406), .A3(n50483), .ZN(n50445) );
  NAND3_X1 U50566 ( .A1(n50445), .A2(n50408), .A3(n50482), .ZN(n50409) );
  NAND3_X1 U50567 ( .A1(n50485), .A2(n50452), .A3(n50483), .ZN(n50441) );
  AND2_X1 U50568 ( .A1(n50466), .A2(n50479), .ZN(n50417) );
  NAND2_X1 U50569 ( .A1(n50459), .A2(n50483), .ZN(n50469) );
  INV_X1 U50570 ( .A(n50412), .ZN(n50413) );
  NAND2_X1 U50571 ( .A1(n50413), .A2(n50482), .ZN(n50414) );
  OAI211_X1 U50572 ( .C1(n50451), .C2(n50469), .A(n50414), .B(n50486), .ZN(
        n50416) );
  NOR2_X1 U50573 ( .A1(n50459), .A2(n50483), .ZN(n50478) );
  OAI21_X1 U50574 ( .B1(n50417), .B2(n50416), .A(n50415), .ZN(n50421) );
  NAND2_X1 U50575 ( .A1(n50470), .A2(n50433), .ZN(n50418) );
  NOR2_X1 U50576 ( .A1(n50418), .A2(n50486), .ZN(n50419) );
  OAI22_X1 U50577 ( .A1(n50419), .A2(n50457), .B1(n50436), .B2(n50458), .ZN(
        n50420) );
  INV_X1 U50578 ( .A(n4788), .ZN(n50424) );
  INV_X1 U50579 ( .A(n50468), .ZN(n50425) );
  NAND2_X1 U50580 ( .A1(n50425), .A2(n50466), .ZN(n50426) );
  NAND3_X1 U50581 ( .A1(n50440), .A2(n50445), .A3(n50426), .ZN(n50430) );
  AND2_X1 U50582 ( .A1(n50485), .A2(n50486), .ZN(n50481) );
  OAI211_X1 U50583 ( .C1(n50481), .C2(n50466), .A(n7139), .B(n50433), .ZN(
        n50429) );
  INV_X1 U50584 ( .A(n50458), .ZN(n50427) );
  NAND4_X1 U50585 ( .A1(n50427), .A2(n50436), .A3(n50459), .A4(n50433), .ZN(
        n50428) );
  AND2_X1 U50588 ( .A1(n50433), .A2(n50483), .ZN(n50471) );
  AND2_X1 U50589 ( .A1(n7114), .A2(n50471), .ZN(n50434) );
  NAND2_X1 U50590 ( .A1(n50435), .A2(n7139), .ZN(n50439) );
  INV_X1 U50591 ( .A(n50469), .ZN(n50437) );
  NAND3_X1 U50592 ( .A1(n50437), .A2(n50479), .A3(n50436), .ZN(n50438) );
  INV_X1 U50593 ( .A(n50440), .ZN(n50444) );
  NAND3_X1 U50594 ( .A1(n50445), .A2(n50479), .A3(n50452), .ZN(n50442) );
  NAND2_X1 U50595 ( .A1(n50442), .A2(n50441), .ZN(n50443) );
  AOI21_X1 U50596 ( .B1(n50458), .B2(n50444), .A(n50443), .ZN(n50448) );
  NOR2_X1 U50597 ( .A1(n50451), .A2(n50482), .ZN(n50446) );
  NAND2_X1 U50598 ( .A1(n50446), .A2(n50445), .ZN(n50460) );
  INV_X1 U50599 ( .A(n4638), .ZN(n50450) );
  AOI21_X1 U50600 ( .B1(n7139), .B2(n50451), .A(n50481), .ZN(n50456) );
  INV_X1 U50601 ( .A(n50473), .ZN(n50476) );
  INV_X1 U50602 ( .A(n50453), .ZN(n50454) );
  OAI21_X1 U50603 ( .B1(n50460), .B2(n50459), .A(n50477), .ZN(n50461) );
  NAND3_X1 U50606 ( .A1(n50479), .A2(n7139), .A3(n50482), .ZN(n50467) );
  INV_X1 U50607 ( .A(n50471), .ZN(n50474) );
  NAND3_X1 U50608 ( .A1(n7114), .A2(n50471), .A3(n50470), .ZN(n50472) );
  OAI21_X1 U50609 ( .B1(n50474), .B2(n50473), .A(n50472), .ZN(n50475) );
  OAI21_X1 U50610 ( .B1(n50479), .B2(n50482), .A(n50478), .ZN(n50480) );
  XNOR2_X1 U50611 ( .A(n50482), .B(n50486), .ZN(n50484) );
  OAI211_X1 U50612 ( .C1(n50486), .C2(n50485), .A(n50484), .B(n50483), .ZN(
        n50487) );
  INV_X1 U50613 ( .A(n4487), .ZN(n50488) );
  NAND2_X1 U50614 ( .A1(n50542), .A2(n50550), .ZN(n50536) );
  AOI21_X1 U50615 ( .B1(n50536), .B2(n50541), .A(n50533), .ZN(n50502) );
  INV_X1 U50616 ( .A(n50495), .ZN(n50489) );
  OAI211_X1 U50617 ( .C1(n50489), .C2(n50552), .A(n50497), .B(n50562), .ZN(
        n50501) );
  AND2_X1 U50618 ( .A1(n50555), .A2(n50550), .ZN(n50565) );
  AND2_X1 U50619 ( .A1(n50553), .A2(n50533), .ZN(n50504) );
  AOI22_X1 U50620 ( .A1(n50504), .A2(n50555), .B1(n50490), .B2(n50533), .ZN(
        n50493) );
  NOR2_X1 U50621 ( .A1(n50562), .A2(n50552), .ZN(n50491) );
  NAND4_X1 U50622 ( .A1(n50491), .A2(n50554), .A3(n50520), .A4(n50564), .ZN(
        n50492) );
  NAND4_X1 U50623 ( .A1(n50495), .A2(n50553), .A3(n50554), .A4(n50552), .ZN(
        n50496) );
  OR2_X1 U50624 ( .A1(n50552), .A2(n50520), .ZN(n50561) );
  OAI21_X1 U50625 ( .B1(n50561), .B2(n50555), .A(n50562), .ZN(n50500) );
  INV_X1 U50627 ( .A(n4712), .ZN(n50503) );
  AND2_X1 U50628 ( .A1(n1151), .A2(n50527), .ZN(n50506) );
  INV_X1 U50629 ( .A(n50548), .ZN(n50505) );
  AOI21_X1 U50630 ( .B1(n50506), .B2(n50505), .A(n50504), .ZN(n50514) );
  NAND2_X1 U50631 ( .A1(n50526), .A2(n50554), .ZN(n50543) );
  OR2_X1 U50632 ( .A1(n50543), .A2(n50555), .ZN(n50513) );
  INV_X1 U50633 ( .A(n50536), .ZN(n50507) );
  OAI21_X1 U50634 ( .B1(n50539), .B2(n50534), .A(n50507), .ZN(n50512) );
  OAI21_X1 U50635 ( .B1(n50555), .B2(n50508), .A(n50533), .ZN(n50509) );
  NAND2_X1 U50636 ( .A1(n50509), .A2(n50564), .ZN(n50510) );
  NAND2_X1 U50637 ( .A1(n50510), .A2(n50526), .ZN(n50511) );
  NAND4_X1 U50638 ( .A1(n50514), .A2(n50513), .A3(n50512), .A4(n50511), .ZN(
        n50516) );
  INV_X1 U50639 ( .A(n4641), .ZN(n50515) );
  XNOR2_X1 U50640 ( .A(n50516), .B(n50515), .ZN(Plaintext[158]) );
  OAI21_X1 U50641 ( .B1(n50551), .B2(n50552), .A(n50533), .ZN(n50519) );
  NAND2_X1 U50642 ( .A1(n50521), .A2(n50553), .ZN(n50523) );
  NAND2_X1 U50643 ( .A1(n50550), .A2(n50554), .ZN(n50522) );
  OAI22_X1 U50644 ( .A1(n50563), .A2(n50523), .B1(n50541), .B2(n50522), .ZN(
        n50524) );
  INV_X1 U50645 ( .A(n50524), .ZN(n50531) );
  NAND3_X1 U50646 ( .A1(n50526), .A2(n50555), .A3(n50525), .ZN(n50530) );
  INV_X1 U50647 ( .A(n50527), .ZN(n50528) );
  NAND3_X1 U50648 ( .A1(n50528), .A2(n50554), .A3(n50551), .ZN(n50529) );
  INV_X1 U50649 ( .A(n3367), .ZN(n50532) );
  NAND2_X1 U50650 ( .A1(n50563), .A2(n50562), .ZN(n50535) );
  NAND2_X1 U50651 ( .A1(n51349), .A2(n50564), .ZN(n50558) );
  OAI21_X1 U50652 ( .B1(n50535), .B2(n50548), .A(n50558), .ZN(n50538) );
  NOR2_X1 U50653 ( .A1(n50538), .A2(n50537), .ZN(n50545) );
  OAI21_X1 U50654 ( .B1(n50540), .B2(n50565), .A(n50539), .ZN(n50549) );
  OR3_X1 U50655 ( .A1(n50543), .A2(n50542), .A3(n50541), .ZN(n50544) );
  XNOR2_X1 U50656 ( .A(n50547), .B(n50546), .ZN(Plaintext[160]) );
  NOR2_X1 U50657 ( .A1(n50551), .A2(n50550), .ZN(n50560) );
  OAI21_X1 U50658 ( .B1(n50555), .B2(n50552), .A(n50562), .ZN(n50559) );
  NOR2_X1 U50659 ( .A1(n50553), .A2(n50552), .ZN(n50556) );
  OAI21_X1 U50660 ( .B1(n50556), .B2(n50555), .A(n50554), .ZN(n50557) );
  NAND4_X1 U50661 ( .A1(n50560), .A2(n50559), .A3(n50558), .A4(n50557), .ZN(
        n50568) );
  AND3_X1 U50662 ( .A1(n50563), .A2(n50562), .A3(n50561), .ZN(n50566) );
  OAI21_X1 U50663 ( .B1(n50566), .B2(n50565), .A(n50564), .ZN(n50567) );
  INV_X1 U50664 ( .A(n4612), .ZN(n50570) );
  XNOR2_X1 U50665 ( .A(n50571), .B(n50570), .ZN(Plaintext[161]) );
  INV_X1 U50666 ( .A(n50588), .ZN(n50572) );
  OAI21_X1 U50667 ( .B1(n50573), .B2(n50633), .A(n50572), .ZN(n50574) );
  NAND3_X1 U50668 ( .A1(n50574), .A2(n50642), .A3(n51029), .ZN(n50585) );
  AOI21_X1 U50669 ( .B1(n8018), .B2(n52226), .A(n50641), .ZN(n50577) );
  OR2_X1 U50670 ( .A1(n50588), .A2(n51029), .ZN(n50576) );
  AND2_X1 U50671 ( .A1(n52225), .A2(n52081), .ZN(n50643) );
  AOI22_X1 U50672 ( .A1(n50577), .A2(n50576), .B1(n50575), .B2(n50643), .ZN(
        n50584) );
  NAND3_X1 U50673 ( .A1(n50642), .A2(n50579), .A3(n50615), .ZN(n50580) );
  NAND2_X1 U50674 ( .A1(n50638), .A2(n52082), .ZN(n50621) );
  NAND4_X1 U50675 ( .A1(n50580), .A2(n50618), .A3(n52061), .A4(n50622), .ZN(
        n50583) );
  INV_X1 U50676 ( .A(n50624), .ZN(n50581) );
  INV_X1 U50677 ( .A(n50621), .ZN(n50632) );
  NAND3_X1 U50678 ( .A1(n50581), .A2(n50632), .A3(n51029), .ZN(n50582) );
  NAND4_X1 U50679 ( .A1(n50585), .A2(n50584), .A3(n50583), .A4(n50582), .ZN(
        n50587) );
  XNOR2_X1 U50680 ( .A(n50587), .B(n50586), .ZN(Plaintext[162]) );
  NAND3_X1 U50681 ( .A1(n50588), .A2(n50638), .A3(n50615), .ZN(n50590) );
  MUX2_X1 U50682 ( .A(n50590), .B(n50589), .S(n50644), .Z(n50606) );
  INV_X1 U50683 ( .A(n50591), .ZN(n50592) );
  NAND4_X1 U50684 ( .A1(n50592), .A2(n50611), .A3(n50638), .A4(n50641), .ZN(
        n50594) );
  OAI21_X1 U50685 ( .B1(n50594), .B2(n50618), .A(n50593), .ZN(n50597) );
  OR2_X1 U50686 ( .A1(n50622), .A2(n51029), .ZN(n50595) );
  NAND2_X1 U50687 ( .A1(n50643), .A2(n50630), .ZN(n50617) );
  OAI211_X1 U50688 ( .C1(n50624), .C2(n52061), .A(n50595), .B(n50617), .ZN(
        n50596) );
  NOR2_X1 U50689 ( .A1(n50597), .A2(n50596), .ZN(n50605) );
  AND2_X1 U50690 ( .A1(n50610), .A2(n8018), .ZN(n50603) );
  INV_X1 U50691 ( .A(n50599), .ZN(n50600) );
  AOI21_X1 U50692 ( .B1(n50615), .B2(n50600), .A(n50638), .ZN(n50602) );
  AND2_X1 U50693 ( .A1(n50618), .A2(n52225), .ZN(n50601) );
  OAI22_X1 U50694 ( .A1(n50603), .A2(n50602), .B1(n50633), .B2(n50601), .ZN(
        n50604) );
  INV_X1 U50695 ( .A(n4930), .ZN(n50607) );
  XNOR2_X1 U50696 ( .A(n50608), .B(n50607), .ZN(Plaintext[163]) );
  NAND2_X1 U50697 ( .A1(n50630), .A2(n51029), .ZN(n50612) );
  OAI21_X1 U50698 ( .B1(n50615), .B2(n50611), .A(n50642), .ZN(n50614) );
  OAI21_X1 U50699 ( .B1(n50612), .B2(n52082), .A(n50638), .ZN(n50613) );
  OR2_X1 U50700 ( .A1(n50615), .A2(n50621), .ZN(n50616) );
  AND2_X1 U50701 ( .A1(n50617), .A2(n50616), .ZN(n50627) );
  OAI211_X1 U50702 ( .C1(n50638), .C2(n52081), .A(n50619), .B(n50618), .ZN(
        n50626) );
  NAND2_X1 U50703 ( .A1(n50622), .A2(n50621), .ZN(n50623) );
  NAND3_X1 U50704 ( .A1(n50624), .A2(n50641), .A3(n50623), .ZN(n50625) );
  INV_X1 U50705 ( .A(n4579), .ZN(n50628) );
  XNOR2_X1 U50706 ( .A(n50629), .B(n50628), .ZN(Plaintext[165]) );
  OR2_X1 U50707 ( .A1(n50631), .A2(n50630), .ZN(n50636) );
  MUX2_X1 U50708 ( .A(n50636), .B(n50635), .S(n50634), .Z(n50647) );
  NAND2_X1 U50709 ( .A1(n50638), .A2(n51029), .ZN(n50639) );
  AOI21_X1 U50710 ( .B1(n50641), .B2(n52225), .A(n50639), .ZN(n50645) );
  AOI22_X1 U50711 ( .A1(n50645), .A2(n50644), .B1(n50643), .B2(n50642), .ZN(
        n50646) );
  INV_X1 U50712 ( .A(n4471), .ZN(n50648) );
  XNOR2_X1 U50713 ( .A(n50649), .B(n50648), .ZN(Plaintext[166]) );
  OAI21_X1 U50714 ( .B1(n51367), .B2(n50721), .A(n50680), .ZN(n50686) );
  INV_X1 U50715 ( .A(n50710), .ZN(n50652) );
  NAND3_X1 U50716 ( .A1(n50686), .A2(n50652), .A3(n50731), .ZN(n50659) );
  NAND2_X1 U50717 ( .A1(n50721), .A2(n50716), .ZN(n50732) );
  NAND2_X1 U50718 ( .A1(n50732), .A2(n50705), .ZN(n50654) );
  NAND2_X1 U50719 ( .A1(n50727), .A2(n50679), .ZN(n50663) );
  OAI21_X1 U50720 ( .B1(n50727), .B2(n50700), .A(n50663), .ZN(n50653) );
  NAND2_X1 U50721 ( .A1(n50654), .A2(n50653), .ZN(n50658) );
  AND2_X1 U50722 ( .A1(n50721), .A2(n50708), .ZN(n50656) );
  NOR2_X1 U50723 ( .A1(n50681), .A2(n50679), .ZN(n50709) );
  AOI22_X1 U50724 ( .A1(n50656), .A2(n50709), .B1(n50727), .B2(n50655), .ZN(
        n50657) );
  NAND4_X1 U50725 ( .A1(n50660), .A2(n50659), .A3(n50658), .A4(n50657), .ZN(
        n50662) );
  INV_X1 U50726 ( .A(n4706), .ZN(n50661) );
  XNOR2_X1 U50727 ( .A(n50662), .B(n50661), .ZN(Plaintext[168]) );
  AND2_X1 U50728 ( .A1(n50709), .A2(n50708), .ZN(n50687) );
  OAI211_X1 U50729 ( .C1(n50727), .C2(n50716), .A(n50663), .B(n50721), .ZN(
        n50664) );
  AOI22_X1 U50730 ( .A1(n50687), .A2(n51367), .B1(n50664), .B2(n50728), .ZN(
        n50672) );
  INV_X1 U50731 ( .A(n50717), .ZN(n50666) );
  NAND3_X1 U50732 ( .A1(n50666), .A2(n50680), .A3(n50665), .ZN(n50671) );
  INV_X1 U50733 ( .A(n50723), .ZN(n50670) );
  INV_X1 U50734 ( .A(n50732), .ZN(n50668) );
  OAI21_X1 U50735 ( .B1(n50668), .B2(n50718), .A(n50667), .ZN(n50669) );
  NAND4_X1 U50736 ( .A1(n50672), .A2(n50671), .A3(n50670), .A4(n50669), .ZN(
        n50674) );
  INV_X1 U50737 ( .A(n4295), .ZN(n50673) );
  XNOR2_X1 U50738 ( .A(n50674), .B(n50673), .ZN(Plaintext[170]) );
  NAND2_X1 U50739 ( .A1(n50727), .A2(n50681), .ZN(n50678) );
  NAND2_X1 U50740 ( .A1(n50676), .A2(n50716), .ZN(n50677) );
  AND2_X1 U50741 ( .A1(n50679), .A2(n50708), .ZN(n50694) );
  NAND2_X1 U50742 ( .A1(n50694), .A2(n50680), .ZN(n50733) );
  OAI21_X1 U50743 ( .B1(n50733), .B2(n50721), .A(n1224), .ZN(n50683) );
  NAND2_X1 U50744 ( .A1(n50681), .A2(n50708), .ZN(n50722) );
  NOR2_X1 U50745 ( .A1(n50722), .A2(n50704), .ZN(n50682) );
  NOR2_X1 U50746 ( .A1(n50683), .A2(n50682), .ZN(n50684) );
  AND2_X1 U50747 ( .A1(n50721), .A2(n50734), .ZN(n50685) );
  AND2_X1 U50749 ( .A1(n50687), .A2(n50686), .ZN(n50691) );
  INV_X1 U50750 ( .A(n50691), .ZN(n50688) );
  OAI21_X1 U50751 ( .B1(n50693), .B2(n50689), .A(n50688), .ZN(n50699) );
  INV_X1 U50752 ( .A(n1224), .ZN(n50696) );
  OAI21_X1 U50753 ( .B1(n50691), .B2(n50690), .A(n50696), .ZN(n50698) );
  NOR2_X1 U50755 ( .A1(n50721), .A2(n50716), .ZN(n50701) );
  INV_X1 U50756 ( .A(n50701), .ZN(n50703) );
  NAND3_X1 U50757 ( .A1(n50703), .A2(n50731), .A3(n50694), .ZN(n50695) );
  NAND2_X1 U50758 ( .A1(n50701), .A2(n50700), .ZN(n50719) );
  NAND2_X1 U50759 ( .A1(n50719), .A2(n50718), .ZN(n50713) );
  NAND2_X1 U50760 ( .A1(n50704), .A2(n50727), .ZN(n50702) );
  AOI21_X1 U50761 ( .B1(n51367), .B2(n50705), .A(n50704), .ZN(n50706) );
  NAND2_X1 U50762 ( .A1(n50707), .A2(n50706), .ZN(n50712) );
  NAND4_X1 U50763 ( .A1(n50710), .A2(n50727), .A3(n50709), .A4(n50708), .ZN(
        n50711) );
  INV_X1 U50764 ( .A(n4864), .ZN(n50714) );
  XNOR2_X1 U50765 ( .A(n50715), .B(n50714), .ZN(Plaintext[172]) );
  NAND2_X1 U50766 ( .A1(n50733), .A2(n1467), .ZN(n50725) );
  NAND2_X1 U50767 ( .A1(n50722), .A2(n50721), .ZN(n50724) );
  NAND3_X1 U50768 ( .A1(n50728), .A2(n50727), .A3(n50726), .ZN(n50729) );
  NOR2_X1 U50769 ( .A1(n50732), .A2(n50731), .ZN(n50736) );
  INV_X1 U50770 ( .A(n50733), .ZN(n50735) );
  MUX2_X1 U50771 ( .A(n50736), .B(n50735), .S(n51367), .Z(n50737) );
  XNOR2_X1 U50772 ( .A(n50779), .B(n50809), .ZN(n50738) );
  AOI21_X1 U50773 ( .B1(n50739), .B2(n50761), .A(n2095), .ZN(n50742) );
  NAND2_X1 U50774 ( .A1(n50787), .A2(n51353), .ZN(n50740) );
  NAND2_X1 U50775 ( .A1(n50751), .A2(n50809), .ZN(n50812) );
  NAND2_X1 U50776 ( .A1(n50744), .A2(n51730), .ZN(n50743) );
  OAI22_X1 U50777 ( .A1(n50740), .A2(n50812), .B1(n50743), .B2(n50779), .ZN(
        n50741) );
  NOR2_X1 U50778 ( .A1(n50742), .A2(n50741), .ZN(n50757) );
  NOR2_X1 U50779 ( .A1(n51354), .A2(n50773), .ZN(n50745) );
  OAI21_X1 U50780 ( .B1(n50745), .B2(n50751), .A(n50743), .ZN(n50746) );
  NAND2_X1 U50781 ( .A1(n51353), .A2(n2095), .ZN(n50765) );
  NAND2_X1 U50782 ( .A1(n50746), .A2(n50765), .ZN(n50749) );
  AND2_X1 U50783 ( .A1(n50809), .A2(n51296), .ZN(n50788) );
  OAI21_X1 U50784 ( .B1(n50747), .B2(n51353), .A(n50783), .ZN(n50748) );
  AOI22_X1 U50785 ( .A1(n50749), .A2(n50788), .B1(n50748), .B2(n50804), .ZN(
        n50756) );
  INV_X1 U50786 ( .A(n50765), .ZN(n50750) );
  NAND3_X1 U50787 ( .A1(n50750), .A2(n51730), .A3(n50809), .ZN(n50754) );
  NAND4_X1 U50788 ( .A1(n50752), .A2(n52076), .A3(n50751), .A4(n50808), .ZN(
        n50753) );
  AND2_X1 U50789 ( .A1(n50754), .A2(n50753), .ZN(n50755) );
  NAND2_X1 U50792 ( .A1(n50763), .A2(n50804), .ZN(n50769) );
  INV_X1 U50793 ( .A(n50764), .ZN(n50799) );
  AOI21_X1 U50794 ( .B1(n50765), .B2(n50812), .A(n50799), .ZN(n50767) );
  OAI211_X1 U50795 ( .C1(n50781), .C2(n51730), .A(n50797), .B(n50808), .ZN(
        n50766) );
  INV_X1 U50796 ( .A(n4746), .ZN(n50770) );
  NAND2_X1 U50797 ( .A1(n50798), .A2(n50787), .ZN(n50807) );
  NAND2_X1 U50798 ( .A1(n51354), .A2(n50773), .ZN(n50777) );
  AND2_X1 U50799 ( .A1(n51353), .A2(n51296), .ZN(n50800) );
  NOR2_X1 U50800 ( .A1(n50773), .A2(n2095), .ZN(n50805) );
  OAI21_X1 U50802 ( .B1(n50797), .B2(n50809), .A(n50774), .ZN(n50775) );
  OAI211_X1 U50803 ( .C1(n50807), .C2(n50777), .A(n50776), .B(n50775), .ZN(
        n50778) );
  INV_X1 U50804 ( .A(n50778), .ZN(n50794) );
  NAND2_X1 U50805 ( .A1(n50807), .A2(n50779), .ZN(n50782) );
  NAND4_X1 U50806 ( .A1(n50782), .A2(n52076), .A3(n51296), .A4(n51730), .ZN(
        n50793) );
  NOR2_X1 U50807 ( .A1(n50798), .A2(n50783), .ZN(n50785) );
  OAI21_X1 U50808 ( .B1(n50786), .B2(n50785), .A(n51730), .ZN(n50792) );
  OR2_X1 U50809 ( .A1(n50788), .A2(n50787), .ZN(n50790) );
  NAND4_X1 U50810 ( .A1(n50807), .A2(n50790), .A3(n50773), .A4(n50812), .ZN(
        n50791) );
  INV_X1 U50811 ( .A(n4565), .ZN(n50795) );
  AOI21_X1 U50812 ( .B1(n50799), .B2(n50798), .A(n50797), .ZN(n50803) );
  INV_X1 U50813 ( .A(n50800), .ZN(n50801) );
  OAI21_X1 U50814 ( .B1(n50807), .B2(n50801), .A(n50804), .ZN(n50802) );
  OAI21_X1 U50815 ( .B1(n50804), .B2(n50803), .A(n50802), .ZN(n50816) );
  INV_X1 U50816 ( .A(n50805), .ZN(n50806) );
  NAND2_X1 U50817 ( .A1(n50807), .A2(n50806), .ZN(n50810) );
  NAND3_X1 U50818 ( .A1(n50810), .A2(n50809), .A3(n50808), .ZN(n50814) );
  OR2_X1 U50819 ( .A1(n50812), .A2(n50811), .ZN(n50813) );
  INV_X1 U50820 ( .A(n4687), .ZN(n50817) );
  AND2_X1 U50821 ( .A1(n50850), .A2(n50826), .ZN(n50880) );
  NAND2_X1 U50822 ( .A1(n50863), .A2(n50837), .ZN(n50819) );
  NAND2_X1 U50823 ( .A1(n50819), .A2(n51312), .ZN(n50889) );
  OAI21_X1 U50824 ( .B1(n50864), .B2(n52098), .A(n50889), .ZN(n50820) );
  NOR2_X1 U50825 ( .A1(n50837), .A2(n50886), .ZN(n50855) );
  AND2_X1 U50826 ( .A1(n50855), .A2(n50894), .ZN(n50870) );
  INV_X1 U50827 ( .A(n50892), .ZN(n50839) );
  NOR2_X1 U50828 ( .A1(n50894), .A2(n50837), .ZN(n50821) );
  NOR2_X1 U50829 ( .A1(n52097), .A2(n52098), .ZN(n50822) );
  NOR2_X1 U50830 ( .A1(n50863), .A2(n50837), .ZN(n50835) );
  INV_X1 U50831 ( .A(n1326), .ZN(n50825) );
  AOI22_X1 U50833 ( .A1(n50869), .A2(n50855), .B1(n50831), .B2(n50829), .ZN(
        n50827) );
  MUX2_X1 U50834 ( .A(n50828), .B(n50827), .S(n50850), .Z(n50844) );
  NAND2_X1 U50836 ( .A1(n52063), .A2(n601), .ZN(n50830) );
  NAND2_X1 U50837 ( .A1(n50853), .A2(n50830), .ZN(n50833) );
  NAND3_X1 U50838 ( .A1(n50887), .A2(n50848), .A3(n50883), .ZN(n50832) );
  AND3_X1 U50839 ( .A1(n50833), .A2(n50832), .A3(n50897), .ZN(n50843) );
  INV_X1 U50840 ( .A(n50869), .ZN(n50834) );
  NAND4_X1 U50841 ( .A1(n50836), .A2(n50835), .A3(n50834), .A4(n50886), .ZN(
        n50842) );
  NAND2_X1 U50842 ( .A1(n52097), .A2(n50890), .ZN(n50840) );
  NAND2_X1 U50843 ( .A1(n50837), .A2(n50886), .ZN(n50862) );
  NAND4_X1 U50844 ( .A1(n50840), .A2(n50839), .A3(n52063), .A4(n50862), .ZN(
        n50841) );
  NAND4_X1 U50845 ( .A1(n50844), .A2(n50843), .A3(n50842), .A4(n50841), .ZN(
        n50846) );
  INV_X1 U50846 ( .A(n4667), .ZN(n50845) );
  XNOR2_X1 U50847 ( .A(n50846), .B(n50845), .ZN(Plaintext[181]) );
  OAI211_X1 U50848 ( .C1(n5295), .C2(n50883), .A(n50849), .B(n601), .ZN(n50858) );
  NAND2_X1 U50849 ( .A1(n50864), .A2(n50850), .ZN(n50852) );
  OAI22_X1 U50850 ( .A1(n50882), .A2(n50853), .B1(n50852), .B2(n50851), .ZN(
        n50857) );
  NAND2_X1 U50851 ( .A1(n50855), .A2(n601), .ZN(n50871) );
  NAND2_X1 U50852 ( .A1(n50887), .A2(n50880), .ZN(n50856) );
  NAND4_X1 U50853 ( .A1(n50858), .A2(n50857), .A3(n344), .A4(n50856), .ZN(
        n50860) );
  INV_X1 U50854 ( .A(n4909), .ZN(n50859) );
  XNOR2_X1 U50855 ( .A(n50860), .B(n50859), .ZN(Plaintext[182]) );
  OR2_X1 U50856 ( .A1(n50873), .A2(n50861), .ZN(n50877) );
  AND3_X1 U50857 ( .A1(n50892), .A2(n50894), .A3(n50862), .ZN(n50868) );
  OAI21_X1 U50858 ( .B1(n52093), .B2(n52098), .A(n51312), .ZN(n50867) );
  OAI22_X1 U50859 ( .A1(n50864), .A2(n50894), .B1(n50890), .B2(n50863), .ZN(
        n50866) );
  AOI22_X1 U50860 ( .A1(n50868), .A2(n50867), .B1(n50866), .B2(n52098), .ZN(
        n50876) );
  NAND2_X1 U50861 ( .A1(n50870), .A2(n50869), .ZN(n50875) );
  NAND3_X1 U50862 ( .A1(n50873), .A2(n50872), .A3(n50871), .ZN(n50874) );
  NAND4_X1 U50863 ( .A1(n50877), .A2(n50876), .A3(n50875), .A4(n50874), .ZN(
        n50879) );
  INV_X1 U50864 ( .A(n4940), .ZN(n50878) );
  XNOR2_X1 U50865 ( .A(n50879), .B(n50878), .ZN(Plaintext[183]) );
  INV_X1 U50866 ( .A(n50880), .ZN(n50881) );
  NAND2_X1 U50867 ( .A1(n50882), .A2(n50881), .ZN(n50885) );
  INV_X1 U50868 ( .A(n50883), .ZN(n50884) );
  OAI211_X1 U50869 ( .C1(n50887), .C2(n50886), .A(n50885), .B(n50884), .ZN(
        n50898) );
  NAND2_X1 U50870 ( .A1(n6817), .A2(n50889), .ZN(n50895) );
  OAI21_X1 U50871 ( .B1(n50892), .B2(n52093), .A(n50890), .ZN(n50893) );
  NAND3_X1 U50872 ( .A1(n50895), .A2(n50894), .A3(n50893), .ZN(n50896) );
  NAND3_X1 U50873 ( .A1(n50898), .A2(n50897), .A3(n50896), .ZN(n50900) );
  XNOR2_X1 U50874 ( .A(n50900), .B(n50899), .ZN(Plaintext[184]) );
  NOR2_X1 U50875 ( .A1(n50928), .A2(n50913), .ZN(n50927) );
  AOI22_X1 U50876 ( .A1(n50927), .A2(n50929), .B1(n50925), .B2(n50955), .ZN(
        n50904) );
  OR2_X1 U50877 ( .A1(n50950), .A2(n51486), .ZN(n50902) );
  AND2_X1 U50878 ( .A1(n50904), .A2(n50944), .ZN(n50922) );
  NAND2_X1 U50879 ( .A1(n50953), .A2(n50950), .ZN(n50908) );
  NAND4_X1 U50880 ( .A1(n50949), .A2(n50934), .A3(n50913), .A4(n50906), .ZN(
        n50907) );
  OAI21_X1 U50881 ( .B1(n50909), .B2(n50908), .A(n50907), .ZN(n50912) );
  INV_X1 U50882 ( .A(n50910), .ZN(n50911) );
  NOR3_X1 U50883 ( .A1(n50925), .A2(n50934), .A3(n50955), .ZN(n50919) );
  INV_X1 U50884 ( .A(n50950), .ZN(n50914) );
  NAND4_X1 U50885 ( .A1(n50914), .A2(n51486), .A3(n50929), .A4(n50913), .ZN(
        n50915) );
  NAND2_X1 U50886 ( .A1(n50916), .A2(n50915), .ZN(n50918) );
  AOI22_X1 U50887 ( .A1(n50919), .A2(n50918), .B1(n50917), .B2(n50916), .ZN(
        n50921) );
  INV_X1 U50888 ( .A(n4934), .ZN(n50923) );
  NOR2_X1 U50889 ( .A1(n50955), .A2(n50958), .ZN(n50924) );
  MUX2_X1 U50890 ( .A(n50925), .B(n50924), .S(n50953), .Z(n50926) );
  NAND2_X1 U50891 ( .A1(n50926), .A2(n5365), .ZN(n50942) );
  NAND2_X1 U50892 ( .A1(n50927), .A2(n50958), .ZN(n50931) );
  NAND3_X1 U50893 ( .A1(n50928), .A2(n51486), .A3(n50950), .ZN(n50930) );
  MUX2_X1 U50894 ( .A(n50931), .B(n50930), .S(n50929), .Z(n50941) );
  OAI211_X1 U50895 ( .C1(n50935), .C2(n50934), .A(n50933), .B(n50932), .ZN(
        n50936) );
  INV_X1 U50896 ( .A(n50936), .ZN(n50940) );
  NAND4_X1 U50898 ( .A1(n50942), .A2(n50941), .A3(n50940), .A4(n50939), .ZN(
        n50943) );
  XNOR2_X1 U50899 ( .A(n50943), .B(n3111), .ZN(Plaintext[189]) );
  NOR2_X1 U50900 ( .A1(n50946), .A2(n50950), .ZN(n50948) );
  AOI21_X1 U50901 ( .B1(n50949), .B2(n50948), .A(n50947), .ZN(n50962) );
  XNOR2_X1 U50902 ( .A(n50950), .B(n50955), .ZN(n50952) );
  NAND2_X1 U50903 ( .A1(n50952), .A2(n51486), .ZN(n50954) );
  AOI22_X1 U50904 ( .A1(n50956), .A2(n50955), .B1(n50954), .B2(n50953), .ZN(
        n50961) );
  OAI21_X1 U50905 ( .B1(n50959), .B2(n50958), .A(n50957), .ZN(n50960) );
  INV_X1 U50906 ( .A(n4668), .ZN(n50964) );
  OR2_X2 U60 ( .A1(n52054), .A2(n37781), .ZN(n39342) );
  AND2_X2 U2609 ( .A1(n6218), .A2(n51077), .ZN(n2043) );
  BUF_X2 U4853 ( .A(n12740), .Z(n15770) );
  BUF_X1 U3320 ( .A(n45560), .Z(n48522) );
  AND2_X2 U3644 ( .A1(n37988), .A2(n37974), .ZN(n37991) );
  BUF_X1 U4110 ( .A(n27278), .Z(n30407) );
  BUF_X2 U185 ( .A(n19277), .Z(n20441) );
  INV_X2 U605 ( .A(n24001), .ZN(n23986) );
  NAND4_X2 U5119 ( .A1(n38883), .A2(n38884), .A3(n38882), .A4(n38881), .ZN(
        n44061) );
  AND2_X2 U2872 ( .A1(n11601), .A2(n9083), .ZN(n11593) );
  OAI21_X2 U4914 ( .B1(n12437), .B2(n12436), .A(n12435), .ZN(n12449) );
  BUF_X2 U2753 ( .A(n20787), .Z(n23090) );
  INV_X1 U3700 ( .A(n35939), .ZN(n37775) );
  BUF_X2 U4565 ( .A(n17740), .Z(n21463) );
  OR2_X2 U3214 ( .A1(n49977), .A2(n49982), .ZN(n49626) );
  OR2_X2 U4258 ( .A1(n22230), .A2(n22229), .ZN(n24792) );
  INV_X1 U582 ( .A(n32701), .ZN(n31658) );
  BUF_X2 U4402 ( .A(n21016), .Z(n22864) );
  OAI21_X2 U4904 ( .B1(n11214), .B2(n9496), .A(n11204), .ZN(n9505) );
  NAND2_X2 U2801 ( .A1(n6074), .A2(n2873), .ZN(n18749) );
  OAI211_X2 U9224 ( .C1(n20160), .C2(n20166), .A(n20165), .B(n20164), .ZN(
        n23409) );
  BUF_X2 U4268 ( .A(n25771), .Z(n750) );
  AND2_X2 U4792 ( .A1(n14455), .A2(n14453), .ZN(n14434) );
  AND2_X2 U33081 ( .A1(n24570), .A2(n27732), .ZN(n27719) );
  BUF_X2 U4544 ( .A(n21212), .Z(n2229) );
  OR2_X2 U10370 ( .A1(n6967), .A2(n23982), .ZN(n23028) );
  INV_X1 U20511 ( .A(n39194), .ZN(n39386) );
  BUF_X2 U23052 ( .A(n10858), .Z(n15177) );
  BUF_X1 U44802 ( .A(n43059), .Z(n46060) );
  OAI21_X2 U3839 ( .B1(n31943), .B2(n31944), .A(n8330), .ZN(n35544) );
  BUF_X2 U50 ( .A(n42054), .Z(n480) );
  BUF_X1 U2914 ( .A(Key[86]), .Z(n4208) );
  BUF_X1 U5095 ( .A(Key[115]), .Z(n4721) );
  CLKBUF_X1 U2886 ( .A(Key[88]), .Z(n4823) );
  CLKBUF_X1 U3021 ( .A(Key[26]), .Z(n4353) );
  BUF_X1 U3037 ( .A(Key[31]), .Z(n2203) );
  CLKBUF_X1 U2994 ( .A(Key[67]), .Z(n4247) );
  CLKBUF_X1 U2909 ( .A(Key[0]), .Z(n4515) );
  BUF_X1 U2923 ( .A(Key[71]), .Z(n4744) );
  CLKBUF_X1 U2897 ( .A(Key[140]), .Z(n4568) );
  CLKBUF_X1 U2966 ( .A(Key[36]), .Z(n4454) );
  CLKBUF_X1 U3009 ( .A(Key[24]), .Z(n4659) );
  CLKBUF_X1 U2974 ( .A(Key[48]), .Z(n4035) );
  CLKBUF_X1 U2976 ( .A(Key[75]), .Z(n4451) );
  BUF_X1 U3004 ( .A(Key[162]), .Z(n4847) );
  CLKBUF_X1 U2888 ( .A(Key[170]), .Z(n4295) );
  CLKBUF_X1 U2989 ( .A(Key[9]), .Z(n4312) );
  CLKBUF_X1 U2982 ( .A(Key[163]), .Z(n4930) );
  CLKBUF_X1 U194 ( .A(Key[30]), .Z(n75) );
  CLKBUF_X1 U2992 ( .A(Key[85]), .Z(n4065) );
  BUF_X1 U2916 ( .A(Key[11]), .Z(n4649) );
  CLKBUF_X1 U2908 ( .A(Key[2]), .Z(n4517) );
  BUF_X1 U16689 ( .A(Key[134]), .Z(n4932) );
  CLKBUF_X1 U3019 ( .A(Key[12]), .Z(n4578) );
  CLKBUF_X1 U2904 ( .A(Key[146]), .Z(n3014) );
  CLKBUF_X1 U3032 ( .A(Key[6]), .Z(n842) );
  CLKBUF_X1 U2958 ( .A(Key[118]), .Z(n4204) );
  CLKBUF_X1 U2915 ( .A(Key[131]), .Z(n1354) );
  CLKBUF_X1 U2996 ( .A(Key[3]), .Z(n4564) );
  CLKBUF_X1 U2949 ( .A(Key[111]), .Z(n4316) );
  XNOR2_X1 U14542 ( .A(Key[177]), .B(Ciphertext[164]), .ZN(n12325) );
  CLKBUF_X1 U2930 ( .A(Key[129]), .Z(n4343) );
  CLKBUF_X1 U2902 ( .A(Key[128]), .Z(n3276) );
  BUF_X1 U2882 ( .A(n10790), .Z(n12480) );
  XNOR2_X1 U14255 ( .A(n8983), .B(Key[83]), .ZN(n9417) );
  CLKBUF_X1 U5066 ( .A(n9186), .Z(n11984) );
  XNOR2_X1 U21452 ( .A(n8989), .B(Key[186]), .ZN(n9647) );
  XNOR2_X1 U585 ( .A(n9199), .B(Key[143]), .ZN(n9203) );
  AND2_X1 U2423 ( .A1(n10143), .A2(n10147), .ZN(n10219) );
  INV_X1 U5112 ( .A(n10572), .ZN(n7185) );
  AND2_X1 U5040 ( .A1(n11393), .A2(n9384), .ZN(n10362) );
  AND2_X1 U1727 ( .A1(n10669), .A2(n12340), .ZN(n10676) );
  INV_X1 U1119 ( .A(n9647), .ZN(n12263) );
  OR2_X1 U19091 ( .A1(n12278), .A2(n9015), .ZN(n10234) );
  INV_X1 U1449 ( .A(n9056), .ZN(n12314) );
  NAND2_X1 U2869 ( .A1(n11611), .A2(n11608), .ZN(n11598) );
  AND2_X1 U4973 ( .A1(n10120), .A2(n10959), .ZN(n10054) );
  AND2_X1 U4968 ( .A1(n6465), .A2(n10361), .ZN(n10664) );
  AND2_X1 U4972 ( .A1(n6465), .A2(n9384), .ZN(n12045) );
  AND2_X1 U1427 ( .A1(n10594), .A2(n9340), .ZN(n11269) );
  AND2_X1 U21960 ( .A1(n11352), .A2(n12381), .ZN(n12097) );
  AND2_X1 U804 ( .A1(n11367), .A2(n11376), .ZN(n9636) );
  AND2_X1 U4995 ( .A1(n9142), .A2(n9932), .ZN(n9500) );
  AND2_X1 U1786 ( .A1(n11641), .A2(n10563), .ZN(n11655) );
  AND2_X1 U1765 ( .A1(n11014), .A2(n51762), .ZN(n11001) );
  NOR2_X1 U459 ( .A1(n7444), .A2(n2452), .ZN(n7443) );
  NAND4_X2 U637 ( .A1(n12365), .A2(n12368), .A3(n12367), .A4(n12366), .ZN(
        n14711) );
  NAND4_X1 U213 ( .A1(n10484), .A2(n10483), .A3(n10481), .A4(n10482), .ZN(
        n14257) );
  NOR2_X1 U1861 ( .A1(n10937), .A2(n297), .ZN(n12403) );
  AND2_X2 U1550 ( .A1(n7562), .A2(n7561), .ZN(n14318) );
  AND3_X1 U1683 ( .A1(n11677), .A2(n11678), .A3(n6181), .ZN(n11694) );
  NAND2_X1 U12446 ( .A1(n9228), .A2(n2261), .ZN(n13885) );
  OR2_X2 U6369 ( .A1(n1421), .A2(n10171), .ZN(n13148) );
  BUF_X1 U4875 ( .A(n10499), .Z(n15126) );
  INV_X1 U2828 ( .A(n14178), .ZN(n13135) );
  INV_X1 U22664 ( .A(n13131), .ZN(n13152) );
  OR2_X1 U9987 ( .A1(n13306), .A2(n13729), .ZN(n13736) );
  AND2_X1 U23396 ( .A1(n14408), .A2(n14410), .ZN(n14068) );
  OR2_X1 U4805 ( .A1(n12228), .A2(n14344), .ZN(n13006) );
  OR2_X1 U1896 ( .A1(n14285), .A2(n14287), .ZN(n13015) );
  OR2_X1 U453 ( .A1(n14311), .A2(n14317), .ZN(n13824) );
  NOR2_X1 U4775 ( .A1(n483), .A2(n2072), .ZN(n14652) );
  OR2_X1 U376 ( .A1(n13856), .A2(n13550), .ZN(n13843) );
  NOR2_X1 U22373 ( .A1(n13971), .A2(n14228), .ZN(n13214) );
  NOR2_X1 U1515 ( .A1(n14664), .A2(n13632), .ZN(n13622) );
  AOI21_X1 U869 ( .B1(n12394), .B2(n12393), .A(n14088), .ZN(n12400) );
  OR2_X1 U4692 ( .A1(n3395), .A2(n12016), .ZN(n17847) );
  NAND4_X1 U4716 ( .A1(n12025), .A2(n12024), .A3(n12026), .A4(n5732), .ZN(
        n16661) );
  NOR2_X1 U17153 ( .A1(n5344), .A2(n5343), .ZN(n15542) );
  NAND3_X1 U2439 ( .A1(n12036), .A2(n12030), .A3(n3359), .ZN(n17177) );
  OAI211_X1 U4699 ( .C1(n14483), .C2(n14482), .A(n14887), .B(n14886), .ZN(
        n18169) );
  AND3_X1 U4696 ( .A1(n8146), .A2(n13725), .A3(n8147), .ZN(n8145) );
  NAND4_X1 U963 ( .A1(n15453), .A2(n15452), .A3(n15451), .A4(n15450), .ZN(
        n17288) );
  NAND4_X1 U14865 ( .A1(n11437), .A2(n11438), .A3(n11435), .A4(n11436), .ZN(
        n16064) );
  INV_X1 U860 ( .A(n18747), .ZN(n18135) );
  BUF_X1 U2297 ( .A(n948), .Z(n484) );
  XNOR2_X1 U5467 ( .A(n15542), .B(n948), .ZN(n16781) );
  OR2_X2 U10107 ( .A1(n3083), .A2(n5190), .ZN(n19199) );
  XNOR2_X1 U1493 ( .A(n16186), .B(n49109), .ZN(n18828) );
  XNOR2_X1 U13553 ( .A(n16186), .B(n16435), .ZN(n17178) );
  XNOR2_X1 U25794 ( .A(n355), .B(n15018), .ZN(n18605) );
  XNOR2_X1 U25793 ( .A(n15017), .B(n15016), .ZN(n17522) );
  XNOR2_X1 U1464 ( .A(n19273), .B(n19272), .ZN(n20334) );
  XNOR2_X1 U20604 ( .A(n17114), .B(n17113), .ZN(n19834) );
  INV_X1 U27090 ( .A(n19141), .ZN(n16218) );
  OR2_X1 U1086 ( .A1(n18888), .A2(n19795), .ZN(n19797) );
  BUF_X1 U1241 ( .A(n51385), .Z(n19643) );
  XNOR2_X1 U4640 ( .A(n16734), .B(n16733), .ZN(n18313) );
  NAND2_X1 U7172 ( .A1(n20230), .A2(n20684), .ZN(n20678) );
  OR2_X1 U2771 ( .A1(n18313), .A2(n17059), .ZN(n20101) );
  BUF_X1 U979 ( .A(n15928), .Z(n20682) );
  INV_X1 U4603 ( .A(n17639), .ZN(n20477) );
  BUF_X2 U7639 ( .A(n21484), .Z(n2221) );
  BUF_X1 U2454 ( .A(n18357), .Z(n574) );
  CLKBUF_X1 U4597 ( .A(n15399), .Z(n19425) );
  AND2_X1 U324 ( .A1(n20638), .A2(n51485), .ZN(n20752) );
  NAND2_X1 U27428 ( .A1(n20114), .A2(n19534), .ZN(n20166) );
  AND2_X1 U4564 ( .A1(n21369), .A2(n21389), .ZN(n21398) );
  NOR2_X1 U12787 ( .A1(n5519), .A2(n18063), .ZN(n18332) );
  INV_X1 U509 ( .A(n21544), .ZN(n20738) );
  NAND2_X2 U7657 ( .A1(n51755), .A2(n21584), .ZN(n21569) );
  INV_X1 U1440 ( .A(n21494), .ZN(n20812) );
  AND2_X1 U696 ( .A1(n3370), .A2(n21654), .ZN(n16891) );
  NOR2_X1 U682 ( .A1(n19482), .A2(n19477), .ZN(n18969) );
  OR2_X1 U6491 ( .A1(n20815), .A2(n20448), .ZN(n21479) );
  AND4_X1 U260 ( .A1(n14386), .A2(n14387), .A3(n14388), .A4(n18338), .ZN(
        n14389) );
  MUX2_X1 U427 ( .A(n18339), .B(n14385), .S(n18342), .Z(n14390) );
  OAI21_X1 U28793 ( .B1(n20802), .B2(n21398), .A(n17980), .ZN(n17986) );
  NAND2_X1 U4417 ( .A1(n8717), .A2(n8703), .ZN(n21744) );
  BUF_X1 U162 ( .A(n20161), .Z(n22037) );
  OR2_X2 U15414 ( .A1(n6174), .A2(n6178), .ZN(n23981) );
  NAND3_X1 U1654 ( .A1(n267), .A2(n2453), .A3(n21192), .ZN(n23177) );
  NAND3_X1 U12878 ( .A1(n8309), .A2(n3089), .A3(n3085), .ZN(n23810) );
  INV_X1 U11421 ( .A(n20161), .ZN(n23412) );
  NAND4_X2 U17910 ( .A1(n16310), .A2(n16312), .A3(n16313), .A4(n16311), .ZN(
        n21948) );
  INV_X1 U1974 ( .A(n22144), .ZN(n22142) );
  AND2_X1 U739 ( .A1(n23157), .A2(n21948), .ZN(n23147) );
  NOR2_X1 U1211 ( .A1(n22471), .A2(n22464), .ZN(n22476) );
  NOR2_X1 U770 ( .A1(n23020), .A2(n22856), .ZN(n21880) );
  INV_X1 U4410 ( .A(n22176), .ZN(n21106) );
  INV_X1 U160 ( .A(n22946), .ZN(n23049) );
  NOR2_X1 U5356 ( .A1(n23336), .A2(n17510), .ZN(n21731) );
  OR2_X1 U1598 ( .A1(n51001), .A2(n23129), .ZN(n24119) );
  INV_X1 U563 ( .A(n24334), .ZN(n23695) );
  OR2_X1 U4356 ( .A1(n22995), .A2(n22557), .ZN(n22990) );
  AND2_X1 U806 ( .A1(n21731), .A2(n21730), .ZN(n21736) );
  AND2_X1 U20899 ( .A1(n21961), .A2(n23469), .ZN(n21966) );
  AND4_X1 U31318 ( .A1(n21815), .A2(n21817), .A3(n21816), .A4(n21814), .ZN(
        n21826) );
  AND2_X1 U608 ( .A1(n22532), .A2(n5114), .ZN(n5115) );
  NOR3_X1 U4294 ( .A1(n22396), .A2(n22395), .A3(n22394), .ZN(n22397) );
  AND3_X1 U4279 ( .A1(n20946), .A2(n20947), .A3(n2108), .ZN(n20950) );
  NAND3_X1 U144 ( .A1(n22206), .A2(n22205), .A3(n22204), .ZN(n26610) );
  NAND4_X2 U1121 ( .A1(n21787), .A2(n21790), .A3(n21788), .A4(n21789), .ZN(
        n27250) );
  NAND4_X1 U888 ( .A1(n22028), .A2(n22030), .A3(n22027), .A4(n22029), .ZN(
        n25494) );
  BUF_X1 U2081 ( .A(n27459), .Z(n370) );
  OR2_X1 U746 ( .A1(n6309), .A2(n6310), .ZN(n26425) );
  BUF_X1 U32874 ( .A(n25508), .Z(n26581) );
  XNOR2_X1 U493 ( .A(n8119), .B(n26614), .ZN(n29029) );
  CLKBUF_X1 U4197 ( .A(n23809), .Z(n30662) );
  INV_X1 U2709 ( .A(n28862), .ZN(n28951) );
  BUF_X1 U1395 ( .A(n23301), .Z(n30790) );
  BUF_X1 U2719 ( .A(n23112), .Z(n2169) );
  BUF_X1 U903 ( .A(n30718), .Z(n2205) );
  XNOR2_X1 U19632 ( .A(n7612), .B(n24875), .ZN(n7614) );
  BUF_X1 U1599 ( .A(n27783), .Z(n377) );
  BUF_X1 U7499 ( .A(n2109), .Z(n30716) );
  NAND2_X1 U1030 ( .A1(n30273), .A2(n27918), .ZN(n30263) );
  XNOR2_X1 U238 ( .A(n27343), .B(n27342), .ZN(n27379) );
  XNOR2_X1 U2333 ( .A(n26539), .B(n26538), .ZN(n28155) );
  INV_X1 U2699 ( .A(n51722), .ZN(n23658) );
  AND2_X1 U595 ( .A1(n2774), .A2(n30780), .ZN(n26828) );
  OR2_X1 U4090 ( .A1(n30707), .A2(n30721), .ZN(n30710) );
  NOR2_X1 U2712 ( .A1(n2774), .A2(n30780), .ZN(n30789) );
  OR2_X1 U11825 ( .A1(n7438), .A2(n447), .ZN(n27067) );
  BUF_X2 U2122 ( .A(n29533), .Z(n398) );
  NAND2_X1 U244 ( .A1(n27379), .A2(n30374), .ZN(n30733) );
  AND2_X1 U1298 ( .A1(n29747), .A2(n29737), .ZN(n28996) );
  NOR2_X1 U1078 ( .A1(n7909), .A2(n27783), .ZN(n28713) );
  AND2_X1 U480 ( .A1(n27056), .A2(n8455), .ZN(n29543) );
  NAND2_X1 U708 ( .A1(n626), .A2(n52165), .ZN(n29172) );
  BUF_X1 U1633 ( .A(n24984), .Z(n30245) );
  BUF_X1 U2680 ( .A(n28138), .Z(n28950) );
  CLKBUF_X1 U1470 ( .A(n26973), .Z(n29525) );
  INV_X1 U1089 ( .A(n26667), .ZN(n29496) );
  OR2_X1 U778 ( .A1(n30263), .A2(n1964), .ZN(n29233) );
  OR2_X1 U884 ( .A1(n7042), .A2(n28007), .ZN(n28568) );
  AND4_X1 U35864 ( .A1(n27969), .A2(n27970), .A3(n27971), .A4(n29240), .ZN(
        n27974) );
  AND4_X1 U3997 ( .A1(n29792), .A2(n4265), .A3(n29791), .A4(n4264), .ZN(n8738)
         );
  AND3_X1 U18237 ( .A1(n6284), .A2(n27693), .A3(n6283), .ZN(n30601) );
  AND4_X1 U1242 ( .A1(n28185), .A2(n28186), .A3(n28184), .A4(n28183), .ZN(
        n28193) );
  NAND2_X1 U12304 ( .A1(n30255), .A2(n2866), .ZN(n31558) );
  OR2_X1 U38298 ( .A1(n32402), .A2(n51519), .ZN(n32062) );
  AND4_X2 U892 ( .A1(n7335), .A2(n7336), .A3(n8185), .A4(n8184), .ZN(n29622)
         );
  BUF_X1 U2104 ( .A(n31748), .Z(n386) );
  INV_X1 U8667 ( .A(n31383), .ZN(n3241) );
  AND3_X1 U1485 ( .A1(n28706), .A2(n28707), .A3(n28705), .ZN(n232) );
  NOR2_X1 U37049 ( .A1(n32074), .A2(n32402), .ZN(n33155) );
  INV_X1 U12533 ( .A(n32876), .ZN(n33034) );
  NOR2_X1 U488 ( .A1(n32509), .A2(n31986), .ZN(n30879) );
  OR2_X2 U3906 ( .A1(n30750), .A2(n30749), .ZN(n31454) );
  NOR2_X1 U805 ( .A1(n32725), .A2(n32316), .ZN(n32318) );
  INV_X1 U2650 ( .A(n32407), .ZN(n714) );
  OR2_X1 U1136 ( .A1(n30853), .A2(n31624), .ZN(n30558) );
  OR2_X1 U3865 ( .A1(n31566), .A2(n7627), .ZN(n1890) );
  INV_X1 U394 ( .A(n31630), .ZN(n31625) );
  MUX2_X1 U2267 ( .A(n32979), .B(n32978), .S(n32977), .Z(n32995) );
  NAND4_X1 U1123 ( .A1(n30923), .A2(n30921), .A3(n30922), .A4(n30920), .ZN(
        n31923) );
  NAND4_X1 U14529 ( .A1(n5439), .A2(n5440), .A3(n30869), .A4(n30870), .ZN(
        n32310) );
  NAND4_X1 U1194 ( .A1(n31183), .A2(n31186), .A3(n31184), .A4(n31185), .ZN(
        n34412) );
  NAND4_X1 U20491 ( .A1(n30480), .A2(n2281), .A3(n8537), .A4(n8535), .ZN(
        n34594) );
  INV_X1 U418 ( .A(n33212), .ZN(n37111) );
  XNOR2_X1 U16665 ( .A(n34293), .B(n34292), .ZN(n36429) );
  XNOR2_X1 U13413 ( .A(n7126), .B(n34131), .ZN(n36571) );
  CLKBUF_X1 U1930 ( .A(n37519), .Z(n618) );
  BUF_X2 U72 ( .A(n33648), .Z(n37557) );
  CLKBUF_X1 U2615 ( .A(n36772), .Z(n39019) );
  XNOR2_X1 U242 ( .A(n36816), .B(n36815), .ZN(n37901) );
  CLKBUF_X1 U2289 ( .A(n36105), .Z(n481) );
  OR2_X1 U1106 ( .A1(n34908), .A2(n1698), .ZN(n39393) );
  AND2_X1 U65 ( .A1(n34984), .A2(n37974), .ZN(n37977) );
  AND2_X1 U1438 ( .A1(n34908), .A2(n1698), .ZN(n39397) );
  OR2_X1 U748 ( .A1(n4512), .A2(n38270), .ZN(n38290) );
  INV_X1 U2610 ( .A(n39272), .ZN(n39258) );
  AND2_X1 U1216 ( .A1(n39258), .A2(n8429), .ZN(n2571) );
  AND2_X1 U6876 ( .A1(n36312), .A2(n38094), .ZN(n38073) );
  BUF_X1 U2485 ( .A(n5711), .Z(n594) );
  NOR2_X1 U7110 ( .A1(n5711), .A2(n37983), .ZN(n36522) );
  AND2_X1 U9597 ( .A1(n39234), .A2(n3874), .ZN(n4674) );
  AOI21_X1 U1417 ( .B1(n38734), .B2(n8077), .A(n222), .ZN(n6150) );
  NOR3_X1 U1667 ( .A1(n35169), .A2(n38557), .A3(n5846), .ZN(n38542) );
  AND4_X1 U3577 ( .A1(n37029), .A2(n37030), .A3(n37027), .A4(n37028), .ZN(
        n37034) );
  NAND3_X1 U492 ( .A1(n2887), .A2(n34645), .A3(n34643), .ZN(n41079) );
  NAND4_X2 U16616 ( .A1(n38208), .A2(n38209), .A3(n38207), .A4(n38206), .ZN(
        n40972) );
  AND4_X2 U17690 ( .A1(n37412), .A2(n5806), .A3(n5805), .A4(n37413), .ZN(
        n40778) );
  AND2_X1 U355 ( .A1(n34805), .A2(n34803), .ZN(n1) );
  AND4_X1 U1294 ( .A1(n37700), .A2(n37703), .A3(n37699), .A4(n3734), .ZN(n7697) );
  AND2_X2 U5911 ( .A1(n7697), .A2(n37705), .ZN(n40822) );
  AND2_X1 U8749 ( .A1(n36009), .A2(n36008), .ZN(n4070) );
  NOR2_X1 U5965 ( .A1(n41083), .A2(n41079), .ZN(n39707) );
  OR2_X1 U1547 ( .A1(n35203), .A2(n35202), .ZN(n39103) );
  OR2_X1 U568 ( .A1(n7848), .A2(n40565), .ZN(n40315) );
  INV_X1 U13710 ( .A(n41489), .ZN(n42049) );
  NOR2_X1 U3488 ( .A1(n40609), .A2(n41647), .ZN(n41986) );
  AND2_X1 U1487 ( .A1(n6617), .A2(n41939), .ZN(n233) );
  OR2_X1 U1409 ( .A1(n41356), .A2(n41355), .ZN(n41342) );
  INV_X1 U1697 ( .A(n2855), .ZN(n40450) );
  OR2_X1 U998 ( .A1(n431), .A2(n40785), .ZN(n40067) );
  AND2_X1 U7376 ( .A1(n610), .A2(n2016), .ZN(n41053) );
  NAND4_X1 U41926 ( .A1(n37348), .A2(n37349), .A3(n37351), .A4(n37350), .ZN(
        n44879) );
  NAND4_X1 U12351 ( .A1(n41092), .A2(n41091), .A3(n41090), .A4(n41089), .ZN(
        n41956) );
  NAND2_X1 U1100 ( .A1(n4187), .A2(n41990), .ZN(n44176) );
  BUF_X1 U7616 ( .A(n45101), .Z(n2206) );
  CLKBUF_X1 U2445 ( .A(n44972), .Z(n569) );
  XNOR2_X1 U13561 ( .A(n7005), .B(n43519), .ZN(n6172) );
  BUF_X1 U2167 ( .A(n50382), .Z(n423) );
  XNOR2_X1 U14650 ( .A(n43260), .B(n43259), .ZN(n49662) );
  XNOR2_X1 U46506 ( .A(n44228), .B(n44227), .ZN(n46322) );
  XOR2_X1 U7486 ( .A(n44519), .B(n7900), .Z(n2104) );
  INV_X2 U3340 ( .A(n43797), .ZN(n667) );
  INV_X1 U2546 ( .A(n45560), .ZN(n48505) );
  AND2_X1 U3292 ( .A1(n48201), .A2(n48213), .ZN(n45540) );
  BUF_X1 U2024 ( .A(n50350), .Z(n555) );
  AND2_X1 U2143 ( .A1(n46597), .A2(n45793), .ZN(n46587) );
  INV_X1 U2541 ( .A(n45793), .ZN(n46714) );
  OR2_X1 U18114 ( .A1(n52039), .A2(n46322), .ZN(n46318) );
  NOR2_X1 U5726 ( .A1(n51344), .A2(n50965), .ZN(n46740) );
  AND2_X1 U16041 ( .A1(n46648), .A2(n46844), .ZN(n46840) );
  CLKBUF_X1 U2124 ( .A(n47078), .Z(n399) );
  AND2_X1 U693 ( .A1(n49939), .A2(n50292), .ZN(n50307) );
  NOR2_X1 U1726 ( .A1(n47288), .A2(n50344), .ZN(n49961) );
  AND2_X1 U3219 ( .A1(n3108), .A2(n46589), .ZN(n44845) );
  AND2_X1 U985 ( .A1(n45773), .A2(n46844), .ZN(n46860) );
  AND2_X1 U830 ( .A1(n45773), .A2(n3892), .ZN(n47129) );
  AND2_X1 U3193 ( .A1(n48543), .A2(n45634), .ZN(n48242) );
  AND4_X1 U5207 ( .A1(n50271), .A2(n50273), .A3(n50274), .A4(n50272), .ZN(
        n50286) );
  OR2_X1 U3174 ( .A1(n46768), .A2(n46769), .ZN(n6570) );
  AND3_X2 U1107 ( .A1(n44619), .A2(n49971), .A3(n44620), .ZN(n50727) );
  NOR2_X1 U1279 ( .A1(n49606), .A2(n49599), .ZN(n49574) );
  BUF_X1 U2435 ( .A(n50115), .Z(n562) );
  INV_X1 U318 ( .A(n48365), .ZN(n48382) );
  OR2_X1 U18892 ( .A1(n1501), .A2(n49114), .ZN(n44798) );
  AND2_X1 U477 ( .A1(n49706), .A2(n49644), .ZN(n49823) );
  BUF_X1 U2901 ( .A(Key[122]), .Z(n2183) );
  CLKBUF_X1 U3006 ( .A(Key[156]), .Z(n4482) );
  CLKBUF_X1 U2940 ( .A(Key[27]), .Z(n4045) );
  CLKBUF_X1 U5083 ( .A(Key[153]), .Z(n4638) );
  CLKBUF_X1 U2951 ( .A(Key[70]), .Z(n4845) );
  CLKBUF_X1 U3016 ( .A(Key[56]), .Z(n48597) );
  INV_X1 U21565 ( .A(n11590), .ZN(n11601) );
  INV_X1 U21517 ( .A(n12325), .ZN(n10669) );
  INV_X1 U21846 ( .A(n10065), .ZN(n10069) );
  BUF_X1 U2059 ( .A(n11136), .Z(n357) );
  INV_X2 U1145 ( .A(n10527), .ZN(n9482) );
  NAND2_X1 U2865 ( .A1(n12470), .A2(n12480), .ZN(n12478) );
  INV_X1 U21286 ( .A(n11485), .ZN(n12481) );
  NAND2_X2 U13101 ( .A1(n3250), .A2(n10816), .ZN(n11600) );
  NAND2_X2 U959 ( .A1(n12663), .A2(n9188), .ZN(n11973) );
  NAND2_X2 U560 ( .A1(n12282), .A2(n12280), .ZN(n10715) );
  INV_X1 U1894 ( .A(n13822), .ZN(n13826) );
  INV_X2 U1895 ( .A(n13779), .ZN(n12419) );
  INV_X2 U968 ( .A(n14234), .ZN(n16221) );
  INV_X1 U4826 ( .A(n15425), .ZN(n1556) );
  BUF_X1 U2830 ( .A(n11293), .Z(n12963) );
  NAND2_X2 U6239 ( .A1(n10898), .A2(n10899), .ZN(n13782) );
  INV_X2 U1626 ( .A(n51670), .ZN(n14717) );
  AND3_X1 U2288 ( .A1(n7371), .A2(n14676), .A3(n14675), .ZN(n15014) );
  BUF_X1 U2418 ( .A(n16373), .Z(n557) );
  INV_X1 U9158 ( .A(n21181), .ZN(n17201) );
  INV_X1 U25849 ( .A(n17522), .ZN(n20021) );
  INV_X1 U25512 ( .A(n20478), .ZN(n20466) );
  XNOR2_X1 U333 ( .A(n17946), .B(n17945), .ZN(n20376) );
  INV_X2 U2786 ( .A(n20326), .ZN(n21424) );
  XNOR2_X1 U29163 ( .A(n18493), .B(n18492), .ZN(n20642) );
  AND2_X2 U4578 ( .A1(n19671), .A2(n51006), .ZN(n20217) );
  XNOR2_X1 U14775 ( .A(n16263), .B(n16262), .ZN(n17081) );
  NAND2_X1 U12156 ( .A1(n2773), .A2(n20244), .ZN(n5541) );
  BUF_X2 U4585 ( .A(n17195), .Z(n19826) );
  AND2_X1 U510 ( .A1(n20627), .A2(n18495), .ZN(n21544) );
  NAND2_X1 U17943 ( .A1(n21495), .A2(n2221), .ZN(n20811) );
  NAND2_X1 U7171 ( .A1(n5373), .A2(n20678), .ZN(n18875) );
  NAND2_X1 U7090 ( .A1(n19820), .A2(n19822), .ZN(n21196) );
  INV_X2 U1584 ( .A(n21744), .ZN(n629) );
  INV_X1 U1911 ( .A(n23314), .ZN(n23310) );
  INV_X1 U10312 ( .A(n22989), .ZN(n22985) );
  NOR2_X1 U2751 ( .A1(n23827), .A2(n3520), .ZN(n23834) );
  INV_X1 U14267 ( .A(n22521), .ZN(n23143) );
  INV_X1 U9202 ( .A(n24034), .ZN(n24025) );
  INV_X1 U9181 ( .A(n23171), .ZN(n23183) );
  INV_X1 U7991 ( .A(n21756), .ZN(n22262) );
  AND2_X2 U1693 ( .A1(n8205), .A2(n1648), .ZN(n22275) );
  INV_X1 U2752 ( .A(n24000), .ZN(n23983) );
  INV_X2 U7169 ( .A(n22287), .ZN(n22701) );
  INV_X1 U6285 ( .A(n24211), .ZN(n23066) );
  NOR2_X2 U1350 ( .A1(n6167), .A2(n21782), .ZN(n21778) );
  XNOR2_X1 U9317 ( .A(n24795), .B(n28352), .ZN(n27477) );
  XNOR2_X1 U2203 ( .A(n25029), .B(n22973), .ZN(n25934) );
  INV_X1 U32863 ( .A(n30769), .ZN(n30771) );
  XNOR2_X1 U277 ( .A(n25491), .B(n24940), .ZN(n30248) );
  XNOR2_X1 U889 ( .A(n23108), .B(n25965), .ZN(n28809) );
  INV_X1 U33183 ( .A(n29413), .ZN(n26989) );
  INV_X1 U4208 ( .A(n30171), .ZN(n1771) );
  INV_X1 U307 ( .A(n27668), .ZN(n2642) );
  INV_X1 U1921 ( .A(n29278), .ZN(n28715) );
  INV_X1 U2646 ( .A(n30912), .ZN(n30602) );
  INV_X2 U6575 ( .A(n1428), .ZN(n7430) );
  INV_X1 U8608 ( .A(n30873), .ZN(n32004) );
  INV_X1 U37439 ( .A(n31377), .ZN(n33002) );
  NOR2_X2 U1722 ( .A1(n31369), .A2(n711), .ZN(n32300) );
  INV_X2 U2622 ( .A(n38275), .ZN(n38272) );
  INV_X1 U280 ( .A(n38630), .ZN(n38637) );
  INV_X1 U6376 ( .A(n35923), .ZN(n37750) );
  BUF_X1 U374 ( .A(n39272), .Z(n551) );
  INV_X1 U3766 ( .A(n38659), .ZN(n700) );
  INV_X1 U8127 ( .A(n36248), .ZN(n3650) );
  INV_X2 U1447 ( .A(n39464), .ZN(n39035) );
  NAND2_X2 U619 ( .A1(n36029), .A2(n34090), .ZN(n36542) );
  AND2_X1 U1142 ( .A1(n37901), .A2(n38946), .ZN(n39423) );
  INV_X1 U7833 ( .A(n35010), .ZN(n38146) );
  AND2_X1 U1313 ( .A1(n51102), .A2(n39195), .ZN(n39367) );
  INV_X1 U2422 ( .A(n39834), .ZN(n677) );
  INV_X1 U2587 ( .A(n43327), .ZN(n41008) );
  INV_X1 U3487 ( .A(n41581), .ZN(n42010) );
  INV_X1 U16724 ( .A(n4954), .ZN(n4950) );
  INV_X1 U2534 ( .A(n49662), .ZN(n6116) );
  NAND2_X1 U13014 ( .A1(n46591), .A2(n46708), .ZN(n46580) );
  INV_X1 U11031 ( .A(n43798), .ZN(n50370) );
  INV_X1 U45110 ( .A(n48462), .ZN(n46448) );
  INV_X1 U306 ( .A(n46519), .ZN(n46511) );
  INV_X2 U44623 ( .A(n41908), .ZN(n48200) );
  INV_X1 U2514 ( .A(n50486), .ZN(n7114) );
  INV_X1 U3160 ( .A(n49070), .ZN(n1502) );
  INV_X2 U11181 ( .A(n2192), .ZN(n49510) );
  NAND2_X1 U1834 ( .A1(n49443), .A2(n49445), .ZN(n49461) );
  AND4_X2 U2428 ( .A1(n5544), .A2(n26073), .A3(n5545), .A4(n26072), .ZN(n1685)
         );
  NAND4_X2 U12514 ( .A1(n12930), .A2(n12931), .A3(n12929), .A4(n12928), .ZN(
        n16743) );
  BUF_X2 U1517 ( .A(n45995), .Z(n49707) );
  NOR2_X2 U309 ( .A1(n49793), .A2(n49862), .ZN(n49829) );
  INV_X2 U2744 ( .A(n22129), .ZN(n22658) );
  AND3_X2 U3547 ( .A1(n39188), .A2(n39187), .A3(n39186), .ZN(n41238) );
  NAND2_X2 U14920 ( .A1(n10423), .A2(n10428), .ZN(n11943) );
  OR2_X2 U880 ( .A1(n8044), .A2(n31275), .ZN(n35085) );
  NAND4_X2 U36210 ( .A1(n28477), .A2(n28476), .A3(n28475), .A4(n28474), .ZN(
        n34546) );
  XNOR2_X2 U2437 ( .A(n16294), .B(n18689), .ZN(n16658) );
  OR2_X2 U1315 ( .A1(n6715), .A2(n28527), .ZN(n32327) );
  NOR2_X2 U358 ( .A1(n8291), .A2(n41029), .ZN(n41025) );
  OR2_X2 U1631 ( .A1(n5037), .A2(n36133), .ZN(n38152) );
  OR2_X2 U1188 ( .A1(n668), .A2(n48180), .ZN(n48166) );
  NAND2_X2 U15918 ( .A1(n13543), .A2(n13544), .ZN(n21780) );
  BUF_X2 U40660 ( .A(n35406), .Z(n36468) );
  NAND2_X2 U13913 ( .A1(n36029), .A2(n36547), .ZN(n37964) );
  OR2_X2 U1634 ( .A1(n47044), .A2(n47341), .ZN(n47335) );
  BUF_X2 U3327 ( .A(n42883), .Z(n49397) );
  OR2_X2 U1185 ( .A1(n40862), .A2(n40868), .ZN(n5747) );
  NAND2_X2 U14604 ( .A1(n29597), .A2(n4059), .ZN(n33195) );
  XNOR2_X2 U4688 ( .A(n16919), .B(n18443), .ZN(n15519) );
  AND3_X2 U2326 ( .A1(n45627), .A2(n45626), .A3(n45625), .ZN(n48853) );
  OR2_X2 U19560 ( .A1(n26465), .A2(n26464), .ZN(n30534) );
  INV_X2 U2739 ( .A(n22386), .ZN(n5371) );
  AND4_X2 U4724 ( .A1(n14438), .A2(n14439), .A3(n14437), .A4(n14436), .ZN(
        n14462) );
  NAND2_X2 U18464 ( .A1(n15465), .A2(n15464), .ZN(n21767) );
  OR2_X2 U13536 ( .A1(n23410), .A2(n20890), .ZN(n23408) );
  INV_X2 U1760 ( .A(n41702), .ZN(n41697) );
  INV_X2 U11995 ( .A(n18519), .ZN(n16720) );
  AND4_X2 U14871 ( .A1(n7281), .A2(n7280), .A3(n7284), .A4(n2437), .ZN(n6481)
         );
  OR2_X2 U1452 ( .A1(n22479), .A2(n22306), .ZN(n21130) );
  NAND4_X2 U2586 ( .A1(n5327), .A2(n4474), .A3(n33176), .A4(n33177), .ZN(
        n39834) );
  AND2_X2 U532 ( .A1(n95), .A2(n29501), .ZN(n30925) );
  AND2_X2 U15331 ( .A1(n15206), .A2(n14767), .ZN(n15235) );
  OR2_X2 U13317 ( .A1(n26770), .A2(n26769), .ZN(n29998) );
  OR2_X2 U1740 ( .A1(n5199), .A2(n28333), .ZN(n30434) );
  BUF_X2 U2361 ( .A(n15851), .Z(n511) );
  NOR2_X2 U900 ( .A1(n10765), .A2(n7195), .ZN(n14239) );
  AND2_X2 U695 ( .A1(n21652), .A2(n20658), .ZN(n21654) );
  BUF_X2 U2557 ( .A(n42685), .Z(n44752) );
  NOR2_X2 U957 ( .A1(n22832), .A2(n22826), .ZN(n22503) );
  AND4_X2 U1817 ( .A1(n3618), .A2(n3620), .A3(n3617), .A4(n3613), .ZN(n14106)
         );
  AND2_X2 U1653 ( .A1(n38694), .A2(n38695), .ZN(n41352) );
  INV_X2 U2654 ( .A(n32559), .ZN(n32566) );
  NOR2_X2 U5648 ( .A1(n1050), .A2(n6607), .ZN(n32559) );
  XNOR2_X2 U17259 ( .A(n36696), .B(n36695), .ZN(n39273) );
  BUF_X2 U21099 ( .A(n50744), .Z(n50751) );
  NAND2_X2 U4708 ( .A1(n4717), .A2(n12941), .ZN(n17906) );
  XNOR2_X2 U5076 ( .A(n8800), .B(Key[70]), .ZN(n10055) );
  BUF_X2 U2465 ( .A(n21392), .Z(n581) );
  OR2_X2 U1535 ( .A1(n41117), .A2(n39600), .ZN(n43928) );
  NAND3_X2 U2804 ( .A1(n4326), .A2(n4146), .A3(n9533), .ZN(n16904) );
  OR2_X2 U15524 ( .A1(n15380), .A2(n787), .ZN(n15363) );
  BUF_X2 U2094 ( .A(n31545), .Z(n381) );
  OR2_X2 U16742 ( .A1(n4967), .A2(n34649), .ZN(n36606) );
  BUF_X2 U3255 ( .A(n44985), .Z(n46614) );
  NAND4_X2 U1766 ( .A1(n8873), .A2(n8875), .A3(n8874), .A4(n8876), .ZN(n13683)
         );
  BUF_X2 U2127 ( .A(n29930), .Z(n402) );
  XNOR2_X2 U7076 ( .A(n33113), .B(n329), .ZN(n38040) );
  NOR2_X2 U16597 ( .A1(n660), .A2(n48273), .ZN(n45590) );
  AND2_X2 U3075 ( .A1(n7139), .A2(n50486), .ZN(n50458) );
  XNOR2_X2 U42124 ( .A(n42659), .B(n42907), .ZN(n44207) );
  NAND3_X2 U1595 ( .A1(n259), .A2(n7479), .A3(n258), .ZN(n33711) );
  AND3_X2 U15350 ( .A1(n4344), .A2(n4441), .A3(n10411), .ZN(n15185) );
  BUF_X2 U2213 ( .A(n7558), .Z(n444) );
  BUF_X2 U1673 ( .A(n14738), .Z(n19370) );
  BUF_X2 U1371 ( .A(n27379), .Z(n30379) );
  XNOR2_X2 U14852 ( .A(n4154), .B(n17739), .ZN(n20493) );
  NOR2_X2 U7534 ( .A1(n30931), .A2(n29642), .ZN(n30936) );
  AND2_X2 U1671 ( .A1(n5473), .A2(n8882), .ZN(n10431) );
  NAND2_X2 U1548 ( .A1(n4785), .A2(n5123), .ZN(n35059) );
  AND2_X2 U8731 ( .A1(n37885), .A2(n3735), .ZN(n37892) );
  NAND2_X2 U1421 ( .A1(n6379), .A2(n11459), .ZN(n15380) );
  NAND3_X2 U3388 ( .A1(n3463), .A2(n38610), .A3(n38609), .ZN(n44190) );
  BUF_X2 U2304 ( .A(n30426), .Z(n487) );
  NAND4_X2 U4919 ( .A1(n6444), .A2(n6443), .A3(n6446), .A4(n9025), .ZN(n13822)
         );
  NAND3_X2 U3810 ( .A1(n2449), .A2(n32550), .A3(n4234), .ZN(n37303) );
  AND2_X2 U3191 ( .A1(n45652), .A2(n45651), .ZN(n5691) );
  AND2_X2 U3164 ( .A1(n49747), .A2(n49748), .ZN(n49854) );
  BUF_X2 U3306 ( .A(n42606), .Z(n45697) );
  NAND3_X2 U296 ( .A1(n5899), .A2(n5900), .A3(n40206), .ZN(n43920) );
  XNOR2_X2 U3801 ( .A(n36841), .B(n35512), .ZN(n34471) );
  OR2_X2 U1630 ( .A1(n38005), .A2(n38018), .ZN(n38190) );
  BUF_X2 U950 ( .A(n9074), .Z(n11613) );
  AND3_X2 U1887 ( .A1(n16580), .A2(n16581), .A3(n5455), .ZN(n21945) );
  BUF_X2 U21645 ( .A(n9139), .Z(n11209) );
  XNOR2_X2 U6208 ( .A(Key[152]), .B(Ciphertext[37]), .ZN(n8881) );
  NAND2_X2 U40789 ( .A1(n38514), .A2(n37489), .ZN(n38517) );
  AND4_X2 U1876 ( .A1(n28756), .A2(n28754), .A3(n28755), .A4(n28753), .ZN(
        n5977) );
  XNOR2_X2 U20858 ( .A(n18430), .B(n17127), .ZN(n16707) );
  OR3_X2 U10 ( .A1(n5288), .A2(n44606), .A3(n44605), .ZN(n50681) );
  AND2_X2 U3686 ( .A1(n37587), .A2(n37591), .ZN(n37592) );
  AND2_X2 U2025 ( .A1(n6741), .A2(n44652), .ZN(n45763) );
  NOR2_X2 U9999 ( .A1(n14664), .A2(n11315), .ZN(n12952) );
  AND2_X2 U3478 ( .A1(n41671), .A2(n4400), .ZN(n41227) );
  AND3_X2 U17708 ( .A1(n17538), .A2(n17540), .A3(n17539), .ZN(n22145) );
  XNOR2_X2 U17122 ( .A(n43214), .B(n43215), .ZN(n46028) );
  OR2_X2 U473 ( .A1(n28543), .A2(n28544), .ZN(n32691) );
  XNOR2_X2 U2484 ( .A(n27224), .B(n24047), .ZN(n28410) );
  BUF_X1 U7504 ( .A(n9124), .Z(n11582) );
  BUF_X1 U2881 ( .A(n8871), .Z(n12470) );
  NAND2_X1 U7889 ( .A1(n11035), .A2(n10008), .ZN(n10578) );
  BUF_X1 U1335 ( .A(n11723), .Z(n16044) );
  OR2_X1 U298 ( .A1(n13322), .A2(n14605), .ZN(n14010) );
  INV_X1 U13487 ( .A(n19868), .ZN(n19647) );
  AND2_X1 U707 ( .A1(n19482), .A2(n21248), .ZN(n21253) );
  NAND3_X1 U13310 ( .A1(n3333), .A2(n21333), .A3(n21332), .ZN(n25047) );
  NOR2_X1 U15457 ( .A1(n20719), .A2(n20718), .ZN(n22973) );
  NAND2_X1 U16040 ( .A1(n28882), .A2(n28870), .ZN(n29032) );
  OR2_X1 U1767 ( .A1(n30280), .A2(n24878), .ZN(n30292) );
  INV_X1 U4119 ( .A(n30461), .ZN(n29737) );
  INV_X1 U10590 ( .A(n31311), .ZN(n30824) );
  NAND4_X1 U2156 ( .A1(n29957), .A2(n31123), .A3(n29956), .A4(n29955), .ZN(
        n36764) );
  NAND4_X1 U430 ( .A1(n29610), .A2(n29612), .A3(n5680), .A4(n29611), .ZN(
        n36671) );
  AND2_X1 U37891 ( .A1(n51524), .A2(n31355), .ZN(n38214) );
  AND2_X1 U16220 ( .A1(n38732), .A2(n39299), .ZN(n38314) );
  AND2_X1 U1944 ( .A1(n40525), .A2(n6525), .ZN(n40873) );
  AND2_X1 U1681 ( .A1(n41083), .A2(n8316), .ZN(n41077) );
  OR2_X1 U265 ( .A1(n40119), .A2(n51352), .ZN(n40113) );
  INV_X1 U2532 ( .A(n46730), .ZN(n46753) );
  OR2_X1 U43627 ( .A1(n45589), .A2(n48259), .ZN(n48267) );
  AND2_X1 U5539 ( .A1(n2688), .A2(n988), .ZN(n46494) );
  INV_X1 U21 ( .A(n48213), .ZN(n45538) );
  AND2_X1 U19 ( .A1(n49707), .A2(n49710), .ZN(n45898) );
  NOR2_X2 U45945 ( .A1(n43486), .A2(n43485), .ZN(n49503) );
  NOR2_X2 U6 ( .A1(n48392), .A2(n8104), .ZN(n48369) );
  AND2_X1 U8916 ( .A1(n649), .A2(n50708), .ZN(n50728) );
  AND2_X1 U12 ( .A1(n51515), .A2(n46288), .ZN(n46292) );
  BUF_X1 U28 ( .A(n46519), .Z(n51068) );
  NAND4_X1 U29 ( .A1(n39498), .A2(n39496), .A3(n39495), .A4(n39497), .ZN(
        n45354) );
  OAI21_X2 U57 ( .B1(n40256), .B2(n42201), .A(n40255), .ZN(n44130) );
  AND4_X2 U79 ( .A1(n7404), .A2(n7405), .A3(n39006), .A4(n7406), .ZN(n41690)
         );
  OR2_X1 U95 ( .A1(n6869), .A2(n38565), .ZN(n38572) );
  BUF_X1 U96 ( .A(n36035), .Z(n51077) );
  XNOR2_X1 U116 ( .A(n32606), .B(n32605), .ZN(n34611) );
  AND2_X1 U134 ( .A1(n32608), .A2(n7064), .ZN(n31566) );
  OR2_X1 U137 ( .A1(n32251), .A2(n32252), .ZN(n32247) );
  AND2_X1 U139 ( .A1(n2956), .A2(n51110), .ZN(n29495) );
  NAND3_X1 U154 ( .A1(n7219), .A2(n7221), .A3(n7220), .ZN(n50990) );
  AND2_X1 U156 ( .A1(n19647), .A2(n19648), .ZN(n19848) );
  BUF_X1 U180 ( .A(n19868), .Z(n51039) );
  OR2_X1 U227 ( .A1(n13089), .A2(n13102), .ZN(n13104) );
  INV_X1 U252 ( .A(n11496), .ZN(n12675) );
  AND2_X2 U255 ( .A1(n23052), .A2(n23054), .ZN(n22943) );
  OR2_X2 U257 ( .A1(n49119), .A2(n49126), .ZN(n49101) );
  OAI211_X2 U327 ( .C1(n5064), .C2(n5063), .A(n5062), .B(n5059), .ZN(n51406)
         );
  XNOR2_X2 U362 ( .A(n44134), .B(n43155), .ZN(n42822) );
  OR2_X2 U372 ( .A1(n49274), .A2(n5783), .ZN(n49265) );
  BUF_X1 U412 ( .A(n15167), .Z(n51452) );
  INV_X2 U479 ( .A(n48792), .ZN(n48808) );
  NAND4_X2 U487 ( .A1(n39152), .A2(n39153), .A3(n39151), .A4(n39150), .ZN(
        n44501) );
  AND2_X2 U508 ( .A1(n22462), .A2(n22464), .ZN(n22721) );
  AND4_X2 U513 ( .A1(n48447), .A2(n48446), .A3(n48445), .A4(n48444), .ZN(
        n51382) );
  OR2_X2 U543 ( .A1(n28916), .A2(n28926), .ZN(n28915) );
  AND4_X2 U550 ( .A1(n19366), .A2(n19367), .A3(n19368), .A4(n19369), .ZN(
        n22329) );
  NAND2_X2 U559 ( .A1(n8633), .A2(n878), .ZN(n35255) );
  NAND4_X2 U566 ( .A1(n22613), .A2(n22612), .A3(n22610), .A4(n22611), .ZN(
        n27382) );
  XNOR2_X2 U594 ( .A(n23880), .B(n23879), .ZN(n28242) );
  AND3_X2 U599 ( .A1(n5556), .A2(n39218), .A3(n39217), .ZN(n41245) );
  BUF_X2 U633 ( .A(n34544), .Z(n376) );
  XNOR2_X1 U662 ( .A(n45304), .B(n46042), .ZN(n45454) );
  NAND2_X1 U664 ( .A1(n29346), .A2(n967), .ZN(n30210) );
  INV_X1 U683 ( .A(n24180), .ZN(n23756) );
  INV_X1 U684 ( .A(n43490), .ZN(n49539) );
  INV_X1 U694 ( .A(n50553), .ZN(n50564) );
  NAND2_X1 U714 ( .A1(n32509), .A2(n31986), .ZN(n32500) );
  INV_X1 U717 ( .A(n41685), .ZN(n41234) );
  BUF_X1 U724 ( .A(n36306), .Z(n51524) );
  INV_X1 U725 ( .A(n41323), .ZN(n41317) );
  INV_X1 U726 ( .A(n41083), .ZN(n39713) );
  NAND2_X1 U743 ( .A1(n39350), .A2(n37781), .ZN(n36186) );
  AND2_X2 U758 ( .A1(n20050), .A2(n20051), .ZN(n452) );
  NAND4_X2 U794 ( .A1(n39572), .A2(n39574), .A3(n39573), .A4(n39571), .ZN(
        n51398) );
  NAND2_X2 U795 ( .A1(n4083), .A2(n38194), .ZN(n40967) );
  NAND3_X2 U800 ( .A1(n3435), .A2(n36357), .A3(n3434), .ZN(n39767) );
  NAND4_X2 U814 ( .A1(n41070), .A2(n41069), .A3(n41068), .A4(n41067), .ZN(
        n44153) );
  INV_X2 U817 ( .A(n49990), .ZN(n47360) );
  XOR2_X1 U821 ( .A(n41757), .B(n41756), .Z(n50965) );
  OR2_X2 U832 ( .A1(n3890), .A2(n3887), .ZN(n50950) );
  AND3_X2 U833 ( .A1(n46195), .A2(n8473), .A3(n46194), .ZN(n49029) );
  NOR2_X2 U843 ( .A1(n1981), .A2(n486), .ZN(n29869) );
  NAND2_X1 U847 ( .A1(n9228), .A2(n2261), .ZN(n50966) );
  INV_X1 U859 ( .A(n13885), .ZN(n7245) );
  INV_X1 U865 ( .A(n13590), .ZN(n13583) );
  NAND4_X1 U871 ( .A1(n4740), .A2(n40392), .A3(n40391), .A4(n40390), .ZN(
        n45459) );
  INV_X2 U872 ( .A(n22488), .ZN(n22462) );
  NAND4_X1 U894 ( .A1(n26482), .A2(n26479), .A3(n26480), .A4(n26481), .ZN(
        n31377) );
  NAND3_X2 U916 ( .A1(n14301), .A2(n14302), .A3(n51269), .ZN(n18599) );
  NAND2_X2 U929 ( .A1(n35898), .A2(n5738), .ZN(n39907) );
  OAI211_X2 U930 ( .C1(n43459), .C2(n43458), .A(n43457), .B(n2802), .ZN(n2192)
         );
  OR2_X2 U936 ( .A1(n30296), .A2(n30283), .ZN(n28560) );
  CLKBUF_X1 U954 ( .A(n21063), .Z(n50976) );
  AOI21_X1 U960 ( .B1(n19741), .B2(n19740), .A(n19739), .ZN(n21063) );
  BUF_X2 U978 ( .A(n31768), .Z(n50981) );
  NAND2_X1 U982 ( .A1(n24890), .A2(n24889), .ZN(n31768) );
  XNOR2_X1 U1000 ( .A(n5234), .B(n34412), .ZN(n37020) );
  XNOR2_X1 U1002 ( .A(n33269), .B(n33268), .ZN(n38084) );
  NAND4_X1 U1016 ( .A1(n26704), .A2(n26701), .A3(n26702), .A4(n26703), .ZN(
        n31040) );
  NAND2_X2 U1060 ( .A1(n38151), .A2(n38150), .ZN(n41374) );
  NAND3_X1 U1063 ( .A1(n7219), .A2(n7221), .A3(n7220), .ZN(n23706) );
  XNOR2_X2 U1065 ( .A(n17711), .B(n17710), .ZN(n20314) );
  NAND4_X1 U1077 ( .A1(n6359), .A2(n6360), .A3(n6358), .A4(n6361), .ZN(n21925)
         );
  CLKBUF_X1 U1108 ( .A(n11496), .Z(n50997) );
  XNOR2_X1 U1110 ( .A(Key[147]), .B(Ciphertext[50]), .ZN(n11496) );
  NAND4_X2 U1122 ( .A1(n12784), .A2(n12783), .A3(n12782), .A4(n12781), .ZN(
        n16016) );
  XNOR2_X1 U1156 ( .A(n42475), .B(n43828), .ZN(n48462) );
  NAND3_X1 U1161 ( .A1(n21588), .A2(n94), .A3(n21587), .ZN(n51001) );
  CLKBUF_X1 U1183 ( .A(n12325), .Z(n51004) );
  XNOR2_X1 U1196 ( .A(n4506), .B(n15722), .ZN(n51521) );
  XNOR2_X2 U1198 ( .A(n9214), .B(Key[181]), .ZN(n12057) );
  NAND4_X1 U1245 ( .A1(n5119), .A2(n5115), .A3(n5117), .A4(n5642), .ZN(n28358)
         );
  NAND4_X1 U1261 ( .A1(n31361), .A2(n2948), .A3(n31362), .A4(n31360), .ZN(
        n41149) );
  BUF_X1 U1280 ( .A(n5668), .Z(n51016) );
  CLKBUF_X1 U1282 ( .A(n5668), .Z(n51017) );
  XNOR2_X1 U1284 ( .A(n43312), .B(n43311), .ZN(n5668) );
  NAND2_X2 U1290 ( .A1(n31900), .A2(n31901), .ZN(n35095) );
  NAND2_X1 U1303 ( .A1(n419), .A2(n2066), .ZN(n39176) );
  OR2_X2 U1311 ( .A1(n37924), .A2(n419), .ZN(n38667) );
  BUF_X2 U1326 ( .A(n16037), .Z(n51019) );
  NAND2_X1 U1327 ( .A1(n11694), .A2(n11693), .ZN(n16037) );
  XNOR2_X2 U1347 ( .A(n16666), .B(n17280), .ZN(n18697) );
  XNOR2_X1 U1356 ( .A(n15490), .B(n15489), .ZN(n20501) );
  NAND4_X2 U1358 ( .A1(n18099), .A2(n18098), .A3(n21101), .A4(n18097), .ZN(
        n25161) );
  NAND3_X1 U1359 ( .A1(n1739), .A2(n36650), .A3(n1742), .ZN(n51022) );
  AND2_X2 U1372 ( .A1(n51219), .A2(n8497), .ZN(n14137) );
  NAND4_X2 U1378 ( .A1(n31861), .A2(n31858), .A3(n31860), .A4(n31859), .ZN(
        n33550) );
  NAND4_X2 U1408 ( .A1(n14728), .A2(n14729), .A3(n14727), .A4(n14726), .ZN(
        n18134) );
  CLKBUF_X1 U1415 ( .A(n50339), .Z(n51025) );
  XNOR2_X1 U1430 ( .A(n43814), .B(n43813), .ZN(n50339) );
  BUF_X2 U1458 ( .A(n50637), .Z(n51029) );
  OAI211_X1 U1463 ( .C1(n47293), .C2(n47023), .A(n43903), .B(n43902), .ZN(
        n50637) );
  OR2_X2 U1482 ( .A1(n7163), .A2(n9792), .ZN(n14220) );
  BUF_X1 U1507 ( .A(n16337), .Z(n51031) );
  BUF_X1 U1509 ( .A(n16337), .Z(n51032) );
  XNOR2_X1 U1529 ( .A(n16105), .B(n18777), .ZN(n16337) );
  XNOR2_X2 U1530 ( .A(n16672), .B(n16671), .ZN(n19504) );
  INV_X1 U1546 ( .A(n15068), .ZN(n15307) );
  OR2_X2 U1566 ( .A1(n7228), .A2(n12615), .ZN(n15068) );
  BUF_X2 U1572 ( .A(n35849), .Z(n38313) );
  NAND2_X2 U1573 ( .A1(n4662), .A2(n19804), .ZN(n23101) );
  XNOR2_X2 U1594 ( .A(n43384), .B(n45120), .ZN(n46288) );
  OR2_X2 U1596 ( .A1(n3233), .A2(n6403), .ZN(n6916) );
  NAND3_X1 U1612 ( .A1(n4001), .A2(n21400), .A3(n318), .ZN(n51033) );
  NAND3_X1 U1615 ( .A1(n4001), .A2(n21400), .A3(n318), .ZN(n51034) );
  NAND3_X1 U1616 ( .A1(n4001), .A2(n21400), .A3(n318), .ZN(n23902) );
  INV_X1 U1619 ( .A(n23902), .ZN(n23926) );
  OR2_X1 U1629 ( .A1(n29782), .A2(n28772), .ZN(n29780) );
  XNOR2_X1 U1685 ( .A(n16940), .B(n16939), .ZN(n19868) );
  AND4_X2 U1686 ( .A1(n927), .A2(n923), .A3(n922), .A4(n921), .ZN(n32935) );
  NAND4_X1 U1711 ( .A1(n8000), .A2(n22925), .A3(n22924), .A4(n22923), .ZN(
        n27210) );
  AND3_X2 U1712 ( .A1(n6214), .A2(n8992), .A3(n6213), .ZN(n13820) );
  INV_X2 U1734 ( .A(n16142), .ZN(n17365) );
  AND3_X2 U1754 ( .A1(n4988), .A2(n7677), .A3(n4989), .ZN(n21885) );
  BUF_X1 U1772 ( .A(n19213), .Z(n51046) );
  XNOR2_X1 U1780 ( .A(n17901), .B(n15649), .ZN(n19213) );
  CLKBUF_X1 U1782 ( .A(n16126), .Z(n51048) );
  BUF_X1 U1793 ( .A(n16126), .Z(n51050) );
  XNOR2_X1 U1794 ( .A(n16124), .B(n2081), .ZN(n16126) );
  XNOR2_X2 U1800 ( .A(n4956), .B(n43914), .ZN(n44056) );
  AND2_X1 U1801 ( .A1(n19965), .A2(n20334), .ZN(n21494) );
  OR2_X2 U1808 ( .A1(n2923), .A2(n3319), .ZN(n37241) );
  NAND4_X1 U1839 ( .A1(n36111), .A2(n36109), .A3(n36110), .A4(n36108), .ZN(
        n41208) );
  NAND4_X2 U1856 ( .A1(n30115), .A2(n30114), .A3(n30113), .A4(n30112), .ZN(
        n36805) );
  NAND4_X1 U1870 ( .A1(n14328), .A2(n13053), .A3(n13051), .A4(n13052), .ZN(
        n18168) );
  NAND2_X2 U1872 ( .A1(n5419), .A2(n7374), .ZN(n32105) );
  BUF_X1 U1883 ( .A(n28040), .Z(n51057) );
  XNOR2_X1 U1884 ( .A(n23042), .B(n26378), .ZN(n28040) );
  XNOR2_X1 U1899 ( .A(n46157), .B(n46158), .ZN(n50374) );
  XNOR2_X1 U1920 ( .A(n5623), .B(Key[137]), .ZN(n11515) );
  NAND2_X1 U1955 ( .A1(n51244), .A2(n9038), .ZN(n51064) );
  CLKBUF_X1 U1980 ( .A(n13504), .Z(n51067) );
  NAND4_X1 U1983 ( .A1(n11238), .A2(n7516), .A3(n8295), .A4(n9329), .ZN(n13504) );
  XNOR2_X1 U1990 ( .A(n45457), .B(n45456), .ZN(n46519) );
  NAND4_X2 U2013 ( .A1(n12956), .A2(n4252), .A3(n12957), .A4(n12955), .ZN(
        n17212) );
  BUF_X2 U2020 ( .A(n25198), .Z(n30181) );
  NAND4_X1 U2042 ( .A1(n48243), .A2(n48241), .A3(n48242), .A4(n48240), .ZN(
        n48365) );
  XNOR2_X1 U2063 ( .A(n25007), .B(n25006), .ZN(n30273) );
  XNOR2_X1 U2076 ( .A(n2617), .B(n34083), .ZN(n36035) );
  NAND4_X2 U2092 ( .A1(n39936), .A2(n39935), .A3(n39934), .A4(n39933), .ZN(
        n42715) );
  AND2_X2 U2098 ( .A1(n27525), .A2(n30393), .ZN(n30688) );
  OR2_X2 U2099 ( .A1(n41945), .A2(n6544), .ZN(n43596) );
  XNOR2_X1 U2119 ( .A(n1887), .B(n1888), .ZN(n37721) );
  AND3_X2 U2125 ( .A1(n6198), .A2(n6200), .A3(n37472), .ZN(n41850) );
  NAND4_X1 U2129 ( .A1(n14392), .A2(n14391), .A3(n14390), .A4(n14389), .ZN(
        n51080) );
  NAND4_X1 U2133 ( .A1(n14392), .A2(n14391), .A3(n14390), .A4(n14389), .ZN(
        n51081) );
  NAND4_X2 U2178 ( .A1(n7069), .A2(n35030), .A3(n7071), .A4(n7068), .ZN(n41292) );
  XNOR2_X2 U2183 ( .A(n15977), .B(n15976), .ZN(n21613) );
  XNOR2_X2 U2196 ( .A(n16346), .B(n51703), .ZN(n16568) );
  XNOR2_X2 U2212 ( .A(n9453), .B(Key[122]), .ZN(n9830) );
  BUF_X2 U2216 ( .A(n47382), .Z(n50233) );
  XNOR2_X2 U2218 ( .A(n6974), .B(n35230), .ZN(n38259) );
  BUF_X2 U2222 ( .A(n31307), .Z(n51085) );
  NAND2_X1 U2225 ( .A1(n6110), .A2(n24568), .ZN(n31307) );
  XNOR2_X2 U2233 ( .A(n16414), .B(n16415), .ZN(n19535) );
  NAND4_X2 U2236 ( .A1(n31319), .A2(n31318), .A3(n31317), .A4(n31316), .ZN(
        n35115) );
  XNOR2_X2 U2256 ( .A(n8026), .B(n8028), .ZN(n1417) );
  NOR2_X2 U2257 ( .A1(n33173), .A2(n34945), .ZN(n36381) );
  XNOR2_X2 U2259 ( .A(n35280), .B(n6937), .ZN(n34945) );
  AND2_X1 U2268 ( .A1(n48382), .A2(n51728), .ZN(n48341) );
  INV_X1 U2273 ( .A(n8104), .ZN(n51087) );
  CLKBUF_X2 U2283 ( .A(n49695), .Z(n51095) );
  BUF_X1 U2284 ( .A(n45399), .Z(n51101) );
  BUF_X1 U2308 ( .A(n31883), .Z(n51479) );
  INV_X1 U2325 ( .A(n7064), .ZN(n32616) );
  NAND2_X2 U2328 ( .A1(n2677), .A2(n748), .ZN(n27669) );
  BUF_X1 U2331 ( .A(n29488), .Z(n51110) );
  INV_X1 U2350 ( .A(n3143), .ZN(n28897) );
  INV_X1 U2359 ( .A(n22509), .ZN(n22831) );
  AND2_X1 U2363 ( .A1(n51125), .A2(n23316), .ZN(n22954) );
  BUF_X1 U2382 ( .A(n21391), .Z(n358) );
  BUF_X1 U2386 ( .A(n17822), .Z(n51134) );
  INV_X1 U2394 ( .A(n10068), .ZN(n10617) );
  CLKBUF_X1 U2395 ( .A(Key[42]), .Z(n274) );
  INV_X2 U2396 ( .A(n49347), .ZN(n49367) );
  OR2_X1 U2401 ( .A1(n43486), .A2(n43485), .ZN(n51395) );
  OR2_X1 U2408 ( .A1(n45507), .A2(n45506), .ZN(n51328) );
  OR2_X1 U2410 ( .A1(n46237), .A2(n46238), .ZN(n51321) );
  AND2_X2 U2414 ( .A1(n7500), .A2(n7502), .ZN(n49923) );
  AND4_X1 U2416 ( .A1(n47330), .A2(n47332), .A3(n47329), .A4(n47331), .ZN(
        n51480) );
  NAND4_X1 U2421 ( .A1(n47330), .A2(n47332), .A3(n47329), .A4(n47331), .ZN(
        n50234) );
  INV_X1 U2425 ( .A(n49465), .ZN(n51091) );
  AND4_X1 U2427 ( .A1(n8761), .A2(n46809), .A3(n46807), .A4(n46808), .ZN(
        n51312) );
  AND3_X1 U2429 ( .A1(n46761), .A2(n1233), .A3(n46764), .ZN(n51346) );
  NOR2_X1 U2432 ( .A1(n42514), .A2(n42513), .ZN(n42515) );
  AND3_X1 U2436 ( .A1(n7309), .A2(n45912), .A3(n7310), .ZN(n7311) );
  INV_X1 U2448 ( .A(n48033), .ZN(n51092) );
  NOR2_X1 U2449 ( .A1(n2422), .A2(n4625), .ZN(n8761) );
  AOI21_X1 U2467 ( .B1(n2805), .B2(n2806), .A(n2804), .ZN(n8006) );
  INV_X1 U2468 ( .A(n43281), .ZN(n45962) );
  BUF_X1 U2470 ( .A(n46989), .Z(n51421) );
  BUF_X2 U2475 ( .A(n44786), .Z(n46255) );
  OR2_X1 U2477 ( .A1(n50343), .A2(n47026), .ZN(n47294) );
  BUF_X1 U2492 ( .A(n46708), .Z(n51396) );
  INV_X1 U2493 ( .A(n49629), .ZN(n51093) );
  BUF_X1 U2497 ( .A(n50293), .Z(n51313) );
  CLKBUF_X1 U2498 ( .A(n49720), .Z(n51295) );
  BUF_X1 U2506 ( .A(n46899), .Z(n51513) );
  INV_X1 U2515 ( .A(n49720), .ZN(n51094) );
  BUF_X2 U2535 ( .A(n43575), .Z(n43141) );
  BUF_X2 U2552 ( .A(n43059), .Z(n43196) );
  AND2_X1 U2563 ( .A1(n37363), .A2(n37362), .ZN(n51371) );
  AND3_X1 U2596 ( .A1(n41019), .A2(n41020), .A3(n41021), .ZN(n51283) );
  BUF_X2 U2597 ( .A(n46042), .Z(n51097) );
  NAND2_X1 U2614 ( .A1(n39559), .A2(n7122), .ZN(n7121) );
  NAND4_X1 U2634 ( .A1(n40077), .A2(n40076), .A3(n40079), .A4(n40078), .ZN(
        n51460) );
  AND3_X1 U2665 ( .A1(n38426), .A2(n38427), .A3(n38432), .ZN(n51569) );
  BUF_X2 U2667 ( .A(n46121), .Z(n51100) );
  AOI21_X1 U2675 ( .B1(n7367), .B2(n7638), .A(n4646), .ZN(n7366) );
  AND3_X1 U2696 ( .A1(n42086), .A2(n42092), .A3(n5824), .ZN(n7646) );
  OR2_X1 U2706 ( .A1(n6551), .A2(n6550), .ZN(n6548) );
  INV_X2 U2708 ( .A(n43669), .ZN(n41797) );
  AND2_X1 U2713 ( .A1(n38401), .A2(n40672), .ZN(n38404) );
  NAND4_X1 U2717 ( .A1(n36024), .A2(n36026), .A3(n36025), .A4(n36023), .ZN(
        n51325) );
  NAND3_X1 U2729 ( .A1(n36140), .A2(n36139), .A3(n36138), .ZN(n51430) );
  AND4_X1 U2741 ( .A1(n35411), .A2(n35414), .A3(n35413), .A4(n35412), .ZN(
        n51297) );
  AND4_X1 U2763 ( .A1(n7507), .A2(n7505), .A3(n7506), .A4(n36049), .ZN(n40110)
         );
  NAND4_X1 U2767 ( .A1(n7507), .A2(n7505), .A3(n7506), .A4(n36049), .ZN(n51352) );
  MUX2_X1 U2812 ( .A(n37487), .B(n37486), .S(n38522), .Z(n37494) );
  AND2_X1 U2814 ( .A1(n38009), .A2(n38176), .ZN(n51217) );
  AOI22_X1 U2816 ( .A1(n36136), .A2(n36135), .B1(n37576), .B2(n36134), .ZN(
        n36139) );
  OAI211_X1 U2827 ( .C1(n39403), .C2(n39402), .A(n5049), .B(n39405), .ZN(n5048) );
  AOI21_X1 U2829 ( .B1(n36046), .B2(n4279), .A(n2369), .ZN(n7507) );
  AND2_X1 U2832 ( .A1(n39389), .A2(n39368), .ZN(n51258) );
  AND2_X1 U2839 ( .A1(n37228), .A2(n6456), .ZN(n38632) );
  BUF_X1 U2878 ( .A(n37484), .Z(n51411) );
  BUF_X2 U3060 ( .A(n33173), .Z(n38043) );
  BUF_X1 U3061 ( .A(n34906), .Z(n39399) );
  INV_X1 U3090 ( .A(n38957), .ZN(n51102) );
  CLKBUF_X1 U3112 ( .A(n33983), .Z(n51495) );
  INV_X1 U3139 ( .A(n32717), .ZN(n32311) );
  OR2_X1 U3151 ( .A1(n31546), .A2(n31538), .ZN(n31549) );
  INV_X1 U3159 ( .A(n30982), .ZN(n708) );
  INV_X1 U3243 ( .A(n32507), .ZN(n51105) );
  NOR2_X1 U3267 ( .A1(n1641), .A2(n51557), .ZN(n1841) );
  NAND4_X1 U3273 ( .A1(n25848), .A2(n25853), .A3(n25849), .A4(n25850), .ZN(
        n31883) );
  NAND4_X1 U3280 ( .A1(n26662), .A2(n26663), .A3(n26664), .A4(n26665), .ZN(
        n26711) );
  NAND4_X1 U3286 ( .A1(n29197), .A2(n29196), .A3(n846), .A4(n29195), .ZN(
        n51520) );
  AND2_X1 U3303 ( .A1(n398), .A2(n29535), .ZN(n28615) );
  OR2_X1 U3323 ( .A1(n29462), .A2(n29459), .ZN(n29455) );
  BUF_X2 U3366 ( .A(n29347), .Z(n51109) );
  INV_X1 U3369 ( .A(n26158), .ZN(n51111) );
  INV_X1 U3373 ( .A(n29421), .ZN(n51112) );
  INV_X1 U3379 ( .A(n29933), .ZN(n51113) );
  BUF_X2 U3383 ( .A(n28659), .Z(n51114) );
  BUF_X2 U3387 ( .A(n28919), .Z(n51115) );
  INV_X1 U3406 ( .A(n29182), .ZN(n51116) );
  BUF_X2 U3410 ( .A(n27663), .Z(n51117) );
  XNOR2_X1 U3462 ( .A(n28228), .B(n28227), .ZN(n28348) );
  XNOR2_X1 U3474 ( .A(n25935), .B(n25934), .ZN(n27217) );
  BUF_X2 U3511 ( .A(n23772), .Z(n28214) );
  NAND4_X1 U3548 ( .A1(n51157), .A2(n22808), .A3(n22807), .A4(n22806), .ZN(
        n24976) );
  AOI21_X1 U3559 ( .B1(n7774), .B2(n23617), .A(n51548), .ZN(n7773) );
  INV_X1 U3575 ( .A(n24936), .ZN(n51122) );
  OAI211_X1 U3578 ( .C1(n23194), .C2(n23196), .A(n18861), .B(n18860), .ZN(
        n25903) );
  OR3_X2 U3615 ( .A1(n18386), .A2(n6576), .A3(n18372), .ZN(n1377) );
  NOR2_X1 U3641 ( .A1(n24023), .A2(n24024), .ZN(n2068) );
  OR2_X1 U3645 ( .A1(n23037), .A2(n22531), .ZN(n23993) );
  AND2_X1 U3650 ( .A1(n22944), .A2(n424), .ZN(n51603) );
  AND2_X1 U3687 ( .A1(n3778), .A2(n23702), .ZN(n23707) );
  INV_X1 U3704 ( .A(n21755), .ZN(n1024) );
  NAND2_X1 U3711 ( .A1(n3907), .A2(n23895), .ZN(n23923) );
  INV_X1 U3780 ( .A(n51580), .ZN(n2232) );
  INV_X1 U3812 ( .A(n23314), .ZN(n51125) );
  OR2_X1 U3814 ( .A1(n14383), .A2(n18327), .ZN(n51218) );
  AND2_X1 U3817 ( .A1(n20630), .A2(n21533), .ZN(n51551) );
  OR2_X1 U3842 ( .A1(n20473), .A2(n17639), .ZN(n19382) );
  OR2_X1 U3907 ( .A1(n21544), .A2(n20628), .ZN(n20741) );
  INV_X1 U3927 ( .A(n19048), .ZN(n51126) );
  INV_X1 U3944 ( .A(n20209), .ZN(n51128) );
  INV_X1 U3979 ( .A(n20745), .ZN(n51129) );
  INV_X1 U4017 ( .A(n20472), .ZN(n51130) );
  XNOR2_X1 U4131 ( .A(n51174), .B(n13572), .ZN(n17576) );
  BUF_X2 U4154 ( .A(n21251), .Z(n51132) );
  XNOR2_X1 U4162 ( .A(n51251), .B(n15938), .ZN(n15941) );
  XNOR2_X1 U4168 ( .A(n15940), .B(n16057), .ZN(n51251) );
  XNOR2_X1 U4186 ( .A(n15883), .B(n14698), .ZN(n15018) );
  BUF_X2 U4194 ( .A(n16926), .Z(n51482) );
  BUF_X2 U4215 ( .A(n18196), .Z(n51133) );
  AND2_X1 U4232 ( .A1(n14695), .A2(n14694), .ZN(n51237) );
  NOR2_X1 U4242 ( .A1(n15241), .A2(n13273), .ZN(n13286) );
  BUF_X2 U4292 ( .A(n18431), .Z(n51135) );
  INV_X1 U4298 ( .A(n7361), .ZN(n14826) );
  INV_X1 U4314 ( .A(n780), .ZN(n14247) );
  OR2_X1 U4338 ( .A1(n13711), .A2(n51579), .ZN(n13705) );
  AND2_X1 U4349 ( .A1(n7802), .A2(n14982), .ZN(n780) );
  INV_X1 U4366 ( .A(n5099), .ZN(n14516) );
  NOR2_X1 U4376 ( .A1(n14107), .A2(n14453), .ZN(n14441) );
  AND2_X1 U4377 ( .A1(n14863), .A2(n15448), .ZN(n51575) );
  INV_X1 U4412 ( .A(n13819), .ZN(n14321) );
  AND2_X1 U4422 ( .A1(n13306), .A2(n14022), .ZN(n13299) );
  INV_X1 U4485 ( .A(n15244), .ZN(n15204) );
  OR2_X1 U4487 ( .A1(n14472), .A2(n11737), .ZN(n9719) );
  AND2_X1 U4515 ( .A1(n13797), .A2(n13800), .ZN(n13480) );
  AND4_X1 U4539 ( .A1(n12468), .A2(n12469), .A3(n12466), .A4(n12467), .ZN(
        n51500) );
  AOI21_X1 U4568 ( .B1(n11461), .B2(n51150), .A(n51238), .ZN(n11238) );
  AND2_X1 U4569 ( .A1(n2236), .A2(n51612), .ZN(n51611) );
  AND4_X1 U4602 ( .A1(n11117), .A2(n11114), .A3(n11116), .A4(n11115), .ZN(
        n15244) );
  AOI21_X1 U4607 ( .B1(n51550), .B2(n10369), .A(n51549), .ZN(n10380) );
  OR2_X1 U4608 ( .A1(n10921), .A2(n10147), .ZN(n9735) );
  OR2_X1 U4614 ( .A1(n10182), .A2(n10555), .ZN(n51535) );
  AND2_X1 U4620 ( .A1(n11958), .A2(n12728), .ZN(n51171) );
  OR2_X1 U4646 ( .A1(n11346), .A2(n6267), .ZN(n9646) );
  AND2_X1 U4661 ( .A1(n12120), .A2(n10368), .ZN(n51549) );
  OR2_X1 U4671 ( .A1(n12111), .A2(n10367), .ZN(n10706) );
  OR2_X1 U4684 ( .A1(n9743), .A2(n8781), .ZN(n2703) );
  INV_X1 U4687 ( .A(n11695), .ZN(n51182) );
  NAND2_X2 U4709 ( .A1(n2680), .A2(n9667), .ZN(n10288) );
  INV_X1 U4713 ( .A(n9785), .ZN(n51137) );
  BUF_X1 U4732 ( .A(n11028), .Z(n580) );
  AND2_X1 U4736 ( .A1(n11581), .A2(n11515), .ZN(n11579) );
  BUF_X2 U4769 ( .A(n12084), .Z(n51138) );
  BUF_X2 U4782 ( .A(n12612), .Z(n51140) );
  OR2_X1 U4833 ( .A1(n10431), .A2(n11942), .ZN(n51577) );
  INV_X1 U4855 ( .A(n795), .ZN(n12604) );
  AND2_X1 U4862 ( .A1(n12640), .A2(n12638), .ZN(n51621) );
  AND2_X1 U4877 ( .A1(n11066), .A2(n12481), .ZN(n51554) );
  AND2_X1 U4915 ( .A1(n12635), .A2(n9208), .ZN(n12620) );
  XNOR2_X1 U4921 ( .A(n9255), .B(Key[7]), .ZN(n12610) );
  AND2_X1 U4948 ( .A1(n11920), .A2(n11914), .ZN(n12594) );
  INV_X1 U4967 ( .A(n12451), .ZN(n12672) );
  OR2_X1 U4988 ( .A1(n9433), .A2(n10398), .ZN(n8050) );
  INV_X1 U5026 ( .A(n12170), .ZN(n10417) );
  OR2_X1 U5041 ( .A1(n6911), .A2(n9573), .ZN(n51584) );
  OR2_X1 U5043 ( .A1(n10985), .A2(n10991), .ZN(n12367) );
  NAND2_X1 U5045 ( .A1(n2584), .A2(n2156), .ZN(n12711) );
  CLKBUF_X1 U5048 ( .A(n12555), .Z(n51491) );
  OR2_X1 U5052 ( .A1(n12577), .A2(n11568), .ZN(n2962) );
  AND2_X1 U5054 ( .A1(n9752), .A2(n10245), .ZN(n11003) );
  INV_X1 U5068 ( .A(n10195), .ZN(n9748) );
  AOI22_X1 U5069 ( .A1(n10452), .A2(n10453), .B1(n10454), .B2(n11976), .ZN(
        n10459) );
  AND3_X1 U5078 ( .A1(n12439), .A2(n12438), .A3(n3711), .ZN(n12448) );
  AND4_X1 U5122 ( .A1(n9457), .A2(n9458), .A3(n9964), .A4(n9456), .ZN(n9470)
         );
  OR2_X1 U5124 ( .A1(n9933), .A2(n11210), .ZN(n1078) );
  AND3_X1 U5142 ( .A1(n51167), .A2(n10202), .A3(n6841), .ZN(n3329) );
  AND3_X1 U5147 ( .A1(n9572), .A2(n9570), .A3(n9565), .ZN(n51219) );
  INV_X1 U5149 ( .A(n14720), .ZN(n14088) );
  AND3_X1 U5158 ( .A1(n9040), .A2(n9039), .A3(n9041), .ZN(n51244) );
  NOR2_X1 U5159 ( .A1(n11938), .A2(n11939), .ZN(n11940) );
  AOI22_X1 U5166 ( .A1(n7464), .A2(n13853), .B1(n13844), .B2(n2522), .ZN(
        n11735) );
  AND2_X1 U5190 ( .A1(n12101), .A2(n12100), .ZN(n51264) );
  AND2_X1 U5194 ( .A1(n8664), .A2(n11909), .ZN(n127) );
  AND4_X1 U5195 ( .A1(n9887), .A2(n9886), .A3(n9885), .A4(n9884), .ZN(n14837)
         );
  INV_X1 U5209 ( .A(n12755), .ZN(n14641) );
  OR2_X1 U5221 ( .A1(n9829), .A2(n10556), .ZN(n10537) );
  AOI21_X1 U5231 ( .B1(n15244), .B2(n14761), .A(n14760), .ZN(n14774) );
  NAND2_X2 U5235 ( .A1(n51244), .A2(n9038), .ZN(n13819) );
  INV_X1 U5251 ( .A(n15081), .ZN(n15302) );
  NAND4_X1 U5253 ( .A1(n13736), .A2(n1873), .A3(n13737), .A4(n11049), .ZN(
        n6724) );
  AND2_X1 U5255 ( .A1(n7688), .A2(n12205), .ZN(n13575) );
  NOR2_X1 U5339 ( .A1(n14411), .A2(n14393), .ZN(n12869) );
  AND2_X1 U5363 ( .A1(n14317), .A2(n14311), .ZN(n14322) );
  OR2_X1 U5364 ( .A1(n12981), .A2(n14533), .ZN(n12187) );
  BUF_X1 U5387 ( .A(n17913), .Z(n2214) );
  CLKBUF_X1 U5399 ( .A(n16535), .Z(n51402) );
  AND2_X1 U5421 ( .A1(n20460), .A2(n51130), .ZN(n51246) );
  OR2_X1 U5439 ( .A1(n20685), .A2(n1621), .ZN(n20674) );
  OR2_X1 U5498 ( .A1(n17576), .A2(n17484), .ZN(n17567) );
  XNOR2_X1 U5547 ( .A(n4635), .B(n15156), .ZN(n17873) );
  OR2_X1 U5548 ( .A1(n20016), .A2(n20015), .ZN(n51206) );
  NOR2_X1 U5562 ( .A1(n17859), .A2(n19330), .ZN(n19322) );
  AND2_X1 U5614 ( .A1(n5953), .A2(n51710), .ZN(n21566) );
  INV_X1 U5618 ( .A(n20157), .ZN(n5058) );
  INV_X1 U5667 ( .A(n19814), .ZN(n19734) );
  INV_X1 U5669 ( .A(n20118), .ZN(n20125) );
  AND2_X1 U5675 ( .A1(n20322), .A2(n19956), .ZN(n20321) );
  AND2_X1 U5684 ( .A1(n6875), .A2(n21948), .ZN(n51250) );
  OR2_X1 U5689 ( .A1(n21479), .A2(n4174), .ZN(n21500) );
  INV_X1 U5694 ( .A(n18937), .ZN(n18936) );
  BUF_X1 U5721 ( .A(n19839), .Z(n51434) );
  OR2_X1 U5730 ( .A1(n22129), .A2(n23257), .ZN(n20932) );
  INV_X1 U5731 ( .A(n18966), .ZN(n21242) );
  AND2_X1 U5768 ( .A1(n21946), .A2(n23467), .ZN(n51558) );
  AND2_X1 U5797 ( .A1(n5415), .A2(n23535), .ZN(n23379) );
  OR2_X1 U5803 ( .A1(n24211), .A2(n23068), .ZN(n22635) );
  OR2_X1 U5811 ( .A1(n20849), .A2(n23955), .ZN(n51623) );
  AND3_X1 U5812 ( .A1(n18066), .A2(n14379), .A3(n51218), .ZN(n14392) );
  AND2_X1 U5824 ( .A1(n22509), .A2(n22506), .ZN(n22490) );
  AND2_X1 U5830 ( .A1(n21589), .A2(n21590), .ZN(n94) );
  OR2_X1 U5840 ( .A1(n5370), .A2(n22375), .ZN(n22379) );
  OR2_X1 U5844 ( .A1(n22919), .A2(n22363), .ZN(n22909) );
  NOR2_X1 U5852 ( .A1(n23832), .A2(n630), .ZN(n1450) );
  OR2_X1 U5853 ( .A1(n22144), .A2(n22155), .ZN(n21919) );
  AND3_X1 U5865 ( .A1(n20848), .A2(n51623), .A3(n20847), .ZN(n4449) );
  INV_X1 U5910 ( .A(n22490), .ZN(n20297) );
  AND3_X1 U5917 ( .A1(n24005), .A2(n24006), .A3(n24004), .ZN(n250) );
  INV_X1 U5918 ( .A(n23316), .ZN(n756) );
  AND2_X1 U5923 ( .A1(n22188), .A2(n21714), .ZN(n22191) );
  INV_X1 U5936 ( .A(n21820), .ZN(n24250) );
  AND2_X1 U5937 ( .A1(n23616), .A2(n23615), .ZN(n51548) );
  NOR2_X1 U5955 ( .A1(n23833), .A2(n630), .ZN(n24161) );
  OR2_X1 U5959 ( .A1(n22701), .A2(n21782), .ZN(n22291) );
  NOR2_X1 U5986 ( .A1(n22182), .A2(n22181), .ZN(n22194) );
  AND4_X1 U5989 ( .A1(n851), .A2(n20524), .A3(n20525), .A4(n20526), .ZN(n20530) );
  OAI21_X1 U6031 ( .B1(n22721), .B2(n22722), .A(n22720), .ZN(n22723) );
  XNOR2_X1 U6074 ( .A(n28259), .B(n28258), .ZN(n28260) );
  NAND2_X1 U6075 ( .A1(n2004), .A2(n24455), .ZN(n25385) );
  XOR2_X1 U6084 ( .A(n24857), .B(n26273), .Z(n8723) );
  OR2_X1 U6088 ( .A1(n30709), .A2(n30705), .ZN(n1052) );
  OR2_X1 U6097 ( .A1(n30165), .A2(n30162), .ZN(n227) );
  XNOR2_X1 U6131 ( .A(n6659), .B(n25803), .ZN(n25479) );
  OR2_X1 U6133 ( .A1(n51514), .A2(n29159), .ZN(n29156) );
  OR2_X1 U6146 ( .A1(n28032), .A2(n29141), .ZN(n237) );
  OR2_X1 U6197 ( .A1(n25106), .A2(n5564), .ZN(n29115) );
  AND2_X1 U6199 ( .A1(n8681), .A2(n32917), .ZN(n51608) );
  OR2_X1 U6202 ( .A1(n31040), .A2(n26711), .ZN(n1682) );
  INV_X1 U6218 ( .A(n29734), .ZN(n30448) );
  OAI21_X1 U6219 ( .B1(n26324), .B2(n26325), .A(n29321), .ZN(n8209) );
  AND2_X1 U6234 ( .A1(n26781), .A2(n27765), .ZN(n29457) );
  OR2_X1 U6235 ( .A1(n24984), .A2(n29155), .ZN(n8082) );
  AND2_X1 U6262 ( .A1(n27782), .A2(n29283), .ZN(n29181) );
  NOR2_X1 U6275 ( .A1(n32136), .A2(n31699), .ZN(n51546) );
  INV_X1 U6281 ( .A(n31010), .ZN(n51223) );
  AND2_X1 U6313 ( .A1(n1428), .A2(n32402), .ZN(n51177) );
  AND2_X1 U6326 ( .A1(n24573), .A2(n24575), .ZN(n281) );
  AND2_X1 U6335 ( .A1(n27909), .A2(n27971), .ZN(n27911) );
  INV_X1 U6340 ( .A(n31747), .ZN(n51532) );
  AND3_X1 U6352 ( .A1(n29500), .A2(n51568), .A3(n51567), .ZN(n6362) );
  CLKBUF_X1 U6353 ( .A(n24092), .Z(n30687) );
  OR2_X1 U6355 ( .A1(n33013), .A2(n33005), .ZN(n30539) );
  AND2_X1 U6377 ( .A1(n33009), .A2(n51223), .ZN(n26638) );
  INV_X1 U6394 ( .A(n32214), .ZN(n716) );
  NOR2_X1 U6399 ( .A1(n32356), .A2(n1385), .ZN(n32051) );
  OR2_X1 U6435 ( .A1(n27528), .A2(n51257), .ZN(n27530) );
  OAI21_X1 U6458 ( .B1(n26484), .B2(n26485), .A(n29174), .ZN(n26492) );
  OR2_X1 U6485 ( .A1(n30982), .A2(n31684), .ZN(n31676) );
  AND2_X1 U6498 ( .A1(n32687), .A2(n31670), .ZN(n51564) );
  XNOR2_X1 U6528 ( .A(n36703), .B(n36700), .ZN(n242) );
  OAI21_X1 U6543 ( .B1(n32816), .B2(n51617), .A(n51616), .ZN(n30477) );
  AND3_X1 U6610 ( .A1(n32413), .A2(n32414), .A3(n32405), .ZN(n51220) );
  AOI22_X1 U6651 ( .A1(n31451), .A2(n31455), .B1(n31449), .B2(n31450), .ZN(
        n51533) );
  AND2_X1 U6675 ( .A1(n7477), .A2(n29997), .ZN(n258) );
  XNOR2_X1 U6705 ( .A(n5616), .B(n34361), .ZN(n51366) );
  XNOR2_X1 U6711 ( .A(n36722), .B(n32859), .ZN(n35618) );
  XNOR2_X1 U6725 ( .A(n5234), .B(n36829), .ZN(n35286) );
  XNOR2_X1 U6734 ( .A(n35543), .B(n32310), .ZN(n51449) );
  CLKBUF_X1 U6740 ( .A(n34122), .Z(n51501) );
  AND2_X1 U6741 ( .A1(n31084), .A2(n32373), .ZN(n51537) );
  XNOR2_X1 U6751 ( .A(n34566), .B(n34565), .ZN(n51573) );
  OR2_X1 U6761 ( .A1(n39300), .A2(n39307), .ZN(n51273) );
  XNOR2_X1 U6786 ( .A(n33240), .B(n8321), .ZN(n35402) );
  AND3_X1 U6797 ( .A1(n51282), .A2(n35986), .A3(n51281), .ZN(n7348) );
  XNOR2_X1 U6869 ( .A(n37111), .B(n35231), .ZN(n36730) );
  INV_X1 U6877 ( .A(n36000), .ZN(n37640) );
  AND2_X1 U6898 ( .A1(n35443), .A2(n35444), .ZN(n35) );
  OR2_X1 U6905 ( .A1(n38590), .A2(n38593), .ZN(n38596) );
  INV_X1 U6928 ( .A(n39478), .ZN(n36215) );
  AND2_X1 U6967 ( .A1(n38728), .A2(n38722), .ZN(n39288) );
  OAI21_X1 U6994 ( .B1(n39938), .B2(n39754), .A(n39955), .ZN(n39764) );
  CLKBUF_X1 U7010 ( .A(n34908), .Z(n37731) );
  AND2_X1 U7013 ( .A1(n39346), .A2(n35946), .ZN(n104) );
  OR2_X1 U7049 ( .A1(n41212), .A2(n51052), .ZN(n39499) );
  AND3_X1 U7063 ( .A1(n7377), .A2(n34678), .A3(n34680), .ZN(n51190) );
  AND3_X1 U7065 ( .A1(n35143), .A2(n35144), .A3(n35145), .ZN(n254) );
  NOR2_X1 U7074 ( .A1(n35), .A2(n51241), .ZN(n35449) );
  AND3_X1 U7091 ( .A1(n35569), .A2(n51632), .A3(n38538), .ZN(n7847) );
  INV_X1 U7144 ( .A(n40388), .ZN(n135) );
  INV_X1 U7158 ( .A(n51620), .ZN(n51619) );
  OR2_X1 U7183 ( .A1(n39908), .A2(n39912), .ZN(n38449) );
  INV_X1 U7191 ( .A(n675), .ZN(n2065) );
  INV_X1 U7220 ( .A(n40910), .ZN(n40901) );
  BUF_X1 U7237 ( .A(n40272), .Z(n2224) );
  INV_X1 U7435 ( .A(n674), .ZN(n41327) );
  AND2_X1 U7465 ( .A1(n40817), .A2(n40818), .ZN(n675) );
  AND3_X1 U7471 ( .A1(n36390), .A2(n7208), .A3(n36391), .ZN(n36394) );
  AND2_X1 U7474 ( .A1(n2063), .A2(n675), .ZN(n40138) );
  AND3_X1 U7479 ( .A1(n845), .A2(n38873), .A3(n38874), .ZN(n38883) );
  AND4_X1 U7516 ( .A1(n35886), .A2(n35885), .A3(n35884), .A4(n35883), .ZN(
        n38445) );
  AND2_X1 U7527 ( .A1(n52198), .A2(n3861), .ZN(n41231) );
  OAI21_X1 U7535 ( .B1(n38780), .B2(n40124), .A(n40126), .ZN(n7240) );
  NOR2_X1 U7537 ( .A1(n41038), .A2(n41037), .ZN(n41043) );
  XNOR2_X1 U7542 ( .A(n41629), .B(n6573), .ZN(n42869) );
  XNOR2_X1 U7551 ( .A(n42962), .B(n45459), .ZN(n44098) );
  XNOR2_X1 U7558 ( .A(n42626), .B(n43522), .ZN(n44553) );
  OR2_X1 U7567 ( .A1(n49218), .A2(n49216), .ZN(n132) );
  NAND2_X1 U7601 ( .A1(n46276), .A2(n45237), .ZN(n46342) );
  AND2_X1 U7605 ( .A1(n44708), .A2(n44840), .ZN(n7127) );
  AND2_X1 U7607 ( .A1(n41923), .A2(n918), .ZN(n917) );
  OR2_X1 U7624 ( .A1(n45868), .A2(n45869), .ZN(n45871) );
  NOR2_X1 U7632 ( .A1(n47831), .A2(n51470), .ZN(n47855) );
  NAND4_X1 U7741 ( .A1(n44284), .A2(n44285), .A3(n3054), .A4(n3051), .ZN(
        n51343) );
  OR2_X1 U7775 ( .A1(n47199), .A2(n51315), .ZN(n51274) );
  AND2_X1 U7793 ( .A1(n46180), .A2(n46181), .ZN(n51276) );
  AND2_X1 U7807 ( .A1(n5444), .A2(n14257), .ZN(n51142) );
  INV_X1 U7855 ( .A(n13930), .ZN(n13206) );
  OR2_X1 U7909 ( .A1(n14133), .A2(n14573), .ZN(n51143) );
  NOR3_X1 U7932 ( .A1(n14296), .A2(n14295), .A3(n14294), .ZN(n51144) );
  AND3_X1 U8037 ( .A1(n5415), .A2(n457), .A3(n23531), .ZN(n51145) );
  AND4_X1 U8051 ( .A1(n37495), .A2(n37494), .A3(n37493), .A4(n37492), .ZN(
        n51146) );
  NOR2_X1 U8077 ( .A1(n40149), .A2(n52160), .ZN(n51147) );
  AND2_X1 U8098 ( .A1(n20487), .A2(n21465), .ZN(n51148) );
  AND3_X1 U8144 ( .A1(n14298), .A2(n5411), .A3(n14297), .ZN(n51149) );
  AND2_X1 U8156 ( .A1(n11470), .A2(n11466), .ZN(n51150) );
  NAND2_X1 U8216 ( .A1(n18863), .A2(n15872), .ZN(n20685) );
  NAND4_X1 U8229 ( .A1(n35411), .A2(n35414), .A3(n35413), .A4(n35412), .ZN(
        n39667) );
  INV_X1 U8233 ( .A(n29325), .ZN(n29319) );
  INV_X1 U8249 ( .A(n10673), .ZN(n51194) );
  INV_X1 U8318 ( .A(n11379), .ZN(n51256) );
  OR2_X1 U8321 ( .A1(n10068), .A2(n10065), .ZN(n51151) );
  AND2_X1 U8335 ( .A1(n13352), .A2(n14542), .ZN(n51152) );
  NOR2_X1 U8365 ( .A1(n9178), .A2(n9186), .ZN(n10451) );
  NAND4_X1 U8385 ( .A1(n10679), .A2(n10681), .A3(n10680), .A4(n10682), .ZN(
        n13323) );
  INV_X1 U8508 ( .A(n13323), .ZN(n51534) );
  INV_X1 U8531 ( .A(n9), .ZN(n14095) );
  INV_X1 U8552 ( .A(n20013), .ZN(n51208) );
  AND2_X1 U8561 ( .A1(n8401), .A2(n8159), .ZN(n51153) );
  INV_X1 U8587 ( .A(n19086), .ZN(n51222) );
  OR2_X1 U8599 ( .A1(n22799), .A2(n5143), .ZN(n51154) );
  INV_X1 U8644 ( .A(n23336), .ZN(n51200) );
  NAND3_X1 U8709 ( .A1(n18961), .A2(n17078), .A3(n17077), .ZN(n51155) );
  AND3_X1 U8720 ( .A1(n25056), .A2(n23101), .A3(n22875), .ZN(n51156) );
  AND3_X1 U8745 ( .A1(n51191), .A2(n22798), .A3(n51154), .ZN(n51157) );
  NAND2_X1 U8773 ( .A1(n21145), .A2(n20868), .ZN(n51158) );
  AND2_X1 U8819 ( .A1(n27854), .A2(n2956), .ZN(n51159) );
  INV_X1 U8930 ( .A(n32815), .ZN(n8542) );
  INV_X1 U8960 ( .A(n8542), .ZN(n51618) );
  AND4_X1 U8975 ( .A1(n30397), .A2(n4216), .A3(n4217), .A4(n30396), .ZN(n51160) );
  AND2_X1 U9028 ( .A1(n38949), .A2(n38651), .ZN(n51161) );
  AND2_X1 U9168 ( .A1(n39299), .A2(n2436), .ZN(n51162) );
  AND2_X1 U9208 ( .A1(n34706), .A2(n36208), .ZN(n51163) );
  AND2_X1 U9297 ( .A1(n51234), .A2(n51232), .ZN(n51164) );
  NOR2_X1 U9340 ( .A1(n50497), .A2(n50536), .ZN(n51165) );
  AND3_X1 U9352 ( .A1(n47543), .A2(n51287), .A3(n47575), .ZN(n51166) );
  NOR2_X1 U9379 ( .A1(n32063), .A2(n32062), .ZN(n51179) );
  NAND3_X1 U9391 ( .A1(n7627), .A2(n31556), .A3(n31557), .ZN(n6394) );
  OAI21_X1 U9419 ( .B1(n10200), .B2(n10241), .A(n11006), .ZN(n51167) );
  AND2_X2 U9440 ( .A1(n51168), .A2(n8691), .ZN(n30058) );
  NAND3_X1 U9541 ( .A1(n19352), .A2(n21466), .A3(n19357), .ZN(n17743) );
  NAND2_X1 U9542 ( .A1(n11005), .A2(n11011), .ZN(n8782) );
  NAND2_X1 U9562 ( .A1(n8776), .A2(n10240), .ZN(n11005) );
  NAND4_X1 U9601 ( .A1(n15002), .A2(n5346), .A3(n14996), .A4(n15001), .ZN(
        n5344) );
  XNOR2_X1 U9639 ( .A(n51169), .B(n45866), .ZN(Plaintext[15]) );
  NAND3_X1 U9676 ( .A1(n45863), .A2(n45865), .A3(n45864), .ZN(n51169) );
  NAND2_X1 U9677 ( .A1(n27408), .A2(n29905), .ZN(n1374) );
  NAND2_X1 U9699 ( .A1(n1375), .A2(n30790), .ZN(n27408) );
  NAND2_X1 U9724 ( .A1(n51793), .A2(n29325), .ZN(n26323) );
  XNOR2_X2 U9754 ( .A(n7834), .B(n7833), .ZN(n29325) );
  OAI21_X1 U9771 ( .B1(n14967), .B2(n14966), .A(n51170), .ZN(n14971) );
  INV_X1 U9793 ( .A(n14968), .ZN(n51170) );
  NAND2_X1 U9794 ( .A1(n11105), .A2(n51171), .ZN(n11106) );
  AOI22_X2 U9908 ( .A1(n8862), .A2(n51172), .B1(n14291), .B2(n13587), .ZN(
        n13984) );
  NAND2_X1 U9963 ( .A1(n8860), .A2(n5411), .ZN(n51172) );
  NAND2_X1 U9974 ( .A1(n5408), .A2(n10251), .ZN(n9030) );
  OAI211_X1 U10046 ( .C1(n23271), .C2(n23270), .A(n23269), .B(n51173), .ZN(
        n23272) );
  NAND2_X1 U10093 ( .A1(n24160), .A2(n23267), .ZN(n51173) );
  NAND2_X1 U10134 ( .A1(n3344), .A2(n21654), .ZN(n3343) );
  NAND2_X1 U10179 ( .A1(n15233), .A2(n15244), .ZN(n15196) );
  XNOR2_X1 U10202 ( .A(n5136), .B(n13536), .ZN(n51174) );
  INV_X1 U10239 ( .A(n17478), .ZN(n17580) );
  NAND2_X1 U10252 ( .A1(n29028), .A2(n28530), .ZN(n28160) );
  NAND2_X1 U10256 ( .A1(n20422), .A2(n17838), .ZN(n20423) );
  NAND2_X1 U10300 ( .A1(n22191), .A2(n21710), .ZN(n2554) );
  AND2_X1 U10362 ( .A1(n14155), .A2(n51175), .ZN(n818) );
  OR2_X2 U10403 ( .A1(n5926), .A2(n5929), .ZN(n14155) );
  NAND2_X1 U10428 ( .A1(n20296), .A2(n22490), .ZN(n22496) );
  INV_X1 U10481 ( .A(n51176), .ZN(n11506) );
  OAI211_X1 U10492 ( .C1(n11494), .C2(n11888), .A(n11492), .B(n11493), .ZN(
        n51176) );
  NAND3_X1 U10507 ( .A1(n29173), .A2(n30251), .A3(n29157), .ZN(n29162) );
  NAND2_X1 U10510 ( .A1(n32082), .A2(n51177), .ZN(n32083) );
  NAND2_X1 U10636 ( .A1(n1425), .A2(n51179), .ZN(n8711) );
  INV_X1 U10712 ( .A(n51180), .ZN(n20635) );
  OAI21_X1 U10713 ( .B1(n20632), .B2(n21538), .A(n20631), .ZN(n51180) );
  NAND3_X1 U10783 ( .A1(n22855), .A2(n22854), .A3(n23021), .ZN(n22871) );
  AOI21_X1 U10819 ( .B1(n13660), .B2(n13659), .A(n51181), .ZN(n13671) );
  NAND2_X1 U10906 ( .A1(n13658), .A2(n14644), .ZN(n51181) );
  NAND2_X1 U10932 ( .A1(n4411), .A2(n32009), .ZN(n31196) );
  NAND2_X1 U10988 ( .A1(n22253), .A2(n22252), .ZN(n7028) );
  AOI21_X1 U11024 ( .B1(n51183), .B2(n51182), .A(n11697), .ZN(n11703) );
  NAND2_X1 U11089 ( .A1(n11696), .A2(n11705), .ZN(n51183) );
  AND2_X1 U11145 ( .A1(n19298), .A2(n19299), .ZN(n51186) );
  NAND2_X1 U11207 ( .A1(n31995), .A2(n32507), .ZN(n31194) );
  XNOR2_X1 U11224 ( .A(n51185), .B(n23123), .ZN(n23190) );
  XNOR2_X1 U11260 ( .A(n23121), .B(n23120), .ZN(n51185) );
  NOR2_X1 U11277 ( .A1(n9081), .A2(n9082), .ZN(n9093) );
  NAND2_X1 U11313 ( .A1(n19662), .A2(n19891), .ZN(n18937) );
  NAND2_X2 U11314 ( .A1(n19300), .A2(n51186), .ZN(n23982) );
  NAND2_X1 U11318 ( .A1(n12066), .A2(n9203), .ZN(n12618) );
  NAND4_X2 U11360 ( .A1(n10022), .A2(n10024), .A3(n10025), .A4(n10023), .ZN(
        n13173) );
  NAND2_X1 U11457 ( .A1(n3381), .A2(n19695), .ZN(n19696) );
  INV_X1 U11476 ( .A(n39376), .ZN(n39387) );
  OAI21_X1 U11543 ( .B1(n39389), .B2(n39388), .A(n51187), .ZN(n3985) );
  NAND2_X1 U11608 ( .A1(n39376), .A2(n39194), .ZN(n51187) );
  AND2_X2 U11710 ( .A1(n7026), .A2(n39377), .ZN(n39376) );
  NAND2_X1 U11771 ( .A1(n11461), .A2(n11460), .ZN(n11463) );
  AND2_X2 U11799 ( .A1(n11229), .A2(n11468), .ZN(n11461) );
  NAND3_X1 U11818 ( .A1(n30745), .A2(n3967), .A3(n30744), .ZN(n30750) );
  NAND3_X1 U11821 ( .A1(n38264), .A2(n38252), .A3(n38262), .ZN(n38644) );
  NAND2_X1 U11847 ( .A1(n51189), .A2(n3042), .ZN(n22215) );
  NOR2_X1 U11915 ( .A1(n23100), .A2(n22763), .ZN(n51189) );
  NAND2_X1 U11998 ( .A1(n49836), .A2(n49841), .ZN(n49775) );
  INV_X1 U12006 ( .A(n10288), .ZN(n10286) );
  NAND2_X1 U12023 ( .A1(n19307), .A2(n51148), .ZN(n19313) );
  NAND3_X1 U12036 ( .A1(n23914), .A2(n23895), .A3(n8149), .ZN(n51191) );
  INV_X1 U12054 ( .A(n26994), .ZN(n26996) );
  NAND2_X1 U12101 ( .A1(n29424), .A2(n29422), .ZN(n26994) );
  NAND2_X1 U12114 ( .A1(n51193), .A2(n51192), .ZN(n2553) );
  NAND2_X1 U12134 ( .A1(n10673), .A2(n12328), .ZN(n51192) );
  NAND2_X1 U12143 ( .A1(n10288), .A2(n51194), .ZN(n51193) );
  NAND2_X1 U12144 ( .A1(n22690), .A2(n22522), .ZN(n22528) );
  NAND2_X1 U12193 ( .A1(n1148), .A2(n22520), .ZN(n22690) );
  INV_X1 U12233 ( .A(n31166), .ZN(n32664) );
  NAND2_X1 U12312 ( .A1(n31454), .A2(n31545), .ZN(n31166) );
  NAND3_X1 U12396 ( .A1(n51197), .A2(n20301), .A3(n20303), .ZN(n51196) );
  NOR2_X1 U12408 ( .A1(n51198), .A2(n20294), .ZN(n51197) );
  INV_X1 U12411 ( .A(n20300), .ZN(n51198) );
  AOI22_X1 U12414 ( .A1(n21459), .A2(n21460), .B1(n21462), .B2(n21461), .ZN(
        n21477) );
  NAND2_X1 U12429 ( .A1(n38721), .A2(n51162), .ZN(n37179) );
  NAND2_X1 U12449 ( .A1(n6748), .A2(n39300), .ZN(n38721) );
  NAND2_X1 U12468 ( .A1(n51233), .A2(n38380), .ZN(n6186) );
  NAND2_X1 U12558 ( .A1(n51200), .A2(n21755), .ZN(n23333) );
  NAND2_X2 U12570 ( .A1(n51199), .A2(n51153), .ZN(n21755) );
  NAND3_X1 U12611 ( .A1(n13214), .A2(n5830), .A3(n14229), .ZN(n9801) );
  NAND2_X1 U12622 ( .A1(n37647), .A2(n35732), .ZN(n6262) );
  NAND2_X1 U12637 ( .A1(n3093), .A2(n39551), .ZN(n3092) );
  OR2_X2 U12660 ( .A1(n30346), .A2(n28298), .ZN(n28300) );
  NAND2_X1 U12665 ( .A1(n7650), .A2(n7651), .ZN(n7649) );
  NAND3_X1 U12700 ( .A1(n45245), .A2(n46346), .A3(n46267), .ZN(n44760) );
  NAND2_X1 U12721 ( .A1(n42605), .A2(n46356), .ZN(n45686) );
  NAND3_X2 U12728 ( .A1(n28818), .A2(n28816), .A3(n28817), .ZN(n32634) );
  XNOR2_X1 U12733 ( .A(n51201), .B(n42533), .ZN(n42547) );
  XNOR2_X1 U12759 ( .A(n43742), .B(n42762), .ZN(n51201) );
  NAND2_X1 U12821 ( .A1(n40118), .A2(n40110), .ZN(n38781) );
  OAI211_X1 U12843 ( .C1(n35873), .C2(n36056), .A(n35206), .B(n51202), .ZN(
        n35207) );
  NAND2_X1 U12867 ( .A1(n22037), .A2(n3506), .ZN(n23420) );
  NAND2_X1 U12882 ( .A1(n590), .A2(n18288), .ZN(n20012) );
  XNOR2_X1 U12884 ( .A(n51203), .B(n14858), .ZN(n3508) );
  XNOR2_X1 U12888 ( .A(n2298), .B(n17912), .ZN(n51203) );
  NAND3_X2 U12898 ( .A1(n24253), .A2(n51204), .A3(n51205), .ZN(n26544) );
  NAND2_X1 U12910 ( .A1(n24243), .A2(n24242), .ZN(n51204) );
  NAND2_X1 U12917 ( .A1(n24241), .A2(n24250), .ZN(n51205) );
  OAI211_X1 U12974 ( .C1(n20018), .C2(n20019), .A(n51207), .B(n51206), .ZN(
        n2649) );
  INV_X1 U13022 ( .A(n20014), .ZN(n51209) );
  NAND4_X1 U13023 ( .A1(n51210), .A2(n5837), .A3(n50627), .A4(n50626), .ZN(
        n50629) );
  NAND2_X1 U13036 ( .A1(n50644), .A2(n5835), .ZN(n51210) );
  NAND3_X1 U13084 ( .A1(n39381), .A2(n39386), .A3(n39380), .ZN(n51211) );
  NAND2_X1 U13118 ( .A1(n18071), .A2(n403), .ZN(n18339) );
  NAND3_X1 U13121 ( .A1(n51213), .A2(n10620), .A3(n51212), .ZN(n10622) );
  INV_X1 U13138 ( .A(n10617), .ZN(n51212) );
  NAND2_X1 U13143 ( .A1(n10618), .A2(n10619), .ZN(n51213) );
  NAND2_X1 U13154 ( .A1(n10995), .A2(n51214), .ZN(n7810) );
  OAI21_X1 U13164 ( .B1(n3001), .B2(n10989), .A(n10988), .ZN(n51214) );
  AND3_X2 U13184 ( .A1(n5848), .A2(n5847), .A3(n43690), .ZN(n50638) );
  NOR2_X1 U13205 ( .A1(n32457), .A2(n32311), .ZN(n32314) );
  NAND3_X2 U13206 ( .A1(n40813), .A2(n40811), .A3(n40812), .ZN(n8515) );
  XNOR2_X1 U13213 ( .A(n51215), .B(n45708), .ZN(Plaintext[79]) );
  NAND3_X1 U13363 ( .A1(n5076), .A2(n40098), .A3(n40081), .ZN(n5075) );
  XNOR2_X1 U13366 ( .A(n51216), .B(n42600), .ZN(n42606) );
  XNOR2_X1 U13368 ( .A(n42599), .B(n42598), .ZN(n51216) );
  NAND3_X1 U13377 ( .A1(n38011), .A2(n38010), .A3(n51217), .ZN(n38026) );
  NAND2_X1 U13394 ( .A1(n6184), .A2(n34993), .ZN(n1036) );
  NAND3_X1 U13400 ( .A1(n22904), .A2(n22908), .A3(n22918), .ZN(n22905) );
  NAND4_X4 U13430 ( .A1(n12449), .A2(n12446), .A3(n12447), .A4(n12448), .ZN(
        n14962) );
  NAND3_X1 U13438 ( .A1(n11057), .A2(n311), .A3(n816), .ZN(n4074) );
  NAND3_X2 U13450 ( .A1(n51220), .A2(n8252), .A3(n8250), .ZN(n34811) );
  INV_X1 U13466 ( .A(n18961), .ZN(n19101) );
  NAND2_X1 U13490 ( .A1(n21250), .A2(n21253), .ZN(n18961) );
  NAND2_X1 U13521 ( .A1(n31011), .A2(n8517), .ZN(n33009) );
  NAND2_X1 U13574 ( .A1(n14454), .A2(n14106), .ZN(n9) );
  NOR2_X1 U13575 ( .A1(n12811), .A2(n12805), .ZN(n12806) );
  NAND3_X1 U13591 ( .A1(n16044), .A2(n51019), .A3(n13384), .ZN(n12811) );
  XNOR2_X2 U13596 ( .A(n17763), .B(n19196), .ZN(n5670) );
  NAND4_X2 U13611 ( .A1(n14425), .A2(n14423), .A3(n14426), .A4(n14424), .ZN(
        n19196) );
  NAND2_X1 U13618 ( .A1(n8032), .A2(n39853), .ZN(n8031) );
  NAND2_X1 U13622 ( .A1(n6591), .A2(n6592), .ZN(n6590) );
  NAND2_X1 U13646 ( .A1(n12757), .A2(n13659), .ZN(n12758) );
  NAND3_X1 U13685 ( .A1(n38167), .A2(n38166), .A3(n38156), .ZN(n35688) );
  XNOR2_X1 U13715 ( .A(n51224), .B(n41407), .ZN(n41409) );
  XNOR2_X1 U13731 ( .A(n41371), .B(n41370), .ZN(n51224) );
  NAND2_X2 U13751 ( .A1(n51225), .A2(n4821), .ZN(n14030) );
  NOR2_X1 U13765 ( .A1(n7810), .A2(n51784), .ZN(n51225) );
  NAND2_X1 U13828 ( .A1(n48041), .A2(n48077), .ZN(n48068) );
  NAND2_X1 U13838 ( .A1(n32988), .A2(n32974), .ZN(n28608) );
  NAND2_X1 U13851 ( .A1(n46575), .A2(n46699), .ZN(n45788) );
  NAND2_X1 U13867 ( .A1(n10246), .A2(n8781), .ZN(n8784) );
  XNOR2_X1 U13868 ( .A(n51226), .B(n49063), .ZN(Plaintext[96]) );
  NAND3_X1 U13905 ( .A1(n49061), .A2(n49062), .A3(n49060), .ZN(n51226) );
  NAND2_X1 U13927 ( .A1(n39110), .A2(n39937), .ZN(n51227) );
  AND2_X1 U14018 ( .A1(n6272), .A2(n39113), .ZN(n51228) );
  NAND3_X1 U14029 ( .A1(n39653), .A2(n37465), .A3(n37464), .ZN(n37466) );
  NAND2_X1 U14036 ( .A1(n28995), .A2(n29749), .ZN(n4102) );
  AND2_X1 U14073 ( .A1(n47655), .A2(n47686), .ZN(n47699) );
  XOR2_X1 U14127 ( .A(n34022), .B(n34021), .Z(n51578) );
  NAND3_X1 U14151 ( .A1(n19831), .A2(n19829), .A3(n19830), .ZN(n19833) );
  NOR2_X2 U14201 ( .A1(n13566), .A2(n13567), .ZN(n17879) );
  OR2_X1 U14212 ( .A1(n9650), .A2(n9649), .ZN(n51572) );
  NAND3_X1 U14262 ( .A1(n46329), .A2(n46327), .A3(n46328), .ZN(n51229) );
  NAND2_X1 U14273 ( .A1(n28144), .A2(n28563), .ZN(n27118) );
  NAND2_X1 U14277 ( .A1(n28145), .A2(n26494), .ZN(n24882) );
  NAND3_X1 U14283 ( .A1(n162), .A2(n3605), .A3(n21299), .ZN(n22544) );
  NOR2_X1 U14295 ( .A1(n26976), .A2(n5183), .ZN(n5182) );
  NAND2_X1 U14330 ( .A1(n27795), .A2(n28626), .ZN(n26976) );
  INV_X1 U14346 ( .A(n19254), .ZN(n18430) );
  XNOR2_X1 U14392 ( .A(n17644), .B(n15186), .ZN(n19254) );
  NAND2_X1 U14394 ( .A1(n32208), .A2(n32193), .ZN(n4489) );
  XNOR2_X1 U14404 ( .A(n51230), .B(n23286), .ZN(n23108) );
  XNOR2_X1 U14418 ( .A(n23018), .B(n23017), .ZN(n51230) );
  NAND2_X1 U14455 ( .A1(n1390), .A2(n1391), .ZN(n1389) );
  INV_X1 U14463 ( .A(n39764), .ZN(n8072) );
  NAND2_X1 U14480 ( .A1(n3564), .A2(n14139), .ZN(n4007) );
  XNOR2_X1 U14528 ( .A(n51231), .B(n43196), .ZN(n42625) );
  XNOR2_X1 U14540 ( .A(n42623), .B(n42622), .ZN(n51231) );
  NAND2_X1 U14577 ( .A1(n38770), .A2(n51233), .ZN(n51232) );
  INV_X1 U14578 ( .A(n2153), .ZN(n51233) );
  NAND2_X1 U14610 ( .A1(n39552), .A2(n2153), .ZN(n51234) );
  NOR2_X1 U14611 ( .A1(n38784), .A2(n51325), .ZN(n39552) );
  NAND2_X1 U14623 ( .A1(n3612), .A2(n30848), .ZN(n999) );
  NAND2_X2 U14659 ( .A1(n1646), .A2(n7869), .ZN(n41212) );
  AOI22_X1 U14660 ( .A1(n21377), .A2(n21376), .B1(n21378), .B2(n7836), .ZN(
        n21380) );
  NAND2_X1 U14667 ( .A1(n1861), .A2(n776), .ZN(n21377) );
  NAND2_X1 U14682 ( .A1(n3198), .A2(n48958), .ZN(n46950) );
  NOR2_X1 U14700 ( .A1(n3209), .A2(n48957), .ZN(n3198) );
  OAI211_X1 U14714 ( .C1(n413), .C2(n23209), .A(n51235), .B(n51355), .ZN(
        n20306) );
  OR2_X1 U14717 ( .A1(n23223), .A2(n23207), .ZN(n51235) );
  NAND2_X1 U14735 ( .A1(n7572), .A2(n14911), .ZN(n15081) );
  INV_X1 U14736 ( .A(n51236), .ZN(n5402) );
  OAI21_X1 U14773 ( .B1(n38415), .B2(n39929), .A(n40679), .ZN(n51236) );
  NAND4_X2 U14774 ( .A1(n11301), .A2(n11300), .A3(n11299), .A4(n11302), .ZN(
        n15883) );
  NOR2_X1 U14781 ( .A1(n10852), .A2(n11630), .ZN(n51238) );
  INV_X1 U14805 ( .A(n11632), .ZN(n51239) );
  NAND2_X1 U14812 ( .A1(n14750), .A2(n20484), .ZN(n20400) );
  NAND3_X1 U14813 ( .A1(n20405), .A2(n22090), .A3(n22085), .ZN(n3498) );
  OR2_X1 U14901 ( .A1(n47841), .A2(n42192), .ZN(n47814) );
  NAND2_X2 U15090 ( .A1(n265), .A2(n7785), .ZN(n30982) );
  AND3_X2 U15097 ( .A1(n6844), .A2(n17096), .A3(n6845), .ZN(n17420) );
  NAND3_X1 U15109 ( .A1(n4097), .A2(n27584), .A3(n2400), .ZN(n3997) );
  NOR2_X1 U15112 ( .A1(n6318), .A2(n38117), .ZN(n51241) );
  NAND2_X1 U15186 ( .A1(n21050), .A2(n2138), .ZN(n51242) );
  NAND2_X1 U15198 ( .A1(n51243), .A2(n12771), .ZN(n7716) );
  NAND3_X1 U15265 ( .A1(n12769), .A2(n13521), .A3(n13522), .ZN(n51243) );
  OR3_X1 U15285 ( .A1(n40558), .A2(n40316), .A3(n40572), .ZN(n40151) );
  XNOR2_X2 U15303 ( .A(n7999), .B(n25813), .ZN(n27420) );
  NAND4_X2 U15317 ( .A1(n22894), .A2(n22892), .A3(n22893), .A4(n22895), .ZN(
        n25813) );
  OAI21_X1 U15417 ( .B1(n14145), .B2(n51245), .A(n10310), .ZN(n1063) );
  NAND3_X1 U15430 ( .A1(n14150), .A2(n51175), .A3(n13761), .ZN(n51245) );
  NAND2_X1 U15446 ( .A1(n20461), .A2(n51246), .ZN(n19376) );
  NAND2_X1 U15510 ( .A1(n22874), .A2(n51156), .ZN(n22878) );
  XNOR2_X1 U15511 ( .A(n51247), .B(n48885), .ZN(Plaintext[81]) );
  NAND4_X1 U15513 ( .A1(n5887), .A2(n5886), .A3(n48883), .A4(n5888), .ZN(
        n51247) );
  NAND2_X1 U15514 ( .A1(n36547), .A2(n34089), .ZN(n36552) );
  OAI211_X1 U15522 ( .C1(n49226), .C2(n49203), .A(n51248), .B(n49212), .ZN(
        n43440) );
  NAND2_X1 U15578 ( .A1(n49222), .A2(n46215), .ZN(n51248) );
  NAND2_X1 U15582 ( .A1(n30606), .A2(n30605), .ZN(n150) );
  NAND2_X1 U15589 ( .A1(n755), .A2(n24290), .ZN(n2712) );
  XNOR2_X1 U15592 ( .A(n35339), .B(n36730), .ZN(n51249) );
  NAND2_X1 U15607 ( .A1(n21957), .A2(n51250), .ZN(n21164) );
  NAND2_X1 U15661 ( .A1(n23041), .A2(n4935), .ZN(n1170) );
  NAND2_X1 U15674 ( .A1(n20441), .A2(n19280), .ZN(n20826) );
  INV_X1 U15681 ( .A(n5176), .ZN(n13322) );
  NAND3_X1 U15682 ( .A1(n4950), .A2(n40558), .A3(n40156), .ZN(n40570) );
  OAI211_X2 U15690 ( .C1(n30838), .C2(n31302), .A(n30837), .B(n51252), .ZN(
        n35224) );
  INV_X1 U15700 ( .A(n31296), .ZN(n51252) );
  XNOR2_X1 U15711 ( .A(n51253), .B(n25084), .ZN(n25086) );
  XNOR2_X1 U15761 ( .A(n25083), .B(n25082), .ZN(n51253) );
  NAND2_X2 U15764 ( .A1(n51254), .A2(n20407), .ZN(n26395) );
  OAI22_X1 U15807 ( .A1(n3496), .A2(n3497), .B1(n424), .B2(n22943), .ZN(n51254) );
  NAND2_X1 U15810 ( .A1(n11378), .A2(n51255), .ZN(n11380) );
  NAND2_X1 U15814 ( .A1(n51256), .A2(n10702), .ZN(n51255) );
  INV_X1 U15841 ( .A(n30389), .ZN(n51257) );
  NAND2_X1 U15849 ( .A1(n28757), .A2(n51113), .ZN(n27528) );
  NAND2_X1 U15859 ( .A1(n14660), .A2(n12799), .ZN(n13996) );
  NAND2_X1 U15908 ( .A1(n51258), .A2(n39361), .ZN(n39362) );
  NOR2_X1 U15946 ( .A1(n1351), .A2(n13294), .ZN(n51259) );
  NAND2_X1 U16023 ( .A1(n31724), .A2(n32791), .ZN(n32782) );
  INV_X1 U16048 ( .A(n51261), .ZN(n5952) );
  OAI21_X1 U16052 ( .B1(n7144), .B2(n23732), .A(n24068), .ZN(n51261) );
  AND4_X2 U16053 ( .A1(n10275), .A2(n10260), .A3(n10276), .A4(n7594), .ZN(
        n14159) );
  NAND2_X1 U16066 ( .A1(n51262), .A2(n6332), .ZN(n15465) );
  NAND4_X1 U16078 ( .A1(n15403), .A2(n15402), .A3(n15401), .A4(n17471), .ZN(
        n51262) );
  NAND2_X1 U16080 ( .A1(n21543), .A2(n51485), .ZN(n20746) );
  NAND3_X1 U16148 ( .A1(n5054), .A2(n28952), .A3(n28497), .ZN(n28499) );
  NAND2_X1 U16170 ( .A1(n22262), .A2(n21730), .ZN(n21143) );
  NAND2_X1 U16197 ( .A1(n7422), .A2(n36896), .ZN(n37716) );
  INV_X1 U16227 ( .A(n17510), .ZN(n5528) );
  NAND2_X1 U16232 ( .A1(n847), .A2(n5529), .ZN(n17510) );
  NOR2_X1 U16250 ( .A1(n14441), .A2(n14440), .ZN(n14449) );
  XNOR2_X2 U16252 ( .A(n35255), .B(n33894), .ZN(n34535) );
  NAND3_X1 U16253 ( .A1(n51265), .A2(n12102), .A3(n51264), .ZN(n12103) );
  NAND2_X1 U16264 ( .A1(n4790), .A2(n4283), .ZN(n51265) );
  NAND2_X2 U16279 ( .A1(n5872), .A2(n38006), .ZN(n38015) );
  XNOR2_X1 U16294 ( .A(n43573), .B(n43574), .ZN(n51266) );
  NAND3_X1 U16314 ( .A1(n1), .A2(n2), .A3(n34802), .ZN(n34809) );
  NAND3_X1 U16321 ( .A1(n22261), .A2(n22263), .A3(n20868), .ZN(n42) );
  XNOR2_X1 U16330 ( .A(n51267), .B(n16246), .ZN(n16249) );
  XNOR2_X1 U16338 ( .A(n16240), .B(n16239), .ZN(n51267) );
  NAND3_X1 U16368 ( .A1(n21254), .A2(n19474), .A3(n18966), .ZN(n18967) );
  NAND2_X1 U16370 ( .A1(n3335), .A2(n19086), .ZN(n18966) );
  NOR2_X1 U16423 ( .A1(n51149), .A2(n51144), .ZN(n51269) );
  INV_X1 U16424 ( .A(n30584), .ZN(n31038) );
  NAND2_X1 U16454 ( .A1(n31039), .A2(n6107), .ZN(n30584) );
  NAND3_X1 U16465 ( .A1(n26669), .A2(n29486), .A3(n51159), .ZN(n26670) );
  NAND2_X2 U16499 ( .A1(n51270), .A2(n37215), .ZN(n40446) );
  AND3_X1 U16526 ( .A1(n37217), .A2(n37216), .A3(n37214), .ZN(n51270) );
  NAND2_X1 U16550 ( .A1(n51271), .A2(n39744), .ZN(n7662) );
  NAND2_X1 U16570 ( .A1(n51272), .A2(n41670), .ZN(n40714) );
  NAND2_X1 U16572 ( .A1(n40709), .A2(n40708), .ZN(n51272) );
  NAND3_X1 U16576 ( .A1(n38310), .A2(n38311), .A3(n51273), .ZN(n38312) );
  NAND2_X1 U16584 ( .A1(n37659), .A2(n38317), .ZN(n38310) );
  NAND2_X1 U16587 ( .A1(n47198), .A2(n51274), .ZN(n2694) );
  NAND2_X1 U16590 ( .A1(n49521), .A2(n43490), .ZN(n45022) );
  NAND3_X1 U16607 ( .A1(n3739), .A2(n46175), .A3(n46176), .ZN(n46177) );
  XNOR2_X1 U16636 ( .A(n51278), .B(n42585), .ZN(n42589) );
  XNOR2_X1 U16669 ( .A(n42577), .B(n42578), .ZN(n51278) );
  NAND3_X1 U16698 ( .A1(n22135), .A2(n23242), .A3(n23255), .ZN(n22136) );
  NAND4_X2 U16735 ( .A1(n12209), .A2(n12210), .A3(n12208), .A4(n12207), .ZN(
        n18447) );
  NAND2_X1 U16738 ( .A1(n1168), .A2(n32717), .ZN(n31977) );
  XNOR2_X1 U16745 ( .A(n24792), .B(n23879), .ZN(n23794) );
  XNOR2_X2 U16753 ( .A(n7939), .B(n24791), .ZN(n23879) );
  NOR2_X1 U16826 ( .A1(n12676), .A2(n11872), .ZN(n12455) );
  NAND2_X1 U16836 ( .A1(n12675), .A2(n592), .ZN(n11872) );
  NAND3_X1 U16842 ( .A1(n15343), .A2(n15438), .A3(n15341), .ZN(n14864) );
  NAND2_X1 U16847 ( .A1(n21293), .A2(n509), .ZN(n19716) );
  AND2_X2 U16857 ( .A1(n19711), .A2(n3685), .ZN(n21293) );
  BUF_X1 U16929 ( .A(n12338), .Z(n51462) );
  NAND2_X1 U16968 ( .A1(n35981), .A2(n35980), .ZN(n51281) );
  NAND2_X1 U16978 ( .A1(n35982), .A2(n37597), .ZN(n51282) );
  XNOR2_X1 U16990 ( .A(n43890), .B(n44963), .ZN(n43598) );
  NAND3_X1 U17073 ( .A1(n39891), .A2(n40737), .A3(n40740), .ZN(n6475) );
  NAND3_X1 U17074 ( .A1(n3823), .A2(n23378), .A3(n3821), .ZN(n22238) );
  NAND3_X1 U17151 ( .A1(n10704), .A2(n51256), .A3(n51391), .ZN(n9641) );
  NAND2_X1 U17154 ( .A1(n3254), .A2(n12750), .ZN(n13646) );
  NAND2_X1 U17160 ( .A1(n903), .A2(n23560), .ZN(n23561) );
  NOR2_X1 U17176 ( .A1(n9743), .A2(n11005), .ZN(n51605) );
  XNOR2_X1 U17268 ( .A(n51284), .B(n28249), .ZN(n25477) );
  XNOR2_X1 U17269 ( .A(n25466), .B(n25465), .ZN(n51284) );
  BUF_X1 U17294 ( .A(n47868), .Z(n372) );
  XNOR2_X1 U17383 ( .A(n1512), .B(n35761), .ZN(n35488) );
  NOR2_X1 U17447 ( .A1(n46684), .A2(n46683), .ZN(n51286) );
  NOR2_X1 U17456 ( .A1(n46684), .A2(n46683), .ZN(n51287) );
  NOR2_X1 U17483 ( .A1(n46684), .A2(n46683), .ZN(n414) );
  OR2_X1 U17541 ( .A1(n5443), .A2(n38132), .ZN(n38053) );
  NAND2_X1 U17694 ( .A1(n5787), .A2(n3473), .ZN(n51290) );
  NAND3_X1 U17716 ( .A1(n46718), .A2(n5410), .A3(n7127), .ZN(n47554) );
  AND3_X1 U17722 ( .A1(n26820), .A2(n26822), .A3(n26821), .ZN(n26848) );
  NOR2_X1 U17723 ( .A1(n41049), .A2(n41058), .ZN(n40494) );
  NAND4_X1 U17728 ( .A1(n914), .A2(n2949), .A3(n919), .A4(n917), .ZN(n51469)
         );
  NOR2_X1 U17745 ( .A1(n32985), .A2(n32984), .ZN(n32994) );
  INV_X1 U17746 ( .A(n31497), .ZN(n31488) );
  AND3_X1 U17747 ( .A1(n46470), .A2(n46469), .A3(n46468), .ZN(n51291) );
  XNOR2_X1 U17794 ( .A(n52196), .B(n44084), .ZN(n51292) );
  XNOR2_X1 U17796 ( .A(n52196), .B(n44084), .ZN(n46816) );
  AND2_X1 U17853 ( .A1(n14633), .A2(n12755), .ZN(n12753) );
  NAND4_X1 U17863 ( .A1(n6575), .A2(n6574), .A3(n2260), .A4(n47348), .ZN(
        n50744) );
  XNOR2_X1 U17929 ( .A(n42916), .B(n42917), .ZN(n49720) );
  AND4_X1 U17939 ( .A1(n8628), .A2(n47148), .A3(n47147), .A4(n8668), .ZN(
        n50780) );
  XNOR2_X1 U17941 ( .A(n39849), .B(n44164), .ZN(n44960) );
  AND2_X1 U18028 ( .A1(n46034), .A2(n50292), .ZN(n50299) );
  NAND4_X1 U18055 ( .A1(n45152), .A2(n45151), .A3(n45149), .A4(n45150), .ZN(
        n51298) );
  NAND4_X1 U18060 ( .A1(n45152), .A2(n45151), .A3(n45149), .A4(n45150), .ZN(
        n51299) );
  XNOR2_X1 U18063 ( .A(n43038), .B(n43037), .ZN(n51300) );
  CLKBUF_X1 U18089 ( .A(n48481), .Z(n51301) );
  XNOR2_X1 U18103 ( .A(n44346), .B(n44345), .ZN(n48481) );
  NAND2_X1 U18105 ( .A1(n41378), .A2(n41375), .ZN(n40924) );
  NAND4_X1 U18119 ( .A1(n46727), .A2(n46728), .A3(n46729), .A4(n46726), .ZN(
        n51302) );
  NAND4_X1 U18122 ( .A1(n46727), .A2(n46728), .A3(n46729), .A4(n46726), .ZN(
        n51303) );
  NAND4_X1 U18125 ( .A1(n46727), .A2(n46728), .A3(n46729), .A4(n46726), .ZN(
        n47547) );
  OR2_X1 U18129 ( .A1(n50486), .A2(n50483), .ZN(n50401) );
  NAND4_X2 U18150 ( .A1(n2567), .A2(n2566), .A3(n2565), .A4(n44593), .ZN(
        n50679) );
  INV_X1 U18151 ( .A(n661), .ZN(n51304) );
  XNOR2_X1 U18211 ( .A(n44036), .B(n44037), .ZN(n46828) );
  NOR2_X1 U18223 ( .A1(n36533), .A2(n51305), .ZN(n2389) );
  NAND2_X1 U18225 ( .A1(n51306), .A2(n36348), .ZN(n51305) );
  OR2_X1 U18226 ( .A1(n37982), .A2(n36524), .ZN(n51306) );
  NOR2_X2 U18276 ( .A1(n46647), .A2(n46646), .ZN(n46668) );
  AND2_X1 U18284 ( .A1(n49365), .A2(n49370), .ZN(n51308) );
  AND2_X1 U18305 ( .A1(n4903), .A2(n49343), .ZN(n51309) );
  AND2_X1 U18332 ( .A1(n49365), .A2(n49370), .ZN(n1879) );
  OAI21_X1 U18364 ( .B1(n49805), .B2(n49753), .A(n49853), .ZN(n51314) );
  NAND2_X1 U18399 ( .A1(n7311), .A2(n3300), .ZN(n51315) );
  NAND2_X1 U18498 ( .A1(n7311), .A2(n3300), .ZN(n51316) );
  NAND2_X1 U18512 ( .A1(n7311), .A2(n3300), .ZN(n49457) );
  INV_X1 U18519 ( .A(n3155), .ZN(n51317) );
  XNOR2_X1 U18525 ( .A(n4888), .B(n41307), .ZN(n46597) );
  AND2_X1 U18591 ( .A1(n49126), .A2(n44772), .ZN(n51320) );
  INV_X1 U18615 ( .A(n51102), .ZN(n51322) );
  XNOR2_X1 U18624 ( .A(n36937), .B(n36938), .ZN(n38957) );
  AND2_X1 U18700 ( .A1(n1312), .A2(n50487), .ZN(n51598) );
  AND2_X1 U18701 ( .A1(n14962), .A2(n15278), .ZN(n15273) );
  NAND4_X1 U18711 ( .A1(n39498), .A2(n39496), .A3(n39495), .A4(n39497), .ZN(
        n51323) );
  AND3_X1 U18721 ( .A1(n32083), .A2(n4261), .A3(n32069), .ZN(n5778) );
  XOR2_X1 U18740 ( .A(n7126), .B(n34131), .Z(n51324) );
  NAND4_X1 U18792 ( .A1(n36024), .A2(n36026), .A3(n36025), .A4(n36023), .ZN(
        n40121) );
  OR2_X1 U18815 ( .A1(n49850), .A2(n49854), .ZN(n49793) );
  XNOR2_X1 U18893 ( .A(n43129), .B(n43128), .ZN(n51326) );
  NOR2_X1 U18946 ( .A1(n50462), .A2(n50461), .ZN(n51327) );
  NAND3_X1 U18977 ( .A1(n6549), .A2(n6548), .A3(n41154), .ZN(n51329) );
  NAND3_X1 U18994 ( .A1(n6549), .A2(n6548), .A3(n41154), .ZN(n51330) );
  AND2_X1 U19016 ( .A1(n51382), .A2(n48633), .ZN(n51331) );
  NAND2_X1 U19034 ( .A1(n49915), .A2(n51332), .ZN(n1077) );
  AND2_X1 U19075 ( .A1(n49923), .A2(n49916), .ZN(n51332) );
  INV_X1 U19078 ( .A(n37219), .ZN(n38257) );
  AND2_X1 U19117 ( .A1(n37741), .A2(n37742), .ZN(n148) );
  NAND4_X2 U19142 ( .A1(n47117), .A2(n8766), .A3(n47116), .A4(n47115), .ZN(
        n50772) );
  XNOR2_X1 U19177 ( .A(n42066), .B(n43123), .ZN(n43833) );
  XNOR2_X1 U19238 ( .A(n34612), .B(n34611), .ZN(n51334) );
  XNOR2_X1 U19376 ( .A(n34612), .B(n34611), .ZN(n36405) );
  AND2_X1 U19383 ( .A1(n45670), .A2(n49272), .ZN(n51335) );
  AND2_X1 U19414 ( .A1(n45670), .A2(n49272), .ZN(n45667) );
  XOR2_X1 U19425 ( .A(n13893), .B(n18193), .Z(n51336) );
  OAI21_X1 U19430 ( .B1(n40672), .B2(n39674), .A(n39673), .ZN(n51620) );
  OR2_X1 U19432 ( .A1(n36528), .A2(n36527), .ZN(n1740) );
  NAND2_X1 U19443 ( .A1(n42089), .A2(n7646), .ZN(n51337) );
  NAND2_X1 U19476 ( .A1(n42089), .A2(n7646), .ZN(n51338) );
  NAND2_X1 U19485 ( .A1(n42089), .A2(n7646), .ZN(n44042) );
  XNOR2_X1 U19517 ( .A(n34502), .B(n34501), .ZN(n51339) );
  OR2_X1 U19525 ( .A1(n50224), .A2(n50225), .ZN(n51565) );
  XOR2_X1 U19561 ( .A(n27311), .B(n26021), .Z(n26023) );
  XNOR2_X1 U19608 ( .A(n242), .B(n36701), .ZN(n36705) );
  NOR2_X1 U19609 ( .A1(n47744), .A2(n47782), .ZN(n47754) );
  AND4_X1 U19657 ( .A1(n38220), .A2(n38216), .A3(n38215), .A4(n38219), .ZN(
        n38224) );
  BUF_X1 U19659 ( .A(n5262), .Z(n2100) );
  INV_X1 U19660 ( .A(n5262), .ZN(n8480) );
  INV_X1 U19672 ( .A(n7044), .ZN(n51341) );
  XNOR2_X1 U19682 ( .A(n44553), .B(n44552), .ZN(n46869) );
  BUF_X1 U19689 ( .A(n29719), .Z(n51342) );
  INV_X1 U19731 ( .A(n36405), .ZN(n37649) );
  NAND4_X1 U19794 ( .A1(n44284), .A2(n44285), .A3(n3054), .A4(n3051), .ZN(
        n48033) );
  INV_X1 U19889 ( .A(n14666), .ZN(n51347) );
  INV_X1 U19914 ( .A(n14666), .ZN(n14665) );
  INV_X1 U19959 ( .A(n41063), .ZN(n51348) );
  AND2_X1 U19971 ( .A1(n50533), .A2(n50552), .ZN(n51349) );
  NOR2_X1 U19993 ( .A1(n51297), .A2(n40014), .ZN(n40002) );
  OAI21_X1 U20009 ( .B1(n48422), .B2(n48421), .A(n48420), .ZN(n51350) );
  OAI21_X1 U20023 ( .B1(n48422), .B2(n48421), .A(n48420), .ZN(n48606) );
  CLKBUF_X1 U20041 ( .A(n24675), .Z(n51351) );
  NAND2_X1 U20049 ( .A1(n6564), .A2(n47084), .ZN(n51353) );
  NAND2_X1 U20059 ( .A1(n6564), .A2(n47084), .ZN(n51354) );
  NAND2_X1 U20079 ( .A1(n6564), .A2(n47084), .ZN(n50771) );
  INV_X1 U20157 ( .A(n8104), .ZN(n51356) );
  OR2_X1 U20228 ( .A1(n1835), .A2(n19535), .ZN(n17021) );
  OR2_X1 U20277 ( .A1(n41352), .A2(n41354), .ZN(n40749) );
  AND2_X1 U20391 ( .A1(n654), .A2(n49932), .ZN(n49905) );
  AND2_X1 U20410 ( .A1(n31536), .A2(n32666), .ZN(n51588) );
  NAND4_X1 U20459 ( .A1(n37495), .A2(n37494), .A3(n37493), .A4(n37492), .ZN(
        n51357) );
  NAND4_X1 U20472 ( .A1(n37495), .A2(n37494), .A3(n37493), .A4(n37492), .ZN(
        n51358) );
  XNOR2_X1 U20475 ( .A(n44898), .B(n44897), .ZN(n51359) );
  XNOR2_X1 U20498 ( .A(n44898), .B(n44897), .ZN(n46686) );
  OR2_X1 U20559 ( .A1(n32909), .A2(n32895), .ZN(n31603) );
  XNOR2_X1 U20586 ( .A(n35245), .B(n35244), .ZN(n51360) );
  BUF_X1 U20649 ( .A(n44826), .Z(n45534) );
  CLKBUF_X1 U20656 ( .A(n6603), .Z(n51361) );
  XNOR2_X1 U20673 ( .A(n46150), .B(n42961), .ZN(n7592) );
  AND2_X1 U20719 ( .A1(n40447), .A2(n40450), .ZN(n40404) );
  INV_X1 U20811 ( .A(n37439), .ZN(n51363) );
  OR2_X1 U20843 ( .A1(n41328), .A2(n41332), .ZN(n51364) );
  NAND2_X1 U20901 ( .A1(n46905), .A2(n51365), .ZN(n4996) );
  AND2_X1 U20906 ( .A1(n46693), .A2(n51359), .ZN(n51365) );
  XNOR2_X1 U20918 ( .A(n3966), .B(n28263), .ZN(n28298) );
  INV_X1 U20922 ( .A(n50727), .ZN(n51367) );
  XNOR2_X1 U20932 ( .A(n5616), .B(n34361), .ZN(n35678) );
  BUF_X1 U20969 ( .A(n46153), .Z(n51368) );
  XNOR2_X1 U21036 ( .A(n44176), .B(n41875), .ZN(n46153) );
  NAND4_X1 U21063 ( .A1(n51611), .A2(n10840), .A3(n10839), .A4(n51610), .ZN(
        n51369) );
  NAND4_X1 U21074 ( .A1(n51611), .A2(n10840), .A3(n10839), .A4(n51610), .ZN(
        n51370) );
  NAND4_X1 U21132 ( .A1(n51611), .A2(n10840), .A3(n10839), .A4(n51610), .ZN(
        n14123) );
  AND2_X1 U21134 ( .A1(n12514), .A2(n12516), .ZN(n10832) );
  OR2_X1 U21135 ( .A1(n12057), .A2(n10662), .ZN(n12059) );
  AOI21_X1 U21136 ( .B1(n29280), .B2(n5522), .A(n871), .ZN(n29197) );
  BUF_X1 U21217 ( .A(n50270), .Z(n51372) );
  XNOR2_X1 U21261 ( .A(n15272), .B(n15271), .ZN(n51374) );
  NAND4_X2 U21262 ( .A1(n37769), .A2(n37771), .A3(n37772), .A4(n37770), .ZN(
        n51375) );
  AND2_X1 U21389 ( .A1(n49177), .A2(n539), .ZN(n51376) );
  NAND4_X2 U21570 ( .A1(n35886), .A2(n35885), .A3(n35884), .A4(n35883), .ZN(
        n51377) );
  NAND2_X1 U21571 ( .A1(n4961), .A2(n11770), .ZN(n51378) );
  NAND2_X1 U21700 ( .A1(n4961), .A2(n11770), .ZN(n51379) );
  NOR2_X2 U21807 ( .A1(n4963), .A2(n4962), .ZN(n4961) );
  NAND2_X1 U21809 ( .A1(n4961), .A2(n11770), .ZN(n18738) );
  XNOR2_X1 U22064 ( .A(n27419), .B(n25947), .ZN(n26567) );
  INV_X1 U22134 ( .A(n6481), .ZN(n51383) );
  OAI21_X1 U22178 ( .B1(n14100), .B2(n14453), .A(n14096), .ZN(n51384) );
  INV_X1 U22236 ( .A(n6481), .ZN(n14100) );
  NAND3_X2 U22237 ( .A1(n7003), .A2(n6478), .A3(n11397), .ZN(n14453) );
  INV_X1 U22302 ( .A(n14342), .ZN(n13417) );
  XOR2_X1 U22316 ( .A(n16984), .B(n16983), .Z(n51385) );
  XOR2_X1 U22322 ( .A(n51663), .B(n33583), .Z(n35603) );
  NAND4_X2 U22478 ( .A1(n17986), .A2(n17985), .A3(n5920), .A4(n5921), .ZN(
        n22901) );
  NOR2_X1 U22651 ( .A1(n33026), .A2(n32874), .ZN(n32877) );
  XNOR2_X1 U22721 ( .A(n43861), .B(n43860), .ZN(n50343) );
  OR2_X1 U22736 ( .A1(n50906), .A2(n51299), .ZN(n51388) );
  NAND4_X1 U22767 ( .A1(n36182), .A2(n36185), .A3(n36184), .A4(n36183), .ZN(
        n45399) );
  INV_X1 U22822 ( .A(n39035), .ZN(n51389) );
  XNOR2_X1 U22839 ( .A(n3526), .B(n45408), .ZN(n51390) );
  XNOR2_X1 U22931 ( .A(n3526), .B(n45408), .ZN(n43856) );
  NOR2_X1 U22932 ( .A1(n29221), .A2(n1708), .ZN(n27913) );
  NAND4_X1 U22969 ( .A1(n39961), .A2(n5476), .A3(n39959), .A4(n39960), .ZN(
        n51392) );
  NAND4_X1 U23002 ( .A1(n39961), .A2(n5476), .A3(n39959), .A4(n39960), .ZN(
        n51393) );
  XNOR2_X1 U23023 ( .A(n9402), .B(Key[167]), .ZN(n11361) );
  NAND4_X1 U23039 ( .A1(n39961), .A2(n5476), .A3(n39959), .A4(n39960), .ZN(
        n5108) );
  INV_X1 U23158 ( .A(n40967), .ZN(n40963) );
  XNOR2_X1 U23182 ( .A(n41468), .B(n41467), .ZN(n46708) );
  INV_X1 U23351 ( .A(n49029), .ZN(n653) );
  NAND4_X1 U23406 ( .A1(n46621), .A2(n46618), .A3(n46619), .A4(n46620), .ZN(
        n51400) );
  NAND4_X1 U23448 ( .A1(n46621), .A2(n46618), .A3(n46619), .A4(n46620), .ZN(
        n51401) );
  XNOR2_X1 U23468 ( .A(n44970), .B(n44969), .ZN(n46691) );
  NAND4_X1 U23525 ( .A1(n46621), .A2(n46618), .A3(n46619), .A4(n46620), .ZN(
        n47596) );
  OR2_X1 U23556 ( .A1(n49932), .A2(n49916), .ZN(n49877) );
  INV_X1 U23613 ( .A(n16546), .ZN(n51403) );
  AND2_X1 U23614 ( .A1(n44583), .A2(n47058), .ZN(n50276) );
  NOR2_X1 U23807 ( .A1(n31749), .A2(n31740), .ZN(n31849) );
  BUF_X1 U23842 ( .A(n46810), .Z(n51404) );
  XNOR2_X1 U23868 ( .A(n44023), .B(n44022), .ZN(n46810) );
  OAI211_X1 U23985 ( .C1(n5064), .C2(n5063), .A(n5062), .B(n5059), .ZN(n43000)
         );
  XNOR2_X1 U23990 ( .A(n15668), .B(n15669), .ZN(n51407) );
  NAND3_X1 U24098 ( .A1(n270), .A2(n1185), .A3(n8721), .ZN(n45386) );
  NOR2_X1 U24183 ( .A1(n50710), .A2(n50685), .ZN(n50693) );
  BUF_X2 U24204 ( .A(n50383), .Z(n2198) );
  XNOR2_X1 U24260 ( .A(n43918), .B(n43919), .ZN(n51410) );
  XNOR2_X1 U24295 ( .A(n45426), .B(n45284), .ZN(n46069) );
  XNOR2_X1 U24385 ( .A(n43918), .B(n43919), .ZN(n50265) );
  XNOR2_X1 U24493 ( .A(n35758), .B(n4492), .ZN(n37484) );
  OAI211_X1 U24619 ( .C1(n31593), .C2(n31592), .A(n31591), .B(n31590), .ZN(
        n51413) );
  OAI211_X1 U24645 ( .C1(n31593), .C2(n31592), .A(n31591), .B(n31590), .ZN(
        n34812) );
  NAND4_X1 U24883 ( .A1(n2069), .A2(n2068), .A3(n24045), .A4(n24044), .ZN(
        n51415) );
  NAND4_X1 U24884 ( .A1(n2069), .A2(n2068), .A3(n24045), .A4(n24044), .ZN(
        n51416) );
  XNOR2_X1 U24948 ( .A(n51415), .B(n26147), .ZN(n26292) );
  AND2_X1 U25135 ( .A1(n49126), .A2(n1501), .ZN(n49113) );
  XNOR2_X1 U25187 ( .A(n19260), .B(n17972), .ZN(n51417) );
  XNOR2_X1 U25283 ( .A(n19260), .B(n17972), .ZN(n560) );
  XNOR2_X1 U25284 ( .A(n33603), .B(n51381), .ZN(n51418) );
  INV_X1 U25313 ( .A(n7047), .ZN(n51419) );
  XNOR2_X1 U25314 ( .A(n7870), .B(n44054), .ZN(n44109) );
  XNOR2_X1 U25318 ( .A(n43357), .B(n46138), .ZN(n51420) );
  XNOR2_X1 U25341 ( .A(n43357), .B(n46138), .ZN(n43725) );
  XNOR2_X1 U25360 ( .A(n25464), .B(n27197), .ZN(n25680) );
  INV_X1 U25676 ( .A(n34067), .ZN(n51422) );
  XNOR2_X1 U25750 ( .A(n33943), .B(n36991), .ZN(n37323) );
  XNOR2_X1 U25751 ( .A(n35488), .B(n37323), .ZN(n35404) );
  NAND2_X1 U25857 ( .A1(n4658), .A2(n4447), .ZN(n51423) );
  NAND2_X1 U25906 ( .A1(n4658), .A2(n4447), .ZN(n51424) );
  NAND2_X1 U25907 ( .A1(n4658), .A2(n4447), .ZN(n28060) );
  CLKBUF_X1 U25974 ( .A(n46648), .Z(n51425) );
  NOR2_X1 U26066 ( .A1(n38998), .A2(n34906), .ZN(n38995) );
  INV_X1 U26104 ( .A(n45219), .ZN(n51426) );
  XNOR2_X1 U26425 ( .A(n42888), .B(n4704), .ZN(n46498) );
  NAND4_X1 U27623 ( .A1(n30548), .A2(n30547), .A3(n30546), .A4(n30545), .ZN(
        n3524) );
  XNOR2_X1 U27633 ( .A(n35631), .B(n35630), .ZN(n51429) );
  XNOR2_X1 U27717 ( .A(n35630), .B(n35631), .ZN(n38587) );
  NAND3_X1 U27758 ( .A1(n36140), .A2(n36139), .A3(n36138), .ZN(n41195) );
  OAI21_X1 U27798 ( .B1(n8109), .B2(n8107), .A(n7366), .ZN(n51431) );
  OAI21_X1 U27851 ( .B1(n8109), .B2(n8107), .A(n7366), .ZN(n46120) );
  AND2_X1 U27899 ( .A1(n11501), .A2(n11884), .ZN(n12673) );
  AND2_X1 U27998 ( .A1(n12458), .A2(n11501), .ZN(n12671) );
  XNOR2_X1 U28001 ( .A(Key[115]), .B(Ciphertext[18]), .ZN(n51432) );
  XNOR2_X1 U28006 ( .A(Key[115]), .B(Ciphertext[18]), .ZN(n51433) );
  XNOR2_X1 U28009 ( .A(Key[115]), .B(Ciphertext[18]), .ZN(n12626) );
  XNOR2_X1 U28374 ( .A(n17193), .B(n17192), .ZN(n19839) );
  NAND4_X1 U28411 ( .A1(n13287), .A2(n13285), .A3(n13286), .A4(n13284), .ZN(
        n51435) );
  NAND4_X1 U28672 ( .A1(n13287), .A2(n13285), .A3(n13286), .A4(n13284), .ZN(
        n51436) );
  XNOR2_X1 U28728 ( .A(n18404), .B(n17707), .ZN(n51437) );
  XNOR2_X1 U29020 ( .A(n18404), .B(n17707), .ZN(n51438) );
  NAND4_X1 U29058 ( .A1(n13287), .A2(n13285), .A3(n13286), .A4(n13284), .ZN(
        n18404) );
  XNOR2_X1 U29446 ( .A(n44535), .B(n44189), .ZN(n51439) );
  XNOR2_X1 U29466 ( .A(n44535), .B(n44189), .ZN(n43914) );
  NOR2_X1 U29482 ( .A1(n18376), .A2(n20037), .ZN(n51440) );
  BUF_X1 U29520 ( .A(n25131), .Z(n51441) );
  NOR2_X1 U29540 ( .A1(n18376), .A2(n20037), .ZN(n18374) );
  XNOR2_X1 U29544 ( .A(n26285), .B(n28257), .ZN(n25131) );
  AND3_X1 U29584 ( .A1(n50018), .A2(n6413), .A3(n50017), .ZN(n50128) );
  XNOR2_X1 U29780 ( .A(n43063), .B(n44534), .ZN(n51444) );
  NAND4_X1 U29798 ( .A1(n32892), .A2(n32893), .A3(n32891), .A4(n32890), .ZN(
        n51445) );
  NAND4_X1 U29816 ( .A1(n32892), .A2(n32893), .A3(n32891), .A4(n32890), .ZN(
        n35240) );
  NAND4_X1 U29914 ( .A1(n28946), .A2(n28945), .A3(n28944), .A4(n28943), .ZN(
        n51446) );
  NAND4_X1 U30014 ( .A1(n28946), .A2(n28945), .A3(n28944), .A4(n28943), .ZN(
        n51447) );
  XOR2_X1 U30041 ( .A(n41629), .B(n6573), .Z(n51448) );
  XNOR2_X1 U30255 ( .A(n35543), .B(n32310), .ZN(n35635) );
  XNOR2_X1 U30292 ( .A(n51099), .B(n43950), .ZN(n51450) );
  BUF_X1 U30330 ( .A(n52039), .Z(n51451) );
  INV_X1 U30341 ( .A(n31816), .ZN(n31034) );
  INV_X1 U30387 ( .A(n49465), .ZN(n51453) );
  XNOR2_X1 U30388 ( .A(n15619), .B(n17954), .ZN(n51454) );
  XNOR2_X1 U30391 ( .A(n15619), .B(n17954), .ZN(n18480) );
  OR3_X2 U30401 ( .A1(n4420), .A2(n2238), .A3(n2380), .ZN(n15619) );
  OR2_X1 U30409 ( .A1(n12450), .A2(n50997), .ZN(n12469) );
  XNOR2_X1 U30592 ( .A(n8293), .B(n44055), .ZN(n46830) );
  XNOR2_X1 U30980 ( .A(n16011), .B(n16711), .ZN(n17671) );
  INV_X1 U31134 ( .A(n33470), .ZN(n51463) );
  NAND4_X1 U31233 ( .A1(n38858), .A2(n6713), .A3(n38857), .A4(n38856), .ZN(
        n51465) );
  INV_X1 U31480 ( .A(n47795), .ZN(n51467) );
  INV_X1 U31600 ( .A(n47795), .ZN(n51468) );
  INV_X1 U31770 ( .A(n47795), .ZN(n47778) );
  NAND4_X1 U31897 ( .A1(n914), .A2(n2949), .A3(n919), .A4(n917), .ZN(n51470)
         );
  NAND4_X1 U31938 ( .A1(n914), .A2(n2949), .A3(n919), .A4(n917), .ZN(n47869)
         );
  AND4_X1 U31939 ( .A1(n51542), .A2(n30276), .A3(n51541), .A4(n30275), .ZN(
        n51471) );
  XNOR2_X1 U31966 ( .A(n7624), .B(n36672), .ZN(n51472) );
  XNOR2_X1 U31973 ( .A(n7624), .B(n36672), .ZN(n34829) );
  INV_X1 U31986 ( .A(n51726), .ZN(n51473) );
  XNOR2_X1 U31989 ( .A(n1499), .B(n1498), .ZN(n29159) );
  XNOR2_X1 U32012 ( .A(n5474), .B(n34840), .ZN(n51474) );
  NAND4_X1 U32515 ( .A1(n6029), .A2(n42406), .A3(n6030), .A4(n6028), .ZN(
        n48944) );
  BUF_X1 U32867 ( .A(n16926), .Z(n51481) );
  XNOR2_X1 U33194 ( .A(n25494), .B(n23525), .ZN(n51483) );
  XNOR2_X1 U33386 ( .A(n25494), .B(n23525), .ZN(n51484) );
  XNOR2_X1 U33944 ( .A(n16016), .B(n16450), .ZN(n16926) );
  XNOR2_X1 U33945 ( .A(n25494), .B(n23525), .ZN(n27257) );
  NOR2_X1 U34362 ( .A1(n47786), .A2(n45877), .ZN(n644) );
  XOR2_X1 U34367 ( .A(n7813), .B(n18417), .Z(n51485) );
  INV_X1 U34368 ( .A(n50958), .ZN(n51486) );
  INV_X1 U34411 ( .A(n50958), .ZN(n50951) );
  AND2_X1 U34412 ( .A1(n27638), .A2(n27633), .ZN(n26888) );
  XNOR2_X1 U34636 ( .A(n35564), .B(n35565), .ZN(n51487) );
  BUF_X1 U34766 ( .A(n45804), .Z(n51488) );
  XNOR2_X1 U34769 ( .A(n35564), .B(n35565), .ZN(n37488) );
  XNOR2_X1 U34835 ( .A(n41595), .B(n41594), .ZN(n45804) );
  XNOR2_X1 U34836 ( .A(n28229), .B(n28348), .ZN(n51489) );
  XNOR2_X1 U34888 ( .A(n28229), .B(n28348), .ZN(n51490) );
  XNOR2_X1 U34912 ( .A(n28348), .B(n28229), .ZN(n30344) );
  XNOR2_X1 U34914 ( .A(n5612), .B(n8087), .ZN(n51493) );
  NAND4_X1 U35149 ( .A1(n37615), .A2(n37614), .A3(n37613), .A4(n41020), .ZN(
        n51498) );
  XNOR2_X1 U35166 ( .A(n33702), .B(n33973), .ZN(n37277) );
  XNOR2_X1 U35293 ( .A(n27177), .B(n7103), .ZN(n51502) );
  XNOR2_X1 U35310 ( .A(n42822), .B(n42819), .ZN(n51503) );
  XNOR2_X1 U35481 ( .A(n27177), .B(n7103), .ZN(n25215) );
  XNOR2_X1 U35586 ( .A(n42819), .B(n42822), .ZN(n45321) );
  NAND2_X1 U35587 ( .A1(n3479), .A2(n39027), .ZN(n39453) );
  INV_X1 U35630 ( .A(n52131), .ZN(n51504) );
  XNOR2_X1 U35817 ( .A(n43066), .B(n43067), .ZN(n49635) );
  INV_X1 U36000 ( .A(n51736), .ZN(n51507) );
  XNOR2_X1 U36042 ( .A(n3061), .B(n37282), .ZN(n39235) );
  XNOR2_X1 U36235 ( .A(n37312), .B(n37313), .ZN(n39224) );
  CLKBUF_X1 U36274 ( .A(n42662), .Z(n51509) );
  NAND2_X1 U36368 ( .A1(n42515), .A2(n42516), .ZN(n51510) );
  NAND2_X1 U36372 ( .A1(n42515), .A2(n42516), .ZN(n51511) );
  NAND2_X1 U36452 ( .A1(n42515), .A2(n42516), .ZN(n48975) );
  OR2_X1 U36527 ( .A1(n50314), .A2(n50317), .ZN(n50316) );
  BUF_X1 U36551 ( .A(n25352), .Z(n51512) );
  XOR2_X1 U36599 ( .A(n24914), .B(n24913), .Z(n51514) );
  XNOR2_X1 U36626 ( .A(n193), .B(n43396), .ZN(n51515) );
  OR2_X1 U36653 ( .A1(n52107), .A2(n49442), .ZN(n51516) );
  XNOR2_X1 U36678 ( .A(n193), .B(n43396), .ZN(n49154) );
  XNOR2_X1 U36859 ( .A(n6808), .B(n6807), .ZN(n51517) );
  XNOR2_X1 U37116 ( .A(n6808), .B(n6807), .ZN(n51518) );
  XNOR2_X1 U37161 ( .A(n6808), .B(n6807), .ZN(n29288) );
  NAND4_X1 U37310 ( .A1(n29197), .A2(n29196), .A3(n846), .A4(n29195), .ZN(
        n51519) );
  NAND4_X1 U37312 ( .A1(n29197), .A2(n29196), .A3(n846), .A4(n29195), .ZN(
        n32401) );
  XNOR2_X1 U37317 ( .A(n31508), .B(n34476), .ZN(n51522) );
  XNOR2_X1 U37399 ( .A(n16913), .B(n12401), .ZN(n18196) );
  XNOR2_X1 U37400 ( .A(n34476), .B(n31508), .ZN(n38135) );
  BUF_X2 U37507 ( .A(n43558), .Z(n51525) );
  XNOR2_X1 U37513 ( .A(n43562), .B(n2371), .ZN(n51526) );
  OAI211_X1 U37711 ( .C1(n31353), .C2(n36147), .A(n31352), .B(n3586), .ZN(
        n31354) );
  NAND3_X1 U37913 ( .A1(n38550), .A2(n38549), .A3(n38228), .ZN(n3586) );
  NAND3_X1 U38051 ( .A1(n12099), .A2(n12098), .A3(n10687), .ZN(n10689) );
  INV_X1 U38078 ( .A(n8782), .ZN(n10200) );
  XNOR2_X1 U38254 ( .A(n41879), .B(n41878), .ZN(n51529) );
  NAND2_X1 U38268 ( .A1(n6274), .A2(n6275), .ZN(n13631) );
  NAND2_X1 U38413 ( .A1(n20120), .A2(n20121), .ZN(n20127) );
  NAND3_X1 U38426 ( .A1(n11593), .A2(n11600), .A3(n9279), .ZN(n10805) );
  NAND2_X1 U38517 ( .A1(n51530), .A2(n21296), .ZN(n18892) );
  NAND3_X1 U38560 ( .A1(n21290), .A2(n19715), .A3(n18883), .ZN(n51530) );
  NAND2_X1 U38700 ( .A1(n5099), .A2(n13377), .ZN(n13371) );
  AND2_X1 U38709 ( .A1(n11723), .A2(n16036), .ZN(n5099) );
  NAND3_X2 U39023 ( .A1(n39068), .A2(n4748), .A3(n7417), .ZN(n46068) );
  INV_X1 U39031 ( .A(n644), .ZN(n47780) );
  NAND2_X1 U39039 ( .A1(n1331), .A2(n644), .ZN(n1330) );
  NAND2_X1 U39065 ( .A1(n3446), .A2(n51531), .ZN(n31755) );
  NAND2_X1 U39255 ( .A1(n51532), .A2(n31743), .ZN(n51531) );
  INV_X1 U39482 ( .A(n35974), .ZN(n36227) );
  NAND2_X1 U39483 ( .A1(n37592), .A2(n35973), .ZN(n35974) );
  AND2_X1 U39605 ( .A1(n19675), .A2(n51006), .ZN(n19690) );
  NAND3_X1 U39612 ( .A1(n14932), .A2(n3730), .A3(n14933), .ZN(n17887) );
  NAND2_X1 U39722 ( .A1(n31143), .A2(n31142), .ZN(n1551) );
  NAND3_X1 U40167 ( .A1(n1740), .A2(n36526), .A3(n36520), .ZN(n1288) );
  NAND2_X1 U40378 ( .A1(n6490), .A2(n5083), .ZN(n19871) );
  OAI21_X1 U40379 ( .B1(n38404), .B2(n51022), .A(n51622), .ZN(n7779) );
  NAND2_X1 U40392 ( .A1(n11361), .A2(n11376), .ZN(n10695) );
  NAND4_X2 U40568 ( .A1(n10729), .A2(n10730), .A3(n10727), .A4(n10728), .ZN(
        n5176) );
  NAND3_X1 U40615 ( .A1(n31294), .A2(n30642), .A3(n4607), .ZN(n30828) );
  NAND3_X1 U40842 ( .A1(n1942), .A2(n23822), .A3(n24157), .ZN(n20590) );
  NAND2_X1 U40850 ( .A1(n51534), .A2(n5176), .ZN(n14001) );
  NAND3_X1 U40910 ( .A1(n9957), .A2(n9956), .A3(n51535), .ZN(n9958) );
  XNOR2_X2 U40936 ( .A(n17917), .B(n18787), .ZN(n20375) );
  NAND2_X1 U41041 ( .A1(n1367), .A2(n1366), .ZN(n1361) );
  NAND2_X1 U41116 ( .A1(n43474), .A2(n49690), .ZN(n49683) );
  NAND2_X1 U41155 ( .A1(n41728), .A2(n41256), .ZN(n41258) );
  NAND2_X1 U41184 ( .A1(n4796), .A2(n49386), .ZN(n4795) );
  NAND2_X1 U41198 ( .A1(n51536), .A2(n10554), .ZN(n9464) );
  XNOR2_X2 U41200 ( .A(n9452), .B(Key[47]), .ZN(n10554) );
  INV_X1 U41284 ( .A(n9830), .ZN(n51536) );
  XNOR2_X1 U41308 ( .A(n18540), .B(n17900), .ZN(n17904) );
  OAI211_X2 U41402 ( .C1(n13792), .C2(n13793), .A(n13790), .B(n13791), .ZN(
        n18540) );
  NAND2_X1 U41809 ( .A1(n2905), .A2(n12315), .ZN(n9656) );
  XNOR2_X2 U41845 ( .A(Key[121]), .B(Ciphertext[156]), .ZN(n12315) );
  NAND3_X2 U41847 ( .A1(n2310), .A2(n31085), .A3(n51537), .ZN(n36748) );
  XNOR2_X1 U41904 ( .A(n51538), .B(n47388), .ZN(Plaintext[144]) );
  NAND3_X1 U41931 ( .A1(n47386), .A2(n50157), .A3(n47387), .ZN(n51538) );
  OR2_X2 U41996 ( .A1(n51539), .A2(n8658), .ZN(n16532) );
  NAND3_X1 U42013 ( .A1(n14834), .A2(n14830), .A3(n14833), .ZN(n51539) );
  NAND2_X1 U42016 ( .A1(n51129), .A2(n20752), .ZN(n51540) );
  OR2_X1 U42051 ( .A1(n10554), .A2(n9830), .ZN(n9952) );
  INV_X1 U42228 ( .A(n10882), .ZN(n1545) );
  NAND2_X1 U42327 ( .A1(n13514), .A2(n51067), .ZN(n10882) );
  NAND4_X1 U42368 ( .A1(n30259), .A2(n30260), .A3(n30261), .A4(n30262), .ZN(
        n51541) );
  NAND2_X1 U42402 ( .A1(n30266), .A2(n52102), .ZN(n51542) );
  NAND3_X2 U42409 ( .A1(n808), .A2(n3519), .A3(n13428), .ZN(n18668) );
  AOI21_X1 U42431 ( .B1(n49669), .B2(n49672), .A(n49668), .ZN(n49676) );
  NAND3_X1 U42471 ( .A1(n31882), .A2(n31886), .A3(n31792), .ZN(n30127) );
  XNOR2_X1 U42530 ( .A(n51543), .B(n47725), .ZN(Plaintext[18]) );
  NAND3_X1 U42534 ( .A1(n1297), .A2(n1299), .A3(n47724), .ZN(n51543) );
  OR2_X1 U42545 ( .A1(n20157), .A2(n17018), .ZN(n20122) );
  NAND2_X1 U42554 ( .A1(n18010), .A2(n18015), .ZN(n17478) );
  NAND2_X1 U42665 ( .A1(n964), .A2(n39339), .ZN(n51544) );
  XNOR2_X1 U42675 ( .A(n34001), .B(n33334), .ZN(n33340) );
  XNOR2_X1 U42684 ( .A(n34823), .B(n33325), .ZN(n34001) );
  OAI22_X1 U42685 ( .A1(n1568), .A2(n38759), .B1(n41008), .B2(n39614), .ZN(
        n37610) );
  OAI21_X1 U42732 ( .B1(n10993), .B2(n10994), .A(n10992), .ZN(n10995) );
  AND2_X2 U42772 ( .A1(n28723), .A2(n51545), .ZN(n31636) );
  OAI21_X1 U42778 ( .B1(n51547), .B2(n51546), .A(n3096), .ZN(n29091) );
  INV_X1 U42928 ( .A(n29087), .ZN(n51547) );
  NAND2_X1 U43068 ( .A1(n7627), .A2(n31158), .ZN(n31475) );
  NAND2_X1 U43077 ( .A1(n36248), .A2(n37765), .ZN(n37764) );
  XNOR2_X2 U43115 ( .A(n33342), .B(n33341), .ZN(n37765) );
  NAND3_X1 U43279 ( .A1(n9906), .A2(n9907), .A3(n51151), .ZN(n9473) );
  INV_X1 U43373 ( .A(n10706), .ZN(n51550) );
  OR2_X1 U43554 ( .A1(n21820), .A2(n20876), .ZN(n24244) );
  NAND2_X1 U43564 ( .A1(n20193), .A2(n51551), .ZN(n20744) );
  XNOR2_X2 U43601 ( .A(n44353), .B(n43374), .ZN(n42819) );
  NAND3_X2 U43603 ( .A1(n6827), .A2(n39742), .A3(n39743), .ZN(n44353) );
  NAND2_X1 U43604 ( .A1(n46649), .A2(n45771), .ZN(n47123) );
  AND3_X2 U43657 ( .A1(n1859), .A2(n1857), .A3(n1858), .ZN(n22481) );
  NAND2_X1 U43692 ( .A1(n7057), .A2(n48718), .ZN(n87) );
  NAND3_X1 U43817 ( .A1(n13122), .A2(n13124), .A3(n13761), .ZN(n10771) );
  NAND2_X1 U43830 ( .A1(n38644), .A2(n37221), .ZN(n37222) );
  NAND3_X1 U43921 ( .A1(n29724), .A2(n28982), .A3(n28179), .ZN(n3067) );
  AOI22_X1 U43945 ( .A1(n20551), .A2(n20550), .B1(n22476), .B2(n51552), .ZN(
        n7718) );
  NAND2_X1 U44018 ( .A1(n51553), .A2(n51124), .ZN(n51552) );
  INV_X1 U44090 ( .A(n20547), .ZN(n51553) );
  INV_X1 U44125 ( .A(n40749), .ZN(n39891) );
  OR3_X1 U44245 ( .A1(n38237), .A2(n39176), .A3(n51496), .ZN(n38673) );
  OAI211_X1 U44326 ( .C1(n51556), .C2(n11908), .A(n10793), .B(n51554), .ZN(
        n10803) );
  INV_X1 U44427 ( .A(n11063), .ZN(n51556) );
  OAI21_X1 U44514 ( .B1(n30753), .B2(n27557), .A(n1640), .ZN(n51557) );
  NAND2_X1 U44920 ( .A1(n157), .A2(n937), .ZN(n935) );
  NOR2_X1 U45096 ( .A1(n32014), .A2(n32015), .ZN(n32471) );
  NAND2_X1 U45152 ( .A1(n51559), .A2(n51558), .ZN(n16695) );
  NAND2_X1 U45154 ( .A1(n5829), .A2(n23463), .ZN(n51559) );
  XNOR2_X1 U45175 ( .A(n51560), .B(n50173), .ZN(Plaintext[145]) );
  NAND4_X1 U45207 ( .A1(n50172), .A2(n50170), .A3(n50169), .A4(n51570), .ZN(
        n51560) );
  OAI21_X1 U45775 ( .B1(n8510), .B2(n13031), .A(n14264), .ZN(n8511) );
  NAND2_X1 U45841 ( .A1(n15139), .A2(n51142), .ZN(n14264) );
  NAND2_X1 U45896 ( .A1(n2749), .A2(n19534), .ZN(n20118) );
  NAND2_X2 U45897 ( .A1(n6596), .A2(n6597), .ZN(n41085) );
  XNOR2_X1 U45930 ( .A(n27257), .B(n25495), .ZN(n22114) );
  OR2_X2 U45947 ( .A1(n27902), .A2(n6872), .ZN(n32299) );
  NAND3_X1 U46043 ( .A1(n38833), .A2(n38832), .A3(n38831), .ZN(n38835) );
  NAND2_X1 U46204 ( .A1(n52073), .A2(n39751), .ZN(n38831) );
  INV_X1 U46223 ( .A(n27913), .ZN(n27917) );
  INV_X1 U46224 ( .A(n19384), .ZN(n51562) );
  NAND2_X1 U46232 ( .A1(n39272), .A2(n39019), .ZN(n39284) );
  NAND3_X1 U46269 ( .A1(n27639), .A2(n27628), .A3(n27627), .ZN(n26885) );
  NAND3_X1 U46361 ( .A1(n40720), .A2(n41247), .A3(n40719), .ZN(n7889) );
  NAND3_X1 U46567 ( .A1(n50242), .A2(n50240), .A3(n50241), .ZN(n50243) );
  NAND2_X1 U46859 ( .A1(n50223), .A2(n51565), .ZN(n50242) );
  NAND2_X1 U46974 ( .A1(n5602), .A2(n18065), .ZN(n14379) );
  INV_X1 U47038 ( .A(n3645), .ZN(n13153) );
  XNOR2_X1 U47055 ( .A(n51566), .B(n44320), .ZN(n43861) );
  XNOR2_X1 U47058 ( .A(n43846), .B(n44321), .ZN(n51566) );
  NAND2_X1 U47500 ( .A1(n1328), .A2(n44815), .ZN(n44816) );
  NAND2_X1 U47694 ( .A1(n26675), .A2(n27856), .ZN(n51567) );
  NAND2_X1 U47760 ( .A1(n3105), .A2(n2294), .ZN(n51568) );
  NAND3_X1 U47762 ( .A1(n14925), .A2(n15307), .A3(n2189), .ZN(n13789) );
  NOR2_X1 U47770 ( .A1(n15066), .A2(n15309), .ZN(n14925) );
  NAND3_X2 U47771 ( .A1(n38435), .A2(n38434), .A3(n51569), .ZN(n44541) );
  NAND3_X1 U47783 ( .A1(n861), .A2(n37649), .A3(n35731), .ZN(n35740) );
  NAND3_X1 U47785 ( .A1(n10467), .A2(n12630), .A3(n12620), .ZN(n10322) );
  NAND3_X1 U47962 ( .A1(n4570), .A2(n50214), .A3(n50213), .ZN(n51570) );
  NAND2_X1 U48086 ( .A1(n21117), .A2(n22701), .ZN(n21769) );
  OR2_X1 U48293 ( .A1(n51571), .A2(n41034), .ZN(n41294) );
  AOI21_X1 U48299 ( .B1(n40421), .B2(n40417), .A(n5086), .ZN(n51571) );
  NAND2_X1 U48332 ( .A1(n44990), .A2(n41912), .ZN(n45547) );
  NAND2_X1 U48362 ( .A1(n12363), .A2(n10978), .ZN(n7164) );
  OR2_X2 U48617 ( .A1(n51572), .A2(n9651), .ZN(n13849) );
  XNOR2_X2 U48678 ( .A(n51573), .B(n34568), .ZN(n37636) );
  OAI22_X1 U48717 ( .A1(n20122), .A2(n19055), .B1(n5058), .B2(n20116), .ZN(
        n5971) );
  NAND3_X1 U48794 ( .A1(n27683), .A2(n27575), .A3(n27681), .ZN(n26959) );
  NAND2_X1 U48917 ( .A1(n38652), .A2(n51161), .ZN(n38655) );
  NAND3_X1 U48918 ( .A1(n1604), .A2(n35906), .A3(n39781), .ZN(n35913) );
  NOR2_X1 U49023 ( .A1(n14065), .A2(n14394), .ZN(n14403) );
  NAND2_X1 U49024 ( .A1(n14408), .A2(n14412), .ZN(n14065) );
  NAND3_X1 U49078 ( .A1(n27580), .A2(n27581), .A3(n8481), .ZN(n27583) );
  NAND2_X1 U49080 ( .A1(n19966), .A2(n21486), .ZN(n20448) );
  NAND2_X1 U49081 ( .A1(n18032), .A2(n6332), .ZN(n6331) );
  NAND2_X1 U49324 ( .A1(n3459), .A2(n10325), .ZN(n51574) );
  NAND3_X1 U49437 ( .A1(n47535), .A2(n47537), .A3(n47536), .ZN(Plaintext[3])
         );
  NAND2_X1 U49541 ( .A1(n14980), .A2(n780), .ZN(n13677) );
  INV_X1 U49697 ( .A(n13902), .ZN(n129) );
  NAND2_X1 U49796 ( .A1(n15343), .A2(n51575), .ZN(n13902) );
  OAI21_X1 U49950 ( .B1(n51166), .B2(n51576), .A(n47530), .ZN(n47532) );
  NOR2_X1 U50197 ( .A1(n47575), .A2(n52044), .ZN(n51576) );
  NAND2_X1 U50289 ( .A1(n6116), .A2(n43282), .ZN(n43281) );
  XNOR2_X1 U50538 ( .A(n34012), .B(n51578), .ZN(n34056) );
  XNOR2_X1 U50604 ( .A(n8022), .B(n35350), .ZN(n34012) );
  NAND3_X1 U50605 ( .A1(n14998), .A2(n13701), .A3(n15136), .ZN(n51579) );
  OAI21_X1 U50754 ( .B1(n18237), .B2(n18236), .A(n18235), .ZN(n51580) );
  INV_X1 U50907 ( .A(n48927), .ZN(n42805) );
  NAND2_X1 U50908 ( .A1(n52137), .A2(n48975), .ZN(n48927) );
  AOI21_X1 U50909 ( .B1(n21552), .B2(n20643), .A(n20642), .ZN(n20644) );
  NAND2_X1 U50911 ( .A1(n45801), .A2(n46747), .ZN(n44853) );
  NAND2_X1 U50912 ( .A1(n44854), .A2(n44855), .ZN(n44863) );
  NAND2_X1 U50913 ( .A1(n8663), .A2(n14827), .ZN(n15433) );
  NAND2_X1 U50914 ( .A1(n47754), .A2(n47745), .ZN(n47722) );
  NAND2_X1 U50916 ( .A1(n23703), .A2(n51145), .ZN(n51581) );
  NAND2_X1 U50917 ( .A1(n15324), .A2(n15438), .ZN(n7361) );
  XNOR2_X2 U50918 ( .A(n18690), .B(n18126), .ZN(n16431) );
  NAND3_X1 U50920 ( .A1(n22931), .A2(n23044), .A3(n22932), .ZN(n22933) );
  NAND2_X1 U50921 ( .A1(n31116), .A2(n30057), .ZN(n30072) );
  NAND2_X1 U50922 ( .A1(n38159), .A2(n51429), .ZN(n37580) );
  NAND2_X1 U50923 ( .A1(n51582), .A2(n37921), .ZN(n3707) );
  NAND2_X1 U50924 ( .A1(n38663), .A2(n38667), .ZN(n51582) );
  NAND3_X1 U50926 ( .A1(n51583), .A2(n40067), .A3(n39797), .ZN(n39806) );
  NAND2_X1 U50927 ( .A1(n39795), .A2(n39796), .ZN(n51583) );
  NAND3_X1 U50928 ( .A1(n26084), .A2(n28701), .A3(n26650), .ZN(n3740) );
  NAND2_X1 U50929 ( .A1(n51585), .A2(n51584), .ZN(n6907) );
  NAND2_X1 U50930 ( .A1(n9581), .A2(n10422), .ZN(n51585) );
  NAND2_X1 U50932 ( .A1(n2178), .A2(n43688), .ZN(n45164) );
  AND4_X2 U50933 ( .A1(n46991), .A2(n46992), .A3(n46990), .A4(n46993), .ZN(
        n50553) );
  NAND2_X1 U50935 ( .A1(n31625), .A2(n30558), .ZN(n28720) );
  NAND2_X1 U50936 ( .A1(n50693), .A2(n50692), .ZN(n50697) );
  NAND2_X1 U50937 ( .A1(n51587), .A2(n51586), .ZN(n19465) );
  NAND2_X1 U50938 ( .A1(n19463), .A2(n21269), .ZN(n51586) );
  NAND2_X1 U50939 ( .A1(n19462), .A2(n19777), .ZN(n51587) );
  NAND2_X1 U50940 ( .A1(n31537), .A2(n51588), .ZN(n30806) );
  NAND2_X1 U50941 ( .A1(n30967), .A2(n31448), .ZN(n31537) );
  NAND2_X1 U50942 ( .A1(n51589), .A2(n23785), .ZN(n20286) );
  OAI22_X1 U50943 ( .A1(n23454), .A2(n24242), .B1(n20872), .B2(n21823), .ZN(
        n51589) );
  NAND4_X4 U50944 ( .A1(n36500), .A2(n36502), .A3(n36501), .A4(n36499), .ZN(
        n39943) );
  NAND2_X1 U50945 ( .A1(n32298), .A2(n31368), .ZN(n2087) );
  NOR2_X1 U50946 ( .A1(n4299), .A2(n31366), .ZN(n32298) );
  NAND4_X2 U50947 ( .A1(n22432), .A2(n4484), .A3(n22433), .A4(n22431), .ZN(
        n5785) );
  NAND3_X1 U50948 ( .A1(n39340), .A2(n37780), .A3(n39351), .ZN(n39346) );
  NAND2_X1 U50949 ( .A1(n36552), .A2(n7851), .ZN(n5688) );
  NAND2_X1 U50950 ( .A1(n41355), .A2(n40740), .ZN(n41353) );
  OR2_X2 U50951 ( .A1(n4626), .A2(n6148), .ZN(n41355) );
  NOR2_X2 U50952 ( .A1(n21137), .A2(n21136), .ZN(n25050) );
  NAND3_X1 U50953 ( .A1(n6590), .A2(n6593), .A3(n21132), .ZN(n21137) );
  INV_X1 U50954 ( .A(n26882), .ZN(n30997) );
  NAND2_X1 U50955 ( .A1(n31497), .A2(n30102), .ZN(n26882) );
  XNOR2_X1 U50956 ( .A(n25664), .B(n26160), .ZN(n25665) );
  XNOR2_X2 U50959 ( .A(n33541), .B(n34369), .ZN(n35133) );
  NAND2_X2 U50960 ( .A1(n51590), .A2(n1397), .ZN(n34369) );
  NAND3_X1 U50961 ( .A1(n19313), .A2(n6175), .A3(n19312), .ZN(n6174) );
  NAND3_X1 U50962 ( .A1(n4877), .A2(n23752), .A3(n51591), .ZN(n23868) );
  NAND3_X1 U50963 ( .A1(n23191), .A2(n23203), .A3(n2210), .ZN(n51591) );
  NAND4_X2 U50964 ( .A1(n12468), .A2(n12469), .A3(n12466), .A4(n12467), .ZN(
        n14957) );
  NAND2_X1 U50965 ( .A1(n3242), .A2(n33004), .ZN(n33011) );
  NAND3_X1 U50967 ( .A1(n51592), .A2(n28574), .A3(n28934), .ZN(n28575) );
  NAND3_X1 U50968 ( .A1(n28572), .A2(n29020), .A3(n28571), .ZN(n51592) );
  XNOR2_X1 U50969 ( .A(n51593), .B(n35747), .ZN(n35755) );
  XNOR2_X1 U50970 ( .A(n35750), .B(n35746), .ZN(n51593) );
  NAND2_X1 U50971 ( .A1(n9212), .A2(n9211), .ZN(n6037) );
  XNOR2_X1 U50972 ( .A(n51594), .B(n4648), .ZN(n16673) );
  XNOR2_X1 U50973 ( .A(n16591), .B(n17942), .ZN(n51594) );
  NAND2_X1 U50974 ( .A1(n36216), .A2(n39478), .ZN(n34698) );
  NAND2_X1 U50975 ( .A1(n473), .A2(n33870), .ZN(n39478) );
  INV_X1 U50976 ( .A(n51595), .ZN(n3901) );
  OAI211_X1 U50977 ( .C1(n4984), .C2(n51395), .A(n1032), .B(n51596), .ZN(
        n51595) );
  INV_X1 U50978 ( .A(n45022), .ZN(n51596) );
  XNOR2_X1 U50979 ( .A(n50488), .B(n51597), .ZN(Plaintext[155]) );
  NAND3_X1 U50980 ( .A1(n51598), .A2(n8245), .A3(n1311), .ZN(n51597) );
  XNOR2_X1 U50981 ( .A(n51599), .B(n26577), .ZN(n26579) );
  XNOR2_X1 U50982 ( .A(n27418), .B(n26576), .ZN(n51599) );
  NOR2_X1 U50985 ( .A1(n51147), .A2(n51601), .ZN(n40161) );
  OAI21_X1 U50986 ( .B1(n40570), .B2(n40157), .A(n40151), .ZN(n51601) );
  XNOR2_X1 U50987 ( .A(n51602), .B(n45884), .ZN(Plaintext[21]) );
  NAND4_X4 U50989 ( .A1(n31374), .A2(n1083), .A3(n31373), .A4(n31372), .ZN(
        n34219) );
  NAND2_X1 U50990 ( .A1(n3498), .A2(n51603), .ZN(n3497) );
  NAND4_X2 U50995 ( .A1(n51606), .A2(n40217), .A3(n40216), .A4(n41241), .ZN(
        n41518) );
  INV_X1 U50996 ( .A(n40219), .ZN(n51606) );
  NAND2_X1 U50997 ( .A1(n1656), .A2(n23049), .ZN(n23060) );
  NAND2_X1 U50998 ( .A1(n51607), .A2(n32918), .ZN(n32921) );
  NAND2_X1 U50999 ( .A1(n32915), .A2(n51608), .ZN(n51607) );
  NAND2_X1 U51000 ( .A1(n3238), .A2(n32313), .ZN(n31971) );
  XNOR2_X1 U51001 ( .A(n51609), .B(n6327), .ZN(Plaintext[87]) );
  NAND3_X1 U51002 ( .A1(n47486), .A2(n7277), .A3(n3206), .ZN(n51609) );
  NAND3_X2 U51003 ( .A1(n42309), .A2(n42308), .A3(n7067), .ZN(n48935) );
  NAND2_X2 U51004 ( .A1(n38313), .A2(n39289), .ZN(n39300) );
  NAND2_X1 U51005 ( .A1(n10828), .A2(n5268), .ZN(n51610) );
  NAND2_X1 U51006 ( .A1(n12495), .A2(n10827), .ZN(n51612) );
  NAND2_X1 U51007 ( .A1(n45828), .A2(n44646), .ZN(n44826) );
  XNOR2_X1 U51008 ( .A(n51613), .B(n33708), .ZN(n45) );
  XNOR2_X1 U51009 ( .A(n6205), .B(n33706), .ZN(n51613) );
  NAND2_X1 U51010 ( .A1(n30392), .A2(n30391), .ZN(n4216) );
  OR2_X2 U51011 ( .A1(n51614), .A2(n3651), .ZN(n45877) );
  NAND4_X1 U51012 ( .A1(n44833), .A2(n44821), .A3(n44818), .A4(n51637), .ZN(
        n51614) );
  OAI211_X1 U51015 ( .C1(n17623), .C2(n17624), .A(n17622), .B(n4346), .ZN(
        n17632) );
  NAND2_X1 U51016 ( .A1(n32421), .A2(n32830), .ZN(n51616) );
  NAND2_X1 U51017 ( .A1(n51618), .A2(n32823), .ZN(n51617) );
  NAND2_X1 U51019 ( .A1(n40674), .A2(n51619), .ZN(n38408) );
  NAND2_X1 U51021 ( .A1(n12639), .A2(n51621), .ZN(n12641) );
  NAND2_X1 U51022 ( .A1(n39929), .A2(n38402), .ZN(n51622) );
  AND2_X1 U51023 ( .A1(n18863), .A2(n20686), .ZN(n51624) );
  AND3_X1 U51024 ( .A1(n7420), .A2(n6903), .A3(n52210), .ZN(n51625) );
  OR2_X1 U51025 ( .A1(n24334), .A2(n20711), .ZN(n51626) );
  XNOR2_X1 U51026 ( .A(n25739), .B(n26049), .ZN(n51627) );
  OR2_X1 U51027 ( .A1(n32771), .A2(n32175), .ZN(n51628) );
  OR3_X1 U51028 ( .A1(n32175), .A2(n32965), .A3(n32760), .ZN(n51629) );
  AND2_X1 U51029 ( .A1(n32815), .A2(n31401), .ZN(n51630) );
  AND3_X1 U51030 ( .A1(n32526), .A2(n32525), .A3(n32966), .ZN(n51631) );
  XNOR2_X2 U51031 ( .A(n35503), .B(n34533), .ZN(n36869) );
  OR2_X1 U51032 ( .A1(n35566), .A2(n37480), .ZN(n51632) );
  BUF_X1 U51033 ( .A(n35890), .Z(n38341) );
  NAND3_X2 U51034 ( .A1(n35715), .A2(n35716), .A3(n35717), .ZN(n4954) );
  AND3_X1 U51035 ( .A1(n40690), .A2(n40692), .A3(n40675), .ZN(n51633) );
  AND2_X1 U51037 ( .A1(n41714), .A2(n41716), .ZN(n51634) );
  XNOR2_X2 U51038 ( .A(n42683), .B(n42682), .ZN(n45967) );
  BUF_X2 U51039 ( .A(n46880), .Z(n2159) );
  NOR2_X1 U51041 ( .A1(n49956), .A2(n49940), .ZN(n51635) );
  AND4_X1 U51042 ( .A1(n50387), .A2(n50390), .A3(n49742), .A4(n47321), .ZN(
        n51636) );
  AND2_X1 U51043 ( .A1(n112), .A2(n3933), .ZN(n51637) );
  NAND2_X2 U18666 ( .A1(n6674), .A2(n660), .ZN(n48437) );
  INV_X2 U626 ( .A(n40338), .ZN(n40328) );
  BUF_X1 U2214 ( .A(n7558), .Z(n445) );
  AND2_X2 U4977 ( .A1(n11931), .A2(n12705), .ZN(n12696) );
  OR2_X2 U4723 ( .A1(n13753), .A2(n13752), .ZN(n18175) );
  AND2_X2 U1478 ( .A1(n11621), .A2(n11634), .ZN(n11464) );
  BUF_X2 U5075 ( .A(n8775), .Z(n10240) );
  AND2_X2 U3623 ( .A1(n39474), .A2(n37805), .ZN(n39488) );
  BUF_X2 U7590 ( .A(n13945), .Z(n2173) );
  INV_X2 U12686 ( .A(n9074), .ZN(n3250) );
  NAND2_X2 U13755 ( .A1(n27613), .A2(n3502), .ZN(n32473) );
  AND2_X2 U1381 ( .A1(n18726), .A2(n21351), .ZN(n21356) );
  AND2_X2 U31692 ( .A1(n22416), .A2(n23987), .ZN(n23032) );
  AND4_X2 U790 ( .A1(n25401), .A2(n25402), .A3(n25399), .A4(n25400), .ZN(n6969) );
  AND2_X2 U41889 ( .A1(n39235), .A2(n38704), .ZN(n39245) );
  INV_X1 U16475 ( .A(n40446), .ZN(n40403) );
  XNOR2_X2 U1193 ( .A(n37131), .B(n37132), .ZN(n38241) );
  BUF_X1 U2097 ( .A(n28638), .Z(n383) );
  XNOR2_X1 U2431 ( .A(n21681), .B(n24531), .ZN(n27638) );
  OR2_X2 U2693 ( .A1(n24563), .A2(n29467), .ZN(n29461) );
  BUF_X2 U2549 ( .A(n46069), .Z(n51409) );
  OR2_X2 U8431 ( .A1(n23832), .A2(n24158), .ZN(n24146) );
  NAND4_X4 U29271 ( .A1(n18614), .A2(n18613), .A3(n18612), .A4(n18611), .ZN(
        n24187) );
  INV_X2 U15901 ( .A(n41770), .ZN(n42145) );
  NOR2_X2 U6171 ( .A1(n51671), .A2(n14712), .ZN(n14718) );
  AND3_X2 U5967 ( .A1(n307), .A2(n308), .A3(n10088), .ZN(n10899) );
  NAND4_X4 U2405 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n44848), .ZN(n47786) );
  XNOR2_X2 U2790 ( .A(n18454), .B(n18453), .ZN(n20201) );
  OR2_X2 U2781 ( .A1(n3230), .A2(n38598), .ZN(n41332) );
  AND2_X2 U2670 ( .A1(n27794), .A2(n3125), .ZN(n31418) );
  AND2_X2 U16875 ( .A1(n22714), .A2(n22470), .ZN(n22308) );
  XNOR2_X2 U3741 ( .A(n33647), .B(n5809), .ZN(n37560) );
  BUF_X2 U2594 ( .A(n38258), .Z(n2188) );
  OR2_X2 U5515 ( .A1(n661), .A2(n46810), .ZN(n47069) );
  OR2_X2 U1828 ( .A1(n27644), .A2(n27643), .ZN(n32485) );
  INV_X2 U3974 ( .A(n29616), .ZN(n32600) );
  AND3_X2 U4012 ( .A1(n28162), .A2(n7334), .A3(n7333), .ZN(n29616) );
  OR2_X2 U4889 ( .A1(n11530), .A2(n7340), .ZN(n12572) );
  BUF_X2 U2237 ( .A(n24333), .Z(n457) );
  AND2_X2 U744 ( .A1(n6538), .A2(n36141), .ZN(n38549) );
  XNOR2_X2 U44492 ( .A(n41721), .B(n41722), .ZN(n45188) );
  BUF_X1 U1312 ( .A(n16037), .Z(n51018) );
  NAND2_X2 U16628 ( .A1(n8423), .A2(n8425), .ZN(n30853) );
  BUF_X2 U2381 ( .A(n37403), .Z(n525) );
  OR2_X2 U4499 ( .A1(n17081), .A2(n21248), .ZN(n18963) );
  OR2_X2 U1823 ( .A1(n40579), .A2(n40578), .ZN(n41187) );
  OR2_X2 U9139 ( .A1(n5150), .A2(n21355), .ZN(n21360) );
  CLKBUF_X3 U1085 ( .A(n33709), .Z(n2204) );
  BUF_X2 U2160 ( .A(n39181), .Z(n419) );
  OR2_X2 U4193 ( .A1(n25734), .A2(n3059), .ZN(n28688) );
  BUF_X2 U7 ( .A(n47857), .Z(n508) );
  INV_X2 U2664 ( .A(n32874), .ZN(n33041) );
  BUF_X1 U4672 ( .A(n18819), .Z(n2216) );
  OR2_X2 U46 ( .A1(n216), .A2(n33068), .ZN(n40377) );
  INV_X2 U1097 ( .A(n41735), .ZN(n41256) );
  NOR2_X2 U36525 ( .A1(n32851), .A2(n32377), .ZN(n31920) );
  AND2_X2 U4553 ( .A1(n18039), .A2(n8378), .ZN(n19424) );
  OAI21_X2 U4880 ( .B1(n10011), .B2(n10012), .A(n11027), .ZN(n10898) );
  NAND3_X2 U3284 ( .A1(n51160), .A2(n30388), .A3(n30400), .ZN(n32420) );
  BUF_X2 U7481 ( .A(n50772), .Z(n2095) );
  AND2_X2 U12065 ( .A1(n45659), .A2(n46395), .ZN(n46503) );
  BUF_X1 U1790 ( .A(n16126), .Z(n51049) );
  OAI211_X2 U14317 ( .C1(n21438), .C2(n8148), .A(n18608), .B(n18609), .ZN(
        n18614) );
  BUF_X2 U2241 ( .A(n36575), .Z(n458) );
  AND2_X2 U8451 ( .A1(n18563), .A2(n20326), .ZN(n21438) );
  BUF_X2 U6058 ( .A(n8886), .Z(n8882) );
  BUF_X1 U3364 ( .A(n45400), .Z(n2185) );
  CLKBUF_X3 U3330 ( .A(n42271), .Z(n49163) );
  XNOR2_X2 U4287 ( .A(n25240), .B(n28370), .ZN(n24855) );
  OR2_X4 U456 ( .A1(n38646), .A2(n38645), .ZN(n41348) );
  AND4_X2 U1996 ( .A1(n27151), .A2(n27150), .A3(n8580), .A4(n8579), .ZN(n30873) );
  BUF_X1 U4562 ( .A(n15093), .Z(n17489) );
  AND2_X2 U14286 ( .A1(n11015), .A2(n11011), .ZN(n11004) );
  INV_X2 U3799 ( .A(n33397), .ZN(n35534) );
  XNOR2_X2 U14456 ( .A(n4015), .B(Key[191]), .ZN(n9049) );
  OR2_X2 U4601 ( .A1(n16792), .A2(n17057), .ZN(n20097) );
  AND2_X2 U7302 ( .A1(n50951), .A2(n45194), .ZN(n50949) );
  AND2_X2 U118 ( .A1(n8423), .A2(n8425), .ZN(n51545) );
  OR2_X2 U3376 ( .A1(n40699), .A2(n40698), .ZN(n44217) );
  OR2_X2 U1281 ( .A1(n373), .A2(n19869), .ZN(n19865) );
  OR2_X2 U3165 ( .A1(n32251), .A2(n32242), .ZN(n31240) );
  BUF_X1 U349 ( .A(n5454), .Z(n2154) );
  BUF_X2 U2644 ( .A(n717), .Z(n31413) );
  NAND4_X4 U4419 ( .A1(n7994), .A2(n20318), .A3(n20319), .A4(n7995), .ZN(
        n23044) );
  NAND4_X4 U7663 ( .A1(n7095), .A2(n7096), .A3(n19003), .A4(n19004), .ZN(
        n22989) );
  XNOR2_X2 U35097 ( .A(n33702), .B(n33973), .ZN(n51497) );
  NOR2_X2 U10091 ( .A1(n14207), .A2(n14206), .ZN(n17281) );
  INV_X1 U8221 ( .A(n51688), .ZN(n5081) );
  XNOR2_X2 U1080 ( .A(n36792), .B(n33104), .ZN(n34753) );
  NAND2_X2 U12585 ( .A1(n21424), .A2(n20325), .ZN(n21420) );
  OR2_X4 U13537 ( .A1(n38026), .A2(n38025), .ZN(n40903) );
  CLKBUF_X3 U4667 ( .A(n18804), .Z(n2226) );
  AND3_X2 U2619 ( .A1(n39586), .A2(n39588), .A3(n5460), .ZN(n42458) );
  AND2_X2 U3256 ( .A1(n43460), .A2(n43464), .ZN(n49191) );
  BUF_X1 U3010 ( .A(Key[165]), .Z(n4579) );
  INV_X2 U5736 ( .A(n32463), .ZN(n1085) );
  AND2_X2 U29862 ( .A1(n8796), .A2(n8795), .ZN(n9785) );
  INV_X1 U22499 ( .A(n22901), .ZN(n22916) );
  OR2_X2 U747 ( .A1(n29454), .A2(n29453), .ZN(n30930) );
  BUF_X2 U2198 ( .A(n31850), .Z(n435) );
  AND3_X2 U5928 ( .A1(n34200), .A2(n5523), .A3(n5524), .ZN(n5525) );
  NAND4_X2 U31537 ( .A1(n22162), .A2(n22161), .A3(n22160), .A4(n22159), .ZN(
        n24791) );
  AND2_X2 U1575 ( .A1(n30683), .A2(n30687), .ZN(n28757) );
  OR2_X2 U1454 ( .A1(n27987), .A2(n27121), .ZN(n28579) );
  BUF_X2 U7553 ( .A(n30459), .Z(n2143) );
  BUF_X2 U2192 ( .A(n40781), .Z(n431) );
  AND2_X2 U3617 ( .A1(n37806), .A2(n39479), .ZN(n39486) );
  AND2_X2 U9717 ( .A1(n596), .A2(n42061), .ZN(n40293) );
  OR2_X2 U4873 ( .A1(n15279), .A2(n15278), .ZN(n15285) );
  NAND4_X2 U2269 ( .A1(n19766), .A2(n19767), .A3(n19765), .A4(n19764), .ZN(
        n25320) );
  NOR2_X2 U1025 ( .A1(n22701), .A2(n51080), .ZN(n21114) );
  INV_X1 U49008 ( .A(n33221), .ZN(n47708) );
  NAND2_X2 U1392 ( .A1(n6405), .A2(n6410), .ZN(n15278) );
  NAND3_X2 U419 ( .A1(n31348), .A2(n31349), .A3(n8292), .ZN(n37137) );
  NOR2_X2 U520 ( .A1(n14958), .A2(n14962), .ZN(n14059) );
  NAND4_X4 U7623 ( .A1(n27598), .A2(n27596), .A3(n27597), .A4(n27595), .ZN(
        n32478) );
  BUF_X2 U30 ( .A(n45127), .Z(n671) );
  AND2_X2 U1505 ( .A1(n36232), .A2(n37591), .ZN(n37597) );
  XNOR2_X2 U45811 ( .A(n43350), .B(n43349), .ZN(n46095) );
  AND2_X2 U528 ( .A1(n40556), .A2(n40316), .ZN(n40566) );
  NAND2_X2 U7239 ( .A1(n48180), .A2(n48404), .ZN(n48410) );
  OR2_X2 U1414 ( .A1(n614), .A2(n33174), .ZN(n35159) );
  NAND2_X2 U3782 ( .A1(n8483), .A2(n8484), .ZN(n36685) );
  OAI22_X2 U8629 ( .A1(n30715), .A2(n30713), .B1(n27594), .B2(n29855), .ZN(
        n27597) );
  CLKBUF_X3 U2015 ( .A(n36509), .Z(n39751) );
  NAND3_X2 U4238 ( .A1(n21317), .A2(n22068), .A3(n21316), .ZN(n24047) );
  NAND4_X4 U1304 ( .A1(n20263), .A2(n20264), .A3(n20262), .A4(n20265), .ZN(
        n23785) );
  AND2_X2 U15731 ( .A1(n50270), .A2(n51410), .ZN(n50281) );
  XNOR2_X2 U3361 ( .A(n51307), .B(n51100), .ZN(n45269) );
  AND2_X2 U3616 ( .A1(n33174), .A2(n614), .ZN(n36376) );
  NAND4_X2 U36186 ( .A1(n28454), .A2(n28453), .A3(n28452), .A4(n28451), .ZN(
        n32965) );
  AND2_X2 U8299 ( .A1(n12198), .A2(n12204), .ZN(n13587) );
  AND2_X2 U2843 ( .A1(n35310), .A2(n38638), .ZN(n38252) );
  BUF_X2 U3370 ( .A(n42659), .Z(n44296) );
  OR2_X4 U10015 ( .A1(n9019), .A2(n9018), .ZN(n14311) );
  NAND3_X2 U4266 ( .A1(n19319), .A2(n19318), .A3(n2264), .ZN(n26529) );
  AND2_X2 U35569 ( .A1(n487), .A2(n51746), .ZN(n29873) );
  OR2_X2 U19730 ( .A1(n39470), .A2(n39469), .ZN(n41587) );
  BUF_X2 U4625 ( .A(n18610), .Z(n21427) );
  INV_X2 U4872 ( .A(n51712), .ZN(n14515) );
  INV_X1 U1904 ( .A(n18495), .ZN(n21547) );
  BUF_X1 U1787 ( .A(n33981), .Z(n2167) );
  INV_X1 U7331 ( .A(n32254), .ZN(n32243) );
  OR3_X4 U149 ( .A1(n1452), .A2(n1451), .A3(n1453), .ZN(n23832) );
  NAND4_X2 U2520 ( .A1(n44791), .A2(n44790), .A3(n44789), .A4(n45214), .ZN(
        n49070) );
  AND2_X2 U18738 ( .A1(n8260), .A2(n30534), .ZN(n30528) );
  NAND4_X2 U30683 ( .A1(n40077), .A2(n40076), .A3(n40079), .A4(n40078), .ZN(
        n51461) );
  AND2_X2 U8300 ( .A1(n12125), .A2(n9405), .ZN(n11379) );
  AND2_X2 U263 ( .A1(n48778), .A2(n995), .ZN(n48750) );
  OR3_X2 U3362 ( .A1(n6144), .A2(n6145), .A3(n40036), .ZN(n7608) );
  XNOR2_X1 U19212 ( .A(n23780), .B(n23781), .ZN(n30663) );
  BUF_X2 U21883 ( .A(n26567), .Z(n51380) );
  BUF_X1 U3537 ( .A(n26567), .Z(n51120) );
  BUF_X2 U3287 ( .A(n50383), .Z(n2199) );
  AND4_X2 U41811 ( .A1(n37181), .A2(n37180), .A3(n37179), .A4(n37178), .ZN(
        n37186) );
  BUF_X2 U30620 ( .A(n17671), .Z(n51459) );
  BUF_X1 U988 ( .A(n37020), .Z(n50982) );
  BUF_X2 U3279 ( .A(n31567), .Z(n51106) );
  OR2_X2 U3152 ( .A1(n50641), .A2(n51029), .ZN(n50615) );
  BUF_X1 U3757 ( .A(n34911), .Z(n37745) );
  NAND4_X4 U18283 ( .A1(n49196), .A2(n49195), .A3(n49194), .A4(n49193), .ZN(
        n49376) );
  NAND2_X2 U107 ( .A1(n28938), .A2(n4141), .ZN(n31911) );
  NOR2_X2 U46972 ( .A1(n24187), .A2(n24180), .ZN(n4462) );
  AND2_X2 U10982 ( .A1(n45693), .A2(n46358), .ZN(n46346) );
  INV_X2 U2235 ( .A(n41912), .ZN(n48205) );
  AOI21_X1 U1788 ( .B1(n19031), .B2(n19030), .A(n4242), .ZN(n4241) );
  BUF_X2 U206 ( .A(n12205), .Z(n14280) );
  BUF_X1 U39978 ( .A(n34528), .Z(n38282) );
  AND2_X2 U9797 ( .A1(n48722), .A2(n48769), .ZN(n48760) );
  OR3_X2 U3829 ( .A1(n862), .A2(n29377), .A3(n29376), .ZN(n37062) );
  AND4_X1 U4275 ( .A1(n21994), .A2(n21993), .A3(n21985), .A4(n1559), .ZN(n1345) );
  NOR2_X1 U9065 ( .A1(n13947), .A2(n13945), .ZN(n12882) );
  BUF_X2 U1252 ( .A(n8824), .Z(n11027) );
  OR2_X2 U2260 ( .A1(n26973), .A2(n51747), .ZN(n27795) );
  OR2_X2 U41703 ( .A1(n39377), .A2(n39369), .ZN(n39388) );
  NAND4_X4 U11225 ( .A1(n9611), .A2(n9612), .A3(n9613), .A4(n9610), .ZN(n15256) );
  OR2_X2 U5046 ( .A1(n9104), .A2(n9103), .ZN(n11635) );
  BUF_X2 U2079 ( .A(n28301), .Z(n369) );
  AND2_X2 U1552 ( .A1(n20082), .A2(n19141), .ZN(n20063) );
  NAND2_X2 U3168 ( .A1(n50407), .A2(n50406), .ZN(n50486) );
  XNOR2_X2 U12526 ( .A(n18750), .B(n16485), .ZN(n17976) );
  XNOR2_X2 U4195 ( .A(n18602), .B(n18712), .ZN(n16485) );
  OR2_X2 U13 ( .A1(n45988), .A2(n45987), .ZN(n49195) );
  NAND2_X2 U14843 ( .A1(n29290), .A2(n28695), .ZN(n29306) );
  BUF_X1 U2078 ( .A(n28301), .Z(n368) );
  NOR2_X2 U334 ( .A1(n3243), .A2(n51050), .ZN(n18903) );
  BUF_X2 U4106 ( .A(n23861), .Z(n27604) );
  BUF_X1 U3685 ( .A(n31358), .Z(n38226) );
  AND2_X1 U584 ( .A1(n15435), .A2(n15448), .ZN(n15342) );
  BUF_X2 U1260 ( .A(n41149), .Z(n51012) );
  NAND4_X2 U37814 ( .A1(n31213), .A2(n31212), .A3(n31211), .A4(n31210), .ZN(
        n33142) );
  BUF_X1 U2703 ( .A(n27093), .Z(n30200) );
  AND3_X2 U48815 ( .A1(n47423), .A2(n7345), .A3(n47424), .ZN(n49903) );
  BUF_X1 U129 ( .A(n5228), .Z(n459) );
  BUF_X2 U239 ( .A(n13504), .Z(n51066) );
  NAND4_X4 U5556 ( .A1(n1919), .A2(n1918), .A3(n46341), .A4(n46340), .ZN(
        n48751) );
  XNOR2_X1 U13475 ( .A(Key[178]), .B(Ciphertext[123]), .ZN(n10519) );
  XNOR2_X1 U1039 ( .A(Key[166]), .B(Ciphertext[39]), .ZN(n8885) );
  XNOR2_X1 U1291 ( .A(Key[35]), .B(Ciphertext[34]), .ZN(n9547) );
  XNOR2_X1 U21865 ( .A(Key[38]), .B(Ciphertext[103]), .ZN(n11639) );
  XNOR2_X1 U377 ( .A(n9055), .B(Key[46]), .ZN(n9057) );
  XNOR2_X1 U20770 ( .A(n8785), .B(Key[18]), .ZN(n9786) );
  XNOR2_X1 U14795 ( .A(n8986), .B(Key[172]), .ZN(n12266) );
  XNOR2_X1 U4764 ( .A(n1594), .B(Key[130]), .ZN(n9015) );
  XNOR2_X1 U21142 ( .A(n8786), .B(Key[93]), .ZN(n10268) );
  XNOR2_X1 U1600 ( .A(n8867), .B(Key[100]), .ZN(n11900) );
  XNOR2_X2 U26030 ( .A(n4793), .B(n4579), .ZN(n42816) );
  XNOR2_X1 U885 ( .A(n9400), .B(Key[139]), .ZN(n9406) );
  XNOR2_X1 U5061 ( .A(n9332), .B(Key[10]), .ZN(n9339) );
  INV_X1 U1037 ( .A(n8849), .ZN(n10529) );
  INV_X1 U11148 ( .A(n11530), .ZN(n7341) );
  XNOR2_X1 U624 ( .A(n9245), .B(Key[148]), .ZN(n9433) );
  INV_X1 U5022 ( .A(n9140), .ZN(n11704) );
  INV_X1 U21723 ( .A(n9210), .ZN(n12630) );
  INV_X1 U21118 ( .A(n11011), .ZN(n10192) );
  INV_X1 U1338 ( .A(n9336), .ZN(n9341) );
  AND2_X1 U5014 ( .A1(n9510), .A2(n9306), .ZN(n11663) );
  INV_X1 U1127 ( .A(n8773), .ZN(n11015) );
  INV_X1 U21156 ( .A(n8790), .ZN(n9782) );
  NAND2_X1 U268 ( .A1(n10519), .A2(n10031), .ZN(n10633) );
  INV_X1 U4773 ( .A(n12610), .ZN(n51139) );
  BUF_X1 U4835 ( .A(n9001), .Z(n12280) );
  BUF_X1 U687 ( .A(n8803), .Z(n10121) );
  AND2_X1 U220 ( .A1(n8853), .A2(n10109), .ZN(n10513) );
  AND2_X1 U5047 ( .A1(n9278), .A2(n11611), .ZN(n9279) );
  OR2_X1 U1168 ( .A1(n8909), .A2(n12464), .ZN(n11874) );
  NAND2_X1 U1453 ( .A1(n10781), .A2(n11443), .ZN(n12534) );
  NAND2_X1 U2393 ( .A1(n9109), .A2(n11091), .ZN(n12546) );
  AND2_X1 U5029 ( .A1(n10138), .A2(n8839), .ZN(n10926) );
  AND2_X1 U4974 ( .A1(n9855), .A2(n10052), .ZN(n10964) );
  NAND2_X2 U18771 ( .A1(n51138), .A2(n11354), .ZN(n12389) );
  AND2_X1 U5002 ( .A1(n12573), .A2(n9129), .ZN(n12556) );
  NAND2_X1 U454 ( .A1(n9015), .A2(n3444), .ZN(n7823) );
  NOR2_X1 U5003 ( .A1(n8987), .A2(n10742), .ZN(n12243) );
  AND2_X1 U7689 ( .A1(n9341), .A2(n10594), .ZN(n9973) );
  AND2_X1 U9960 ( .A1(n11276), .A2(n11687), .ZN(n11683) );
  AND2_X1 U1717 ( .A1(n10589), .A2(n11276), .ZN(n11669) );
  AND2_X1 U5006 ( .A1(n9939), .A2(n11639), .ZN(n11658) );
  OR2_X1 U472 ( .A1(n2197), .A2(n8639), .ZN(n11031) );
  BUF_X1 U4971 ( .A(n11077), .Z(n12676) );
  AND2_X1 U15444 ( .A1(n51140), .A2(n357), .ZN(n795) );
  NAND2_X1 U7236 ( .A1(n51139), .A2(n11914), .ZN(n9539) );
  OR2_X1 U2854 ( .A1(n51139), .A2(n11914), .ZN(n11137) );
  NAND2_X1 U7860 ( .A1(n51650), .A2(n11695), .ZN(n11210) );
  AND2_X1 U1199 ( .A1(n10250), .A2(n11011), .ZN(n10195) );
  AND2_X1 U4960 ( .A1(n12323), .A2(n12333), .ZN(n12339) );
  AND2_X1 U12722 ( .A1(n8840), .A2(n10148), .ZN(n10134) );
  NAND2_X1 U13150 ( .A1(n9806), .A2(n8840), .ZN(n10218) );
  AND2_X1 U4996 ( .A1(n11077), .A2(n11884), .ZN(n12454) );
  AND2_X1 U9968 ( .A1(n12173), .A2(n11322), .ZN(n9585) );
  AND2_X1 U4976 ( .A1(n12702), .A2(n11931), .ZN(n12435) );
  AND2_X1 U4985 ( .A1(n11229), .A2(n11226), .ZN(n11234) );
  NOR2_X1 U9063 ( .A1(n6672), .A2(n10601), .ZN(n9878) );
  AOI21_X1 U23813 ( .B1(n12673), .B2(n12672), .A(n12675), .ZN(n11882) );
  AND2_X1 U5244 ( .A1(n10277), .A2(n10673), .ZN(n5776) );
  AND2_X1 U4911 ( .A1(n7178), .A2(n10058), .ZN(n9867) );
  AND4_X1 U214 ( .A1(n9873), .A2(n9881), .A3(n9872), .A4(n6119), .ZN(n4285) );
  AND2_X1 U23364 ( .A1(n11260), .A2(n11259), .ZN(n11266) );
  NOR2_X1 U22427 ( .A1(n9854), .A2(n9853), .ZN(n9868) );
  AND4_X1 U2846 ( .A1(n9312), .A2(n9311), .A3(n9310), .A4(n9309), .ZN(n9315)
         );
  NAND3_X1 U811 ( .A1(n5253), .A2(n5255), .A3(n11490), .ZN(n15358) );
  AND4_X1 U4898 ( .A1(n7554), .A2(n11075), .A3(n11074), .A4(n4915), .ZN(n7555)
         );
  NAND4_X1 U17832 ( .A1(n8726), .A2(n11666), .A3(n11664), .A4(n11665), .ZN(
        n13378) );
  NAND3_X1 U6248 ( .A1(n12148), .A2(n12150), .A3(n3674), .ZN(n14552) );
  NAND4_X2 U23236 ( .A1(n11104), .A2(n11103), .A3(n11102), .A4(n11101), .ZN(
        n15189) );
  NAND4_X2 U12689 ( .A1(n9868), .A2(n9866), .A3(n9865), .A4(n9867), .ZN(n13947) );
  AND4_X1 U552 ( .A1(n8382), .A2(n8383), .A3(n9134), .A4(n9133), .ZN(n12750)
         );
  AND3_X1 U7902 ( .A1(n4372), .A2(n10237), .A3(n10236), .ZN(n7390) );
  AND3_X1 U1662 ( .A1(n12078), .A2(n12077), .A3(n12076), .ZN(n12083) );
  INV_X1 U8334 ( .A(n15341), .ZN(n15335) );
  NAND3_X2 U20501 ( .A1(n12083), .A2(n12082), .A3(n12081), .ZN(n14550) );
  INV_X1 U1738 ( .A(n14472), .ZN(n13845) );
  INV_X1 U6425 ( .A(n13410), .ZN(n14344) );
  NAND2_X1 U4854 ( .A1(n7536), .A2(n9196), .ZN(n14880) );
  INV_X1 U2834 ( .A(n14644), .ZN(n3254) );
  OR2_X1 U1344 ( .A1(n9988), .A2(n9987), .ZN(n12787) );
  NAND2_X1 U4841 ( .A1(n14813), .A2(n14812), .ZN(n15386) );
  BUF_X1 U4598 ( .A(n13131), .Z(n51136) );
  INV_X1 U375 ( .A(n9721), .ZN(n14473) );
  INV_X1 U4864 ( .A(n14345), .ZN(n14331) );
  AND3_X1 U4870 ( .A1(n9736), .A2(n5963), .A3(n5962), .ZN(n14228) );
  OR2_X1 U4817 ( .A1(n13667), .A2(n12755), .ZN(n14635) );
  NAND2_X1 U4431 ( .A1(n3552), .A2(n12893), .ZN(n14660) );
  INV_X1 U17706 ( .A(n13968), .ZN(n13970) );
  INV_X1 U540 ( .A(n13667), .ZN(n14642) );
  INV_X1 U4832 ( .A(n51682), .ZN(n13505) );
  AND2_X1 U1684 ( .A1(n11694), .A2(n11693), .ZN(n6192) );
  AND2_X1 U13667 ( .A1(n3254), .A2(n2114), .ZN(n12757) );
  NOR2_X1 U17688 ( .A1(n15335), .A2(n15440), .ZN(n15337) );
  INV_X1 U2109 ( .A(n15132), .ZN(n15136) );
  INV_X1 U11335 ( .A(n14370), .ZN(n14544) );
  INV_X1 U22210 ( .A(n15256), .ZN(n15263) );
  INV_X1 U897 ( .A(n14533), .ZN(n14553) );
  NAND2_X1 U1180 ( .A1(n154), .A2(n11086), .ZN(n14767) );
  AND2_X1 U5386 ( .A1(n13277), .A2(n15189), .ZN(n14761) );
  AND2_X1 U1822 ( .A1(n13949), .A2(n13930), .ZN(n13934) );
  OR2_X1 U1758 ( .A1(n2970), .A2(n7151), .ZN(n14870) );
  INV_X1 U4886 ( .A(n11558), .ZN(n787) );
  OR2_X2 U4408 ( .A1(n10327), .A2(n51574), .ZN(n15034) );
  AND2_X1 U19065 ( .A1(n7054), .A2(n7053), .ZN(n12205) );
  INV_X1 U4844 ( .A(n13504), .ZN(n13501) );
  NOR2_X1 U478 ( .A1(n13782), .A2(n13161), .ZN(n10904) );
  NOR2_X1 U1099 ( .A1(n3678), .A2(n51136), .ZN(n12903) );
  NOR2_X1 U14876 ( .A1(n3679), .A2(n14186), .ZN(n13139) );
  NOR2_X1 U4806 ( .A1(n12963), .A2(n14412), .ZN(n14400) );
  OR2_X1 U23134 ( .A1(n13166), .A2(n12017), .ZN(n13778) );
  NOR2_X1 U10243 ( .A1(n2151), .A2(n14950), .ZN(n15275) );
  OR4_X1 U656 ( .A1(n13202), .A2(n13201), .A3(n13207), .A4(n13934), .ZN(n13205) );
  NAND4_X1 U15571 ( .A1(n12999), .A2(n12998), .A3(n12997), .A4(n12996), .ZN(
        n15649) );
  NAND3_X1 U6402 ( .A1(n4011), .A2(n12240), .A3(n7927), .ZN(n18547) );
  AND4_X1 U4712 ( .A1(n12225), .A2(n7442), .A3(n14351), .A4(n12226), .ZN(
        n13816) );
  NAND4_X1 U13306 ( .A1(n12970), .A2(n14406), .A3(n12971), .A4(n12969), .ZN(
        n16980) );
  AND3_X1 U5168 ( .A1(n12432), .A2(n12434), .A3(n12433), .ZN(n4170) );
  NAND4_X1 U24019 ( .A1(n12221), .A2(n12220), .A3(n12219), .A4(n12218), .ZN(
        n17793) );
  NAND4_X1 U2199 ( .A1(n11818), .A2(n11815), .A3(n11816), .A4(n11817), .ZN(
        n16662) );
  OR2_X2 U13568 ( .A1(n7884), .A2(n7885), .ZN(n17364) );
  OR2_X1 U921 ( .A1(n12887), .A2(n1302), .ZN(n15956) );
  OR2_X1 U861 ( .A1(n14275), .A2(n14274), .ZN(n18747) );
  NAND2_X1 U4674 ( .A1(n6279), .A2(n10909), .ZN(n18712) );
  NAND3_X1 U428 ( .A1(n51277), .A2(n14131), .A3(n51143), .ZN(n17280) );
  NAND4_X1 U12685 ( .A1(n12919), .A2(n12918), .A3(n12920), .A4(n13099), .ZN(
        n16105) );
  NAND2_X1 U4698 ( .A1(n12980), .A2(n2953), .ZN(n17218) );
  AND4_X1 U24689 ( .A1(n13391), .A2(n13390), .A3(n16035), .A4(n13389), .ZN(
        n13394) );
  NAND2_X1 U12642 ( .A1(n2972), .A2(n11868), .ZN(n17954) );
  NAND2_X1 U465 ( .A1(n1338), .A2(n10092), .ZN(n18643) );
  AND2_X1 U5295 ( .A1(n12839), .A2(n12838), .ZN(n14619) );
  NOR3_X1 U5701 ( .A1(n4196), .A2(n1066), .A3(n3462), .ZN(n4195) );
  NAND3_X1 U757 ( .A1(n1845), .A2(n4520), .A3(n11171), .ZN(n17972) );
  XNOR2_X1 U26561 ( .A(n17925), .B(n16016), .ZN(n18446) );
  NAND4_X1 U15011 ( .A1(n16054), .A2(n16053), .A3(n51763), .A4(n16051), .ZN(
        n18790) );
  INV_X1 U25713 ( .A(n18756), .ZN(n18153) );
  XNOR2_X1 U12016 ( .A(n19248), .B(n2690), .ZN(n16372) );
  BUF_X1 U1777 ( .A(n19213), .Z(n51047) );
  BUF_X2 U2441 ( .A(n18692), .Z(n566) );
  NAND2_X1 U846 ( .A1(n4195), .A2(n13534), .ZN(n17764) );
  CLKBUF_X1 U2010 ( .A(n17212), .Z(n51373) );
  XNOR2_X1 U4670 ( .A(n18669), .B(n18399), .ZN(n16412) );
  BUF_X1 U24591 ( .A(n16624), .Z(n18408) );
  BUF_X1 U1272 ( .A(n17178), .Z(n51014) );
  BUF_X1 U7636 ( .A(n2217), .Z(n2218) );
  XNOR2_X1 U2340 ( .A(n16161), .B(n16160), .ZN(n20062) );
  XNOR2_X1 U2383 ( .A(n16444), .B(n16443), .ZN(n19534) );
  XNOR2_X1 U12368 ( .A(n3766), .B(n8731), .ZN(n16490) );
  XNOR2_X1 U2209 ( .A(n280), .B(n8715), .ZN(n20641) );
  XNOR2_X1 U4651 ( .A(n15817), .B(n15816), .ZN(n20658) );
  BUF_X2 U5561 ( .A(n17526), .Z(n590) );
  XNOR2_X1 U18786 ( .A(n8175), .B(n16517), .ZN(n18063) );
  INV_X2 U27092 ( .A(n16214), .ZN(n20082) );
  XNOR2_X1 U2782 ( .A(n14625), .B(n8728), .ZN(n20393) );
  XNOR2_X1 U4158 ( .A(n17270), .B(n17271), .ZN(n19452) );
  BUF_X2 U1192 ( .A(n51521), .Z(n51006) );
  INV_X1 U26612 ( .A(n20266), .ZN(n21660) );
  BUF_X1 U1620 ( .A(n16546), .Z(n16807) );
  BUF_X1 U750 ( .A(n16395), .Z(n16821) );
  XNOR2_X1 U1871 ( .A(n5956), .B(n6989), .ZN(n1715) );
  OR2_X1 U11438 ( .A1(n18377), .A2(n16820), .ZN(n6515) );
  AND2_X1 U1419 ( .A1(n21186), .A2(n21181), .ZN(n19837) );
  AND2_X1 U793 ( .A1(n17569), .A2(n18009), .ZN(n18012) );
  INV_X1 U4587 ( .A(n17195), .ZN(n21173) );
  BUF_X1 U173 ( .A(n19016), .Z(n19023) );
  AND2_X1 U16168 ( .A1(n21579), .A2(n21578), .ZN(n21407) );
  AND2_X1 U4600 ( .A1(n19344), .A2(n18085), .ZN(n20513) );
  INV_X2 U2474 ( .A(n16678), .ZN(n770) );
  OR2_X1 U248 ( .A1(n1417), .A2(n20147), .ZN(n20144) );
  AND2_X1 U29167 ( .A1(n18495), .A2(n20642), .ZN(n21533) );
  INV_X1 U2773 ( .A(n20375), .ZN(n1860) );
  NAND2_X1 U16105 ( .A1(n20393), .A2(n20383), .ZN(n20473) );
  AND2_X1 U1783 ( .A1(n51385), .A2(n374), .ZN(n19853) );
  AND2_X1 U1324 ( .A1(n19678), .A2(n19679), .ZN(n19681) );
  NAND2_X1 U5750 ( .A1(n16821), .A2(n20029), .ZN(n20027) );
  NAND2_X1 U1661 ( .A1(n7431), .A2(n21530), .ZN(n21525) );
  AND2_X1 U4570 ( .A1(n19675), .A2(n19685), .ZN(n20221) );
  AND2_X1 U4508 ( .A1(n21601), .A2(n21351), .ZN(n21349) );
  OR2_X1 U4514 ( .A1(n21663), .A2(n21664), .ZN(n21648) );
  INV_X1 U18079 ( .A(n20026), .ZN(n18287) );
  OR2_X1 U2761 ( .A1(n20230), .A2(n51090), .ZN(n20670) );
  NAND2_X2 U12673 ( .A1(n770), .A2(n21233), .ZN(n19520) );
  OR2_X1 U6809 ( .A1(n1715), .A2(n772), .ZN(n18064) );
  NAND2_X1 U7731 ( .A1(n21480), .A2(n21495), .ZN(n4174) );
  AND2_X1 U20603 ( .A1(n21173), .A2(n19834), .ZN(n19702) );
  NOR2_X1 U406 ( .A1(n8624), .A2(n20095), .ZN(n20093) );
  NOR2_X1 U26731 ( .A1(n20231), .A2(n20677), .ZN(n20688) );
  INV_X1 U7962 ( .A(n20737), .ZN(n21548) );
  INV_X1 U4513 ( .A(n20670), .ZN(n20679) );
  NOR2_X1 U10188 ( .A1(n19955), .A2(n19943), .ZN(n21430) );
  NAND2_X1 U448 ( .A1(n3222), .A2(n16986), .ZN(n19870) );
  AND2_X1 U378 ( .A1(n19870), .A2(n19871), .ZN(n19650) );
  AND2_X1 U2759 ( .A1(n18051), .A2(n20362), .ZN(n19181) );
  AND3_X1 U7755 ( .A1(n16845), .A2(n19386), .A3(n8486), .ZN(n8485) );
  OR2_X1 U4465 ( .A1(n19467), .A2(n19466), .ZN(n19468) );
  AND4_X1 U12490 ( .A1(n19457), .A2(n2931), .A3(n19456), .A4(n19458), .ZN(
        n19471) );
  AND2_X1 U30294 ( .A1(n20127), .A2(n20126), .ZN(n20164) );
  NAND4_X1 U16183 ( .A1(n15731), .A2(n15732), .A3(n15730), .A4(n15729), .ZN(
        n23825) );
  AND2_X1 U30286 ( .A1(n20113), .A2(n20112), .ZN(n20165) );
  OR2_X2 U3758 ( .A1(n18925), .A2(n18924), .ZN(n23316) );
  INV_X1 U2756 ( .A(n23825), .ZN(n24158) );
  AND2_X1 U1682 ( .A1(n8079), .A2(n4505), .ZN(n8078) );
  AND3_X1 U4445 ( .A1(n1536), .A2(n1533), .A3(n1535), .ZN(n1243) );
  AND2_X1 U1330 ( .A1(n18226), .A2(n18225), .ZN(n22823) );
  AND4_X1 U4462 ( .A1(n5970), .A2(n5973), .A3(n5972), .A4(n5974), .ZN(n17022)
         );
  NAND3_X1 U2051 ( .A1(n8309), .A2(n3089), .A3(n3085), .ZN(n353) );
  NAND4_X2 U45931 ( .A1(n19471), .A2(n19468), .A3(n19470), .A4(n19469), .ZN(
        n23436) );
  NAND2_X1 U1581 ( .A1(n20280), .A2(n6745), .ZN(n21810) );
  AND2_X1 U4392 ( .A1(n21499), .A2(n6206), .ZN(n23135) );
  BUF_X1 U7626 ( .A(n23755), .Z(n2210) );
  CLKBUF_X1 U2145 ( .A(n23208), .Z(n412) );
  INV_X2 U161 ( .A(n22186), .ZN(n21700) );
  OR2_X1 U4447 ( .A1(n17316), .A2(n17315), .ZN(n17417) );
  OR2_X2 U20091 ( .A1(n20965), .A2(n20966), .ZN(n51355) );
  BUF_X2 U29662 ( .A(n19149), .Z(n23238) );
  INV_X1 U157 ( .A(n23149), .ZN(n23153) );
  BUF_X1 U2172 ( .A(n22946), .Z(n424) );
  BUF_X1 U3784 ( .A(n23149), .Z(n51123) );
  OR3_X2 U18076 ( .A1(n6166), .A2(n6164), .A3(n21522), .ZN(n24105) );
  OR2_X2 U8491 ( .A1(n8555), .A2(n4973), .ZN(n23833) );
  OR2_X1 U512 ( .A1(n23414), .A2(n23412), .ZN(n22034) );
  CLKBUF_X2 U148 ( .A(n23177), .Z(n51021) );
  INV_X1 U17645 ( .A(n23473), .ZN(n23467) );
  AND2_X1 U20408 ( .A1(n8416), .A2(n23149), .ZN(n23472) );
  OR2_X1 U10296 ( .A1(n23924), .A2(n22521), .ZN(n5143) );
  OR2_X1 U5987 ( .A1(n8695), .A2(n51660), .ZN(n22149) );
  NOR2_X1 U455 ( .A1(n354), .A2(n5203), .ZN(n24028) );
  OR2_X1 U706 ( .A1(n16688), .A2(n6010), .ZN(n21946) );
  NOR2_X1 U4378 ( .A1(n23955), .A2(n559), .ZN(n23953) );
  AND2_X1 U3731 ( .A1(n21987), .A2(n23479), .ZN(n21983) );
  NOR2_X1 U12365 ( .A1(n22876), .A2(n22769), .ZN(n22874) );
  AND2_X1 U962 ( .A1(n3062), .A2(n23336), .ZN(n22257) );
  OR2_X1 U29880 ( .A1(n24157), .A2(n23821), .ZN(n23276) );
  AND2_X1 U1244 ( .A1(n19625), .A2(n8518), .ZN(n5025) );
  AND2_X1 U4320 ( .A1(n21341), .A2(n20999), .ZN(n8522) );
  INV_X1 U10329 ( .A(n23276), .ZN(n23835) );
  AND2_X1 U1143 ( .A1(n23274), .A2(n23275), .ZN(n23281) );
  AND4_X1 U302 ( .A1(n20724), .A2(n20725), .A3(n20723), .A4(n20722), .ZN(
        n20735) );
  NAND4_X1 U17899 ( .A1(n6690), .A2(n23491), .A3(n6693), .A4(n2258), .ZN(
        n26448) );
  OAI211_X1 U2457 ( .C1(n24249), .C2(n23459), .A(n23458), .B(n23457), .ZN(
        n26531) );
  AND4_X1 U386 ( .A1(n4453), .A2(n20992), .A3(n20999), .A4(n4452), .ZN(n4922)
         );
  AND3_X1 U3643 ( .A1(n51242), .A2(n21056), .A3(n21057), .ZN(n3442) );
  AND4_X1 U4297 ( .A1(n4696), .A2(n6381), .A3(n23918), .A4(n23928), .ZN(n6380)
         );
  NAND4_X1 U15617 ( .A1(n22760), .A2(n22759), .A3(n22758), .A4(n22757), .ZN(
        n26402) );
  AND2_X1 U20480 ( .A1(n8521), .A2(n8520), .ZN(n8519) );
  NAND4_X1 U17876 ( .A1(n23429), .A2(n23432), .A3(n23430), .A4(n23431), .ZN(
        n24548) );
  AND4_X1 U4308 ( .A1(n22112), .A2(n7492), .A3(n22111), .A4(n7491), .ZN(n7493)
         );
  NAND4_X1 U31607 ( .A1(n22270), .A2(n23609), .A3(n22271), .A4(n23602), .ZN(
        n28359) );
  NAND3_X1 U15561 ( .A1(n4765), .A2(n4766), .A3(n22336), .ZN(n25365) );
  NAND4_X1 U145 ( .A1(n146), .A2(n23328), .A3(n22259), .A4(n22265), .ZN(n24616) );
  NAND2_X1 U1462 ( .A1(n3346), .A2(n1279), .ZN(n25927) );
  NAND4_X1 U14740 ( .A1(n22582), .A2(n22581), .A3(n22580), .A4(n22579), .ZN(
        n26600) );
  OR2_X1 U4289 ( .A1(n19440), .A2(n19439), .ZN(n25540) );
  NAND4_X1 U16342 ( .A1(n22694), .A2(n22692), .A3(n22693), .A4(n22691), .ZN(
        n27450) );
  NAND4_X1 U16159 ( .A1(n20008), .A2(n20007), .A3(n20009), .A4(n20006), .ZN(
        n26509) );
  NAND4_X1 U1650 ( .A1(n22680), .A2(n2481), .A3(n22679), .A4(n3820), .ZN(
        n25740) );
  NAND4_X1 U31623 ( .A1(n22305), .A2(n22304), .A3(n22303), .A4(n22302), .ZN(
        n25703) );
  XNOR2_X1 U32727 ( .A(n27250), .B(n42291), .ZN(n25360) );
  NAND3_X1 U4270 ( .A1(n2622), .A2(n22792), .A3(n2621), .ZN(n25445) );
  XNOR2_X1 U1103 ( .A(n27374), .B(n27373), .ZN(n25726) );
  NAND4_X1 U1019 ( .A1(n903), .A2(n20735), .A3(n20733), .A4(n20734), .ZN(n2667) );
  BUF_X1 U802 ( .A(n27393), .Z(n2164) );
  XNOR2_X1 U2148 ( .A(n22727), .B(n25229), .ZN(n28398) );
  NAND2_X1 U4269 ( .A1(n20530), .A2(n20529), .ZN(n28104) );
  BUF_X1 U4273 ( .A(n27393), .Z(n751) );
  NOR2_X1 U4255 ( .A1(n20288), .A2(n20287), .ZN(n26092) );
  XNOR2_X1 U8516 ( .A(n26395), .B(n26044), .ZN(n25590) );
  XNOR2_X1 U2185 ( .A(n26175), .B(n25703), .ZN(n25610) );
  CLKBUF_X1 U1226 ( .A(n28358), .Z(n51009) );
  XNOR2_X1 U7630 ( .A(n24344), .B(n28291), .ZN(n26536) );
  BUF_X2 U3521 ( .A(n25131), .Z(n51119) );
  BUF_X1 U37449 ( .A(n5713), .Z(n51523) );
  XNOR2_X1 U9330 ( .A(n25494), .B(n25493), .ZN(n28223) );
  BUF_X1 U31760 ( .A(n25762), .Z(n27256) );
  BUF_X1 U1590 ( .A(n28312), .Z(n2209) );
  BUF_X1 U1880 ( .A(n28040), .Z(n51056) );
  XNOR2_X1 U33432 ( .A(n24908), .B(n26304), .ZN(n28041) );
  XNOR2_X1 U33024 ( .A(n28250), .B(n24511), .ZN(n24512) );
  XNOR2_X1 U16807 ( .A(n24722), .B(n22695), .ZN(n27183) );
  XNOR2_X1 U1855 ( .A(n7075), .B(n28438), .ZN(n25639) );
  XNOR2_X1 U15579 ( .A(n25552), .B(n25551), .ZN(n29247) );
  XNOR2_X1 U4201 ( .A(n27195), .B(n27194), .ZN(n28971) );
  XNOR2_X1 U1386 ( .A(n25713), .B(n25714), .ZN(n27847) );
  XNOR2_X1 U6769 ( .A(n23461), .B(n23462), .ZN(n30780) );
  XNOR2_X1 U438 ( .A(n7295), .B(n51627), .ZN(n2956) );
  XNOR2_X1 U4204 ( .A(n26001), .B(n26000), .ZN(n26039) );
  INV_X1 U10524 ( .A(n24649), .ZN(n26905) );
  INV_X1 U19143 ( .A(n29443), .ZN(n26068) );
  BUF_X1 U1991 ( .A(n28764), .Z(n29882) );
  INV_X1 U4216 ( .A(n23109), .ZN(n30706) );
  BUF_X1 U133 ( .A(n29443), .Z(n2213) );
  OR2_X1 U4128 ( .A1(n28333), .A2(n28738), .ZN(n29703) );
  BUF_X1 U774 ( .A(n30180), .Z(n2201) );
  BUF_X1 U4214 ( .A(n25603), .Z(n29123) );
  INV_X2 U618 ( .A(n29260), .ZN(n30234) );
  XNOR2_X1 U1483 ( .A(n26383), .B(n26384), .ZN(n28916) );
  XNOR2_X1 U1640 ( .A(n7898), .B(n1270), .ZN(n2707) );
  AND2_X1 U1994 ( .A1(n28708), .A2(n27783), .ZN(n28710) );
  AND2_X1 U33862 ( .A1(n29343), .A2(n30209), .ZN(n27886) );
  AND2_X1 U2686 ( .A1(n29443), .A2(n29447), .ZN(n27835) );
  CLKBUF_X1 U2190 ( .A(n29442), .Z(n430) );
  BUF_X1 U2702 ( .A(n28449), .Z(n29736) );
  INV_X1 U1114 ( .A(n28298), .ZN(n5389) );
  AND2_X1 U4191 ( .A1(n25410), .A2(n52144), .ZN(n30268) );
  INV_X1 U3339 ( .A(n24265), .ZN(n30754) );
  AND2_X1 U1924 ( .A1(n25410), .A2(n25107), .ZN(n30269) );
  INV_X1 U9342 ( .A(n29853), .ZN(n30711) );
  NAND2_X2 U33796 ( .A1(n28578), .A2(n51118), .ZN(n27991) );
  AND2_X1 U132 ( .A1(n51112), .A2(n29413), .ZN(n27706) );
  BUF_X2 U2176 ( .A(n30442), .Z(n427) );
  OR2_X1 U2690 ( .A1(n738), .A2(n24265), .ZN(n30757) );
  AND2_X1 U658 ( .A1(n30754), .A2(n738), .ZN(n30773) );
  BUF_X2 U130 ( .A(n25840), .Z(n28666) );
  OR2_X1 U4174 ( .A1(n26077), .A2(n26083), .ZN(n27844) );
  OR2_X1 U1135 ( .A1(n2677), .A2(n27652), .ZN(n24776) );
  BUF_X2 U2684 ( .A(n28177), .Z(n30419) );
  OR2_X1 U657 ( .A1(n28874), .A2(n29029), .ZN(n29027) );
  NAND2_X2 U4120 ( .A1(n5563), .A2(n25107), .ZN(n2158) );
  AND2_X1 U1329 ( .A1(n28497), .A2(n28965), .ZN(n29796) );
  OR2_X1 U4112 ( .A1(n30179), .A2(n30182), .ZN(n30168) );
  OR2_X1 U4085 ( .A1(n29532), .A2(n28622), .ZN(n28618) );
  AND2_X1 U2342 ( .A1(n30285), .A2(n26494), .ZN(n28545) );
  NAND2_X1 U33384 ( .A1(n28148), .A2(n30296), .ZN(n30291) );
  AND2_X1 U2678 ( .A1(n29418), .A2(n27711), .ZN(n29428) );
  OR2_X1 U10486 ( .A1(n2815), .A2(n30163), .ZN(n28022) );
  INV_X1 U2337 ( .A(n30376), .ZN(n1121) );
  OR2_X1 U6777 ( .A1(n748), .A2(n2677), .ZN(n27665) );
  AND2_X1 U9386 ( .A1(n30723), .A2(n30719), .ZN(n30715) );
  OR2_X1 U8612 ( .A1(n24882), .A2(n28147), .ZN(n28557) );
  NOR2_X1 U1669 ( .A1(n24882), .A2(n30282), .ZN(n28563) );
  AND2_X1 U3305 ( .A1(n28138), .A2(n28497), .ZN(n28865) );
  AND2_X1 U120 ( .A1(n28867), .A2(n3827), .ZN(n28866) );
  BUF_X1 U33688 ( .A(n30159), .Z(n30306) );
  NOR2_X1 U1240 ( .A1(n27097), .A2(n51109), .ZN(n30203) );
  NOR2_X1 U4083 ( .A1(n27097), .A2(n30202), .ZN(n27881) );
  OR2_X1 U4048 ( .A1(n26723), .A2(n27034), .ZN(n29450) );
  OR2_X1 U20924 ( .A1(n27859), .A2(n27858), .ZN(n28672) );
  OR2_X1 U11663 ( .A1(n737), .A2(n27623), .ZN(n27629) );
  AOI22_X1 U15026 ( .A1(n25630), .A2(n25629), .B1(n28664), .B2(n29264), .ZN(
        n25848) );
  OR2_X1 U3988 ( .A1(n26813), .A2(n27577), .ZN(n26961) );
  OAI21_X1 U4032 ( .B1(n29067), .B2(n29770), .A(n29769), .ZN(n28818) );
  AND4_X1 U16132 ( .A1(n30276), .A2(n51541), .A3(n30275), .A4(n51542), .ZN(
        n7064) );
  AND4_X1 U1046 ( .A1(n5472), .A2(n28299), .A3(n5471), .A4(n30342), .ZN(n5470)
         );
  AND4_X1 U3965 ( .A1(n27843), .A2(n1180), .A3(n27842), .A4(n1546), .ZN(n1548)
         );
  AND3_X1 U4014 ( .A1(n27574), .A2(n29895), .A3(n23655), .ZN(n7006) );
  NAND3_X1 U14179 ( .A1(n6524), .A2(n3869), .A3(n3867), .ZN(n32590) );
  AND4_X1 U792 ( .A1(n27817), .A2(n27816), .A3(n27815), .A4(n27814), .ZN(
        n27825) );
  NAND3_X1 U4033 ( .A1(n24780), .A2(n24779), .A3(n6866), .ZN(n31300) );
  AND3_X1 U33208 ( .A1(n24682), .A2(n26853), .A3(n24681), .ZN(n24690) );
  INV_X1 U423 ( .A(n31075), .ZN(n30484) );
  AND4_X1 U7265 ( .A1(n30704), .A2(n30701), .A3(n30702), .A4(n30703), .ZN(
        n31544) );
  OR3_X2 U342 ( .A1(n1977), .A2(n22347), .A3(n1978), .ZN(n32254) );
  NAND3_X1 U1542 ( .A1(n26845), .A2(n26847), .A3(n26846), .ZN(n31489) );
  INV_X1 U4005 ( .A(n32560), .ZN(n32089) );
  AND4_X2 U6301 ( .A1(n29913), .A2(n29914), .A3(n29912), .A4(n29911), .ZN(
        n32056) );
  BUF_X1 U1741 ( .A(n26711), .Z(n30846) );
  OR2_X2 U3968 ( .A1(n3914), .A2(n29307), .ZN(n32107) );
  NOR2_X1 U37606 ( .A1(n32254), .A2(n31778), .ZN(n32231) );
  CLKBUF_X2 U2301 ( .A(n26202), .Z(n32130) );
  NAND2_X1 U1860 ( .A1(n6057), .A2(n1154), .ZN(n32125) );
  OR2_X1 U99 ( .A1(n32719), .A2(n32724), .ZN(n32457) );
  INV_X1 U3993 ( .A(n31418), .ZN(n725) );
  INV_X1 U591 ( .A(n32960), .ZN(n8390) );
  AND3_X1 U440 ( .A1(n25846), .A2(n2442), .A3(n25845), .ZN(n28487) );
  NOR2_X1 U3952 ( .A1(n30924), .A2(n31512), .ZN(n30935) );
  OR2_X1 U35227 ( .A1(n31346), .A2(n29602), .ZN(n29959) );
  INV_X1 U2658 ( .A(n32957), .ZN(n32771) );
  OR2_X1 U5735 ( .A1(n32716), .A2(n1085), .ZN(n32315) );
  NOR2_X1 U2643 ( .A1(n26795), .A2(n30983), .ZN(n2098) );
  OR2_X1 U9436 ( .A1(n32883), .A2(n7231), .ZN(n33032) );
  AND2_X1 U1811 ( .A1(n31749), .A2(n31740), .ZN(n32302) );
  INV_X2 U3950 ( .A(n32595), .ZN(n712) );
  OR2_X1 U3890 ( .A1(n30853), .A2(n1672), .ZN(n31639) );
  NOR2_X1 U3870 ( .A1(n32829), .A2(n32815), .ZN(n32424) );
  AND2_X2 U541 ( .A1(n26849), .A2(n26848), .ZN(n31497) );
  OR2_X1 U37515 ( .A1(n4434), .A2(n31749), .ZN(n32297) );
  NOR2_X1 U36676 ( .A1(n32407), .A2(n32066), .ZN(n32081) );
  BUF_X1 U2224 ( .A(n31307), .Z(n51086) );
  NAND2_X1 U3161 ( .A1(n7430), .A2(n32407), .ZN(n32409) );
  AND2_X1 U970 ( .A1(n8542), .A2(n32420), .ZN(n32825) );
  OR2_X1 U7803 ( .A1(n27075), .A2(n31340), .ZN(n31935) );
  INV_X1 U11237 ( .A(n30593), .ZN(n31087) );
  NAND2_X1 U3145 ( .A1(n32080), .A2(n32401), .ZN(n33151) );
  AND4_X1 U549 ( .A1(n30088), .A2(n30089), .A3(n30090), .A4(n30087), .ZN(
        n30096) );
  NOR2_X1 U9509 ( .A1(n7066), .A2(n31932), .ZN(n27078) );
  OR3_X1 U28375 ( .A1(n32305), .A2(n32300), .A3(n2334), .ZN(n31757) );
  AND4_X1 U2349 ( .A1(n31604), .A2(n8635), .A3(n31605), .A4(n8634), .ZN(n8633)
         );
  NAND4_X2 U37063 ( .A1(n29834), .A2(n29835), .A3(n29836), .A4(n32568), .ZN(
        n36999) );
  NAND4_X1 U2130 ( .A1(n32061), .A2(n32058), .A3(n32059), .A4(n32060), .ZN(
        n36722) );
  NOR2_X1 U2440 ( .A1(n31909), .A2(n31908), .ZN(n36703) );
  AND3_X1 U1165 ( .A1(n30616), .A2(n151), .A3(n150), .ZN(n149) );
  AND2_X1 U1743 ( .A1(n2843), .A2(n6322), .ZN(n32997) );
  AND3_X1 U1556 ( .A1(n32668), .A2(n6785), .A3(n4573), .ZN(n33943) );
  BUF_X1 U3809 ( .A(n32952), .Z(n35633) );
  XNOR2_X1 U3820 ( .A(n35762), .B(n37318), .ZN(n36873) );
  NAND2_X1 U2320 ( .A1(n5044), .A2(n31806), .ZN(n7199) );
  NAND2_X1 U935 ( .A1(n4684), .A2(n4685), .ZN(n33894) );
  NAND3_X1 U15283 ( .A1(n4319), .A2(n32221), .A3(n4318), .ZN(n33848) );
  NAND2_X1 U2639 ( .A1(n3139), .A2(n29092), .ZN(n35522) );
  XNOR2_X1 U39892 ( .A(n34360), .B(n4847), .ZN(n35669) );
  XNOR2_X1 U17928 ( .A(n37261), .B(n33336), .ZN(n34491) );
  INV_X1 U2636 ( .A(n33894), .ZN(n35501) );
  BUF_X2 U78 ( .A(n33703), .Z(n35625) );
  XNOR2_X1 U2629 ( .A(n7611), .B(n35086), .ZN(n37284) );
  XNOR2_X1 U6465 ( .A(n34811), .B(n34812), .ZN(n34392) );
  BUF_X1 U999 ( .A(n37020), .Z(n50983) );
  XNOR2_X1 U1840 ( .A(n35064), .B(n35063), .ZN(n38464) );
  XNOR2_X1 U1391 ( .A(n36716), .B(n36715), .ZN(n39007) );
  XNOR2_X1 U625 ( .A(n36990), .B(n36989), .ZN(n37790) );
  XNOR2_X1 U2319 ( .A(n34358), .B(n7732), .ZN(n36458) );
  BUF_X1 U1277 ( .A(n36429), .Z(n51015) );
  XNOR2_X1 U2018 ( .A(n36834), .B(n2277), .ZN(n38953) );
  XNOR2_X1 U3103 ( .A(n33239), .B(n33238), .ZN(n34958) );
  XNOR2_X1 U2626 ( .A(n5531), .B(n33209), .ZN(n34189) );
  XNOR2_X1 U2346 ( .A(n35044), .B(n35043), .ZN(n35103) );
  BUF_X1 U2616 ( .A(n35693), .Z(n38585) );
  XNOR2_X1 U3755 ( .A(n34584), .B(n32275), .ZN(n34971) );
  AND2_X1 U22820 ( .A1(n34629), .A2(n37633), .ZN(n35728) );
  AND2_X1 U5170 ( .A1(n39195), .A2(n38957), .ZN(n39194) );
  AND2_X1 U243 ( .A1(n7083), .A2(n37765), .ZN(n37749) );
  OR2_X1 U1863 ( .A1(n38057), .A2(n5464), .ZN(n38054) );
  INV_X1 U670 ( .A(n36015), .ZN(n63) );
  BUF_X1 U10684 ( .A(n35666), .Z(n36133) );
  XNOR2_X1 U2255 ( .A(n33518), .B(n35551), .ZN(n37385) );
  BUF_X1 U2479 ( .A(n38575), .Z(n591) );
  AND2_X1 U3737 ( .A1(n37406), .A2(n33650), .ZN(n37553) );
  XNOR2_X1 U105 ( .A(n8611), .B(n31966), .ZN(n35010) );
  AND2_X1 U3708 ( .A1(n34528), .A2(n34529), .ZN(n38284) );
  NOR2_X1 U3736 ( .A1(n34656), .A2(n36428), .ZN(n36616) );
  XNOR2_X1 U3080 ( .A(n37312), .B(n37313), .ZN(n51508) );
  NOR2_X1 U3712 ( .A1(n36428), .A2(n8089), .ZN(n36426) );
  NAND2_X1 U345 ( .A1(n3248), .A2(n34987), .ZN(n37990) );
  OR2_X1 U23526 ( .A1(n37596), .A2(n37378), .ZN(n36225) );
  AND2_X1 U3681 ( .A1(n7483), .A2(n37633), .ZN(n37637) );
  NAND2_X1 U6969 ( .A1(n8480), .A2(n39273), .ZN(n39271) );
  BUF_X2 U767 ( .A(n33871), .Z(n39472) );
  OR2_X1 U297 ( .A1(n37488), .A2(n8315), .ZN(n37430) );
  OR2_X1 U1504 ( .A1(n39429), .A2(n5151), .ZN(n39422) );
  AND2_X1 U2602 ( .A1(n38941), .A2(n38950), .ZN(n39204) );
  AND2_X1 U3627 ( .A1(n38027), .A2(n614), .ZN(n34948) );
  XNOR2_X1 U2132 ( .A(n35759), .B(n35758), .ZN(n38728) );
  AND2_X1 U692 ( .A1(n37750), .A2(n37745), .ZN(n37766) );
  NAND2_X1 U6841 ( .A1(n36372), .A2(n38040), .ZN(n38031) );
  NAND2_X1 U15272 ( .A1(n38273), .A2(n38271), .ZN(n38283) );
  OR2_X1 U1739 ( .A1(n38005), .A2(n36359), .ZN(n37997) );
  OR2_X1 U3717 ( .A1(n7004), .A2(n37385), .ZN(n38493) );
  AND2_X1 U11581 ( .A1(n37385), .A2(n7004), .ZN(n35953) );
  OR2_X1 U2254 ( .A1(n37385), .A2(n37519), .ZN(n35951) );
  OR2_X1 U1574 ( .A1(n3927), .A2(n36454), .ZN(n35214) );
  OR2_X2 U8679 ( .A1(n52191), .A2(n8509), .ZN(n36115) );
  INV_X1 U15162 ( .A(n35102), .ZN(n38477) );
  AND2_X1 U39040 ( .A1(n37756), .A2(n37496), .ZN(n36247) );
  AND2_X1 U2848 ( .A1(n38543), .A2(n36141), .ZN(n38212) );
  BUF_X1 U337 ( .A(n38273), .Z(n37629) );
  OR2_X1 U3720 ( .A1(n616), .A2(n38728), .ZN(n37654) );
  BUF_X1 U68 ( .A(n33994), .Z(n37985) );
  NAND2_X1 U338 ( .A1(n33994), .A2(n37976), .ZN(n37975) );
  AND2_X1 U1528 ( .A1(n39262), .A2(n39268), .ZN(n39285) );
  AND2_X1 U1544 ( .A1(n39262), .A2(n39007), .ZN(n39264) );
  NAND2_X2 U1938 ( .A1(n36468), .A2(n37665), .ZN(n38337) );
  AND2_X1 U1518 ( .A1(n3255), .A2(n38340), .ZN(n2714) );
  AND2_X1 U11796 ( .A1(n2188), .A2(n38638), .ZN(n38629) );
  INV_X1 U11668 ( .A(n37810), .ZN(n39471) );
  OR2_X1 U2590 ( .A1(n689), .A2(n38572), .ZN(n36103) );
  NOR2_X1 U41452 ( .A1(n36588), .A2(n36587), .ZN(n36601) );
  AND4_X1 U40984 ( .A1(n35865), .A2(n35864), .A3(n35863), .A4(n35862), .ZN(
        n35870) );
  AND4_X1 U39950 ( .A1(n34431), .A2(n36600), .A3(n36580), .A4(n34430), .ZN(
        n34432) );
  AND4_X1 U3568 ( .A1(n35697), .A2(n35696), .A3(n35699), .A4(n37582), .ZN(
        n5031) );
  NAND4_X2 U42450 ( .A1(n38269), .A2(n38266), .A3(n38268), .A4(n38267), .ZN(
        n40868) );
  AND4_X1 U3572 ( .A1(n34983), .A2(n34982), .A3(n34981), .A4(n34980), .ZN(
        n34991) );
  AND3_X1 U43099 ( .A1(n39346), .A2(n39345), .A3(n39344), .ZN(n39356) );
  AND4_X1 U1803 ( .A1(n37795), .A2(n37794), .A3(n37796), .A4(n37797), .ZN(
        n8332) );
  OR2_X1 U1503 ( .A1(n33681), .A2(n33682), .ZN(n43666) );
  NAND4_X1 U3535 ( .A1(n36154), .A2(n36153), .A3(n36152), .A4(n36151), .ZN(
        n40029) );
  AND3_X1 U8797 ( .A1(n37540), .A2(n37564), .A3(n37541), .ZN(n8539) );
  NAND2_X1 U791 ( .A1(n1191), .A2(n2441), .ZN(n39712) );
  OR2_X2 U1833 ( .A1(n35463), .A2(n35462), .ZN(n40558) );
  AND2_X1 U609 ( .A1(n35302), .A2(n35301), .ZN(n35429) );
  AND3_X1 U40805 ( .A1(n35585), .A2(n35584), .A3(n35583), .ZN(n40572) );
  NAND3_X1 U457 ( .A1(n7224), .A2(n6540), .A3(n7223), .ZN(n41446) );
  BUF_X1 U2488 ( .A(n41489), .Z(n596) );
  INV_X2 U43160 ( .A(n40029), .ZN(n41202) );
  OR3_X2 U2142 ( .A1(n36204), .A2(n42055), .A3(n42056), .ZN(n40295) );
  AND4_X1 U3517 ( .A1(n34954), .A2(n34956), .A3(n34957), .A4(n34955), .ZN(
        n40500) );
  INV_X1 U3554 ( .A(n41211), .ZN(n685) );
  INV_X1 U3491 ( .A(n41207), .ZN(n41210) );
  BUF_X2 U42100 ( .A(n39077), .Z(n40815) );
  INV_X1 U17874 ( .A(n41442), .ZN(n41433) );
  NOR2_X1 U12290 ( .A1(n37342), .A2(n4064), .ZN(n2855) );
  OR2_X2 U12803 ( .A1(n7349), .A2(n2492), .ZN(n42205) );
  AND2_X1 U3461 ( .A1(n4302), .A2(n40558), .ZN(n40573) );
  BUF_X1 U2584 ( .A(n38812), .Z(n43665) );
  INV_X1 U15868 ( .A(n39857), .ZN(n40341) );
  AND4_X2 U13748 ( .A1(n37899), .A2(n37898), .A3(n37896), .A4(n37897), .ZN(
        n40943) );
  BUF_X2 U1838 ( .A(n41208), .Z(n51052) );
  INV_X1 U314 ( .A(n38812), .ZN(n41800) );
  NAND2_X1 U14631 ( .A1(n4070), .A2(n4367), .ZN(n40125) );
  NAND4_X1 U41158 ( .A1(n36091), .A2(n36090), .A3(n36089), .A4(n36088), .ZN(
        n38782) );
  INV_X1 U3494 ( .A(n39899), .ZN(n37356) );
  AND3_X1 U10795 ( .A1(n3775), .A2(n40960), .A3(n41374), .ZN(n40957) );
  OR2_X1 U14138 ( .A1(n39409), .A2(n5048), .ZN(n41581) );
  INV_X2 U3509 ( .A(n38764), .ZN(n43329) );
  AND2_X1 U3496 ( .A1(n39543), .A2(n40250), .ZN(n3514) );
  OR2_X1 U11844 ( .A1(n41671), .A2(n41685), .ZN(n40210) );
  INV_X1 U2574 ( .A(n40330), .ZN(n7117) );
  OR2_X1 U8166 ( .A1(n575), .A2(n39955), .ZN(n39111) );
  OR2_X1 U1144 ( .A1(n41356), .A2(n41348), .ZN(n41358) );
  INV_X1 U35186 ( .A(n40081), .ZN(n40906) );
  BUF_X2 U2193 ( .A(n40781), .Z(n432) );
  AND2_X1 U3475 ( .A1(n41702), .A2(n41693), .ZN(n41163) );
  OR2_X1 U3484 ( .A1(n40558), .A2(n3043), .ZN(n40549) );
  AND2_X1 U7324 ( .A1(n42201), .A2(n41938), .ZN(n41932) );
  OR2_X1 U1545 ( .A1(n6468), .A2(n41348), .ZN(n39632) );
  AND2_X1 U1208 ( .A1(n41751), .A2(n687), .ZN(n42144) );
  NOR2_X1 U315 ( .A1(n43329), .A2(n43327), .ZN(n38763) );
  NOR2_X1 U6923 ( .A1(n432), .A2(n40774), .ZN(n40600) );
  OR2_X1 U1479 ( .A1(n42441), .A2(n679), .ZN(n42048) );
  NOR2_X1 U474 ( .A1(n3597), .A2(n40730), .ZN(n41900) );
  OR2_X1 U12669 ( .A1(n7702), .A2(n7701), .ZN(n36395) );
  AND4_X1 U1668 ( .A1(n41335), .A2(n41321), .A3(n41334), .A4(n41322), .ZN(n859) );
  NAND3_X1 U3411 ( .A1(n6508), .A2(n39698), .A3(n2064), .ZN(n45097) );
  AND3_X1 U3417 ( .A1(n37708), .A2(n37713), .A3(n37707), .ZN(n3417) );
  NAND2_X1 U281 ( .A1(n6503), .A2(n40994), .ZN(n43584) );
  NAND4_X1 U316 ( .A1(n40103), .A2(n40102), .A3(n40101), .A4(n40100), .ZN(
        n42316) );
  NAND4_X1 U51036 ( .A1(n40323), .A2(n40321), .A3(n40322), .A4(n40324), .ZN(
        n44182) );
  NAND4_X1 U3391 ( .A1(n39328), .A2(n39327), .A3(n40696), .A4(n39326), .ZN(
        n45467) );
  NAND4_X1 U1725 ( .A1(n40406), .A2(n1403), .A3(n40407), .A4(n1381), .ZN(
        n43357) );
  AND3_X1 U1416 ( .A1(n41044), .A2(n41042), .A3(n41295), .ZN(n5017) );
  NAND3_X1 U895 ( .A1(n7461), .A2(n4280), .A3(n40129), .ZN(n42500) );
  NAND4_X1 U2348 ( .A1(n40629), .A2(n40628), .A3(n40627), .A4(n40626), .ZN(
        n44327) );
  NAND4_X1 U2618 ( .A1(n41423), .A2(n41422), .A3(n41421), .A4(n7039), .ZN(
        n51294) );
  NAND4_X2 U622 ( .A1(n39717), .A2(n39715), .A3(n314), .A4(n1183), .ZN(n44944)
         );
  NAND2_X1 U18554 ( .A1(n6595), .A2(n8337), .ZN(n45445) );
  XNOR2_X1 U2066 ( .A(n44240), .B(n44314), .ZN(n1673) );
  NAND4_X1 U3368 ( .A1(n39137), .A2(n39136), .A3(n39135), .A4(n39134), .ZN(
        n43723) );
  NAND3_X1 U33 ( .A1(n1723), .A2(n39333), .A3(n39332), .ZN(n44374) );
  NAND3_X1 U16629 ( .A1(n42023), .A2(n42024), .A3(n42022), .ZN(n45408) );
  BUF_X1 U2641 ( .A(n45400), .Z(n51099) );
  NAND4_X1 U2266 ( .A1(n40435), .A2(n40434), .A3(n40432), .A4(n40433), .ZN(
        n6345) );
  XNOR2_X1 U6178 ( .A(n52096), .B(n41308), .ZN(n44525) );
  XNOR2_X1 U3371 ( .A(n43619), .B(n44237), .ZN(n45274) );
  BUF_X1 U19163 ( .A(n43833), .Z(n51333) );
  XNOR2_X1 U1191 ( .A(n40757), .B(n42863), .ZN(n45252) );
  BUF_X1 U34949 ( .A(n44081), .Z(n51494) );
  BUF_X2 U51040 ( .A(n43180), .Z(n49980) );
  BUF_X1 U1601 ( .A(n41908), .Z(n44990) );
  BUF_X1 U3309 ( .A(n42605), .Z(n46353) );
  CLKBUF_X2 U2082 ( .A(n39811), .Z(n48433) );
  BUF_X1 U24 ( .A(n50374), .Z(n51058) );
  INV_X1 U47381 ( .A(n46463), .ZN(n48239) );
  AND2_X1 U20571 ( .A1(n44673), .A2(n48479), .ZN(n913) );
  BUF_X2 U1979 ( .A(n40174), .Z(n48436) );
  NAND2_X1 U293 ( .A1(n667), .A2(n6811), .ZN(n50363) );
  CLKBUF_X1 U2510 ( .A(n46691), .Z(n51399) );
  NAND2_X1 U237 ( .A1(n49731), .A2(n423), .ZN(n50378) );
  BUF_X1 U44754 ( .A(n42180), .Z(n45827) );
  BUF_X2 U1184 ( .A(n42305), .Z(n49162) );
  BUF_X1 U2555 ( .A(n45771), .Z(n46842) );
  AND2_X1 U2313 ( .A1(n47152), .A2(n46888), .ZN(n47150) );
  INV_X1 U27 ( .A(n44118), .ZN(n50277) );
  OR2_X1 U18614 ( .A1(n51526), .A2(n7616), .ZN(n50322) );
  BUF_X1 U1579 ( .A(n45922), .Z(n587) );
  BUF_X2 U23 ( .A(n45922), .Z(n588) );
  AND2_X1 U14530 ( .A1(n48462), .A2(n48461), .ZN(n46441) );
  AND2_X1 U13535 ( .A1(n669), .A2(n46872), .ZN(n47104) );
  OR2_X1 U46526 ( .A1(n46475), .A2(n52066), .ZN(n48498) );
  BUF_X1 U2471 ( .A(n47078), .Z(n400) );
  OR2_X1 U17013 ( .A1(n51094), .A2(n42990), .ZN(n49717) );
  AND2_X1 U20276 ( .A1(n46627), .A2(n44873), .ZN(n45761) );
  OR2_X1 U3227 ( .A1(n48546), .A2(n45628), .ZN(n48550) );
  AND2_X1 U3236 ( .A1(n45589), .A2(n44431), .ZN(n48438) );
  BUF_X1 U1439 ( .A(n43795), .Z(n50366) );
  OR2_X1 U1614 ( .A1(n4274), .A2(n44873), .ZN(n46632) );
  AND2_X1 U16104 ( .A1(n44996), .A2(n48213), .ZN(n48210) );
  AND2_X1 U19639 ( .A1(n50315), .A2(n52143), .ZN(n50329) );
  AND2_X1 U1561 ( .A1(n48206), .A2(n44992), .ZN(n45539) );
  OR2_X1 U45246 ( .A1(n49201), .A2(n49197), .ZN(n46231) );
  AND2_X1 U12464 ( .A1(n46903), .A2(n46691), .ZN(n46919) );
  AND2_X1 U3254 ( .A1(n45551), .A2(n44992), .ZN(n45545) );
  OR2_X1 U3250 ( .A1(n46475), .A2(n52039), .ZN(n48521) );
  OR2_X1 U2487 ( .A1(n46201), .A2(n46203), .ZN(n49267) );
  NAND2_X1 U16115 ( .A1(n42703), .A2(n44752), .ZN(n49209) );
  AND2_X1 U3220 ( .A1(n44765), .A2(n46358), .ZN(n46355) );
  OR2_X1 U45210 ( .A1(n46352), .A2(n42602), .ZN(n45232) );
  CLKBUF_X1 U1885 ( .A(n44765), .Z(n46345) );
  AND2_X1 U320 ( .A1(n46905), .A2(n46693), .ZN(n46912) );
  AND2_X1 U44651 ( .A1(n52161), .A2(n44693), .ZN(n48214) );
  AND3_X1 U3188 ( .A1(n47912), .A2(n47913), .A3(n47914), .ZN(n44655) );
  NOR2_X1 U8846 ( .A1(n6536), .A2(n539), .ZN(n46258) );
  AND3_X1 U1524 ( .A1(n46482), .A2(n46481), .A3(n46480), .ZN(n48697) );
  NAND3_X1 U12389 ( .A1(n42803), .A2(n42802), .A3(n2898), .ZN(n48957) );
  INV_X1 U2519 ( .A(n47403), .ZN(n48698) );
  MUX2_X1 U26462 ( .A(n46516), .B(n46515), .S(n48416), .Z(n46527) );
  AND2_X1 U273 ( .A1(n44112), .A2(n5742), .ZN(n50641) );
  NAND3_X1 U49465 ( .A1(n48495), .A2(n48496), .A3(n48494), .ZN(n48647) );
  OAI21_X1 U1087 ( .B1(n49221), .B2(n49220), .A(n131), .ZN(n6685) );
  NOR2_X1 U7622 ( .A1(n48697), .A2(n48714), .ZN(n48685) );
  AND3_X1 U46655 ( .A1(n44416), .A2(n44415), .A3(n44414), .ZN(n48083) );
  NAND4_X1 U32346 ( .A1(n6029), .A2(n42406), .A3(n6030), .A4(n6028), .ZN(
        n51478) );
  OAI211_X1 U20122 ( .C1(n49986), .C2(n47360), .A(n49991), .B(n8114), .ZN(
        n50127) );
  OR2_X1 U3115 ( .A1(n48659), .A2(n48703), .ZN(n48687) );
  BUF_X1 U2023 ( .A(n48365), .Z(n51072) );
  INV_X1 U644 ( .A(n50716), .ZN(n50680) );
  NOR2_X1 U815 ( .A1(n3075), .A2(n48077), .ZN(n48059) );
  AND2_X1 U48533 ( .A1(n50521), .A2(n50520), .ZN(n50526) );
  NOR2_X2 U48586 ( .A1(n50809), .A2(n50773), .ZN(n50804) );
  CLKBUF_X1 U392 ( .A(n48730), .Z(n48768) );
  BUF_X2 U2400 ( .A(n45859), .Z(n47665) );
  OR2_X1 U11046 ( .A1(n47683), .A2(n47667), .ZN(n5966) );
  BUF_X1 U2997 ( .A(Key[114]), .Z(n3383) );
  BUF_X1 U2890 ( .A(Key[188]), .Z(n47401) );
  BUF_X2 U2906 ( .A(Key[167]), .Z(n4694) );
  BUF_X2 U2911 ( .A(Key[60]), .Z(n4931) );
  CLKBUF_X1 U2952 ( .A(Key[34]), .Z(n4317) );
  INV_X1 U21404 ( .A(n8949), .ZN(n9109) );
  INV_X2 U21849 ( .A(n9289), .ZN(n10074) );
  INV_X2 U373 ( .A(n51652), .ZN(n12514) );
  INV_X1 U2862 ( .A(n10831), .ZN(n5180) );
  BUF_X1 U5034 ( .A(n9045), .Z(n12333) );
  INV_X1 U2867 ( .A(n10302), .ZN(n12313) );
  NAND2_X2 U735 ( .A1(n10525), .A2(n10529), .ZN(n10508) );
  INV_X1 U1890 ( .A(n12301), .ZN(n12317) );
  INV_X2 U5017 ( .A(n12659), .ZN(n12649) );
  INV_X2 U21693 ( .A(n11978), .ZN(n9188) );
  INV_X2 U2861 ( .A(n12285), .ZN(n12291) );
  INV_X2 U21312 ( .A(n12728), .ZN(n11964) );
  INV_X2 U2870 ( .A(n12373), .ZN(n12380) );
  INV_X2 U5023 ( .A(n10161), .ZN(n8639) );
  INV_X2 U21208 ( .A(n10162), .ZN(n10584) );
  NAND2_X2 U2853 ( .A1(n11359), .A2(n10375), .ZN(n12107) );
  BUF_X1 U409 ( .A(n9429), .Z(n12129) );
  NAND2_X2 U2857 ( .A1(n11275), .A2(n9969), .ZN(n11279) );
  NAND2_X2 U6035 ( .A1(n9419), .A2(n11341), .ZN(n11346) );
  NAND2_X2 U4969 ( .A1(n51762), .A2(n9744), .ZN(n11008) );
  INV_X2 U4879 ( .A(n1571), .ZN(n13207) );
  INV_X1 U1897 ( .A(n13091), .ZN(n13103) );
  INV_X1 U4851 ( .A(n13633), .ZN(n785) );
  INV_X1 U1998 ( .A(n12834), .ZN(n783) );
  INV_X2 U4868 ( .A(n12750), .ZN(n13669) );
  INV_X1 U7899 ( .A(n13086), .ZN(n13090) );
  INV_X2 U2831 ( .A(n14070), .ZN(n14408) );
  INV_X2 U2818 ( .A(n14011), .ZN(n13316) );
  INV_X2 U4878 ( .A(n14601), .ZN(n14170) );
  INV_X2 U2841 ( .A(n13102), .ZN(n13092) );
  INV_X2 U2388 ( .A(n13173), .ZN(n13161) );
  INV_X2 U6389 ( .A(n15309), .ZN(n15300) );
  INV_X1 U208 ( .A(n13801), .ZN(n277) );
  INV_X2 U18169 ( .A(n13820), .ZN(n14307) );
  INV_X2 U10359 ( .A(n14155), .ZN(n14150) );
  INV_X2 U2822 ( .A(n14318), .ZN(n14320) );
  NAND2_X1 U2813 ( .A1(n14228), .A2(n14224), .ZN(n13960) );
  INV_X2 U2819 ( .A(n15046), .ZN(n15044) );
  INV_X2 U4830 ( .A(n13761), .ZN(n14966) );
  INV_X1 U22697 ( .A(n14160), .ZN(n14156) );
  NAND2_X1 U13965 ( .A1(n14550), .A2(n14545), .ZN(n14368) );
  INV_X1 U1755 ( .A(n14870), .ZN(n15421) );
  CLKBUF_X2 U4774 ( .A(n2149), .Z(n2150) );
  NAND2_X2 U4396 ( .A1(n13061), .A2(n14137), .ZN(n15257) );
  INV_X1 U20083 ( .A(n14984), .ZN(n15103) );
  NAND3_X2 U1831 ( .A1(n14837), .A2(n14836), .A3(n15758), .ZN(n16701) );
  INV_X2 U2287 ( .A(n15014), .ZN(n18119) );
  BUF_X1 U7633 ( .A(n17913), .Z(n2215) );
  INV_X2 U2783 ( .A(n20493), .ZN(n21465) );
  INV_X1 U11214 ( .A(n21198), .ZN(n6078) );
  INV_X1 U1072 ( .A(n20641), .ZN(n6929) );
  INV_X1 U1903 ( .A(n19504), .ZN(n19503) );
  INV_X1 U16701 ( .A(n19112), .ZN(n6226) );
  INV_X1 U2792 ( .A(n18942), .ZN(n19894) );
  INV_X1 U7668 ( .A(n18063), .ZN(n17553) );
  INV_X1 U26657 ( .A(n15872), .ZN(n20677) );
  INV_X1 U2384 ( .A(n20684), .ZN(n51090) );
  NOR2_X1 U5783 ( .A1(n21484), .A2(n19969), .ZN(n21492) );
  INV_X1 U2785 ( .A(n19969), .ZN(n21495) );
  INV_X2 U26821 ( .A(n15997), .ZN(n21614) );
  INV_X2 U2227 ( .A(n19535), .ZN(n20158) );
  NAND2_X1 U6665 ( .A1(n6226), .A2(n19510), .ZN(n21234) );
  NAND2_X1 U4538 ( .A1(n19007), .A2(n19725), .ZN(n19819) );
  NOR2_X2 U2765 ( .A1(n771), .A2(n18376), .ZN(n20046) );
  NAND2_X1 U2775 ( .A1(n19016), .A2(n2182), .ZN(n19785) );
  NAND2_X2 U13637 ( .A1(n52210), .A2(n21530), .ZN(n21521) );
  OAI21_X1 U18853 ( .B1(n19465), .B2(n51013), .A(n6868), .ZN(n19469) );
  INV_X2 U653 ( .A(n23546), .ZN(n23563) );
  INV_X1 U10279 ( .A(n21885), .ZN(n21887) );
  INV_X1 U3798 ( .A(n22470), .ZN(n51124) );
  INV_X2 U2750 ( .A(n21947), .ZN(n23157) );
  OR2_X1 U4372 ( .A1(n24191), .A2(n24187), .ZN(n23871) );
  NAND2_X2 U29046 ( .A1(n21725), .A2(n23229), .ZN(n23213) );
  INV_X1 U4424 ( .A(n23961), .ZN(n754) );
  INV_X2 U5802 ( .A(n23981), .ZN(n23987) );
  BUF_X1 U2743 ( .A(n19901), .Z(n23092) );
  INV_X2 U6921 ( .A(n23785), .ZN(n24238) );
  INV_X1 U2749 ( .A(n23489), .ZN(n23485) );
  INV_X1 U5845 ( .A(n22390), .ZN(n753) );
  INV_X2 U676 ( .A(n23178), .ZN(n23184) );
  INV_X2 U2746 ( .A(n20298), .ZN(n22826) );
  INV_X2 U4390 ( .A(n22481), .ZN(n22714) );
  INV_X1 U5276 ( .A(n20876), .ZN(n24245) );
  INV_X2 U13680 ( .A(n24332), .ZN(n23703) );
  INV_X2 U2354 ( .A(n23833), .ZN(n24150) );
  INV_X2 U14128 ( .A(n23374), .ZN(n5415) );
  INV_X1 U30582 ( .A(n22736), .ZN(n23811) );
  INV_X1 U9310 ( .A(n25365), .ZN(n27473) );
  INV_X1 U4222 ( .A(n27652), .ZN(n748) );
  INV_X1 U2718 ( .A(n26668), .ZN(n27852) );
  INV_X1 U8023 ( .A(n6730), .ZN(n29155) );
  XNOR2_X1 U1292 ( .A(n25167), .B(n25166), .ZN(n30171) );
  INV_X1 U14928 ( .A(n28923), .ZN(n29011) );
  INV_X1 U19671 ( .A(n2956), .ZN(n27858) );
  NAND2_X1 U13560 ( .A1(n51490), .A2(n29764), .ZN(n30349) );
  INV_X1 U699 ( .A(n30191), .ZN(n30202) );
  NAND2_X2 U3337 ( .A1(n29325), .A2(n52217), .ZN(n29332) );
  NAND2_X2 U964 ( .A1(n8455), .A2(n29545), .ZN(n27697) );
  BUF_X1 U2681 ( .A(n24878), .Z(n30295) );
  NAND2_X2 U15077 ( .A1(n6080), .A2(n27860), .ZN(n26676) );
  INV_X1 U34188 ( .A(n26651), .ZN(n29290) );
  NAND2_X2 U1256 ( .A1(n27635), .A2(n22344), .ZN(n27627) );
  INV_X2 U7393 ( .A(n31033), .ZN(n6107) );
  INV_X1 U5349 ( .A(n32784), .ZN(n32157) );
  INV_X2 U2327 ( .A(n31684), .ZN(n31680) );
  BUF_X1 U2067 ( .A(n31113), .Z(n362) );
  NAND3_X1 U3961 ( .A1(n6079), .A2(n26339), .A3(n26338), .ZN(n31700) );
  INV_X1 U12505 ( .A(n32194), .ZN(n32215) );
  INV_X1 U12636 ( .A(n31876), .ZN(n31798) );
  INV_X1 U10553 ( .A(n29591), .ZN(n31106) );
  INV_X1 U10596 ( .A(n32691), .ZN(n30140) );
  INV_X2 U3946 ( .A(n32724), .ZN(n32720) );
  BUF_X1 U2666 ( .A(n31110), .Z(n623) );
  INV_X2 U13909 ( .A(n5111), .ZN(n32540) );
  INV_X2 U5226 ( .A(n32634), .ZN(n32915) );
  NOR2_X2 U3921 ( .A1(n32356), .A2(n32439), .ZN(n32347) );
  INV_X2 U1672 ( .A(n31815), .ZN(n31039) );
  INV_X2 U20503 ( .A(n32883), .ZN(n8544) );
  INV_X1 U36201 ( .A(n32760), .ZN(n32765) );
  INV_X1 U10573 ( .A(n31911), .ZN(n32385) );
  NOR2_X2 U36601 ( .A1(n30982), .A2(n31679), .ZN(n30007) );
  OR2_X2 U13440 ( .A1(n717), .A2(n31425), .ZN(n31420) );
  NAND2_X1 U5265 ( .A1(n30592), .A2(n30601), .ZN(n30590) );
  INV_X1 U10616 ( .A(n30058), .ZN(n31116) );
  INV_X1 U9499 ( .A(n32830), .ZN(n32823) );
  INV_X1 U511 ( .A(n31746), .ZN(n31369) );
  INV_X2 U2645 ( .A(n31385), .ZN(n33017) );
  NOR2_X1 U1331 ( .A1(n26968), .A2(n51742), .ZN(n30946) );
  CLKBUF_X1 U2087 ( .A(n34544), .Z(n375) );
  BUF_X2 U3824 ( .A(n33709), .Z(n703) );
  INV_X1 U3793 ( .A(n7828), .ZN(n37017) );
  INV_X1 U2620 ( .A(n34911), .ZN(n36251) );
  INV_X1 U38604 ( .A(n36359), .ZN(n38018) );
  OR2_X1 U1756 ( .A1(n39429), .A2(n38937), .ZN(n39208) );
  INV_X1 U8112 ( .A(n38035), .ZN(n36372) );
  NAND2_X1 U15013 ( .A1(n38057), .A2(n51522), .ZN(n36167) );
  INV_X1 U2613 ( .A(n36027), .ZN(n6218) );
  INV_X1 U39664 ( .A(n34089), .ZN(n36029) );
  AND2_X1 U3646 ( .A1(n36545), .A2(n37969), .ZN(n36553) );
  NAND2_X1 U18749 ( .A1(n36186), .A2(n39342), .ZN(n39349) );
  INV_X2 U3690 ( .A(n37496), .ZN(n37757) );
  INV_X1 U11496 ( .A(n36051), .ZN(n36459) );
  INV_X1 U11142 ( .A(n36141), .ZN(n35175) );
  OR2_X1 U3702 ( .A1(n37593), .A2(n37378), .ZN(n36233) );
  NAND2_X2 U5827 ( .A1(n5364), .A2(n33562), .ZN(n37520) );
  INV_X1 U1936 ( .A(n38496), .ZN(n38504) );
  AND4_X1 U601 ( .A1(n8013), .A2(n8009), .A3(n37966), .A4(n34091), .ZN(n6286)
         );
  INV_X2 U2579 ( .A(n39768), .ZN(n41436) );
  INV_X1 U20318 ( .A(n39712), .ZN(n8316) );
  INV_X2 U2576 ( .A(n41123), .ZN(n41265) );
  AND2_X2 U8772 ( .A1(n40029), .A2(n41211), .ZN(n5060) );
  INV_X1 U7451 ( .A(n42209), .ZN(n41939) );
  INV_X2 U20533 ( .A(n39906), .ZN(n39908) );
  INV_X1 U14996 ( .A(n40683), .ZN(n40672) );
  INV_X2 U1942 ( .A(n40377), .ZN(n40385) );
  INV_X2 U18618 ( .A(n42018), .ZN(n41588) );
  NOR2_X1 U20003 ( .A1(n41539), .A2(n40986), .ZN(n7985) );
  INV_X1 U9659 ( .A(n41997), .ZN(n42011) );
  INV_X2 U2291 ( .A(n39907), .ZN(n39565) );
  BUF_X1 U870 ( .A(n45459), .Z(n50967) );
  AND4_X1 U3414 ( .A1(n42142), .A2(n42143), .A3(n42141), .A4(n42140), .ZN(
        n42166) );
  NAND3_X2 U45 ( .A1(n270), .A2(n1185), .A3(n8721), .ZN(n51408) );
  XNOR2_X1 U18969 ( .A(n45089), .B(n42458), .ZN(n42534) );
  INV_X1 U17524 ( .A(n46196), .ZN(n49272) );
  INV_X1 U705 ( .A(n48248), .ZN(n48487) );
  INV_X1 U7573 ( .A(n5924), .ZN(n50386) );
  INV_X1 U2553 ( .A(n46693), .ZN(n46901) );
  INV_X1 U45082 ( .A(n48456), .ZN(n46446) );
  INV_X1 U11209 ( .A(n46028), .ZN(n49663) );
  INV_X1 U2525 ( .A(n49667), .ZN(n49659) );
  INV_X2 U1559 ( .A(n42990), .ZN(n49721) );
  NAND2_X1 U673 ( .A1(n52131), .A2(n50294), .ZN(n49956) );
  INV_X1 U20 ( .A(n51690), .ZN(n28) );
  BUF_X1 U7596 ( .A(n7777), .Z(n2178) );
  AND2_X1 U834 ( .A1(n43187), .A2(n43179), .ZN(n1624) );
  INV_X1 U661 ( .A(n49376), .ZN(n49365) );
  INV_X1 U2415 ( .A(n45872), .ZN(n47763) );
  AND2_X1 U1172 ( .A1(n47194), .A2(n47193), .ZN(n49445) );
  INV_X1 U19159 ( .A(n50485), .ZN(n50465) );
  INV_X1 U23239 ( .A(n49029), .ZN(n51397) );
  INV_X2 U15772 ( .A(n50542), .ZN(n50555) );
  NAND4_X2 U2462 ( .A1(n8007), .A2(n8006), .A3(n47047), .A4(n47048), .ZN(
        n50552) );
  INV_X1 U620 ( .A(n47573), .ZN(n47542) );
  INV_X1 U9782 ( .A(n47831), .ZN(n47883) );
  INV_X2 U497 ( .A(n45711), .ZN(n2034) );
  INV_X1 U11150 ( .A(n47745), .ZN(n47797) );
  INV_X2 U2033 ( .A(n45739), .ZN(n1585) );
  INV_X1 U18641 ( .A(n50521), .ZN(n50562) );
  NAND2_X1 U635 ( .A1(n602), .A2(n50235), .ZN(n50227) );
  AND2_X2 U5050 ( .A1(n11489), .A2(n12488), .ZN(n11908) );
  AND3_X2 U13573 ( .A1(n26836), .A2(n26838), .A3(n26837), .ZN(n30102) );
  BUF_X2 U1632 ( .A(n13540), .Z(n17569) );
  AND2_X2 U2293 ( .A1(n5519), .A2(n18063), .ZN(n18071) );
  OR2_X2 U230 ( .A1(n10055), .A2(n8803), .ZN(n9856) );
  AND3_X2 U6204 ( .A1(n1268), .A2(n13212), .A3(n13213), .ZN(n17754) );
  BUF_X2 U3348 ( .A(n44925), .Z(n670) );
  OR2_X2 U6567 ( .A1(n1420), .A2(n372), .ZN(n47858) );
  AND4_X2 U22628 ( .A1(n10156), .A2(n10155), .A3(n10154), .A4(n10153), .ZN(
        n12211) );
  XNOR2_X2 U267 ( .A(n35589), .B(n36685), .ZN(n34238) );
  OR2_X2 U20362 ( .A1(n19619), .A2(n19618), .ZN(n25213) );
  OR2_X2 U19733 ( .A1(n39450), .A2(n39027), .ZN(n39032) );
  NAND2_X2 U7706 ( .A1(n9806), .A2(n52189), .ZN(n10921) );
  INV_X2 U9688 ( .A(n41275), .ZN(n41286) );
  INV_X2 U1628 ( .A(n23020), .ZN(n4413) );
  OR2_X2 U15931 ( .A1(n6906), .A2(n44742), .ZN(n49114) );
  XNOR2_X2 U1664 ( .A(n25481), .B(n26610), .ZN(n24171) );
  OR2_X2 U346 ( .A1(n33026), .A2(n32876), .ZN(n32645) );
  AND2_X2 U8811 ( .A1(n677), .A2(n40377), .ZN(n38612) );
  AND4_X2 U18093 ( .A1(n21786), .A2(n22292), .A3(n21785), .A4(n21784), .ZN(
        n21787) );
  OR2_X2 U1001 ( .A1(n18270), .A2(n18269), .ZN(n22509) );
  BUF_X2 U2649 ( .A(n31608), .Z(n32561) );
  BUF_X2 U1578 ( .A(n21484), .Z(n2220) );
  OR2_X2 U12376 ( .A1(n51196), .A2(n20295), .ZN(n25429) );
  BUF_X2 U234 ( .A(n9234), .Z(n11322) );
  NOR2_X2 U399 ( .A1(n46501), .A2(n46492), .ZN(n46396) );
  OR2_X2 U2112 ( .A1(n6152), .A2(n6151), .ZN(n15132) );
  NAND2_X2 U1299 ( .A1(n3565), .A2(n4229), .ZN(n14139) );
  XNOR2_X2 U4262 ( .A(n25554), .B(n27211), .ZN(n28371) );
  NOR2_X2 U1648 ( .A1(n31302), .A2(n31300), .ZN(n30830) );
  BUF_X2 U2569 ( .A(n44972), .Z(n51096) );
  XNOR2_X2 U14786 ( .A(n4126), .B(n18744), .ZN(n21578) );
  AND3_X2 U18086 ( .A1(n39736), .A2(n41028), .A3(n39735), .ZN(n43374) );
  XNOR2_X2 U7550 ( .A(n43244), .B(n42643), .ZN(n43027) );
  OR2_X2 U4555 ( .A1(n18014), .A2(n19396), .ZN(n18024) );
  AND2_X2 U4991 ( .A1(n9932), .A2(n51650), .ZN(n11707) );
  AND2_X2 U1514 ( .A1(n37667), .A2(n35405), .ZN(n37195) );
  AND3_X2 U20380 ( .A1(n21478), .A2(n21476), .A3(n8395), .ZN(n22521) );
  XNOR2_X2 U19653 ( .A(n25047), .B(n26152), .ZN(n25798) );
  XNOR2_X2 U2163 ( .A(n36885), .B(n35774), .ZN(n38722) );
  NAND2_X2 U787 ( .A1(n10961), .A2(n10055), .ZN(n10955) );
  INV_X2 U2513 ( .A(n47381), .ZN(n602) );
  AND2_X2 U829 ( .A1(n9235), .A2(n10333), .ZN(n10418) );
  BUF_X2 U926 ( .A(n25734), .Z(n28699) );
  CLKBUF_X3 U2085 ( .A(n18261), .Z(n374) );
  INV_X2 U1677 ( .A(n10722), .ZN(n12282) );
  NAND2_X2 U1484 ( .A1(n232), .A2(n2995), .ZN(n30855) );
  OR2_X2 U3386 ( .A1(n39509), .A2(n39510), .ZN(n43354) );
  AND4_X2 U740 ( .A1(n38327), .A2(n38326), .A3(n38325), .A4(n38324), .ZN(
        n38351) );
  AND2_X2 U2253 ( .A1(n38005), .A2(n38018), .ZN(n38173) );
  OR2_X2 U3662 ( .A1(n38587), .A2(n38159), .ZN(n37569) );
  AND4_X2 U1351 ( .A1(n3364), .A2(n24408), .A3(n24407), .A4(n24419), .ZN(n6554) );
  AND2_X2 U9843 ( .A1(n50906), .A2(n51298), .ZN(n50953) );
  AND3_X2 U18241 ( .A1(n6288), .A2(n6289), .A3(n6287), .ZN(n32560) );
  BUF_X2 U5080 ( .A(n9407), .Z(n12112) );
  INV_X2 U4391 ( .A(n22145), .ZN(n22154) );
  BUF_X2 U1084 ( .A(n47013), .Z(n50390) );
  AND2_X2 U18652 ( .A1(n10077), .A2(n9289), .ZN(n10601) );
  AND2_X2 U1228 ( .A1(n37032), .A2(n39369), .ZN(n39381) );
  INV_X2 U2391 ( .A(n13800), .ZN(n13483) );
  AND2_X2 U12104 ( .A1(n10365), .A2(n10366), .ZN(n13800) );
  NAND2_X2 U3949 ( .A1(n28005), .A2(n28006), .ZN(n32974) );
  NOR2_X2 U1130 ( .A1(n50386), .A2(n2199), .ZN(n49742) );
  INV_X2 U3792 ( .A(n6240), .ZN(n35124) );
  OR2_X2 U1257 ( .A1(n3683), .A2(n18888), .ZN(n18992) );
  AND3_X2 U852 ( .A1(n7188), .A2(n7187), .A3(n7186), .ZN(n22434) );
  OAI21_X2 U1480 ( .B1(n38388), .B2(n38387), .A(n38386), .ZN(n43219) );
  AND2_X2 U2852 ( .A1(n799), .A2(n10360), .ZN(n11387) );
  BUF_X2 U4641 ( .A(n19119), .Z(n2182) );
  NOR2_X2 U11096 ( .A1(n50145), .A2(n51727), .ZN(n50113) );
  AND2_X2 U789 ( .A1(n31799), .A2(n31873), .ZN(n31801) );
  AND3_X2 U1262 ( .A1(n10627), .A2(n10626), .A3(n10625), .ZN(n13410) );
  OR2_X2 U14182 ( .A1(n30692), .A2(n51113), .ZN(n30387) );
  NOR2_X2 U1274 ( .A1(n13462), .A2(n51369), .ZN(n15159) );
  NAND2_X2 U15249 ( .A1(n35937), .A2(n35936), .ZN(n41938) );
  OR2_X2 U896 ( .A1(n51107), .A2(n28641), .ZN(n27808) );
  NAND4_X2 U5952 ( .A1(n31278), .A2(n31277), .A3(n31276), .A4(n31279), .ZN(
        n5612) );
  OR2_X2 U4958 ( .A1(n7264), .A2(n12545), .ZN(n12544) );
  AND2_X2 U1499 ( .A1(n5465), .A2(n17878), .ZN(n22359) );
  XNOR2_X2 U20620 ( .A(n18827), .B(n19186), .ZN(n18123) );
  NOR2_X2 U7665 ( .A1(n18988), .A2(n7097), .ZN(n7096) );
  XNOR2_X2 U3805 ( .A(n36747), .B(n33938), .ZN(n34425) );
  AND2_X2 U3836 ( .A1(n2087), .A2(n2088), .ZN(n31374) );
  NAND3_X2 U3385 ( .A1(n41177), .A2(n41176), .A3(n41175), .ZN(n44937) );
  AND2_X2 U3651 ( .A1(n1087), .A2(n37396), .ZN(n37559) );
  OR2_X2 U1708 ( .A1(n27882), .A2(n30209), .ZN(n27097) );
  OR2_X2 U42899 ( .A1(n41695), .A2(n41706), .ZN(n41166) );
  OR2_X2 U8505 ( .A1(n24115), .A2(n24409), .ZN(n24420) );
  OR2_X2 U12005 ( .A1(n2680), .A2(n9667), .ZN(n12338) );
  AND2_X2 U15390 ( .A1(n11352), .A2(n10687), .ZN(n12087) );
  AND2_X2 U1818 ( .A1(n17059), .A2(n18313), .ZN(n20092) );
  AND2_X2 U14154 ( .A1(n49207), .A2(n49197), .ZN(n46226) );
  OR2_X2 U4181 ( .A1(n28187), .A2(n27281), .ZN(n30412) );
  NAND2_X2 U6922 ( .A1(n776), .A2(n20376), .ZN(n20805) );
  NAND3_X2 U1096 ( .A1(n5489), .A2(n38625), .A3(n4510), .ZN(n44198) );
  OR2_X2 U7559 ( .A1(n31358), .A2(n51738), .ZN(n38552) );
  INV_X2 U20110 ( .A(n45763), .ZN(n46633) );
  AND2_X2 U391 ( .A1(n5482), .A2(n37667), .ZN(n38322) );
  AND2_X2 U1888 ( .A1(n10026), .A2(n8853), .ZN(n9484) );
  NAND2_X2 U2353 ( .A1(n6450), .A2(n36579), .ZN(n39674) );
  AND2_X2 U5004 ( .A1(n11662), .A2(n10563), .ZN(n10018) );
  BUF_X2 U1889 ( .A(n10639), .Z(n14346) );
  AND2_X2 U1641 ( .A1(n18921), .A2(n20211), .ZN(n19675) );
  INV_X2 U28169 ( .A(n17287), .ZN(n21276) );
  INV_X2 U48217 ( .A(n46542), .ZN(n48136) );
  XNOR2_X2 U636 ( .A(n8847), .B(Key[75]), .ZN(n10527) );
  AND2_X2 U20357 ( .A1(n8360), .A2(n8359), .ZN(n32027) );
  AND4_X2 U1320 ( .A1(n4686), .A2(n3732), .A3(n13187), .A4(n13188), .ZN(n3313)
         );
  OR2_X2 U2296 ( .A1(n23301), .A2(n27566), .ZN(n29905) );
  CLKBUF_X3 U3040 ( .A(Key[154]), .Z(n4613) );
  NAND4_X2 U37042 ( .A1(n29822), .A2(n29820), .A3(n32687), .A4(n29821), .ZN(
        n35683) );
  BUF_X2 U2244 ( .A(n36881), .Z(n460) );
  AND2_X2 U3925 ( .A1(n1417), .A2(n20147), .ZN(n17065) );
  OR2_X2 U2343 ( .A1(n26494), .A2(n2195), .ZN(n30279) );
  NAND3_X2 U3977 ( .A1(n6772), .A2(n6769), .A3(n30439), .ZN(n31398) );
  AND3_X2 U4443 ( .A1(n18844), .A2(n18845), .A3(n18843), .ZN(n23866) );
  INV_X2 U628 ( .A(n33104), .ZN(n35800) );
  OR2_X2 U8380 ( .A1(n18823), .A2(n777), .ZN(n20600) );
  AND2_X2 U48236 ( .A1(n47620), .A2(n47617), .ZN(n47608) );
  BUF_X2 U4821 ( .A(n11409), .Z(n51141) );
  NAND3_X2 U12333 ( .A1(n29659), .A2(n4697), .A3(n29660), .ZN(n34156) );
  XNOR2_X2 U20168 ( .A(n33835), .B(n34553), .ZN(n36934) );
  XNOR2_X2 U43435 ( .A(n42492), .B(n40998), .ZN(n44076) );
  OAI21_X2 U43426 ( .B1(n39868), .B2(n39869), .A(n39867), .ZN(n42492) );
  AND2_X2 U9711 ( .A1(n40250), .A2(n42205), .ZN(n41942) );
  XNOR2_X2 U1120 ( .A(n25508), .B(n27250), .ZN(n25005) );
  NAND3_X2 U759 ( .A1(n15291), .A2(n1226), .A3(n15289), .ZN(n16660) );
  NOR2_X2 U22197 ( .A1(n9604), .A2(n11411), .ZN(n12138) );
  AND2_X2 U5044 ( .A1(n10968), .A2(n9855), .ZN(n10960) );
  AND2_X2 U2731 ( .A1(n5528), .A2(n23341), .ZN(n22263) );
  OR2_X2 U6018 ( .A1(n22908), .A2(n22367), .ZN(n22165) );
  OR2_X2 U4081 ( .A1(n26039), .A2(n1022), .ZN(n29446) );
  CLKBUF_X3 U1502 ( .A(n33649), .Z(n37545) );
  XNOR2_X2 U1071 ( .A(n8932), .B(Key[39]), .ZN(n12532) );
  NOR2_X4 U531 ( .A1(n10574), .A2(n10573), .ZN(n14339) );
  AND2_X2 U2014 ( .A1(n3352), .A2(n35870), .ZN(n39899) );
  AND2_X2 U266 ( .A1(n38273), .A2(n51339), .ZN(n38291) );
  BUF_X2 U35308 ( .A(n27158), .Z(n30721) );
  AND4_X2 U3837 ( .A1(n6156), .A2(n31962), .A3(n1566), .A4(n6155), .ZN(n33104)
         );
  BUF_X2 U4846 ( .A(n10208), .Z(n14186) );
  XNOR2_X2 U12560 ( .A(n46058), .B(n42284), .ZN(n44338) );
  NAND3_X2 U4894 ( .A1(n12666), .A2(n4560), .A3(n4559), .ZN(n15309) );
  AND2_X2 U614 ( .A1(n21392), .A2(n20375), .ZN(n20416) );
  XNOR2_X2 U21197 ( .A(n8817), .B(Key[14]), .ZN(n10161) );
  NAND2_X2 U9761 ( .A1(n4066), .A2(n22634), .ZN(n27451) );
  BUF_X1 U975 ( .A(n31768), .Z(n50980) );
  CLKBUF_X3 U41920 ( .A(n37345), .Z(n40458) );
  BUF_X2 U2095 ( .A(n31545), .Z(n382) );
  BUF_X2 U3300 ( .A(n42886), .Z(n49689) );
  NAND2_X2 U2556 ( .A1(n51283), .A2(n41022), .ZN(n43890) );
  BUF_X2 U50143 ( .A(n49766), .Z(n49871) );
  AND4_X2 U1050 ( .A1(n24986), .A2(n2830), .A3(n8136), .A4(n24987), .ZN(n32214) );
  NAND4_X2 U2844 ( .A1(n9832), .A2(n9834), .A3(n9831), .A4(n9833), .ZN(n1571)
         );
  OR2_X2 U12055 ( .A1(n17003), .A2(n17004), .ZN(n23513) );
  NAND2_X2 U4703 ( .A1(n4106), .A2(n5551), .ZN(n16571) );
  BUF_X2 U35919 ( .A(n28082), .Z(n29797) );
  NAND2_X2 U808 ( .A1(n5800), .A2(n8254), .ZN(n25825) );
  OR2_X2 U19095 ( .A1(n37765), .A2(n7083), .ZN(n37501) );
  AND2_X2 U3742 ( .A1(n20704), .A2(n20705), .ZN(n23374) );
  XNOR2_X2 U1342 ( .A(n35345), .B(n32952), .ZN(n515) );
  NOR2_X2 U23109 ( .A1(n51683), .A2(n13525), .ZN(n13512) );
  AND4_X2 U4434 ( .A1(n20485), .A2(n8594), .A3(n8593), .A4(n8591), .ZN(n8590)
         );
  AND2_X2 U485 ( .A1(n6853), .A2(n25198), .ZN(n28025) );
  INV_X2 U1714 ( .A(n11049), .ZN(n14036) );
  AND2_X2 U16902 ( .A1(n5111), .A2(n8681), .ZN(n32899) );
  NAND4_X2 U1379 ( .A1(n15268), .A2(n15269), .A3(n15267), .A4(n15270), .ZN(
        n16749) );
  NAND2_X2 U1571 ( .A1(n7710), .A2(n12772), .ZN(n16919) );
  NAND4_X2 U14633 ( .A1(n21552), .A2(n21553), .A3(n21554), .A4(n21551), .ZN(
        n23129) );
  NAND2_X2 U6038 ( .A1(n1207), .A2(n41636), .ZN(n44901) );
  NAND3_X2 U19273 ( .A1(n31228), .A2(n31227), .A3(n7251), .ZN(n35745) );
  AND2_X2 U5037 ( .A1(n10069), .A2(n9476), .ZN(n9908) );
  AND2_X2 U5673 ( .A1(n21547), .A2(n20642), .ZN(n21541) );
  AND2_X2 U3648 ( .A1(n34676), .A2(n37543), .ZN(n37554) );
  NAND4_X2 U1385 ( .A1(n11847), .A2(n11849), .A3(n11848), .A4(n11850), .ZN(
        n17730) );
  AND2_X2 U8083 ( .A1(n37191), .A2(n35409), .ZN(n35894) );
  OAI21_X2 U2796 ( .B1(n38346), .B2(n38347), .A(n38345), .ZN(n38348) );
  AND3_X2 U38445 ( .A1(n32349), .A2(n32350), .A3(n32348), .ZN(n32364) );
  BUF_X1 U30413 ( .A(n40838), .Z(n51455) );
  OR2_X4 U1465 ( .A1(n7257), .A2(n7260), .ZN(n25064) );
  BUF_X2 U20665 ( .A(n7592), .Z(n51362) );
  XNOR2_X2 U958 ( .A(n8822), .B(Key[117]), .ZN(n10579) );
  NAND2_X2 U1764 ( .A1(n3266), .A2(n3175), .ZN(n26304) );
  NAND2_X2 U1293 ( .A1(n4814), .A2(n7154), .ZN(n45339) );
  BUF_X2 U2271 ( .A(n38972), .Z(n473) );
  OR2_X2 U907 ( .A1(n6343), .A2(n38701), .ZN(n38706) );
  BUF_X2 U2309 ( .A(n19336), .Z(n489) );
  OR2_X2 U4871 ( .A1(n10691), .A2(n10690), .ZN(n14011) );
  NOR2_X2 U3915 ( .A1(n32701), .A2(n32324), .ZN(n32704) );
  OR2_X2 U10181 ( .A1(n21199), .A2(n19819), .ZN(n21218) );
  NOR2_X2 U17774 ( .A1(n5875), .A2(n20432), .ZN(n20349) );
  OR2_X2 U1137 ( .A1(n10628), .A2(n10535), .ZN(n10639) );
  INV_X2 U2621 ( .A(n37646), .ZN(n36410) );
  INV_X2 U18413 ( .A(n40740), .ZN(n6469) );
  AND2_X2 U729 ( .A1(n38701), .A2(n6343), .ZN(n39236) );
  OR2_X2 U43968 ( .A1(n40756), .A2(n40755), .ZN(n41629) );
  INV_X2 U21662 ( .A(n9148), .ZN(n11705) );
  OR2_X2 U12668 ( .A1(n664), .A2(n49163), .ZN(n46244) );
  BUF_X2 U4994 ( .A(n9142), .Z(n11696) );
  OR2_X2 U7209 ( .A1(n46446), .A2(n42508), .ZN(n46449) );
  XNOR2_X2 U17301 ( .A(n37137), .B(n36829), .ZN(n5445) );
  INV_X2 U104 ( .A(n32867), .ZN(n32882) );
  NOR2_X2 U4442 ( .A1(n17473), .A2(n17472), .ZN(n21748) );
  AND2_X2 U10066 ( .A1(n13514), .A2(n11841), .ZN(n13509) );
  NAND4_X2 U2188 ( .A1(n22743), .A2(n22746), .A3(n22744), .A4(n22745), .ZN(
        n24556) );
  NAND4_X2 U20695 ( .A1(n45169), .A2(n47010), .A3(n45168), .A4(n45167), .ZN(
        n45194) );
  NOR2_X2 U11824 ( .A1(n51117), .A2(n26944), .ZN(n27660) );
  NOR2_X2 U12405 ( .A1(n6469), .A2(n41348), .ZN(n40736) );
  XNOR2_X2 U4786 ( .A(n9402), .B(Key[167]), .ZN(n51391) );
  INV_X2 U38035 ( .A(n32732), .ZN(n31648) );
  XNOR2_X2 U1029 ( .A(n9401), .B(Key[64]), .ZN(n9405) );
  AND2_X2 U16021 ( .A1(n5056), .A2(n28862), .ZN(n5054) );
  NAND4_X2 U3394 ( .A1(n40735), .A2(n3682), .A3(n40734), .A4(n3681), .ZN(
        n44208) );
  BUF_X2 U80 ( .A(n33336), .Z(n619) );
  NOR2_X2 U37024 ( .A1(n32724), .A2(n32316), .ZN(n32464) );
  NOR2_X1 U1255 ( .A1(n8224), .A2(n23547), .ZN(n23551) );
  AND2_X2 U1174 ( .A1(n18010), .A2(n17479), .ZN(n19395) );
  AND3_X2 U45136 ( .A1(n16493), .A2(n16495), .A3(n7987), .ZN(n21947) );
  BUF_X2 U5412 ( .A(n16470), .Z(n485) );
  AND2_X2 U403 ( .A1(n36604), .A2(n36429), .ZN(n36425) );
  AND2_X2 U9918 ( .A1(n52185), .A2(n10074), .ZN(n9915) );
  AND2_X2 U1623 ( .A1(n783), .A2(n13633), .ZN(n14672) );
  AND3_X2 U3423 ( .A1(n38848), .A2(n38850), .A3(n38847), .ZN(n6713) );
  OR2_X2 U10775 ( .A1(n40003), .A2(n39101), .ZN(n6965) );
  INV_X2 U4394 ( .A(n16849), .ZN(n21970) );
  XNOR2_X2 U31412 ( .A(n51465), .B(n41187), .ZN(n45432) );
  AND2_X2 U1521 ( .A1(n49770), .A2(n49771), .ZN(n49782) );
  NAND2_X2 U18109 ( .A1(n30096), .A2(n30095), .ZN(n35325) );
  BUF_X2 U1422 ( .A(n50339), .Z(n51026) );
  XNOR2_X2 U1412 ( .A(n24667), .B(n24666), .ZN(n29413) );
  NOR2_X2 U6405 ( .A1(n30924), .A2(n30930), .ZN(n31055) );
  AND2_X4 U7804 ( .A1(n3037), .A2(n3753), .ZN(n32175) );
  NOR2_X2 U4172 ( .A1(n29413), .A2(n51679), .ZN(n26985) );
  NOR2_X2 U5773 ( .A1(n21186), .A2(n21181), .ZN(n19703) );
  AND3_X2 U2583 ( .A1(n34214), .A2(n34213), .A3(n6714), .ZN(n39855) );
  AND4_X2 U1730 ( .A1(n13360), .A2(n13359), .A3(n13358), .A4(n13357), .ZN(
        n13365) );
  NAND2_X2 U16012 ( .A1(n11940), .A2(n8470), .ZN(n15434) );
  NAND2_X2 U32256 ( .A1(n23383), .A2(n23384), .ZN(n28423) );
  XNOR2_X2 U7515 ( .A(n34448), .B(n34449), .ZN(n2123) );
  BUF_X2 U26242 ( .A(n16201), .Z(n18505) );
  BUF_X2 U27924 ( .A(n17005), .Z(n24290) );
  AND2_X2 U46265 ( .A1(n51725), .A2(n555), .ZN(n47291) );
  INV_X2 U25891 ( .A(n15154), .ZN(n18437) );
  OR2_X4 U12116 ( .A1(n35970), .A2(n35969), .ZN(n40250) );
  NOR2_X2 U26950 ( .A1(n21521), .A2(n20614), .ZN(n20175) );
  NOR2_X2 U50535 ( .A1(n50459), .A2(n50485), .ZN(n50470) );
  NAND4_X4 U7149 ( .A1(n10353), .A2(n10352), .A3(n10350), .A4(n10351), .ZN(
        n13801) );
  CLKBUF_X3 U38501 ( .A(n32801), .Z(n34835) );
  BUF_X2 U7519 ( .A(n34844), .Z(n2129) );
  AND2_X2 U20582 ( .A1(n8629), .A2(n18250), .ZN(n20298) );
  OR2_X2 U20991 ( .A1(n37901), .A2(n39410), .ZN(n37907) );
  BUF_X2 U2228 ( .A(n26458), .Z(n28918) );
  INV_X2 U4433 ( .A(n20787), .ZN(n23641) );
  NOR2_X2 U9216 ( .A1(n22736), .A2(n22386), .ZN(n22742) );
  XNOR2_X2 U16999 ( .A(n5201), .B(n5200), .ZN(n17057) );
  XNOR2_X2 U6250 ( .A(n44027), .B(n5032), .ZN(n43575) );
  NAND2_X2 U6316 ( .A1(n23809), .A2(n30667), .ZN(n27608) );
  XNOR2_X2 U3359 ( .A(n44547), .B(n43781), .ZN(n43642) );
  OR2_X2 U10826 ( .A1(n41702), .A2(n41692), .ZN(n41689) );
  INV_X2 U452 ( .A(n14341), .ZN(n6073) );
  BUF_X2 U2084 ( .A(n18261), .Z(n373) );
  NOR2_X2 U36006 ( .A1(n28174), .A2(n28173), .ZN(n32741) );
  OR2_X2 U9334 ( .A1(n27139), .A2(n2568), .ZN(n27995) );
  OR2_X2 U9663 ( .A1(n37892), .A2(n6825), .ZN(n39407) );
  BUF_X2 U235 ( .A(n9335), .Z(n9969) );
  NAND4_X4 U35588 ( .A1(n27532), .A2(n27530), .A3(n27531), .A4(n27533), .ZN(
        n32788) );
  NAND2_X2 U849 ( .A1(n5377), .A2(n27779), .ZN(n37262) );
  INV_X2 U20001 ( .A(n26804), .ZN(n27732) );
  BUF_X2 U2102 ( .A(n13323), .Z(n14600) );
  XNOR2_X2 U7846 ( .A(n7608), .B(n44963), .ZN(n43349) );
  AND2_X2 U836 ( .A1(n12323), .A2(n9668), .ZN(n12344) );
  OR2_X2 U2599 ( .A1(n695), .A2(n34189), .ZN(n34963) );
  OR2_X2 U14375 ( .A1(n39765), .A2(n3979), .ZN(n43547) );
  BUF_X2 U226 ( .A(n12145), .Z(n438) );
  INV_X2 U6387 ( .A(n48834), .ZN(n48817) );
  OR2_X2 U4595 ( .A1(n51130), .A2(n20474), .ZN(n17999) );
  INV_X2 U7983 ( .A(n23175), .ZN(n5269) );
  NAND4_X2 U1892 ( .A1(n28648), .A2(n28649), .A3(n28647), .A4(n28646), .ZN(
        n31637) );
  OR2_X2 U395 ( .A1(n28723), .A2(n30856), .ZN(n31630) );
  XNOR2_X2 U521 ( .A(n25318), .B(n25317), .ZN(n29346) );
  NOR2_X2 U10960 ( .A1(n40458), .A2(n40403), .ZN(n39990) );
  AOI22_X2 U9593 ( .A1(n9381), .A2(n9382), .B1(n9383), .B2(n11390), .ZN(n9392)
         );
  OR2_X2 U30926 ( .A1(n21071), .A2(n21070), .ZN(n24256) );
  AND2_X2 U10478 ( .A1(n29332), .A2(n29315), .ZN(n27896) );
  BUF_X2 U2247 ( .A(n18535), .Z(n462) );
  NAND4_X4 U4892 ( .A1(n11267), .A2(n11264), .A3(n11266), .A4(n11265), .ZN(
        n14410) );
  XNOR2_X2 U1169 ( .A(n8896), .B(Key[58]), .ZN(n8909) );
  AND2_X2 U4990 ( .A1(n10831), .A2(n12502), .ZN(n11550) );
  OAI211_X2 U7581 ( .C1(n47134), .C2(n46677), .A(n46663), .B(n46662), .ZN(
        n47599) );
  NAND3_X2 U1443 ( .A1(n30989), .A2(n30988), .A3(n2974), .ZN(n7787) );
  NAND2_X2 U7047 ( .A1(n18000), .A2(n19370), .ZN(n1789) );
  BUF_X2 U2116 ( .A(n7877), .Z(n395) );
  XNOR2_X2 U2360 ( .A(n3669), .B(n7351), .ZN(n24319) );
  AND4_X2 U20879 ( .A1(n16806), .A2(n16805), .A3(n18358), .A4(n19074), .ZN(
        n16813) );
  INV_X2 U20045 ( .A(n23479), .ZN(n21981) );
  OR2_X2 U4098 ( .A1(n28139), .A2(n5056), .ZN(n28458) );
  AND2_X4 U20456 ( .A1(n8492), .A2(n8491), .ZN(n24190) );
  MUX2_X2 U26735 ( .A(n20670), .B(n20678), .S(n1597), .Z(n20239) );
  BUF_X2 U2049 ( .A(n15102), .Z(n352) );
  BUF_X2 U1383 ( .A(n12542), .Z(n442) );
  BUF_X2 U4249 ( .A(n28312), .Z(n749) );
  OR2_X2 U12764 ( .A1(n3005), .A2(n9053), .ZN(n14317) );
  INV_X2 U3913 ( .A(n32974), .ZN(n2037) );
  OR2_X2 U4109 ( .A1(n30179), .A2(n2201), .ZN(n29140) );
  OR2_X2 U4865 ( .A1(n805), .A2(n8796), .ZN(n12359) );
  INV_X2 U14071 ( .A(n19277), .ZN(n20825) );
  OR2_X2 U7886 ( .A1(n51683), .A2(n13514), .ZN(n13529) );
  NAND2_X2 U7173 ( .A1(n15928), .A2(n51090), .ZN(n5373) );
  XNOR2_X2 U2453 ( .A(n16392), .B(n16391), .ZN(n18377) );
  NAND2_X2 U517 ( .A1(n21656), .A2(n1704), .ZN(n20650) );
  AND2_X2 U3669 ( .A1(n33562), .A2(n38495), .ZN(n37517) );
  BUF_X2 U5025 ( .A(n9140), .Z(n9499) );
  NAND4_X2 U33896 ( .A1(n25409), .A2(n25408), .A3(n25407), .A4(n25406), .ZN(
        n35835) );
  AND2_X2 U47994 ( .A1(n9598), .A2(n10398), .ZN(n12141) );
  NAND2_X2 U28328 ( .A1(n19823), .A2(n2229), .ZN(n21215) );
  BUF_X2 U5012 ( .A(n9308), .Z(n11641) );
  AND2_X2 U700 ( .A1(n35923), .A2(n34911), .ZN(n37762) );
  NOR2_X2 U1534 ( .A1(n24213), .A2(n24214), .ZN(n1778) );
  AND3_X2 U4206 ( .A1(n14697), .A2(n14696), .A3(n51237), .ZN(n14698) );
  BUF_X2 U174 ( .A(n15997), .Z(n21630) );
  OR2_X2 U22424 ( .A1(n9847), .A2(n9846), .ZN(n13948) );
  BUF_X2 U15232 ( .A(n15400), .Z(n18039) );
  INV_X2 U31 ( .A(n41518), .ZN(n42938) );
  OR2_X2 U2817 ( .A1(n14033), .A2(n13291), .ZN(n13296) );
  OR2_X2 U1733 ( .A1(n17466), .A2(n18032), .ZN(n19408) );
  NAND2_X2 U5144 ( .A1(n26972), .A2(n814), .ZN(n34533) );
  OR2_X2 U41088 ( .A1(n42201), .A2(n41938), .ZN(n41925) );
  NOR2_X2 U5700 ( .A1(n3745), .A2(n17639), .ZN(n20483) );
  AND2_X2 U3680 ( .A1(n39299), .A2(n39291), .ZN(n39293) );
  AND2_X2 U6497 ( .A1(n30982), .A2(n51240), .ZN(n31690) );
  INV_X2 U2323 ( .A(n29998), .ZN(n51240) );
  AND2_X2 U319 ( .A1(n40670), .A2(n40671), .ZN(n5062) );
  OR2_X2 U4748 ( .A1(n14445), .A2(n14433), .ZN(n14438) );
  NAND4_X2 U1052 ( .A1(n23236), .A2(n23234), .A3(n23235), .A4(n23233), .ZN(
        n26375) );
  NAND4_X2 U2727 ( .A1(n23740), .A2(n23739), .A3(n23738), .A4(n23737), .ZN(
        n25444) );
  AND3_X4 U4449 ( .A1(n980), .A2(n8324), .A3(n17563), .ZN(n22140) );
  NAND2_X2 U641 ( .A1(n12695), .A2(n12690), .ZN(n12710) );
  AND2_X2 U348 ( .A1(n52198), .A2(n3490), .ZN(n41246) );
  OR2_X2 U4981 ( .A1(n10097), .A2(n10096), .ZN(n9835) );
  NAND4_X2 U36 ( .A1(n38904), .A2(n38905), .A3(n38902), .A4(n38903), .ZN(n5379) );
  XNOR2_X2 U20675 ( .A(n34874), .B(n34873), .ZN(n34906) );
  OR2_X2 U33891 ( .A1(n50981), .A2(n32211), .ZN(n30893) );
  NOR2_X2 U8904 ( .A1(n50222), .A2(n50235), .ZN(n50187) );
  XNOR2_X2 U2144 ( .A(n9202), .B(Key[26]), .ZN(n9207) );
  AND2_X2 U22748 ( .A1(n15034), .A2(n13804), .ZN(n13798) );
  XNOR2_X2 U21784 ( .A(n9243), .B(Key[45]), .ZN(n11403) );
  INV_X2 U12870 ( .A(n10563), .ZN(n11660) );
  XNOR2_X2 U533 ( .A(n9304), .B(Key[66]), .ZN(n10563) );
  XNOR2_X2 U4241 ( .A(n25346), .B(n24849), .ZN(n25805) );
  NAND2_X2 U2412 ( .A1(n834), .A2(n20979), .ZN(n24849) );
  AOI22_X2 U2676 ( .A1(n40068), .A2(n40067), .B1(n40586), .B2(n40066), .ZN(
        n40079) );
  NAND4_X2 U2151 ( .A1(n22726), .A2(n22723), .A3(n22724), .A4(n22725), .ZN(
        n25229) );
  AND2_X2 U22303 ( .A1(n26288), .A2(n28623), .ZN(n28614) );
  BUF_X2 U2505 ( .A(n47381), .Z(n50196) );
  OR2_X2 U1713 ( .A1(n14030), .A2(n14022), .ZN(n11049) );
  INV_X2 U2806 ( .A(n13221), .ZN(n13971) );
  OAI21_X1 U945 ( .B1(n38343), .B2(n38344), .A(n38342), .ZN(n38349) );
  AND2_X2 U34713 ( .A1(n28923), .A2(n28926), .ZN(n28566) );
  XNOR2_X2 U467 ( .A(n9361), .B(Key[36]), .ZN(n10686) );
  INV_X2 U4421 ( .A(n23895), .ZN(n23913) );
  XNOR2_X2 U21168 ( .A(n8799), .B(Key[145]), .ZN(n8803) );
  NAND2_X2 U19179 ( .A1(n4012), .A2(n7327), .ZN(n14149) );
  AND2_X2 U4963 ( .A1(n10925), .A2(n10147), .ZN(n10222) );
  INV_X2 U7666 ( .A(n20095), .ZN(n16788) );
  XNOR2_X2 U2195 ( .A(n1138), .B(n16764), .ZN(n20095) );
  BUF_X2 U34216 ( .A(n25789), .Z(n29478) );
  NAND2_X2 U1233 ( .A1(n51726), .A2(n51514), .ZN(n29174) );
  XNOR2_X2 U38859 ( .A(n35106), .B(n33145), .ZN(n33729) );
  OR2_X2 U16937 ( .A1(n50611), .A2(n50618), .ZN(n50624) );
  OR2_X2 U10045 ( .A1(n2189), .A2(n15770), .ZN(n15073) );
  AND2_X2 U17135 ( .A1(n21975), .A2(n23480), .ZN(n21987) );
  INV_X2 U3229 ( .A(n50980), .ZN(n51103) );
  INV_X2 U6380 ( .A(n11028), .ZN(n11035) );
  AND2_X2 U4823 ( .A1(n15161), .A2(n6384), .ZN(n15168) );
  NAND4_X4 U25103 ( .A1(n14014), .A2(n14013), .A3(n14016), .A4(n14015), .ZN(
        n17938) );
  AND2_X2 U4979 ( .A1(n9641), .A2(n10694), .ZN(n9696) );
  AND4_X2 U413 ( .A1(n15099), .A2(n4867), .A3(n15098), .A4(n2644), .ZN(n4866)
         );
  INV_X2 U2789 ( .A(n6952), .ZN(n633) );
  OR2_X2 U3791 ( .A1(n6518), .A2(n6519), .ZN(n34514) );
  INV_X2 U2657 ( .A(n29618), .ZN(n32988) );
  NAND3_X2 U16379 ( .A1(n2292), .A2(n4807), .A3(n19920), .ZN(n27177) );
  NAND2_X2 U1652 ( .A1(n12297), .A2(n12298), .ZN(n14712) );
  NAND2_X2 U18140 ( .A1(n7020), .A2(n12278), .ZN(n12276) );
  NAND2_X2 U2849 ( .A1(n12630), .A2(n5220), .ZN(n12616) );
  BUF_X2 U5062 ( .A(n8949), .Z(n11443) );
  OR2_X2 U1959 ( .A1(n15394), .A2(n15393), .ZN(n305) );
  NAND2_X2 U2392 ( .A1(n5180), .A2(n12502), .ZN(n12504) );
  XNOR2_X2 U2239 ( .A(Key[106]), .B(Ciphertext[3]), .ZN(n10662) );
  INV_X2 U14687 ( .A(n13148), .ZN(n14179) );
  AND4_X2 U4907 ( .A1(n12552), .A2(n6406), .A3(n12551), .A4(n6407), .ZN(n6405)
         );
  BUF_X2 U12450 ( .A(n23858), .Z(n51492) );
  NAND4_X2 U18272 ( .A1(n34329), .A2(n34328), .A3(n34327), .A4(n34326), .ZN(
        n51307) );
  OAI21_X2 U12667 ( .B1(n15043), .B2(n15042), .A(n15047), .ZN(n2981) );
  INV_X2 U1336 ( .A(n9308), .ZN(n11662) );
  NAND2_X1 U13732 ( .A1(n10077), .A2(n10074), .ZN(n10618) );
  AND2_X1 U13186 ( .A1(n10004), .A2(n11028), .ZN(n11032) );
  NAND2_X1 U240 ( .A1(n10662), .A2(n12057), .ZN(n12051) );
  BUF_X1 U2261 ( .A(n14029), .Z(n469) );
  BUF_X1 U2823 ( .A(n12788), .Z(n12894) );
  BUF_X1 U1251 ( .A(n9721), .Z(n13855) );
  INV_X1 U4836 ( .A(n14149), .ZN(n13122) );
  OR2_X1 U18121 ( .A1(n10877), .A2(n15173), .ZN(n15178) );
  AND2_X1 U9007 ( .A1(n14170), .A2(n14006), .ZN(n14175) );
  BUF_X1 U3035 ( .A(Key[171]), .Z(n1224) );
  NOR2_X2 U980 ( .A1(n15206), .A2(n14767), .ZN(n14769) );
  OAI21_X1 U10122 ( .B1(n9167), .B2(n14642), .A(n13645), .ZN(n14561) );
  OR2_X1 U22435 ( .A1(n9870), .A2(n9869), .ZN(n15758) );
  AND2_X1 U1737 ( .A1(n14092), .A2(n14093), .ZN(n16142) );
  AOI22_X1 U5139 ( .A1(n14449), .A2(n14448), .B1(n14447), .B2(n14446), .ZN(
        n14461) );
  AND3_X1 U4679 ( .A1(n7852), .A2(n13120), .A3(n13121), .ZN(n18669) );
  NAND3_X1 U18235 ( .A1(n6278), .A2(n11053), .A3(n11054), .ZN(n18602) );
  BUF_X1 U245 ( .A(n16162), .Z(n15957) );
  INV_X1 U6440 ( .A(n17526), .ZN(n16798) );
  BUF_X1 U16094 ( .A(n15871), .Z(n18863) );
  NAND2_X1 U507 ( .A1(n20201), .A2(n20641), .ZN(n20745) );
  BUF_X1 U1583 ( .A(n17401), .Z(n19823) );
  NAND2_X1 U26658 ( .A1(n20683), .A2(n20677), .ZN(n18101) );
  NOR2_X1 U26160 ( .A1(n17627), .A2(n18085), .ZN(n19348) );
  INV_X1 U8414 ( .A(n21620), .ZN(n21629) );
  NAND2_X1 U13746 ( .A1(n19156), .A2(n52139), .ZN(n19957) );
  NAND4_X1 U466 ( .A1(n19964), .A2(n19963), .A3(n19962), .A4(n19961), .ZN(
        n22101) );
  MUX2_X1 U4468 ( .A(n18918), .B(n18228), .S(n51006), .Z(n18242) );
  INV_X1 U8433 ( .A(n22506), .ZN(n22492) );
  BUF_X1 U812 ( .A(n22101), .Z(n24033) );
  NAND4_X1 U4278 ( .A1(n19585), .A2(n19584), .A3(n19583), .A4(n19582), .ZN(
        n28427) );
  BUF_X1 U33369 ( .A(n24842), .Z(n26571) );
  OR2_X1 U853 ( .A1(n8640), .A2(n51721), .ZN(n29899) );
  NAND2_X1 U19879 ( .A1(n29028), .A2(n28882), .ZN(n28875) );
  OR2_X1 U5981 ( .A1(n51118), .A2(n28588), .ZN(n28577) );
  AND2_X1 U125 ( .A1(n26671), .A2(n27858), .ZN(n28671) );
  NAND4_X2 U2141 ( .A1(n28595), .A2(n28594), .A3(n28593), .A4(n28592), .ZN(
        n32705) );
  NAND4_X2 U7589 ( .A1(n27144), .A2(n27141), .A3(n27143), .A4(n27142), .ZN(
        n31986) );
  AND2_X2 U17756 ( .A1(n30680), .A2(n30681), .ZN(n31452) );
  INV_X1 U3956 ( .A(n31995), .ZN(n32511) );
  INV_X1 U3963 ( .A(n32056), .ZN(n718) );
  INV_X1 U677 ( .A(n33252), .ZN(n35386) );
  XNOR2_X1 U1481 ( .A(n35749), .B(n5997), .ZN(n36818) );
  XNOR2_X1 U3725 ( .A(n2691), .B(n5448), .ZN(n36051) );
  BUF_X1 U11241 ( .A(n33067), .Z(n38196) );
  AND2_X1 U39750 ( .A1(n36473), .A2(n36567), .ZN(n35315) );
  BUF_X1 U35090 ( .A(n38664), .Z(n51496) );
  BUF_X1 U3751 ( .A(n35409), .Z(n37665) );
  NAND3_X1 U3596 ( .A1(n37602), .A2(n8339), .A3(n37600), .ZN(n39576) );
  BUF_X1 U2455 ( .A(n39944), .Z(n575) );
  INV_X1 U18702 ( .A(n39855), .ZN(n40340) );
  BUF_X2 U2298 ( .A(n40792), .Z(n426) );
  OR2_X1 U9704 ( .A1(n41195), .A2(n41212), .ZN(n40662) );
  AND2_X1 U42 ( .A1(n39316), .A2(n41670), .ZN(n41683) );
  OR2_X1 U7536 ( .A1(n40327), .A2(n40330), .ZN(n40337) );
  BUF_X1 U1508 ( .A(n42778), .Z(n44562) );
  BUF_X1 U1604 ( .A(n41875), .Z(n43113) );
  BUF_X1 U26 ( .A(n42684), .Z(n49207) );
  NAND2_X1 U518 ( .A1(n45772), .A2(n45138), .ZN(n47118) );
  AND2_X1 U47303 ( .A1(n45614), .A2(n51732), .ZN(n48450) );
  NOR2_X2 U32403 ( .A1(n666), .A2(n49263), .ZN(n49275) );
  AND2_X1 U45926 ( .A1(n588), .A2(n49684), .ZN(n49251) );
  AND3_X1 U3 ( .A1(n50018), .A2(n6413), .A3(n50017), .ZN(n51442) );
  BUF_X1 U4 ( .A(n48904), .Z(n51688) );
  AND2_X1 U5 ( .A1(n44813), .A2(n44640), .ZN(n45524) );
  AND2_X1 U11 ( .A1(n45631), .A2(n46464), .ZN(n48535) );
  AND2_X1 U18 ( .A1(n52136), .A2(n45661), .ZN(n46492) );
  BUF_X2 U22 ( .A(n42590), .Z(n43380) );
  NAND3_X1 U47 ( .A1(n6480), .A2(n39535), .A3(n39536), .ZN(n43254) );
  AND2_X1 U62 ( .A1(n6468), .A2(n41348), .ZN(n41345) );
  NOR2_X1 U66 ( .A1(n41374), .A2(n40960), .ZN(n40970) );
  NAND2_X2 U67 ( .A1(n8553), .A2(n8554), .ZN(n52120) );
  BUF_X1 U70 ( .A(n41800), .Z(n51684) );
  AND2_X1 U77 ( .A1(n35026), .A2(n36362), .ZN(n38177) );
  INV_X1 U98 ( .A(n35531), .ZN(n38514) );
  XNOR2_X2 U127 ( .A(n7827), .B(n34178), .ZN(n36567) );
  BUF_X1 U131 ( .A(n37135), .Z(n518) );
  NOR2_X2 U136 ( .A1(n26967), .A2(n26966), .ZN(n52121) );
  BUF_X1 U140 ( .A(n29278), .Z(n51706) );
  NOR2_X1 U155 ( .A1(n30178), .A2(n25198), .ZN(n547) );
  XNOR2_X1 U158 ( .A(n25732), .B(n25731), .ZN(n26651) );
  BUF_X1 U163 ( .A(n25770), .Z(n51720) );
  BUF_X1 U175 ( .A(n23957), .Z(n559) );
  BUF_X2 U178 ( .A(n23564), .Z(n51676) );
  NAND4_X1 U182 ( .A1(n14392), .A2(n14391), .A3(n14390), .A4(n14389), .ZN(
        n21122) );
  BUF_X1 U187 ( .A(n15630), .Z(n19663) );
  BUF_X1 U196 ( .A(n16662), .Z(n51703) );
  BUF_X2 U209 ( .A(n11543), .Z(n51709) );
  AND2_X2 U210 ( .A1(n39400), .A2(n39395), .ZN(n37890) );
  BUF_X1 U211 ( .A(n12534), .Z(n51672) );
  NAND2_X2 U218 ( .A1(n48534), .A2(n46463), .ZN(n48526) );
  OR2_X4 U224 ( .A1(n52267), .A2(n15930), .ZN(n24157) );
  AND2_X2 U241 ( .A1(n38628), .A2(n51360), .ZN(n38641) );
  NAND2_X2 U251 ( .A1(n3493), .A2(n21425), .ZN(n20838) );
  AND2_X2 U253 ( .A1(n8803), .A2(n10967), .ZN(n10965) );
  INV_X2 U261 ( .A(n47989), .ZN(n47988) );
  OR2_X2 U262 ( .A1(n1075), .A2(n33870), .ZN(n37810) );
  BUF_X2 U264 ( .A(n9235), .Z(n10328) );
  AND2_X2 U270 ( .A1(n26973), .A2(n29532), .ZN(n29521) );
  OR2_X2 U275 ( .A1(n51111), .A2(n27695), .ZN(n29563) );
  BUF_X1 U282 ( .A(n9806), .Z(n10920) );
  AND4_X2 U284 ( .A1(n8325), .A2(n8326), .A3(n9494), .A4(n9355), .ZN(n4056) );
  NAND3_X2 U286 ( .A1(n25203), .A2(n25204), .A3(n51790), .ZN(n32211) );
  OR2_X2 U290 ( .A1(n7625), .A2(n51106), .ZN(n32622) );
  NAND2_X2 U292 ( .A1(n20825), .A2(n19280), .ZN(n21480) );
  OR2_X2 U295 ( .A1(n45209), .A2(n44784), .ZN(n45649) );
  NAND2_X2 U299 ( .A1(n36647), .A2(n36648), .ZN(n40683) );
  OR2_X4 U304 ( .A1(n5932), .A2(n5931), .ZN(n32595) );
  AND2_X2 U305 ( .A1(n18362), .A2(n1417), .ZN(n19070) );
  OR2_X2 U311 ( .A1(n22908), .A2(n22918), .ZN(n22360) );
  AND4_X4 U312 ( .A1(n35903), .A2(n52342), .A3(n35902), .A4(n35901), .ZN(
        n38448) );
  AND2_X2 U317 ( .A1(n5593), .A2(n38732), .ZN(n37659) );
  AND2_X2 U325 ( .A1(n22701), .A2(n21780), .ZN(n3553) );
  AND2_X2 U330 ( .A1(n49366), .A2(n51729), .ZN(n49342) );
  NAND2_X2 U343 ( .A1(n37371), .A2(n35457), .ZN(n37377) );
  AND3_X2 U344 ( .A1(n27878), .A2(n27879), .A3(n27877), .ZN(n27903) );
  NOR2_X2 U347 ( .A1(n45559), .A2(n48517), .ZN(n48512) );
  AND2_X2 U351 ( .A1(n48084), .A2(n48033), .ZN(n48020) );
  AND2_X2 U352 ( .A1(n41442), .A2(n41435), .ZN(n40643) );
  NAND2_X2 U353 ( .A1(n6869), .A2(n38565), .ZN(n38204) );
  OR2_X2 U354 ( .A1(n3189), .A2(n20641), .ZN(n20630) );
  AND4_X2 U361 ( .A1(n27606), .A2(n27611), .A3(n27612), .A4(n30672), .ZN(n3502) );
  AND2_X2 U364 ( .A1(n38259), .A2(n35305), .ZN(n37219) );
  NAND2_X2 U367 ( .A1(n3447), .A2(n1051), .ZN(n39077) );
  BUF_X4 U369 ( .A(n50338), .Z(n51725) );
  CLKBUF_X3 U370 ( .A(n31940), .Z(n51744) );
  AND2_X2 U371 ( .A1(n30924), .A2(n30930), .ZN(n31058) );
  NAND2_X2 U382 ( .A1(n48534), .A2(n48239), .ZN(n48551) );
  AND2_X2 U396 ( .A1(n4555), .A2(n11687), .ZN(n11673) );
  NAND2_X2 U397 ( .A1(n5385), .A2(n18380), .ZN(n20044) );
  NAND4_X2 U398 ( .A1(n23450), .A2(n23447), .A3(n23448), .A4(n23449), .ZN(
        n28288) );
  OR2_X2 U410 ( .A1(n43464), .A2(n43460), .ZN(n45987) );
  INV_X2 U411 ( .A(n6961), .ZN(n40003) );
  NAND4_X2 U422 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n17389) );
  BUF_X2 U429 ( .A(n45065), .Z(n47122) );
  BUF_X1 U431 ( .A(n26519), .Z(n52201) );
  INV_X2 U433 ( .A(n20903), .ZN(n23442) );
  BUF_X2 U436 ( .A(n30432), .Z(n51746) );
  XNOR2_X2 U437 ( .A(n17177), .B(n15896), .ZN(n16782) );
  NOR2_X2 U439 ( .A1(n48919), .A2(n48888), .ZN(n48911) );
  INV_X2 U441 ( .A(n18755), .ZN(n16498) );
  OR2_X2 U444 ( .A1(n38401), .A2(n40684), .ZN(n39931) );
  CLKBUF_X3 U447 ( .A(n15631), .Z(n51127) );
  OR2_X4 U458 ( .A1(n5189), .A2(n52358), .ZN(n17891) );
  OR2_X2 U462 ( .A1(n7990), .A2(n51868), .ZN(n40689) );
  XNOR2_X2 U463 ( .A(n28213), .B(n27291), .ZN(n24945) );
  AND2_X2 U468 ( .A1(n46691), .A2(n51513), .ZN(n46692) );
  NAND4_X2 U481 ( .A1(n29981), .A2(n29980), .A3(n29979), .A4(n29978), .ZN(
        n34361) );
  AND3_X2 U483 ( .A1(n281), .A2(n24576), .A3(n24574), .ZN(n31311) );
  AND2_X2 U484 ( .A1(n40295), .A2(n42062), .ZN(n40294) );
  NAND2_X2 U489 ( .A1(n12350), .A2(n805), .ZN(n8791) );
  BUF_X1 U491 ( .A(n33151), .Z(n51638) );
  BUF_X2 U494 ( .A(n21441), .Z(n52139) );
  INV_X2 U498 ( .A(n41004), .ZN(n40807) );
  BUF_X1 U499 ( .A(n20497), .Z(n52146) );
  INV_X2 U504 ( .A(n12756), .ZN(n14633) );
  BUF_X2 U505 ( .A(n28809), .Z(n52218) );
  BUF_X2 U514 ( .A(n47771), .Z(n52149) );
  NOR2_X2 U519 ( .A1(n17546), .A2(n18331), .ZN(n403) );
  AND2_X2 U523 ( .A1(n6486), .A2(n30265), .ZN(n29242) );
  NOR2_X2 U526 ( .A1(n8687), .A2(n51704), .ZN(n20508) );
  NOR2_X2 U527 ( .A1(n41110), .A2(n41268), .ZN(n41734) );
  XNOR2_X2 U529 ( .A(Key[110]), .B(Ciphertext[31]), .ZN(n52140) );
  INV_X2 U542 ( .A(n45189), .ZN(n46738) );
  XNOR2_X2 U551 ( .A(n4993), .B(n51850), .ZN(n37804) );
  AND2_X2 U555 ( .A1(n30665), .A2(n23861), .ZN(n27601) );
  OR2_X2 U558 ( .A1(n44800), .A2(n49127), .ZN(n49083) );
  AND2_X2 U567 ( .A1(n30696), .A2(n30389), .ZN(n30391) );
  OR2_X2 U569 ( .A1(n20805), .A2(n7835), .ZN(n21373) );
  NOR2_X2 U570 ( .A1(n14454), .A2(n14106), .ZN(n14450) );
  BUF_X2 U571 ( .A(n27210), .Z(n51751) );
  INV_X2 U572 ( .A(n49854), .ZN(n49863) );
  CLKBUF_X3 U576 ( .A(n49375), .Z(n51729) );
  AND2_X2 U577 ( .A1(n38514), .A2(n37437), .ZN(n38535) );
  XNOR2_X2 U580 ( .A(n45386), .B(n43219), .ZN(n44288) );
  NAND3_X2 U581 ( .A1(n1863), .A2(n1862), .A3(n52334), .ZN(n31995) );
  AND2_X2 U592 ( .A1(n3996), .A2(n8911), .ZN(n14984) );
  OR2_X2 U600 ( .A1(n2143), .A2(n51693), .ZN(n29000) );
  INV_X2 U602 ( .A(n41292), .ZN(n40417) );
  NAND4_X2 U610 ( .A1(n38858), .A2(n38857), .A3(n6713), .A4(n38856), .ZN(
        n51464) );
  AND2_X2 U611 ( .A1(n1085), .A2(n32716), .ZN(n32717) );
  AND2_X2 U629 ( .A1(n49242), .A2(n49397), .ZN(n49248) );
  OR2_X2 U630 ( .A1(n49521), .A2(n49511), .ZN(n49491) );
  AND2_X2 U643 ( .A1(n51093), .A2(n49983), .ZN(n47349) );
  XNOR2_X2 U647 ( .A(n40283), .B(n40282), .ZN(n43148) );
  OR3_X1 U652 ( .A1(n2895), .A2(n2421), .A3(n38632), .ZN(n38646) );
  OR2_X1 U654 ( .A1(n650), .A2(n48074), .ZN(n48069) );
  INV_X1 U665 ( .A(n28796), .ZN(n28970) );
  BUF_X1 U671 ( .A(n46830), .Z(n51456) );
  NAND4_X1 U672 ( .A1(n40977), .A2(n40978), .A3(n40976), .A4(n40975), .ZN(
        n52125) );
  INV_X1 U675 ( .A(n36575), .ZN(n4246) );
  INV_X1 U681 ( .A(n46356), .ZN(n46274) );
  OR2_X1 U688 ( .A1(n21425), .A2(n3493), .ZN(n19943) );
  AND4_X1 U712 ( .A1(n8523), .A2(n47090), .A3(n47092), .A4(n47091), .ZN(n47117) );
  OR2_X1 U715 ( .A1(n17584), .A2(n19336), .ZN(n17619) );
  INV_X1 U716 ( .A(n49782), .ZN(n49862) );
  NAND2_X1 U718 ( .A1(n36122), .A2(n35666), .ZN(n38584) );
  BUF_X1 U728 ( .A(n39813), .Z(n44431) );
  INV_X1 U732 ( .A(n37624), .ZN(n38279) );
  AND2_X1 U741 ( .A1(n31302), .A2(n31311), .ZN(n31298) );
  INV_X1 U745 ( .A(n27609), .ZN(n30665) );
  OR2_X1 U753 ( .A1(n21425), .A2(n19947), .ZN(n20327) );
  INV_X1 U762 ( .A(n49580), .ZN(n51088) );
  AND2_X1 U763 ( .A1(n10562), .A2(n11640), .ZN(n11649) );
  AOI22_X1 U765 ( .A1(n14652), .A2(n13434), .B1(n13439), .B2(n14656), .ZN(
        n12898) );
  INV_X1 U766 ( .A(n40269), .ZN(n40900) );
  BUF_X1 U768 ( .A(n11713), .Z(n51649) );
  AND2_X1 U773 ( .A1(n39290), .A2(n38731), .ZN(n38317) );
  XNOR2_X2 U776 ( .A(n52326), .B(n18526), .ZN(n21425) );
  NAND4_X2 U777 ( .A1(n16838), .A2(n16837), .A3(n16836), .A4(n16839), .ZN(
        n23481) );
  NAND3_X2 U779 ( .A1(n3408), .A2(n17207), .A3(n17205), .ZN(n52155) );
  NAND4_X2 U780 ( .A1(n22597), .A2(n22596), .A3(n22595), .A4(n22594), .ZN(
        n25775) );
  NAND4_X2 U784 ( .A1(n23839), .A2(n23836), .A3(n23838), .A4(n23837), .ZN(
        n28106) );
  XNOR2_X1 U796 ( .A(n6208), .B(n8498), .ZN(n26494) );
  AND3_X2 U798 ( .A1(n3109), .A2(n6622), .A3(n23162), .ZN(n52100) );
  NAND4_X2 U838 ( .A1(n29083), .A2(n29082), .A3(n29081), .A4(n29080), .ZN(
        n33759) );
  AND4_X2 U840 ( .A1(n38129), .A2(n38130), .A3(n38128), .A4(n38127), .ZN(
        n41375) );
  INV_X2 U841 ( .A(n41375), .ZN(n51853) );
  NAND3_X2 U845 ( .A1(n38711), .A2(n38713), .A3(n38712), .ZN(n40740) );
  INV_X2 U850 ( .A(n36509), .ZN(n39938) );
  NOR2_X2 U856 ( .A1(n6533), .A2(n37842), .ZN(n42863) );
  CLKBUF_X3 U866 ( .A(n44891), .Z(n51681) );
  NAND3_X2 U868 ( .A1(n36515), .A2(n36514), .A3(n4574), .ZN(n52096) );
  XNOR2_X2 U875 ( .A(n5362), .B(n6717), .ZN(n51344) );
  BUF_X2 U876 ( .A(n48698), .Z(n51659) );
  NAND2_X2 U877 ( .A1(n4348), .A2(n52415), .ZN(n48140) );
  NAND4_X2 U881 ( .A1(n31890), .A2(n31887), .A3(n31888), .A4(n31889), .ZN(
        n35543) );
  XNOR2_X2 U886 ( .A(n8247), .B(n33505), .ZN(n33562) );
  NAND4_X2 U893 ( .A1(n31248), .A2(n31246), .A3(n31247), .A4(n31245), .ZN(
        n34503) );
  BUF_X2 U904 ( .A(n7877), .Z(n396) );
  BUF_X1 U908 ( .A(n33151), .Z(n51639) );
  BUF_X1 U909 ( .A(n33151), .Z(n51640) );
  NAND4_X2 U910 ( .A1(n27972), .A2(n27922), .A3(n27921), .A4(n27923), .ZN(
        n32295) );
  AND4_X2 U912 ( .A1(n8314), .A2(n2718), .A3(n4221), .A4(n2717), .ZN(n13277)
         );
  BUF_X2 U913 ( .A(n17510), .Z(n21758) );
  CLKBUF_X1 U914 ( .A(n18547), .Z(n51641) );
  BUF_X2 U915 ( .A(n18547), .Z(n51642) );
  CLKBUF_X1 U920 ( .A(n50127), .Z(n51643) );
  BUF_X1 U924 ( .A(n50127), .Z(n51644) );
  BUF_X1 U925 ( .A(n50127), .Z(n51645) );
  XNOR2_X2 U934 ( .A(n34400), .B(n36681), .ZN(n34720) );
  OR2_X2 U938 ( .A1(n7750), .A2(n27978), .ZN(n36681) );
  OAI21_X2 U943 ( .B1(n36583), .B2(n36582), .A(n36581), .ZN(n36602) );
  CLKBUF_X1 U949 ( .A(n28416), .Z(n51646) );
  CLKBUF_X3 U955 ( .A(n28416), .Z(n51647) );
  NAND4_X1 U961 ( .A1(n23281), .A2(n23282), .A3(n23280), .A4(n23279), .ZN(
        n28416) );
  NAND4_X2 U965 ( .A1(n11309), .A2(n11308), .A3(n5584), .A4(n5580), .ZN(n18464) );
  BUF_X2 U966 ( .A(n28359), .Z(n51648) );
  NAND2_X1 U967 ( .A1(n36045), .A2(n36052), .ZN(n36595) );
  BUF_X2 U969 ( .A(n11713), .Z(n51650) );
  XNOR2_X1 U971 ( .A(n9138), .B(Key[71]), .ZN(n11713) );
  XNOR2_X1 U972 ( .A(n17821), .B(n51378), .ZN(n15876) );
  AND2_X1 U974 ( .A1(n29924), .A2(n27558), .ZN(n26842) );
  BUF_X2 U981 ( .A(n15396), .Z(n19198) );
  XNOR2_X2 U984 ( .A(n16743), .B(n18780), .ZN(n18181) );
  NAND2_X2 U986 ( .A1(n45186), .A2(n45188), .ZN(n46756) );
  CLKBUF_X1 U997 ( .A(n12505), .Z(n51652) );
  CLKBUF_X3 U1005 ( .A(n12505), .Z(n51653) );
  XNOR2_X1 U1015 ( .A(Key[95]), .B(Ciphertext[70]), .ZN(n12505) );
  CLKBUF_X3 U1017 ( .A(n23094), .Z(n51654) );
  BUF_X2 U1018 ( .A(n28127), .Z(n51121) );
  AND2_X2 U1020 ( .A1(n46305), .A2(n46304), .ZN(n52179) );
  CLKBUF_X3 U1031 ( .A(n47868), .Z(n51285) );
  CLKBUF_X1 U1040 ( .A(n13929), .Z(n51655) );
  BUF_X1 U1041 ( .A(n13929), .Z(n51656) );
  BUF_X1 U1045 ( .A(n13929), .Z(n51657) );
  NAND3_X1 U1048 ( .A1(n4427), .A2(n9816), .A3(n9817), .ZN(n13929) );
  BUF_X1 U1051 ( .A(n47403), .Z(n48714) );
  XNOR2_X2 U1053 ( .A(n52075), .B(n43973), .ZN(n44512) );
  OR2_X2 U1054 ( .A1(n18504), .A2(n18503), .ZN(n22605) );
  OR2_X2 U1070 ( .A1(n38057), .A2(n51522), .ZN(n38050) );
  CLKBUF_X1 U1075 ( .A(n48698), .Z(n51658) );
  AND2_X2 U1076 ( .A1(n8687), .A2(n51705), .ZN(n18086) );
  BUF_X1 U1088 ( .A(n15553), .Z(n51705) );
  XNOR2_X2 U1094 ( .A(n51329), .B(n44559), .ZN(n45304) );
  NAND2_X2 U1098 ( .A1(n39779), .A2(n39780), .ZN(n44559) );
  BUF_X2 U1102 ( .A(n29718), .Z(n51108) );
  INV_X1 U1104 ( .A(n27711), .ZN(n29424) );
  CLKBUF_X1 U1105 ( .A(n33607), .Z(n36960) );
  NAND2_X2 U1129 ( .A1(n29732), .A2(n29731), .ZN(n32732) );
  NAND4_X1 U1131 ( .A1(n17593), .A2(n6357), .A3(n17591), .A4(n17592), .ZN(
        n51660) );
  NAND4_X1 U1134 ( .A1(n17593), .A2(n6357), .A3(n17591), .A4(n17592), .ZN(
        n51661) );
  NAND4_X2 U1141 ( .A1(n17593), .A2(n6357), .A3(n17591), .A4(n17592), .ZN(
        n22157) );
  BUF_X1 U1150 ( .A(n34727), .Z(n51662) );
  BUF_X1 U1154 ( .A(n34727), .Z(n51663) );
  BUF_X1 U1166 ( .A(n34727), .Z(n51664) );
  XNOR2_X1 U1171 ( .A(n33195), .B(n36671), .ZN(n34727) );
  NAND2_X2 U1175 ( .A1(n886), .A2(n22773), .ZN(n7254) );
  XNOR2_X2 U1176 ( .A(n26579), .B(n26580), .ZN(n28882) );
  NAND2_X2 U1178 ( .A1(n4181), .A2(n4180), .ZN(n12914) );
  OR2_X2 U1179 ( .A1(n38969), .A2(n38970), .ZN(n41693) );
  INV_X2 U1186 ( .A(n41187), .ZN(n43168) );
  OAI211_X2 U1202 ( .C1(n32291), .C2(n32290), .A(n32289), .B(n32288), .ZN(
        n37292) );
  OAI211_X2 U1204 ( .C1(n43459), .C2(n43458), .A(n43457), .B(n2802), .ZN(n2193) );
  AND3_X2 U1218 ( .A1(n47351), .A2(n43454), .A3(n2803), .ZN(n2802) );
  CLKBUF_X1 U1222 ( .A(n28050), .Z(n51665) );
  CLKBUF_X1 U1225 ( .A(n28050), .Z(n51666) );
  BUF_X2 U1229 ( .A(n28050), .Z(n51667) );
  NAND4_X1 U1231 ( .A1(n20570), .A2(n5132), .A3(n5133), .A4(n20569), .ZN(
        n28050) );
  CLKBUF_X3 U1243 ( .A(n40951), .Z(n46642) );
  CLKBUF_X3 U1247 ( .A(n14687), .Z(n2151) );
  BUF_X2 U1259 ( .A(n17889), .Z(n51668) );
  XNOR2_X1 U1263 ( .A(n17764), .B(n7115), .ZN(n17889) );
  AND2_X2 U1264 ( .A1(n51480), .A2(n50192), .ZN(n50232) );
  NAND2_X2 U1273 ( .A1(n2886), .A2(n47345), .ZN(n50192) );
  XNOR2_X2 U1289 ( .A(n51249), .B(n35327), .ZN(n37667) );
  CLKBUF_X1 U1322 ( .A(n14702), .Z(n51669) );
  BUF_X1 U1337 ( .A(n14702), .Z(n51670) );
  CLKBUF_X1 U1345 ( .A(n14702), .Z(n51671) );
  NAND4_X1 U1346 ( .A1(n12274), .A2(n12273), .A3(n12275), .A4(n12272), .ZN(
        n14702) );
  BUF_X2 U1348 ( .A(n31573), .Z(n37252) );
  OAI21_X2 U1352 ( .B1(n27157), .B2(n27156), .A(n27155), .ZN(n31573) );
  XNOR2_X2 U1353 ( .A(n1513), .B(n7722), .ZN(n7721) );
  BUF_X1 U1354 ( .A(n12534), .Z(n51673) );
  BUF_X1 U1355 ( .A(n12534), .Z(n51674) );
  XNOR2_X2 U1357 ( .A(n33818), .B(n35835), .ZN(n33335) );
  NAND4_X2 U1360 ( .A1(n31617), .A2(n31616), .A3(n31615), .A4(n31614), .ZN(
        n33818) );
  INV_X1 U1369 ( .A(n17546), .ZN(n17542) );
  INV_X1 U1373 ( .A(n13874), .ZN(n14871) );
  NAND3_X2 U1382 ( .A1(n8653), .A2(n9252), .A3(n8651), .ZN(n13874) );
  XNOR2_X2 U1387 ( .A(n42173), .B(n42174), .ZN(n44640) );
  OR2_X2 U1388 ( .A1(n52263), .A2(n5944), .ZN(n32463) );
  AND2_X2 U1389 ( .A1(n49263), .A2(n52079), .ZN(n49273) );
  XNOR2_X2 U1399 ( .A(n42392), .B(n42391), .ZN(n49263) );
  CLKBUF_X1 U1411 ( .A(n23564), .Z(n51675) );
  BUF_X2 U1433 ( .A(n23564), .Z(n51677) );
  NAND2_X1 U1435 ( .A1(n1265), .A2(n17063), .ZN(n23564) );
  CLKBUF_X1 U1437 ( .A(n29421), .Z(n51678) );
  BUF_X1 U1442 ( .A(n29421), .Z(n51679) );
  XNOR2_X1 U1456 ( .A(n24624), .B(n24803), .ZN(n29421) );
  NAND2_X1 U1457 ( .A1(n2677), .A2(n27652), .ZN(n27671) );
  CLKBUF_X1 U1467 ( .A(n44891), .Z(n51680) );
  NAND2_X1 U1469 ( .A1(n3389), .A2(n6211), .ZN(n44891) );
  NOR2_X1 U1475 ( .A1(n39011), .A2(n3973), .ZN(n39025) );
  AND2_X2 U1489 ( .A1(n51991), .A2(n23875), .ZN(n25708) );
  XNOR2_X2 U1495 ( .A(n45323), .B(n45322), .ZN(n46464) );
  CLKBUF_X1 U1500 ( .A(n13520), .Z(n51682) );
  CLKBUF_X3 U1501 ( .A(n13520), .Z(n51683) );
  NAND4_X1 U1510 ( .A1(n3077), .A2(n3078), .A3(n8329), .A4(n9315), .ZN(n13520)
         );
  INV_X1 U1531 ( .A(n15259), .ZN(n51685) );
  INV_X1 U1532 ( .A(n15259), .ZN(n51686) );
  INV_X1 U1533 ( .A(n15259), .ZN(n15264) );
  AND2_X2 U1554 ( .A1(n2096), .A2(n2097), .ZN(n26100) );
  INV_X2 U1558 ( .A(n41646), .ZN(n40617) );
  OR2_X2 U1563 ( .A1(n7118), .A2(n2325), .ZN(n52101) );
  XNOR2_X2 U1580 ( .A(n41758), .B(n42715), .ZN(n45490) );
  NAND2_X2 U1585 ( .A1(n1457), .A2(n8288), .ZN(n13780) );
  XNOR2_X2 U1587 ( .A(n9287), .B(Key[108]), .ZN(n10068) );
  NAND2_X1 U1588 ( .A1(n489), .A2(n17584), .ZN(n20512) );
  XNOR2_X1 U1589 ( .A(n52308), .B(n15803), .ZN(n20656) );
  AND2_X2 U1606 ( .A1(n47037), .A2(n47038), .ZN(n50521) );
  OR4_X1 U1611 ( .A1(n36233), .A2(n37591), .A3(n37372), .A4(n36232), .ZN(
        n37367) );
  OR2_X2 U1627 ( .A1(n29439), .A2(n29442), .ZN(n26722) );
  NAND2_X1 U1637 ( .A1(n747), .A2(n29439), .ZN(n27830) );
  NOR2_X1 U1643 ( .A1(n44752), .A2(n45966), .ZN(n46232) );
  XNOR2_X2 U1644 ( .A(Key[52]), .B(Ciphertext[105]), .ZN(n10562) );
  XNOR2_X2 U1645 ( .A(n33777), .B(n2304), .ZN(n35457) );
  NOR2_X2 U1649 ( .A1(n4057), .A2(n39287), .ZN(n39316) );
  CLKBUF_X1 U1663 ( .A(n48904), .Z(n51687) );
  CLKBUF_X1 U1665 ( .A(n48904), .Z(n51689) );
  NAND4_X1 U1666 ( .A1(n45639), .A2(n45637), .A3(n48242), .A4(n45638), .ZN(
        n48904) );
  XNOR2_X2 U1676 ( .A(n15601), .B(n15600), .ZN(n15630) );
  NAND2_X2 U1688 ( .A1(n5605), .A2(n5608), .ZN(n41796) );
  CLKBUF_X1 U1689 ( .A(n50300), .Z(n51690) );
  CLKBUF_X3 U1690 ( .A(n50300), .Z(n51691) );
  XNOR2_X1 U1698 ( .A(n43085), .B(n43084), .ZN(n50300) );
  NAND4_X2 U1701 ( .A1(n6001), .A2(n6002), .A3(n23475), .A4(n23476), .ZN(
        n28238) );
  XNOR2_X2 U1703 ( .A(n18831), .B(n19186), .ZN(n16176) );
  AND2_X2 U1704 ( .A1(n28772), .A2(n29782), .ZN(n30375) );
  AND2_X2 U1705 ( .A1(n52181), .A2(n29782), .ZN(n30734) );
  XNOR2_X2 U1706 ( .A(n27332), .B(n27331), .ZN(n29782) );
  BUF_X1 U1709 ( .A(n30455), .Z(n51692) );
  BUF_X2 U1716 ( .A(n30455), .Z(n51693) );
  XNOR2_X1 U1721 ( .A(n28421), .B(n28422), .ZN(n30455) );
  NAND2_X2 U1724 ( .A1(n8741), .A2(n32582), .ZN(n33145) );
  INV_X1 U1728 ( .A(n21122), .ZN(n51694) );
  INV_X1 U1732 ( .A(n21122), .ZN(n51695) );
  BUF_X1 U1745 ( .A(n30754), .Z(n51696) );
  CLKBUF_X1 U1750 ( .A(n30754), .Z(n51697) );
  BUF_X2 U1759 ( .A(n51062), .Z(n51063) );
  XNOR2_X2 U1761 ( .A(n28106), .B(n26090), .ZN(n26393) );
  OR2_X2 U1775 ( .A1(n23819), .A2(n23820), .ZN(n26090) );
  CLKBUF_X1 U1781 ( .A(n15337), .Z(n51698) );
  BUF_X1 U1796 ( .A(n15337), .Z(n51699) );
  BUF_X1 U1806 ( .A(n15337), .Z(n51700) );
  BUF_X2 U1816 ( .A(n34392), .Z(n51702) );
  AND2_X2 U1825 ( .A1(n1061), .A2(n1062), .ZN(n2690) );
  AND4_X2 U1826 ( .A1(n4458), .A2(n2493), .A3(n4457), .A4(n3186), .ZN(n23414)
         );
  XNOR2_X2 U1827 ( .A(n43761), .B(n43762), .ZN(n50364) );
  BUF_X2 U1845 ( .A(n50343), .Z(n51386) );
  BUF_X1 U1854 ( .A(n15553), .Z(n51704) );
  XNOR2_X1 U1858 ( .A(n15477), .B(n779), .ZN(n15553) );
  NAND4_X2 U1866 ( .A1(n11181), .A2(n1844), .A3(n11180), .A4(n11182), .ZN(
        n19260) );
  NAND2_X2 U1867 ( .A1(n3420), .A2(n26799), .ZN(n35589) );
  NAND3_X2 U1868 ( .A1(n35429), .A2(n35432), .A3(n5987), .ZN(n39101) );
  NAND2_X2 U1877 ( .A1(n1090), .A2(n1091), .ZN(n16039) );
  OAI21_X2 U1879 ( .B1(n24259), .B2(n24258), .A(n24257), .ZN(n26547) );
  AND2_X2 U1886 ( .A1(n5619), .A2(n5620), .ZN(n15163) );
  OR2_X1 U1893 ( .A1(n15553), .A2(n20501), .ZN(n17627) );
  XNOR2_X2 U1900 ( .A(n45382), .B(n44208), .ZN(n42067) );
  BUF_X2 U1909 ( .A(n31040), .Z(n50986) );
  XNOR2_X2 U1913 ( .A(Key[154]), .B(Ciphertext[147]), .ZN(n10199) );
  XNOR2_X2 U1914 ( .A(n44373), .B(n51323), .ZN(n7387) );
  AND2_X2 U1916 ( .A1(n12128), .A2(n12127), .ZN(n14533) );
  XNOR2_X2 U1931 ( .A(n18635), .B(n18634), .ZN(n21354) );
  CLKBUF_X1 U1933 ( .A(n11543), .Z(n51708) );
  XNOR2_X1 U1939 ( .A(n8638), .B(Key[81]), .ZN(n11543) );
  AND3_X2 U1943 ( .A1(n3721), .A2(n3720), .A3(n3726), .ZN(n32725) );
  XNOR2_X2 U1949 ( .A(n8866), .B(Key[114]), .ZN(n11485) );
  OR2_X2 U1956 ( .A1(n36072), .A2(n36071), .ZN(n584) );
  NAND4_X2 U1957 ( .A1(n4134), .A2(n29100), .A3(n29098), .A4(n29099), .ZN(
        n37065) );
  OR2_X2 U1964 ( .A1(n18040), .A2(n15398), .ZN(n18032) );
  XNOR2_X2 U1984 ( .A(n15397), .B(n5672), .ZN(n18040) );
  BUF_X2 U2001 ( .A(n40686), .Z(n39929) );
  BUF_X2 U2002 ( .A(n21579), .Z(n51710) );
  CLKBUF_X1 U2006 ( .A(n21579), .Z(n51711) );
  XNOR2_X1 U2007 ( .A(n18839), .B(n18838), .ZN(n21579) );
  OAI211_X2 U2011 ( .C1(n20927), .C2(n20926), .A(n20925), .B(n20924), .ZN(
        n27424) );
  XNOR2_X2 U2016 ( .A(n18201), .B(n18200), .ZN(n18888) );
  AND2_X2 U2026 ( .A1(n39410), .A2(n37901), .ZN(n39426) );
  XNOR2_X2 U2027 ( .A(n36799), .B(n36798), .ZN(n39410) );
  BUF_X1 U2035 ( .A(n13378), .Z(n51712) );
  BUF_X1 U2041 ( .A(n13378), .Z(n51713) );
  BUF_X1 U2043 ( .A(n13378), .Z(n51714) );
  CLKBUF_X1 U2044 ( .A(n36621), .Z(n51715) );
  BUF_X2 U2046 ( .A(n36621), .Z(n51716) );
  CLKBUF_X1 U2047 ( .A(n36621), .Z(n51717) );
  XNOR2_X1 U2052 ( .A(n34230), .B(n34231), .ZN(n36621) );
  XNOR2_X2 U2058 ( .A(n9097), .B(Key[76]), .ZN(n9104) );
  AND2_X2 U2061 ( .A1(n15399), .A2(n18041), .ZN(n19404) );
  CLKBUF_X1 U2064 ( .A(n25770), .Z(n51719) );
  NOR2_X2 U2068 ( .A1(n1414), .A2(n1417), .ZN(n18352) );
  CLKBUF_X1 U2069 ( .A(n5714), .Z(n51721) );
  CLKBUF_X1 U2071 ( .A(n5714), .Z(n51722) );
  BUF_X1 U2072 ( .A(n5714), .Z(n51723) );
  BUF_X2 U2073 ( .A(n15275), .Z(n51724) );
  INV_X1 U2074 ( .A(n48769), .ZN(n48729) );
  INV_X1 U2075 ( .A(n46173), .ZN(n49933) );
  BUF_X1 U2089 ( .A(n46542), .Z(n48155) );
  BUF_X2 U2090 ( .A(n50784), .Z(n51730) );
  NAND2_X2 U2093 ( .A1(n49978), .A2(n2790), .ZN(n49987) );
  INV_X1 U2106 ( .A(n46203), .ZN(n49278) );
  INV_X2 U2111 ( .A(n45597), .ZN(n48478) );
  BUF_X1 U2114 ( .A(n49662), .Z(n51733) );
  BUF_X2 U2115 ( .A(n44206), .Z(n48517) );
  BUF_X1 U2117 ( .A(n49276), .Z(n52086) );
  INV_X2 U2135 ( .A(n41054), .ZN(n41057) );
  AND4_X1 U2138 ( .A1(n38654), .A2(n38655), .A3(n38657), .A4(n38656), .ZN(
        n41356) );
  NAND2_X2 U2139 ( .A1(n1075), .A2(n7159), .ZN(n36216) );
  INV_X1 U2140 ( .A(n36200), .ZN(n37778) );
  INV_X1 U2152 ( .A(n38561), .ZN(n38201) );
  CLKBUF_X2 U2164 ( .A(n38084), .Z(n50984) );
  INV_X1 U2165 ( .A(n38547), .ZN(n31355) );
  INV_X1 U2166 ( .A(n36473), .ZN(n36493) );
  BUF_X1 U2173 ( .A(n35768), .Z(n52071) );
  INV_X1 U2174 ( .A(n29211), .ZN(n32080) );
  BUF_X1 U2179 ( .A(n31377), .Z(n51740) );
  INV_X2 U2181 ( .A(n31398), .ZN(n32829) );
  NAND3_X1 U2200 ( .A1(n25846), .A2(n2442), .A3(n25845), .ZN(n52047) );
  INV_X2 U2204 ( .A(n31821), .ZN(n31826) );
  INV_X2 U2211 ( .A(n32345), .ZN(n723) );
  AND2_X1 U2217 ( .A1(n5417), .A2(n29147), .ZN(n29153) );
  NAND2_X2 U2219 ( .A1(n28666), .A2(n6346), .ZN(n26677) );
  NAND2_X1 U2226 ( .A1(n5522), .A2(n29192), .ZN(n29269) );
  BUF_X1 U2232 ( .A(n7614), .Z(n51748) );
  BUF_X1 U2243 ( .A(n26306), .Z(n51747) );
  INV_X1 U2246 ( .A(n29159), .ZN(n51726) );
  BUF_X2 U2250 ( .A(n28358), .Z(n51749) );
  INV_X1 U2251 ( .A(n22434), .ZN(n22982) );
  INV_X1 U2263 ( .A(n23955), .ZN(n23638) );
  NAND2_X1 U2270 ( .A1(n23483), .A2(n21981), .ZN(n21991) );
  INV_X2 U2274 ( .A(n23135), .ZN(n23906) );
  INV_X2 U2276 ( .A(n24412), .ZN(n24117) );
  BUF_X1 U2277 ( .A(n23810), .Z(n51753) );
  INV_X1 U2278 ( .A(n22184), .ZN(n5683) );
  INV_X2 U2282 ( .A(n22856), .ZN(n23021) );
  INV_X2 U2285 ( .A(n22861), .ZN(n22849) );
  NAND2_X2 U2300 ( .A1(n6929), .A2(n20623), .ZN(n20197) );
  INV_X2 U2311 ( .A(n19777), .ZN(n21269) );
  BUF_X1 U2312 ( .A(n21303), .Z(n509) );
  BUF_X1 U2314 ( .A(n15723), .Z(n19685) );
  INV_X1 U2329 ( .A(n20232), .ZN(n1597) );
  CLKBUF_X1 U2332 ( .A(n20613), .Z(n52213) );
  INV_X2 U2334 ( .A(n14542), .ZN(n14536) );
  INV_X1 U2335 ( .A(n14285), .ZN(n5411) );
  INV_X1 U2336 ( .A(n14164), .ZN(n51175) );
  INV_X1 U2339 ( .A(n14103), .ZN(n14107) );
  NAND3_X1 U2341 ( .A1(n52291), .A2(n9106), .A3(n7485), .ZN(n12755) );
  NAND2_X2 U2344 ( .A1(n9499), .A2(n9495), .ZN(n11697) );
  INV_X2 U2351 ( .A(n12161), .ZN(n12173) );
  INV_X2 U2352 ( .A(n9895), .ZN(n9083) );
  AND2_X1 U2364 ( .A1(n48754), .A2(n48753), .ZN(n51865) );
  AND4_X1 U2365 ( .A1(n5148), .A2(n45880), .A3(n2451), .A4(n45878), .ZN(n52029) );
  OR2_X1 U2373 ( .A1(n46421), .A2(n994), .ZN(n48786) );
  NOR2_X1 U2374 ( .A1(n47234), .A2(n51388), .ZN(n50938) );
  NOR2_X1 U2375 ( .A1(n46936), .A2(n49025), .ZN(n52258) );
  AND3_X1 U2379 ( .A1(n2635), .A2(n48877), .A3(n2636), .ZN(n45707) );
  AOI22_X1 U2380 ( .A1(n50633), .A2(n51994), .B1(n44124), .B2(n50588), .ZN(
        n44128) );
  AND2_X1 U2385 ( .A1(n50429), .A2(n50435), .ZN(n52015) );
  NOR2_X1 U2389 ( .A1(n50906), .A2(n50950), .ZN(n47396) );
  BUF_X2 U2390 ( .A(n46279), .Z(n51310) );
  AND2_X1 U2397 ( .A1(n48729), .A2(n48747), .ZN(n48749) );
  OR2_X1 U2398 ( .A1(n49579), .A2(n49569), .ZN(n49605) );
  BUF_X2 U2402 ( .A(n7459), .Z(n50705) );
  BUF_X1 U2413 ( .A(n45886), .Z(n47698) );
  INV_X1 U2426 ( .A(n50143), .ZN(n51727) );
  NOR2_X1 U2430 ( .A1(n46237), .A2(n46238), .ZN(n46279) );
  BUF_X2 U2438 ( .A(n48391), .Z(n51728) );
  OR2_X1 U2444 ( .A1(n46647), .A2(n46646), .ZN(n51340) );
  AND4_X1 U2446 ( .A1(n46887), .A2(n46886), .A3(n46885), .A4(n46884), .ZN(
        n52093) );
  NAND3_X1 U2450 ( .A1(n46761), .A2(n1233), .A3(n46764), .ZN(n47570) );
  NAND2_X1 U2460 ( .A1(n47194), .A2(n47193), .ZN(n47195) );
  AND4_X1 U2463 ( .A1(n7167), .A2(n43449), .A3(n6126), .A4(n43450), .ZN(n6125)
         );
  INV_X1 U2472 ( .A(n48604), .ZN(n48649) );
  NAND2_X1 U2476 ( .A1(n1662), .A2(n52393), .ZN(n47937) );
  AND3_X2 U2490 ( .A1(n5814), .A2(n7300), .A3(n7301), .ZN(n49580) );
  OR2_X1 U2491 ( .A1(n51229), .A2(n52287), .ZN(n48747) );
  AND2_X1 U2496 ( .A1(n45556), .A2(n5320), .ZN(n51881) );
  AND2_X1 U2509 ( .A1(n47403), .A2(n48697), .ZN(n47407) );
  NOR2_X1 U2512 ( .A1(n1339), .A2(n50025), .ZN(n47194) );
  NAND4_X1 U2518 ( .A1(n45956), .A2(n45955), .A3(n45954), .A4(n45953), .ZN(
        n52107) );
  NAND3_X1 U2527 ( .A1(n46718), .A2(n5410), .A3(n7127), .ZN(n51289) );
  AND4_X1 U2528 ( .A1(n8628), .A2(n47148), .A3(n47147), .A4(n8668), .ZN(n51296) );
  AND3_X1 U2533 ( .A1(n48495), .A2(n48496), .A3(n48494), .ZN(n52042) );
  AND3_X1 U2536 ( .A1(n5171), .A2(n47131), .A3(n47130), .ZN(n6251) );
  NOR2_X1 U2539 ( .A1(n45941), .A2(n45940), .ZN(n45956) );
  OR2_X1 U2540 ( .A1(n49955), .A2(n51691), .ZN(n27) );
  INV_X1 U2543 ( .A(n49233), .ZN(n51731) );
  OR2_X1 U2544 ( .A1(n46376), .A2(n48233), .ZN(n51997) );
  AND2_X1 U2547 ( .A1(n46901), .A2(n46905), .ZN(n46607) );
  INV_X1 U2548 ( .A(n52003), .ZN(n48507) );
  INV_X1 U2550 ( .A(n49148), .ZN(n46299) );
  OAI21_X1 U2551 ( .B1(n7110), .B2(n46471), .A(n48196), .ZN(n52003) );
  CLKBUF_X1 U2554 ( .A(n45231), .Z(n52187) );
  INV_X2 U2558 ( .A(n43479), .ZN(n49242) );
  AND2_X1 U2565 ( .A1(n7426), .A2(n43797), .ZN(n47139) );
  INV_X1 U2570 ( .A(n46492), .ZN(n46502) );
  NOR2_X1 U2581 ( .A1(n6132), .A2(n50280), .ZN(n50251) );
  AND2_X1 U2585 ( .A1(n46709), .A2(n46708), .ZN(n46575) );
  OR2_X1 U2592 ( .A1(n48456), .A2(n42508), .ZN(n48455) );
  XNOR2_X1 U2604 ( .A(n43934), .B(n41186), .ZN(n45790) );
  BUF_X2 U2605 ( .A(n50317), .Z(n52224) );
  OR2_X1 U2630 ( .A1(n46565), .A2(n46721), .ZN(n47111) );
  NOR2_X1 U2637 ( .A1(n663), .A2(n47152), .ZN(n45165) );
  XNOR2_X1 U2656 ( .A(n41842), .B(n41841), .ZN(n44992) );
  BUF_X1 U2661 ( .A(n48201), .Z(n52070) );
  BUF_X2 U2662 ( .A(n48462), .Z(n51732) );
  INV_X1 U2668 ( .A(n46888), .ZN(n663) );
  XNOR2_X1 U2672 ( .A(n43602), .B(n45344), .ZN(n47152) );
  INV_X2 U2685 ( .A(n49170), .ZN(n49161) );
  BUF_X1 U2689 ( .A(n46463), .Z(n2207) );
  BUF_X1 U2691 ( .A(n46197), .Z(n52079) );
  XNOR2_X1 U2697 ( .A(n41871), .B(n41870), .ZN(n48213) );
  XNOR2_X1 U2714 ( .A(n42280), .B(n43812), .ZN(n42487) );
  BUF_X1 U2740 ( .A(n43638), .Z(n45299) );
  CLKBUF_X1 U2748 ( .A(n43740), .Z(n52084) );
  CLKBUF_X1 U2754 ( .A(n45101), .Z(n607) );
  NAND4_X2 U2755 ( .A1(n1237), .A2(n41386), .A3(n41384), .A4(n41385), .ZN(
        n45355) );
  NAND4_X1 U2764 ( .A1(n39688), .A2(n39687), .A3(n39686), .A4(n39685), .ZN(
        n43014) );
  OAI21_X1 U2769 ( .B1(n51847), .B2(n40664), .A(n41207), .ZN(n41220) );
  NOR2_X1 U2772 ( .A1(n4040), .A2(n40965), .ZN(n40977) );
  AND2_X1 U2779 ( .A1(n39129), .A2(n40493), .ZN(n52357) );
  AND2_X1 U2788 ( .A1(n41535), .A2(n40938), .ZN(n41526) );
  NOR2_X1 U2795 ( .A1(n39908), .A2(n39907), .ZN(n39918) );
  AND2_X1 U2805 ( .A1(n41049), .A2(n40502), .ZN(n40499) );
  AND2_X1 U2811 ( .A1(n8500), .A2(n7818), .ZN(n40049) );
  AND2_X1 U2815 ( .A1(n40341), .A2(n40327), .ZN(n39853) );
  NOR2_X1 U2820 ( .A1(n38782), .A2(n40110), .ZN(n40192) );
  INV_X1 U2847 ( .A(n38810), .ZN(n51734) );
  NAND4_X1 U2856 ( .A1(n812), .A2(n37676), .A3(n37674), .A4(n37675), .ZN(
        n52151) );
  AND2_X1 U2858 ( .A1(n6451), .A2(n51918), .ZN(n6450) );
  NAND2_X1 U2863 ( .A1(n35570), .A2(n7847), .ZN(n40565) );
  NAND3_X1 U2879 ( .A1(n1864), .A2(n6552), .A3(n2272), .ZN(n52083) );
  OR2_X1 U2883 ( .A1(n35428), .A2(n35427), .ZN(n6961) );
  AND3_X1 U3020 ( .A1(n5397), .A2(n5396), .A3(n51952), .ZN(n1196) );
  AND2_X1 U3051 ( .A1(n38223), .A2(n2720), .ZN(n52329) );
  AOI21_X1 U3062 ( .B1(n51810), .B2(n37884), .A(n51809), .ZN(n39405) );
  OAI21_X1 U3066 ( .B1(n36583), .B2(n36453), .A(n36458), .ZN(n36466) );
  AND3_X1 U3069 ( .A1(n38254), .A2(n5990), .A3(n38253), .ZN(n38269) );
  AND2_X1 U3086 ( .A1(n39397), .A2(n39003), .ZN(n51810) );
  OR2_X1 U3098 ( .A1(n38512), .A2(n35530), .ZN(n35960) );
  OR2_X1 U3113 ( .A1(n36233), .A2(n52372), .ZN(n36234) );
  OR2_X1 U3121 ( .A1(n36225), .A2(n35452), .ZN(n35971) );
  AND2_X1 U3125 ( .A1(n35458), .A2(n37378), .ZN(n35980) );
  INV_X1 U3126 ( .A(n38962), .ZN(n51872) );
  AND2_X1 U3128 ( .A1(n38962), .A2(n37790), .ZN(n39361) );
  NOR2_X1 U3133 ( .A1(n6367), .A2(n35010), .ZN(n36325) );
  AND2_X1 U3136 ( .A1(n37420), .A2(n38475), .ZN(n38116) );
  INV_X1 U3142 ( .A(n38529), .ZN(n51735) );
  AND2_X1 U3144 ( .A1(n33456), .A2(n35939), .ZN(n37780) );
  NOR2_X1 U3153 ( .A1(n35939), .A2(n36196), .ZN(n39335) );
  NAND2_X1 U3163 ( .A1(n39429), .A2(n38937), .ZN(n38949) );
  BUF_X1 U3172 ( .A(n34084), .Z(n36541) );
  INV_X1 U3183 ( .A(n39235), .ZN(n51736) );
  XNOR2_X1 U3186 ( .A(n35138), .B(n35137), .ZN(n37420) );
  AND2_X2 U3189 ( .A1(n36299), .A2(n31358), .ZN(n38550) );
  NOR2_X1 U3194 ( .A1(n36473), .A2(n51874), .ZN(n51873) );
  BUF_X2 U3211 ( .A(n37721), .Z(n51737) );
  XNOR2_X1 U3237 ( .A(n35349), .B(n35348), .ZN(n35405) );
  INV_X1 U3238 ( .A(n36299), .ZN(n51738) );
  XNOR2_X1 U3257 ( .A(n51942), .B(n33868), .ZN(n2176) );
  INV_X1 U3265 ( .A(n702), .ZN(n36992) );
  NAND2_X1 U3268 ( .A1(n51882), .A2(n31072), .ZN(n33938) );
  BUF_X2 U3274 ( .A(n37112), .Z(n51739) );
  NAND2_X1 U3275 ( .A1(n52412), .A2(n52411), .ZN(n36758) );
  NOR2_X1 U3277 ( .A1(n32624), .A2(n32625), .ZN(n702) );
  NAND4_X1 U3289 ( .A1(n31672), .A2(n31673), .A3(n31667), .A4(n51564), .ZN(
        n34605) );
  NAND4_X1 U3291 ( .A1(n30548), .A2(n30547), .A3(n30546), .A4(n30545), .ZN(
        n51427) );
  OR2_X1 U3294 ( .A1(n31776), .A2(n31775), .ZN(n52411) );
  NAND4_X1 U3304 ( .A1(n52278), .A2(n29948), .A3(n1762), .A4(n1761), .ZN(
        n33806) );
  AND3_X1 U3321 ( .A1(n32167), .A2(n32168), .A3(n32169), .ZN(n52241) );
  AND2_X1 U3324 ( .A1(n32469), .A2(n51840), .ZN(n52262) );
  AOI22_X1 U3326 ( .A1(n1701), .A2(n29104), .B1(n1702), .B2(n29103), .ZN(n1700) );
  NOR2_X1 U3332 ( .A1(n31885), .A2(n31797), .ZN(n1823) );
  AND2_X1 U3350 ( .A1(n6157), .A2(n32609), .ZN(n32614) );
  INV_X1 U3352 ( .A(n31553), .ZN(n31159) );
  AOI21_X1 U3367 ( .B1(n32358), .B2(n32359), .A(n32357), .ZN(n32362) );
  OR2_X1 U3377 ( .A1(n7626), .A2(n51106), .ZN(n31155) );
  AND2_X1 U3398 ( .A1(n3754), .A2(n32175), .ZN(n32967) );
  NOR2_X1 U3404 ( .A1(n31638), .A2(n30855), .ZN(n31632) );
  OR2_X1 U3429 ( .A1(n31546), .A2(n382), .ZN(n2699) );
  OR2_X1 U3451 ( .A1(n32830), .A2(n32815), .ZN(n32426) );
  NOR2_X1 U3456 ( .A1(n30861), .A2(n51545), .ZN(n31626) );
  AND2_X1 U3459 ( .A1(n32057), .A2(n32056), .ZN(n32360) );
  OR2_X1 U3467 ( .A1(n30872), .A2(n30873), .ZN(n29675) );
  AND2_X1 U3472 ( .A1(n32882), .A2(n32879), .ZN(n32887) );
  NOR2_X1 U3486 ( .A1(n3099), .A2(n30925), .ZN(n31519) );
  OR2_X1 U3498 ( .A1(n28515), .A2(n28516), .ZN(n32701) );
  AND3_X2 U3507 ( .A1(n52250), .A2(n52249), .A3(n28968), .ZN(n32883) );
  AND3_X1 U3512 ( .A1(n28845), .A2(n28844), .A3(n28846), .ZN(n51822) );
  OR2_X2 U3522 ( .A1(n8272), .A2(n8361), .ZN(n32486) );
  NOR2_X1 U3526 ( .A1(n32761), .A2(n32960), .ZN(n32956) );
  OR2_X1 U3539 ( .A1(n28515), .A2(n28516), .ZN(n52182) );
  INV_X1 U3544 ( .A(n32795), .ZN(n32286) );
  INV_X1 U3545 ( .A(n30073), .ZN(n51742) );
  INV_X1 U3550 ( .A(n31873), .ZN(n51743) );
  OR2_X1 U3551 ( .A1(n32785), .A2(n32784), .ZN(n32795) );
  AND3_X1 U3557 ( .A1(n28665), .A2(n2458), .A3(n7573), .ZN(n7392) );
  AND2_X1 U3561 ( .A1(n27117), .A2(n27118), .ZN(n52334) );
  AND3_X1 U3563 ( .A1(n27028), .A2(n27027), .A3(n51910), .ZN(n27046) );
  AOI21_X1 U3566 ( .B1(n28152), .B2(n51842), .A(n51767), .ZN(n6524) );
  AND3_X1 U3582 ( .A1(n25978), .A2(n25970), .A3(n25977), .ZN(n6877) );
  AND2_X1 U3583 ( .A1(n28197), .A2(n28196), .ZN(n52370) );
  AND2_X1 U3586 ( .A1(n29219), .A2(n27916), .ZN(n51974) );
  NOR2_X1 U3589 ( .A1(n29342), .A2(n29204), .ZN(n30208) );
  OR2_X1 U3640 ( .A1(n27030), .A2(n27029), .ZN(n51910) );
  OR2_X1 U3657 ( .A1(n29248), .A2(n29263), .ZN(n52023) );
  AND2_X1 U3659 ( .A1(n28860), .A2(n2707), .ZN(n28508) );
  AND2_X1 U3661 ( .A1(n28669), .A2(n26668), .ZN(n27859) );
  AND2_X1 U3665 ( .A1(n29747), .A2(n29749), .ZN(n30452) );
  INV_X1 U3667 ( .A(n29068), .ZN(n29760) );
  BUF_X2 U3672 ( .A(n28638), .Z(n51107) );
  NAND2_X2 U3675 ( .A1(n1484), .A2(n26954), .ZN(n27685) );
  BUF_X1 U3688 ( .A(n26455), .Z(n29007) );
  OR2_X1 U3695 ( .A1(n30209), .A2(n29343), .ZN(n29200) );
  XNOR2_X1 U3701 ( .A(n23653), .B(n23654), .ZN(n5714) );
  XNOR2_X1 U3707 ( .A(n51927), .B(n25819), .ZN(n27860) );
  CLKBUF_X1 U3710 ( .A(n26552), .Z(n52163) );
  OAI211_X1 U3715 ( .C1(n4847), .C2(n23007), .A(n23011), .B(n51787), .ZN(
        n26548) );
  XNOR2_X1 U3732 ( .A(n3110), .B(n24403), .ZN(n25816) );
  BUF_X2 U3739 ( .A(n26607), .Z(n51750) );
  OR3_X2 U3750 ( .A1(n23699), .A2(n7215), .A3(n7214), .ZN(n25724) );
  AND3_X1 U3760 ( .A1(n23010), .A2(n23008), .A3(n23332), .ZN(n23007) );
  NAND3_X1 U3773 ( .A1(n21966), .A2(n4619), .A3(n21965), .ZN(n2080) );
  OAI211_X1 U3777 ( .C1(n22324), .C2(n22323), .A(n22322), .B(n22321), .ZN(
        n25770) );
  BUF_X2 U3808 ( .A(n26519), .Z(n51752) );
  AND2_X1 U3816 ( .A1(n22094), .A2(n51901), .ZN(n51900) );
  OR2_X1 U3821 ( .A1(n2025), .A2(n23595), .ZN(n23594) );
  NOR2_X1 U3822 ( .A1(n23294), .A2(n23095), .ZN(n51923) );
  AND2_X1 U3825 ( .A1(n23029), .A2(n24001), .ZN(n23036) );
  AND2_X1 U3856 ( .A1(n23539), .A2(n23703), .ZN(n52310) );
  INV_X1 U3871 ( .A(n1024), .ZN(n51832) );
  OR2_X1 U3873 ( .A1(n22320), .A2(n23411), .ZN(n22033) );
  CLKBUF_X1 U3878 ( .A(n20876), .Z(n24239) );
  AND2_X1 U3889 ( .A1(n7440), .A2(n52343), .ZN(n20876) );
  AND3_X1 U3894 ( .A1(n19878), .A2(n2929), .A3(n19879), .ZN(n7357) );
  BUF_X2 U3899 ( .A(n22915), .Z(n2175) );
  OR2_X1 U3957 ( .A1(n23445), .A2(n20903), .ZN(n22589) );
  NAND4_X1 U3967 ( .A1(n5782), .A2(n16397), .A3(n16399), .A4(n16398), .ZN(
        n23149) );
  NOR2_X1 U3976 ( .A1(n17632), .A2(n17631), .ZN(n22356) );
  AND2_X1 U3999 ( .A1(n18342), .A2(n18059), .ZN(n17428) );
  OR2_X1 U4008 ( .A1(n19059), .A2(n20122), .ZN(n4185) );
  NOR2_X1 U4016 ( .A1(n20449), .A2(n21490), .ZN(n51829) );
  NOR2_X1 U4034 ( .A1(n20812), .A2(n1365), .ZN(n51828) );
  AOI21_X1 U4043 ( .B1(n20193), .B2(n20628), .A(n51993), .ZN(n19941) );
  AND2_X1 U4056 ( .A1(n21533), .A2(n7484), .ZN(n51993) );
  INV_X1 U4082 ( .A(n21492), .ZN(n51754) );
  OR2_X1 U4093 ( .A1(n19663), .A2(n19636), .ZN(n51928) );
  AND2_X1 U4113 ( .A1(n19404), .A2(n2222), .ZN(n51946) );
  OR2_X1 U4121 ( .A1(n1763), .A2(n20428), .ZN(n20357) );
  NOR2_X1 U4123 ( .A1(n18999), .A2(n19796), .ZN(n19721) );
  BUF_X2 U4130 ( .A(n20026), .Z(n2166) );
  BUF_X2 U4142 ( .A(n19019), .Z(n51013) );
  OR2_X1 U4152 ( .A1(n52271), .A2(n20656), .ZN(n21663) );
  NOR2_X1 U4156 ( .A1(n774), .A2(n20493), .ZN(n19357) );
  INV_X2 U4180 ( .A(n19892), .ZN(n19662) );
  NAND2_X2 U4225 ( .A1(n15094), .A2(n18294), .ZN(n18282) );
  BUF_X1 U4244 ( .A(n18897), .Z(n52210) );
  OR2_X1 U4247 ( .A1(n634), .A2(n19359), .ZN(n20497) );
  BUF_X2 U4253 ( .A(n15872), .Z(n18873) );
  INV_X1 U4259 ( .A(n19947), .ZN(n3493) );
  OR2_X1 U4263 ( .A1(n20428), .A2(n20432), .ZN(n20343) );
  NAND2_X1 U4274 ( .A1(n21464), .A2(n634), .ZN(n21449) );
  XNOR2_X1 U4277 ( .A(n18545), .B(n18544), .ZN(n19947) );
  BUF_X2 U4285 ( .A(n21414), .Z(n51755) );
  NAND2_X2 U4286 ( .A1(n20062), .A2(n20052), .ZN(n19143) );
  INV_X1 U4324 ( .A(n20133), .ZN(n51756) );
  CLKBUF_X1 U4335 ( .A(n15846), .Z(n52194) );
  BUF_X2 U4360 ( .A(n18628), .Z(n51757) );
  OR2_X2 U4382 ( .A1(n7712), .A2(n7713), .ZN(n18443) );
  AND3_X1 U4413 ( .A1(n10867), .A2(n13456), .A3(n10868), .ZN(n12992) );
  BUF_X2 U4428 ( .A(n18168), .Z(n51758) );
  OAI21_X1 U4435 ( .B1(n13670), .B2(n13671), .A(n13669), .ZN(n13672) );
  AND3_X1 U4451 ( .A1(n11856), .A2(n11857), .A3(n11855), .ZN(n3958) );
  OR2_X1 U4456 ( .A1(n2871), .A2(n13376), .ZN(n13033) );
  AOI22_X1 U4484 ( .A1(n13973), .A2(n14231), .B1(n13974), .B2(n13975), .ZN(
        n16222) );
  OAI21_X1 U4486 ( .B1(n13671), .B2(n2763), .A(n8128), .ZN(n13673) );
  NOR2_X1 U4490 ( .A1(n13963), .A2(n12927), .ZN(n13967) );
  OR2_X1 U4524 ( .A1(n14303), .A2(n13832), .ZN(n52248) );
  OR2_X1 U4529 ( .A1(n15069), .A2(n15309), .ZN(n15071) );
  AND2_X1 U4547 ( .A1(n14296), .A2(n14294), .ZN(n52337) );
  INV_X1 U4554 ( .A(n7735), .ZN(n51984) );
  AND2_X1 U4567 ( .A1(n13948), .A2(n13930), .ZN(n11865) );
  INV_X2 U4584 ( .A(n14709), .ZN(n14719) );
  NAND2_X1 U4596 ( .A1(n2287), .A2(n8830), .ZN(n12204) );
  OR2_X1 U4606 ( .A1(n15384), .A2(n15358), .ZN(n14484) );
  NAND4_X2 U4609 ( .A1(n7148), .A2(n9240), .A3(n9241), .A4(n7149), .ZN(n15425)
         );
  AND2_X1 U4610 ( .A1(n12184), .A2(n12183), .ZN(n52423) );
  AND3_X1 U4626 ( .A1(n9107), .A2(n9101), .A3(n9100), .ZN(n52291) );
  OR3_X2 U4635 ( .A1(n9115), .A2(n9121), .A3(n9116), .ZN(n12756) );
  AND3_X1 U4645 ( .A1(n9518), .A2(n3583), .A3(n5658), .ZN(n52420) );
  OAI21_X1 U4658 ( .B1(n9861), .B2(n9862), .A(n10964), .ZN(n9866) );
  INV_X1 U4665 ( .A(n12090), .ZN(n52327) );
  OR2_X1 U4685 ( .A1(n11261), .A2(n12498), .ZN(n51971) );
  OR2_X1 U4695 ( .A1(n11499), .A2(n11496), .ZN(n11878) );
  AND2_X1 U4718 ( .A1(n12300), .A2(n10940), .ZN(n9655) );
  INV_X1 U4766 ( .A(n11209), .ZN(n51969) );
  NAND2_X1 U4801 ( .A1(n9305), .A2(n11640), .ZN(n11644) );
  INV_X1 U4808 ( .A(n10959), .ZN(n51988) );
  BUF_X2 U4812 ( .A(n11515), .Z(n51760) );
  INV_X1 U4822 ( .A(n10552), .ZN(n51761) );
  XNOR2_X1 U4842 ( .A(n9288), .B(Key[169]), .ZN(n52185) );
  INV_X1 U4843 ( .A(n11016), .ZN(n51762) );
  BUF_X2 U4845 ( .A(n11907), .Z(n2211) );
  INV_X1 U4849 ( .A(n9186), .ZN(n10457) );
  XNOR2_X1 U4881 ( .A(Ciphertext[24]), .B(Key[157]), .ZN(n9186) );
  OR2_X1 U4883 ( .A1(n11445), .A2(n12545), .ZN(n51883) );
  NAND2_X1 U4897 ( .A1(n11705), .A2(n9932), .ZN(n51968) );
  OR2_X1 U4902 ( .A1(n10134), .A2(n9807), .ZN(n9808) );
  AND2_X1 U4931 ( .A1(n12058), .A2(n10662), .ZN(n51936) );
  INV_X1 U4934 ( .A(n10143), .ZN(n10925) );
  OR2_X1 U4998 ( .A1(n12631), .A2(n12635), .ZN(n52319) );
  AND2_X1 U5010 ( .A1(n12532), .A2(n12545), .ZN(n11446) );
  INV_X1 U5099 ( .A(n12590), .ZN(n51846) );
  AND2_X1 U5103 ( .A1(n9973), .A2(n11268), .ZN(n11682) );
  OR2_X1 U5104 ( .A1(n10444), .A2(n52152), .ZN(n11977) );
  OR2_X1 U5118 ( .A1(n15279), .A2(n14950), .ZN(n14939) );
  BUF_X1 U5131 ( .A(n8908), .Z(n12680) );
  INV_X1 U5136 ( .A(n10127), .ZN(n10120) );
  AND2_X1 U5153 ( .A1(n9279), .A2(n9280), .ZN(n9087) );
  INV_X1 U5160 ( .A(n15046), .ZN(n51966) );
  OR2_X1 U5169 ( .A1(n11324), .A2(n12175), .ZN(n12152) );
  NOR2_X1 U5178 ( .A1(n52293), .A2(n52292), .ZN(n12273) );
  INV_X1 U5179 ( .A(n10346), .ZN(n52275) );
  BUF_X1 U5198 ( .A(n8818), .Z(n2197) );
  OR2_X1 U5208 ( .A1(n11605), .A2(n11600), .ZN(n9282) );
  AND4_X1 U5216 ( .A1(n8812), .A2(n8813), .A3(n10051), .A4(n8811), .ZN(n8814)
         );
  OR2_X1 U5222 ( .A1(n10884), .A2(n13525), .ZN(n12769) );
  OR2_X1 U5227 ( .A1(n2640), .A2(n13874), .ZN(n13257) );
  OAI21_X1 U5237 ( .B1(n10044), .B2(n9466), .A(n9953), .ZN(n9468) );
  AND2_X1 U5238 ( .A1(n14294), .A2(n14287), .ZN(n13573) );
  INV_X1 U5243 ( .A(n13172), .ZN(n10905) );
  AND2_X1 U5263 ( .A1(n14307), .A2(n13822), .ZN(n14319) );
  AND2_X1 U5277 ( .A1(n7711), .A2(n7717), .ZN(n51856) );
  NOR2_X1 U5281 ( .A1(n3679), .A2(n13148), .ZN(n3645) );
  OR2_X1 U5282 ( .A1(n51683), .A2(n955), .ZN(n11840) );
  AND2_X1 U5290 ( .A1(n13795), .A2(n51965), .ZN(n51964) );
  OR2_X1 U5294 ( .A1(n13256), .A2(n13257), .ZN(n52265) );
  OR2_X1 U5303 ( .A1(n14345), .A2(n14339), .ZN(n13418) );
  NOR2_X1 U5306 ( .A1(n14911), .A2(n15309), .ZN(n15063) );
  OR2_X1 U5334 ( .A1(n13449), .A2(n12787), .ZN(n13994) );
  OR2_X1 U5342 ( .A1(n13839), .A2(n13552), .ZN(n51861) );
  OR2_X1 U5343 ( .A1(n14605), .A2(n14011), .ZN(n12995) );
  XNOR2_X1 U5344 ( .A(n16980), .B(n15229), .ZN(n52388) );
  BUF_X1 U5345 ( .A(n17671), .Z(n51458) );
  OR2_X1 U5367 ( .A1(n11311), .A2(n12949), .ZN(n11314) );
  NOR2_X1 U5374 ( .A1(n51948), .A2(n13003), .ZN(n13401) );
  AND2_X1 U5375 ( .A1(n14289), .A2(n14285), .ZN(n14291) );
  AND3_X1 U5383 ( .A1(n13694), .A2(n13691), .A3(n13693), .ZN(n52419) );
  AND3_X1 U5385 ( .A1(n9692), .A2(n9691), .A3(n51861), .ZN(n9728) );
  OR2_X1 U5401 ( .A1(n13884), .A2(n13883), .ZN(n51939) );
  INV_X1 U5403 ( .A(n2640), .ZN(n14875) );
  NAND4_X1 U5433 ( .A1(n12911), .A2(n12909), .A3(n12908), .A4(n12910), .ZN(
        n18777) );
  AND2_X1 U5438 ( .A1(n14100), .A2(n14103), .ZN(n14097) );
  CLKBUF_X1 U5449 ( .A(n18815), .Z(n51414) );
  BUF_X1 U5451 ( .A(n18628), .Z(n52209) );
  OR3_X1 U5463 ( .A1(n20628), .A2(n20201), .A3(n20624), .ZN(n18455) );
  OR2_X1 U5486 ( .A1(n19535), .A2(n16490), .ZN(n20116) );
  INV_X1 U5502 ( .A(n16490), .ZN(n20156) );
  OR2_X1 U5542 ( .A1(n17576), .A2(n7956), .ZN(n18023) );
  AND2_X1 U5567 ( .A1(n20014), .A2(n20013), .ZN(n51207) );
  AND2_X1 U5633 ( .A1(n20389), .A2(n17639), .ZN(n52005) );
  INV_X1 U5637 ( .A(n18024), .ZN(n51934) );
  OR2_X1 U5643 ( .A1(n51021), .A2(n23167), .ZN(n52289) );
  NOR2_X1 U5651 ( .A1(n18938), .A2(n19663), .ZN(n51906) );
  AND2_X1 U5655 ( .A1(n20104), .A2(n17059), .ZN(n18316) );
  AND2_X1 U5660 ( .A1(n20427), .A2(n20435), .ZN(n19326) );
  OR3_X1 U5670 ( .A1(n18318), .A2(n16788), .A3(n16787), .ZN(n16789) );
  AND2_X1 U5671 ( .A1(n20135), .A2(n52037), .ZN(n51816) );
  OR2_X1 U5678 ( .A1(n18316), .A2(n20097), .ZN(n17605) );
  AND2_X1 U5679 ( .A1(n21491), .A2(n21480), .ZN(n51827) );
  NAND2_X1 U5683 ( .A1(n19678), .A2(n18921), .ZN(n20210) );
  OR2_X1 U5691 ( .A1(n17503), .A2(n17056), .ZN(n20089) );
  AND2_X1 U5704 ( .A1(n52037), .A2(n20132), .ZN(n19061) );
  AND2_X1 U5716 ( .A1(n17997), .A2(n17639), .ZN(n19380) );
  AND2_X1 U5740 ( .A1(n19994), .A2(n19995), .ZN(n52255) );
  XNOR2_X1 U5810 ( .A(n16359), .B(n16358), .ZN(n17047) );
  OAI21_X1 U5822 ( .B1(n17070), .B2(n51817), .A(n51816), .ZN(n17072) );
  INV_X1 U5823 ( .A(n21872), .ZN(n51859) );
  OR2_X1 U5826 ( .A1(n22593), .A2(n20903), .ZN(n22009) );
  AND3_X1 U5831 ( .A1(n20229), .A2(n8095), .A3(n8094), .ZN(n20237) );
  AND2_X1 U5835 ( .A1(n51222), .A2(n51132), .ZN(n19472) );
  NOR2_X1 U5842 ( .A1(n3167), .A2(n18848), .ZN(n20667) );
  OR2_X1 U5848 ( .A1(n23924), .A2(n23895), .ZN(n3904) );
  AND2_X1 U5854 ( .A1(n22978), .A2(n22989), .ZN(n52247) );
  AND2_X1 U5878 ( .A1(n52155), .A2(n17420), .ZN(n51930) );
  OR2_X1 U5879 ( .A1(n19609), .A2(n22864), .ZN(n22328) );
  OR2_X1 U5893 ( .A1(n21895), .A2(n23504), .ZN(n51836) );
  OR2_X1 U5898 ( .A1(n19693), .A2(n51954), .ZN(n18920) );
  OAI211_X1 U5905 ( .C1(n18337), .C2(n18336), .A(n18335), .B(n18334), .ZN(
        n20965) );
  OR3_X1 U5907 ( .A1(n21950), .A2(n51123), .A3(n2076), .ZN(n21955) );
  AND2_X1 U5913 ( .A1(n23306), .A2(n23314), .ZN(n51875) );
  OR2_X1 U5927 ( .A1(n22354), .A2(n22901), .ZN(n3022) );
  AND2_X1 U5940 ( .A1(n23080), .A2(n22268), .ZN(n23599) );
  BUF_X1 U5976 ( .A(n21925), .Z(n50991) );
  AND2_X1 U5977 ( .A1(n23531), .A2(n457), .ZN(n24330) );
  AND4_X1 U5982 ( .A1(n5103), .A2(n22531), .A3(n22420), .A4(n24002), .ZN(n5102) );
  OR2_X1 U5985 ( .A1(n23338), .A2(n21755), .ZN(n21140) );
  AOI21_X1 U5990 ( .B1(n21025), .B2(n17614), .A(n52381), .ZN(n3665) );
  INV_X1 U5991 ( .A(n20270), .ZN(n1704) );
  INV_X1 U5993 ( .A(n24111), .ZN(n24414) );
  AND2_X1 U6004 ( .A1(n6621), .A2(n23161), .ZN(n3109) );
  NOR2_X1 U6019 ( .A1(n23876), .A2(n23877), .ZN(n51992) );
  OR2_X1 U6032 ( .A1(n23700), .A2(n23533), .ZN(n52295) );
  OR2_X1 U6052 ( .A1(n23603), .A2(n23595), .ZN(n51960) );
  AND3_X1 U6056 ( .A1(n21004), .A2(n18959), .A3(n18926), .ZN(n52276) );
  AND2_X1 U6062 ( .A1(n22969), .A2(n22971), .ZN(n52277) );
  AOI22_X1 U6066 ( .A1(n19999), .A2(n24033), .B1(n20000), .B2(n20001), .ZN(
        n20008) );
  OR2_X1 U6072 ( .A1(n22601), .A2(n24188), .ZN(n23196) );
  NOR2_X1 U6082 ( .A1(n22149), .A2(n21919), .ZN(n21030) );
  INV_X1 U6107 ( .A(n22576), .ZN(n22578) );
  AND3_X1 U6108 ( .A1(n52295), .A2(n51581), .A3(n52294), .ZN(n23544) );
  XNOR2_X1 U6113 ( .A(n1377), .B(n28287), .ZN(n26221) );
  XNOR2_X1 U6128 ( .A(n25510), .B(n25354), .ZN(n25355) );
  XNOR2_X1 U6151 ( .A(n51955), .B(n27196), .ZN(n27417) );
  XNOR2_X1 U6152 ( .A(n51119), .B(n52238), .ZN(n24220) );
  AND2_X1 U6153 ( .A1(n2956), .A2(n26668), .ZN(n51821) );
  XNOR2_X1 U6162 ( .A(n25936), .B(n25820), .ZN(n51927) );
  XOR2_X1 U6189 ( .A(n24516), .B(n24515), .Z(n2401) );
  OR2_X1 U6191 ( .A1(n27628), .A2(n27629), .ZN(n8273) );
  AND2_X1 U6192 ( .A1(n28636), .A2(n459), .ZN(n51958) );
  OR2_X1 U6193 ( .A1(n27711), .A2(n26998), .ZN(n27709) );
  AND2_X1 U6215 ( .A1(n26901), .A2(n51768), .ZN(n52360) );
  BUF_X1 U6224 ( .A(n27525), .Z(n30698) );
  OR2_X1 U6225 ( .A1(n29264), .A2(n30218), .ZN(n28663) );
  OR2_X1 U6259 ( .A1(n27820), .A2(n27821), .ZN(n27894) );
  AND2_X1 U6265 ( .A1(n32240), .A2(n32231), .ZN(n51961) );
  NAND2_X1 U6310 ( .A1(n27162), .A2(n30706), .ZN(n30709) );
  OR2_X1 U6311 ( .A1(n27706), .A2(n51772), .ZN(n29423) );
  INV_X1 U6321 ( .A(n29289), .ZN(n29300) );
  NAND2_X1 U6323 ( .A1(n27162), .A2(n2109), .ZN(n30712) );
  NOR2_X1 U6327 ( .A1(n52418), .A2(n27163), .ZN(n27542) );
  BUF_X1 U6328 ( .A(n28145), .Z(n2195) );
  AND2_X1 U6347 ( .A1(n28998), .A2(n29736), .ZN(n30444) );
  OR2_X1 U6357 ( .A1(n51489), .A2(n29764), .ZN(n29068) );
  AND2_X1 U6358 ( .A1(n30791), .A2(n23658), .ZN(n29909) );
  AND2_X1 U6368 ( .A1(n31106), .A2(n30058), .ZN(n51863) );
  CLKBUF_X1 U6378 ( .A(n27729), .Z(n2144) );
  AND2_X1 U6381 ( .A1(n29156), .A2(n30245), .ZN(n52352) );
  AND2_X1 U6406 ( .A1(n459), .A2(n51107), .ZN(n29317) );
  OAI211_X1 U6416 ( .C1(n26961), .C2(n26960), .A(n26959), .B(n26958), .ZN(
        n26967) );
  INV_X1 U6419 ( .A(n28155), .ZN(n29035) );
  OR2_X1 U6451 ( .A1(n26679), .A2(n26676), .ZN(n29498) );
  AND2_X1 U6461 ( .A1(n28547), .A2(n30291), .ZN(n51842) );
  OR2_X1 U6462 ( .A1(n27562), .A2(n5769), .ZN(n1637) );
  OR2_X1 U6464 ( .A1(n31489), .A2(n31484), .ZN(n29837) );
  AND3_X1 U6476 ( .A1(n27823), .A2(n27826), .A3(n27824), .ZN(n838) );
  INV_X1 U6479 ( .A(n31158), .ZN(n52364) );
  INV_X1 U6489 ( .A(n33155), .ZN(n52390) );
  OR2_X1 U6516 ( .A1(n28959), .A2(n5056), .ZN(n52249) );
  INV_X1 U6518 ( .A(n28896), .ZN(n28905) );
  AND2_X1 U6519 ( .A1(n51106), .A2(n7064), .ZN(n31553) );
  AOI22_X1 U6525 ( .A1(n24990), .A2(n30249), .B1(n24988), .B2(n52352), .ZN(
        n2830) );
  NOR2_X1 U6526 ( .A1(n51178), .A2(n4082), .ZN(n8710) );
  AND2_X1 U6535 ( .A1(n27966), .A2(n27965), .ZN(n52315) );
  NAND4_X1 U6536 ( .A1(n26470), .A2(n26471), .A3(n26469), .A4(n26472), .ZN(
        n31384) );
  OR2_X1 U6562 ( .A1(n29677), .A2(n7667), .ZN(n31991) );
  INV_X1 U6563 ( .A(n30642), .ZN(n30640) );
  NOR2_X1 U6565 ( .A1(n31155), .A2(n52364), .ZN(n8746) );
  NOR2_X1 U6585 ( .A1(n5278), .A2(n30593), .ZN(n31093) );
  AND2_X1 U6603 ( .A1(n52407), .A2(n31297), .ZN(n52333) );
  AND2_X1 U6615 ( .A1(n31699), .A2(n31700), .ZN(n32119) );
  INV_X1 U6616 ( .A(n31749), .ZN(n31743) );
  AND3_X1 U6617 ( .A1(n8239), .A2(n8238), .A3(n31629), .ZN(n51590) );
  OR2_X1 U6639 ( .A1(n28487), .A2(n31873), .ZN(n31879) );
  AOI22_X1 U6645 ( .A1(n31180), .A2(n32671), .B1(n31181), .B2(n31182), .ZN(
        n31183) );
  OR2_X1 U6661 ( .A1(n30882), .A2(n31991), .ZN(n32003) );
  MUX2_X1 U6662 ( .A(n31587), .B(n31582), .S(n31581), .Z(n31591) );
  OR2_X1 U6683 ( .A1(n32409), .A2(n32394), .ZN(n32065) );
  AND3_X1 U6688 ( .A1(n32705), .A2(n31668), .A3(n52301), .ZN(n30144) );
  AND2_X1 U6695 ( .A1(n711), .A2(n32299), .ZN(n31845) );
  NOR2_X1 U6697 ( .A1(n5935), .A2(n6239), .ZN(n51841) );
  AND2_X1 U6708 ( .A1(n31389), .A2(n33021), .ZN(n6422) );
  OAI21_X1 U6709 ( .B1(n31494), .B2(n31495), .A(n31493), .ZN(n31505) );
  NOR2_X1 U6716 ( .A1(n2994), .A2(n2993), .ZN(n28946) );
  XNOR2_X1 U6717 ( .A(n37278), .B(n37276), .ZN(n52405) );
  AOI22_X1 U6720 ( .A1(n51976), .A2(n32871), .B1(n32873), .B2(n5498), .ZN(
        n32892) );
  INV_X1 U6726 ( .A(n32843), .ZN(n31914) );
  AOI22_X1 U6739 ( .A1(n31745), .A2(n32295), .B1(n32302), .B2(n31845), .ZN(
        n31756) );
  CLKBUF_X1 U6749 ( .A(n35603), .Z(n51381) );
  XNOR2_X1 U6758 ( .A(n35586), .B(n34549), .ZN(n35494) );
  XNOR2_X1 U6759 ( .A(n34821), .B(n34815), .ZN(n51862) );
  INV_X1 U6779 ( .A(n34122), .ZN(n36858) );
  XNOR2_X1 U6780 ( .A(n7199), .B(n702), .ZN(n33540) );
  AND2_X1 U6784 ( .A1(n6825), .A2(n39399), .ZN(n37730) );
  INV_X1 U6785 ( .A(n51324), .ZN(n51874) );
  INV_X1 U6801 ( .A(n52156), .ZN(n51909) );
  AND2_X1 U6802 ( .A1(n39399), .A2(n39400), .ZN(n51809) );
  INV_X1 U6821 ( .A(n38007), .ZN(n34970) );
  OR2_X1 U6824 ( .A1(n39208), .A2(n38950), .ZN(n52242) );
  AND2_X1 U6829 ( .A1(n34692), .A2(n37781), .ZN(n36199) );
  XNOR2_X1 U6830 ( .A(n1113), .B(n32339), .ZN(n36364) );
  XNOR2_X1 U6833 ( .A(n3061), .B(n7385), .ZN(n37881) );
  NOR2_X1 U6834 ( .A1(n34692), .A2(n37781), .ZN(n33461) );
  INV_X1 U6842 ( .A(n33871), .ZN(n39479) );
  NOR2_X1 U6881 ( .A1(n38075), .A2(n34960), .ZN(n38089) );
  AND2_X1 U6889 ( .A1(n36574), .A2(n2443), .ZN(n51918) );
  AND2_X1 U6904 ( .A1(n36492), .A2(n36473), .ZN(n36572) );
  AND2_X1 U6909 ( .A1(n37809), .A2(n37805), .ZN(n37798) );
  AND2_X1 U6911 ( .A1(n37779), .A2(n37782), .ZN(n51830) );
  OR2_X1 U6914 ( .A1(n34976), .A2(n38007), .ZN(n52279) );
  NOR2_X1 U6918 ( .A1(n41057), .A2(n41049), .ZN(n40510) );
  AND2_X1 U6958 ( .A1(n33062), .A2(n38561), .ZN(n38576) );
  INV_X1 U6959 ( .A(n2571), .ZN(n51956) );
  OR2_X1 U6970 ( .A1(n6637), .A2(n38475), .ZN(n36112) );
  OR2_X1 U6971 ( .A1(n37976), .A2(n37983), .ZN(n36529) );
  INV_X1 U6972 ( .A(n37882), .ZN(n39390) );
  AND2_X1 U6976 ( .A1(n5312), .A2(n38573), .ZN(n35709) );
  XNOR2_X1 U6978 ( .A(n33369), .B(n33368), .ZN(n35923) );
  AND2_X1 U6991 ( .A1(n37815), .A2(n8332), .ZN(n40258) );
  AND2_X1 U7000 ( .A1(n34965), .A2(n34966), .ZN(n51995) );
  AND2_X1 U7001 ( .A1(n38628), .A2(n35305), .ZN(n37689) );
  AND2_X1 U7039 ( .A1(n36414), .A2(n37648), .ZN(n36396) );
  OR2_X1 U7068 ( .A1(n38947), .A2(n39210), .ZN(n52000) );
  OR2_X1 U7072 ( .A1(n197), .A2(n38630), .ZN(n38262) );
  NOR2_X1 U7089 ( .A1(n42061), .A2(n41489), .ZN(n41482) );
  OR2_X1 U7098 ( .A1(n39286), .A2(n51956), .ZN(n4069) );
  NAND2_X1 U7099 ( .A1(n6317), .A2(n35103), .ZN(n38478) );
  AND3_X1 U7115 ( .A1(n39434), .A2(n39420), .A3(n39421), .ZN(n52244) );
  NOR2_X1 U7117 ( .A1(n4954), .A2(n40572), .ZN(n35718) );
  AND2_X1 U7128 ( .A1(n37871), .A2(n40340), .ZN(n52011) );
  AND2_X1 U7146 ( .A1(n37768), .A2(n37767), .ZN(n37769) );
  AOI22_X1 U7192 ( .A1(n37669), .A2(n38339), .B1(n37671), .B2(n37668), .ZN(
        n37676) );
  AND2_X1 U7207 ( .A1(n37532), .A2(n33557), .ZN(n38510) );
  AND2_X1 U7210 ( .A1(n41263), .A2(n40477), .ZN(n52413) );
  OR2_X1 U7224 ( .A1(n39949), .A2(n51879), .ZN(n6370) );
  AND2_X1 U7228 ( .A1(n40525), .A2(n1984), .ZN(n51891) );
  OR2_X1 U7229 ( .A1(n41065), .A2(n40502), .ZN(n40506) );
  AND2_X1 U7248 ( .A1(n40088), .A2(n40087), .ZN(n51972) );
  CLKBUF_X1 U7249 ( .A(n41978), .Z(n52080) );
  AND2_X1 U7254 ( .A1(n35858), .A2(n39314), .ZN(n52237) );
  INV_X1 U7263 ( .A(n40967), .ZN(n51394) );
  AND2_X1 U7293 ( .A1(n43334), .A2(n43331), .ZN(n51855) );
  OR2_X1 U7294 ( .A1(n52198), .A2(n41245), .ZN(n41673) );
  OR2_X2 U7312 ( .A1(n37908), .A2(n37909), .ZN(n41540) );
  AND2_X1 U7340 ( .A1(n1984), .A2(n40869), .ZN(n40876) );
  INV_X1 U7341 ( .A(n39101), .ZN(n40015) );
  AND2_X1 U7350 ( .A1(n43329), .A2(n43327), .ZN(n41010) );
  OR2_X2 U7359 ( .A1(n6085), .A2(n6086), .ZN(n41646) );
  AND3_X1 U7365 ( .A1(n51990), .A2(n40823), .A3(n40818), .ZN(n39692) );
  XNOR2_X1 U7386 ( .A(n40307), .B(n43943), .ZN(n40308) );
  AND2_X1 U7388 ( .A1(n6961), .A2(n51297), .ZN(n38416) );
  AND2_X1 U7389 ( .A1(n38804), .A2(n38793), .ZN(n52299) );
  AND2_X1 U7414 ( .A1(n41052), .A2(n52357), .ZN(n2345) );
  OR2_X1 U7432 ( .A1(n41390), .A2(n41391), .ZN(n6506) );
  INV_X1 U7433 ( .A(n40823), .ZN(n40835) );
  OR2_X1 U7466 ( .A1(n40373), .A2(n41902), .ZN(n39628) );
  OR2_X1 U7467 ( .A1(n41702), .A2(n41693), .ZN(n41168) );
  AOI22_X1 U7475 ( .A1(n51889), .A2(n42109), .B1(n51734), .B2(n42107), .ZN(
        n42115) );
  AND2_X1 U7477 ( .A1(n40838), .A2(n40823), .ZN(n40831) );
  AND4_X1 U7496 ( .A1(n41550), .A2(n51819), .A3(n41548), .A4(n51818), .ZN(
        n41558) );
  OAI21_X1 U7509 ( .B1(n2363), .B2(n40182), .A(n40663), .ZN(n40191) );
  AND4_X1 U7518 ( .A1(n6506), .A2(n6504), .A3(n40992), .A4(n40993), .ZN(n6503)
         );
  OAI21_X1 U7540 ( .B1(n37861), .B2(n41606), .A(n41604), .ZN(n41302) );
  AND3_X1 U7544 ( .A1(n35005), .A2(n35008), .A3(n6212), .ZN(n6211) );
  NOR2_X1 U7545 ( .A1(n41779), .A2(n41778), .ZN(n43496) );
  XNOR2_X1 U7548 ( .A(n43219), .B(n42450), .ZN(n45390) );
  CLKBUF_X1 U7552 ( .A(n45091), .Z(n52123) );
  OR2_X1 U7561 ( .A1(n49209), .A2(n49201), .ZN(n52259) );
  OR2_X1 U7563 ( .A1(n46201), .A2(n52079), .ZN(n51957) );
  CLKBUF_X1 U7564 ( .A(n45067), .Z(n52135) );
  XNOR2_X1 U7566 ( .A(n52013), .B(n51529), .ZN(n41908) );
  OR2_X1 U7577 ( .A1(n2207), .A2(n48546), .ZN(n51844) );
  BUF_X1 U7578 ( .A(n46510), .Z(n668) );
  OR2_X1 U7580 ( .A1(n49177), .A2(n539), .ZN(n45653) );
  CLKBUF_X1 U7587 ( .A(n43479), .Z(n43474) );
  INV_X1 U7588 ( .A(n49146), .ZN(n2695) );
  AND2_X1 U7638 ( .A1(n49740), .A2(n50035), .ZN(n51963) );
  INV_X1 U7645 ( .A(n2806), .ZN(n47342) );
  CLKBUF_X1 U7681 ( .A(n44085), .Z(n52196) );
  INV_X1 U7687 ( .A(n45138), .ZN(n47128) );
  AND2_X1 U7719 ( .A1(n46522), .A2(n51068), .ZN(n46521) );
  NOR2_X1 U7725 ( .A1(n49278), .A2(n49265), .ZN(n6026) );
  NAND2_X1 U7733 ( .A1(n46163), .A2(n50034), .ZN(n50387) );
  BUF_X1 U7735 ( .A(n43687), .Z(n46999) );
  XNOR2_X1 U7747 ( .A(n43617), .B(n43616), .ZN(n46888) );
  AND2_X1 U7791 ( .A1(n44850), .A2(n46730), .ZN(n46743) );
  INV_X1 U7816 ( .A(n47841), .ZN(n51941) );
  AND2_X1 U7828 ( .A1(n48522), .A2(n46471), .ZN(n48510) );
  AND3_X1 U7888 ( .A1(n1643), .A2(n45596), .A3(n45595), .ZN(n52415) );
  AND3_X1 U7919 ( .A1(n52032), .A2(n46453), .A3(n46451), .ZN(n52031) );
  OAI21_X1 U7978 ( .B1(n49204), .B2(n49203), .A(n52304), .ZN(n49221) );
  OR2_X1 U7980 ( .A1(n47368), .A2(n49993), .ZN(n50328) );
  AND2_X1 U7993 ( .A1(n1567), .A2(n47120), .ZN(n47133) );
  INV_X1 U7997 ( .A(n50935), .ZN(n47397) );
  AND2_X1 U8017 ( .A1(n51916), .A2(n45692), .ZN(n2306) );
  OAI211_X1 U8019 ( .C1(n45647), .C2(n45646), .A(n49162), .B(n45645), .ZN(
        n5689) );
  AND2_X1 U8054 ( .A1(n46954), .A2(n46951), .ZN(n51824) );
  AND4_X1 U8093 ( .A1(n45956), .A2(n45955), .A3(n45954), .A4(n45953), .ZN(
        n49432) );
  NOR2_X1 U8102 ( .A1(n50640), .A2(n50638), .ZN(n50610) );
  BUF_X1 U8167 ( .A(n48083), .Z(n52127) );
  INV_X1 U8186 ( .A(n48112), .ZN(n48157) );
  AND4_X1 U8202 ( .A1(n4787), .A2(n46460), .A3(n336), .A4(n46461), .ZN(n52157)
         );
  AND3_X1 U8220 ( .A1(n2898), .A2(n42802), .A3(n42803), .ZN(n52137) );
  OR2_X1 U8232 ( .A1(n49433), .A2(n49461), .ZN(n51893) );
  NOR2_X1 U8243 ( .A1(n49960), .A2(n49959), .ZN(n52055) );
  AND2_X1 U8293 ( .A1(n5365), .A2(n50958), .ZN(n50901) );
  CLKBUF_X2 U8338 ( .A(Key[37]), .Z(n4754) );
  INV_X1 U8353 ( .A(n48353), .ZN(n48380) );
  AOI22_X1 U8375 ( .A1(n50551), .A2(n5263), .B1(n5264), .B2(n50539), .ZN(
        n47055) );
  BUF_X1 U8427 ( .A(Key[62]), .Z(n4886) );
  AND3_X1 U8443 ( .A1(n16046), .A2(n16047), .A3(n52303), .ZN(n51763) );
  AND2_X1 U8458 ( .A1(n15259), .A2(n14137), .ZN(n51764) );
  AND2_X1 U8474 ( .A1(n3700), .A2(n3694), .ZN(n51765) );
  AND2_X1 U8487 ( .A1(n48259), .A2(n48260), .ZN(n51766) );
  AND2_X1 U8501 ( .A1(n28146), .A2(n2195), .ZN(n51767) );
  OR2_X1 U8512 ( .A1(n26989), .A2(n29422), .ZN(n51768) );
  AND2_X1 U8515 ( .A1(n10978), .A2(n9782), .ZN(n51769) );
  OR2_X1 U8551 ( .A1(n27623), .A2(n27638), .ZN(n51770) );
  AND2_X1 U8555 ( .A1(n27056), .A2(n29568), .ZN(n51771) );
  AND2_X1 U8563 ( .A1(n51351), .A2(n51112), .ZN(n51772) );
  NAND2_X1 U8586 ( .A1(n18961), .A2(n51132), .ZN(n51773) );
  AND3_X1 U8635 ( .A1(n19062), .A2(n19066), .A3(n574), .ZN(n51774) );
  OR2_X1 U8673 ( .A1(n40633), .A2(n51950), .ZN(n51775) );
  AND4_X1 U8682 ( .A1(n20388), .A2(n20387), .A3(n20386), .A4(n20477), .ZN(
        n51776) );
  AND2_X1 U8712 ( .A1(n40486), .A2(n39598), .ZN(n51777) );
  AND2_X1 U8789 ( .A1(n37426), .A2(n35445), .ZN(n51778) );
  AND3_X1 U8812 ( .A1(n37415), .A2(n38471), .A3(n35446), .ZN(n51779) );
  AND3_X1 U8864 ( .A1(n51980), .A2(n23644), .A3(n51788), .ZN(n51780) );
  AND2_X1 U8889 ( .A1(n27146), .A2(n30245), .ZN(n51781) );
  OR2_X1 U8890 ( .A1(n10526), .A2(n10525), .ZN(n51782) );
  OR2_X1 U8938 ( .A1(n10100), .A2(n10101), .ZN(n51783) );
  AND2_X1 U8969 ( .A1(n52007), .A2(n52006), .ZN(n51784) );
  INV_X1 U8979 ( .A(n12976), .ZN(n52312) );
  INV_X1 U9018 ( .A(n20114), .ZN(n51815) );
  INV_X1 U9057 ( .A(n19676), .ZN(n51954) );
  XOR2_X1 U9058 ( .A(n16759), .B(n16758), .Z(n51785) );
  AND2_X1 U9082 ( .A1(n22053), .A2(n22051), .ZN(n51786) );
  OR2_X1 U9112 ( .A1(n23013), .A2(n4847), .ZN(n51787) );
  OR2_X1 U9142 ( .A1(n23645), .A2(n5068), .ZN(n51788) );
  AND3_X1 U9194 ( .A1(n23593), .A2(n23594), .A3(n51960), .ZN(n51789) );
  OR2_X1 U9235 ( .A1(n30174), .A2(n30178), .ZN(n51790) );
  AND2_X1 U9255 ( .A1(n7604), .A2(n7605), .ZN(n51791) );
  NAND2_X1 U9269 ( .A1(n26888), .A2(n27732), .ZN(n51792) );
  INV_X1 U9308 ( .A(n5056), .ZN(n52251) );
  XOR2_X1 U9418 ( .A(n7560), .B(n25966), .Z(n51793) );
  AND2_X1 U9422 ( .A1(n31503), .A2(n31504), .ZN(n51794) );
  OR2_X1 U9465 ( .A1(n32075), .A2(n32402), .ZN(n51795) );
  AND2_X1 U9472 ( .A1(n32075), .A2(n32396), .ZN(n51796) );
  AND3_X1 U9520 ( .A1(n32589), .A2(n30502), .A3(n32987), .ZN(n51797) );
  INV_X1 U9564 ( .A(n36035), .ZN(n37957) );
  XOR2_X1 U9612 ( .A(n35504), .B(n35837), .Z(n51798) );
  AND2_X1 U9631 ( .A1(n39191), .A2(n37037), .ZN(n51799) );
  AND2_X1 U9634 ( .A1(n1742), .A2(n36520), .ZN(n51800) );
  AND3_X1 U9665 ( .A1(n38436), .A2(n6645), .A3(n39914), .ZN(n51801) );
  INV_X1 U9675 ( .A(n41792), .ZN(n51950) );
  OR2_X1 U9689 ( .A1(n49232), .A2(n49231), .ZN(n51802) );
  AND2_X1 U9742 ( .A1(n46685), .A2(n46606), .ZN(n51803) );
  OR2_X1 U9773 ( .A1(n48127), .A2(n48159), .ZN(n51804) );
  AND4_X1 U9829 ( .A1(n44690), .A2(n44688), .A3(n44689), .A4(n44687), .ZN(
        n51805) );
  AND2_X1 U9874 ( .A1(n46919), .A2(n46912), .ZN(n51806) );
  NAND2_X1 U9876 ( .A1(n29442), .A2(n29439), .ZN(n27034) );
  XNOR2_X2 U9916 ( .A(n26024), .B(n26023), .ZN(n29439) );
  NAND2_X1 U9932 ( .A1(n29063), .A2(n29062), .ZN(n29773) );
  AND2_X2 U9939 ( .A1(n30354), .A2(n29764), .ZN(n29063) );
  BUF_X1 U9958 ( .A(n1946), .Z(n52069) );
  NAND2_X1 U10003 ( .A1(n51895), .A2(n1088), .ZN(n1626) );
  NAND2_X1 U10018 ( .A1(n51807), .A2(n41683), .ZN(n8124) );
  NAND4_X1 U10023 ( .A1(n41673), .A2(n41685), .A3(n40037), .A4(n41680), .ZN(
        n51807) );
  AND4_X2 U10033 ( .A1(n36479), .A2(n36477), .A3(n36476), .A4(n36478), .ZN(
        n36502) );
  NOR2_X1 U10069 ( .A1(n40700), .A2(n51808), .ZN(n40707) );
  OAI21_X1 U10110 ( .B1(n6235), .B2(n42008), .A(n41583), .ZN(n51808) );
  NAND2_X1 U10125 ( .A1(n51814), .A2(n51811), .ZN(n19548) );
  NAND2_X1 U10133 ( .A1(n51813), .A2(n51812), .ZN(n51811) );
  AOI21_X1 U10152 ( .B1(n19536), .B2(n16490), .A(n51815), .ZN(n51812) );
  NAND2_X1 U10170 ( .A1(n19540), .A2(n20155), .ZN(n51813) );
  NAND2_X1 U10253 ( .A1(n19539), .A2(n51815), .ZN(n51814) );
  XNOR2_X1 U10301 ( .A(n6368), .B(n26064), .ZN(n52394) );
  NAND2_X1 U10309 ( .A1(n2870), .A2(n51803), .ZN(n46621) );
  NAND2_X1 U10339 ( .A1(n7839), .A2(n20145), .ZN(n51817) );
  NAND2_X1 U10358 ( .A1(n41542), .A2(n41543), .ZN(n51818) );
  NAND2_X1 U10389 ( .A1(n41541), .A2(n41540), .ZN(n51819) );
  AOI22_X1 U10393 ( .A1(n19945), .A2(n19946), .B1(n316), .B2(n19947), .ZN(
        n19964) );
  NAND2_X1 U10444 ( .A1(n6397), .A2(n6396), .ZN(n811) );
  NAND3_X1 U10495 ( .A1(n23904), .A2(n51033), .A3(n23903), .ZN(n23918) );
  NAND4_X1 U10496 ( .A1(n51820), .A2(n11191), .A3(n11185), .A4(n11570), .ZN(
        n11197) );
  NAND2_X1 U10550 ( .A1(n11189), .A2(n11186), .ZN(n51820) );
  XNOR2_X2 U10579 ( .A(n42850), .B(n44237), .ZN(n43143) );
  NAND4_X2 U10584 ( .A1(n35996), .A2(n7171), .A3(n7173), .A4(n38926), .ZN(
        n42850) );
  NAND2_X1 U10595 ( .A1(n28831), .A2(n28832), .ZN(n28833) );
  NAND2_X1 U10602 ( .A1(n26666), .A2(n28674), .ZN(n25836) );
  NAND2_X1 U10606 ( .A1(n29478), .A2(n51821), .ZN(n28674) );
  NAND2_X2 U10630 ( .A1(n28847), .A2(n51822), .ZN(n32843) );
  XNOR2_X1 U10688 ( .A(n35496), .B(n51798), .ZN(n35507) );
  XNOR2_X1 U10750 ( .A(n33817), .B(n37040), .ZN(n35496) );
  NAND2_X1 U10779 ( .A1(n31155), .A2(n51823), .ZN(n31157) );
  OAI21_X1 U10844 ( .B1(n31463), .B2(n51106), .A(n32610), .ZN(n51823) );
  NAND2_X1 U10912 ( .A1(n46952), .A2(n51824), .ZN(n46960) );
  OAI211_X1 U10925 ( .C1(n39251), .C2(n39250), .A(n51825), .B(n39249), .ZN(
        n39252) );
  NAND2_X1 U10948 ( .A1(n4258), .A2(n4257), .ZN(n51825) );
  AND2_X1 U10974 ( .A1(n38549), .A2(n38547), .ZN(n35171) );
  INV_X1 U10977 ( .A(n13907), .ZN(n15447) );
  NAND2_X1 U10978 ( .A1(n15435), .A2(n15437), .ZN(n13907) );
  NAND2_X1 U10985 ( .A1(n19798), .A2(n19802), .ZN(n19805) );
  NAND2_X1 U10986 ( .A1(n46348), .A2(n46347), .ZN(n46351) );
  OR2_X2 U11009 ( .A1(n51826), .A2(n36166), .ZN(n41211) );
  NAND4_X1 U11029 ( .A1(n36164), .A2(n36162), .A3(n36163), .A4(n36165), .ZN(
        n51826) );
  AND2_X1 U11075 ( .A1(n23992), .A2(n24001), .ZN(n2008) );
  NAND3_X1 U11154 ( .A1(n32877), .A2(n8544), .A3(n32876), .ZN(n32878) );
  NAND2_X1 U11164 ( .A1(n18990), .A2(n19715), .ZN(n18890) );
  OAI21_X1 U11165 ( .B1(n51829), .B2(n51828), .A(n51827), .ZN(n19282) );
  AOI21_X1 U11190 ( .B1(n34684), .B2(n34685), .A(n51830), .ZN(n34697) );
  NOR2_X2 U11217 ( .A1(n945), .A2(n944), .ZN(n26160) );
  NAND2_X1 U11223 ( .A1(n51833), .A2(n51831), .ZN(n23349) );
  NAND2_X1 U11317 ( .A1(n23329), .A2(n51832), .ZN(n51831) );
  NAND2_X1 U11322 ( .A1(n23328), .A2(n1024), .ZN(n51833) );
  NAND3_X1 U11330 ( .A1(n22257), .A2(n21758), .A3(n629), .ZN(n23328) );
  NAND2_X1 U11410 ( .A1(n51834), .A2(n9186), .ZN(n11986) );
  INV_X1 U11488 ( .A(n9178), .ZN(n51834) );
  INV_X1 U11491 ( .A(n21010), .ZN(n51858) );
  NAND2_X1 U11544 ( .A1(n3219), .A2(n49453), .ZN(n51890) );
  NAND3_X1 U11673 ( .A1(n51835), .A2(n26503), .A3(n7601), .ZN(n26504) );
  NAND2_X1 U11709 ( .A1(n51791), .A2(n28152), .ZN(n51835) );
  NAND2_X1 U11716 ( .A1(n51837), .A2(n51836), .ZN(n21918) );
  NAND2_X1 U11727 ( .A1(n3488), .A2(n23509), .ZN(n21895) );
  NAND2_X1 U11729 ( .A1(n21897), .A2(n23504), .ZN(n51837) );
  INV_X1 U11742 ( .A(n39816), .ZN(n41331) );
  NAND2_X1 U11815 ( .A1(n41319), .A2(n4703), .ZN(n39816) );
  NAND4_X1 U11830 ( .A1(n41897), .A2(n39827), .A3(n39828), .A4(n39829), .ZN(
        n39849) );
  NAND3_X1 U11837 ( .A1(n39824), .A2(n4341), .A3(n4342), .ZN(n41897) );
  OR2_X1 U11842 ( .A1(n32503), .A2(n32507), .ZN(n30882) );
  NAND3_X1 U11893 ( .A1(n1730), .A2(n1729), .A3(n1734), .ZN(n52426) );
  NAND3_X1 U11947 ( .A1(n39697), .A2(n40835), .A3(n40143), .ZN(n37708) );
  NAND3_X1 U11955 ( .A1(n4598), .A2(n30292), .A3(n24880), .ZN(n24890) );
  OR2_X2 U11980 ( .A1(n3026), .A2(n20835), .ZN(n23955) );
  NOR2_X1 U11996 ( .A1(n1215), .A2(n51838), .ZN(n1213) );
  NAND2_X1 U12022 ( .A1(n30301), .A2(n30299), .ZN(n51838) );
  NAND3_X2 U12026 ( .A1(n5450), .A2(n39356), .A3(n51839), .ZN(n41997) );
  NAND3_X1 U12027 ( .A1(n39341), .A2(n51544), .A3(n39340), .ZN(n51839) );
  NAND2_X1 U12029 ( .A1(n12198), .A2(n13573), .ZN(n13577) );
  NAND2_X1 U12045 ( .A1(n41381), .A2(n41380), .ZN(n1237) );
  NAND2_X1 U12049 ( .A1(n35573), .A2(n38495), .ZN(n37521) );
  NAND2_X1 U12070 ( .A1(n1798), .A2(n2979), .ZN(n1920) );
  NAND3_X1 U12103 ( .A1(n32464), .A2(n32715), .A3(n32732), .ZN(n51840) );
  NAND3_X1 U12141 ( .A1(n46269), .A2(n46343), .A3(n46277), .ZN(n45240) );
  NAND2_X1 U12147 ( .A1(n32590), .A2(n32595), .ZN(n29621) );
  NAND3_X1 U12155 ( .A1(n51841), .A2(n6243), .A3(n51797), .ZN(n6240) );
  AND3_X4 U12172 ( .A1(n5877), .A2(n44260), .A3(n44259), .ZN(n48084) );
  NOR2_X1 U12204 ( .A1(n10968), .A2(n9855), .ZN(n10047) );
  INV_X1 U12208 ( .A(n22033), .ZN(n22315) );
  NOR2_X1 U12209 ( .A1(n18041), .A2(n15399), .ZN(n19423) );
  NAND3_X1 U12229 ( .A1(n42512), .A2(n45614), .A3(n46448), .ZN(n5521) );
  AND4_X4 U12231 ( .A1(n49260), .A2(n49258), .A3(n49257), .A4(n49259), .ZN(
        n49347) );
  NAND4_X1 U12232 ( .A1(n33008), .A2(n3487), .A3(n31383), .A4(n31385), .ZN(
        n33021) );
  OR2_X1 U12309 ( .A1(n24569), .A2(n51792), .ZN(n26889) );
  NAND4_X2 U12311 ( .A1(n32643), .A2(n32641), .A3(n32642), .A4(n32640), .ZN(
        n37324) );
  NOR2_X1 U12317 ( .A1(n40494), .A2(n51843), .ZN(n40498) );
  NAND2_X1 U12326 ( .A1(n40493), .A2(n41057), .ZN(n51843) );
  INV_X1 U12331 ( .A(n38677), .ZN(n38660) );
  NAND2_X1 U12332 ( .A1(n38241), .A2(n38670), .ZN(n38677) );
  NAND2_X1 U12339 ( .A1(n48526), .A2(n51844), .ZN(n48236) );
  NAND4_X4 U12342 ( .A1(n5179), .A2(n12528), .A3(n12530), .A4(n12529), .ZN(
        n15279) );
  OR2_X1 U12346 ( .A1(n41063), .A2(n41058), .ZN(n40513) );
  NAND2_X1 U12356 ( .A1(n32486), .A2(n32025), .ZN(n31205) );
  OAI211_X1 U12358 ( .C1(n11922), .C2(n11139), .A(n51846), .B(n51845), .ZN(
        n11140) );
  NAND2_X1 U12369 ( .A1(n11137), .A2(n357), .ZN(n51845) );
  NAND2_X1 U12374 ( .A1(n11368), .A2(n11367), .ZN(n8161) );
  OAI211_X1 U12375 ( .C1(n719), .C2(n29025), .A(n33034), .B(n29023), .ZN(n4438) );
  INV_X1 U12380 ( .A(n41206), .ZN(n51847) );
  NAND3_X1 U12383 ( .A1(n41196), .A2(n40032), .A3(n41195), .ZN(n41206) );
  NOR2_X1 U12391 ( .A1(n7389), .A2(n51848), .ZN(n7388) );
  OAI211_X1 U12402 ( .C1(n39383), .C2(n39384), .A(n51211), .B(n39382), .ZN(
        n51848) );
  AND2_X2 U12439 ( .A1(n442), .A2(n12536), .ZN(n12549) );
  XNOR2_X1 U12454 ( .A(n51849), .B(n47708), .ZN(Plaintext[17]) );
  NAND4_X1 U12455 ( .A1(n47705), .A2(n47706), .A3(n47704), .A4(n47707), .ZN(
        n51849) );
  XNOR2_X1 U12457 ( .A(n4995), .B(n33815), .ZN(n51850) );
  NAND2_X1 U12461 ( .A1(n51851), .A2(n46211), .ZN(n46221) );
  NAND3_X1 U12469 ( .A1(n46209), .A2(n52259), .A3(n51852), .ZN(n51851) );
  INV_X1 U12472 ( .A(n49218), .ZN(n51852) );
  NAND2_X1 U12517 ( .A1(n51854), .A2(n51853), .ZN(n4566) );
  NAND2_X1 U12523 ( .A1(n3469), .A2(n41377), .ZN(n51854) );
  NAND2_X1 U12547 ( .A1(n8937), .A2(n8938), .ZN(n8939) );
  NAND3_X1 U12580 ( .A1(n40639), .A2(n38816), .A3(n41796), .ZN(n8346) );
  NAND3_X1 U12583 ( .A1(n43333), .A2(n43332), .A3(n51855), .ZN(n43346) );
  NOR2_X1 U12588 ( .A1(n3273), .A2(n2354), .ZN(n27079) );
  NAND3_X1 U12599 ( .A1(n36917), .A2(n7644), .A3(n6089), .ZN(n6085) );
  NAND4_X2 U12632 ( .A1(n11223), .A2(n11221), .A3(n11222), .A4(n11220), .ZN(
        n14412) );
  NAND3_X2 U12644 ( .A1(n104), .A2(n4205), .A3(n3049), .ZN(n42209) );
  NAND3_X1 U12647 ( .A1(n9507), .A2(n11663), .A3(n9317), .ZN(n9312) );
  NAND3_X1 U12657 ( .A1(n51802), .A2(n51731), .A3(n49238), .ZN(n1252) );
  NAND2_X1 U12675 ( .A1(n49242), .A2(n49690), .ZN(n49233) );
  NAND2_X1 U12676 ( .A1(n12111), .A2(n10368), .ZN(n11372) );
  NAND3_X1 U12693 ( .A1(n30092), .A2(n31511), .A3(n31066), .ZN(n30094) );
  NAND2_X1 U12732 ( .A1(n32618), .A2(n31553), .ZN(n30323) );
  NOR2_X1 U12738 ( .A1(n7716), .A2(n51856), .ZN(n7710) );
  NAND2_X1 U12747 ( .A1(n21009), .A2(n51857), .ZN(n24017) );
  NAND2_X1 U12793 ( .A1(n51859), .A2(n51858), .ZN(n51857) );
  OR2_X2 U12813 ( .A1(n25113), .A2(n52231), .ZN(n32194) );
  NAND2_X1 U12846 ( .A1(n40676), .A2(n51860), .ZN(n36653) );
  NAND2_X1 U12847 ( .A1(n36650), .A2(n51800), .ZN(n51860) );
  NAND2_X2 U12859 ( .A1(n9694), .A2(n1073), .ZN(n13841) );
  INV_X1 U12860 ( .A(n36611), .ZN(n36612) );
  NAND2_X1 U12862 ( .A1(n34928), .A2(n8090), .ZN(n36611) );
  XNOR2_X1 U12864 ( .A(n51862), .B(n704), .ZN(n34826) );
  NAND3_X1 U12889 ( .A1(n23027), .A2(n23029), .A3(n23028), .ZN(n5034) );
  NAND3_X1 U12895 ( .A1(n3436), .A2(n48038), .A3(n650), .ZN(n44436) );
  OR2_X4 U12909 ( .A1(n5812), .A2(n8494), .ZN(n42441) );
  NAND2_X1 U12911 ( .A1(n36263), .A2(n51932), .ZN(n5812) );
  OR2_X1 U12946 ( .A1(n52147), .A2(n27918), .ZN(n25106) );
  NAND2_X1 U12950 ( .A1(n26927), .A2(n26928), .ZN(n26932) );
  NAND3_X1 U12962 ( .A1(n40533), .A2(n678), .A3(n1984), .ZN(n51271) );
  NAND2_X1 U12984 ( .A1(n26905), .A2(n29422), .ZN(n26731) );
  OAI21_X1 U12985 ( .B1(n30072), .B2(n30949), .A(n30071), .ZN(n30074) );
  NAND2_X1 U13000 ( .A1(n31117), .A2(n51863), .ZN(n30071) );
  NAND2_X1 U13003 ( .A1(n30944), .A2(n30945), .ZN(n31109) );
  NAND3_X1 U13004 ( .A1(n30063), .A2(n31115), .A3(n31106), .ZN(n30944) );
  XNOR2_X2 U13015 ( .A(n4592), .B(n16146), .ZN(n20052) );
  XNOR2_X1 U13037 ( .A(n51864), .B(n48757), .ZN(Plaintext[68]) );
  OAI21_X1 U13040 ( .B1(n48756), .B2(n48755), .A(n51865), .ZN(n51864) );
  NAND2_X1 U13049 ( .A1(n45949), .A2(n49138), .ZN(n43428) );
  NAND3_X1 U13050 ( .A1(n21548), .A2(n21547), .A3(n51129), .ZN(n21552) );
  NAND3_X1 U13051 ( .A1(n36572), .A2(n36490), .A3(n36491), .ZN(n6396) );
  XNOR2_X2 U13052 ( .A(n28069), .B(n27322), .ZN(n27467) );
  NAND4_X2 U13067 ( .A1(n22248), .A2(n22247), .A3(n22246), .A4(n22245), .ZN(
        n27322) );
  NOR2_X2 U13088 ( .A1(n3180), .A2(n22240), .ZN(n28069) );
  NOR2_X2 U13127 ( .A1(n7306), .A2(n42205), .ZN(n41934) );
  NAND2_X1 U13132 ( .A1(n39931), .A2(n40672), .ZN(n39930) );
  AND2_X2 U13135 ( .A1(n5746), .A2(n51866), .ZN(n33306) );
  NOR2_X1 U13149 ( .A1(n5745), .A2(n31200), .ZN(n51866) );
  NAND4_X1 U13153 ( .A1(n20868), .A2(n21758), .A3(n21755), .A4(n21756), .ZN(
        n21739) );
  NAND2_X1 U13159 ( .A1(n3062), .A2(n21744), .ZN(n20868) );
  NAND4_X2 U13185 ( .A1(n37954), .A2(n37955), .A3(n37952), .A4(n37953), .ZN(
        n43973) );
  NAND2_X1 U13193 ( .A1(n51867), .A2(n51777), .ZN(n7630) );
  NAND2_X1 U13232 ( .A1(n40487), .A2(n41118), .ZN(n51867) );
  NAND3_X1 U13251 ( .A1(n36555), .A2(n36556), .A3(n36554), .ZN(n51868) );
  NAND3_X2 U13252 ( .A1(n37034), .A2(n51869), .A3(n51799), .ZN(n41113) );
  NAND2_X1 U13276 ( .A1(n37036), .A2(n39369), .ZN(n51869) );
  NAND2_X1 U13318 ( .A1(n4840), .A2(n51870), .ZN(n49280) );
  OR2_X1 U13319 ( .A1(n49279), .A2(n49278), .ZN(n51870) );
  OAI21_X1 U13320 ( .B1(n39367), .B2(n51872), .A(n51871), .ZN(n8625) );
  NAND2_X1 U13325 ( .A1(n39367), .A2(n39375), .ZN(n51871) );
  NAND4_X1 U13329 ( .A1(n37357), .A2(n37358), .A3(n38436), .A4(n39560), .ZN(
        n4538) );
  NAND3_X1 U13344 ( .A1(n47653), .A2(n47654), .A3(n4223), .ZN(n47659) );
  NAND2_X1 U13349 ( .A1(n27881), .A2(n27875), .ZN(n27878) );
  NAND2_X1 U13351 ( .A1(n36471), .A2(n51873), .ZN(n36479) );
  NAND2_X1 U13352 ( .A1(n22250), .A2(n21861), .ZN(n4514) );
  NAND2_X1 U13359 ( .A1(n23318), .A2(n51875), .ZN(n22250) );
  NAND3_X1 U13381 ( .A1(n51876), .A2(n29366), .A3(n29368), .ZN(n29377) );
  NAND2_X1 U13398 ( .A1(n32232), .A2(n32257), .ZN(n51876) );
  NAND2_X1 U13405 ( .A1(n30173), .A2(n30174), .ZN(n30175) );
  NAND4_X2 U13417 ( .A1(n51765), .A2(n13265), .A3(n2990), .A4(n13264), .ZN(
        n17232) );
  OAI211_X1 U13433 ( .C1(n40830), .C2(n40826), .A(n51877), .B(n39081), .ZN(
        n39082) );
  NAND3_X1 U13436 ( .A1(n39079), .A2(n39078), .A3(n40822), .ZN(n51877) );
  NAND2_X1 U13449 ( .A1(n38272), .A2(n38282), .ZN(n2741) );
  NAND2_X1 U13486 ( .A1(n38043), .A2(n36372), .ZN(n38030) );
  NAND4_X2 U13489 ( .A1(n34531), .A2(n4416), .A3(n34526), .A4(n34530), .ZN(
        n41082) );
  OR2_X1 U13527 ( .A1(n51050), .A2(n16125), .ZN(n20616) );
  XNOR2_X2 U13544 ( .A(n35656), .B(n34504), .ZN(n34078) );
  AND4_X2 U13564 ( .A1(n1552), .A2(n1549), .A3(n31152), .A4(n1550), .ZN(n35656) );
  NAND3_X1 U13572 ( .A1(n41643), .A2(n41642), .A3(n41638), .ZN(n5090) );
  AOI21_X1 U13608 ( .B1(n50191), .B2(n50209), .A(n51878), .ZN(n50165) );
  AND2_X1 U13609 ( .A1(n50188), .A2(n7201), .ZN(n51878) );
  INV_X1 U13627 ( .A(n38828), .ZN(n51879) );
  NAND2_X1 U13631 ( .A1(n8150), .A2(n39754), .ZN(n39949) );
  NAND2_X1 U13650 ( .A1(n51880), .A2(n22251), .ZN(n3115) );
  NAND2_X1 U13658 ( .A1(n22254), .A2(n8303), .ZN(n51880) );
  NAND2_X1 U13713 ( .A1(n51125), .A2(n21873), .ZN(n22254) );
  NAND4_X4 U13716 ( .A1(n5321), .A2(n5437), .A3(n51881), .A4(n45555), .ZN(
        n48156) );
  MUX2_X1 U13723 ( .A(n31509), .B(n31071), .S(n31513), .Z(n51882) );
  NAND3_X1 U13725 ( .A1(n10787), .A2(n12546), .A3(n51883), .ZN(n10788) );
  NAND3_X1 U13726 ( .A1(n19665), .A2(n19666), .A3(n19667), .ZN(n19668) );
  NAND2_X1 U13750 ( .A1(n51884), .A2(n1080), .ZN(n47857) );
  NOR2_X1 U13813 ( .A1(n51886), .A2(n51885), .ZN(n51884) );
  NAND3_X1 U13815 ( .A1(n41813), .A2(n45191), .A3(n41812), .ZN(n51885) );
  OAI21_X1 U13843 ( .B1(n46555), .B2(n45810), .A(n41816), .ZN(n51886) );
  NAND3_X1 U13846 ( .A1(n51888), .A2(n5968), .A3(n51887), .ZN(n2918) );
  NAND2_X1 U13848 ( .A1(n46912), .A2(n45848), .ZN(n51887) );
  NAND2_X1 U13900 ( .A1(n46904), .A2(n45845), .ZN(n51888) );
  OR3_X1 U13901 ( .A1(n47827), .A2(n372), .A3(n47828), .ZN(n47833) );
  NAND2_X1 U13918 ( .A1(n933), .A2(n42104), .ZN(n51889) );
  NAND3_X1 U13920 ( .A1(n19499), .A2(n20078), .A3(n19491), .ZN(n19496) );
  OAI21_X1 U13940 ( .B1(n3220), .B2(n51890), .A(n49455), .ZN(n3216) );
  NAND2_X1 U13945 ( .A1(n40872), .A2(n51891), .ZN(n39525) );
  INV_X1 U13951 ( .A(n29773), .ZN(n29767) );
  XNOR2_X1 U13956 ( .A(n51892), .B(n46184), .ZN(Plaintext[133]) );
  NAND3_X1 U13992 ( .A1(n46182), .A2(n46183), .A3(n51276), .ZN(n51892) );
  NAND2_X1 U14023 ( .A1(n47396), .A2(n47397), .ZN(n50933) );
  NAND2_X1 U14048 ( .A1(n51894), .A2(n51893), .ZN(n3220) );
  NAND3_X1 U14059 ( .A1(n49435), .A2(n47195), .A3(n49449), .ZN(n51894) );
  NAND3_X2 U14077 ( .A1(n8412), .A2(n14892), .A3(n14897), .ZN(n18519) );
  NOR2_X2 U14094 ( .A1(n14894), .A2(n14895), .ZN(n8412) );
  NAND2_X1 U14191 ( .A1(n12363), .A2(n51769), .ZN(n10979) );
  NAND2_X1 U14214 ( .A1(n48703), .A2(n48674), .ZN(n48701) );
  NAND2_X1 U14219 ( .A1(n39361), .A2(n39386), .ZN(n51895) );
  BUF_X2 U14245 ( .A(n41675), .Z(n52198) );
  NAND3_X1 U14250 ( .A1(n13781), .A2(n13779), .A3(n13780), .ZN(n13784) );
  NAND2_X1 U14251 ( .A1(n788), .A2(n13173), .ZN(n13781) );
  OR2_X2 U14275 ( .A1(n51896), .A2(n8511), .ZN(n17117) );
  NAND4_X1 U14278 ( .A1(n10502), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n51896) );
  NAND2_X1 U14284 ( .A1(n52020), .A2(n51801), .ZN(n38444) );
  NOR2_X1 U14288 ( .A1(n23473), .A2(n23160), .ZN(n19589) );
  OR2_X2 U14314 ( .A1(n10061), .A2(n10062), .ZN(n13172) );
  NAND3_X1 U14331 ( .A1(n52322), .A2(n6399), .A3(n6400), .ZN(n6398) );
  NAND2_X1 U14332 ( .A1(n51897), .A2(n41925), .ZN(n41944) );
  NAND2_X1 U14380 ( .A1(n6617), .A2(n6980), .ZN(n51897) );
  NAND3_X1 U14388 ( .A1(n46448), .A2(n48449), .A3(n46446), .ZN(n46447) );
  NAND4_X1 U14393 ( .A1(n45706), .A2(n45704), .A3(n45707), .A4(n51898), .ZN(
        n51215) );
  AOI22_X1 U14406 ( .A1(n45703), .A2(n45702), .B1(n48873), .B2(n48915), .ZN(
        n51898) );
  NAND2_X1 U14407 ( .A1(n50455), .A2(n50454), .ZN(n7113) );
  INV_X1 U14471 ( .A(n45653), .ZN(n49167) );
  NAND4_X2 U14491 ( .A1(n22095), .A2(n22093), .A3(n51900), .A4(n51899), .ZN(
        n25493) );
  NAND2_X1 U14492 ( .A1(n22089), .A2(n22752), .ZN(n51899) );
  NAND2_X1 U14495 ( .A1(n22091), .A2(n22090), .ZN(n51901) );
  XNOR2_X1 U14517 ( .A(n51327), .B(n4613), .ZN(Plaintext[154]) );
  NAND3_X1 U14536 ( .A1(n21660), .A2(n20658), .A3(n20660), .ZN(n20272) );
  NAND3_X1 U14547 ( .A1(n21143), .A2(n21140), .A3(n6), .ZN(n23010) );
  NAND3_X1 U14581 ( .A1(n29153), .A2(n29154), .A3(n29155), .ZN(n29163) );
  NAND2_X1 U14584 ( .A1(n51902), .A2(n6488), .ZN(n3153) );
  OAI21_X1 U14585 ( .B1(n1432), .B2(n30257), .A(n1964), .ZN(n51902) );
  NAND2_X1 U14626 ( .A1(n51903), .A2(n29003), .ZN(n29004) );
  NAND3_X1 U14629 ( .A1(n28997), .A2(n4102), .A3(n30448), .ZN(n51903) );
  INV_X2 U14641 ( .A(n47674), .ZN(n47687) );
  NAND2_X1 U14653 ( .A1(n47651), .A2(n47674), .ZN(n47642) );
  AND4_X2 U14679 ( .A1(n45840), .A2(n45841), .A3(n45838), .A4(n45839), .ZN(
        n47674) );
  NAND2_X1 U14699 ( .A1(n7014), .A2(n23301), .ZN(n30783) );
  NAND3_X1 U14709 ( .A1(n27928), .A2(n27929), .A3(n27927), .ZN(n27935) );
  NAND3_X1 U14724 ( .A1(n48905), .A2(n5081), .A3(n48912), .ZN(n45700) );
  NOR2_X1 U14730 ( .A1(n28985), .A2(n51904), .ZN(n28986) );
  NAND2_X1 U14731 ( .A1(n28980), .A2(n28981), .ZN(n51904) );
  INV_X1 U14744 ( .A(n14681), .ZN(n15283) );
  NAND2_X1 U14745 ( .A1(n14962), .A2(n14950), .ZN(n14681) );
  NOR2_X1 U14751 ( .A1(n51905), .A2(n24269), .ZN(n20172) );
  OAI21_X1 U14771 ( .B1(n23424), .B2(n23425), .A(n20170), .ZN(n24269) );
  AND2_X1 U14794 ( .A1(n24266), .A2(n20171), .ZN(n51905) );
  OAI21_X1 U14801 ( .B1(n51907), .B2(n51906), .A(n19887), .ZN(n52281) );
  INV_X1 U14808 ( .A(n18935), .ZN(n51907) );
  INV_X1 U14862 ( .A(n11794), .ZN(n13049) );
  NAND3_X1 U14880 ( .A1(n44623), .A2(n44621), .A3(n44622), .ZN(n44637) );
  NAND2_X1 U14894 ( .A1(n27829), .A2(n29438), .ZN(n27827) );
  NAND2_X1 U14917 ( .A1(n5589), .A2(n5587), .ZN(n3261) );
  NAND3_X1 U14922 ( .A1(n36543), .A2(n36544), .A3(n51908), .ZN(n36546) );
  NAND2_X1 U14938 ( .A1(n51077), .A2(n51909), .ZN(n51908) );
  NAND2_X2 U14944 ( .A1(n770), .A2(n19518), .ZN(n21232) );
  NOR2_X1 U14945 ( .A1(n47876), .A2(n51911), .ZN(n47816) );
  NAND3_X1 U14948 ( .A1(n47883), .A2(n47873), .A3(n51941), .ZN(n51911) );
  XNOR2_X1 U14966 ( .A(n51912), .B(n34737), .ZN(n34740) );
  XNOR2_X1 U14967 ( .A(n34736), .B(n34735), .ZN(n51912) );
  NAND2_X1 U14971 ( .A1(n51123), .A2(n23157), .ZN(n23466) );
  NAND3_X1 U14988 ( .A1(n51913), .A2(n3984), .A3(n33163), .ZN(n36998) );
  NAND2_X1 U15006 ( .A1(n52389), .A2(n33154), .ZN(n51913) );
  INV_X2 U15030 ( .A(n32879), .ZN(n719) );
  NAND2_X1 U15051 ( .A1(n32879), .A2(n51914), .ZN(n29023) );
  INV_X1 U15053 ( .A(n29026), .ZN(n51914) );
  AND3_X2 U15067 ( .A1(n28986), .A2(n28987), .A3(n28988), .ZN(n32879) );
  XNOR2_X1 U15073 ( .A(n51915), .B(n50450), .ZN(Plaintext[153]) );
  NAND3_X1 U15079 ( .A1(n50449), .A2(n50448), .A3(n4690), .ZN(n51915) );
  OAI21_X1 U15106 ( .B1(n45698), .B2(n46360), .A(n657), .ZN(n51916) );
  NAND4_X4 U15107 ( .A1(n11038), .A2(n11039), .A3(n11040), .A4(n51917), .ZN(
        n13729) );
  NOR2_X2 U15108 ( .A1(n11034), .A2(n8641), .ZN(n51917) );
  NAND3_X1 U15123 ( .A1(n52029), .A2(n45881), .A3(n45882), .ZN(n51602) );
  OR3_X1 U15139 ( .A1(n35214), .A2(n35215), .A3(n36045), .ZN(n36584) );
  NAND3_X1 U15145 ( .A1(n7056), .A2(n7058), .A3(n46529), .ZN(n6639) );
  NAND2_X1 U15151 ( .A1(n4933), .A2(n50), .ZN(n19180) );
  NAND3_X2 U15157 ( .A1(n46470), .A2(n46468), .A3(n46469), .ZN(n48703) );
  NOR2_X2 U15158 ( .A1(n3668), .A2(n51919), .ZN(n7351) );
  NAND4_X1 U15161 ( .A1(n5310), .A2(n1522), .A3(n1523), .A4(n17992), .ZN(
        n51919) );
  NAND3_X1 U15184 ( .A1(n5743), .A2(n30168), .A3(n30167), .ZN(n102) );
  NAND2_X1 U15185 ( .A1(n37593), .A2(n37378), .ZN(n36222) );
  XNOR2_X2 U15187 ( .A(n45), .B(n33714), .ZN(n37378) );
  INV_X1 U15191 ( .A(n51920), .ZN(n30745) );
  OAI211_X1 U15229 ( .C1(n52173), .C2(n30737), .A(n30735), .B(n30736), .ZN(
        n51920) );
  OAI21_X1 U15243 ( .B1(n2425), .B2(n40146), .A(n40159), .ZN(n5771) );
  NAND3_X1 U15281 ( .A1(n37468), .A2(n40549), .A3(n40567), .ZN(n40146) );
  NAND3_X1 U15311 ( .A1(n27852), .A2(n26677), .A3(n26676), .ZN(n27863) );
  NAND2_X1 U15330 ( .A1(n8276), .A2(n8743), .ZN(n30322) );
  XNOR2_X1 U15341 ( .A(n51921), .B(n41253), .ZN(n41470) );
  XNOR2_X1 U15346 ( .A(n41252), .B(n41254), .ZN(n51921) );
  NAND3_X1 U15349 ( .A1(n25052), .A2(n25053), .A3(n51922), .ZN(n24904) );
  NOR2_X1 U15357 ( .A1(n51924), .A2(n51923), .ZN(n51922) );
  INV_X1 U15360 ( .A(n25061), .ZN(n51924) );
  NAND3_X2 U15368 ( .A1(n35450), .A2(n35449), .A3(n51925), .ZN(n40316) );
  NOR2_X1 U15370 ( .A1(n51778), .A2(n51779), .ZN(n51925) );
  AND2_X2 U15381 ( .A1(n46595), .A2(n45790), .ZN(n46705) );
  NAND4_X4 U15384 ( .A1(n1722), .A2(n6523), .A3(n1721), .A4(n7127), .ZN(n47989) );
  NAND2_X1 U15416 ( .A1(n35893), .A2(n51926), .ZN(n35897) );
  AOI21_X1 U15422 ( .B1(n6615), .B2(n38345), .A(n6614), .ZN(n51926) );
  NAND2_X1 U15423 ( .A1(n18944), .A2(n51928), .ZN(n18945) );
  NAND2_X1 U15433 ( .A1(n14398), .A2(n14394), .ZN(n14396) );
  NAND2_X1 U15439 ( .A1(n14408), .A2(n14393), .ZN(n14398) );
  NAND2_X1 U15463 ( .A1(n10328), .A2(n12161), .ZN(n11330) );
  NAND3_X1 U15466 ( .A1(n22642), .A2(n17419), .A3(n51929), .ZN(n17423) );
  NAND2_X1 U15490 ( .A1(n23066), .A2(n51930), .ZN(n51929) );
  NAND2_X1 U15529 ( .A1(n50542), .A2(n50553), .ZN(n50548) );
  NAND2_X1 U15564 ( .A1(n38018), .A2(n5872), .ZN(n38007) );
  NAND2_X1 U15565 ( .A1(n51931), .A2(n38566), .ZN(n5503) );
  NAND2_X1 U15566 ( .A1(n35147), .A2(n5505), .ZN(n51931) );
  INV_X1 U15570 ( .A(n19721), .ZN(n19799) );
  NAND3_X1 U15580 ( .A1(n26329), .A2(n25839), .A3(n25838), .ZN(n51981) );
  NOR2_X1 U15603 ( .A1(n52367), .A2(n52366), .ZN(n51932) );
  NAND2_X1 U15620 ( .A1(n39335), .A2(n37782), .ZN(n39336) );
  NAND2_X1 U15678 ( .A1(n9539), .A2(n9542), .ZN(n12611) );
  NAND2_X1 U15679 ( .A1(n16803), .A2(n16804), .ZN(n16806) );
  NAND2_X2 U15698 ( .A1(n37185), .A2(n37186), .ZN(n40456) );
  NAND3_X1 U15704 ( .A1(n4278), .A2(n46221), .A3(n46218), .ZN(n46238) );
  NAND3_X1 U15710 ( .A1(n24040), .A2(n24038), .A3(n24039), .ZN(n2069) );
  NOR2_X1 U15730 ( .A1(n48258), .A2(n51766), .ZN(n48266) );
  XNOR2_X1 U15738 ( .A(n51933), .B(n47244), .ZN(Plaintext[186]) );
  NAND4_X1 U15748 ( .A1(n47242), .A2(n47240), .A3(n47241), .A4(n47243), .ZN(
        n51933) );
  NAND3_X1 U15749 ( .A1(n18012), .A2(n17574), .A3(n51934), .ZN(n17583) );
  NAND2_X1 U15759 ( .A1(n51935), .A2(n10527), .ZN(n10534) );
  NAND2_X1 U15762 ( .A1(n10632), .A2(n51782), .ZN(n51935) );
  NAND2_X1 U15767 ( .A1(n9836), .A2(n10513), .ZN(n10632) );
  NOR2_X1 U15776 ( .A1(n5307), .A2(n51936), .ZN(n4975) );
  NAND3_X1 U15817 ( .A1(n31863), .A2(n32157), .A3(n32778), .ZN(n32291) );
  NOR2_X1 U15829 ( .A1(n29114), .A2(n51937), .ZN(n29118) );
  OAI22_X1 U15837 ( .A1(n29239), .A2(n29226), .B1(n625), .B2(n30267), .ZN(
        n51937) );
  NAND3_X1 U15861 ( .A1(n49278), .A2(n45668), .A3(n46196), .ZN(n44776) );
  NAND2_X1 U15871 ( .A1(n51938), .A2(n28803), .ZN(n3622) );
  NAND3_X1 U15881 ( .A1(n5638), .A2(n28800), .A3(n28799), .ZN(n51938) );
  NAND2_X1 U15885 ( .A1(n19725), .A2(n17405), .ZN(n21214) );
  NAND4_X2 U15906 ( .A1(n51939), .A2(n13892), .A3(n13891), .A4(n13889), .ZN(
        n18193) );
  NAND2_X1 U15934 ( .A1(n1319), .A2(n19824), .ZN(n1318) );
  NOR2_X2 U15960 ( .A1(n8437), .A2(n2640), .ZN(n51023) );
  NAND3_X1 U15962 ( .A1(n3545), .A2(n49819), .A3(n49815), .ZN(n3544) );
  NAND3_X1 U15972 ( .A1(n47819), .A2(n47818), .A3(n51940), .ZN(n47820) );
  NAND2_X1 U15974 ( .A1(n51285), .A2(n51941), .ZN(n51940) );
  XNOR2_X1 U15975 ( .A(n33866), .B(n33865), .ZN(n51942) );
  NAND3_X1 U15976 ( .A1(n31002), .A2(n31001), .A3(n31000), .ZN(n8044) );
  NAND3_X1 U15979 ( .A1(n51943), .A2(n10416), .A3(n10415), .ZN(n6151) );
  NAND3_X1 U15980 ( .A1(n3451), .A2(n10420), .A3(n10421), .ZN(n51943) );
  AOI22_X2 U15993 ( .A1(n29938), .A2(n28751), .B1(n28750), .B2(n28752), .ZN(
        n28763) );
  NAND2_X1 U16000 ( .A1(n1604), .A2(n39787), .ZN(n37360) );
  NAND3_X1 U16005 ( .A1(n19512), .A2(n19511), .A3(n51944), .ZN(n19515) );
  OR2_X1 U16014 ( .A1(n19513), .A2(n21233), .ZN(n51944) );
  INV_X1 U16017 ( .A(n35579), .ZN(n35578) );
  NAND2_X1 U16020 ( .A1(n37520), .A2(n38494), .ZN(n35579) );
  NAND3_X1 U16028 ( .A1(n50730), .A2(n7745), .A3(n7746), .ZN(n7739) );
  NAND3_X1 U16030 ( .A1(n50720), .A2(n50718), .A3(n50719), .ZN(n50730) );
  XNOR2_X1 U16049 ( .A(n51945), .B(n42815), .ZN(Plaintext[89]) );
  NAND3_X1 U16129 ( .A1(n30), .A2(n42814), .A3(n42813), .ZN(n51945) );
  OAI21_X1 U16130 ( .B1(n25106), .B2(n30272), .A(n29240), .ZN(n25108) );
  NAND2_X1 U16131 ( .A1(n51978), .A2(n51259), .ZN(n5189) );
  OAI21_X1 U16136 ( .B1(n17470), .B2(n19427), .A(n17867), .ZN(n17473) );
  NAND2_X1 U16144 ( .A1(n19411), .A2(n51946), .ZN(n17867) );
  NAND2_X1 U16155 ( .A1(n38955), .A2(n51947), .ZN(n5142) );
  NAND2_X1 U16167 ( .A1(n247), .A2(n248), .ZN(n51947) );
  INV_X1 U16176 ( .A(n32525), .ZN(n31835) );
  NAND2_X1 U16177 ( .A1(n6042), .A2(n32962), .ZN(n32525) );
  NAND3_X1 U16219 ( .A1(n16993), .A2(n4710), .A3(n20983), .ZN(n4709) );
  NAND3_X1 U16221 ( .A1(n25110), .A2(n25111), .A3(n25109), .ZN(n52231) );
  NAND2_X1 U16237 ( .A1(n9429), .A2(n9433), .ZN(n12137) );
  NAND2_X1 U16249 ( .A1(n14331), .A2(n14344), .ZN(n51948) );
  NAND3_X1 U16266 ( .A1(n615), .A2(n36252), .A3(n37762), .ZN(n35915) );
  NAND3_X1 U16271 ( .A1(n40351), .A2(n40349), .A3(n40350), .ZN(n5125) );
  NAND3_X1 U16280 ( .A1(n42807), .A2(n1255), .A3(n1256), .ZN(n4259) );
  NAND3_X1 U16291 ( .A1(n22238), .A2(n22237), .A3(n22239), .ZN(n3180) );
  OR2_X2 U16303 ( .A1(n51949), .A2(n52386), .ZN(n24332) );
  OR2_X1 U16324 ( .A1(n20644), .A2(n20645), .ZN(n51949) );
  NAND2_X1 U16325 ( .A1(n32486), .A2(n32484), .ZN(n32014) );
  NAND2_X1 U16331 ( .A1(n48744), .A2(n48760), .ZN(n48736) );
  NAND2_X1 U16400 ( .A1(n27620), .A2(n27719), .ZN(n1162) );
  NAND2_X1 U16407 ( .A1(n48269), .A2(n48268), .ZN(n48261) );
  NAND2_X1 U16418 ( .A1(n51951), .A2(n51775), .ZN(n39329) );
  NAND2_X1 U16428 ( .A1(n43667), .A2(n40633), .ZN(n51951) );
  OAI21_X1 U16452 ( .B1(n35171), .B2(n38551), .A(n35180), .ZN(n51952) );
  OAI21_X1 U16456 ( .B1(n27147), .B2(n27148), .A(n51781), .ZN(n27151) );
  OR2_X2 U16462 ( .A1(n473), .A2(n7159), .ZN(n37802) );
  NAND4_X4 U16466 ( .A1(n14461), .A2(n14462), .A3(n14459), .A4(n14460), .ZN(
        n17763) );
  AOI22_X1 U16473 ( .A1(n728), .A2(n29704), .B1(n29705), .B2(n29707), .ZN(
        n29710) );
  NAND3_X1 U16489 ( .A1(n50606), .A2(n50605), .A3(n50604), .ZN(n50608) );
  NAND3_X1 U16497 ( .A1(n19423), .A2(n17469), .A3(n19424), .ZN(n19429) );
  NAND2_X1 U16534 ( .A1(n48762), .A2(n52067), .ZN(n1933) );
  NAND3_X1 U16538 ( .A1(n19073), .A2(n16804), .A3(n1418), .ZN(n17071) );
  NAND2_X1 U16549 ( .A1(n1415), .A2(n19066), .ZN(n19073) );
  NAND2_X2 U16569 ( .A1(n1086), .A2(n29787), .ZN(n32716) );
  NAND4_X2 U16595 ( .A1(n8672), .A2(n41592), .A3(n41591), .A4(n8671), .ZN(
        n44535) );
  NAND3_X1 U16600 ( .A1(n22012), .A2(n22593), .A3(n22011), .ZN(n22013) );
  NAND2_X1 U16601 ( .A1(n11268), .A2(n9974), .ZN(n11686) );
  OAI22_X1 U16611 ( .A1(n44727), .A2(n46299), .B1(n49150), .B2(n49138), .ZN(
        n44728) );
  AND2_X2 U16644 ( .A1(n43427), .A2(n51017), .ZN(n49148) );
  XNOR2_X1 U16654 ( .A(n51953), .B(n50759), .ZN(Plaintext[175]) );
  NAND4_X1 U16691 ( .A1(n50757), .A2(n50756), .A3(n50758), .A4(n50755), .ZN(
        n51953) );
  NAND2_X1 U16714 ( .A1(n20221), .A2(n51006), .ZN(n19693) );
  NAND2_X1 U16719 ( .A1(n36137), .A2(n3211), .ZN(n38582) );
  NAND3_X2 U16725 ( .A1(n31505), .A2(n31506), .A3(n51794), .ZN(n34553) );
  NAND2_X1 U16734 ( .A1(n47109), .A2(n47111), .ZN(n7918) );
  XNOR2_X2 U16737 ( .A(n17389), .B(n16660), .ZN(n18696) );
  XNOR2_X1 U16788 ( .A(n1778), .B(n27197), .ZN(n51955) );
  NAND3_X1 U16808 ( .A1(n23556), .A2(n23555), .A3(n23554), .ZN(n23558) );
  NAND2_X1 U16809 ( .A1(n39271), .A2(n39014), .ZN(n39286) );
  NAND2_X1 U16823 ( .A1(n45928), .A2(n51957), .ZN(n44779) );
  NAND2_X1 U16851 ( .A1(n49265), .A2(n45668), .ZN(n45928) );
  INV_X1 U16864 ( .A(n51126), .ZN(n52401) );
  NAND2_X1 U16865 ( .A1(n28637), .A2(n51958), .ZN(n27817) );
  NAND3_X1 U16867 ( .A1(n13760), .A2(n13125), .A3(n13761), .ZN(n13126) );
  NOR2_X1 U16868 ( .A1(n2556), .A2(n13124), .ZN(n13760) );
  XNOR2_X2 U16880 ( .A(n51959), .B(n52022), .ZN(n30393) );
  XNOR2_X1 U16881 ( .A(n24054), .B(n7934), .ZN(n51959) );
  NAND2_X1 U16885 ( .A1(n6019), .A2(n12054), .ZN(n12056) );
  NAND2_X1 U16921 ( .A1(n32232), .A2(n51961), .ZN(n32235) );
  OAI21_X1 U16922 ( .B1(n51962), .B2(n1296), .A(n19283), .ZN(n6432) );
  NAND2_X1 U16926 ( .A1(n19274), .A2(n19275), .ZN(n51962) );
  OAI21_X1 U16931 ( .B1(n49739), .B2(n51963), .A(n49738), .ZN(n49746) );
  NAND4_X1 U16932 ( .A1(n43419), .A2(n43417), .A3(n43413), .A4(n43414), .ZN(
        n3962) );
  AOI21_X1 U16980 ( .B1(n20958), .B2(n22154), .A(n20957), .ZN(n20960) );
  NOR2_X1 U16983 ( .A1(n3423), .A2(n50992), .ZN(n20958) );
  NAND2_X1 U16985 ( .A1(n15054), .A2(n51964), .ZN(n13478) );
  NAND2_X1 U16991 ( .A1(n51967), .A2(n51966), .ZN(n51965) );
  INV_X1 U17048 ( .A(n13797), .ZN(n51967) );
  NAND2_X1 U17064 ( .A1(n30058), .A2(n52121), .ZN(n30941) );
  AOI21_X1 U17072 ( .B1(n51970), .B2(n51969), .A(n51968), .ZN(n9935) );
  INV_X1 U17147 ( .A(n9933), .ZN(n51970) );
  NAND2_X1 U17148 ( .A1(n12523), .A2(n51971), .ZN(n11262) );
  NAND3_X1 U17182 ( .A1(n13257), .A2(n12028), .A3(n7245), .ZN(n12029) );
  NAND3_X1 U17245 ( .A1(n49275), .A2(n49278), .A3(n46199), .ZN(n7212) );
  INV_X2 U17247 ( .A(n48888), .ZN(n48905) );
  NAND4_X2 U17249 ( .A1(n3592), .A2(n2306), .A3(n3632), .A4(n45691), .ZN(
        n48888) );
  AND2_X2 U17250 ( .A1(n45697), .A2(n46267), .ZN(n46344) );
  NAND2_X1 U17255 ( .A1(n39553), .A2(n40125), .ZN(n40195) );
  BUF_X2 U17307 ( .A(n47599), .Z(n2163) );
  NAND3_X1 U17312 ( .A1(n1739), .A2(n1742), .A3(n36650), .ZN(n40686) );
  NOR2_X1 U17334 ( .A1(n1288), .A2(n1289), .ZN(n1739) );
  AND4_X2 U17342 ( .A1(n7486), .A2(n9152), .A3(n9150), .A4(n9151), .ZN(n14644)
         );
  AND3_X1 U17358 ( .A1(n2651), .A2(n2646), .A3(n2649), .ZN(n52417) );
  NAND2_X1 U17406 ( .A1(n19896), .A2(n18932), .ZN(n19898) );
  NAND2_X1 U17417 ( .A1(n51973), .A2(n51972), .ZN(n40093) );
  NAND2_X1 U17438 ( .A1(n40085), .A2(n40903), .ZN(n51973) );
  NAND2_X1 U17479 ( .A1(n27917), .A2(n51974), .ZN(n27920) );
  OAI21_X1 U17480 ( .B1(n51372), .B2(n50277), .A(n51975), .ZN(n47040) );
  NAND2_X1 U17495 ( .A1(n50277), .A2(n47333), .ZN(n51975) );
  NAND3_X1 U17496 ( .A1(n5337), .A2(n9069), .A3(n9070), .ZN(n6435) );
  INV_X1 U17510 ( .A(n32868), .ZN(n51976) );
  NAND2_X1 U17523 ( .A1(n32879), .A2(n8544), .ZN(n32868) );
  NAND2_X1 U17525 ( .A1(n20320), .A2(n20321), .ZN(n20324) );
  NAND3_X1 U17529 ( .A1(n21559), .A2(n5167), .A3(n21578), .ZN(n21576) );
  NAND2_X1 U17530 ( .A1(n46987), .A2(n46988), .ZN(n46991) );
  OAI21_X1 U17573 ( .B1(n48085), .B2(n48084), .A(n48005), .ZN(n3436) );
  NAND2_X1 U17591 ( .A1(n48020), .A2(n3075), .ZN(n48005) );
  NAND2_X1 U17603 ( .A1(n5937), .A2(n43427), .ZN(n43429) );
  NAND2_X1 U17639 ( .A1(n45944), .A2(n44733), .ZN(n5937) );
  NAND2_X1 U17652 ( .A1(n7348), .A2(n35988), .ZN(n7349) );
  NAND2_X1 U17668 ( .A1(n51977), .A2(n47989), .ZN(n47979) );
  INV_X1 U17711 ( .A(n47991), .ZN(n51977) );
  OR2_X1 U17766 ( .A1(n49683), .A2(n49232), .ZN(n49250) );
  NOR2_X1 U17773 ( .A1(n13302), .A2(n13728), .ZN(n51978) );
  NAND3_X1 U17779 ( .A1(n14295), .A2(n5411), .A3(n14287), .ZN(n13586) );
  NAND3_X1 U17780 ( .A1(n47211), .A2(n47265), .A3(n47617), .ZN(n47213) );
  XNOR2_X1 U17787 ( .A(n51979), .B(n49612), .ZN(Plaintext[125]) );
  NAND2_X1 U17789 ( .A1(n6007), .A2(n6006), .ZN(n51979) );
  XNOR2_X2 U17805 ( .A(n4591), .B(n33683), .ZN(n36200) );
  OAI21_X1 U17808 ( .B1(n50938), .B2(n50937), .A(n50958), .ZN(n50939) );
  NAND2_X1 U17812 ( .A1(n23640), .A2(n23639), .ZN(n51980) );
  NAND2_X1 U17818 ( .A1(n51981), .A2(n26677), .ZN(n25846) );
  NAND3_X1 U17820 ( .A1(n30452), .A2(n29748), .A3(n29000), .ZN(n28832) );
  NAND2_X1 U17824 ( .A1(n51983), .A2(n51982), .ZN(n15394) );
  NAND2_X1 U17840 ( .A1(n15370), .A2(n7735), .ZN(n51982) );
  NAND2_X1 U17885 ( .A1(n15371), .A2(n51984), .ZN(n51983) );
  OAI21_X1 U17921 ( .B1(n51985), .B2(n45153), .A(n4780), .ZN(n45169) );
  INV_X1 U17931 ( .A(n2708), .ZN(n51985) );
  NAND3_X2 U17937 ( .A1(n8858), .A2(n7687), .A3(n8859), .ZN(n14294) );
  NAND2_X1 U17938 ( .A1(n20328), .A2(n21426), .ZN(n3491) );
  NOR2_X1 U17945 ( .A1(n31793), .A2(n31792), .ZN(n31027) );
  NAND2_X1 U17949 ( .A1(n5912), .A2(n31886), .ZN(n31793) );
  NAND4_X1 U17977 ( .A1(n31470), .A2(n31471), .A3(n51471), .A4(n32609), .ZN(
        n8743) );
  NAND3_X1 U18005 ( .A1(n31770), .A2(n30890), .A3(n30889), .ZN(n30891) );
  XNOR2_X1 U18016 ( .A(n51986), .B(n19258), .ZN(n19277) );
  XNOR2_X1 U18022 ( .A(n19257), .B(n19256), .ZN(n51986) );
  NAND2_X1 U18035 ( .A1(n23871), .A2(n51987), .ZN(n23874) );
  INV_X1 U18048 ( .A(n23869), .ZN(n51987) );
  NAND2_X1 U18050 ( .A1(n23756), .A2(n22605), .ZN(n23869) );
  NAND2_X1 U18057 ( .A1(n51988), .A2(n10127), .ZN(n10956) );
  XNOR2_X2 U18095 ( .A(n7140), .B(Key[173]), .ZN(n10127) );
  INV_X1 U18108 ( .A(n13952), .ZN(n13946) );
  NAND2_X1 U18110 ( .A1(n12882), .A2(n13941), .ZN(n13952) );
  NOR2_X1 U18123 ( .A1(n51774), .A2(n51989), .ZN(n18366) );
  OAI21_X1 U18178 ( .B1(n18360), .B2(n19065), .A(n18358), .ZN(n51989) );
  INV_X1 U18192 ( .A(n39077), .ZN(n51990) );
  NOR2_X1 U18200 ( .A1(n51992), .A2(n23868), .ZN(n51991) );
  OAI21_X1 U18254 ( .B1(n47217), .B2(n52226), .A(n50622), .ZN(n51994) );
  NAND2_X1 U18260 ( .A1(n46395), .A2(n46488), .ZN(n46392) );
  XNOR2_X2 U18316 ( .A(n42796), .B(n42797), .ZN(n46488) );
  AND2_X2 U18318 ( .A1(n18873), .A2(n20683), .ZN(n20672) );
  NAND2_X1 U18342 ( .A1(n20467), .A2(n8232), .ZN(n20384) );
  NAND3_X1 U18349 ( .A1(n1789), .A2(n51130), .A3(n20473), .ZN(n20467) );
  NAND2_X1 U18414 ( .A1(n7916), .A2(n36632), .ZN(n36320) );
  NAND2_X1 U18418 ( .A1(n30711), .A2(n27164), .ZN(n30707) );
  INV_X1 U18460 ( .A(n40510), .ZN(n40514) );
  NAND2_X1 U18461 ( .A1(n49113), .A2(n49054), .ZN(n49107) );
  AND3_X2 U18462 ( .A1(n51995), .A2(n34967), .A3(n34968), .ZN(n41054) );
  INV_X1 U18524 ( .A(n9558), .ZN(n11976) );
  NAND2_X1 U18532 ( .A1(n11986), .A2(n10444), .ZN(n9558) );
  NAND3_X1 U18543 ( .A1(n2786), .A2(n2785), .A3(n38279), .ZN(n2781) );
  NAND2_X1 U18547 ( .A1(n23020), .A2(n23021), .ZN(n22851) );
  NAND4_X2 U18563 ( .A1(n19385), .A2(n19379), .A3(n5862), .A4(n51562), .ZN(
        n22856) );
  OAI21_X1 U18580 ( .B1(n14127), .B2(n14126), .A(n14125), .ZN(n51277) );
  NAND3_X1 U18581 ( .A1(n1686), .A2(n24271), .A3(n24270), .ZN(n26093) );
  XNOR2_X1 U18582 ( .A(n51996), .B(n26050), .ZN(n5020) );
  XNOR2_X1 U18663 ( .A(n26049), .B(n26051), .ZN(n51996) );
  NAND3_X1 U18665 ( .A1(n48749), .A2(n48762), .A3(n48730), .ZN(n48721) );
  NAND2_X1 U18674 ( .A1(n51998), .A2(n51997), .ZN(n46377) );
  NAND2_X1 U18730 ( .A1(n48538), .A2(n46462), .ZN(n51998) );
  NAND4_X2 U18732 ( .A1(n3471), .A2(n4764), .A3(n40266), .A4(n42142), .ZN(
        n50987) );
  INV_X1 U18737 ( .A(n12321), .ZN(n12334) );
  NAND3_X1 U18745 ( .A1(n12342), .A2(n12322), .A3(n51999), .ZN(n4351) );
  AND2_X1 U18759 ( .A1(n52199), .A2(n12321), .ZN(n51999) );
  NAND2_X1 U18847 ( .A1(n12336), .A2(n10669), .ZN(n12321) );
  NAND2_X1 U18864 ( .A1(n9476), .A2(n10065), .ZN(n9921) );
  NAND2_X1 U18865 ( .A1(n463), .A2(n22184), .ZN(n21095) );
  NAND3_X1 U18874 ( .A1(n21178), .A2(n19702), .A3(n21181), .ZN(n19700) );
  NAND2_X1 U18911 ( .A1(n27786), .A2(n27788), .ZN(n27787) );
  NAND4_X1 U18928 ( .A1(n899), .A2(n5565), .A3(n39420), .A4(n52000), .ZN(n897)
         );
  NAND2_X1 U18934 ( .A1(n40259), .A2(n52001), .ZN(n4763) );
  INV_X1 U18940 ( .A(n42149), .ZN(n52001) );
  NOR2_X2 U18944 ( .A1(n42154), .A2(n41770), .ZN(n42149) );
  NAND2_X1 U18948 ( .A1(n22575), .A2(n24026), .ZN(n22576) );
  XNOR2_X1 U18973 ( .A(n42248), .B(n52002), .ZN(n52325) );
  XNOR2_X1 U19004 ( .A(n42247), .B(n45317), .ZN(n52002) );
  NAND2_X1 U19019 ( .A1(n8042), .A2(n8043), .ZN(n8041) );
  NAND2_X1 U19077 ( .A1(n45804), .A2(n46730), .ZN(n45189) );
  OR2_X2 U19101 ( .A1(n22544), .A2(n22543), .ZN(n23178) );
  NAND2_X1 U19124 ( .A1(n48667), .A2(n47407), .ZN(n46530) );
  INV_X1 U19178 ( .A(n48702), .ZN(n52004) );
  AOI21_X1 U19189 ( .B1(n20390), .B2(n52005), .A(n51776), .ZN(n20402) );
  NAND2_X1 U19192 ( .A1(n10984), .A2(n10983), .ZN(n52006) );
  OR2_X1 U19226 ( .A1(n12359), .A2(n9780), .ZN(n10984) );
  NAND2_X1 U19227 ( .A1(n10985), .A2(n52008), .ZN(n52007) );
  INV_X1 U19235 ( .A(n10983), .ZN(n52008) );
  NAND3_X1 U19250 ( .A1(n46491), .A2(n46488), .A3(n46487), .ZN(n46490) );
  NAND3_X1 U19305 ( .A1(n52009), .A2(n21987), .A3(n2130), .ZN(n4277) );
  INV_X1 U19316 ( .A(n21991), .ZN(n52009) );
  NAND2_X2 U19317 ( .A1(n52010), .A2(n16894), .ZN(n24287) );
  AND3_X1 U19330 ( .A1(n16895), .A2(n3268), .A3(n16893), .ZN(n52010) );
  NAND2_X1 U19331 ( .A1(n24283), .A2(n21900), .ZN(n3100) );
  AOI22_X1 U19360 ( .A1(n32360), .A2(n32347), .B1(n32455), .B2(n32441), .ZN(
        n32058) );
  NAND2_X1 U19402 ( .A1(n35211), .A2(n35875), .ZN(n6129) );
  NAND2_X1 U19426 ( .A1(n12668), .A2(n12669), .ZN(n12670) );
  NAND3_X1 U19428 ( .A1(n38851), .A2(n37870), .A3(n52011), .ZN(n37872) );
  OR2_X2 U19439 ( .A1(n37283), .A2(n38701), .ZN(n39240) );
  XNOR2_X2 U19442 ( .A(n37248), .B(n37249), .ZN(n38701) );
  AOI22_X1 U19450 ( .A1(n39442), .A2(n39443), .B1(n52012), .B2(n39441), .ZN(
        n39459) );
  NOR2_X1 U19454 ( .A1(n39439), .A2(n39438), .ZN(n52012) );
  XNOR2_X1 U19474 ( .A(n8757), .B(n41881), .ZN(n52013) );
  XNOR2_X1 U19481 ( .A(n52014), .B(n50431), .ZN(Plaintext[152]) );
  NAND3_X1 U19502 ( .A1(n50428), .A2(n50430), .A3(n52015), .ZN(n52014) );
  NOR2_X2 U19504 ( .A1(n49606), .A2(n49579), .ZN(n49600) );
  NAND2_X1 U19507 ( .A1(n23986), .A2(n23982), .ZN(n22428) );
  AND2_X2 U19531 ( .A1(n23245), .A2(n23257), .ZN(n23241) );
  NOR2_X2 U19533 ( .A1(n7953), .A2(n52016), .ZN(n14164) );
  NAND2_X1 U19576 ( .A1(n2696), .A2(n7952), .ZN(n52016) );
  NAND2_X1 U19587 ( .A1(n18388), .A2(n21726), .ZN(n18389) );
  NAND3_X1 U19605 ( .A1(n44125), .A2(n4941), .A3(n44128), .ZN(n8499) );
  NAND2_X1 U19627 ( .A1(n4284), .A2(n40185), .ZN(n39501) );
  NAND3_X1 U19629 ( .A1(n44432), .A2(n44433), .A3(n44434), .ZN(n3521) );
  NAND2_X1 U19652 ( .A1(n23127), .A2(n24111), .ZN(n24416) );
  AND3_X2 U19714 ( .A1(n94), .A2(n21588), .A3(n21587), .ZN(n24111) );
  NAND2_X2 U19734 ( .A1(n7555), .A2(n11076), .ZN(n15206) );
  NAND3_X1 U19745 ( .A1(n37524), .A2(n37522), .A3(n37523), .ZN(n6994) );
  OAI21_X1 U19757 ( .B1(n51175), .B2(n14149), .A(n14156), .ZN(n2659) );
  NAND4_X1 U19850 ( .A1(n52017), .A2(n13748), .A3(n14198), .A4(n13746), .ZN(
        n13753) );
  NAND3_X1 U19854 ( .A1(n13745), .A2(n14717), .A3(n13744), .ZN(n52017) );
  NAND3_X1 U19855 ( .A1(n1044), .A2(n37802), .A3(n39481), .ZN(n36218) );
  NAND3_X1 U19861 ( .A1(n18974), .A2(n5271), .A3(n17201), .ZN(n18977) );
  NAND2_X1 U19904 ( .A1(n14574), .A2(n14577), .ZN(n14133) );
  NAND2_X1 U19907 ( .A1(n9698), .A2(n10722), .ZN(n12286) );
  XNOR2_X2 U19932 ( .A(n8998), .B(Key[116]), .ZN(n10722) );
  INV_X1 U19938 ( .A(n45648), .ZN(n45650) );
  NAND2_X1 U19947 ( .A1(n46244), .A2(n49161), .ZN(n45648) );
  NAND2_X1 U19964 ( .A1(n52248), .A2(n8612), .ZN(n9070) );
  AND2_X1 U19965 ( .A1(n23473), .A2(n23160), .ZN(n21166) );
  NOR2_X2 U19970 ( .A1(n50680), .A2(n50721), .ZN(n50710) );
  AOI21_X2 U19986 ( .B1(n18984), .B2(n18983), .A(n18982), .ZN(n22978) );
  NAND2_X1 U19992 ( .A1(n48205), .A2(n52161), .ZN(n44998) );
  NAND3_X1 U19994 ( .A1(n32091), .A2(n32560), .A3(n31609), .ZN(n31616) );
  XNOR2_X1 U20013 ( .A(n52018), .B(n17756), .ZN(n17760) );
  XNOR2_X1 U20024 ( .A(n17755), .B(n17754), .ZN(n52018) );
  OAI211_X1 U20044 ( .C1(n5416), .C2(n52049), .A(n52019), .B(n40752), .ZN(
        n40364) );
  NAND2_X1 U20054 ( .A1(n40357), .A2(n41342), .ZN(n52019) );
  NAND2_X1 U20077 ( .A1(n3631), .A2(n48888), .ZN(n7607) );
  NAND2_X1 U20097 ( .A1(n4111), .A2(n1931), .ZN(n39843) );
  INV_X1 U20109 ( .A(n39918), .ZN(n52020) );
  NAND4_X1 U20132 ( .A1(n9011), .A2(n52021), .A3(n9010), .A4(n9012), .ZN(n9019) );
  OAI211_X1 U20158 ( .C1(n9003), .C2(n9703), .A(n12294), .B(n12291), .ZN(
        n52021) );
  NAND2_X1 U20170 ( .A1(n37648), .A2(n7483), .ZN(n36401) );
  NAND2_X1 U20189 ( .A1(n24092), .A2(n24091), .ZN(n30699) );
  XNOR2_X2 U20196 ( .A(n5954), .B(n23939), .ZN(n24091) );
  INV_X2 U20198 ( .A(n14311), .ZN(n13827) );
  NAND2_X1 U20236 ( .A1(n12568), .A2(n12569), .ZN(n12571) );
  NAND3_X1 U20260 ( .A1(n42103), .A2(n41795), .A3(n8346), .ZN(n201) );
  NAND2_X1 U20288 ( .A1(n41793), .A2(n889), .ZN(n42103) );
  XNOR2_X1 U20289 ( .A(n2327), .B(n7933), .ZN(n52022) );
  NAND3_X1 U20296 ( .A1(n15636), .A2(n19896), .A3(n19887), .ZN(n19635) );
  NAND2_X1 U20299 ( .A1(n29252), .A2(n28650), .ZN(n29125) );
  NAND2_X1 U20343 ( .A1(n29257), .A2(n52023), .ZN(n28651) );
  OR2_X2 U20370 ( .A1(n52024), .A2(n43440), .ZN(n49514) );
  NAND4_X1 U20383 ( .A1(n43437), .A2(n43438), .A3(n43436), .A4(n43435), .ZN(
        n52024) );
  NAND3_X1 U20385 ( .A1(n52025), .A2(n26943), .A3(n26940), .ZN(n51263) );
  NAND2_X1 U20401 ( .A1(n26951), .A2(n26950), .ZN(n52025) );
  NAND4_X2 U20452 ( .A1(n11385), .A2(n11384), .A3(n11386), .A4(n11383), .ZN(
        n14103) );
  NAND2_X1 U20458 ( .A1(n5180), .A2(n12515), .ZN(n11539) );
  NAND2_X1 U20497 ( .A1(n36155), .A2(n38523), .ZN(n36166) );
  XNOR2_X1 U20509 ( .A(n52026), .B(n45439), .ZN(n45497) );
  XNOR2_X1 U20510 ( .A(n45440), .B(n45438), .ZN(n52026) );
  XNOR2_X1 U20526 ( .A(n52027), .B(n35557), .ZN(n35559) );
  XNOR2_X1 U20547 ( .A(n37114), .B(n35556), .ZN(n52027) );
  NAND2_X1 U20554 ( .A1(n28793), .A2(n28971), .ZN(n29714) );
  OR2_X2 U20563 ( .A1(n49606), .A2(n49608), .ZN(n49585) );
  AND2_X2 U20568 ( .A1(n7729), .A2(n38659), .ZN(n38663) );
  NAND2_X1 U20576 ( .A1(n52028), .A2(n32765), .ZN(n32190) );
  NAND2_X1 U20591 ( .A1(n3339), .A2(n32182), .ZN(n52028) );
  NAND3_X1 U20593 ( .A1(n48437), .A2(n48269), .A3(n48433), .ZN(n52178) );
  NAND3_X1 U20635 ( .A1(n45595), .A2(n44664), .A3(n2390), .ZN(n3570) );
  NAND3_X2 U20645 ( .A1(n52240), .A2(n2282), .A3(n14061), .ZN(n3710) );
  XNOR2_X2 U20650 ( .A(n33549), .B(n33550), .ZN(n37001) );
  NAND4_X2 U20684 ( .A1(n29681), .A2(n29680), .A3(n29679), .A4(n29678), .ZN(
        n33549) );
  AND2_X2 U20744 ( .A1(n38575), .A2(n38200), .ZN(n38566) );
  XNOR2_X1 U20775 ( .A(n27467), .B(n25889), .ZN(n22282) );
  NAND3_X1 U20802 ( .A1(n173), .A2(n47932), .A3(n172), .ZN(n4913) );
  NAND2_X1 U20809 ( .A1(n52030), .A2(n49146), .ZN(n7842) );
  XNOR2_X2 U20810 ( .A(n43351), .B(n46095), .ZN(n49146) );
  INV_X1 U20823 ( .A(n49137), .ZN(n52030) );
  NAND2_X1 U20837 ( .A1(n47990), .A2(n47938), .ZN(n47939) );
  NAND2_X2 U20950 ( .A1(n52031), .A2(n46454), .ZN(n48659) );
  AOI22_X1 U20952 ( .A1(n5429), .A2(n48448), .B1(n48469), .B2(n46445), .ZN(
        n52032) );
  NAND4_X1 U20966 ( .A1(n47431), .A2(n52033), .A3(n47429), .A4(n47430), .ZN(
        n47432) );
  NAND3_X1 U20967 ( .A1(n47427), .A2(n49908), .A3(n49877), .ZN(n52033) );
  NAND2_X1 U20992 ( .A1(n8039), .A2(n14175), .ZN(n4584) );
  NAND2_X2 U21004 ( .A1(n6347), .A2(n4652), .ZN(n16450) );
  XNOR2_X1 U21052 ( .A(n52064), .B(n4931), .ZN(Plaintext[60]) );
  XNOR2_X1 U21069 ( .A(n52034), .B(n24489), .ZN(n24490) );
  XNOR2_X1 U21072 ( .A(n52331), .B(n24762), .ZN(n52034) );
  XNOR2_X2 U21090 ( .A(n52035), .B(n46107), .ZN(n49731) );
  XNOR2_X1 U21095 ( .A(n46110), .B(n6210), .ZN(n52035) );
  OAI211_X1 U21102 ( .C1(n52036), .C2(n47953), .A(n47952), .B(n47951), .ZN(
        n47956) );
  NOR2_X1 U21106 ( .A1(n47942), .A2(n47943), .ZN(n52036) );
  NOR2_X1 U21110 ( .A1(n41055), .A2(n41064), .ZN(n40496) );
  NAND2_X1 U21123 ( .A1(n41049), .A2(n41063), .ZN(n41055) );
  NAND2_X2 U21161 ( .A1(n36557), .A2(n36571), .ZN(n36490) );
  AND2_X2 U21162 ( .A1(n45237), .A2(n46359), .ZN(n45231) );
  INV_X2 U21193 ( .A(n48751), .ZN(n48759) );
  AND2_X2 U21195 ( .A1(n48451), .A2(n46444), .ZN(n48448) );
  XOR2_X1 U21221 ( .A(n48694), .B(n4886), .Z(Plaintext[62]) );
  XNOR2_X1 U21264 ( .A(n16563), .B(n16564), .ZN(n52037) );
  CLKBUF_X1 U21269 ( .A(n5724), .Z(n52038) );
  XNOR2_X1 U21374 ( .A(n42170), .B(n45293), .ZN(n5724) );
  NOR2_X1 U21375 ( .A1(n24105), .A2(n24098), .ZN(n24113) );
  OAI21_X1 U21391 ( .B1(n1001), .B2(n8271), .A(n39331), .ZN(n1723) );
  XOR2_X1 U21469 ( .A(n44245), .B(n44244), .Z(n52039) );
  AND2_X1 U21474 ( .A1(n52040), .A2(n23592), .ZN(n23593) );
  NAND4_X1 U21485 ( .A1(n52155), .A2(n17418), .A3(n23591), .A4(n23590), .ZN(
        n52040) );
  AND2_X1 U21541 ( .A1(n46901), .A2(n3999), .ZN(n52041) );
  NAND4_X2 U21544 ( .A1(n1961), .A2(n14144), .A3(n14787), .A4(n1962), .ZN(
        n18126) );
  NAND3_X2 U21547 ( .A1(n34707), .A2(n34708), .A3(n51163), .ZN(n41650) );
  AND2_X2 U21554 ( .A1(n6941), .A2(n51190), .ZN(n41642) );
  XNOR2_X1 U21579 ( .A(n44533), .B(n44532), .ZN(n46721) );
  AND2_X1 U21597 ( .A1(n2742), .A2(n48416), .ZN(n48179) );
  OAI211_X2 U21615 ( .C1(n42447), .C2(n42446), .A(n42445), .B(n42444), .ZN(
        n44216) );
  AND3_X1 U21616 ( .A1(n48156), .A2(n52344), .A3(n48100), .ZN(n48141) );
  XNOR2_X2 U21655 ( .A(n4771), .B(Key[56]), .ZN(n10959) );
  NAND4_X2 U21761 ( .A1(n8761), .A2(n46809), .A3(n46807), .A4(n46808), .ZN(
        n50886) );
  BUF_X1 U21767 ( .A(n45101), .Z(n52043) );
  NAND4_X1 U21776 ( .A1(n46698), .A2(n46697), .A3(n46696), .A4(n46695), .ZN(
        n52044) );
  NAND4_X1 U21795 ( .A1(n46698), .A2(n46697), .A3(n46696), .A4(n46695), .ZN(
        n52045) );
  NAND4_X1 U21838 ( .A1(n46698), .A2(n46697), .A3(n46696), .A4(n46695), .ZN(
        n47563) );
  BUF_X2 U21839 ( .A(n46245), .Z(n539) );
  BUF_X2 U21840 ( .A(n46245), .Z(n540) );
  AND2_X1 U21871 ( .A1(n19673), .A2(n19680), .ZN(n20209) );
  XNOR2_X1 U21900 ( .A(n25248), .B(n28388), .ZN(n3143) );
  AND2_X1 U21901 ( .A1(n32595), .A2(n32590), .ZN(n52046) );
  OR3_X1 U21915 ( .A1(n36112), .A2(n36115), .A3(n35103), .ZN(n38120) );
  INV_X1 U21994 ( .A(n36112), .ZN(n38485) );
  OR4_X2 U22057 ( .A1(n7753), .A2(n18069), .A3(n7752), .A4(n18073), .ZN(n52048) );
  NOR2_X1 U22073 ( .A1(n41356), .A2(n41355), .ZN(n52049) );
  OR4_X1 U22140 ( .A1(n7753), .A2(n18069), .A3(n7752), .A4(n18073), .ZN(n22176) );
  BUF_X2 U22141 ( .A(n16849), .Z(n23483) );
  AND2_X1 U22154 ( .A1(n39060), .A2(n52314), .ZN(n39068) );
  OR2_X1 U22190 ( .A1(n7119), .A2(n52048), .ZN(n52414) );
  OR2_X1 U22223 ( .A1(n21223), .A2(n19518), .ZN(n17415) );
  INV_X1 U22247 ( .A(n16673), .ZN(n21233) );
  AND2_X1 U22248 ( .A1(n47795), .A2(n45872), .ZN(n1902) );
  XNOR2_X1 U22265 ( .A(n41907), .B(n8760), .ZN(n52050) );
  NAND2_X1 U22285 ( .A1(n48778), .A2(n48759), .ZN(n52051) );
  INV_X1 U22286 ( .A(n49719), .ZN(n52052) );
  BUF_X2 U22327 ( .A(n42971), .Z(n49719) );
  NOR2_X1 U22412 ( .A1(n45237), .A2(n46276), .ZN(n46357) );
  INV_X1 U22413 ( .A(n38638), .ZN(n68) );
  CLKBUF_X1 U22431 ( .A(n47122), .Z(n52053) );
  AND2_X1 U22485 ( .A1(n52093), .A2(n52098), .ZN(n50869) );
  XNOR2_X1 U22486 ( .A(n33415), .B(n33414), .ZN(n52054) );
  XNOR2_X1 U22527 ( .A(n33415), .B(n33414), .ZN(n39350) );
  AND2_X1 U22544 ( .A1(n42106), .A2(n41796), .ZN(n41794) );
  NOR2_X1 U22547 ( .A1(n49960), .A2(n49959), .ZN(n50144) );
  NAND4_X1 U22577 ( .A1(n44690), .A2(n44688), .A3(n44689), .A4(n44687), .ZN(
        n52056) );
  NAND4_X1 U22607 ( .A1(n44690), .A2(n44688), .A3(n44689), .A4(n44687), .ZN(
        n52057) );
  NAND4_X1 U22702 ( .A1(n38398), .A2(n38397), .A3(n38396), .A4(n38395), .ZN(
        n52058) );
  NAND4_X1 U22784 ( .A1(n38398), .A2(n38397), .A3(n38396), .A4(n38395), .ZN(
        n42450) );
  CLKBUF_X1 U22785 ( .A(n48531), .Z(n52059) );
  OR2_X1 U22786 ( .A1(n48531), .A2(n2207), .ZN(n52060) );
  BUF_X1 U22842 ( .A(n50621), .Z(n52061) );
  INV_X1 U22882 ( .A(n51386), .ZN(n52062) );
  OR2_X1 U22893 ( .A1(n47957), .A2(n52057), .ZN(n47961) );
  NAND2_X1 U22894 ( .A1(n50837), .A2(n50826), .ZN(n52063) );
  OR2_X1 U22936 ( .A1(n51015), .A2(n34928), .ZN(n36617) );
  AND4_X1 U22942 ( .A1(n48677), .A2(n48678), .A3(n48679), .A4(n48676), .ZN(
        n52064) );
  INV_X1 U23032 ( .A(n19514), .ZN(n52065) );
  OR2_X1 U23033 ( .A1(n27669), .A2(n3765), .ZN(n1049) );
  XNOR2_X1 U23034 ( .A(n44245), .B(n44244), .ZN(n52066) );
  NOR2_X2 U23040 ( .A1(n51229), .A2(n52287), .ZN(n52067) );
  NOR2_X1 U23053 ( .A1(n31826), .A2(n30846), .ZN(n30580) );
  AND2_X1 U23154 ( .A1(n47122), .A2(n45138), .ZN(n46854) );
  CLKBUF_X1 U23155 ( .A(Key[178]), .Z(n4687) );
  XNOR2_X1 U23209 ( .A(n41655), .B(n51498), .ZN(n52068) );
  XNOR2_X1 U23261 ( .A(n41655), .B(n51498), .ZN(n5775) );
  XNOR2_X1 U23262 ( .A(n1599), .B(n44022), .ZN(n49274) );
  XNOR2_X1 U23313 ( .A(n44030), .B(n43619), .ZN(n1946) );
  XNOR2_X1 U23314 ( .A(n41857), .B(n41856), .ZN(n48201) );
  NOR2_X1 U23338 ( .A1(n41110), .A2(n41112), .ZN(n41269) );
  NOR2_X2 U23365 ( .A1(n8616), .A2(n44122), .ZN(n50633) );
  OR2_X1 U23410 ( .A1(n664), .A2(n44784), .ZN(n46243) );
  NAND4_X1 U23412 ( .A1(n46887), .A2(n46886), .A3(n46885), .A4(n46884), .ZN(
        n50826) );
  AND2_X1 U23413 ( .A1(n45925), .A2(n45924), .ZN(n52072) );
  BUF_X1 U23469 ( .A(n45772), .Z(n46676) );
  NAND2_X1 U23507 ( .A1(n35026), .A2(n36364), .ZN(n38014) );
  AND2_X1 U23629 ( .A1(n45372), .A2(n48531), .ZN(n48540) );
  NAND2_X1 U23676 ( .A1(n2557), .A2(n36435), .ZN(n52073) );
  NAND4_X1 U23677 ( .A1(n38106), .A2(n38105), .A3(n40083), .A4(n38104), .ZN(
        n52074) );
  NAND4_X1 U23710 ( .A1(n38106), .A2(n38105), .A3(n40083), .A4(n38104), .ZN(
        n52075) );
  INV_X1 U23711 ( .A(n50809), .ZN(n52076) );
  INV_X1 U23712 ( .A(n50809), .ZN(n50781) );
  INV_X1 U23809 ( .A(n50143), .ZN(n52077) );
  AND2_X1 U23915 ( .A1(n52077), .A2(n51442), .ZN(n52078) );
  XNOR2_X1 U23941 ( .A(n42379), .B(n42378), .ZN(n46197) );
  NAND4_X1 U23966 ( .A1(n43801), .A2(n43800), .A3(n43799), .A4(n47142), .ZN(
        n52081) );
  NAND4_X1 U23968 ( .A1(n43801), .A2(n43800), .A3(n43799), .A4(n47142), .ZN(
        n52082) );
  NAND4_X1 U23976 ( .A1(n43801), .A2(n43800), .A3(n43799), .A4(n47142), .ZN(
        n50620) );
  NAND3_X1 U23984 ( .A1(n1864), .A2(n6552), .A3(n2272), .ZN(n39836) );
  BUF_X2 U24005 ( .A(n43740), .Z(n52085) );
  XNOR2_X1 U24050 ( .A(n45358), .B(n43254), .ZN(n43740) );
  XNOR2_X1 U24051 ( .A(n42338), .B(n42698), .ZN(n49276) );
  NAND4_X1 U24070 ( .A1(n38654), .A2(n38655), .A3(n38657), .A4(n38656), .ZN(
        n52087) );
  NAND4_X1 U24128 ( .A1(n38654), .A2(n38655), .A3(n38657), .A4(n38656), .ZN(
        n52088) );
  AND2_X1 U24173 ( .A1(n40014), .A2(n39103), .ZN(n39094) );
  XNOR2_X1 U24215 ( .A(n44901), .B(n52058), .ZN(n52089) );
  NAND2_X1 U24221 ( .A1(n3246), .A2(n2266), .ZN(n52090) );
  NAND2_X1 U24322 ( .A1(n3246), .A2(n2266), .ZN(n52091) );
  NAND2_X1 U24349 ( .A1(n3246), .A2(n2266), .ZN(n45749) );
  INV_X1 U24393 ( .A(n43089), .ZN(n49946) );
  INV_X1 U24504 ( .A(n8332), .ZN(n52092) );
  INV_X1 U24530 ( .A(n8332), .ZN(n42156) );
  NAND4_X1 U24608 ( .A1(n36464), .A2(n36465), .A3(n36463), .A4(n36466), .ZN(
        n52094) );
  NAND4_X1 U24627 ( .A1(n36464), .A2(n36465), .A3(n36463), .A4(n36466), .ZN(
        n52095) );
  NAND4_X1 U24641 ( .A1(n36464), .A2(n36465), .A3(n36463), .A4(n36466), .ZN(
        n39752) );
  INV_X1 U24741 ( .A(n50850), .ZN(n52097) );
  INV_X1 U24789 ( .A(n1441), .ZN(n52098) );
  INV_X1 U24831 ( .A(n1441), .ZN(n50865) );
  OR2_X1 U24855 ( .A1(n45749), .A2(n52434), .ZN(n45743) );
  OR2_X2 U24858 ( .A1(n41723), .A2(n45188), .ZN(n46747) );
  AND2_X1 U24860 ( .A1(n47990), .A2(n47991), .ZN(n47960) );
  INV_X1 U24862 ( .A(n49276), .ZN(n46201) );
  AND2_X1 U24871 ( .A1(n47376), .A2(n47377), .ZN(n52099) );
  AND3_X1 U24879 ( .A1(n3109), .A2(n6622), .A3(n23162), .ZN(n24403) );
  OR2_X1 U24895 ( .A1(n7118), .A2(n2325), .ZN(n40342) );
  OR2_X1 U24915 ( .A1(n48600), .A2(n48604), .ZN(n48618) );
  XNOR2_X1 U24918 ( .A(n25089), .B(n25600), .ZN(n52102) );
  BUF_X2 U24946 ( .A(n390), .Z(n52103) );
  XNOR2_X1 U25016 ( .A(n25600), .B(n25089), .ZN(n30265) );
  XNOR2_X1 U25025 ( .A(n43106), .B(n45327), .ZN(n390) );
  INV_X1 U25026 ( .A(n36122), .ZN(n52104) );
  XNOR2_X2 U25056 ( .A(n35602), .B(n35601), .ZN(n36122) );
  NAND2_X1 U25072 ( .A1(n45967), .A2(n49199), .ZN(n52105) );
  NAND2_X1 U25073 ( .A1(n45967), .A2(n49199), .ZN(n52106) );
  NAND2_X1 U25112 ( .A1(n45967), .A2(n49199), .ZN(n46222) );
  NOR2_X1 U25325 ( .A1(n2726), .A2(n6116), .ZN(n49669) );
  XOR2_X1 U25326 ( .A(n34626), .B(n35403), .Z(n33666) );
  INV_X1 U25494 ( .A(n41085), .ZN(n52108) );
  INV_X1 U25515 ( .A(n41085), .ZN(n38870) );
  NAND2_X1 U25605 ( .A1(n8676), .A2(n52112), .ZN(n52109) );
  AND2_X1 U25683 ( .A1(n52109), .A2(n52110), .ZN(n29660) );
  OR2_X1 U25748 ( .A1(n52111), .A2(n2366), .ZN(n52110) );
  INV_X1 U25814 ( .A(n725), .ZN(n52111) );
  AND2_X1 U25831 ( .A1(n29992), .A2(n725), .ZN(n52112) );
  NOR2_X1 U25832 ( .A1(n50539), .A2(n52113), .ZN(n1095) );
  AND2_X1 U25944 ( .A1(n50562), .A2(n50564), .ZN(n52113) );
  AND2_X1 U25957 ( .A1(n45909), .A2(n49710), .ZN(n49722) );
  NOR2_X2 U25983 ( .A1(n271), .A2(n52114), .ZN(n48908) );
  NAND2_X1 U26103 ( .A1(n52115), .A2(n2685), .ZN(n52114) );
  OR2_X1 U26332 ( .A1(n45664), .A2(n2688), .ZN(n52115) );
  NAND2_X1 U26424 ( .A1(n44665), .A2(n48273), .ZN(n48434) );
  AND2_X1 U26565 ( .A1(n1155), .A2(n52116), .ZN(n49118) );
  NOR2_X1 U26571 ( .A1(n49112), .A2(n49127), .ZN(n52116) );
  AND2_X1 U26754 ( .A1(n49702), .A2(n49703), .ZN(n52403) );
  NAND3_X1 U26807 ( .A1(n29406), .A2(n29404), .A3(n29405), .ZN(n52117) );
  INV_X1 U26863 ( .A(n50483), .ZN(n7139) );
  INV_X1 U26864 ( .A(n49205), .ZN(n52304) );
  AND2_X1 U26891 ( .A1(n2091), .A2(n32705), .ZN(n32333) );
  NOR2_X2 U26892 ( .A1(n6715), .A2(n28527), .ZN(n2091) );
  INV_X1 U27267 ( .A(n47777), .ZN(n52118) );
  INV_X1 U27324 ( .A(n47777), .ZN(n47790) );
  OR2_X1 U27630 ( .A1(n1383), .A2(n47790), .ZN(n47785) );
  AOI21_X1 U27631 ( .B1(n48437), .B2(n48264), .A(n48432), .ZN(n44658) );
  INV_X1 U27691 ( .A(n52383), .ZN(n52382) );
  XNOR2_X1 U27793 ( .A(n37292), .B(n35088), .ZN(n52119) );
  NOR2_X1 U27911 ( .A1(n42131), .A2(n41770), .ZN(n42153) );
  NAND2_X1 U27929 ( .A1(n8553), .A2(n8554), .ZN(n41395) );
  AND4_X1 U27971 ( .A1(n40323), .A2(n40321), .A3(n40322), .A4(n40324), .ZN(
        n52122) );
  NOR2_X1 U27992 ( .A1(n26966), .A2(n26967), .ZN(n31114) );
  XNOR2_X1 U28007 ( .A(n44979), .B(n1357), .ZN(n45091) );
  NAND2_X1 U28020 ( .A1(n49198), .A2(n45966), .ZN(n45970) );
  INV_X1 U28306 ( .A(n49993), .ZN(n52124) );
  INV_X1 U28368 ( .A(n50708), .ZN(n52126) );
  NAND4_X1 U28391 ( .A1(n40977), .A2(n40978), .A3(n40976), .A4(n40975), .ZN(
        n43318) );
  NOR2_X1 U28437 ( .A1(n41149), .A2(n39836), .ZN(n40380) );
  NOR2_X1 U28438 ( .A1(n677), .A2(n39836), .ZN(n40382) );
  XNOR2_X2 U28439 ( .A(n6763), .B(n33418), .ZN(n37781) );
  BUF_X1 U28462 ( .A(n42044), .Z(n52128) );
  OR2_X1 U28464 ( .A1(n49534), .A2(n52129), .ZN(n49532) );
  NAND2_X1 U28471 ( .A1(n43490), .A2(n49529), .ZN(n52129) );
  OR2_X1 U28479 ( .A1(n47638), .A2(n47639), .ZN(n47641) );
  XOR2_X1 U28493 ( .A(n19254), .B(n19253), .Z(n19256) );
  OR2_X1 U28633 ( .A1(n38659), .A2(n39184), .ZN(n38237) );
  AND3_X1 U28683 ( .A1(n2053), .A2(n22118), .A3(n2054), .ZN(n2052) );
  XNOR2_X1 U28865 ( .A(n44061), .B(n5379), .ZN(n52130) );
  XOR2_X1 U29055 ( .A(n43066), .B(n43067), .Z(n52131) );
  OR2_X1 U29065 ( .A1(n3100), .A2(n23510), .ZN(n4710) );
  OR2_X1 U29066 ( .A1(n32472), .A2(n32484), .ZN(n32028) );
  OR2_X1 U29067 ( .A1(n46587), .A2(n46709), .ZN(n46596) );
  OR2_X1 U29172 ( .A1(n28960), .A2(n52251), .ZN(n52250) );
  OR2_X1 U29177 ( .A1(n30265), .A2(n30256), .ZN(n30272) );
  AND2_X2 U29179 ( .A1(n2031), .A2(n1920), .ZN(n48834) );
  XOR2_X1 U29193 ( .A(Key[190]), .B(Ciphertext[15]), .Z(n52132) );
  NAND4_X1 U29210 ( .A1(n19084), .A2(n19083), .A3(n19082), .A4(n19081), .ZN(
        n52133) );
  NAND4_X1 U29268 ( .A1(n19084), .A2(n19083), .A3(n19082), .A4(n19081), .ZN(
        n52134) );
  NAND4_X1 U29485 ( .A1(n19084), .A2(n19083), .A3(n19082), .A4(n19081), .ZN(
        n23244) );
  NAND4_X4 U29486 ( .A1(n36601), .A2(n36602), .A3(n8366), .A4(n36599), .ZN(
        n40684) );
  OR2_X1 U29489 ( .A1(n32025), .A2(n32491), .ZN(n32015) );
  INV_X1 U29513 ( .A(n15185), .ZN(n17118) );
  XNOR2_X1 U29526 ( .A(n44074), .B(n45484), .ZN(n45067) );
  XOR2_X1 U29545 ( .A(n6846), .B(n43983), .Z(n52136) );
  CLKBUF_X1 U29555 ( .A(n36841), .Z(n52138) );
  OR2_X1 U29760 ( .A1(n42006), .A2(n41581), .ZN(n41509) );
  XNOR2_X1 U29761 ( .A(n18578), .B(n18577), .ZN(n21441) );
  OR2_X1 U29776 ( .A1(n40820), .A2(n40818), .ZN(n39071) );
  NAND3_X1 U29784 ( .A1(n1834), .A2(n15430), .A3(n15429), .ZN(n52141) );
  NAND3_X1 U29786 ( .A1(n1834), .A2(n15430), .A3(n15429), .ZN(n52142) );
  XNOR2_X1 U29812 ( .A(Key[110]), .B(Ciphertext[31]), .ZN(n12595) );
  NAND3_X1 U29826 ( .A1(n1834), .A2(n15430), .A3(n15429), .ZN(n17169) );
  NAND2_X1 U29865 ( .A1(n46614), .A2(n46693), .ZN(n46913) );
  AND2_X1 U29872 ( .A1(n40081), .A2(n40901), .ZN(n5073) );
  NAND2_X2 U29923 ( .A1(n49156), .A2(n49155), .ZN(n49366) );
  XNOR2_X1 U29934 ( .A(n51266), .B(n6653), .ZN(n52143) );
  XNOR2_X1 U29942 ( .A(n51266), .B(n6653), .ZN(n7616) );
  BUF_X1 U29943 ( .A(n25421), .Z(n52144) );
  XNOR2_X1 U29955 ( .A(n8515), .B(n45399), .ZN(n52145) );
  XNOR2_X1 U29961 ( .A(n8515), .B(n45399), .ZN(n5874) );
  XNOR2_X2 U29986 ( .A(n25007), .B(n25006), .ZN(n52147) );
  NAND4_X2 U29992 ( .A1(n52339), .A2(n31460), .A3(n51533), .A4(n31457), .ZN(
        n52148) );
  NAND4_X1 U30017 ( .A1(n52339), .A2(n31460), .A3(n51533), .A4(n31457), .ZN(
        n36669) );
  INV_X1 U30035 ( .A(n45877), .ZN(n47771) );
  AND2_X1 U30072 ( .A1(n45829), .A2(n45819), .ZN(n45836) );
  OR2_X1 U30110 ( .A1(n27119), .A2(n3143), .ZN(n28907) );
  OR2_X1 U30121 ( .A1(n8397), .A2(n12204), .ZN(n52150) );
  NAND4_X1 U30188 ( .A1(n812), .A2(n37676), .A3(n37674), .A4(n37675), .ZN(
        n39695) );
  INV_X1 U30232 ( .A(n10445), .ZN(n52152) );
  AND2_X1 U30242 ( .A1(n11978), .A2(n11979), .ZN(n10445) );
  AND2_X1 U30299 ( .A1(n26960), .A2(n27576), .ZN(n27578) );
  NAND2_X1 U30300 ( .A1(n27576), .A2(n26823), .ZN(n27580) );
  XNOR2_X1 U30302 ( .A(n40286), .B(n40285), .ZN(n52153) );
  XNOR2_X1 U30320 ( .A(n40286), .B(n40285), .ZN(n52154) );
  XNOR2_X1 U30321 ( .A(n40286), .B(n40285), .ZN(n46636) );
  NAND3_X1 U30426 ( .A1(n3408), .A2(n17207), .A3(n17205), .ZN(n24207) );
  INV_X1 U30463 ( .A(n36541), .ZN(n52156) );
  OR2_X1 U30464 ( .A1(n9656), .A2(n10296), .ZN(n52345) );
  XNOR2_X1 U30465 ( .A(n41824), .B(n42487), .ZN(n52161) );
  INV_X1 U30513 ( .A(n50850), .ZN(n50894) );
  BUF_X1 U30528 ( .A(n47592), .Z(n52158) );
  XNOR2_X1 U30612 ( .A(n16563), .B(n16564), .ZN(n20133) );
  INV_X1 U30619 ( .A(n4951), .ZN(n52159) );
  OR2_X1 U30751 ( .A1(n7848), .A2(n40565), .ZN(n52160) );
  BUF_X1 U30808 ( .A(n47935), .Z(n52162) );
  XNOR2_X1 U30843 ( .A(n41824), .B(n42487), .ZN(n45551) );
  NOR2_X1 U30844 ( .A1(n33023), .A2(n33022), .ZN(n52164) );
  NOR2_X1 U30845 ( .A1(n33023), .A2(n33022), .ZN(n6729) );
  AND2_X1 U30851 ( .A1(n31164), .A2(n5479), .ZN(n52351) );
  BUF_X2 U30873 ( .A(n30248), .Z(n52165) );
  OR2_X1 U30896 ( .A1(n46636), .A2(n44873), .ZN(n46630) );
  AND2_X1 U30986 ( .A1(n43184), .A2(n51326), .ZN(n49979) );
  XNOR2_X1 U30988 ( .A(n51398), .B(n7121), .ZN(n52166) );
  XNOR2_X1 U31071 ( .A(n51398), .B(n7121), .ZN(n1925) );
  NOR2_X1 U31140 ( .A1(n42062), .A2(n686), .ZN(n42044) );
  NAND4_X1 U31154 ( .A1(n14867), .A2(n14869), .A3(n14866), .A4(n14868), .ZN(
        n52167) );
  NAND4_X1 U31162 ( .A1(n14867), .A2(n14869), .A3(n14866), .A4(n14868), .ZN(
        n52168) );
  NOR2_X1 U31186 ( .A1(n45848), .A2(n51359), .ZN(n52169) );
  NAND4_X1 U31187 ( .A1(n14867), .A2(n14869), .A3(n14866), .A4(n14868), .ZN(
        n18534) );
  XNOR2_X1 U31193 ( .A(n6265), .B(n28060), .ZN(n52170) );
  BUF_X2 U31268 ( .A(n46043), .Z(n52171) );
  XNOR2_X1 U31273 ( .A(n6265), .B(n28060), .ZN(n7819) );
  NAND4_X1 U31277 ( .A1(n6120), .A2(n39671), .A3(n39669), .A4(n39670), .ZN(
        n46043) );
  NAND4_X1 U31303 ( .A1(n47134), .A2(n6251), .A3(n47132), .A4(n47133), .ZN(
        n50784) );
  AOI21_X2 U31359 ( .B1(n48257), .B2(n48256), .A(n48308), .ZN(n52172) );
  AOI21_X1 U31382 ( .B1(n48257), .B2(n48256), .A(n48308), .ZN(n51318) );
  CLKBUF_X3 U31451 ( .A(n34905), .Z(n39003) );
  OR2_X1 U31452 ( .A1(n29880), .A2(n30376), .ZN(n52173) );
  NAND2_X1 U31519 ( .A1(n7357), .A2(n19880), .ZN(n52174) );
  NAND2_X1 U31546 ( .A1(n7357), .A2(n19880), .ZN(n52175) );
  NAND2_X1 U31595 ( .A1(n7357), .A2(n19880), .ZN(n22769) );
  INV_X1 U31804 ( .A(n4081), .ZN(n52176) );
  BUF_X1 U31805 ( .A(n29327), .Z(n52177) );
  XNOR2_X1 U31881 ( .A(n25933), .B(n27183), .ZN(n29327) );
  AND2_X1 U32077 ( .A1(n46305), .A2(n46304), .ZN(n49047) );
  BUF_X1 U32078 ( .A(n18820), .Z(n52180) );
  XOR2_X1 U32138 ( .A(n27313), .B(n27444), .Z(n52181) );
  AND2_X1 U32225 ( .A1(n35890), .A2(n38340), .ZN(n38323) );
  OR2_X1 U32248 ( .A1(n30163), .A2(n30171), .ZN(n29137) );
  AND2_X1 U32334 ( .A1(n34971), .A2(n36362), .ZN(n38192) );
  BUF_X1 U32337 ( .A(n563), .Z(n52183) );
  XNOR2_X1 U32338 ( .A(n18827), .B(n18832), .ZN(n563) );
  CLKBUF_X1 U32339 ( .A(n25680), .Z(n52184) );
  XNOR2_X1 U32369 ( .A(n9288), .B(Key[169]), .ZN(n9291) );
  NOR2_X1 U32370 ( .A1(n30602), .A2(n30592), .ZN(n31094) );
  INV_X1 U32397 ( .A(n6721), .ZN(n52186) );
  XNOR2_X1 U32490 ( .A(n15831), .B(n15984), .ZN(n21652) );
  XNOR2_X1 U32531 ( .A(n8834), .B(Key[187]), .ZN(n52188) );
  XNOR2_X1 U32543 ( .A(n8834), .B(Key[187]), .ZN(n52189) );
  XNOR2_X1 U32571 ( .A(n17754), .B(n6098), .ZN(n52190) );
  XNOR2_X1 U32572 ( .A(n8834), .B(Key[187]), .ZN(n10915) );
  XNOR2_X1 U32596 ( .A(n17754), .B(n6098), .ZN(n18162) );
  XNOR2_X1 U32633 ( .A(n35079), .B(n35078), .ZN(n52191) );
  NAND2_X1 U32750 ( .A1(n254), .A2(n4875), .ZN(n52192) );
  NAND2_X1 U32790 ( .A1(n254), .A2(n4875), .ZN(n52193) );
  XNOR2_X1 U32791 ( .A(n35079), .B(n35078), .ZN(n35102) );
  NAND2_X1 U32812 ( .A1(n254), .A2(n4875), .ZN(n41293) );
  XNOR2_X1 U32909 ( .A(n8403), .B(n16952), .ZN(n15846) );
  OR2_X1 U32997 ( .A1(n746), .A2(n52147), .ZN(n52195) );
  BUF_X1 U33085 ( .A(n36962), .Z(n52197) );
  NAND4_X1 U33086 ( .A1(n8393), .A2(n7890), .A3(n39199), .A4(n39200), .ZN(
        n41675) );
  XNOR2_X2 U33134 ( .A(n31573), .B(n27553), .ZN(n37040) );
  INV_X1 U33193 ( .A(n2680), .ZN(n52199) );
  XOR2_X1 U33411 ( .A(n19248), .B(n2690), .Z(n52200) );
  XNOR2_X1 U33514 ( .A(n7775), .B(Key[163]), .ZN(n12324) );
  XNOR2_X1 U33597 ( .A(n44205), .B(n44204), .ZN(n52202) );
  XNOR2_X1 U33616 ( .A(n44205), .B(n44204), .ZN(n52203) );
  XNOR2_X1 U33619 ( .A(n24548), .B(n28288), .ZN(n26519) );
  XNOR2_X1 U33670 ( .A(n44205), .B(n44204), .ZN(n45559) );
  XNOR2_X1 U33695 ( .A(n46112), .B(n46113), .ZN(n52204) );
  XNOR2_X1 U33839 ( .A(n18432), .B(n4979), .ZN(n52205) );
  NAND4_X1 U34090 ( .A1(n16991), .A2(n16990), .A3(n16992), .A4(n16989), .ZN(
        n52206) );
  NAND4_X1 U34171 ( .A1(n16991), .A2(n16990), .A3(n16992), .A4(n16989), .ZN(
        n52207) );
  XNOR2_X1 U34430 ( .A(n18432), .B(n4979), .ZN(n6583) );
  NAND4_X1 U34440 ( .A1(n16991), .A2(n16990), .A3(n16992), .A4(n16989), .ZN(
        n21904) );
  NOR2_X1 U34445 ( .A1(n669), .A2(n46872), .ZN(n47087) );
  INV_X1 U34451 ( .A(n4063), .ZN(n52208) );
  XNOR2_X1 U34544 ( .A(n1480), .B(n18651), .ZN(n21605) );
  XNOR2_X1 U34891 ( .A(n33001), .B(n33000), .ZN(n38200) );
  XNOR2_X1 U34928 ( .A(n18438), .B(n17923), .ZN(n18628) );
  INV_X1 U35112 ( .A(n49657), .ZN(n52211) );
  INV_X1 U35113 ( .A(n49657), .ZN(n52212) );
  NAND4_X1 U35124 ( .A1(n38489), .A2(n7749), .A3(n4103), .A4(n38488), .ZN(
        n52214) );
  NAND4_X1 U35134 ( .A1(n38489), .A2(n7749), .A3(n4103), .A4(n38488), .ZN(
        n52215) );
  NAND4_X1 U35147 ( .A1(n38489), .A2(n7749), .A3(n4103), .A4(n38488), .ZN(
        n41323) );
  XNOR2_X1 U35152 ( .A(n7560), .B(n25966), .ZN(n52216) );
  XNOR2_X1 U35161 ( .A(n7560), .B(n25966), .ZN(n52217) );
  BUF_X1 U35208 ( .A(n35398), .Z(n52219) );
  BUF_X1 U35209 ( .A(n35398), .Z(n52220) );
  BUF_X1 U35224 ( .A(n35398), .Z(n52221) );
  XNOR2_X1 U35248 ( .A(n32628), .B(n33806), .ZN(n35398) );
  AND2_X1 U35266 ( .A1(n29123), .A2(n29263), .ZN(n30231) );
  XNOR2_X1 U35271 ( .A(n5891), .B(n42122), .ZN(n52222) );
  XNOR2_X1 U35275 ( .A(n5891), .B(n42122), .ZN(n43524) );
  INV_X1 U35296 ( .A(n47444), .ZN(n52223) );
  NAND4_X1 U35302 ( .A1(n4552), .A2(n4789), .A3(n6990), .A4(n43583), .ZN(
        n52225) );
  NAND4_X1 U35306 ( .A1(n4552), .A2(n4789), .A3(n6990), .A4(n43583), .ZN(
        n52226) );
  XNOR2_X1 U35307 ( .A(n43550), .B(n43549), .ZN(n50317) );
  NAND4_X1 U35342 ( .A1(n4552), .A2(n4789), .A3(n6990), .A4(n43583), .ZN(
        n50640) );
  OAI211_X1 U35444 ( .C1(n211), .C2(n14774), .A(n14772), .B(n1079), .ZN(n52227) );
  OAI211_X1 U35654 ( .C1(n211), .C2(n14774), .A(n14772), .B(n1079), .ZN(n52228) );
  OAI211_X1 U35725 ( .C1(n211), .C2(n14774), .A(n14772), .B(n1079), .ZN(n18548) );
  XNOR2_X1 U35741 ( .A(n16532), .B(n5256), .ZN(n52229) );
  XNOR2_X1 U35819 ( .A(n16532), .B(n5256), .ZN(n18797) );
  NAND3_X1 U35824 ( .A1(n52230), .A2(n642), .A3(n11547), .ZN(n4881) );
  NAND2_X1 U35829 ( .A1(n11544), .A2(n11545), .ZN(n52230) );
  NAND3_X1 U35839 ( .A1(n1287), .A2(n15377), .A3(n15378), .ZN(n15391) );
  XNOR2_X1 U35861 ( .A(n52232), .B(n7364), .ZN(n282) );
  XNOR2_X1 U35863 ( .A(n33435), .B(n165), .ZN(n52232) );
  AOI21_X1 U35878 ( .B1(n52233), .B2(n28557), .A(n30292), .ZN(n28558) );
  NAND2_X1 U35974 ( .A1(n28555), .A2(n30296), .ZN(n52233) );
  INV_X1 U35985 ( .A(n31041), .ZN(n6809) );
  NAND2_X1 U35988 ( .A1(n31826), .A2(n30846), .ZN(n31041) );
  NOR2_X2 U36026 ( .A1(n39077), .A2(n39695), .ZN(n40820) );
  NAND3_X1 U36027 ( .A1(n43477), .A2(n43478), .A3(n43476), .ZN(n43486) );
  INV_X1 U36227 ( .A(n49250), .ZN(n49246) );
  NAND3_X1 U36264 ( .A1(n2003), .A2(n21483), .A3(n20825), .ZN(n19274) );
  NAND3_X1 U36265 ( .A1(n8381), .A2(n36581), .A3(n35204), .ZN(n51202) );
  NAND2_X1 U36272 ( .A1(n3250), .A2(n9073), .ZN(n11604) );
  NOR2_X1 U36329 ( .A1(n31305), .A2(n31302), .ZN(n31297) );
  NAND2_X1 U36331 ( .A1(n30824), .A2(n30644), .ZN(n31305) );
  NAND2_X1 U36334 ( .A1(n52234), .A2(n26890), .ZN(n24573) );
  NAND2_X1 U36335 ( .A1(n26887), .A2(n51770), .ZN(n52234) );
  OAI21_X1 U36358 ( .B1(n13505), .B2(n13527), .A(n8002), .ZN(n12935) );
  NAND2_X1 U36373 ( .A1(n52235), .A2(n4608), .ZN(n1306) );
  OAI21_X1 U36458 ( .B1(n3560), .B2(n9537), .A(n11921), .ZN(n52235) );
  NAND2_X1 U36467 ( .A1(n20044), .A2(n20027), .ZN(n17446) );
  NAND2_X1 U36620 ( .A1(n47898), .A2(n648), .ZN(n47903) );
  NAND3_X1 U36645 ( .A1(n51805), .A2(n47937), .A3(n47989), .ZN(n47980) );
  NAND4_X1 U36650 ( .A1(n39853), .A2(n40329), .A3(n7117), .A4(n40340), .ZN(
        n38845) );
  NAND2_X1 U36772 ( .A1(n17428), .A2(n403), .ZN(n18337) );
  NAND3_X2 U36891 ( .A1(n2276), .A2(n13582), .A3(n5412), .ZN(n14285) );
  NAND2_X1 U36926 ( .A1(n52236), .A2(n39148), .ZN(n39150) );
  NAND2_X1 U36927 ( .A1(n39711), .A2(n39146), .ZN(n52236) );
  NAND2_X1 U36970 ( .A1(n38870), .A2(n41084), .ZN(n39146) );
  NAND3_X1 U37029 ( .A1(n41935), .A2(n41937), .A3(n41936), .ZN(n41945) );
  NAND3_X2 U37032 ( .A1(n35860), .A2(n35859), .A3(n52237), .ZN(n39912) );
  XNOR2_X2 U37033 ( .A(n35224), .B(n36981), .ZN(n33343) );
  NAND4_X2 U37045 ( .A1(n30844), .A2(n30842), .A3(n30845), .A4(n30843), .ZN(
        n36981) );
  XNOR2_X1 U37203 ( .A(n24218), .B(n28383), .ZN(n52238) );
  NAND4_X2 U37214 ( .A1(n52239), .A2(n24368), .A3(n6118), .A4(n4972), .ZN(
        n35254) );
  NAND2_X1 U37215 ( .A1(n2797), .A2(n32254), .ZN(n52239) );
  NAND3_X1 U37227 ( .A1(n14056), .A2(n14055), .A3(n1309), .ZN(n52240) );
  NAND2_X1 U37280 ( .A1(n36589), .A2(n36045), .ZN(n35209) );
  NAND2_X1 U37333 ( .A1(n37356), .A2(n39912), .ZN(n39782) );
  NAND3_X1 U37334 ( .A1(n12247), .A2(n4532), .A3(n4533), .ZN(n12249) );
  NAND2_X1 U37335 ( .A1(n4759), .A2(n4758), .ZN(n27548) );
  NAND2_X2 U37390 ( .A1(n52241), .A2(n32170), .ZN(n36811) );
  BUF_X1 U37395 ( .A(n21925), .Z(n50992) );
  NAND2_X1 U37456 ( .A1(n8186), .A2(n52242), .ZN(n38954) );
  NAND3_X2 U37482 ( .A1(n39436), .A2(n52244), .A3(n52243), .ZN(n42018) );
  NAND2_X1 U37551 ( .A1(n39431), .A2(n39432), .ZN(n52243) );
  NOR2_X1 U37552 ( .A1(n3060), .A2(n52245), .ZN(n16831) );
  AOI21_X1 U37553 ( .B1(n5880), .B2(n16819), .A(n5879), .ZN(n52245) );
  NAND3_X1 U37577 ( .A1(n32730), .A2(n31972), .A3(n52246), .ZN(n31983) );
  OR2_X1 U37580 ( .A1(n31973), .A2(n32719), .ZN(n52246) );
  NAND2_X1 U37626 ( .A1(n22437), .A2(n52247), .ZN(n22438) );
  NAND3_X1 U37627 ( .A1(n36415), .A2(n36414), .A3(n37649), .ZN(n36416) );
  NAND3_X1 U37628 ( .A1(n5939), .A2(n36246), .A3(n5941), .ZN(n41489) );
  NAND2_X1 U37639 ( .A1(n27600), .A2(n30667), .ZN(n24687) );
  NAND3_X1 U37670 ( .A1(n30313), .A2(n30186), .A3(n30164), .ZN(n29138) );
  AOI21_X1 U37674 ( .B1(n8732), .B2(n20975), .A(n52252), .ZN(n20977) );
  NOR2_X1 U37692 ( .A1(n23212), .A2(n52253), .ZN(n52252) );
  INV_X1 U37718 ( .A(n18369), .ZN(n52253) );
  NAND2_X1 U37734 ( .A1(n418), .A2(n23229), .ZN(n23212) );
  NAND4_X2 U37737 ( .A1(n1922), .A2(n1923), .A3(n47166), .A4(n47165), .ZN(
        n50809) );
  NAND2_X1 U37769 ( .A1(n52254), .A2(n50519), .ZN(n100) );
  NAND2_X1 U37770 ( .A1(n50517), .A2(n50518), .ZN(n52254) );
  INV_X1 U37779 ( .A(n21750), .ZN(n51199) );
  NAND3_X1 U37780 ( .A1(n17495), .A2(n17493), .A3(n17494), .ZN(n21750) );
  NAND3_X1 U37794 ( .A1(n52256), .A2(n52255), .A3(n19997), .ZN(n24029) );
  NAND2_X1 U37888 ( .A1(n19991), .A2(n4825), .ZN(n52256) );
  NOR2_X1 U37909 ( .A1(n52258), .A2(n52257), .ZN(n46939) );
  INV_X1 U37944 ( .A(n49031), .ZN(n52257) );
  NAND3_X1 U37947 ( .A1(n35983), .A2(n37381), .A3(n36233), .ZN(n35985) );
  NAND2_X1 U37951 ( .A1(n47045), .A2(n47044), .ZN(n2806) );
  INV_X1 U37972 ( .A(n1733), .ZN(n1730) );
  NAND3_X1 U37976 ( .A1(n122), .A2(n45740), .A3(n6526), .ZN(n1733) );
  OAI21_X1 U37999 ( .B1(n22388), .B2(n22387), .A(n52260), .ZN(n22396) );
  NAND4_X1 U38022 ( .A1(n23813), .A2(n23811), .A3(n22386), .A4(n23814), .ZN(
        n52260) );
  NAND3_X2 U38023 ( .A1(n52262), .A2(n32470), .A3(n52261), .ZN(n34466) );
  NAND2_X1 U38024 ( .A1(n32466), .A2(n32732), .ZN(n52261) );
  NAND2_X1 U38104 ( .A1(n48817), .A2(n48805), .ZN(n3387) );
  NAND3_X1 U38118 ( .A1(n29742), .A2(n29743), .A3(n191), .ZN(n52263) );
  NAND2_X1 U38148 ( .A1(n9747), .A2(n52264), .ZN(n52368) );
  NAND2_X1 U38166 ( .A1(n9749), .A2(n7942), .ZN(n52264) );
  NAND2_X1 U38170 ( .A1(n1195), .A2(n52265), .ZN(n13265) );
  AOI21_X1 U38178 ( .B1(n50705), .B2(n7460), .A(n52266), .ZN(n51279) );
  NAND2_X1 U38194 ( .A1(n50695), .A2(n7456), .ZN(n52266) );
  AND4_X2 U38236 ( .A1(n27100), .A2(n29353), .A3(n7896), .A4(n27099), .ZN(
        n32507) );
  NAND3_X1 U38246 ( .A1(n33020), .A2(n2924), .A3(n33021), .ZN(n33022) );
  NAND3_X1 U38286 ( .A1(n1518), .A2(n18329), .A3(n18340), .ZN(n7753) );
  NOR2_X1 U38297 ( .A1(n19508), .A2(n17309), .ZN(n19110) );
  NAND2_X1 U38349 ( .A1(n21232), .A2(n17412), .ZN(n19508) );
  NAND3_X1 U38358 ( .A1(n4596), .A2(n15927), .A3(n15926), .ZN(n52267) );
  NAND2_X1 U38411 ( .A1(n21879), .A2(n22854), .ZN(n91) );
  NAND2_X1 U38451 ( .A1(n21887), .A2(n22859), .ZN(n22854) );
  NOR2_X1 U38494 ( .A1(n12472), .A2(n12483), .ZN(n11070) );
  NAND3_X1 U38495 ( .A1(n11065), .A2(n11066), .A3(n12480), .ZN(n12472) );
  NAND2_X2 U38549 ( .A1(n8374), .A2(n8376), .ZN(n40014) );
  NAND2_X1 U38576 ( .A1(n52268), .A2(n10104), .ZN(n9481) );
  OR2_X1 U38580 ( .A1(n9480), .A2(n10529), .ZN(n52268) );
  NAND2_X1 U38607 ( .A1(n5915), .A2(n10018), .ZN(n9516) );
  XNOR2_X1 U38698 ( .A(n43139), .B(n44879), .ZN(n44031) );
  NAND4_X2 U38866 ( .A1(n37174), .A2(n37173), .A3(n37176), .A4(n37175), .ZN(
        n43139) );
  NAND2_X1 U38867 ( .A1(n52269), .A2(n24147), .ZN(n1607) );
  NAND3_X1 U38882 ( .A1(n1609), .A2(n24155), .A3(n24146), .ZN(n52269) );
  AND4_X2 U38885 ( .A1(n10115), .A2(n10117), .A3(n10113), .A4(n10114), .ZN(
        n14178) );
  XNOR2_X2 U38968 ( .A(n52270), .B(n8190), .ZN(n20432) );
  XNOR2_X1 U38970 ( .A(n17782), .B(n17783), .ZN(n52270) );
  INV_X1 U38980 ( .A(n17607), .ZN(n17608) );
  NAND2_X1 U39104 ( .A1(n17603), .A2(n20086), .ZN(n17607) );
  NAND2_X1 U39141 ( .A1(n30718), .A2(n29853), .ZN(n30705) );
  XNOR2_X2 U39184 ( .A(n7945), .B(n7944), .ZN(n29853) );
  INV_X1 U39239 ( .A(n20270), .ZN(n52271) );
  NAND2_X1 U39323 ( .A1(n32356), .A2(n1385), .ZN(n32351) );
  NAND4_X2 U39325 ( .A1(n18058), .A2(n5856), .A3(n3351), .A4(n19181), .ZN(
        n22188) );
  NAND3_X1 U39443 ( .A1(n7165), .A2(n29180), .A3(n29179), .ZN(n29211) );
  INV_X1 U39476 ( .A(n52272), .ZN(n6594) );
  AOI21_X1 U39496 ( .B1(n20494), .B2(n20495), .A(n21468), .ZN(n52272) );
  NAND3_X1 U39557 ( .A1(n34927), .A2(n34928), .A3(n34929), .ZN(n3839) );
  NAND2_X1 U39924 ( .A1(n51504), .A2(n49939), .ZN(n50305) );
  NAND2_X1 U39926 ( .A1(n46822), .A2(n44458), .ZN(n4) );
  AND2_X2 U39927 ( .A1(n51456), .A2(n7046), .ZN(n46822) );
  NAND2_X1 U39947 ( .A1(n23194), .A2(n23751), .ZN(n23752) );
  INV_X1 U39966 ( .A(n30860), .ZN(n30550) );
  NAND2_X1 U40035 ( .A1(n31578), .A2(n30549), .ZN(n30860) );
  OR2_X1 U40073 ( .A1(n14224), .A2(n13968), .ZN(n12927) );
  NAND2_X1 U40147 ( .A1(n38311), .A2(n37654), .ZN(n37656) );
  NAND2_X1 U40185 ( .A1(n38314), .A2(n35852), .ZN(n38311) );
  NAND2_X1 U40186 ( .A1(n43323), .A2(n51146), .ZN(n40800) );
  AND4_X2 U40248 ( .A1(n4997), .A2(n37814), .A3(n37813), .A4(n52273), .ZN(
        n42138) );
  NAND3_X1 U40253 ( .A1(n39488), .A2(n8198), .A3(n39486), .ZN(n52273) );
  XNOR2_X1 U40307 ( .A(n52274), .B(n18506), .ZN(n18525) );
  XNOR2_X1 U40335 ( .A(n18507), .B(n18520), .ZN(n52274) );
  NAND2_X1 U40339 ( .A1(n42153), .A2(n40258), .ZN(n37816) );
  INV_X1 U40351 ( .A(n30580), .ZN(n31042) );
  NAND3_X1 U40359 ( .A1(n52275), .A2(n7529), .A3(n10338), .ZN(n9179) );
  NAND3_X2 U40364 ( .A1(n7490), .A2(n7489), .A3(n37661), .ZN(n40823) );
  NAND3_X2 U40365 ( .A1(n52276), .A2(n18957), .A3(n18958), .ZN(n26530) );
  NAND2_X1 U40369 ( .A1(n31843), .A2(n31367), .ZN(n2088) );
  NAND3_X1 U40478 ( .A1(n22970), .A2(n22972), .A3(n52277), .ZN(n25029) );
  NAND2_X1 U40489 ( .A1(n1387), .A2(n4245), .ZN(n52278) );
  AND4_X1 U40490 ( .A1(n38845), .A2(n38846), .A3(n38844), .A4(n39642), .ZN(
        n38858) );
  NAND2_X1 U40520 ( .A1(n47485), .A2(n48981), .ZN(n2899) );
  NAND2_X1 U40522 ( .A1(n15177), .A2(n15162), .ZN(n15165) );
  NAND2_X1 U40587 ( .A1(n6044), .A2(n7259), .ZN(n18935) );
  NAND3_X1 U40616 ( .A1(n34974), .A2(n52280), .A3(n52279), .ZN(n34978) );
  NAND3_X1 U40710 ( .A1(n38184), .A2(n36362), .A3(n34970), .ZN(n52280) );
  NAND3_X1 U40712 ( .A1(n52281), .A2(n15637), .A3(n15638), .ZN(n8555) );
  NAND2_X1 U40717 ( .A1(n52282), .A2(n29248), .ZN(n28656) );
  INV_X1 U40741 ( .A(n28652), .ZN(n52282) );
  NAND2_X1 U40747 ( .A1(n29263), .A2(n29247), .ZN(n28652) );
  NAND3_X1 U40748 ( .A1(n21149), .A2(n22262), .A3(n21150), .ZN(n23013) );
  OAI21_X1 U40765 ( .B1(n21148), .B2(n22257), .A(n21755), .ZN(n21150) );
  NAND2_X1 U40766 ( .A1(n52283), .A2(n31356), .ZN(n31357) );
  NAND3_X1 U40783 ( .A1(n36300), .A2(n38214), .A3(n38550), .ZN(n52283) );
  XNOR2_X1 U40784 ( .A(n36818), .B(n52284), .ZN(n36822) );
  XNOR2_X1 U40794 ( .A(n36817), .B(n36819), .ZN(n52284) );
  NAND3_X1 U40802 ( .A1(n6457), .A2(n38264), .A3(n38629), .ZN(n38254) );
  NAND2_X2 U40875 ( .A1(n52285), .A2(n10400), .ZN(n15046) );
  NOR2_X1 U40882 ( .A1(n10396), .A2(n10397), .ZN(n52285) );
  NAND3_X1 U40968 ( .A1(n40576), .A2(n40155), .A3(n52160), .ZN(n40160) );
  XNOR2_X1 U40973 ( .A(n52286), .B(n17252), .ZN(n17287) );
  XNOR2_X1 U41029 ( .A(n4263), .B(n17253), .ZN(n52286) );
  NAND2_X1 U41070 ( .A1(n706), .A2(n8241), .ZN(n8240) );
  AOI21_X1 U41073 ( .B1(n46316), .B2(n46317), .A(n46315), .ZN(n52287) );
  NAND2_X1 U41081 ( .A1(n36337), .A2(n35017), .ZN(n38067) );
  NAND2_X1 U41173 ( .A1(n23169), .A2(n52288), .ZN(n8217) );
  NAND3_X1 U41213 ( .A1(n23184), .A2(n5269), .A3(n52289), .ZN(n52288) );
  NAND3_X1 U41237 ( .A1(n13664), .A2(n13663), .A3(n13665), .ZN(n13666) );
  NAND2_X1 U41264 ( .A1(n31613), .A2(n32097), .ZN(n31614) );
  NAND2_X1 U41289 ( .A1(n45842), .A2(n52290), .ZN(n45856) );
  OR2_X1 U41290 ( .A1(n45843), .A2(n47629), .ZN(n52290) );
  NAND2_X1 U41298 ( .A1(n11066), .A2(n12474), .ZN(n11062) );
  NAND3_X1 U41301 ( .A1(n50892), .A2(n50826), .A3(n50855), .ZN(n50828) );
  NAND2_X1 U41376 ( .A1(n50865), .A2(n50863), .ZN(n50892) );
  NAND4_X2 U41395 ( .A1(n29813), .A2(n29811), .A3(n29810), .A4(n29812), .ZN(
        n35483) );
  NAND2_X1 U41407 ( .A1(n39101), .A2(n39667), .ZN(n40009) );
  INV_X1 U41434 ( .A(n28704), .ZN(n28698) );
  NAND2_X1 U41449 ( .A1(n29308), .A2(n26077), .ZN(n28704) );
  NOR2_X1 U41461 ( .A1(n12264), .A2(n12263), .ZN(n52292) );
  NAND2_X1 U41467 ( .A1(n12262), .A2(n12261), .ZN(n52293) );
  NAND2_X1 U41480 ( .A1(n23707), .A2(n24332), .ZN(n52294) );
  XNOR2_X1 U41481 ( .A(n52296), .B(n42036), .ZN(n42038) );
  XNOR2_X1 U41521 ( .A(n42033), .B(n42034), .ZN(n52296) );
  NAND2_X1 U41587 ( .A1(n9339), .A2(n9335), .ZN(n9974) );
  NOR2_X1 U41588 ( .A1(n31069), .A2(n52297), .ZN(n31071) );
  INV_X1 U41707 ( .A(n31065), .ZN(n52297) );
  NAND2_X1 U41805 ( .A1(n30934), .A2(n31510), .ZN(n31065) );
  NAND2_X1 U41834 ( .A1(n29550), .A2(n29545), .ZN(n27058) );
  XNOR2_X2 U41867 ( .A(n26193), .B(n26192), .ZN(n29545) );
  NAND3_X1 U41881 ( .A1(n21362), .A2(n21364), .A3(n21351), .ZN(n21591) );
  NAND3_X1 U41898 ( .A1(n5070), .A2(n52299), .A3(n52298), .ZN(n43635) );
  NAND2_X1 U41899 ( .A1(n5075), .A2(n38799), .ZN(n52298) );
  OAI211_X1 U42052 ( .C1(n21597), .C2(n21596), .A(n52300), .B(n21595), .ZN(
        n21612) );
  NAND2_X1 U42067 ( .A1(n21593), .A2(n21592), .ZN(n52300) );
  INV_X1 U42074 ( .A(n32701), .ZN(n52301) );
  NAND2_X1 U42083 ( .A1(n41488), .A2(n42442), .ZN(n41492) );
  NAND2_X1 U42102 ( .A1(n933), .A2(n42110), .ZN(n934) );
  NAND2_X1 U42122 ( .A1(n52302), .A2(n4148), .ZN(n26432) );
  OAI21_X1 U42146 ( .B1(n1193), .B2(n24097), .A(n24110), .ZN(n52302) );
  NAND2_X1 U42147 ( .A1(n16043), .A2(n16036), .ZN(n52303) );
  INV_X1 U42166 ( .A(n24149), .ZN(n24153) );
  NAND2_X1 U42173 ( .A1(n21795), .A2(n24157), .ZN(n24149) );
  NAND2_X1 U42233 ( .A1(n1043), .A2(n29905), .ZN(n26832) );
  NOR2_X1 U42243 ( .A1(n1042), .A2(n2774), .ZN(n1043) );
  NAND2_X1 U42245 ( .A1(n1194), .A2(n2037), .ZN(n32987) );
  NAND3_X1 U42250 ( .A1(n45685), .A2(n45683), .A3(n45684), .ZN(n1652) );
  NAND3_X1 U42306 ( .A1(n26196), .A2(n26756), .A3(n29557), .ZN(n26199) );
  XNOR2_X1 U42362 ( .A(n52305), .B(n43525), .ZN(n7719) );
  XNOR2_X1 U42424 ( .A(n43534), .B(n52424), .ZN(n52305) );
  NOR2_X1 U42535 ( .A1(n47448), .A2(n52306), .ZN(n47457) );
  NAND2_X1 U42546 ( .A1(n47446), .A2(n48721), .ZN(n52306) );
  NAND2_X1 U42550 ( .A1(n29541), .A2(n51771), .ZN(n27057) );
  OR2_X2 U42574 ( .A1(n20583), .A2(n20582), .ZN(n7971) );
  INV_X1 U42578 ( .A(n30849), .ZN(n31828) );
  NAND2_X1 U42579 ( .A1(n31826), .A2(n31043), .ZN(n30849) );
  AOI21_X1 U42581 ( .B1(n22682), .B2(n52307), .A(n8149), .ZN(n22683) );
  NAND3_X1 U42658 ( .A1(n23906), .A2(n23913), .A3(n23902), .ZN(n52307) );
  NAND2_X1 U42668 ( .A1(n16222), .A2(n16221), .ZN(n836) );
  NAND2_X1 U42731 ( .A1(n4184), .A2(n31519), .ZN(n30083) );
  INV_X1 U42736 ( .A(n8936), .ZN(n11452) );
  NAND2_X1 U42776 ( .A1(n51672), .A2(n12545), .ZN(n8936) );
  XNOR2_X1 U42858 ( .A(n15799), .B(n15798), .ZN(n52308) );
  NAND3_X1 U42915 ( .A1(n52309), .A2(n41670), .A3(n41234), .ZN(n40713) );
  XNOR2_X1 U42921 ( .A(n41671), .B(n41245), .ZN(n52309) );
  NAND2_X1 U42936 ( .A1(n32438), .A2(n1385), .ZN(n31955) );
  NAND2_X1 U42937 ( .A1(n3260), .A2(n14100), .ZN(n11813) );
  NAND2_X1 U42944 ( .A1(n20497), .A2(n21474), .ZN(n19351) );
  NAND2_X1 U42945 ( .A1(n634), .A2(n19359), .ZN(n21474) );
  NAND2_X1 U43005 ( .A1(n23529), .A2(n52310), .ZN(n23545) );
  NAND2_X1 U43008 ( .A1(n3262), .A2(n52311), .ZN(n12975) );
  NAND2_X1 U43020 ( .A1(n52313), .A2(n52312), .ZN(n52311) );
  NOR2_X1 U43021 ( .A1(n12972), .A2(n14454), .ZN(n52313) );
  NAND3_X1 U43042 ( .A1(n1804), .A2(n27541), .A3(n1803), .ZN(n27549) );
  NAND3_X1 U43058 ( .A1(n41440), .A2(n41436), .A3(n41447), .ZN(n39161) );
  NAND2_X1 U43059 ( .A1(n39160), .A2(n39767), .ZN(n41440) );
  AND2_X2 U43090 ( .A1(n3691), .A2(n22995), .ZN(n22999) );
  BUF_X2 U43113 ( .A(n16673), .Z(n19518) );
  OR2_X2 U43124 ( .A1(n35457), .A2(n35973), .ZN(n37585) );
  NAND2_X1 U43128 ( .A1(n23710), .A2(n170), .ZN(n7215) );
  NAND2_X1 U43129 ( .A1(n2726), .A2(n46028), .ZN(n49654) );
  XNOR2_X2 U43130 ( .A(n43198), .B(n44931), .ZN(n2726) );
  NAND4_X1 U43131 ( .A1(n39054), .A2(n39056), .A3(n52128), .A4(n39055), .ZN(
        n52314) );
  NAND3_X2 U43269 ( .A1(n27967), .A2(n27964), .A3(n52315), .ZN(n31749) );
  NAND2_X1 U43280 ( .A1(n52363), .A2(n30929), .ZN(n4386) );
  XNOR2_X2 U43281 ( .A(n17285), .B(n17286), .ZN(n19777) );
  XNOR2_X1 U43287 ( .A(n52316), .B(n16454), .ZN(n16456) );
  XNOR2_X1 U43389 ( .A(n16453), .B(n17348), .ZN(n52316) );
  OR2_X2 U43390 ( .A1(n52317), .A2(n1510), .ZN(n47777) );
  NAND2_X1 U43403 ( .A1(n7698), .A2(n7699), .ZN(n52317) );
  NAND2_X1 U43464 ( .A1(n52318), .A2(n3072), .ZN(n3071) );
  NAND3_X1 U43523 ( .A1(n3070), .A2(n39347), .A3(n37774), .ZN(n52318) );
  NAND3_X1 U43525 ( .A1(n10468), .A2(n12616), .A3(n52319), .ZN(n10469) );
  NAND2_X1 U43573 ( .A1(n12618), .A2(n9208), .ZN(n10468) );
  XNOR2_X1 U43608 ( .A(n51422), .B(n52320), .ZN(n37328) );
  XNOR2_X1 U43634 ( .A(n37320), .B(n37321), .ZN(n52320) );
  NAND2_X1 U43695 ( .A1(n27987), .A2(n28587), .ZN(n28896) );
  XNOR2_X1 U43710 ( .A(n37333), .B(n37332), .ZN(n51062) );
  NAND4_X1 U43711 ( .A1(n869), .A2(n37339), .A3(n37337), .A4(n37338), .ZN(
        n37342) );
  AND2_X2 U43728 ( .A1(n7794), .A2(n4545), .ZN(n49579) );
  NAND2_X1 U43832 ( .A1(n8564), .A2(n45724), .ZN(n45735) );
  NAND2_X1 U43836 ( .A1(n21200), .A2(n21198), .ZN(n19814) );
  XNOR2_X2 U43898 ( .A(n17387), .B(n17388), .ZN(n21200) );
  NAND2_X1 U43946 ( .A1(n8791), .A2(n51137), .ZN(n12363) );
  NAND4_X4 U43947 ( .A1(n9505), .A2(n9504), .A3(n9506), .A4(n9503), .ZN(n13086) );
  OR2_X1 U43950 ( .A1(n33159), .A2(n51795), .ZN(n7908) );
  AND4_X1 U43959 ( .A1(n4623), .A2(n19015), .A3(n19014), .A4(n6497), .ZN(
        n52348) );
  OAI21_X1 U44040 ( .B1(n12332), .B2(n12333), .A(n12331), .ZN(n12335) );
  NAND3_X1 U44077 ( .A1(n12338), .A2(n10288), .A3(n12323), .ZN(n12331) );
  NAND2_X1 U44095 ( .A1(n30670), .A2(n30663), .ZN(n26856) );
  NAND2_X1 U44105 ( .A1(n47698), .A2(n47699), .ZN(n47701) );
  NAND3_X1 U44170 ( .A1(n2893), .A2(n17049), .A3(n17047), .ZN(n17461) );
  NAND2_X1 U44242 ( .A1(n47763), .A2(n47777), .ZN(n47744) );
  NAND2_X1 U44243 ( .A1(n21782), .A2(n51080), .ZN(n20941) );
  XNOR2_X1 U44297 ( .A(n51785), .B(n16760), .ZN(n8622) );
  NAND4_X2 U44369 ( .A1(n24787), .A2(n24788), .A3(n24789), .A4(n24786), .ZN(
        n35833) );
  OAI211_X1 U44401 ( .C1(n40273), .C2(n2223), .A(n52321), .B(n40271), .ZN(
        n40279) );
  NAND2_X1 U44405 ( .A1(n40274), .A2(n40900), .ZN(n52321) );
  NOR2_X2 U44567 ( .A1(n27549), .A2(n27548), .ZN(n32791) );
  NAND3_X2 U44568 ( .A1(n13984), .A2(n7878), .A3(n8865), .ZN(n17936) );
  NAND3_X1 U44585 ( .A1(n8864), .A2(n12198), .A3(n52150), .ZN(n13977) );
  NOR2_X1 U44598 ( .A1(n8397), .A2(n12204), .ZN(n13576) );
  INV_X1 U44644 ( .A(n1823), .ZN(n52322) );
  NAND3_X1 U44667 ( .A1(n12837), .A2(n785), .A3(n14667), .ZN(n12838) );
  NAND2_X1 U44774 ( .A1(n7421), .A2(n7431), .ZN(n20608) );
  NAND3_X1 U44814 ( .A1(n52323), .A2(n1496), .A3(n24246), .ZN(n1493) );
  INV_X1 U44880 ( .A(n24248), .ZN(n52323) );
  INV_X1 U44881 ( .A(n52324), .ZN(n4198) );
  OAI21_X1 U44954 ( .B1(n38724), .B2(n38319), .A(n39295), .ZN(n52324) );
  XNOR2_X1 U44962 ( .A(n52325), .B(n43214), .ZN(n1254) );
  XNOR2_X1 U45077 ( .A(n18525), .B(n18675), .ZN(n52326) );
  NAND2_X1 U45135 ( .A1(n29143), .A2(n29138), .ZN(n51178) );
  NAND2_X1 U45208 ( .A1(n52328), .A2(n52327), .ZN(n4546) );
  NAND2_X1 U45215 ( .A1(n12086), .A2(n12092), .ZN(n52328) );
  NAND3_X1 U45235 ( .A1(n31855), .A2(n31856), .A3(n4299), .ZN(n31857) );
  OAI211_X1 U45331 ( .C1(n10095), .C2(n10526), .A(n10098), .B(n51783), .ZN(
        n10103) );
  NOR2_X1 U45332 ( .A1(n1416), .A2(n18344), .ZN(n1415) );
  NAND2_X1 U45369 ( .A1(n16807), .A2(n20147), .ZN(n1416) );
  AOI22_X1 U45371 ( .A1(n14807), .A2(n15385), .B1(n15386), .B2(n14819), .ZN(
        n14817) );
  AND4_X2 U45372 ( .A1(n52329), .A2(n38224), .A3(n2721), .A4(n38225), .ZN(
        n41380) );
  NAND2_X2 U45442 ( .A1(n52330), .A2(n13861), .ZN(n4979) );
  AND3_X1 U45593 ( .A1(n13860), .A2(n13859), .A3(n13858), .ZN(n52330) );
  NAND3_X1 U45628 ( .A1(n38717), .A2(n2436), .A3(n5571), .ZN(n35850) );
  XNOR2_X1 U45637 ( .A(n24486), .B(n24487), .ZN(n52331) );
  XNOR2_X1 U45699 ( .A(n52332), .B(n34458), .ZN(n34460) );
  XNOR2_X1 U45700 ( .A(n74), .B(n34457), .ZN(n52332) );
  INV_X2 U45717 ( .A(n49514), .ZN(n49521) );
  NOR2_X1 U45803 ( .A1(n52333), .A2(n924), .ZN(n922) );
  AOI21_X1 U45812 ( .B1(n7391), .B2(n30223), .A(n28661), .ZN(n7574) );
  NAND2_X1 U45875 ( .A1(n51114), .A2(n30233), .ZN(n28658) );
  NAND4_X1 U45891 ( .A1(n47257), .A2(n47587), .A3(n52158), .A4(n47617), .ZN(
        n47263) );
  INV_X1 U45941 ( .A(n21512), .ZN(n21517) );
  NAND3_X1 U45949 ( .A1(n21527), .A2(n21525), .A3(n7160), .ZN(n21512) );
  XNOR2_X1 U45950 ( .A(n52335), .B(n16233), .ZN(n16014) );
  XNOR2_X1 U45989 ( .A(n16913), .B(n16012), .ZN(n52335) );
  NAND3_X1 U46001 ( .A1(n30452), .A2(n30451), .A3(n2328), .ZN(n30453) );
  NAND2_X1 U46020 ( .A1(n21355), .A2(n8490), .ZN(n19289) );
  XNOR2_X2 U46028 ( .A(n36852), .B(n36853), .ZN(n39429) );
  NAND2_X1 U46058 ( .A1(n52336), .A2(n10433), .ZN(n10435) );
  NAND3_X1 U46112 ( .A1(n51577), .A2(n11958), .A3(n10430), .ZN(n52336) );
  NAND2_X1 U46195 ( .A1(n13031), .A2(n3510), .ZN(n2766) );
  OR2_X2 U46281 ( .A1(n6737), .A2(n6739), .ZN(n15133) );
  NAND3_X1 U46431 ( .A1(n10442), .A2(n10443), .A3(n10441), .ZN(n6737) );
  OR2_X2 U46432 ( .A1(n21612), .A2(n21611), .ZN(n24412) );
  NAND2_X1 U46489 ( .A1(n52338), .A2(n52337), .ZN(n11790) );
  INV_X1 U46490 ( .A(n14291), .ZN(n52338) );
  NAND2_X1 U46491 ( .A1(n31446), .A2(n32665), .ZN(n52339) );
  INV_X1 U46517 ( .A(n45756), .ZN(n45758) );
  NAND2_X1 U46521 ( .A1(n44873), .A2(n46637), .ZN(n45756) );
  NAND3_X1 U46525 ( .A1(n11325), .A2(n12166), .A3(n12161), .ZN(n9238) );
  NAND3_X1 U46544 ( .A1(n32664), .A2(n31169), .A3(n31538), .ZN(n31445) );
  NAND2_X1 U46669 ( .A1(n9878), .A2(n2517), .ZN(n8174) );
  NAND2_X1 U46770 ( .A1(n41110), .A2(n41111), .ZN(n41728) );
  NAND2_X2 U46827 ( .A1(n36786), .A2(n8644), .ZN(n41110) );
  XNOR2_X2 U46848 ( .A(n25495), .B(n28220), .ZN(n25664) );
  NAND2_X2 U46863 ( .A1(n6380), .A2(n23929), .ZN(n28220) );
  NAND2_X1 U46870 ( .A1(n47990), .A2(n52162), .ZN(n44716) );
  OAI21_X1 U46871 ( .B1(n41235), .B2(n41679), .A(n40040), .ZN(n40717) );
  NAND2_X1 U46897 ( .A1(n3861), .A2(n41685), .ZN(n40040) );
  NAND2_X1 U46930 ( .A1(n52340), .A2(n37974), .ZN(n4356) );
  NAND2_X1 U46932 ( .A1(n36349), .A2(n36073), .ZN(n52340) );
  NAND2_X1 U46940 ( .A1(n2086), .A2(n63), .ZN(n36570) );
  NAND3_X1 U46941 ( .A1(n52425), .A2(n18964), .A3(n18965), .ZN(n18972) );
  XNOR2_X1 U46992 ( .A(n52341), .B(n50923), .ZN(Plaintext[187]) );
  NAND4_X1 U46993 ( .A1(n2863), .A2(n2862), .A3(n50922), .A4(n50921), .ZN(
        n52341) );
  NAND2_X1 U47006 ( .A1(n4582), .A2(n38255), .ZN(n52342) );
  NAND2_X1 U47010 ( .A1(n45749), .A2(n48834), .ZN(n48819) );
  AND2_X2 U47122 ( .A1(n31892), .A2(n31899), .ZN(n29995) );
  NOR2_X1 U47187 ( .A1(n92), .A2(n20184), .ZN(n52343) );
  INV_X1 U47198 ( .A(n48112), .ZN(n52344) );
  NAND2_X1 U47256 ( .A1(n25734), .A2(n27847), .ZN(n29289) );
  NAND2_X1 U47281 ( .A1(n52346), .A2(n52345), .ZN(n9774) );
  NAND2_X1 U47291 ( .A1(n10939), .A2(n10296), .ZN(n52346) );
  NAND3_X2 U47458 ( .A1(n51228), .A2(n39114), .A3(n51227), .ZN(n46150) );
  NAND4_X1 U47494 ( .A1(n44721), .A2(n44718), .A3(n44717), .A4(n44720), .ZN(
        n44723) );
  NAND4_X2 U47502 ( .A1(n52347), .A2(n41127), .A3(n41125), .A4(n41126), .ZN(
        n43889) );
  NAND2_X1 U47554 ( .A1(n41117), .A2(n41116), .ZN(n52347) );
  NAND3_X1 U47593 ( .A1(n5927), .A2(n4820), .A3(n5928), .ZN(n5926) );
  NAND2_X2 U47600 ( .A1(n52348), .A2(n6498), .ZN(n22977) );
  NAND2_X1 U47633 ( .A1(n50805), .A2(n50800), .ZN(n50776) );
  NAND3_X1 U47640 ( .A1(n47093), .A2(n47089), .A3(n47111), .ZN(n47090) );
  NAND2_X1 U47644 ( .A1(n2159), .A2(n46869), .ZN(n47088) );
  XNOR2_X2 U47686 ( .A(n19235), .B(n17925), .ZN(n17798) );
  NAND2_X2 U47742 ( .A1(n52387), .A2(n1908), .ZN(n17925) );
  NAND2_X1 U47748 ( .A1(n35920), .A2(n52349), .ZN(n35921) );
  NAND3_X1 U47749 ( .A1(n692), .A2(n37745), .A3(n691), .ZN(n52349) );
  NAND3_X1 U47781 ( .A1(n10585), .A2(n10584), .A3(n580), .ZN(n10010) );
  NAND2_X1 U47790 ( .A1(n41978), .A2(n39620), .ZN(n39622) );
  NAND2_X1 U47791 ( .A1(n32614), .A2(n31566), .ZN(n31160) );
  XNOR2_X2 U47827 ( .A(n52350), .B(n42682), .ZN(n46203) );
  XNOR2_X1 U47836 ( .A(n42320), .B(n42985), .ZN(n52350) );
  NAND4_X2 U47996 ( .A1(n52351), .A2(n4513), .A3(n31163), .A4(n3363), .ZN(
        n5234) );
  AND2_X2 U48013 ( .A1(n5683), .A2(n21105), .ZN(n21715) );
  NAND2_X1 U48015 ( .A1(n28300), .A2(n30351), .ZN(n28852) );
  NAND2_X1 U48070 ( .A1(n30346), .A2(n28298), .ZN(n30351) );
  NAND2_X1 U48073 ( .A1(n40726), .A2(n3770), .ZN(n3769) );
  XNOR2_X2 U48113 ( .A(n25294), .B(n25293), .ZN(n51118) );
  NAND4_X2 U48116 ( .A1(n19334), .A2(n7451), .A3(n7450), .A4(n19333), .ZN(
        n22861) );
  NAND3_X1 U48141 ( .A1(n46644), .A2(n46645), .A3(n46643), .ZN(n46646) );
  NAND3_X1 U48167 ( .A1(n6026), .A2(n52086), .A3(n49277), .ZN(n4840) );
  NAND2_X1 U48173 ( .A1(n31815), .A2(n31821), .ZN(n3660) );
  AND4_X2 U48190 ( .A1(n26687), .A2(n6336), .A3(n26686), .A4(n26685), .ZN(
        n31821) );
  NAND2_X1 U48191 ( .A1(n38938), .A2(n38949), .ZN(n39418) );
  NAND3_X1 U48195 ( .A1(n1545), .A2(n13506), .A3(n13526), .ZN(n13524) );
  NAND2_X1 U48223 ( .A1(n44424), .A2(n44420), .ZN(n6756) );
  NAND2_X1 U48224 ( .A1(n26915), .A2(n26916), .ZN(n26917) );
  AND2_X1 U48264 ( .A1(n38557), .A2(n36299), .ZN(n36144) );
  NAND2_X1 U48265 ( .A1(n5181), .A2(n31030), .ZN(n31031) );
  NOR2_X1 U48274 ( .A1(n23243), .A2(n52353), .ZN(n22127) );
  NAND2_X1 U48320 ( .A1(n22125), .A2(n23238), .ZN(n52353) );
  NAND2_X1 U48374 ( .A1(n41210), .A2(n51430), .ZN(n40663) );
  XNOR2_X1 U48416 ( .A(n4530), .B(n52354), .ZN(n42684) );
  XNOR2_X1 U48430 ( .A(n44055), .B(n44553), .ZN(n52354) );
  XNOR2_X2 U48450 ( .A(n25457), .B(n26300), .ZN(n8657) );
  NAND4_X2 U48467 ( .A1(n21677), .A2(n21678), .A3(n21679), .A4(n21676), .ZN(
        n26300) );
  NAND2_X1 U48490 ( .A1(n52356), .A2(n52355), .ZN(n34959) );
  NAND2_X1 U48526 ( .A1(n38093), .A2(n38094), .ZN(n52355) );
  NAND2_X1 U48527 ( .A1(n36313), .A2(n34958), .ZN(n38093) );
  NAND2_X1 U48531 ( .A1(n2049), .A2(n50984), .ZN(n52356) );
  NAND3_X1 U48633 ( .A1(n37505), .A2(n37506), .A3(n37504), .ZN(n37515) );
  NAND2_X1 U48665 ( .A1(n40500), .A2(n41054), .ZN(n39604) );
  NAND3_X1 U48721 ( .A1(n1568), .A2(n39615), .A3(n40807), .ZN(n39619) );
  NAND2_X1 U48722 ( .A1(n41008), .A2(n43323), .ZN(n1568) );
  AND2_X2 U48784 ( .A1(n27632), .A2(n26804), .ZN(n27730) );
  NAND2_X1 U48785 ( .A1(n49113), .A2(n5662), .ZN(n7518) );
  NAND3_X1 U48789 ( .A1(n13629), .A2(n14674), .A3(n2150), .ZN(n13637) );
  OAI21_X1 U48826 ( .B1(n30829), .B2(n30830), .A(n30828), .ZN(n31296) );
  NAND3_X1 U48827 ( .A1(n13309), .A2(n13310), .A3(n14038), .ZN(n52358) );
  NAND3_X1 U48845 ( .A1(n3384), .A2(n10922), .A3(n10923), .ZN(n10928) );
  NAND3_X1 U48848 ( .A1(n40717), .A2(n41237), .A3(n40716), .ZN(n40720) );
  OAI21_X1 U48849 ( .B1(n49083), .B2(n49066), .A(n49057), .ZN(n4378) );
  NAND3_X1 U48851 ( .A1(n5661), .A2(n5662), .A3(n1502), .ZN(n49057) );
  NAND2_X1 U48916 ( .A1(n1707), .A2(n29234), .ZN(n25111) );
  NAND2_X1 U48969 ( .A1(n26903), .A2(n52359), .ZN(n26908) );
  NAND2_X1 U49004 ( .A1(n29420), .A2(n52360), .ZN(n52359) );
  OAI21_X1 U49007 ( .B1(n28153), .B2(n28547), .A(n52361), .ZN(n27116) );
  OR2_X1 U49009 ( .A1(n27112), .A2(n30295), .ZN(n52361) );
  OAI21_X1 U49026 ( .B1(n19358), .B2(n21468), .A(n52362), .ZN(n19361) );
  INV_X1 U49041 ( .A(n19357), .ZN(n52362) );
  INV_X1 U49088 ( .A(n31519), .ZN(n52363) );
  NAND3_X2 U49090 ( .A1(n30217), .A2(n5241), .A3(n30215), .ZN(n32609) );
  NAND3_X1 U49091 ( .A1(n9118), .A2(n52365), .A3(n12549), .ZN(n9120) );
  NAND2_X1 U49092 ( .A1(n12544), .A2(n9117), .ZN(n52365) );
  NAND3_X1 U49132 ( .A1(n32531), .A2(n32530), .A3(n32536), .ZN(n175) );
  NAND2_X1 U49136 ( .A1(n35434), .A2(n6881), .ZN(n6880) );
  INV_X1 U49140 ( .A(n36906), .ZN(n52366) );
  OAI21_X1 U49141 ( .B1(n2340), .B2(n36257), .A(n36256), .ZN(n52367) );
  NAND3_X1 U49159 ( .A1(n36209), .A2(n38980), .A3(n38983), .ZN(n36210) );
  NAND2_X1 U49161 ( .A1(n795), .A2(n11137), .ZN(n10471) );
  OAI21_X1 U49169 ( .B1(n52368), .B2(n51605), .A(n51762), .ZN(n3419) );
  OAI21_X1 U49320 ( .B1(n28569), .B2(n28200), .A(n52369), .ZN(n28210) );
  NAND2_X1 U49335 ( .A1(n28198), .A2(n52370), .ZN(n52369) );
  XNOR2_X2 U49493 ( .A(n1274), .B(n42927), .ZN(n42990) );
  OAI21_X1 U49575 ( .B1(n51773), .B2(n52371), .A(n51155), .ZN(n4067) );
  NAND2_X1 U49576 ( .A1(n17080), .A2(n19102), .ZN(n52371) );
  NAND3_X1 U49577 ( .A1(n3020), .A2(n8063), .A3(n8068), .ZN(n1134) );
  INV_X1 U49585 ( .A(n4235), .ZN(n52372) );
  NAND2_X1 U49586 ( .A1(n50958), .A2(n50913), .ZN(n50935) );
  NAND3_X1 U49615 ( .A1(n4692), .A2(n50478), .A3(n50465), .ZN(n50447) );
  NAND3_X1 U49622 ( .A1(n52373), .A2(n23566), .A3(n17074), .ZN(n1246) );
  NAND2_X1 U49624 ( .A1(n23565), .A2(n1648), .ZN(n52373) );
  XNOR2_X1 U49799 ( .A(n6773), .B(n23840), .ZN(n23388) );
  XNOR2_X2 U49838 ( .A(n27451), .B(n26210), .ZN(n6773) );
  NAND4_X4 U49846 ( .A1(n23576), .A2(n23575), .A3(n23578), .A4(n23577), .ZN(
        n26589) );
  XNOR2_X1 U49859 ( .A(n52374), .B(n35119), .ZN(n4133) );
  XNOR2_X1 U49860 ( .A(n35122), .B(n36832), .ZN(n52374) );
  NAND2_X1 U49871 ( .A1(n696), .A2(n36051), .ZN(n36592) );
  NAND3_X1 U49877 ( .A1(n50963), .A2(n50961), .A3(n4504), .ZN(n4503) );
  OAI21_X1 U49979 ( .B1(n51806), .B2(n52169), .A(n52375), .ZN(n46925) );
  NAND2_X1 U50003 ( .A1(n52169), .A2(n46913), .ZN(n52375) );
  NAND2_X1 U50062 ( .A1(n49987), .A2(n49980), .ZN(n49624) );
  NAND3_X1 U50163 ( .A1(n40959), .A2(n40960), .A3(n51853), .ZN(n40961) );
  NAND2_X2 U50164 ( .A1(n1219), .A2(n52376), .ZN(n18475) );
  INV_X1 U50179 ( .A(n14639), .ZN(n52376) );
  NOR2_X1 U50288 ( .A1(n11304), .A2(n14635), .ZN(n14639) );
  NAND3_X2 U50307 ( .A1(n4701), .A2(n8485), .A3(n4700), .ZN(n23480) );
  NAND3_X1 U50341 ( .A1(n52377), .A2(n14273), .A3(n15128), .ZN(n14274) );
  NAND3_X1 U50352 ( .A1(n2986), .A2(n2241), .A3(n14267), .ZN(n52377) );
  NAND2_X1 U50388 ( .A1(n16841), .A2(n16840), .ZN(n16842) );
  NAND2_X1 U50389 ( .A1(n20140), .A2(n52378), .ZN(n20152) );
  NAND2_X1 U50408 ( .A1(n20137), .A2(n20138), .ZN(n52378) );
  NAND2_X1 U50410 ( .A1(n18345), .A2(n18344), .ZN(n20137) );
  NAND3_X1 U50459 ( .A1(n46633), .A2(n52154), .A3(n46628), .ZN(n46625) );
  OAI21_X1 U50478 ( .B1(n31139), .B2(n31140), .A(n52379), .ZN(n31152) );
  NAND2_X1 U50483 ( .A1(n31140), .A2(n31423), .ZN(n52379) );
  NAND2_X1 U50485 ( .A1(n52380), .A2(n36275), .ZN(n36279) );
  NAND2_X1 U50586 ( .A1(n36270), .A2(n36271), .ZN(n52380) );
  NAND3_X1 U50587 ( .A1(n32838), .A2(n31073), .A3(n32385), .ZN(n32846) );
  INV_X1 U50626 ( .A(n19562), .ZN(n52381) );
  OAI22_X1 U50748 ( .A1(n42048), .A2(n42062), .B1(n1332), .B2(n42049), .ZN(
        n42051) );
  NAND3_X1 U50790 ( .A1(n41040), .A2(n40417), .A3(n397), .ZN(n40427) );
  NAND2_X1 U50791 ( .A1(n38589), .A2(n38584), .ZN(n36137) );
  NAND2_X1 U50801 ( .A1(n14974), .A2(n52382), .ZN(n13676) );
  OAI21_X1 U50832 ( .B1(n13688), .B2(n14982), .A(n352), .ZN(n52383) );
  NAND2_X1 U50835 ( .A1(n14984), .A2(n14983), .ZN(n15108) );
  NAND4_X2 U50897 ( .A1(n35021), .A2(n35022), .A3(n35019), .A4(n35020), .ZN(
        n41029) );
  INV_X1 U50910 ( .A(n52384), .ZN(n8073) );
  OAI21_X1 U50915 ( .B1(n12679), .B2(n12672), .A(n11493), .ZN(n52384) );
  NAND3_X1 U50919 ( .A1(n52385), .A2(n11021), .A3(n11033), .ZN(n10007) );
  NAND2_X1 U50925 ( .A1(n10585), .A2(n10005), .ZN(n52385) );
  OAI21_X1 U50931 ( .B1(n13818), .B2(n13819), .A(n14306), .ZN(n13821) );
  NAND2_X1 U50934 ( .A1(n13827), .A2(n25), .ZN(n14306) );
  OR2_X2 U50957 ( .A1(n18048), .A2(n18049), .ZN(n22184) );
  OAI21_X1 U50958 ( .B1(n46539), .B2(n48093), .A(n51804), .ZN(n8069) );
  NAND2_X1 U50966 ( .A1(n5917), .A2(n11648), .ZN(n5916) );
  NAND2_X1 U50983 ( .A1(n21715), .A2(n7119), .ZN(n21100) );
  NAND4_X1 U50984 ( .A1(n20636), .A2(n20637), .A3(n20634), .A4(n20635), .ZN(
        n52386) );
  NAND3_X1 U50988 ( .A1(n12421), .A2(n1911), .A3(n12422), .ZN(n52387) );
  NAND2_X1 U50991 ( .A1(n47798), .A2(n47797), .ZN(n4588) );
  NAND2_X1 U50992 ( .A1(n47741), .A2(n47742), .ZN(n47798) );
  NAND3_X1 U50993 ( .A1(n11463), .A2(n11478), .A3(n11462), .ZN(n11465) );
  XNOR2_X1 U50994 ( .A(n2162), .B(n52388), .ZN(n15231) );
  NAND3_X1 U51013 ( .A1(n3035), .A2(n32962), .A3(n32175), .ZN(n2933) );
  NAND2_X1 U51014 ( .A1(n51540), .A2(n18455), .ZN(n18472) );
  NAND2_X1 U51018 ( .A1(n51796), .A2(n52390), .ZN(n52389) );
  NAND3_X1 U51020 ( .A1(n47301), .A2(n47300), .A3(n50308), .ZN(n47305) );
  NAND3_X1 U51044 ( .A1(n52397), .A2(n29826), .A3(n1396), .ZN(n33541) );
  NAND3_X1 U51045 ( .A1(n18355), .A2(n19066), .A3(n51756), .ZN(n18367) );
  NAND2_X1 U51046 ( .A1(n52391), .A2(n38499), .ZN(n2940) );
  NAND2_X1 U51047 ( .A1(n38490), .A2(n38491), .ZN(n52391) );
  NAND2_X1 U51048 ( .A1(n50208), .A2(n50226), .ZN(n50211) );
  NAND2_X1 U51049 ( .A1(n50222), .A2(n602), .ZN(n50208) );
  NAND2_X1 U51050 ( .A1(n47002), .A2(n47001), .ZN(n47004) );
  AND2_X2 U51051 ( .A1(n52392), .A2(n7206), .ZN(n50189) );
  NAND2_X1 U51052 ( .A1(n7205), .A2(n47308), .ZN(n52392) );
  INV_X1 U51053 ( .A(n39444), .ZN(n39447) );
  NAND2_X1 U51054 ( .A1(n36898), .A2(n39438), .ZN(n39444) );
  NAND3_X1 U51055 ( .A1(n44655), .A2(n1664), .A3(n47908), .ZN(n52393) );
  XNOR2_X2 U51056 ( .A(n52394), .B(n26412), .ZN(n29447) );
  XNOR2_X1 U51057 ( .A(n52395), .B(n50220), .ZN(Plaintext[148]) );
  NAND4_X1 U51058 ( .A1(n50218), .A2(n50216), .A3(n50219), .A4(n50217), .ZN(
        n52395) );
  XNOR2_X2 U51059 ( .A(n43655), .B(n43157), .ZN(n43755) );
  NAND4_X2 U51060 ( .A1(n39630), .A2(n39631), .A3(n39629), .A4(n39820), .ZN(
        n43157) );
  NAND4_X1 U51061 ( .A1(n39459), .A2(n39456), .A3(n39457), .A4(n39458), .ZN(
        n39470) );
  NAND3_X1 U51062 ( .A1(n31364), .A2(n31365), .A3(n31363), .ZN(n1083) );
  XNOR2_X1 U51063 ( .A(n52396), .B(n50107), .ZN(Plaintext[141]) );
  NAND4_X1 U51064 ( .A1(n50106), .A2(n50103), .A3(n50104), .A4(n50105), .ZN(
        n52396) );
  NAND3_X1 U51065 ( .A1(n6270), .A2(n32912), .A3(n6269), .ZN(n3623) );
  NAND2_X1 U51066 ( .A1(n4145), .A2(n1395), .ZN(n52397) );
  OR2_X2 U51067 ( .A1(n52398), .A2(n50045), .ZN(n50143) );
  AOI21_X1 U51068 ( .B1(n50038), .B2(n50039), .A(n50389), .ZN(n52398) );
  NAND3_X1 U51069 ( .A1(n14108), .A2(n14109), .A3(n6495), .ZN(n7884) );
  NAND3_X1 U51070 ( .A1(n50142), .A2(n50098), .A3(n50133), .ZN(n8602) );
  NAND2_X1 U51071 ( .A1(n52077), .A2(n50128), .ZN(n50133) );
  NAND4_X2 U51072 ( .A1(n52399), .A2(n8505), .A3(n13619), .A4(n13618), .ZN(
        n14903) );
  NAND4_X1 U51073 ( .A1(n13615), .A2(n13616), .A3(n13613), .A4(n13614), .ZN(
        n52399) );
  NAND3_X1 U51074 ( .A1(n52400), .A2(n13318), .A3(n13319), .ZN(n13330) );
  NAND3_X1 U51075 ( .A1(n13315), .A2(n13314), .A3(n14006), .ZN(n52400) );
  NAND3_X1 U51076 ( .A1(n27888), .A2(n30194), .A3(n27887), .ZN(n29340) );
  NAND2_X1 U51077 ( .A1(n38947), .A2(n37906), .ZN(n1143) );
  NAND2_X1 U51078 ( .A1(n47936), .A2(n47989), .ZN(n47935) );
  NAND2_X1 U51079 ( .A1(n46478), .A2(n46318), .ZN(n46312) );
  NAND2_X1 U51080 ( .A1(n52402), .A2(n52401), .ZN(n6844) );
  NAND2_X1 U51081 ( .A1(n17101), .A2(n19052), .ZN(n52402) );
  NAND2_X1 U51082 ( .A1(n11697), .A2(n11711), .ZN(n11715) );
  NAND3_X1 U51083 ( .A1(n49701), .A2(n49700), .A3(n52403), .ZN(n49766) );
  NAND2_X1 U51084 ( .A1(n14320), .A2(n13822), .ZN(n11794) );
  NAND3_X2 U51085 ( .A1(n22356), .A2(n22357), .A3(n22355), .ZN(n22908) );
  OAI21_X1 U51086 ( .B1(n19847), .B2(n19846), .A(n3227), .ZN(n3228) );
  NAND4_X1 U51087 ( .A1(n10395), .A2(n11399), .A3(n10394), .A4(n52404), .ZN(
        n10396) );
  NAND3_X1 U51088 ( .A1(n10391), .A2(n10392), .A3(n11423), .ZN(n52404) );
  XNOR2_X1 U51089 ( .A(n51497), .B(n52405), .ZN(n37280) );
  OAI22_X1 U51090 ( .A1(n46490), .A2(n46502), .B1(n46488), .B2(n46501), .ZN(
        n42799) );
  NAND2_X1 U51091 ( .A1(n13065), .A2(n15251), .ZN(n13066) );
  NAND2_X1 U51092 ( .A1(n15254), .A2(n51764), .ZN(n13065) );
  XNOR2_X1 U51093 ( .A(n52406), .B(n42746), .ZN(n42748) );
  XNOR2_X1 U51094 ( .A(n42745), .B(n42869), .ZN(n52406) );
  NAND2_X1 U51095 ( .A1(n47087), .A2(n47098), .ZN(n5986) );
  AND2_X1 U51096 ( .A1(n30652), .A2(n31303), .ZN(n52407) );
  NAND2_X1 U51097 ( .A1(n4945), .A2(n9922), .ZN(n9923) );
  NAND2_X1 U51098 ( .A1(n52408), .A2(n2809), .ZN(n17308) );
  OAI21_X1 U51099 ( .B1(n21272), .B2(n19785), .A(n21269), .ZN(n52408) );
  XNOR2_X1 U51100 ( .A(n52409), .B(n46553), .ZN(Plaintext[47]) );
  NAND2_X1 U51101 ( .A1(n4288), .A2(n46551), .ZN(n52409) );
  NAND2_X1 U51102 ( .A1(n47592), .A2(n47591), .ZN(n47210) );
  NAND2_X1 U51103 ( .A1(n38264), .A2(n37688), .ZN(n35308) );
  OAI211_X1 U51104 ( .C1(n7458), .C2(n50699), .A(n50698), .B(n52410), .ZN(
        Plaintext[171]) );
  NAND2_X1 U51105 ( .A1(n51279), .A2(n50697), .ZN(n52410) );
  OAI21_X1 U51106 ( .B1(n31773), .B2(n31772), .A(n31771), .ZN(n52412) );
  NAND2_X1 U51107 ( .A1(n41269), .A2(n52413), .ZN(n4871) );
  INV_X1 U51108 ( .A(n11605), .ZN(n9900) );
  NAND2_X1 U51109 ( .A1(n9280), .A2(n9281), .ZN(n11605) );
  NAND3_X1 U51110 ( .A1(n38028), .A2(n34939), .A3(n35156), .ZN(n34941) );
  NAND2_X1 U51111 ( .A1(n22175), .A2(n52414), .ZN(n22177) );
  NAND2_X1 U51112 ( .A1(n21106), .A2(n21700), .ZN(n22175) );
  AOI22_X1 U51113 ( .A1(n52416), .A2(n14982), .B1(n14983), .B2(n13681), .ZN(
        n13687) );
  INV_X1 U51114 ( .A(n14976), .ZN(n52416) );
  NAND2_X1 U51115 ( .A1(n5414), .A2(n14252), .ZN(n14976) );
  NAND3_X2 U51116 ( .A1(n22054), .A2(n51786), .A3(n22052), .ZN(n23525) );
  OR2_X2 U51117 ( .A1(n29435), .A2(n29436), .ZN(n30924) );
  NAND2_X1 U51118 ( .A1(n17446), .A2(n20043), .ZN(n18383) );
  NAND2_X1 U51119 ( .A1(n40342), .A2(n40340), .ZN(n37865) );
  INV_X1 U51120 ( .A(n15040), .ZN(n15043) );
  NAND3_X1 U51121 ( .A1(n13480), .A2(n15046), .A3(n277), .ZN(n15040) );
  NAND2_X1 U51122 ( .A1(n2650), .A2(n52417), .ZN(n3506) );
  NAND2_X1 U51123 ( .A1(n30712), .A2(n30723), .ZN(n52418) );
  NAND3_X1 U51124 ( .A1(n5128), .A2(n40376), .A3(n40375), .ZN(n5127) );
  NAND2_X1 U51125 ( .A1(n52419), .A2(n13692), .ZN(n18157) );
  NAND3_X2 U51126 ( .A1(n52420), .A2(n3584), .A3(n5657), .ZN(n13089) );
  NAND3_X1 U51127 ( .A1(n7436), .A2(n35313), .A3(n7437), .ZN(n7435) );
  NAND3_X2 U51128 ( .A1(n37875), .A2(n1216), .A3(n52421), .ZN(n43696) );
  NOR2_X1 U51129 ( .A1(n38849), .A2(n37866), .ZN(n52421) );
  NAND2_X1 U51130 ( .A1(n52422), .A2(n12162), .ZN(n12164) );
  OAI21_X1 U51131 ( .B1(n12157), .B2(n12158), .A(n12169), .ZN(n52422) );
  NAND3_X2 U51132 ( .A1(n12185), .A2(n12182), .A3(n52423), .ZN(n14542) );
  NAND3_X1 U51133 ( .A1(n8144), .A2(n1737), .A3(n3387), .ZN(n122) );
  XNOR2_X1 U51134 ( .A(n43533), .B(n46073), .ZN(n52424) );
  NAND2_X1 U51135 ( .A1(n18961), .A2(n51222), .ZN(n52425) );
  NAND3_X1 U51136 ( .A1(n52426), .A2(n1732), .A3(n1725), .ZN(Plaintext[73]) );
  NAND3_X2 U51137 ( .A1(n28826), .A2(n212), .A3(n28825), .ZN(n34381) );
  NAND3_X1 U51138 ( .A1(n30416), .A2(n28971), .A3(n30417), .ZN(n7690) );
  XNOR2_X1 U51139 ( .A(n52427), .B(n49549), .ZN(Plaintext[119]) );
  NAND4_X1 U51140 ( .A1(n49545), .A2(n49547), .A3(n49546), .A4(n49548), .ZN(
        n52427) );
  NAND3_X1 U51141 ( .A1(n3295), .A2(n18498), .A3(n18497), .ZN(n18504) );
  NOR2_X1 U51142 ( .A1(n50542), .A2(n50553), .ZN(n50551) );
  AND3_X2 U51143 ( .A1(n5508), .A2(n5510), .A3(n5513), .ZN(n13633) );
  NAND2_X1 U51144 ( .A1(n52428), .A2(n20686), .ZN(n1536) );
  OAI22_X1 U51145 ( .A1(n20679), .A2(n20685), .B1(n18105), .B2(n18101), .ZN(
        n52428) );
  NAND2_X2 U51146 ( .A1(n1045), .A2(n12946), .ZN(n18539) );
  OAI22_X1 U51147 ( .A1(n12442), .A2(n12443), .B1(n12712), .B2(n12714), .ZN(
        n12445) );
  NAND3_X1 U51148 ( .A1(n52429), .A2(n17630), .A3(n17628), .ZN(n17631) );
  NAND3_X1 U51149 ( .A1(n17625), .A2(n19344), .A3(n17626), .ZN(n52429) );
  NOR2_X1 U51150 ( .A1(n51263), .A2(n52430), .ZN(n51168) );
  NAND3_X1 U51151 ( .A1(n26953), .A2(n26942), .A3(n26941), .ZN(n52430) );
  NAND2_X1 U51152 ( .A1(n52432), .A2(n52431), .ZN(n30076) );
  NAND2_X1 U51153 ( .A1(n30075), .A2(n51742), .ZN(n52431) );
  NAND2_X1 U51154 ( .A1(n30074), .A2(n30073), .ZN(n52432) );
  NAND2_X1 U51155 ( .A1(n632), .A2(n489), .ZN(n20507) );
  NAND2_X1 U51156 ( .A1(n12099), .A2(n3611), .ZN(n9682) );
  NAND2_X1 U51157 ( .A1(n12379), .A2(n12389), .ZN(n12099) );
  XNOR2_X2 U51158 ( .A(n7556), .B(n33848), .ZN(n5686) );
  OR2_X2 U51159 ( .A1(n5816), .A2(n5818), .ZN(n7556) );
  BUF_X2 U51160 ( .A(n21063), .Z(n50977) );
  NAND2_X1 U51161 ( .A1(n24292), .A2(n24287), .ZN(n52433) );
  NAND4_X2 U51162 ( .A1(n34327), .A2(n34329), .A3(n34328), .A4(n34326), .ZN(
        n46128) );
  NOR2_X2 U51163 ( .A1(n45507), .A2(n45506), .ZN(n52434) );
endmodule


module SPEEDY_Top ( clk, Ciphertext, Key, Plaintext );
  input [191:0] Ciphertext;
  input [191:0] Key;
  output [191:0] Plaintext;
  input clk;

  wire   [191:0] reg_in;
  wire   [191:0] reg_key;
  wire   [191:0] reg_out;

  DFF_X1 \reg_in_reg[191]  ( .D(Ciphertext[191]), .CK(clk), .Q(reg_in[191]) );
  DFF_X1 \reg_in_reg[190]  ( .D(Ciphertext[190]), .CK(clk), .Q(reg_in[190]) );
  DFF_X1 \reg_in_reg[189]  ( .D(Ciphertext[189]), .CK(clk), .Q(reg_in[189]) );
  DFF_X1 \reg_in_reg[188]  ( .D(Ciphertext[188]), .CK(clk), .Q(reg_in[188]) );
  DFF_X1 \reg_in_reg[187]  ( .D(Ciphertext[187]), .CK(clk), .Q(reg_in[187]) );
  DFF_X1 \reg_in_reg[186]  ( .D(Ciphertext[186]), .CK(clk), .Q(reg_in[186]) );
  DFF_X1 \reg_in_reg[185]  ( .D(Ciphertext[185]), .CK(clk), .Q(reg_in[185]) );
  DFF_X1 \reg_in_reg[184]  ( .D(Ciphertext[184]), .CK(clk), .Q(reg_in[184]) );
  DFF_X1 \reg_in_reg[183]  ( .D(Ciphertext[183]), .CK(clk), .Q(reg_in[183]) );
  DFF_X1 \reg_in_reg[182]  ( .D(Ciphertext[182]), .CK(clk), .Q(reg_in[182]) );
  DFF_X1 \reg_in_reg[181]  ( .D(Ciphertext[181]), .CK(clk), .Q(reg_in[181]) );
  DFF_X1 \reg_in_reg[180]  ( .D(Ciphertext[180]), .CK(clk), .Q(reg_in[180]) );
  DFF_X1 \reg_in_reg[179]  ( .D(Ciphertext[179]), .CK(clk), .Q(reg_in[179]) );
  DFF_X1 \reg_in_reg[178]  ( .D(Ciphertext[178]), .CK(clk), .Q(reg_in[178]) );
  DFF_X1 \reg_in_reg[177]  ( .D(Ciphertext[177]), .CK(clk), .Q(reg_in[177]) );
  DFF_X1 \reg_in_reg[176]  ( .D(Ciphertext[176]), .CK(clk), .Q(reg_in[176]) );
  DFF_X1 \reg_in_reg[175]  ( .D(Ciphertext[175]), .CK(clk), .Q(reg_in[175]) );
  DFF_X1 \reg_in_reg[174]  ( .D(Ciphertext[174]), .CK(clk), .Q(reg_in[174]) );
  DFF_X1 \reg_in_reg[173]  ( .D(Ciphertext[173]), .CK(clk), .Q(reg_in[173]) );
  DFF_X1 \reg_in_reg[172]  ( .D(Ciphertext[172]), .CK(clk), .Q(reg_in[172]) );
  DFF_X1 \reg_in_reg[171]  ( .D(Ciphertext[171]), .CK(clk), .Q(reg_in[171]) );
  DFF_X1 \reg_in_reg[170]  ( .D(Ciphertext[170]), .CK(clk), .Q(reg_in[170]) );
  DFF_X1 \reg_in_reg[169]  ( .D(Ciphertext[169]), .CK(clk), .Q(reg_in[169]) );
  DFF_X1 \reg_in_reg[168]  ( .D(Ciphertext[168]), .CK(clk), .Q(reg_in[168]) );
  DFF_X1 \reg_in_reg[167]  ( .D(Ciphertext[167]), .CK(clk), .Q(reg_in[167]) );
  DFF_X1 \reg_in_reg[166]  ( .D(Ciphertext[166]), .CK(clk), .Q(reg_in[166]) );
  DFF_X1 \reg_in_reg[165]  ( .D(Ciphertext[165]), .CK(clk), .Q(reg_in[165]) );
  DFF_X1 \reg_in_reg[164]  ( .D(Ciphertext[164]), .CK(clk), .Q(reg_in[164]) );
  DFF_X1 \reg_in_reg[163]  ( .D(Ciphertext[163]), .CK(clk), .Q(reg_in[163]) );
  DFF_X1 \reg_in_reg[162]  ( .D(Ciphertext[162]), .CK(clk), .Q(reg_in[162]) );
  DFF_X1 \reg_in_reg[161]  ( .D(Ciphertext[161]), .CK(clk), .Q(reg_in[161]) );
  DFF_X1 \reg_in_reg[160]  ( .D(Ciphertext[160]), .CK(clk), .Q(reg_in[160]) );
  DFF_X1 \reg_in_reg[159]  ( .D(Ciphertext[159]), .CK(clk), .Q(reg_in[159]) );
  DFF_X1 \reg_in_reg[158]  ( .D(Ciphertext[158]), .CK(clk), .Q(reg_in[158]) );
  DFF_X1 \reg_in_reg[157]  ( .D(Ciphertext[157]), .CK(clk), .Q(reg_in[157]) );
  DFF_X1 \reg_in_reg[156]  ( .D(Ciphertext[156]), .CK(clk), .Q(reg_in[156]) );
  DFF_X1 \reg_in_reg[155]  ( .D(Ciphertext[155]), .CK(clk), .Q(reg_in[155]) );
  DFF_X1 \reg_in_reg[154]  ( .D(Ciphertext[154]), .CK(clk), .Q(reg_in[154]) );
  DFF_X1 \reg_in_reg[153]  ( .D(Ciphertext[153]), .CK(clk), .Q(reg_in[153]) );
  DFF_X1 \reg_in_reg[152]  ( .D(Ciphertext[152]), .CK(clk), .Q(reg_in[152]) );
  DFF_X1 \reg_in_reg[151]  ( .D(Ciphertext[151]), .CK(clk), .Q(reg_in[151]) );
  DFF_X1 \reg_in_reg[150]  ( .D(Ciphertext[150]), .CK(clk), .Q(reg_in[150]) );
  DFF_X1 \reg_in_reg[149]  ( .D(Ciphertext[149]), .CK(clk), .Q(reg_in[149]) );
  DFF_X1 \reg_in_reg[148]  ( .D(Ciphertext[148]), .CK(clk), .Q(reg_in[148]) );
  DFF_X1 \reg_in_reg[147]  ( .D(Ciphertext[147]), .CK(clk), .Q(reg_in[147]) );
  DFF_X1 \reg_in_reg[146]  ( .D(Ciphertext[146]), .CK(clk), .Q(reg_in[146]) );
  DFF_X1 \reg_in_reg[145]  ( .D(Ciphertext[145]), .CK(clk), .Q(reg_in[145]) );
  DFF_X1 \reg_in_reg[144]  ( .D(Ciphertext[144]), .CK(clk), .Q(reg_in[144]) );
  DFF_X1 \reg_in_reg[143]  ( .D(Ciphertext[143]), .CK(clk), .Q(reg_in[143]) );
  DFF_X1 \reg_in_reg[142]  ( .D(Ciphertext[142]), .CK(clk), .Q(reg_in[142]) );
  DFF_X1 \reg_in_reg[141]  ( .D(Ciphertext[141]), .CK(clk), .Q(reg_in[141]) );
  DFF_X1 \reg_in_reg[140]  ( .D(Ciphertext[140]), .CK(clk), .Q(reg_in[140]) );
  DFF_X1 \reg_in_reg[139]  ( .D(Ciphertext[139]), .CK(clk), .Q(reg_in[139]) );
  DFF_X1 \reg_in_reg[138]  ( .D(Ciphertext[138]), .CK(clk), .Q(reg_in[138]) );
  DFF_X1 \reg_in_reg[137]  ( .D(Ciphertext[137]), .CK(clk), .Q(reg_in[137]) );
  DFF_X1 \reg_in_reg[136]  ( .D(Ciphertext[136]), .CK(clk), .Q(reg_in[136]) );
  DFF_X1 \reg_in_reg[135]  ( .D(Ciphertext[135]), .CK(clk), .Q(reg_in[135]) );
  DFF_X1 \reg_in_reg[134]  ( .D(Ciphertext[134]), .CK(clk), .Q(reg_in[134]) );
  DFF_X1 \reg_in_reg[133]  ( .D(Ciphertext[133]), .CK(clk), .Q(reg_in[133]) );
  DFF_X1 \reg_in_reg[132]  ( .D(Ciphertext[132]), .CK(clk), .Q(reg_in[132]) );
  DFF_X1 \reg_in_reg[131]  ( .D(Ciphertext[131]), .CK(clk), .Q(reg_in[131]) );
  DFF_X1 \reg_in_reg[130]  ( .D(Ciphertext[130]), .CK(clk), .Q(reg_in[130]) );
  DFF_X1 \reg_in_reg[129]  ( .D(Ciphertext[129]), .CK(clk), .Q(reg_in[129]) );
  DFF_X1 \reg_in_reg[128]  ( .D(Ciphertext[128]), .CK(clk), .Q(reg_in[128]) );
  DFF_X1 \reg_in_reg[127]  ( .D(Ciphertext[127]), .CK(clk), .Q(reg_in[127]) );
  DFF_X1 \reg_in_reg[126]  ( .D(Ciphertext[126]), .CK(clk), .Q(reg_in[126]) );
  DFF_X1 \reg_in_reg[125]  ( .D(Ciphertext[125]), .CK(clk), .Q(reg_in[125]) );
  DFF_X1 \reg_in_reg[124]  ( .D(Ciphertext[124]), .CK(clk), .Q(reg_in[124]) );
  DFF_X1 \reg_in_reg[123]  ( .D(Ciphertext[123]), .CK(clk), .Q(reg_in[123]) );
  DFF_X1 \reg_in_reg[122]  ( .D(Ciphertext[122]), .CK(clk), .Q(reg_in[122]) );
  DFF_X1 \reg_in_reg[121]  ( .D(Ciphertext[121]), .CK(clk), .Q(reg_in[121]) );
  DFF_X1 \reg_in_reg[120]  ( .D(Ciphertext[120]), .CK(clk), .Q(reg_in[120]) );
  DFF_X1 \reg_in_reg[119]  ( .D(Ciphertext[119]), .CK(clk), .Q(reg_in[119]) );
  DFF_X1 \reg_in_reg[118]  ( .D(Ciphertext[118]), .CK(clk), .Q(reg_in[118]) );
  DFF_X1 \reg_in_reg[117]  ( .D(Ciphertext[117]), .CK(clk), .Q(reg_in[117]) );
  DFF_X1 \reg_in_reg[116]  ( .D(Ciphertext[116]), .CK(clk), .Q(reg_in[116]) );
  DFF_X1 \reg_in_reg[115]  ( .D(Ciphertext[115]), .CK(clk), .Q(reg_in[115]) );
  DFF_X1 \reg_in_reg[114]  ( .D(Ciphertext[114]), .CK(clk), .Q(reg_in[114]) );
  DFF_X1 \reg_in_reg[113]  ( .D(Ciphertext[113]), .CK(clk), .Q(reg_in[113]) );
  DFF_X1 \reg_in_reg[112]  ( .D(Ciphertext[112]), .CK(clk), .Q(reg_in[112]) );
  DFF_X1 \reg_in_reg[111]  ( .D(Ciphertext[111]), .CK(clk), .Q(reg_in[111]) );
  DFF_X1 \reg_in_reg[110]  ( .D(Ciphertext[110]), .CK(clk), .Q(reg_in[110]) );
  DFF_X1 \reg_in_reg[109]  ( .D(Ciphertext[109]), .CK(clk), .Q(reg_in[109]) );
  DFF_X1 \reg_in_reg[108]  ( .D(Ciphertext[108]), .CK(clk), .Q(reg_in[108]) );
  DFF_X1 \reg_in_reg[107]  ( .D(Ciphertext[107]), .CK(clk), .Q(reg_in[107]) );
  DFF_X1 \reg_in_reg[106]  ( .D(Ciphertext[106]), .CK(clk), .Q(reg_in[106]) );
  DFF_X1 \reg_in_reg[105]  ( .D(Ciphertext[105]), .CK(clk), .Q(reg_in[105]) );
  DFF_X1 \reg_in_reg[104]  ( .D(Ciphertext[104]), .CK(clk), .Q(reg_in[104]) );
  DFF_X1 \reg_in_reg[103]  ( .D(Ciphertext[103]), .CK(clk), .Q(reg_in[103]) );
  DFF_X1 \reg_in_reg[102]  ( .D(Ciphertext[102]), .CK(clk), .Q(reg_in[102]) );
  DFF_X1 \reg_in_reg[101]  ( .D(Ciphertext[101]), .CK(clk), .Q(reg_in[101]) );
  DFF_X1 \reg_in_reg[100]  ( .D(Ciphertext[100]), .CK(clk), .Q(reg_in[100]) );
  DFF_X1 \reg_in_reg[99]  ( .D(Ciphertext[99]), .CK(clk), .Q(reg_in[99]) );
  DFF_X1 \reg_in_reg[98]  ( .D(Ciphertext[98]), .CK(clk), .Q(reg_in[98]) );
  DFF_X1 \reg_in_reg[97]  ( .D(Ciphertext[97]), .CK(clk), .Q(reg_in[97]) );
  DFF_X1 \reg_in_reg[96]  ( .D(Ciphertext[96]), .CK(clk), .Q(reg_in[96]) );
  DFF_X1 \reg_in_reg[95]  ( .D(Ciphertext[95]), .CK(clk), .Q(reg_in[95]) );
  DFF_X1 \reg_in_reg[94]  ( .D(Ciphertext[94]), .CK(clk), .Q(reg_in[94]) );
  DFF_X1 \reg_in_reg[93]  ( .D(Ciphertext[93]), .CK(clk), .Q(reg_in[93]) );
  DFF_X1 \reg_in_reg[92]  ( .D(Ciphertext[92]), .CK(clk), .Q(reg_in[92]) );
  DFF_X1 \reg_in_reg[91]  ( .D(Ciphertext[91]), .CK(clk), .Q(reg_in[91]) );
  DFF_X1 \reg_in_reg[90]  ( .D(Ciphertext[90]), .CK(clk), .Q(reg_in[90]) );
  DFF_X1 \reg_in_reg[89]  ( .D(Ciphertext[89]), .CK(clk), .Q(reg_in[89]) );
  DFF_X1 \reg_in_reg[88]  ( .D(Ciphertext[88]), .CK(clk), .Q(reg_in[88]) );
  DFF_X1 \reg_in_reg[87]  ( .D(Ciphertext[87]), .CK(clk), .Q(reg_in[87]) );
  DFF_X1 \reg_in_reg[86]  ( .D(Ciphertext[86]), .CK(clk), .Q(reg_in[86]) );
  DFF_X1 \reg_in_reg[85]  ( .D(Ciphertext[85]), .CK(clk), .Q(reg_in[85]) );
  DFF_X1 \reg_in_reg[84]  ( .D(Ciphertext[84]), .CK(clk), .Q(reg_in[84]) );
  DFF_X1 \reg_in_reg[83]  ( .D(Ciphertext[83]), .CK(clk), .Q(reg_in[83]) );
  DFF_X1 \reg_in_reg[82]  ( .D(Ciphertext[82]), .CK(clk), .Q(reg_in[82]) );
  DFF_X1 \reg_in_reg[81]  ( .D(Ciphertext[81]), .CK(clk), .Q(reg_in[81]) );
  DFF_X1 \reg_in_reg[80]  ( .D(Ciphertext[80]), .CK(clk), .Q(reg_in[80]) );
  DFF_X1 \reg_in_reg[79]  ( .D(Ciphertext[79]), .CK(clk), .Q(reg_in[79]) );
  DFF_X1 \reg_in_reg[78]  ( .D(Ciphertext[78]), .CK(clk), .Q(reg_in[78]) );
  DFF_X1 \reg_in_reg[77]  ( .D(Ciphertext[77]), .CK(clk), .Q(reg_in[77]) );
  DFF_X1 \reg_in_reg[76]  ( .D(Ciphertext[76]), .CK(clk), .Q(reg_in[76]) );
  DFF_X1 \reg_in_reg[75]  ( .D(Ciphertext[75]), .CK(clk), .Q(reg_in[75]) );
  DFF_X1 \reg_in_reg[74]  ( .D(Ciphertext[74]), .CK(clk), .Q(reg_in[74]) );
  DFF_X1 \reg_in_reg[73]  ( .D(Ciphertext[73]), .CK(clk), .Q(reg_in[73]) );
  DFF_X1 \reg_in_reg[72]  ( .D(Ciphertext[72]), .CK(clk), .Q(reg_in[72]) );
  DFF_X1 \reg_in_reg[71]  ( .D(Ciphertext[71]), .CK(clk), .Q(reg_in[71]) );
  DFF_X1 \reg_in_reg[70]  ( .D(Ciphertext[70]), .CK(clk), .Q(reg_in[70]) );
  DFF_X1 \reg_in_reg[69]  ( .D(Ciphertext[69]), .CK(clk), .Q(reg_in[69]) );
  DFF_X1 \reg_in_reg[68]  ( .D(Ciphertext[68]), .CK(clk), .Q(reg_in[68]) );
  DFF_X1 \reg_in_reg[67]  ( .D(Ciphertext[67]), .CK(clk), .Q(reg_in[67]) );
  DFF_X1 \reg_in_reg[66]  ( .D(Ciphertext[66]), .CK(clk), .Q(reg_in[66]) );
  DFF_X1 \reg_in_reg[65]  ( .D(Ciphertext[65]), .CK(clk), .Q(reg_in[65]) );
  DFF_X1 \reg_in_reg[64]  ( .D(Ciphertext[64]), .CK(clk), .Q(reg_in[64]) );
  DFF_X1 \reg_in_reg[63]  ( .D(Ciphertext[63]), .CK(clk), .Q(reg_in[63]) );
  DFF_X1 \reg_in_reg[62]  ( .D(Ciphertext[62]), .CK(clk), .Q(reg_in[62]) );
  DFF_X1 \reg_in_reg[61]  ( .D(Ciphertext[61]), .CK(clk), .Q(reg_in[61]) );
  DFF_X1 \reg_in_reg[60]  ( .D(Ciphertext[60]), .CK(clk), .Q(reg_in[60]) );
  DFF_X1 \reg_in_reg[59]  ( .D(Ciphertext[59]), .CK(clk), .Q(reg_in[59]) );
  DFF_X1 \reg_in_reg[58]  ( .D(Ciphertext[58]), .CK(clk), .Q(reg_in[58]) );
  DFF_X1 \reg_in_reg[57]  ( .D(Ciphertext[57]), .CK(clk), .Q(reg_in[57]) );
  DFF_X1 \reg_in_reg[56]  ( .D(Ciphertext[56]), .CK(clk), .Q(reg_in[56]) );
  DFF_X1 \reg_in_reg[55]  ( .D(Ciphertext[55]), .CK(clk), .Q(reg_in[55]) );
  DFF_X1 \reg_in_reg[54]  ( .D(Ciphertext[54]), .CK(clk), .Q(reg_in[54]) );
  DFF_X1 \reg_in_reg[53]  ( .D(Ciphertext[53]), .CK(clk), .Q(reg_in[53]) );
  DFF_X1 \reg_in_reg[52]  ( .D(Ciphertext[52]), .CK(clk), .Q(reg_in[52]) );
  DFF_X1 \reg_in_reg[51]  ( .D(Ciphertext[51]), .CK(clk), .Q(reg_in[51]) );
  DFF_X1 \reg_in_reg[50]  ( .D(Ciphertext[50]), .CK(clk), .Q(reg_in[50]) );
  DFF_X1 \reg_in_reg[49]  ( .D(Ciphertext[49]), .CK(clk), .Q(reg_in[49]) );
  DFF_X1 \reg_in_reg[48]  ( .D(Ciphertext[48]), .CK(clk), .Q(reg_in[48]) );
  DFF_X1 \reg_in_reg[47]  ( .D(Ciphertext[47]), .CK(clk), .Q(reg_in[47]) );
  DFF_X1 \reg_in_reg[46]  ( .D(Ciphertext[46]), .CK(clk), .Q(reg_in[46]) );
  DFF_X1 \reg_in_reg[45]  ( .D(Ciphertext[45]), .CK(clk), .Q(reg_in[45]) );
  DFF_X1 \reg_in_reg[44]  ( .D(Ciphertext[44]), .CK(clk), .Q(reg_in[44]) );
  DFF_X1 \reg_in_reg[43]  ( .D(Ciphertext[43]), .CK(clk), .Q(reg_in[43]) );
  DFF_X1 \reg_in_reg[42]  ( .D(Ciphertext[42]), .CK(clk), .Q(reg_in[42]) );
  DFF_X1 \reg_in_reg[41]  ( .D(Ciphertext[41]), .CK(clk), .Q(reg_in[41]) );
  DFF_X1 \reg_in_reg[40]  ( .D(Ciphertext[40]), .CK(clk), .Q(reg_in[40]) );
  DFF_X1 \reg_in_reg[39]  ( .D(Ciphertext[39]), .CK(clk), .Q(reg_in[39]) );
  DFF_X1 \reg_in_reg[38]  ( .D(Ciphertext[38]), .CK(clk), .Q(reg_in[38]) );
  DFF_X1 \reg_in_reg[37]  ( .D(Ciphertext[37]), .CK(clk), .Q(reg_in[37]) );
  DFF_X1 \reg_in_reg[36]  ( .D(Ciphertext[36]), .CK(clk), .Q(reg_in[36]) );
  DFF_X1 \reg_in_reg[35]  ( .D(Ciphertext[35]), .CK(clk), .Q(reg_in[35]) );
  DFF_X1 \reg_in_reg[34]  ( .D(Ciphertext[34]), .CK(clk), .Q(reg_in[34]) );
  DFF_X1 \reg_in_reg[33]  ( .D(Ciphertext[33]), .CK(clk), .Q(reg_in[33]) );
  DFF_X1 \reg_in_reg[32]  ( .D(Ciphertext[32]), .CK(clk), .Q(reg_in[32]) );
  DFF_X1 \reg_in_reg[31]  ( .D(Ciphertext[31]), .CK(clk), .Q(reg_in[31]) );
  DFF_X1 \reg_in_reg[30]  ( .D(Ciphertext[30]), .CK(clk), .Q(reg_in[30]) );
  DFF_X1 \reg_in_reg[29]  ( .D(Ciphertext[29]), .CK(clk), .Q(reg_in[29]) );
  DFF_X1 \reg_in_reg[28]  ( .D(Ciphertext[28]), .CK(clk), .Q(reg_in[28]) );
  DFF_X1 \reg_in_reg[27]  ( .D(Ciphertext[27]), .CK(clk), .Q(reg_in[27]) );
  DFF_X1 \reg_in_reg[26]  ( .D(Ciphertext[26]), .CK(clk), .Q(reg_in[26]) );
  DFF_X1 \reg_in_reg[25]  ( .D(Ciphertext[25]), .CK(clk), .Q(reg_in[25]) );
  DFF_X1 \reg_in_reg[24]  ( .D(Ciphertext[24]), .CK(clk), .Q(reg_in[24]) );
  DFF_X1 \reg_in_reg[23]  ( .D(Ciphertext[23]), .CK(clk), .Q(reg_in[23]) );
  DFF_X1 \reg_in_reg[22]  ( .D(Ciphertext[22]), .CK(clk), .Q(reg_in[22]) );
  DFF_X1 \reg_in_reg[21]  ( .D(Ciphertext[21]), .CK(clk), .Q(reg_in[21]) );
  DFF_X1 \reg_in_reg[20]  ( .D(Ciphertext[20]), .CK(clk), .Q(reg_in[20]) );
  DFF_X1 \reg_in_reg[19]  ( .D(Ciphertext[19]), .CK(clk), .Q(reg_in[19]) );
  DFF_X1 \reg_in_reg[18]  ( .D(Ciphertext[18]), .CK(clk), .Q(reg_in[18]) );
  DFF_X1 \reg_in_reg[17]  ( .D(Ciphertext[17]), .CK(clk), .Q(reg_in[17]) );
  DFF_X1 \reg_in_reg[16]  ( .D(Ciphertext[16]), .CK(clk), .Q(reg_in[16]) );
  DFF_X1 \reg_in_reg[15]  ( .D(Ciphertext[15]), .CK(clk), .Q(reg_in[15]) );
  DFF_X1 \reg_in_reg[14]  ( .D(Ciphertext[14]), .CK(clk), .Q(reg_in[14]) );
  DFF_X1 \reg_in_reg[13]  ( .D(Ciphertext[13]), .CK(clk), .Q(reg_in[13]) );
  DFF_X1 \reg_in_reg[12]  ( .D(Ciphertext[12]), .CK(clk), .Q(reg_in[12]) );
  DFF_X1 \reg_in_reg[11]  ( .D(Ciphertext[11]), .CK(clk), .Q(reg_in[11]) );
  DFF_X1 \reg_in_reg[10]  ( .D(Ciphertext[10]), .CK(clk), .Q(reg_in[10]) );
  DFF_X1 \reg_in_reg[9]  ( .D(Ciphertext[9]), .CK(clk), .Q(reg_in[9]) );
  DFF_X1 \reg_in_reg[8]  ( .D(Ciphertext[8]), .CK(clk), .Q(reg_in[8]) );
  DFF_X1 \reg_in_reg[7]  ( .D(Ciphertext[7]), .CK(clk), .Q(reg_in[7]) );
  DFF_X1 \reg_in_reg[6]  ( .D(Ciphertext[6]), .CK(clk), .Q(reg_in[6]) );
  DFF_X1 \reg_in_reg[5]  ( .D(Ciphertext[5]), .CK(clk), .Q(reg_in[5]) );
  DFF_X1 \reg_in_reg[4]  ( .D(Ciphertext[4]), .CK(clk), .Q(reg_in[4]) );
  DFF_X1 \reg_in_reg[3]  ( .D(Ciphertext[3]), .CK(clk), .Q(reg_in[3]) );
  DFF_X1 \reg_in_reg[2]  ( .D(Ciphertext[2]), .CK(clk), .Q(reg_in[2]) );
  DFF_X1 \reg_in_reg[1]  ( .D(Ciphertext[1]), .CK(clk), .Q(reg_in[1]) );
  DFF_X1 \reg_in_reg[0]  ( .D(Ciphertext[0]), .CK(clk), .Q(reg_in[0]) );
  DFF_X1 \reg_key_reg[160]  ( .D(Key[160]), .CK(clk), .Q(reg_key[160]) );
  DFF_X1 \reg_key_reg[100]  ( .D(Key[100]), .CK(clk), .Q(reg_key[100]) );
  DFF_X1 \reg_key_reg[77]  ( .D(Key[77]), .CK(clk), .Q(reg_key[77]) );
  DFF_X1 \reg_key_reg[67]  ( .D(Key[67]), .CK(clk), .Q(reg_key[67]) );
  DFF_X1 \reg_key_reg[50]  ( .D(Key[50]), .CK(clk), .Q(reg_key[50]) );
  DFF_X1 \reg_key_reg[47]  ( .D(Key[47]), .CK(clk), .Q(reg_key[47]) );
  DFF_X1 \reg_key_reg[17]  ( .D(Key[17]), .CK(clk), .Q(reg_key[17]) );
  DFF_X1 \Plaintext_reg[191]  ( .D(reg_out[191]), .CK(clk), .Q(Plaintext[191])
         );
  DFF_X1 \Plaintext_reg[190]  ( .D(reg_out[190]), .CK(clk), .Q(Plaintext[190])
         );
  DFF_X1 \Plaintext_reg[189]  ( .D(reg_out[189]), .CK(clk), .Q(Plaintext[189])
         );
  DFF_X1 \Plaintext_reg[187]  ( .D(reg_out[187]), .CK(clk), .Q(Plaintext[187])
         );
  DFF_X1 \Plaintext_reg[186]  ( .D(reg_out[186]), .CK(clk), .Q(Plaintext[186])
         );
  DFF_X1 \Plaintext_reg[185]  ( .D(reg_out[185]), .CK(clk), .Q(Plaintext[185])
         );
  DFF_X1 \Plaintext_reg[184]  ( .D(reg_out[184]), .CK(clk), .Q(Plaintext[184])
         );
  DFF_X1 \Plaintext_reg[183]  ( .D(reg_out[183]), .CK(clk), .Q(Plaintext[183])
         );
  DFF_X1 \Plaintext_reg[182]  ( .D(reg_out[182]), .CK(clk), .Q(Plaintext[182])
         );
  DFF_X1 \Plaintext_reg[180]  ( .D(reg_out[180]), .CK(clk), .Q(Plaintext[180])
         );
  DFF_X1 \Plaintext_reg[179]  ( .D(reg_out[179]), .CK(clk), .Q(Plaintext[179])
         );
  DFF_X1 \Plaintext_reg[178]  ( .D(reg_out[178]), .CK(clk), .Q(Plaintext[178])
         );
  DFF_X1 \Plaintext_reg[177]  ( .D(reg_out[177]), .CK(clk), .Q(Plaintext[177])
         );
  DFF_X1 \Plaintext_reg[176]  ( .D(reg_out[176]), .CK(clk), .Q(Plaintext[176])
         );
  DFF_X1 \Plaintext_reg[175]  ( .D(reg_out[175]), .CK(clk), .Q(Plaintext[175])
         );
  DFF_X1 \Plaintext_reg[174]  ( .D(reg_out[174]), .CK(clk), .Q(Plaintext[174])
         );
  DFF_X1 \Plaintext_reg[173]  ( .D(reg_out[173]), .CK(clk), .Q(Plaintext[173])
         );
  DFF_X1 \Plaintext_reg[172]  ( .D(reg_out[172]), .CK(clk), .Q(Plaintext[172])
         );
  DFF_X1 \Plaintext_reg[171]  ( .D(reg_out[171]), .CK(clk), .Q(Plaintext[171])
         );
  DFF_X1 \Plaintext_reg[170]  ( .D(reg_out[170]), .CK(clk), .Q(Plaintext[170])
         );
  DFF_X1 \Plaintext_reg[169]  ( .D(reg_out[169]), .CK(clk), .Q(Plaintext[169])
         );
  DFF_X1 \Plaintext_reg[168]  ( .D(reg_out[168]), .CK(clk), .Q(Plaintext[168])
         );
  DFF_X1 \Plaintext_reg[166]  ( .D(reg_out[166]), .CK(clk), .Q(Plaintext[166])
         );
  DFF_X1 \Plaintext_reg[165]  ( .D(reg_out[165]), .CK(clk), .Q(Plaintext[165])
         );
  DFF_X1 \Plaintext_reg[164]  ( .D(reg_out[164]), .CK(clk), .Q(Plaintext[164])
         );
  DFF_X1 \Plaintext_reg[163]  ( .D(reg_out[163]), .CK(clk), .Q(Plaintext[163])
         );
  DFF_X1 \Plaintext_reg[162]  ( .D(reg_out[162]), .CK(clk), .Q(Plaintext[162])
         );
  DFF_X1 \Plaintext_reg[160]  ( .D(reg_out[160]), .CK(clk), .Q(Plaintext[160])
         );
  DFF_X1 \Plaintext_reg[159]  ( .D(reg_out[159]), .CK(clk), .Q(Plaintext[159])
         );
  DFF_X1 \Plaintext_reg[158]  ( .D(reg_out[158]), .CK(clk), .Q(Plaintext[158])
         );
  DFF_X1 \Plaintext_reg[157]  ( .D(reg_out[157]), .CK(clk), .Q(Plaintext[157])
         );
  DFF_X1 \Plaintext_reg[156]  ( .D(reg_out[156]), .CK(clk), .Q(Plaintext[156])
         );
  DFF_X1 \Plaintext_reg[154]  ( .D(reg_out[154]), .CK(clk), .Q(Plaintext[154])
         );
  DFF_X1 \Plaintext_reg[153]  ( .D(reg_out[153]), .CK(clk), .Q(Plaintext[153])
         );
  DFF_X1 \Plaintext_reg[152]  ( .D(reg_out[152]), .CK(clk), .Q(Plaintext[152])
         );
  DFF_X1 \Plaintext_reg[151]  ( .D(reg_out[151]), .CK(clk), .Q(Plaintext[151])
         );
  DFF_X1 \Plaintext_reg[150]  ( .D(reg_out[150]), .CK(clk), .Q(Plaintext[150])
         );
  DFF_X1 \Plaintext_reg[149]  ( .D(reg_out[149]), .CK(clk), .Q(Plaintext[149])
         );
  DFF_X1 \Plaintext_reg[148]  ( .D(reg_out[148]), .CK(clk), .Q(Plaintext[148])
         );
  DFF_X1 \Plaintext_reg[147]  ( .D(reg_out[147]), .CK(clk), .Q(Plaintext[147])
         );
  DFF_X1 \Plaintext_reg[146]  ( .D(reg_out[146]), .CK(clk), .Q(Plaintext[146])
         );
  DFF_X1 \Plaintext_reg[145]  ( .D(reg_out[145]), .CK(clk), .Q(Plaintext[145])
         );
  DFF_X1 \Plaintext_reg[144]  ( .D(reg_out[144]), .CK(clk), .Q(Plaintext[144])
         );
  DFF_X1 \Plaintext_reg[143]  ( .D(reg_out[143]), .CK(clk), .Q(Plaintext[143])
         );
  DFF_X1 \Plaintext_reg[142]  ( .D(reg_out[142]), .CK(clk), .Q(Plaintext[142])
         );
  DFF_X1 \Plaintext_reg[141]  ( .D(reg_out[141]), .CK(clk), .Q(Plaintext[141])
         );
  DFF_X1 \Plaintext_reg[140]  ( .D(reg_out[140]), .CK(clk), .Q(Plaintext[140])
         );
  DFF_X1 \Plaintext_reg[139]  ( .D(reg_out[139]), .CK(clk), .Q(Plaintext[139])
         );
  DFF_X1 \Plaintext_reg[138]  ( .D(reg_out[138]), .CK(clk), .Q(Plaintext[138])
         );
  DFF_X1 \Plaintext_reg[137]  ( .D(reg_out[137]), .CK(clk), .Q(Plaintext[137])
         );
  DFF_X1 \Plaintext_reg[136]  ( .D(reg_out[136]), .CK(clk), .Q(Plaintext[136])
         );
  DFF_X1 \Plaintext_reg[135]  ( .D(reg_out[135]), .CK(clk), .Q(Plaintext[135])
         );
  DFF_X1 \Plaintext_reg[134]  ( .D(reg_out[134]), .CK(clk), .Q(Plaintext[134])
         );
  DFF_X1 \Plaintext_reg[133]  ( .D(reg_out[133]), .CK(clk), .Q(Plaintext[133])
         );
  DFF_X1 \Plaintext_reg[132]  ( .D(reg_out[132]), .CK(clk), .Q(Plaintext[132])
         );
  DFF_X1 \Plaintext_reg[131]  ( .D(reg_out[131]), .CK(clk), .Q(Plaintext[131])
         );
  DFF_X1 \Plaintext_reg[130]  ( .D(reg_out[130]), .CK(clk), .Q(Plaintext[130])
         );
  DFF_X1 \Plaintext_reg[128]  ( .D(reg_out[128]), .CK(clk), .Q(Plaintext[128])
         );
  DFF_X1 \Plaintext_reg[127]  ( .D(reg_out[127]), .CK(clk), .Q(Plaintext[127])
         );
  DFF_X1 \Plaintext_reg[126]  ( .D(reg_out[126]), .CK(clk), .Q(Plaintext[126])
         );
  DFF_X1 \Plaintext_reg[125]  ( .D(reg_out[125]), .CK(clk), .Q(Plaintext[125])
         );
  DFF_X1 \Plaintext_reg[124]  ( .D(reg_out[124]), .CK(clk), .Q(Plaintext[124])
         );
  DFF_X1 \Plaintext_reg[123]  ( .D(reg_out[123]), .CK(clk), .Q(Plaintext[123])
         );
  DFF_X1 \Plaintext_reg[122]  ( .D(reg_out[122]), .CK(clk), .Q(Plaintext[122])
         );
  DFF_X1 \Plaintext_reg[121]  ( .D(reg_out[121]), .CK(clk), .Q(Plaintext[121])
         );
  DFF_X1 \Plaintext_reg[120]  ( .D(reg_out[120]), .CK(clk), .Q(Plaintext[120])
         );
  DFF_X1 \Plaintext_reg[119]  ( .D(reg_out[119]), .CK(clk), .Q(Plaintext[119])
         );
  DFF_X1 \Plaintext_reg[118]  ( .D(reg_out[118]), .CK(clk), .Q(Plaintext[118])
         );
  DFF_X1 \Plaintext_reg[117]  ( .D(reg_out[117]), .CK(clk), .Q(Plaintext[117])
         );
  DFF_X1 \Plaintext_reg[116]  ( .D(reg_out[116]), .CK(clk), .Q(Plaintext[116])
         );
  DFF_X1 \Plaintext_reg[115]  ( .D(reg_out[115]), .CK(clk), .Q(Plaintext[115])
         );
  DFF_X1 \Plaintext_reg[113]  ( .D(reg_out[113]), .CK(clk), .Q(Plaintext[113])
         );
  DFF_X1 \Plaintext_reg[112]  ( .D(reg_out[112]), .CK(clk), .Q(Plaintext[112])
         );
  DFF_X1 \Plaintext_reg[111]  ( .D(reg_out[111]), .CK(clk), .Q(Plaintext[111])
         );
  DFF_X1 \Plaintext_reg[110]  ( .D(reg_out[110]), .CK(clk), .Q(Plaintext[110])
         );
  DFF_X1 \Plaintext_reg[109]  ( .D(reg_out[109]), .CK(clk), .Q(Plaintext[109])
         );
  DFF_X1 \Plaintext_reg[108]  ( .D(reg_out[108]), .CK(clk), .Q(Plaintext[108])
         );
  DFF_X1 \Plaintext_reg[107]  ( .D(reg_out[107]), .CK(clk), .Q(Plaintext[107])
         );
  DFF_X1 \Plaintext_reg[106]  ( .D(reg_out[106]), .CK(clk), .Q(Plaintext[106])
         );
  DFF_X1 \Plaintext_reg[105]  ( .D(reg_out[105]), .CK(clk), .Q(Plaintext[105])
         );
  DFF_X1 \Plaintext_reg[104]  ( .D(reg_out[104]), .CK(clk), .Q(Plaintext[104])
         );
  DFF_X1 \Plaintext_reg[103]  ( .D(reg_out[103]), .CK(clk), .Q(Plaintext[103])
         );
  DFF_X1 \Plaintext_reg[102]  ( .D(reg_out[102]), .CK(clk), .Q(Plaintext[102])
         );
  DFF_X1 \Plaintext_reg[101]  ( .D(reg_out[101]), .CK(clk), .Q(Plaintext[101])
         );
  DFF_X1 \Plaintext_reg[100]  ( .D(reg_out[100]), .CK(clk), .Q(Plaintext[100])
         );
  DFF_X1 \Plaintext_reg[99]  ( .D(reg_out[99]), .CK(clk), .Q(Plaintext[99]) );
  DFF_X1 \Plaintext_reg[98]  ( .D(reg_out[98]), .CK(clk), .Q(Plaintext[98]) );
  DFF_X1 \Plaintext_reg[97]  ( .D(reg_out[97]), .CK(clk), .Q(Plaintext[97]) );
  DFF_X1 \Plaintext_reg[96]  ( .D(reg_out[96]), .CK(clk), .Q(Plaintext[96]) );
  DFF_X1 \Plaintext_reg[94]  ( .D(reg_out[94]), .CK(clk), .Q(Plaintext[94]) );
  DFF_X1 \Plaintext_reg[93]  ( .D(reg_out[93]), .CK(clk), .Q(Plaintext[93]) );
  DFF_X1 \Plaintext_reg[91]  ( .D(reg_out[91]), .CK(clk), .Q(Plaintext[91]) );
  DFF_X1 \Plaintext_reg[90]  ( .D(reg_out[90]), .CK(clk), .Q(Plaintext[90]) );
  DFF_X1 \Plaintext_reg[89]  ( .D(reg_out[89]), .CK(clk), .Q(Plaintext[89]) );
  DFF_X1 \Plaintext_reg[88]  ( .D(reg_out[88]), .CK(clk), .Q(Plaintext[88]) );
  DFF_X1 \Plaintext_reg[87]  ( .D(reg_out[87]), .CK(clk), .Q(Plaintext[87]) );
  DFF_X1 \Plaintext_reg[86]  ( .D(reg_out[86]), .CK(clk), .Q(Plaintext[86]) );
  DFF_X1 \Plaintext_reg[85]  ( .D(reg_out[85]), .CK(clk), .Q(Plaintext[85]) );
  DFF_X1 \Plaintext_reg[83]  ( .D(reg_out[83]), .CK(clk), .Q(Plaintext[83]) );
  DFF_X1 \Plaintext_reg[82]  ( .D(reg_out[82]), .CK(clk), .Q(Plaintext[82]) );
  DFF_X1 \Plaintext_reg[81]  ( .D(reg_out[81]), .CK(clk), .Q(Plaintext[81]) );
  DFF_X1 \Plaintext_reg[80]  ( .D(reg_out[80]), .CK(clk), .Q(Plaintext[80]) );
  DFF_X1 \Plaintext_reg[79]  ( .D(reg_out[79]), .CK(clk), .Q(Plaintext[79]) );
  DFF_X1 \Plaintext_reg[78]  ( .D(reg_out[78]), .CK(clk), .Q(Plaintext[78]) );
  DFF_X1 \Plaintext_reg[77]  ( .D(reg_out[77]), .CK(clk), .Q(Plaintext[77]) );
  DFF_X1 \Plaintext_reg[76]  ( .D(reg_out[76]), .CK(clk), .Q(Plaintext[76]) );
  DFF_X1 \Plaintext_reg[75]  ( .D(reg_out[75]), .CK(clk), .Q(Plaintext[75]) );
  DFF_X1 \Plaintext_reg[74]  ( .D(reg_out[74]), .CK(clk), .Q(Plaintext[74]) );
  DFF_X1 \Plaintext_reg[73]  ( .D(reg_out[73]), .CK(clk), .Q(Plaintext[73]) );
  DFF_X1 \Plaintext_reg[72]  ( .D(reg_out[72]), .CK(clk), .Q(Plaintext[72]) );
  DFF_X1 \Plaintext_reg[71]  ( .D(reg_out[71]), .CK(clk), .Q(Plaintext[71]) );
  DFF_X1 \Plaintext_reg[70]  ( .D(reg_out[70]), .CK(clk), .Q(Plaintext[70]) );
  DFF_X1 \Plaintext_reg[69]  ( .D(reg_out[69]), .CK(clk), .Q(Plaintext[69]) );
  DFF_X1 \Plaintext_reg[68]  ( .D(reg_out[68]), .CK(clk), .Q(Plaintext[68]) );
  DFF_X1 \Plaintext_reg[67]  ( .D(reg_out[67]), .CK(clk), .Q(Plaintext[67]) );
  DFF_X1 \Plaintext_reg[66]  ( .D(reg_out[66]), .CK(clk), .Q(Plaintext[66]) );
  DFF_X1 \Plaintext_reg[65]  ( .D(reg_out[65]), .CK(clk), .Q(Plaintext[65]) );
  DFF_X1 \Plaintext_reg[64]  ( .D(reg_out[64]), .CK(clk), .Q(Plaintext[64]) );
  DFF_X1 \Plaintext_reg[63]  ( .D(reg_out[63]), .CK(clk), .Q(Plaintext[63]) );
  DFF_X1 \Plaintext_reg[61]  ( .D(reg_out[61]), .CK(clk), .Q(Plaintext[61]) );
  DFF_X1 \Plaintext_reg[60]  ( .D(reg_out[60]), .CK(clk), .Q(Plaintext[60]) );
  DFF_X1 \Plaintext_reg[59]  ( .D(reg_out[59]), .CK(clk), .Q(Plaintext[59]) );
  DFF_X1 \Plaintext_reg[58]  ( .D(reg_out[58]), .CK(clk), .Q(Plaintext[58]) );
  DFF_X1 \Plaintext_reg[57]  ( .D(reg_out[57]), .CK(clk), .Q(Plaintext[57]) );
  DFF_X1 \Plaintext_reg[56]  ( .D(reg_out[56]), .CK(clk), .Q(Plaintext[56]) );
  DFF_X1 \Plaintext_reg[55]  ( .D(reg_out[55]), .CK(clk), .Q(Plaintext[55]) );
  DFF_X1 \Plaintext_reg[54]  ( .D(reg_out[54]), .CK(clk), .Q(Plaintext[54]) );
  DFF_X1 \Plaintext_reg[53]  ( .D(reg_out[53]), .CK(clk), .Q(Plaintext[53]) );
  DFF_X1 \Plaintext_reg[52]  ( .D(reg_out[52]), .CK(clk), .Q(Plaintext[52]) );
  DFF_X1 \Plaintext_reg[51]  ( .D(reg_out[51]), .CK(clk), .Q(Plaintext[51]) );
  DFF_X1 \Plaintext_reg[50]  ( .D(reg_out[50]), .CK(clk), .Q(Plaintext[50]) );
  DFF_X1 \Plaintext_reg[49]  ( .D(reg_out[49]), .CK(clk), .Q(Plaintext[49]) );
  DFF_X1 \Plaintext_reg[48]  ( .D(reg_out[48]), .CK(clk), .Q(Plaintext[48]) );
  DFF_X1 \Plaintext_reg[47]  ( .D(reg_out[47]), .CK(clk), .Q(Plaintext[47]) );
  DFF_X1 \Plaintext_reg[46]  ( .D(reg_out[46]), .CK(clk), .Q(Plaintext[46]) );
  DFF_X1 \Plaintext_reg[45]  ( .D(reg_out[45]), .CK(clk), .Q(Plaintext[45]) );
  DFF_X1 \Plaintext_reg[44]  ( .D(reg_out[44]), .CK(clk), .Q(Plaintext[44]) );
  DFF_X1 \Plaintext_reg[43]  ( .D(reg_out[43]), .CK(clk), .Q(Plaintext[43]) );
  DFF_X1 \Plaintext_reg[42]  ( .D(reg_out[42]), .CK(clk), .Q(Plaintext[42]) );
  DFF_X1 \Plaintext_reg[41]  ( .D(reg_out[41]), .CK(clk), .Q(Plaintext[41]) );
  DFF_X1 \Plaintext_reg[40]  ( .D(reg_out[40]), .CK(clk), .Q(Plaintext[40]) );
  DFF_X1 \Plaintext_reg[39]  ( .D(reg_out[39]), .CK(clk), .Q(Plaintext[39]) );
  DFF_X1 \Plaintext_reg[38]  ( .D(reg_out[38]), .CK(clk), .Q(Plaintext[38]) );
  DFF_X1 \Plaintext_reg[37]  ( .D(reg_out[37]), .CK(clk), .Q(Plaintext[37]) );
  DFF_X1 \Plaintext_reg[36]  ( .D(reg_out[36]), .CK(clk), .Q(Plaintext[36]) );
  DFF_X1 \Plaintext_reg[35]  ( .D(reg_out[35]), .CK(clk), .Q(Plaintext[35]) );
  DFF_X1 \Plaintext_reg[33]  ( .D(reg_out[33]), .CK(clk), .Q(Plaintext[33]) );
  DFF_X1 \Plaintext_reg[32]  ( .D(reg_out[32]), .CK(clk), .Q(Plaintext[32]) );
  DFF_X1 \Plaintext_reg[31]  ( .D(reg_out[31]), .CK(clk), .Q(Plaintext[31]) );
  DFF_X1 \Plaintext_reg[30]  ( .D(reg_out[30]), .CK(clk), .Q(Plaintext[30]) );
  DFF_X1 \Plaintext_reg[29]  ( .D(reg_out[29]), .CK(clk), .Q(Plaintext[29]) );
  DFF_X1 \Plaintext_reg[28]  ( .D(reg_out[28]), .CK(clk), .Q(Plaintext[28]) );
  DFF_X1 \Plaintext_reg[27]  ( .D(reg_out[27]), .CK(clk), .Q(Plaintext[27]) );
  DFF_X1 \Plaintext_reg[26]  ( .D(reg_out[26]), .CK(clk), .Q(Plaintext[26]) );
  DFF_X1 \Plaintext_reg[24]  ( .D(reg_out[24]), .CK(clk), .Q(Plaintext[24]) );
  DFF_X1 \Plaintext_reg[23]  ( .D(reg_out[23]), .CK(clk), .Q(Plaintext[23]) );
  DFF_X1 \Plaintext_reg[22]  ( .D(reg_out[22]), .CK(clk), .Q(Plaintext[22]) );
  DFF_X1 \Plaintext_reg[21]  ( .D(reg_out[21]), .CK(clk), .Q(Plaintext[21]) );
  DFF_X1 \Plaintext_reg[20]  ( .D(reg_out[20]), .CK(clk), .Q(Plaintext[20]) );
  DFF_X1 \Plaintext_reg[19]  ( .D(reg_out[19]), .CK(clk), .Q(Plaintext[19]) );
  DFF_X1 \Plaintext_reg[18]  ( .D(reg_out[18]), .CK(clk), .Q(Plaintext[18]) );
  DFF_X1 \Plaintext_reg[17]  ( .D(reg_out[17]), .CK(clk), .Q(Plaintext[17]) );
  DFF_X1 \Plaintext_reg[16]  ( .D(reg_out[16]), .CK(clk), .Q(Plaintext[16]) );
  DFF_X1 \Plaintext_reg[15]  ( .D(reg_out[15]), .CK(clk), .Q(Plaintext[15]) );
  DFF_X1 \Plaintext_reg[14]  ( .D(reg_out[14]), .CK(clk), .Q(Plaintext[14]) );
  DFF_X1 \Plaintext_reg[13]  ( .D(reg_out[13]), .CK(clk), .Q(Plaintext[13]) );
  DFF_X1 \Plaintext_reg[12]  ( .D(reg_out[12]), .CK(clk), .Q(Plaintext[12]) );
  DFF_X1 \Plaintext_reg[11]  ( .D(reg_out[11]), .CK(clk), .Q(Plaintext[11]) );
  DFF_X1 \Plaintext_reg[10]  ( .D(reg_out[10]), .CK(clk), .Q(Plaintext[10]) );
  DFF_X1 \Plaintext_reg[9]  ( .D(reg_out[9]), .CK(clk), .Q(Plaintext[9]) );
  DFF_X1 \Plaintext_reg[8]  ( .D(reg_out[8]), .CK(clk), .Q(Plaintext[8]) );
  DFF_X1 \Plaintext_reg[7]  ( .D(reg_out[7]), .CK(clk), .Q(Plaintext[7]) );
  DFF_X1 \Plaintext_reg[6]  ( .D(reg_out[6]), .CK(clk), .Q(Plaintext[6]) );
  DFF_X1 \Plaintext_reg[5]  ( .D(reg_out[5]), .CK(clk), .Q(Plaintext[5]) );
  DFF_X1 \Plaintext_reg[4]  ( .D(reg_out[4]), .CK(clk), .Q(Plaintext[4]) );
  DFF_X1 \Plaintext_reg[3]  ( .D(reg_out[3]), .CK(clk), .Q(Plaintext[3]) );
  DFF_X1 \Plaintext_reg[2]  ( .D(reg_out[2]), .CK(clk), .Q(Plaintext[2]) );
  DFF_X1 \Plaintext_reg[1]  ( .D(reg_out[1]), .CK(clk), .Q(Plaintext[1]) );
  DFF_X1 \Plaintext_reg[0]  ( .D(reg_out[0]), .CK(clk), .Q(Plaintext[0]) );
  DFF_X1 \Plaintext_reg[95]  ( .D(reg_out[95]), .CK(clk), .Q(Plaintext[95]) );
  DFF_X1 \reg_key_reg[127]  ( .D(Key[127]), .CK(clk), .Q(reg_key[127]) );
  DFF_X1 \reg_key_reg[121]  ( .D(Key[121]), .CK(clk), .Q(reg_key[121]) );
  DFF_X1 \reg_key_reg[16]  ( .D(Key[16]), .CK(clk), .Q(reg_key[16]) );
  DFF_X1 \reg_key_reg[56]  ( .D(Key[56]), .CK(clk), .Q(reg_key[56]) );
  DFF_X1 \reg_key_reg[104]  ( .D(Key[104]), .CK(clk), .Q(reg_key[104]) );
  DFF_X1 \reg_key_reg[20]  ( .D(Key[20]), .CK(clk), .Q(reg_key[20]) );
  DFF_X1 \reg_key_reg[21]  ( .D(Key[21]), .CK(clk), .Q(reg_key[21]) );
  DFF_X1 \reg_key_reg[7]  ( .D(Key[7]), .CK(clk), .Q(reg_key[7]) );
  DFF_X1 \reg_key_reg[110]  ( .D(Key[110]), .CK(clk), .Q(reg_key[110]) );
  DFF_X1 \reg_key_reg[80]  ( .D(Key[80]), .CK(clk), .Q(reg_key[80]) );
  DFF_X1 \reg_key_reg[134]  ( .D(Key[134]), .CK(clk), .Q(reg_key[134]) );
  DFF_X1 \reg_key_reg[37]  ( .D(Key[37]), .CK(clk), .Q(reg_key[37]) );
  DFF_X1 \reg_key_reg[163]  ( .D(Key[163]), .CK(clk), .Q(reg_key[163]) );
  DFF_X1 \reg_key_reg[187]  ( .D(Key[187]), .CK(clk), .Q(reg_key[187]) );
  DFF_X1 \reg_key_reg[83]  ( .D(Key[83]), .CK(clk), .Q(reg_key[83]) );
  DFF_X1 \reg_key_reg[132]  ( .D(Key[132]), .CK(clk), .Q(reg_key[132]) );
  DFF_X1 \reg_key_reg[164]  ( .D(Key[164]), .CK(clk), .Q(reg_key[164]) );
  DFF_X1 \reg_key_reg[177]  ( .D(Key[177]), .CK(clk), .Q(reg_key[177]) );
  DFF_X1 \reg_key_reg[55]  ( .D(Key[55]), .CK(clk), .Q(reg_key[55]) );
  DFF_X1 \reg_key_reg[103]  ( .D(Key[103]), .CK(clk), .Q(reg_key[103]) );
  DFF_X1 \reg_key_reg[52]  ( .D(Key[52]), .CK(clk), .Q(reg_key[52]) );
  DFF_X1 \reg_key_reg[39]  ( .D(Key[39]), .CK(clk), .Q(reg_key[39]) );
  DFF_X1 \reg_key_reg[62]  ( .D(Key[62]), .CK(clk), .Q(reg_key[62]) );
  DFF_X1 \reg_key_reg[145]  ( .D(Key[145]), .CK(clk), .Q(reg_key[145]) );
  DFF_X1 \reg_key_reg[182]  ( .D(Key[182]), .CK(clk), .Q(reg_key[182]) );
  DFF_X1 \reg_key_reg[73]  ( .D(Key[73]), .CK(clk), .Q(reg_key[73]) );
  DFF_X1 \reg_key_reg[26]  ( .D(Key[26]), .CK(clk), .Q(reg_key[26]) );
  DFF_X1 \reg_key_reg[168]  ( .D(Key[168]), .CK(clk), .Q(reg_key[168]) );
  DFF_X1 \reg_key_reg[169]  ( .D(Key[169]), .CK(clk), .Q(reg_key[169]) );
  DFF_X1 \reg_key_reg[49]  ( .D(Key[49]), .CK(clk), .Q(reg_key[49]) );
  DFF_X1 \reg_key_reg[157]  ( .D(Key[157]), .CK(clk), .Q(reg_key[157]) );
  DFF_X1 \reg_key_reg[178]  ( .D(Key[178]), .CK(clk), .Q(reg_key[178]) );
  DFF_X1 \reg_key_reg[70]  ( .D(Key[70]), .CK(clk), .Q(reg_key[70]) );
  DFF_X1 \reg_key_reg[29]  ( .D(Key[29]), .CK(clk), .Q(reg_key[29]) );
  DFF_X1 \reg_key_reg[141]  ( .D(Key[141]), .CK(clk), .Q(reg_key[141]) );
  DFF_X1 \reg_key_reg[79]  ( .D(Key[79]), .CK(clk), .Q(reg_key[79]) );
  DFF_X1 \reg_key_reg[167]  ( .D(Key[167]), .CK(clk), .Q(reg_key[167]) );
  DFF_X1 \reg_key_reg[115]  ( .D(Key[115]), .CK(clk), .Q(reg_key[115]) );
  DFF_X1 \reg_key_reg[151]  ( .D(Key[151]), .CK(clk), .Q(reg_key[151]) );
  DFF_X1 \reg_key_reg[188]  ( .D(Key[188]), .CK(clk), .Q(reg_key[188]) );
  DFF_X1 \reg_key_reg[61]  ( .D(Key[61]), .CK(clk), .Q(reg_key[61]) );
  DFF_X1 \reg_key_reg[58]  ( .D(Key[58]), .CK(clk), .Q(reg_key[58]) );
  DFF_X1 \reg_key_reg[161]  ( .D(Key[161]), .CK(clk), .Q(reg_key[161]) );
  DFF_X1 \reg_key_reg[44]  ( .D(Key[44]), .CK(clk), .Q(reg_key[44]) );
  DFF_X1 \reg_key_reg[91]  ( .D(Key[91]), .CK(clk), .Q(reg_key[91]) );
  DFF_X1 \reg_key_reg[172]  ( .D(Key[172]), .CK(clk), .Q(reg_key[172]) );
  DFF_X1 \reg_key_reg[116]  ( .D(Key[116]), .CK(clk), .Q(reg_key[116]) );
  DFF_X1 \reg_key_reg[35]  ( .D(Key[35]), .CK(clk), .Q(reg_key[35]) );
  DFF_X1 \reg_key_reg[59]  ( .D(Key[59]), .CK(clk), .Q(reg_key[59]) );
  DFF_X1 \reg_key_reg[154]  ( .D(Key[154]), .CK(clk), .Q(reg_key[154]) );
  DFF_X1 \reg_key_reg[64]  ( .D(Key[64]), .CK(clk), .Q(reg_key[64]) );
  DFF_X1 \reg_key_reg[51]  ( .D(Key[51]), .CK(clk), .Q(reg_key[51]) );
  DFF_X1 \reg_key_reg[13]  ( .D(Key[13]), .CK(clk), .Q(reg_key[13]) );
  DFF_X1 \reg_key_reg[173]  ( .D(Key[173]), .CK(clk), .Q(reg_key[173]) );
  DFF_X1 \reg_key_reg[185]  ( .D(Key[185]), .CK(clk), .Q(reg_key[185]) );
  DFF_X1 \reg_key_reg[130]  ( .D(Key[130]), .CK(clk), .Q(reg_key[130]) );
  DFF_X1 \reg_key_reg[140]  ( .D(Key[140]), .CK(clk), .Q(reg_key[140]) );
  DFF_X1 \reg_key_reg[5]  ( .D(Key[5]), .CK(clk), .Q(reg_key[5]) );
  DFF_X1 \reg_key_reg[65]  ( .D(Key[65]), .CK(clk), .Q(reg_key[65]) );
  DFF_X1 \reg_key_reg[191]  ( .D(Key[191]), .CK(clk), .Q(reg_key[191]) );
  DFF_X1 \reg_key_reg[24]  ( .D(Key[24]), .CK(clk), .Q(reg_key[24]) );
  DFF_X1 \reg_key_reg[89]  ( .D(Key[89]), .CK(clk), .Q(reg_key[89]) );
  DFF_X1 \reg_key_reg[33]  ( .D(Key[33]), .CK(clk), .Q(reg_key[33]) );
  DFF_X1 \reg_key_reg[36]  ( .D(Key[36]), .CK(clk), .Q(reg_key[36]) );
  DFF_X1 \reg_key_reg[63]  ( .D(Key[63]), .CK(clk), .Q(reg_key[63]) );
  DFF_X1 \reg_key_reg[87]  ( .D(Key[87]), .CK(clk), .Q(reg_key[87]) );
  DFF_X1 \reg_key_reg[112]  ( .D(Key[112]), .CK(clk), .Q(reg_key[112]) );
  DFF_X1 \reg_key_reg[71]  ( .D(Key[71]), .CK(clk), .Q(reg_key[71]) );
  DFF_X1 \reg_key_reg[41]  ( .D(Key[41]), .CK(clk), .Q(reg_key[41]) );
  DFF_X1 \reg_key_reg[19]  ( .D(Key[19]), .CK(clk), .Q(reg_key[19]) );
  DFF_X1 \reg_key_reg[8]  ( .D(Key[8]), .CK(clk), .Q(reg_key[8]) );
  DFF_X1 \reg_key_reg[53]  ( .D(Key[53]), .CK(clk), .Q(reg_key[53]) );
  DFF_X1 \reg_key_reg[92]  ( .D(Key[92]), .CK(clk), .Q(reg_key[92]) );
  DFF_X1 \reg_key_reg[90]  ( .D(Key[90]), .CK(clk), .Q(reg_key[90]) );
  DFF_X1 \reg_key_reg[95]  ( .D(Key[95]), .CK(clk), .Q(reg_key[95]) );
  DFF_X1 \reg_key_reg[109]  ( .D(Key[109]), .CK(clk), .Q(reg_key[109]) );
  DFF_X1 \reg_key_reg[133]  ( .D(Key[133]), .CK(clk), .Q(reg_key[133]) );
  DFF_X1 \reg_key_reg[125]  ( .D(Key[125]), .CK(clk), .Q(reg_key[125]) );
  DFF_X1 \reg_key_reg[25]  ( .D(Key[25]), .CK(clk), .Q(reg_key[25]) );
  DFF_X1 \reg_key_reg[68]  ( .D(Key[68]), .CK(clk), .Q(reg_key[68]) );
  DFF_X1 \reg_key_reg[105]  ( .D(Key[105]), .CK(clk), .Q(reg_key[105]) );
  DFF_X1 \reg_key_reg[120]  ( .D(Key[120]), .CK(clk), .Q(reg_key[120]) );
  DFF_X1 \reg_key_reg[175]  ( .D(Key[175]), .CK(clk), .Q(reg_key[175]) );
  DFF_X1 \reg_key_reg[153]  ( .D(Key[153]), .CK(clk), .Q(reg_key[153]) );
  DFF_X1 \reg_key_reg[118]  ( .D(Key[118]), .CK(clk), .Q(reg_key[118]) );
  DFF_X1 \reg_key_reg[94]  ( .D(Key[94]), .CK(clk), .Q(reg_key[94]) );
  DFF_X1 \reg_key_reg[150]  ( .D(Key[150]), .CK(clk), .Q(reg_key[150]) );
  DFF_X1 \reg_key_reg[174]  ( .D(Key[174]), .CK(clk), .Q(reg_key[174]) );
  DFF_X1 \reg_key_reg[93]  ( .D(Key[93]), .CK(clk), .Q(reg_key[93]) );
  DFF_X1 \Plaintext_reg[84]  ( .D(reg_out[84]), .CK(clk), .Q(Plaintext[84]) );
  DFF_X1 \Plaintext_reg[161]  ( .D(reg_out[161]), .CK(clk), .Q(Plaintext[161])
         );
  DFF_X1 \Plaintext_reg[129]  ( .D(reg_out[129]), .CK(clk), .Q(Plaintext[129])
         );
  DFF_X1 \reg_key_reg[190]  ( .D(Key[190]), .CK(clk), .Q(reg_key[190]) );
  DFF_X1 \reg_key_reg[183]  ( .D(Key[183]), .CK(clk), .Q(reg_key[183]) );
  DFF_X1 \reg_key_reg[181]  ( .D(Key[181]), .CK(clk), .Q(reg_key[181]) );
  DFF_X1 \reg_key_reg[179]  ( .D(Key[179]), .CK(clk), .Q(reg_key[179]) );
  DFF_X1 \reg_key_reg[176]  ( .D(Key[176]), .CK(clk), .Q(reg_key[176]) );
  DFF_X1 \reg_key_reg[170]  ( .D(Key[170]), .CK(clk), .Q(reg_key[170]) );
  DFF_X1 \reg_key_reg[166]  ( .D(Key[166]), .CK(clk), .Q(reg_key[166]) );
  DFF_X1 \reg_key_reg[165]  ( .D(Key[165]), .CK(clk), .Q(reg_key[165]) );
  DFF_X1 \reg_key_reg[159]  ( .D(Key[159]), .CK(clk), .Q(reg_key[159]) );
  DFF_X1 \reg_key_reg[158]  ( .D(Key[158]), .CK(clk), .Q(reg_key[158]) );
  DFF_X1 \reg_key_reg[156]  ( .D(Key[156]), .CK(clk), .Q(reg_key[156]) );
  DFF_X1 \reg_key_reg[155]  ( .D(Key[155]), .CK(clk), .Q(reg_key[155]) );
  DFF_X1 \reg_key_reg[152]  ( .D(Key[152]), .CK(clk), .Q(reg_key[152]) );
  DFF_X1 \reg_key_reg[149]  ( .D(Key[149]), .CK(clk), .Q(reg_key[149]) );
  DFF_X1 \reg_key_reg[148]  ( .D(Key[148]), .CK(clk), .Q(reg_key[148]) );
  DFF_X1 \reg_key_reg[147]  ( .D(Key[147]), .CK(clk), .Q(reg_key[147]) );
  DFF_X1 \reg_key_reg[146]  ( .D(Key[146]), .CK(clk), .Q(reg_key[146]) );
  DFF_X1 \reg_key_reg[144]  ( .D(Key[144]), .CK(clk), .Q(reg_key[144]) );
  DFF_X1 \reg_key_reg[143]  ( .D(Key[143]), .CK(clk), .Q(reg_key[143]) );
  DFF_X1 \reg_key_reg[142]  ( .D(Key[142]), .CK(clk), .Q(reg_key[142]) );
  DFF_X1 \reg_key_reg[137]  ( .D(Key[137]), .CK(clk), .Q(reg_key[137]) );
  DFF_X1 \reg_key_reg[135]  ( .D(Key[135]), .CK(clk), .Q(reg_key[135]) );
  DFF_X1 \reg_key_reg[128]  ( .D(Key[128]), .CK(clk), .Q(reg_key[128]) );
  DFF_X1 \reg_key_reg[126]  ( .D(Key[126]), .CK(clk), .Q(reg_key[126]) );
  DFF_X1 \reg_key_reg[119]  ( .D(Key[119]), .CK(clk), .Q(reg_key[119]) );
  DFF_X1 \reg_key_reg[117]  ( .D(Key[117]), .CK(clk), .Q(reg_key[117]) );
  DFF_X1 \reg_key_reg[114]  ( .D(Key[114]), .CK(clk), .Q(reg_key[114]) );
  DFF_X1 \reg_key_reg[113]  ( .D(Key[113]), .CK(clk), .Q(reg_key[113]) );
  DFF_X1 \reg_key_reg[108]  ( .D(Key[108]), .CK(clk), .Q(reg_key[108]) );
  DFF_X1 \reg_key_reg[106]  ( .D(Key[106]), .CK(clk), .Q(reg_key[106]) );
  DFF_X1 \reg_key_reg[102]  ( .D(Key[102]), .CK(clk), .Q(reg_key[102]) );
  DFF_X1 \reg_key_reg[99]  ( .D(Key[99]), .CK(clk), .Q(reg_key[99]) );
  DFF_X1 \reg_key_reg[98]  ( .D(Key[98]), .CK(clk), .Q(reg_key[98]) );
  DFF_X1 \reg_key_reg[97]  ( .D(Key[97]), .CK(clk), .Q(reg_key[97]) );
  DFF_X1 \reg_key_reg[96]  ( .D(Key[96]), .CK(clk), .Q(reg_key[96]) );
  DFF_X1 \reg_key_reg[88]  ( .D(Key[88]), .CK(clk), .Q(reg_key[88]) );
  DFF_X1 \reg_key_reg[86]  ( .D(Key[86]), .CK(clk), .Q(reg_key[86]) );
  DFF_X1 \reg_key_reg[85]  ( .D(Key[85]), .CK(clk), .Q(reg_key[85]) );
  DFF_X1 \reg_key_reg[82]  ( .D(Key[82]), .CK(clk), .Q(reg_key[82]) );
  DFF_X1 \reg_key_reg[76]  ( .D(Key[76]), .CK(clk), .Q(reg_key[76]) );
  DFF_X1 \reg_key_reg[75]  ( .D(Key[75]), .CK(clk), .Q(reg_key[75]) );
  DFF_X1 \reg_key_reg[74]  ( .D(Key[74]), .CK(clk), .Q(reg_key[74]) );
  DFF_X1 \reg_key_reg[66]  ( .D(Key[66]), .CK(clk), .Q(reg_key[66]) );
  DFF_X1 \reg_key_reg[60]  ( .D(Key[60]), .CK(clk), .Q(reg_key[60]) );
  DFF_X1 \reg_key_reg[54]  ( .D(Key[54]), .CK(clk), .Q(reg_key[54]) );
  DFF_X1 \reg_key_reg[43]  ( .D(Key[43]), .CK(clk), .Q(reg_key[43]) );
  DFF_X1 \reg_key_reg[38]  ( .D(Key[38]), .CK(clk), .Q(reg_key[38]) );
  DFF_X1 \reg_key_reg[34]  ( .D(Key[34]), .CK(clk), .Q(reg_key[34]) );
  DFF_X1 \reg_key_reg[28]  ( .D(Key[28]), .CK(clk), .Q(reg_key[28]) );
  DFF_X1 \reg_key_reg[27]  ( .D(Key[27]), .CK(clk), .Q(reg_key[27]) );
  DFF_X1 \reg_key_reg[18]  ( .D(Key[18]), .CK(clk), .Q(reg_key[18]) );
  DFF_X1 \reg_key_reg[15]  ( .D(Key[15]), .CK(clk), .Q(reg_key[15]) );
  DFF_X1 \reg_key_reg[14]  ( .D(Key[14]), .CK(clk), .Q(reg_key[14]) );
  DFF_X1 \reg_key_reg[12]  ( .D(Key[12]), .CK(clk), .Q(reg_key[12]) );
  DFF_X1 \reg_key_reg[10]  ( .D(Key[10]), .CK(clk), .Q(reg_key[10]) );
  DFF_X1 \reg_key_reg[9]  ( .D(Key[9]), .CK(clk), .Q(reg_key[9]) );
  DFF_X1 \reg_key_reg[4]  ( .D(Key[4]), .CK(clk), .Q(reg_key[4]) );
  DFF_X1 \reg_key_reg[1]  ( .D(Key[1]), .CK(clk), .Q(reg_key[1]) );
  DFF_X1 \reg_key_reg[84]  ( .D(Key[84]), .CK(clk), .Q(reg_key[84]) );
  DFF_X1 \reg_key_reg[186]  ( .D(Key[186]), .CK(clk), .Q(reg_key[186]) );
  DFF_X1 \reg_key_reg[184]  ( .D(Key[184]), .CK(clk), .Q(reg_key[184]) );
  DFF_X1 \reg_key_reg[162]  ( .D(Key[162]), .CK(clk), .Q(reg_key[162]) );
  DFF_X1 \reg_key_reg[139]  ( .D(Key[139]), .CK(clk), .Q(reg_key[139]) );
  DFF_X1 \reg_key_reg[138]  ( .D(Key[138]), .CK(clk), .Q(reg_key[138]) );
  DFF_X1 \reg_key_reg[123]  ( .D(Key[123]), .CK(clk), .Q(reg_key[123]) );
  DFF_X1 \reg_key_reg[111]  ( .D(Key[111]), .CK(clk), .Q(reg_key[111]) );
  DFF_X1 \reg_key_reg[107]  ( .D(Key[107]), .CK(clk), .Q(reg_key[107]) );
  DFF_X1 \reg_key_reg[69]  ( .D(Key[69]), .CK(clk), .Q(reg_key[69]) );
  DFF_X1 \reg_key_reg[48]  ( .D(Key[48]), .CK(clk), .Q(reg_key[48]) );
  DFF_X1 \reg_key_reg[32]  ( .D(Key[32]), .CK(clk), .Q(reg_key[32]) );
  DFF_X1 \reg_key_reg[23]  ( .D(Key[23]), .CK(clk), .Q(reg_key[23]) );
  DFF_X1 \reg_key_reg[22]  ( .D(Key[22]), .CK(clk), .Q(reg_key[22]) );
  DFF_X1 \reg_key_reg[11]  ( .D(Key[11]), .CK(clk), .Q(reg_key[11]) );
  DFF_X1 \reg_key_reg[124]  ( .D(Key[124]), .CK(clk), .Q(reg_key[124]) );
  DFF_X1 \reg_key_reg[72]  ( .D(Key[72]), .CK(clk), .Q(reg_key[72]) );
  DFF_X1 \reg_key_reg[46]  ( .D(Key[46]), .CK(clk), .Q(reg_key[46]) );
  DFF_X1 \reg_key_reg[45]  ( .D(Key[45]), .CK(clk), .Q(reg_key[45]) );
  DFF_X1 \reg_key_reg[40]  ( .D(Key[40]), .CK(clk), .Q(reg_key[40]) );
  DFF_X1 \reg_key_reg[2]  ( .D(Key[2]), .CK(clk), .Q(reg_key[2]) );
  DFF_X1 \reg_key_reg[0]  ( .D(Key[0]), .CK(clk), .Q(reg_key[0]) );
  DFF_X1 \reg_key_reg[81]  ( .D(Key[81]), .CK(clk), .Q(reg_key[81]) );
  DFF_X1 \reg_key_reg[129]  ( .D(Key[129]), .CK(clk), .Q(reg_key[129]) );
  DFF_X1 \reg_key_reg[122]  ( .D(Key[122]), .CK(clk), .Q(reg_key[122]) );
  DFF_X1 \reg_key_reg[6]  ( .D(Key[6]), .CK(clk), .Q(reg_key[6]) );
  DFF_X1 \reg_key_reg[136]  ( .D(Key[136]), .CK(clk), .Q(reg_key[136]) );
  DFF_X1 \reg_key_reg[57]  ( .D(Key[57]), .CK(clk), .Q(reg_key[57]) );
  DFF_X1 \reg_key_reg[78]  ( .D(Key[78]), .CK(clk), .Q(reg_key[78]) );
  DFF_X1 \reg_key_reg[101]  ( .D(Key[101]), .CK(clk), .Q(reg_key[101]) );
  DFF_X1 \reg_key_reg[31]  ( .D(Key[31]), .CK(clk), .Q(reg_key[31]) );
  DFF_X1 \reg_key_reg[42]  ( .D(Key[42]), .CK(clk), .Q(reg_key[42]) );
  DFF_X1 \reg_key_reg[131]  ( .D(Key[131]), .CK(clk), .Q(reg_key[131]) );
  DFF_X1 \reg_key_reg[30]  ( .D(Key[30]), .CK(clk), .Q(reg_key[30]) );
  DFF_X1 \reg_key_reg[189]  ( .D(Key[189]), .CK(clk), .Q(reg_key[189]) );
  DFF_X1 \reg_key_reg[3]  ( .D(Key[3]), .CK(clk), .Q(reg_key[3]) );
  DFF_X1 \reg_key_reg[180]  ( .D(Key[180]), .CK(clk), .Q(reg_key[180]) );
  DFF_X1 \reg_key_reg[171]  ( .D(Key[171]), .CK(clk), .Q(reg_key[171]) );
  DFFRS_X1 \Plaintext_reg[188]  ( .D(reg_out[188]), .CK(clk), .RN(1'b1), .SN(
        1'b1), .Q(Plaintext[188]) );
  DFFRS_X1 \Plaintext_reg[25]  ( .D(reg_out[25]), .CK(clk), .RN(1'b1), .SN(
        1'b1), .Q(Plaintext[25]) );
  DFF_X1 \Plaintext_reg[167]  ( .D(reg_out[167]), .CK(clk), .Q(Plaintext[167])
         );
  DFF_X1 \Plaintext_reg[114]  ( .D(reg_out[114]), .CK(clk), .Q(Plaintext[114])
         );
  SPEEDY_Rounds5_0 SPEEDY_instance ( .Ciphertext(reg_in), .Key(reg_key), 
        .Plaintext(reg_out) );
  DFFRS_X1 \Plaintext_reg[62]  ( .D(reg_out[62]), .CK(clk), .RN(1'b1), .SN(
        1'b1), .Q(Plaintext[62]) );
  DFFS_X1 \Plaintext_reg[155]  ( .D(reg_out[155]), .CK(clk), .SN(1'b1), .Q(
        Plaintext[155]) );
  DFFRS_X1 \Plaintext_reg[34]  ( .D(reg_out[34]), .CK(clk), .RN(1'b1), .SN(
        1'b1), .Q(Plaintext[34]) );
  DFF_X1 \Plaintext_reg[181]  ( .D(reg_out[181]), .CK(clk), .Q(Plaintext[181])
         );
  DFF_X1 \Plaintext_reg[92]  ( .D(reg_out[92]), .CK(clk), .Q(Plaintext[92]) );
endmodule

