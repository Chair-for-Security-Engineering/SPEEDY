
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_SPEEDY_Top is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_SPEEDY_Top;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Rounds6_0 is

   port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : out
         std_logic_vector (191 downto 0));

end SPEEDY_Rounds6_0;

architecture SYN_Behavioral of SPEEDY_Rounds6_0 is

   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32
      , n34, n38, n39, n40, n41, n42, n44, n45, n46, n47, n48, n51, n52, n55, 
      n58, n59, n60, n61, n62, n66, n68, n69, n70, n71, n72, n73, n75, n76, n77
      , n78, n79, n81, n82, n85, n87, n88, n89, n92, n95, n96, n97, n98, n100, 
      n101, n102, n103, n104, n107, n108, n109, n111, n112, n113, n114, n115, 
      n118, n119, n120, n121, n122, n123, n125, n126, n127, n128, n129, n131, 
      n133, n135, n136, n137, n138, n139, n140, n141, n142, n144, n145, n146, 
      n147, n148, n149, n151, n152, n153, n155, n156, n158, n159, n160, n161, 
      n162, n164, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n185, n187, n188, n189, n190, n191, n194, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n223, n227, n231, n232, n233, n238, n239, 
      n240, n244, n245, n246, n248, n249, n250, n257, n260, n261, n262, n263, 
      n264, n266, n267, n268, n269, n270, n271, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n287, n288, n290, n291, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n307, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n343, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n361, 
      n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, 
      n374, n376, n377, n379, n380, n381, n382, n383, n385, n386, n387, n388, 
      n389, n391, n392, n394, n395, n396, n397, n398, n399, n400, n401, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n424, n425, n426, n427, n428, 
      n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, 
      n441, n442, n443, n444, n445, n447, n448, n449, n450, n451, n452, n453, 
      n454, n455, n456, n457, n458, n459, n462, n463, n464, n465, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n477, n478, n479, n480, n481, 
      n483, n484, n486, n488, n491, n492, n493, n494, n495, n496, n498, n499, 
      n500, n501, n502, n504, n505, n507, n508, n509, n510, n511, n512, n513, 
      n514, n515, n516, n517, n519, n520, n521, n522, n523, n524, n525, n526, 
      n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, 
      n539, n540, n541, n542, n543, n545, n546, n547, n548, n549, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, 
      n578, n579, n580, n581, n584, n585, n586, n587, n588, n589, n590, n593, 
      n594, n595, n596, n597, n598, n599, n600, n602, n603, n605, n606, n607, 
      n608, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, 
      n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, 
      n634, n635, n636, n637, n638, n640, n641, n642, n644, n645, n646, n647, 
      n648, n649, n650, n651, n652, n654, n655, n656, n657, n658, n659, n660, 
      n661, n662, n663, n664, n665, n667, n668, n669, n670, n671, n672, n673, 
      n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, 
      n686, n687, n688, n689, n690, n692, n693, n695, n696, n697, n698, n699, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n718, n719, n720, n721, n722, n723, n725, n726, n727, n728, 
      n729, n730, n731, n732, n733, n734, n735, n736, n737, n740, n741, n742, 
      n743, n744, n746, n747, n749, n751, n752, n753, n754, n755, n756, n757, 
      n758, n759, n760, n762, n763, n764, n765, n766, n767, n768, n769, n770, 
      n771, n772, n773, n775, n776, n777, n778, n779, n780, n781, n782, n784, 
      n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, 
      n798, n799, n800, n801, n802, n804, n806, n807, n808, n809, n810, n812, 
      n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, 
      n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, 
      n837, n838, n839, n840, n841, n842, n843, n845, n847, n848, n849, n852, 
      n853, n854, n855, n856, n857, n859, n860, n861, n862, n863, n864, n867, 
      n868, n869, n870, n871, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n905, 
      n906, n907, n908, n909, n910, n911, n912, n914, n915, n916, n918, n919, 
      n920, n921, n923, n924, n925, n927, n928, n929, n930, n931, n932, n933, 
      n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, 
      n946, n947, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, 
      n959, n960, n961, n962, n963, n965, n966, n967, n968, n969, n971, n972, 
      n973, n974, n975, n976, n977, n978, n979, n980, n981, n984, n985, n986, 
      n987, n988, n989, n990, n991, n992, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1032, n1033, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1065, n1066, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
      n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
      n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1095, 
      n1096, n1097, n1098, n1099, n1100, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
      n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, 
      n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, 
      n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, 
      n1148, n1149, n1150, n1152, n1153, n1154, n1155, n1156, n1158, n1159, 
      n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
      n1170, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, 
      n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, 
      n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, 
      n1202, n1203, n1204, n1205, n1206, n1208, n1210, n1211, n1212, n1214, 
      n1215, n1216, n1217, n1218, n1219, n1220, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1235, n1237, n1238, 
      n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, 
      n1249, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
      n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, 
      n1272, n1273, n1275, n1276, n1279, n1280, n1281, n1282, n1283, n1284, 
      n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, 
      n1295, n1296, n1297, n1299, n1300, n1301, n1302, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
      n1328, n1329, n1330, n1331, n1332, n1334, n1335, n1336, n1337, n1338, 
      n1339, n1340, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, 
      n1351, n1352, n1353, n1355, n1357, n1358, n1359, n1361, n1362, n1363, 
      n1364, n1365, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, 
      n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, 
      n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, 
      n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, 
      n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, 
      n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
      n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, 
      n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
      n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, 
      n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
      n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, 
      n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, 
      n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, 
      n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, 
      n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, 
      n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1526, n1527, n1528, 
      n1530, n1531, n1532, n1534, n1535, n1536, n1537, n1538, n1539, n1540, 
      n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, 
      n1551, n1552, n1553, n1554, n1556, n1557, n1558, n1559, n1561, n1562, 
      n1563, n1564, n1566, n1568, n1569, n1570, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1604, n1605, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
      n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
      n1649, n1653, n1654, n1655, n1656, n1658, n1660, n1661, n1662, n1663, 
      n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, 
      n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, 
      n1684, n1685, n1686, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1718, 
      n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
      n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
      n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, 
      n1751, n1752, n1753, n1754, n1755, n1757, n1758, n1759, n1760, n1761, 
      n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, 
      n1772, n1773, n1774, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1801, n1802, n1803, 
      n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, 
      n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, 
      n1824, n1825, n1826, n1827, n1828, n1830, n1831, n1832, n1833, n1834, 
      n1835, n1836, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1852, n1854, n1855, n1856, n1857, n1858, 
      n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, 
      n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1879, n1880, 
      n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, 
      n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1899, n1900, n1901, 
      n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, 
      n1912, n1913, n1914, n1915, n1916, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1938, n1939, n1940, n1941, n1943, n1944, 
      n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, 
      n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, 
      n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
      n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, 
      n1985, n1987, n1988, n1990, n1991, n1992, n1993, n1995, n1996, n1999, 
      n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, 
      n2010, n2011, n2012, n2013, n2015, n2016, n2017, n2018, n2020, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2038, n2039, n2040, n2041, n2042, n2043, 
      n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, 
      n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2064, 
      n2066, n2067, n2068, n2069, n2070, n2071, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2104, n2105, n2106, n2107, n2108, 
      n2109, n2110, n2111, n2112, n2113, n2116, n2117, n2118, n2119, n2120, 
      n2121, n2122, n2124, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2183, 
      n2184, n2185, n2186, n2187, n2188, n2190, n2191, n2192, n2193, n2194, 
      n2195, n2196, n2198, n2199, n2202, n2203, n2204, n2206, n2207, n2208, 
      n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, 
      n2219, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, 
      n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2238, n2240, n2241, 
      n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2261, n2262, n2263, 
      n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, 
      n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, 
      n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
      n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, 
      n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, 
      n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, 
      n2324, n2325, n2326, n2327, n2328, n2330, n2331, n2332, n2333, n2334, 
      n2335, n2336, n2338, n2339, n2341, n2342, n2344, n2346, n2347, n2348, 
      n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, 
      n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, 
      n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, 
      n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
      n2389, n2390, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, 
      n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, 
      n2410, n2411, n2412, n2413, n2415, n2416, n2417, n2418, n2419, n2420, 
      n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
      n2431, n2432, n2433, n2435, n2436, n2437, n2438, n2440, n2441, n2442, 
      n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, 
      n2453, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, 
      n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, 
      n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, 
      n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
      n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, 
      n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, 
      n2515, n2516, n2517, n2518, n2520, n2521, n2522, n2523, n2524, n2526, 
      n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, 
      n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, 
      n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, 
      n2578, n2580, n2581, n2583, n2584, n2585, n2586, n2587, n2588, n2589, 
      n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2600, n2601, 
      n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2610, n2611, n2612, 
      n2613, n2614, n2615, n2616, n2617, n2618, n2620, n2621, n2622, n2623, 
      n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, 
      n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, 
      n2644, n2645, n2646, n2648, n2649, n2650, n2651, n2652, n2653, n2657, 
      n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, 
      n2668, n2669, n2670, n2671, n2673, n2674, n2675, n2677, n2679, n2680, 
      n2681, n2682, n2683, n2684, n2685, n2687, n2688, n2689, n2690, n2691, 
      n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2701, n2702, 
      n2703, n2704, n2706, n2708, n2709, n2710, n2711, n2713, n2714, n2715, 
      n2717, n2718, n2720, n2721, n2722, n2724, n2725, n2726, n2727, n2728, 
      n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, 
      n2740, n2741, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, 
      n2751, n2752, n2753, n2754, n2756, n2757, n2758, n2759, n2760, n2761, 
      n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, 
      n2772, n2773, n2774, n2775, n2778, n2779, n2780, n2781, n2782, n2783, 
      n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
      n2794, n2795, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, 
      n2805, n2806, n2807, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
      n2816, n2817, n2818, n2819, n2821, n2823, n2824, n2826, n2827, n2828, 
      n2829, n2830, n2831, n2833, n2834, n2835, n2836, n2837, n2838, n2839, 
      n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, 
      n2850, n2851, n2852, n2853, n2854, n2855, n2857, n2858, n2859, n2861, 
      n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, 
      n2872, n2873, n2874, n2875, n2876, n2878, n2879, n2880, n2881, n2882, 
      n2883, n2884, n2885, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
      n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, 
      n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
      n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, 
      n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, 
      n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, 
      n2944, n2945, n2946, n2947, n2948, n2949, n2951, n2952, n2953, n2955, 
      n2956, n2957, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
      n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2976, n2977, 
      n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, 
      n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, 
      n2998, n2999, n3000, n3002, n3003, n3004, n3005, n3006, n3007, n3008, 
      n3009, n3010, n3011, n3012, n3013, n3014, n3016, n3018, n3022, n3024, 
      n3025, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, 
      n3036, n3037, n3038, n3039, n3040, n3041, n3044, n3045, n3046, n3047, 
      n3048, n3049, n3050, n3052, n3053, n3054, n3055, n3056, n3057, n3058, 
      n3059, n3060, n3061, n3062, n3064, n3065, n3066, n3067, n3068, n3069, 
      n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, 
      n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, 
      n3090, n3091, n3093, n3094, n3095, n3096, n3097, n3098, n3100, n3101, 
      n3102, n3103, n3104, n3105, n3106, n3107, n3109, n3110, n3111, n3112, 
      n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
      n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3133, n3134, 
      n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, 
      n3145, n3146, n3147, n3148, n3149, n3150, n3152, n3153, n3155, n3156, 
      n3157, n3158, n3159, n3160, n3162, n3163, n3164, n3165, n3166, n3167, 
      n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, 
      n3178, n3179, n3180, n3181, n3182, n3183, n3185, n3186, n3187, n3188, 
      n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
      n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, 
      n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, 
      n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
      n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, 
      n3239, n3240, n3241, n3242, n3243, n3244, n3246, n3247, n3248, n3249, 
      n3250, n3251, n3252, n3253, n3255, n3256, n3257, n3258, n3259, n3260, 
      n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, 
      n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3280, n3281, n3282, 
      n3283, n3284, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, 
      n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, 
      n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, 
      n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3324, n3325, 
      n3326, n3327, n3328, n3329, n3330, n3331, n3333, n3334, n3335, n3336, 
      n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, 
      n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3356, n3357, n3358, 
      n3359, n3360, n3361, n3362, n3363, n3365, n3366, n3367, n3368, n3369, 
      n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, 
      n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, 
      n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3400, n3401, 
      n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, 
      n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, 
      n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, 
      n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3441, n3442, n3443, 
      n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, 
      n3454, n3455, n3456, n3457, n3458, n3460, n3461, n3462, n3463, n3464, 
      n3465, n3466, n3467, n3469, n3470, n3471, n3472, n3473, n3475, n3476, 
      n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
      n3487, n3488, n3489, n3491, n3492, n3493, n3494, n3495, n3496, n3497, 
      n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, 
      n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, 
      n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, 
      n3528, n3529, n3530, n3532, n3533, n3534, n3535, n3536, n3538, n3539, 
      n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, 
      n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, 
      n3561, n3562, n3563, n3564, n3565, n3567, n3568, n3569, n3570, n3571, 
      n3572, n3573, n3574, n3575, n3576, n3578, n3579, n3580, n3581, n3583, 
      n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3592, n3593, n3594, 
      n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, 
      n3605, n3606, n3607, n3608, n3611, n3612, n3613, n3614, n3615, n3616, 
      n3617, n3618, n3620, n3622, n3623, n3624, n3625, n3626, n3627, n3628, 
      n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, 
      n3639, n3640, n3641, n3642, n3643, n3645, n3646, n3647, n3648, n3650, 
      n3651, n3652, n3653, n3655, n3656, n3657, n3658, n3660, n3661, n3662, 
      n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, 
      n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, 
      n3684, n3685, n3686, n3688, n3689, n3690, n3691, n3693, n3694, n3695, 
      n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, 
      n3706, n3707, n3708, n3709, n3710, n3712, n3713, n3714, n3715, n3716, 
      n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, 
      n3727, n3728, n3729, n3730, n3732, n3733, n3734, n3735, n3736, n3737, 
      n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3746, n3747, n3748, 
      n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, 
      n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, 
      n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, 
      n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, 
      n3791, n3792, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, 
      n3802, n3804, n3805, n3807, n3808, n3809, n3810, n3811, n3812, n3813, 
      n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, 
      n3826, n3827, n3828, n3829, n3831, n3832, n3833, n3834, n3835, n3836, 
      n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3847, 
      n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, 
      n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, 
      n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, 
      n3878, n3879, n3880, n3881, n3884, n3885, n3886, n3887, n3888, n3889, 
      n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3898, n3899, n3900, 
      n3901, n3903, n3904, n3906, n3907, n3908, n3909, n3910, n3912, n3913, 
      n3914, n3916, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3926, 
      n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3937, 
      n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, 
      n3948, n3949, n3950, n3951, n3952, n3953, n3955, n3956, n3957, n3958, 
      n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, 
      n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, 
      n3979, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, 
      n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n4000, 
      n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, 
      n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, 
      n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, 
      n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, 
      n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4050, n4051, n4052, 
      n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
      n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, 
      n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, 
      n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, 
      n4105, n4106, n4107, n4108, n4109, n4110, n4112, n4113, n4114, n4115, 
      n4116, n4117, n4118, n4120, n4121, n4122, n4123, n4124, n4126, n4127, 
      n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, 
      n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, 
      n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, 
      n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, 
      n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, 
      n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, 
      n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, 
      n4218, n4219, n4221, n4222, n4224, n4225, n4226, n4227, n4229, n4230, 
      n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, 
      n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4249, n4250, n4251, 
      n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, 
      n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4272, 
      n4273, n4274, n4276, n4277, n4278, n4281, n4282, n4283, n4284, n4285, 
      n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, 
      n4296, n4297, n4298, n4299, n4300, n4302, n4303, n4304, n4305, n4306, 
      n4307, n4308, n4309, n4311, n4314, n4315, n4316, n4317, n4318, n4319, 
      n4320, n4321, n4322, n4323, n4324, n4326, n4327, n4328, n4330, n4331, 
      n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, 
      n4342, n4343, n4344, n4345, n4347, n4348, n4349, n4350, n4351, n4352, 
      n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
      n4363, n4364, n4365, n4366, n4369, n4370, n4371, n4372, n4373, n4374, 
      n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, 
      n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, 
      n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, 
      n4405, n4406, n4407, n4411, n4412, n4413, n4414, n4415, n4416, n4417, 
      n4418, n4419, n4420, n4421, n4422, n4424, n4425, n4426, n4427, n4428, 
      n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, 
      n4439, n4440, n4441, n4442, n4443, n4445, n4446, n4447, n4448, n4449, 
      n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, 
      n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, 
      n4470, n4471, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, 
      n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, 
      n4491, n4492, n4493, n4495, n4496, n4497, n4499, n4500, n4501, n4502, 
      n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, 
      n4513, n4514, n4515, n4516, n4517, n4520, n4521, n4522, n4523, n4524, 
      n4525, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4536, 
      n4537, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, 
      n4549, n4550, n4551, n4552, n4553, n4554, n4556, n4557, n4558, n4560, 
      n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, 
      n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, 
      n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, 
      n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4600, n4601, n4602, 
      n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, 
      n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4624, n4625, 
      n4626, n4627, n4628, n4630, n4631, n4632, n4633, n4634, n4635, n4636, 
      n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, 
      n4647, n4648, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, 
      n4658, n4659, n4660, n4661, n4663, n4664, n4665, n4666, n4667, n4668, 
      n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, 
      n4679, n4680, n4681, n4682, n4683, n4684, n4686, n4687, n4688, n4689, 
      n4691, n4692, n4694, n4696, n4697, n4698, n4699, n4700, n4701, n4702, 
      n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, 
      n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, 
      n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, 
      n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, 
      n4743, n4744, n4745, n4746, n4747, n4748, n4750, n4751, n4752, n4753, 
      n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, 
      n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, 
      n4774, n4775, n4777, n4778, n4779, n4780, n4781, n4782, n4784, n4785, 
      n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, 
      n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4806, n4807, 
      n4808, n4809, n4810, n4811, n4812, n4813, n4815, n4816, n4817, n4818, 
      n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, 
      n4829, n4830, n4832, n4833, n4834, n4835, n4837, n4838, n4839, n4840, 
      n4841, n4842, n4843, n4844, n4845, n4846, n4848, n4850, n4851, n4852, 
      n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, 
      n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4873, 
      n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, 
      n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, 
      n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, 
      n4904, n4906, n4907, n4908, n4909, n4910, n4912, n4913, n4914, n4915, 
      n4916, n4917, n4918, n4919, n4921, n4922, n4923, n4924, n4925, n4926, 
      n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4936, n4937, 
      n4938, n4939, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, 
      n4949, n4950, n4951, n4953, n4954, n4956, n4957, n4958, n4960, n4961, 
      n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, 
      n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, 
      n4982, n4983, n4984, n4985, n4986, n4989, n4990, n4991, n4992, n4993, 
      n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, 
      n5004, n5006, n5007, n5009, n5010, n5011, n5012, n5013, n5014, n5015, 
      n5017, n5018, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, 
      n5028, n5029, n5030, n5031, n5032, n5033, n5035, n5036, n5037, n5038, 
      n5039, n5040, n5041, n5042, n5043, n5044, n5046, n5047, n5048, n5049, 
      n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, 
      n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5068, n5070, n5071, 
      n5072, n5073, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, 
      n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, 
      n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, 
      n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, 
      n5113, n5114, n5115, n5116, n5117, n5119, n5120, n5121, n5123, n5124, 
      n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5134, n5135, 
      n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, 
      n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5155, n5156, 
      n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, 
      n5167, n5168, n5169, n5170, n5172, n5173, n5174, n5175, n5176, n5177, 
      n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, 
      n5188, n5189, n5190, n5191, n5192, n5193, n5196, n5197, n5198, n5199, 
      n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, 
      n5210, n5211, n5212, n5213, n5215, n5216, n5217, n5218, n5219, n5220, 
      n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5229, n5230, n5231, 
      n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, 
      n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, 
      n5252, n5253, n5254, n5255, n5256, n5258, n5259, n5260, n5261, n5262, 
      n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, 
      n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, 
      n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, 
      n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, 
      n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, 
      n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, 
      n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, 
      n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, 
      n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, 
      n5353, n5354, n5355, n5356, n5357, n5359, n5360, n5361, n5362, n5363, 
      n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, 
      n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, 
      n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, 
      n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5404, n5405, n5406, 
      n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, 
      n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5427, 
      n5428, n5429, n5432, n5433, n5434, n5436, n5437, n5439, n5440, n5441, 
      n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, 
      n5452, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, 
      n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, 
      n5473, n5474, n5475, n5476, n5477, n5478, n5480, n5481, n5482, n5483, 
      n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, 
      n5494, n5495, n5496, n5497, n5498, n5499, n5501, n5502, n5503, n5504, 
      n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, 
      n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, 
      n5526, n5527, n5528, n5529, n5530, n5531, n5533, n5534, n5535, n5536, 
      n5537, n5538, n5539, n5541, n5542, n5543, n5544, n5545, n5546, n5547, 
      n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, 
      n5558, n5559, n5560, n5561, n5563, n5564, n5565, n5566, n5568, n5569, 
      n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, 
      n5581, n5582, n5583, n5584, n5585, n5586, n5588, n5589, n5590, n5591, 
      n5593, n5594, n5595, n5596, n5598, n5599, n5600, n5601, n5602, n5603, 
      n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, 
      n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, 
      n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, 
      n5634, n5635, n5636, n5637, n5638, n5640, n5641, n5642, n5643, n5644, 
      n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, 
      n5655, n5656, n5658, n5659, n5660, n5662, n5663, n5664, n5665, n5666, 
      n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, 
      n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, 
      n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, 
      n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, 
      n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5719, 
      n5720, n5722, n5723, n5724, n5727, n5728, n5729, n5730, n5731, n5732, 
      n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, 
      n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, 
      n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, 
      n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, 
      n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, 
      n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, 
      n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, 
      n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, 
      n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, 
      n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, 
      n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, 
      n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, 
      n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, 
      n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, 
      n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, 
      n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, 
      n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, 
      n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, 
      n5913, n5914, n5915, n5916, n5917, n5918, n5920, n5921, n5922, n5923, 
      n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, 
      n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, 
      n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, 
      n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, 
      n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, 
      n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, 
      n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, 
      n5994, n5995, n5996, n5997, n5999, n6000, n6001, n6002, n6003, n6004, 
      n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, 
      n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, 
      n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, 
      n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, 
      n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, 
      n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, 
      n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, 
      n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, 
      n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, 
      n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, 
      n6106, n6107, n6108, n6109, n6110, n6112, n6113, n6114, n6115, n6116, 
      n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, 
      n6127, n6128, n6129, n6130, n6131, n6133, n6134, n6135, n6136, n6137, 
      n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, 
      n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6156, n6157, n6158, 
      n6159, n6160, n6161, n6162, n6164, n6165, n6166, n6167, n6168, n6169, 
      n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, 
      n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, 
      n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, 
      n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6211, 
      n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, 
      n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, 
      n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, 
      n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, 
      n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, 
      n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, 
      n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, 
      n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, 
      n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, 
      n6302, n6303, n6304, n6305, n6307, n6308, n6309, n6310, n6311, n6312, 
      n6313, n6314, n6315, n6316, n6317, n6319, n6321, n6322, n6323, n6324, 
      n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, 
      n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, 
      n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6353, n6354, n6355, 
      n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, 
      n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, 
      n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, 
      n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, 
      n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, 
      n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, 
      n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6425, n6426, n6427, 
      n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6436, n6437, n6438, 
      n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, 
      n6449, n6450, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, 
      n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, 
      n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, 
      n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, 
      n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, 
      n6500, n6501, n6502, n6503, n6504, n6506, n6507, n6508, n6509, n6510, 
      n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, 
      n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, 
      n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, 
      n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, 
      n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, 
      n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, 
      n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, 
      n6583, n6584, n6585, n6586, n6587, n6588, n6590, n6591, n6592, n6593, 
      n6594, n6595, n6596, n6597, n6598, n6600, n6601, n6602, n6603, n6604, 
      n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, 
      n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, 
      n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6636, 
      n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, 
      n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, 
      n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, 
      n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, 
      n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, 
      n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, 
      n6698, n6699, n6700, n6701, n6702, n6703, n6705, n6706, n6707, n6708, 
      n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, 
      n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, 
      n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, 
      n6739, n6740, n6742, n6743, n6744, n6746, n6747, n6748, n6749, n6750, 
      n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, 
      n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, 
      n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, 
      n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, 
      n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, 
      n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, 
      n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, 
      n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, 
      n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, 
      n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, 
      n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, 
      n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, 
      n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, 
      n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, 
      n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, 
      n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, 
      n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, 
      n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, 
      n6931, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, 
      n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, 
      n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, 
      n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, 
      n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, 
      n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, 
      n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, 
      n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, 
      n7013, n7014, n7015, n7016, n7018, n7019, n7021, n7022, n7023, n7024, 
      n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, 
      n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, 
      n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, 
      n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, 
      n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, 
      n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, 
      n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, 
      n7095, n7097, n7098, n7099, n7100, n7101, n7103, n7104, n7105, n7106, 
      n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, 
      n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, 
      n7127, n7128, n7129, n7130, n7132, n7133, n7135, n7137, n7138, n7139, 
      n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, 
      n7150, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, 
      n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, 
      n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, 
      n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, 
      n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, 
      n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, 
      n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, 
      n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, 
      n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, 
      n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, 
      n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, 
      n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, 
      n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, 
      n7282, n7283, n7284, n7286, n7287, n7288, n7289, n7290, n7291, n7292, 
      n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, 
      n7303, n7304, n7305, n7306, n7307, n7308, n7310, n7311, n7312, n7313, 
      n7314, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, 
      n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, 
      n7337, n7338, n7339, n7340, n7341, n7343, n7344, n7345, n7346, n7347, 
      n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, 
      n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, 
      n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, 
      n7378, n7379, n7380, n7382, n7383, n7384, n7385, n7386, n7387, n7388, 
      n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, 
      n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, 
      n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, 
      n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, 
      n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, 
      n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, 
      n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, 
      n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, 
      n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, 
      n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, 
      n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, 
      n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7508, n7509, 
      n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, 
      n7520, n7521, n7522, n7524, n7525, n7526, n7527, n7528, n7530, n7531, 
      n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, 
      n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, 
      n7552, n7553, n7554, n7556, n7558, n7559, n7560, n7561, n7562, n7563, 
      n7564, n7565, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, 
      n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, 
      n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, 
      n7595, n7596, n7597, n7598, n7599, n7600, n7602, n7603, n7604, n7605, 
      n7606, n7607, n7608, n7609, n7611, n7612, n7613, n7614, n7615, n7616, 
      n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, 
      n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, 
      n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, 
      n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, 
      n7657, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, 
      n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, 
      n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, 
      n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, 
      n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, 
      n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, 
      n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7727, n7728, 
      n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, 
      n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, 
      n7749, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, 
      n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, 
      n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, 
      n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, 
      n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, 
      n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, 
      n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, 
      n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, 
      n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, 
      n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, 
      n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, 
      n7860, n7861, n7862, n7863, n7864, n7865, n7867, n7868, n7869, n7870, 
      n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7881, 
      n7882, n7883, n7884, n7885, n7887, n7888, n7889, n7890, n7891, n7892, 
      n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7902, n7903, 
      n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, 
      n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, 
      n7924, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, 
      n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, 
      n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, 
      n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, 
      n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, 
      n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, 
      n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, 
      n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, 
      n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, 
      n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, 
      n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8034, n8035, 
      n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, 
      n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, 
      n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, 
      n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, 
      n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, 
      n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, 
      n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, 
      n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, 
      n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, 
      n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, 
      n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, 
      n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, 
      n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, 
      n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, 
      n8176, n8177, n8178, n8179, n8180, n8181, n8183, n8184, n8185, n8186, 
      n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, 
      n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, 
      n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, 
      n8219, n8220, n8221, n8222, n8223, n8225, n8226, n8227, n8228, n8229, 
      n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, 
      n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, 
      n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, 
      n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, 
      n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, 
      n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, 
      n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, 
      n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, 
      n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, 
      n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, 
      n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, 
      n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, 
      n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, 
      n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, 
      n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, 
      n8380, n8381, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, 
      n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, 
      n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, 
      n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, 
      n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, 
      n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, 
      n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, 
      n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, 
      n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, 
      n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, 
      n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, 
      n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, 
      n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, 
      n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, 
      n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, 
      n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, 
      n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, 
      n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, 
      n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, 
      n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, 
      n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, 
      n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, 
      n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, 
      n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, 
      n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, 
      n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, 
      n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, 
      n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, 
      n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, 
      n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8682, 
      n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, 
      n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, 
      n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, 
      n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, 
      n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, 
      n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, 
      n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, 
      n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, 
      n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, 
      n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, 
      n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, 
      n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, 
      n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, 
      n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, 
      n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, 
      n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8841, n8842, n8843, 
      n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, 
      n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, 
      n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, 
      n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, 
      n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, 
      n8894, n8895, n8896, n8897, n8898, n8899, n8901, n8902, n8903, n8904, 
      n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, 
      n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, 
      n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, 
      n8935, n8936, n8937, n8939, n8940, n8941, n8942, n8943, n8944, n8945, 
      n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, 
      n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, 
      n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, 
      n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, 
      n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, 
      n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, 
      n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, 
      n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, 
      n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, 
      n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, 
      n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, 
      n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, 
      n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, 
      n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, 
      n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, 
      n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, 
      n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, 
      n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, 
      n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, 
      n9136, n9137, n9138, n9139, n9140, n9141, n9143, n9144, n9145, n9146, 
      n9147, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, 
      n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, 
      n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, 
      n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, 
      n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, 
      n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9208, n9209, 
      n9210, n9211, n9212, n9213, n9215, n9216, n9217, n9218, n9219, n9220, 
      n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, 
      n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, 
      n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, 
      n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, 
      n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, 
      n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, 
      n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, 
      n9291, n9293, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, 
      n9303, n9304, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, 
      n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, 
      n9325, n9326, n9327, n9328, n9329, n9332, n9333, n9334, n9335, n9336, 
      n9337, n9338, n9339, n9340, n9342, n9343, n9345, n9346, n9348, n9349, 
      n9350, n9351, n9354, n9355, n9357, n9358, n9359, n9360, n9361, n9362, 
      n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, 
      n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, 
      n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, 
      n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, 
      n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, 
      n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, 
      n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, 
      n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, 
      n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, 
      n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, 
      n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9473, n9474, 
      n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, 
      n9485, n9486, n9487, n9488, n9490, n9491, n9493, n9494, n9495, n9496, 
      n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, 
      n9507, n9508, n9509, n9512, n9514, n9515, n9516, n9517, n9518, n9519, 
      n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, 
      n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, 
      n9540, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, 
      n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, 
      n9561, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, 
      n9572, n9573, n9574, n9575, n9577, n9578, n9579, n9580, n9581, n9582, 
      n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, 
      n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, 
      n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, 
      n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, 
      n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9633, 
      n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, 
      n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, 
      n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9663, n9664, 
      n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, 
      n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, 
      n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, 
      n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, 
      n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, 
      n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, 
      n9725, n9726, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, 
      n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, 
      n9746, n9747, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, 
      n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, 
      n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, 
      n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, 
      n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, 
      n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, 
      n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, 
      n9817, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, 
      n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, 
      n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, 
      n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, 
      n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, 
      n9868, n9869, n9870, n9871, n9872, n9874, n9875, n9876, n9877, n9878, 
      n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, 
      n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, 
      n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, 
      n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, 
      n9920, n9921, n9922, n9924, n9925, n9926, n9927, n9928, n9929, n9930, 
      n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, 
      n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, 
      n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, 
      n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, 
      n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, 
      n9982, n9984, n9985, n9986, n9989, n9990, n9991, n9992, n9993, n9994, 
      n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, 
      n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, 
      n10014, n10015, n10016, n10018, n10019, n10020, n10021, n10022, n10023, 
      n10024, n10025, n10026, n10027, n10028, n10029, n10031, n10032, n10033, 
      n10034, n10035, n10037, n10038, n10039, n10040, n10041, n10042, n10043, 
      n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, 
      n10053, n10054, n10055, n10056, n10058, n10059, n10060, n10061, n10062, 
      n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, 
      n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, 
      n10081, n10082, n10084, n10085, n10086, n10087, n10088, n10089, n10090, 
      n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, 
      n10100, n10101, n10103, n10104, n10106, n10107, n10108, n10109, n10110, 
      n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, 
      n10120, n10122, n10124, n10125, n10126, n10127, n10128, n10129, n10130, 
      n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, 
      n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, 
      n10149, n10151, n10152, n10154, n10156, n10157, n10158, n10159, n10160, 
      n10161, n10162, n10163, n10164, n10165, n10166, n10168, n10169, n10170, 
      n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, 
      n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, 
      n10190, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, 
      n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, 
      n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, 
      n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, 
      n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, 
      n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, 
      n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, 
      n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, 
      n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, 
      n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, 
      n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, 
      n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, 
      n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, 
      n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, 
      n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, 
      n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, 
      n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, 
      n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, 
      n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, 
      n10362, n10363, n10364, n10365, n10366, n10368, n10369, n10370, n10371, 
      n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, 
      n10381, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, 
      n10391, n10392, n10394, n10395, n10396, n10397, n10398, n10399, n10400, 
      n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, 
      n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, 
      n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, 
      n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, 
      n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, 
      n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, 
      n10455, n10456, n10457, n10458, n10459, n10460, n10462, n10463, n10464, 
      n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, 
      n10474, n10475, n10476, n10477, n10479, n10480, n10481, n10482, n10483, 
      n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10493, 
      n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, 
      n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, 
      n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, 
      n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, 
      n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10538, n10539, 
      n10540, n10541, n10544, n10545, n10546, n10547, n10548, n10549, n10550, 
      n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, 
      n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, 
      n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, 
      n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, 
      n10587, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, 
      n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, 
      n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, 
      n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, 
      n10624, n10625, n10627, n10628, n10629, n10630, n10632, n10633, n10635, 
      n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, 
      n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, 
      n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, 
      n10663, n10664, n10665, n10666, n10667, n10669, n10670, n10671, n10672, 
      n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, 
      n10682, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, 
      n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, 
      n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, 
      n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, 
      n10719, n10720, n10721, n10722, n10723, n10725, n10726, n10727, n10728, 
      n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, 
      n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, 
      n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, 
      n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, 
      n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, 
      n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, 
      n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10792, 
      n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, 
      n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, 
      n10811, n10812, n10814, n10815, n10816, n10817, n10818, n10819, n10820, 
      n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, 
      n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, 
      n10839, n10840, n10841, n10842, n10843, n10845, n10846, n10847, n10848, 
      n10849, n10850, n10851, n10852, n10854, n10855, n10856, n10857, n10858, 
      n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, 
      n10868, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, 
      n10878, n10879, n10880, n10882, n10883, n10884, n10885, n10886, n10887, 
      n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, 
      n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, 
      n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10914, n10915, 
      n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, 
      n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, 
      n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, 
      n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, 
      n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, 
      n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, 
      n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, 
      n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, 
      n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10996, n10997, 
      n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, 
      n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, 
      n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, 
      n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, 
      n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, 
      n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, 
      n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, 
      n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, 
      n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, 
      n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, 
      n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, 
      n11097, n11098, n11099, n11100, n11101, n11103, n11104, n11106, n11107, 
      n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, 
      n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, 
      n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, 
      n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, 
      n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, 
      n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, 
      n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, 
      n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, 
      n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, 
      n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, 
      n11199, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, 
      n11209, n11210, n11211, n11212, n11214, n11215, n11216, n11217, n11218, 
      n11219, n11220, n11221, n11222, n11224, n11225, n11226, n11227, n11228, 
      n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, 
      n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, 
      n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, 
      n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, 
      n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, 
      n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, 
      n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11291, n11292, 
      n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, 
      n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, 
      n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, 
      n11320, n11321, n11322, n11324, n11326, n11327, n11328, n11329, n11330, 
      n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, 
      n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, 
      n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, 
      n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, 
      n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, 
      n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, 
      n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, 
      n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, 
      n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, 
      n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, 
      n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, 
      n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, 
      n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, 
      n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, 
      n11457, n11458, n11459, n11460, n11461, n11463, n11464, n11465, n11466, 
      n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, 
      n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, 
      n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, 
      n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, 
      n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, 
      n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, 
      n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, 
      n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, 
      n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, 
      n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, 
      n11557, n11558, n11559, n11560, n11561, n11563, n11564, n11565, n11566, 
      n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11575, n11576, 
      n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, 
      n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, 
      n11595, n11596, n11597, n11598, n11600, n11601, n11602, n11603, n11604, 
      n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, 
      n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, 
      n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, 
      n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, 
      n11641, n11642, n11643, n11644, n11646, n11647, n11648, n11649, n11650, 
      n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, 
      n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, 
      n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, 
      n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, 
      n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, 
      n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, 
      n11705, n11706, n11707, n11708, n11709, n11711, n11712, n11713, n11714, 
      n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, 
      n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11733, 
      n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, 
      n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, 
      n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, 
      n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, 
      n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, 
      n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, 
      n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, 
      n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, 
      n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, 
      n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, 
      n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, 
      n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, 
      n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, 
      n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, 
      n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, 
      n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, 
      n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, 
      n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, 
      n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, 
      n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, 
      n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, 
      n11924, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, 
      n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, 
      n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, 
      n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, 
      n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, 
      n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, 
      n11979, n11980, n11981, n11983, n11984, n11985, n11986, n11987, n11988, 
      n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, 
      n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, 
      n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, 
      n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, 
      n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, 
      n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, 
      n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, 
      n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, 
      n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, 
      n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, 
      n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, 
      n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, 
      n12097, n12098, n12099, n12100, n12101, n12102, n12104, n12105, n12106, 
      n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, 
      n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, 
      n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, 
      n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, 
      n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, 
      n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, 
      n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, 
      n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, 
      n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, 
      n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, 
      n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, 
      n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, 
      n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, 
      n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, 
      n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, 
      n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12251, 
      n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, 
      n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, 
      n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, 
      n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, 
      n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, 
      n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, 
      n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, 
      n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, 
      n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, 
      n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, 
      n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, 
      n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, 
      n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, 
      n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, 
      n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, 
      n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, 
      n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, 
      n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, 
      n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, 
      n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, 
      n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, 
      n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, 
      n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, 
      n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, 
      n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, 
      n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, 
      n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, 
      n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, 
      n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12513, n12514, 
      n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, 
      n12526, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, 
      n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, 
      n12546, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, 
      n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12566, 
      n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, 
      n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, 
      n12585, n12586, n12587, n12588, n12589, n12590, n12592, n12593, n12594, 
      n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, 
      n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, 
      n12614, n12615, n12616, n12617, n12619, n12620, n12621, n12622, n12624, 
      n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, 
      n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, 
      n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, 
      n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, 
      n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, 
      n12670, n12671, n12672, n12673, n12674, n12676, n12677, n12678, n12679, 
      n12680, n12681, n12682, n12683, n12684, n12685, n12687, n12688, n12689, 
      n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, 
      n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12707, n12708, 
      n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, 
      n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, 
      n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12736, n12737, 
      n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, 
      n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, 
      n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, 
      n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, 
      n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, 
      n12783, n12784, n12785, n12786, n12787, n12789, n12790, n12791, n12792, 
      n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, 
      n12802, n12803, n12804, n12805, n12807, n12808, n12809, n12810, n12811, 
      n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, 
      n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, 
      n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, 
      n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, 
      n12848, n12849, n12850, n12852, n12853, n12854, n12856, n12857, n12858, 
      n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, 
      n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, 
      n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, 
      n12887, n12888, n12890, n12891, n12892, n12893, n12894, n12895, n12896, 
      n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, 
      n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, 
      n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, 
      n12924, n12925, n12926, n12928, n12929, n12930, n12931, n12932, n12933, 
      n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, 
      n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, 
      n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, 
      n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, 
      n12970, n12971, n12973, n12974, n12975, n12976, n12977, n12979, n12980, 
      n12981, n12982, n12983, n12984, n12986, n12987, n12988, n12991, n12993, 
      n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, 
      n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, 
      n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, 
      n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, 
      n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, 
      n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, 
      n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, 
      n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, 
      n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, 
      n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, 
      n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, 
      n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, 
      n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, 
      n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, 
      n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, 
      n13131, n13132, n13133, n13134, n13136, n13137, n13138, n13139, n13140, 
      n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, 
      n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, 
      n13159, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, 
      n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, 
      n13178, n13179, n13180, n13181, n13182, n13183, n13185, n13186, n13187, 
      n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, 
      n13197, n13198, n13199, n13200, n13202, n13204, n13205, n13206, n13207, 
      n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, 
      n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, 
      n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, 
      n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, 
      n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, 
      n13254, n13255, n13257, n13258, n13259, n13260, n13261, n13262, n13263, 
      n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, 
      n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, 
      n13282, n13283, n13284, n13286, n13287, n13288, n13289, n13291, n13292, 
      n13294, n13295, n13296, n13297, n13298, n13300, n13301, n13302, n13303, 
      n13304, n13305, n13306, n13307, n13309, n13310, n13311, n13312, n13313, 
      n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, 
      n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, 
      n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13341, 
      n13342, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, 
      n13352, n13353, n13354, n13356, n13357, n13358, n13359, n13360, n13361, 
      n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, 
      n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, 
      n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, 
      n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13399, 
      n13400, n13401, n13402, n13403, n13404, n13405, n13407, n13408, n13409, 
      n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, 
      n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, 
      n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13436, n13437, 
      n13438, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13449, 
      n13450, n13453, n13454, n13457, n13458, n13459, n13460, n13462, n13463, 
      n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, 
      n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, 
      n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, 
      n13491, n13492, n13494, n13495, n13496, n13497, n13498, n13499, n13500, 
      n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, 
      n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13518, n13519, 
      n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, 
      n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, 
      n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, 
      n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, 
      n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, 
      n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, 
      n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, 
      n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, 
      n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, 
      n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, 
      n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13619, 
      n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, 
      n13629, n13630, n13631, n13633, n13634, n13635, n13636, n13638, n13639, 
      n13640, n13641, n13642, n13643, n13644, n13646, n13647, n13648, n13649, 
      n13650, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, 
      n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, 
      n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, 
      n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, 
      n13687, n13688, n13690, n13691, n13692, n13693, n13695, n13696, n13697, 
      n13698, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, 
      n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, 
      n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, 
      n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, 
      n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, 
      n13745, n13746, n13747, n13748, n13749, n13751, n13752, n13753, n13754, 
      n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, 
      n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, 
      n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, 
      n13782, n13783, n13784, n13785, n13787, n13788, n13789, n13790, n13791, 
      n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, 
      n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, 
      n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, 
      n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, 
      n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, 
      n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, 
      n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, 
      n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, 
      n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, 
      n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, 
      n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, 
      n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, 
      n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13909, 
      n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, 
      n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, 
      n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, 
      n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, 
      n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, 
      n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, 
      n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, 
      n13973, n13974, n13975, n13977, n13978, n13980, n13981, n13982, n13983, 
      n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, 
      n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, 
      n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, 
      n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, 
      n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, 
      n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, 
      n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, 
      n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14056, 
      n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, 
      n14066, n14067, n14068, n14069, n14070, n14072, n14073, n14074, n14075, 
      n14076, n14077, n14078, n14079, n14080, n14082, n14083, n14084, n14085, 
      n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, 
      n14095, n14097, n14099, n14100, n14101, n14102, n14103, n14104, n14105, 
      n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, 
      n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, 
      n14124, n14125, n14126, n14127, n14129, n14130, n14131, n14132, n14133, 
      n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, 
      n14143, n14144, n14146, n14147, n14148, n14149, n14150, n14151, n14152, 
      n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, 
      n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, 
      n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, 
      n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14188, n14189, 
      n14190, n14191, n14192, n14194, n14196, n14197, n14198, n14199, n14200, 
      n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, 
      n14210, n14211, n14213, n14214, n14215, n14216, n14217, n14218, n14219, 
      n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, 
      n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14238, 
      n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, 
      n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, 
      n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, 
      n14266, n14267, n14268, n14269, n14270, n14271, n14273, n14274, n14276, 
      n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, 
      n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, 
      n14295, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, 
      n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, 
      n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, 
      n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, 
      n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, 
      n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, 
      n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, 
      n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, 
      n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, 
      n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, 
      n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, 
      n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, 
      n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, 
      n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, 
      n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, 
      n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, 
      n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, 
      n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, 
      n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, 
      n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, 
      n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, 
      n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, 
      n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, 
      n14503, n14504, n14505, n14507, n14508, n14509, n14510, n14511, n14512, 
      n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, 
      n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, 
      n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, 
      n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, 
      n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, 
      n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, 
      n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, 
      n14576, n14577, n14579, n14580, n14581, n14582, n14583, n14584, n14585, 
      n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, 
      n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, 
      n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, 
      n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, 
      n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, 
      n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, 
      n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, 
      n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, 
      n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, 
      n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, 
      n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, 
      n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, 
      n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, 
      n14703, n14704, n14705, n14706, n14707, n14708, n14710, n14711, n14712, 
      n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, 
      n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, 
      n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, 
      n14740, n14741, n14742, n14744, n14745, n14747, n14748, n14749, n14750, 
      n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, 
      n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, 
      n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, 
      n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14786, n14787, 
      n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, 
      n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, 
      n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, 
      n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, 
      n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, 
      n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, 
      n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, 
      n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, 
      n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, 
      n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, 
      n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, 
      n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, 
      n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, 
      n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, 
      n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, 
      n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, 
      n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, 
      n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, 
      n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, 
      n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, 
      n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, 
      n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, 
      n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, 
      n14995, n14996, n14997, n14998, n14999, n15000, n15002, n15003, n15004, 
      n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, 
      n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, 
      n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, 
      n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, 
      n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, 
      n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, 
      n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, 
      n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15078, n15079, 
      n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, 
      n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, 
      n15098, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, 
      n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, 
      n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, 
      n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, 
      n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15143, n15144, 
      n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, 
      n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, 
      n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, 
      n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, 
      n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, 
      n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, 
      n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, 
      n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, 
      n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, 
      n15226, n15227, n15228, n15229, n15230, n15232, n15233, n15234, n15235, 
      n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, 
      n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, 
      n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, 
      n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, 
      n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, 
      n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, 
      n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, 
      n15301, n15302, n15303, n15305, n15306, n15307, n15308, n15309, n15310, 
      n15311, n15312, n15313, n15314, n15316, n15317, n15318, n15319, n15321, 
      n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, 
      n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, 
      n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, 
      n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15358, 
      n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, 
      n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, 
      n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, 
      n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, 
      n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15404, 
      n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, 
      n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, 
      n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, 
      n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, 
      n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, 
      n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, 
      n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, 
      n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, 
      n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, 
      n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, 
      n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, 
      n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, 
      n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, 
      n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, 
      n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, 
      n15542, n15543, n15544, n15545, n15546, n15548, n15549, n15550, n15551, 
      n15552, n15553, n15554, n15555, n15556, n15557, n15559, n15560, n15562, 
      n15563, n15564, n15565, n15566, n15568, n15569, n15570, n15571, n15572, 
      n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, 
      n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, 
      n15591, n15592, n15594, n15595, n15596, n15597, n15598, n15599, n15600, 
      n15601, n15602, n15604, n15605, n15606, n15608, n15609, n15610, n15611, 
      n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, 
      n15621, n15622, n15623, n15625, n15626, n15627, n15628, n15629, n15631, 
      n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, 
      n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, 
      n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, 
      n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, 
      n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, 
      n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, 
      n15686, n15687, n15688, n15689, n15690, n15691, n15693, n15694, n15695, 
      n15696, n15697, n15698, n15699, n15700, n15701, n15703, n15704, n15705, 
      n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, 
      n15715, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, 
      n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, 
      n15734, n15735, n15736, n15737, n15739, n15740, n15741, n15742, n15744, 
      n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, 
      n15755, n15757, n15758, n15759, n15760, n15761, n15762, n15764, n15765, 
      n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, 
      n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15785, 
      n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, 
      n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, 
      n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, 
      n15813, n15814, n15815, n15817, n15818, n15819, n15820, n15821, n15822, 
      n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, 
      n15832, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, 
      n15842, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, 
      n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, 
      n15861, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, 
      n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, 
      n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15890, 
      n15891, n15892, n15893, n15894, n15896, n15897, n15898, n15899, n15900, 
      n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, 
      n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, 
      n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, 
      n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, 
      n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, 
      n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, 
      n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, 
      n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, 
      n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, 
      n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, 
      n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, 
      n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, 
      n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, 
      n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, 
      n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, 
      n16036, n16037, n16038, n16041, n16042, n16043, n16045, n16046, n16048, 
      n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, 
      n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, 
      n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, 
      n16076, n16077, n16078, n16080, n16082, n16083, n16084, n16085, n16086, 
      n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, 
      n16096, n16097, n16098, n16100, n16101, n16102, n16103, n16104, n16105, 
      n16106, n16107, n16108, n16109, n16112, n16113, n16114, n16115, n16116, 
      n16117, n16118, n16120, n16121, n16122, n16123, n16124, n16125, n16126, 
      n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, 
      n16136, n16137, n16138, n16140, n16141, n16142, n16143, n16144, n16145, 
      n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16154, n16155, 
      n16156, n16157, n16158, n16159, n16161, n16162, n16163, n16164, n16165, 
      n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, 
      n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, 
      n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, 
      n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, 
      n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, 
      n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, 
      n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, 
      n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, 
      n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, 
      n16247, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, 
      n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, 
      n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16276, n16277, 
      n16278, n16280, n16281, n16283, n16284, n16285, n16286, n16287, n16288, 
      n16290, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, 
      n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, 
      n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, 
      n16319, n16320, n16321, n16322, n16323, n16324, n16326, n16327, n16328, 
      n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, 
      n16339, n16340, n16341, n16342, n16344, n16345, n16346, n16347, n16348, 
      n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, 
      n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, 
      n16368, n16369, n16370, n16371, n16372, n16374, n16375, n16376, n16377, 
      n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, 
      n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, 
      n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, 
      n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, 
      n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, 
      n16423, n16424, n16426, n16427, n16428, n16429, n16430, n16431, n16432, 
      n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, 
      n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, 
      n16451, n16452, n16453, n16455, n16456, n16457, n16458, n16459, n16460, 
      n16461, n16462, n16464, n16465, n16466, n16467, n16468, n16469, n16470, 
      n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, 
      n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, 
      n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, 
      n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, 
      n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, 
      n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, 
      n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, 
      n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, 
      n16544, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, 
      n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, 
      n16563, n16564, n16565, n16566, n16568, n16569, n16570, n16571, n16572, 
      n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, 
      n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, 
      n16591, n16593, n16595, n16597, n16598, n16599, n16600, n16601, n16602, 
      n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, 
      n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, 
      n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, 
      n16630, n16631, n16632, n16634, n16635, n16636, n16637, n16638, n16639, 
      n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, 
      n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, 
      n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, 
      n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, 
      n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, 
      n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16693, n16694, 
      n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, 
      n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16712, n16713, 
      n16714, n16715, n16716, n16717, n16719, n16720, n16721, n16722, n16723, 
      n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, 
      n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, 
      n16742, n16743, n16744, n16745, n16746, n16747, n16749, n16750, n16751, 
      n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, 
      n16761, n16762, n16764, n16765, n16766, n16767, n16768, n16769, n16770, 
      n16771, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, 
      n16782, n16783, n16784, n16785, n16786, n16787, n16789, n16790, n16792, 
      n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, 
      n16802, n16803, n16804, n16806, n16807, n16808, n16809, n16810, n16811, 
      n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, 
      n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, 
      n16831, n16832, n16833, n16834, n16836, n16837, n16838, n16839, n16840, 
      n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, 
      n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, 
      n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, 
      n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, 
      n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, 
      n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, 
      n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, 
      n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, 
      n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, 
      n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, 
      n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, 
      n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, 
      n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, 
      n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, 
      n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, 
      n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, 
      n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, 
      n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, 
      n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, 
      n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, 
      n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, 
      n17032, n17033, n17034, n17035, n17036, n17037, n17039, n17040, n17041, 
      n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, 
      n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, 
      n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, 
      n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, 
      n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, 
      n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, 
      n17096, n17097, n17098, n17099, n17100, n17104, n17105, n17106, n17107, 
      n17108, n17109, n17110, n17112, n17113, n17114, n17115, n17116, n17117, 
      n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, 
      n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, 
      n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, 
      n17145, n17146, n17148, n17150, n17151, n17152, n17153, n17154, n17156, 
      n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, 
      n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, 
      n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, 
      n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, 
      n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, 
      n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, 
      n17211, n17212, n17214, n17215, n17216, n17217, n17218, n17219, n17220, 
      n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17229, n17230, 
      n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, 
      n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, 
      n17249, n17250, n17252, n17253, n17254, n17255, n17256, n17257, n17258, 
      n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, 
      n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, 
      n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, 
      n17286, n17287, n17288, n17289, n17291, n17293, n17294, n17295, n17296, 
      n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, 
      n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, 
      n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, 
      n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, 
      n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, 
      n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, 
      n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, 
      n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, 
      n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, 
      n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, 
      n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, 
      n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, 
      n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, 
      n17414, n17415, n17416, n17418, n17419, n17420, n17421, n17422, n17423, 
      n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, 
      n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17441, n17442, 
      n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, 
      n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, 
      n17463, n17464, n17465, n17467, n17468, n17469, n17470, n17471, n17472, 
      n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, 
      n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, 
      n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, 
      n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, 
      n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, 
      n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, 
      n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, 
      n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, 
      n17545, n17546, n17547, n17548, n17549, n17551, n17552, n17553, n17554, 
      n17555, n17556, n17558, n17559, n17560, n17561, n17562, n17563, n17564, 
      n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, 
      n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, 
      n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, 
      n17592, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, 
      n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, 
      n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, 
      n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, 
      n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, 
      n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, 
      n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, 
      n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, 
      n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, 
      n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17683, 
      n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, 
      n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, 
      n17702, n17703, n17705, n17706, n17708, n17709, n17710, n17711, n17712, 
      n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, 
      n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, 
      n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, 
      n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, 
      n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, 
      n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, 
      n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, 
      n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, 
      n17786, n17787, n17788, n17791, n17792, n17793, n17794, n17795, n17796, 
      n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, 
      n17806, n17807, n17808, n17810, n17811, n17812, n17813, n17814, n17815, 
      n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, 
      n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, 
      n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, 
      n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, 
      n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, 
      n17861, n17862, n17863, n17864, n17865, n17866, n17868, n17869, n17870, 
      n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, 
      n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, 
      n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, 
      n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, 
      n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, 
      n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, 
      n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, 
      n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, 
      n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, 
      n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, 
      n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, 
      n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, 
      n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, 
      n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, 
      n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, 
      n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, 
      n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, 
      n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, 
      n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, 
      n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, 
      n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, 
      n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, 
      n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, 
      n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, 
      n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, 
      n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, 
      n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18116, n18118, 
      n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, 
      n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, 
      n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, 
      n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, 
      n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, 
      n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, 
      n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, 
      n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, 
      n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, 
      n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, 
      n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, 
      n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, 
      n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, 
      n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, 
      n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, 
      n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, 
      n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, 
      n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, 
      n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, 
      n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, 
      n18299, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, 
      n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, 
      n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, 
      n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, 
      n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, 
      n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, 
      n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, 
      n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, 
      n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, 
      n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, 
      n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, 
      n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18407, n18408, 
      n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, 
      n18418, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, 
      n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, 
      n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, 
      n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, 
      n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, 
      n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, 
      n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, 
      n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, 
      n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, 
      n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, 
      n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, 
      n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, 
      n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, 
      n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, 
      n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18555, 
      n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, 
      n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, 
      n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, 
      n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, 
      n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, 
      n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, 
      n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, 
      n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, 
      n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, 
      n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, 
      n18646, n18647, n18648, n18649, n18650, n18651, n18653, n18654, n18655, 
      n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, 
      n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18674, 
      n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, 
      n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, 
      n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, 
      n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, 
      n18711, n18712, n18714, n18716, n18717, n18718, n18719, n18720, n18721, 
      n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, 
      n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, 
      n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, 
      n18749, n18750, n18751, n18752, n18753, n18754, n18756, n18757, n18758, 
      n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, 
      n18768, n18769, n18770, n18772, n18773, n18774, n18775, n18776, n18777, 
      n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, 
      n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, 
      n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, 
      n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, 
      n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, 
      n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, 
      n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, 
      n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, 
      n18850, n18851, n18853, n18854, n18855, n18856, n18857, n18858, n18859, 
      n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18869, 
      n18870, n18871, n18872, n18873, n18874, n18876, n18877, n18879, n18880, 
      n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18889, n18890, 
      n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, 
      n18900, n18901, n18902, n18903, n18904, n18905, n18907, n18908, n18909, 
      n18911, n18912, n18913, n18914, n18916, n18917, n18918, n18919, n18921, 
      n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, 
      n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18940, 
      n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, 
      n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, 
      n18959, n18960, n18961, n18962, n18963, n18964, n18966, n18967, n18968, 
      n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, 
      n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, 
      n18987, n18988, n18990, n18991, n18992, n18993, n18994, n18995, n18996, 
      n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, 
      n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, 
      n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, 
      n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, 
      n19035, n19036, n19037, n19039, n19040, n19041, n19042, n19043, n19044, 
      n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, 
      n19054, n19056, n19057, n19059, n19060, n19061, n19062, n19064, n19065, 
      n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, 
      n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, 
      n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, 
      n19093, n19094, n19095, n19096, n19097, n19098, n19100, n19101, n19102, 
      n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, 
      n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, 
      n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, 
      n19130, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, 
      n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19148, n19149, 
      n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, 
      n19159, n19160, n19161, n19162, n19163, n19164, n19166, n19167, n19168, 
      n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, 
      n19178, n19179, n19180, n19181, n19183, n19184, n19185, n19186, n19187, 
      n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, 
      n19197, n19198, n19199, n19200, n19201, n19202, n19204, n19205, n19206, 
      n19207, n19208, n19209, n19210, n19211, n19213, n19214, n19215, n19217, 
      n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, 
      n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, 
      n19237, n19238, n19239, n19241, n19242, n19243, n19244, n19245, n19246, 
      n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, 
      n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, 
      n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, 
      n19274, n19275, n19276, n19277, n19278, n19279, n19281, n19282, n19283, 
      n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, 
      n19293, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, 
      n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, 
      n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, 
      n19321, n19322, n19323, n19325, n19326, n19327, n19328, n19329, n19330, 
      n19331, n19332, n19334, n19335, n19336, n19337, n19338, n19339, n19340, 
      n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, 
      n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19359, 
      n19360, n19361, n19363, n19364, n19365, n19366, n19367, n19368, n19369, 
      n19370, n19371, n19372, n19373, n19374, n19376, n19377, n19378, n19379, 
      n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, 
      n19389, n19390, n19391, n19392, n19393, n19395, n19396, n19397, n19398, 
      n19399, n19400, n19402, n19403, n19404, n19405, n19406, n19407, n19408, 
      n19409, n19410, n19411, n19412, n19413, n19414, n19416, n19417, n19418, 
      n19419, n19420, n19421, n19422, n19423, n19426, n19427, n19428, n19429, 
      n19430, n19431, n19432, n19433, n19435, n19436, n19437, n19438, n19439, 
      n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, 
      n19449, n19451, n19452, n19456, n19457, n19459, n19460, n19461, n19462, 
      n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, 
      n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, 
      n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19490, n19491, 
      n19492, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, 
      n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, 
      n19511, n19512, n19513, n19514, n19515, n19516, n19518, n19519, n19520, 
      n19521, n19522, n19523, n19525, n19526, n19527, n19528, n19529, n19530, 
      n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, 
      n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, 
      n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, 
      n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, 
      n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, 
      n19576, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, 
      n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19595, 
      n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, 
      n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, 
      n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, 
      n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, 
      n19632, n19633, n19634, n19636, n19637, n19638, n19639, n19640, n19641, 
      n19642, n19645, n19646, n19647, n19648, n19649, n19650, n19652, n19653, 
      n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, 
      n19663, n19664, n19665, n19666, n19667, n19668, n19671, n19672, n19673, 
      n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, 
      n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, 
      n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, 
      n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, 
      n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, 
      n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, 
      n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, 
      n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, 
      n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, 
      n19755, n19756, n19758, n19759, n19760, n19761, n19762, n19764, n19765, 
      n19766, n19767, n19768, n19769, n19772, n19773, n19774, n19776, n19777, 
      n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, 
      n19787, n19788, n19789, n19790, n19791, n19793, n19794, n19795, n19796, 
      n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19806, 
      n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, 
      n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, 
      n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, 
      n19836, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, 
      n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19854, n19855, 
      n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, 
      n19865, n19866, n19867, n19868, n19869, n19870, n19873, n19874, n19875, 
      n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, 
      n19885, n19886, n19887, n19888, n19889, n19892, n19893, n19894, n19895, 
      n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, 
      n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, 
      n19914, n19915, n19916, n19917, n19918, n19920, n19922, n19923, n19924, 
      n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, 
      n19934, n19935, n19936, n19937, n19938, n19939, n19941, n19942, n19943, 
      n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, 
      n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, 
      n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, 
      n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, 
      n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, 
      n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, 
      n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, 
      n20010, n20011, n20013, n20014, n20015, n20016, n20017, n20019, n20020, 
      n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, 
      n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, 
      n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, 
      n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, 
      n20058, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, 
      n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20076, n20077, 
      n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20086, n20087, 
      n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20098, 
      n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20109, 
      n20111, n20112, n20113, n20114, n20116, n20117, n20118, n20119, n20120, 
      n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, 
      n20130, n20131, n20133, n20134, n20135, n20136, n20137, n20138, n20139, 
      n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, 
      n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, 
      n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, 
      n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, 
      n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, 
      n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, 
      n20194, n20195, n20196, n20197, n20199, n20200, n20201, n20203, n20204, 
      n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, 
      n20214, n20215, n20216, n20217, n20218, n20220, n20221, n20222, n20223, 
      n20224, n20225, n20226, n20227, n20229, n20230, n20231, n20232, n20233, 
      n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, 
      n20243, n20244, n20247, n20248, n20249, n20250, n20251, n20252, n20253, 
      n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, 
      n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, 
      n20272, n20273, n20275, n20276, n20277, n20278, n20279, n20280, n20281, 
      n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, 
      n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, 
      n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, 
      n20309, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20319, 
      n20320, n20321, n20322, n20323, n20324, n20326, n20327, n20328, n20329, 
      n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, 
      n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, 
      n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, 
      n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, 
      n20367, n20368, n20369, n20370, n20372, n20373, n20374, n20375, n20376, 
      n20377, n20378, n20379, n20380, n20381, n20383, n20384, n20385, n20386, 
      n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, 
      n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, 
      n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, 
      n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, 
      n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, 
      n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, 
      n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, 
      n20450, n20451, n20452, n20455, n20456, n20457, n20458, n20459, n20460, 
      n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, 
      n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, 
      n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, 
      n20488, n20489, n20490, n20491, n20493, n20494, n20495, n20496, n20497, 
      n20498, n20499, n20501, n20502, n20503, n20504, n20505, n20507, n20508, 
      n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, 
      n20519, n20520, n20521, n20522, n20523, n20525, n20526, n20527, n20528, 
      n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, 
      n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, 
      n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, 
      n20557, n20558, n20559, n20560, n20561, n20562, n20564, n20565, n20566, 
      n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, 
      n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, 
      n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, 
      n20594, n20595, n20597, n20598, n20599, n20600, n20601, n20602, n20603, 
      n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, 
      n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, 
      n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, 
      n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, 
      n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, 
      n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, 
      n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, 
      n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, 
      n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, 
      n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, 
      n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, 
      n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, 
      n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, 
      n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, 
      n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, 
      n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, 
      n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, 
      n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, 
      n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, 
      n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, 
      n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, 
      n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, 
      n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, 
      n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, 
      n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, 
      n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, 
      n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, 
      n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, 
      n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, 
      n20865, n20866, n20867, n20868, n20870, n20871, n20872, n20873, n20874, 
      n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, 
      n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, 
      n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, 
      n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, 
      n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, 
      n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, 
      n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, 
      n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, 
      n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, 
      n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, 
      n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, 
      n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, 
      n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, 
      n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, 
      n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, 
      n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, 
      n21019, n21020, n21023, n21025, n21026, n21027, n21028, n21029, n21030, 
      n21031, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, 
      n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, 
      n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, 
      n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, 
      n21068, n21070, n21071, n21072, n21073, n21074, n21075, n21077, n21078, 
      n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, 
      n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, 
      n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, 
      n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, 
      n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, 
      n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, 
      n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, 
      n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, 
      n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, 
      n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, 
      n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, 
      n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, 
      n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, 
      n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, 
      n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, 
      n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, 
      n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, 
      n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, 
      n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, 
      n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, 
      n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, 
      n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, 
      n21278, n21279, n21281, n21282, n21283, n21284, n21285, n21286, n21287, 
      n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21296, n21297, 
      n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, 
      n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, 
      n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, 
      n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, 
      n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, 
      n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, 
      n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, 
      n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21370, 
      n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, 
      n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21389, n21390, 
      n21391, n21392, n21393, n21395, n21396, n21397, n21398, n21399, n21400, 
      n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, 
      n21410, n21411, n21413, n21414, n21415, n21416, n21417, n21418, n21419, 
      n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, 
      n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, 
      n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, 
      n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, 
      n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, 
      n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, 
      n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, 
      n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21492, 
      n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, 
      n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, 
      n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, 
      n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, 
      n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, 
      n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, 
      n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, 
      n21556, n21557, n21558, n21559, n21561, n21562, n21563, n21564, n21565, 
      n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, 
      n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, 
      n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, 
      n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, 
      n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, 
      n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, 
      n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, 
      n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, 
      n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, 
      n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, 
      n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, 
      n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, 
      n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, 
      n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, 
      n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, 
      n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, 
      n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, 
      n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, 
      n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, 
      n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, 
      n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, 
      n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, 
      n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, 
      n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21781, n21782, 
      n21783, n21784, n21785, n21786, n21788, n21789, n21790, n21791, n21792, 
      n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, 
      n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, 
      n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, 
      n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, 
      n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, 
      n21838, n21839, n21840, n21841, n21842, n21844, n21845, n21846, n21847, 
      n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, 
      n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, 
      n21866, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21876, 
      n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, 
      n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, 
      n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, 
      n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, 
      n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, 
      n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, 
      n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, 
      n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, 
      n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, 
      n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, 
      n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, 
      n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, 
      n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, 
      n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, 
      n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, 
      n22014, n22015, n22016, n22017, n22018, n22019, n22021, n22022, n22023, 
      n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, 
      n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, 
      n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, 
      n22052, n22053, n22054, n22055, n22056, n22058, n22059, n22060, n22061, 
      n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22070, n22071, 
      n22072, n22074, n22075, n22076, n22077, n22079, n22080, n22081, n22082, 
      n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, 
      n22092, n22093, n22095, n22096, n22097, n22099, n22100, n22101, n22102, 
      n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, 
      n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, 
      n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, 
      n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, 
      n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, 
      n22148, n22149, n22150, n22151, n22152, n22153, n22155, n22156, n22157, 
      n22158, n22159, n22161, n22162, n22163, n22164, n22165, n22166, n22168, 
      n22169, n22170, n22172, n22173, n22174, n22175, n22176, n22177, n22178, 
      n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, 
      n22188, n22190, n22191, n22192, n22193, n22194, n22195, n22197, n22198, 
      n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, 
      n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, 
      n22217, n22218, n22219, n22220, n22221, n22222, n22224, n22225, n22226, 
      n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, 
      n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, 
      n22245, n22246, n22247, n22248, n22252, n22253, n22254, n22255, n22257, 
      n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, 
      n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, 
      n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22284, n22285, 
      n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, 
      n22295, n22296, n22297, n22298, n22299, n22301, n22303, n22304, n22305, 
      n22306, n22307, n22308, n22309, n22311, n22312, n22313, n22314, n22315, 
      n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, 
      n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, 
      n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, 
      n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, 
      n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22361, 
      n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, 
      n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, 
      n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, 
      n22389, n22390, n22391, n22393, n22394, n22395, n22396, n22397, n22398, 
      n22399, n22400, n22401, n22403, n22404, n22405, n22406, n22407, n22408, 
      n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, 
      n22418, n22419, n22420, n22421, n22422, n22424, n22426, n22427, n22428, 
      n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, 
      n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22446, n22447, 
      n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, 
      n22458, n22459, n22461, n22462, n22463, n22464, n22465, n22466, n22468, 
      n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, 
      n22478, n22479, n22480, n22482, n22483, n22485, n22486, n22487, n22488, 
      n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, 
      n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, 
      n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, 
      n22516, n22517, n22518, n22519, n22521, n22522, n22523, n22524, n22525, 
      n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, 
      n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, 
      n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, 
      n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, 
      n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, 
      n22571, n22572, n22573, n22574, n22575, n22576, n22578, n22579, n22580, 
      n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, 
      n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, 
      n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, 
      n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, 
      n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, 
      n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, 
      n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, 
      n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, 
      n22654, n22655, n22656, n22657, n22658, n22659, n22661, n22663, n22664, 
      n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, 
      n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22685, n22686, 
      n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, 
      n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22705, 
      n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, 
      n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, 
      n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, 
      n22733, n22734, n22735, n22736, n22737, n22739, n22740, n22741, n22742, 
      n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22752, 
      n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, 
      n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, 
      n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22779, n22780, 
      n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, 
      n22791, n22792, n22794, n22795, n22796, n22797, n22798, n22799, n22800, 
      n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, 
      n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22820, n22821, 
      n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, 
      n22831, n22832, n22834, n22835, n22836, n22837, n22838, n22839, n22840, 
      n22841, n22842, n22846, n22847, n22848, n22849, n22850, n22851, n22852, 
      n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, 
      n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22870, n22872, 
      n22873, n22875, n22877, n22878, n22879, n22880, n22881, n22882, n22883, 
      n22884, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, 
      n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, 
      n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, 
      n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, 
      n22921, n22922, n22923, n22926, n22927, n22928, n22929, n22930, n22931, 
      n22932, n22933, n22934, n22935, n22936, n22938, n22939, n22940, n22941, 
      n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, 
      n22952, n22953, n22954, n22955, n22956, n22958, n22959, n22960, n22961, 
      n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, 
      n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, 
      n22980, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, 
      n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, 
      n22999, n23000, n23001, n23002, n23003, n23005, n23006, n23007, n23008, 
      n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, 
      n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, 
      n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, 
      n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, 
      n23045, n23046, n23047, n23048, n23049, n23050, n23052, n23053, n23054, 
      n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, 
      n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, 
      n23073, n23074, n23076, n23077, n23079, n23080, n23081, n23082, n23085, 
      n23086, n23087, n23088, n23089, n23090, n23091, n23093, n23094, n23095, 
      n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, 
      n23105, n23106, n23107, n23108, n23109, n23110, n23112, n23113, n23114, 
      n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, 
      n23124, n23125, n23126, n23127, n23128, n23129, n23131, n23132, n23133, 
      n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, 
      n23143, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, 
      n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, 
      n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, 
      n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, 
      n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, 
      n23189, n23190, n23191, n23193, n23194, n23195, n23196, n23199, n23200, 
      n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, 
      n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, 
      n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, 
      n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, 
      n23237, n23238, n23239, n23241, n23242, n23243, n23244, n23245, n23247, 
      n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256, 
      n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, 
      n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274, 
      n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, 
      n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, 
      n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, 
      n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, 
      n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, 
      n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, 
      n23329, n23330, n23331, n23332, n23334, n23335, n23336, n23337, n23338, 
      n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, 
      n23348, n23349, n23350, n23353, n23354, n23355, n23356, n23357, n23358, 
      n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, 
      n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, 
      n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, 
      n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, 
      n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, 
      n23405, n23406, n23407, n23408, n23410, n23411, n23413, n23414, n23416, 
      n23417, n23418, n23419, n23420, n23422, n23423, n23424, n23425, n23426, 
      n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435, 
      n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444, 
      n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453, 
      n23454, n23455, n23456, n23458, n23460, n23461, n23462, n23463, n23464, 
      n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473, 
      n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482, 
      n23483, n23484, n23485, n23487, n23488, n23489, n23490, n23491, n23492, 
      n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, 
      n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, 
      n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, 
      n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, 
      n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, 
      n23539, n23540, n23541, n23542, n23543, n23544, n23546, n23547, n23548, 
      n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, 
      n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, 
      n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, 
      n23578, n23579, n23580, n23581, n23582, n23583, n23585, n23586, n23587, 
      n23588, n23589, n23590, n23591, n23592, n23594, n23595, n23596, n23597, 
      n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606, 
      n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615, 
      n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624, 
      n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23634, 
      n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, 
      n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, 
      n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, 
      n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, 
      n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, 
      n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23688, n23689, 
      n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, 
      n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, 
      n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, 
      n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, 
      n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, 
      n23735, n23736, n23737, n23738, n23739, n23740, n23742, n23743, n23744, 
      n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, 
      n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, 
      n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, 
      n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, 
      n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, 
      n23790, n23791, n23792, n23793, n23796, n23798, n23799, n23801, n23802, 
      n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, 
      n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23820, n23821, 
      n23822, n23823, n23824, n23825, n23827, n23828, n23829, n23830, n23831, 
      n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840, 
      n23841, n23842, n23843, n23844, n23846, n23847, n23849, n23850, n23851, 
      n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, 
      n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, 
      n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, 
      n23881, n23882, n23883, n23885, n23886, n23887, n23888, n23889, n23890, 
      n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, 
      n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, 
      n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, 
      n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926, 
      n23927, n23928, n23929, n23930, n23931, n23933, n23934, n23935, n23936, 
      n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945, 
      n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954, 
      n23955, n23956, n23958, n23959, n23960, n23961, n23962, n23963, n23964, 
      n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, 
      n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, 
      n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, 
      n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, 
      n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, 
      n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, 
      n24019, n24020, n24025, n24026, n24027, n24037, n24042, n24043, n24050, 
      n24051, n24054, n24056, n24057, n24059, n24061, n24062, n24063, n24064, 
      n24065, n24067, n24072, n24074, n24075, n24076, n24077, n24078, n24079, 
      n24080, n24082, n24083, n24084, n24085, n24087, n24089, n24090, n24091, 
      n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, 
      n24101, n24103, n24104, n24106, n24107, n24108, n24109, n24110, n24112, 
      n24113, n24114, n24115, n24116, n24118, n24119, n24120, n24121, n24123, 
      n24124, n24125, n24127, n24128, n24130, n24131, n24132, n24133, n24134, 
      n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24143, n24144, 
      n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, 
      n24155, n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, 
      n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24174, n24177, 
      n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, 
      n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, 
      n24196, n24197, n24198, n24199, n24200, n24202, n24203, n24204, n24205, 
      n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24217, n24218, 
      n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, 
      n24229, n24230, n24231, n24233, n24234, n24236, n24237, n24238, n24239, 
      n24240, n24241, n24242, n24243, n24244, n24246, n24247, n24248, n24249, 
      n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, 
      n24259, n24260, n24261, n24262, n24264, n24265, n24267, n24269, n24270, 
      n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, 
      n24281, n24283, n24284, n24285, n24286, n24287, n24288, n24291, n24292, 
      n24293, n24294, n24295, n24296, n24297, n24299, n24300, n24301, n24302, 
      n24303, n24304, n24305, n24306, n24307, n24309, n24310, n24311, n24312, 
      n24313, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, 
      n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24332, 
      n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, 
      n24342, n24343, n24344, n24345, n24346, n24347, n24349, n24350, n24351, 
      n24352, n24353, n24354, n24356, n24357, n24360, n24361, n24362, n24364, 
      n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374, 
      n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24383, n24384, 
      n24385, n24386, n24387, n24389, n24390, n24391, n24392, n24393, n24394, 
      n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, 
      n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, 
      n24413, n24414, n24415, n24416, n24418, n24420, n24421, n24422, n24423, 
      n24424, n24426, n24427, n24428, n24429, n24430, n24431, n24433, n24434, 
      n24435, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, 
      n24447, n24448, n24449, n24451, n24452, n24453, n24454, n24456, n24457, 
      n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, 
      n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475, 
      n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484, 
      n24485, n24486, n24487, n24488, n24490, n24491, n24492, n24493, n24494, 
      n24495, n24496, n24498, n24499, n24500, n24501, n24502, n24503, n24505, 
      n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, 
      n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24525, 
      n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, 
      n24535, n24536, n24537, n24539, n24540, n24542, n24543, n24547, n24549, 
      n24550, n24551, n24552, n24554, n24556, n24558, n24559, n24561, n24565, 
      n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575, 
      n24576, n24577, n24578, n24579, n24581, n24582, n24583, n24584, n24585, 
      n24586, n24587, n24588, n24589, n24591, n24592, n24594, n24595, n24596, 
      n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605, 
      n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24615, 
      n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, 
      n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634, 
      n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643, 
      n24644, n24646, n24647, n24648, n24650, n24652, n24653, n24654, n24655, 
      n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24664, n24665, 
      n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, 
      n24675, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, 
      n24685, n24686, n24687, n24688, n24689, n24691, n24692, n24694, n24697, 
      n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24706, n24707, 
      n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, 
      n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, 
      n24727, n24728, n24729, n24730, n24733, n24734, n24735, n24736, n24737, 
      n24738, n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, 
      n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, 
      n24758, n24759, n24760, n24761, n24763, n24764, n24765, n24767, n24768, 
      n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, 
      n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, 
      n24787, n24788, n24789, n24790, n24791, n24792, n24794, n24795, n24796, 
      n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805, 
      n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814, 
      n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823, 
      n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832, 
      n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24841, n24842, 
      n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24851, n24852, 
      n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, 
      n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, 
      n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, 
      n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, 
      n24889, n24890, n24891, n24892, n24893, n24895, n24896, n24897, n24898, 
      n24899, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, 
      n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917, 
      n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24926, n24927, 
      n24928, n24929, n24930, n24931, n24932, n24933, n24935, n24936, n24937, 
      n24938, n24940, n24941, n24942, n24943, n24944, n24946, n24947, n24948, 
      n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, 
      n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, 
      n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, 
      n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, 
      n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, 
      n24994, n24995, n24996, n24998, n24999, n25000, n25001, n25002, n25003, 
      n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012, 
      n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, 
      n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, 
      n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039, 
      n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048, 
      n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25057, n25058, 
      n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, 
      n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, 
      n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, 
      n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, 
      n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, 
      n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, 
      n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, 
      n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, 
      n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, 
      n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, 
      n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, 
      n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, 
      n25167, n25168, n25169, n25170, n25172, n25173, n25174, n25175, n25176, 
      n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, 
      n25186, n25187, n25188, n25189, n25191, n25192, n25193, n25194, n25195, 
      n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, 
      n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, 
      n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, 
      n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, 
      n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, 
      n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, 
      n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, 
      n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, 
      n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, 
      n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, 
      n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, 
      n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, 
      n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, 
      n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, 
      n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, 
      n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, 
      n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, 
      n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, 
      n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366, 
      n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375, 
      n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384, 
      n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, 
      n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, 
      n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, 
      n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, 
      n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, 
      n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438, 
      n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, 
      n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, 
      n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465, 
      n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474, 
      n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, 
      n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, 
      n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, 
      n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, 
      n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519, 
      n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528, 
      n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537, 
      n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546, 
      n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, 
      n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, 
      n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, 
      n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, 
      n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, 
      n25592, n25593, n25594, n25595, n25596, n25597 : std_logic;

begin
   
   U5 : BUF_X1 port map( A => n22354, Z => n245);
   U8 : XNOR2_X1 port map( A => n21451, B => n21450, ZN => n22962);
   U10 : XNOR2_X1 port map( A => n21980, B => n21745, ZN => n21454);
   U16 : OR2_X1 port map( A1 => n20230, A2 => n20498, ZN => n170);
   U17 : OR2_X1 port map( A1 => n20214, A2 => n20215, ZN => n197);
   U18 : INV_X1 port map( A => n20464, ZN => n20458);
   U19 : INV_X1 port map( A => n20618, ZN => n7);
   U20 : OR2_X1 port map( A1 => n3428, A2 => n20373, ZN => n771);
   U22 : INV_X1 port map( A => n20216, ZN => n100);
   U26 : OR2_X1 port map( A1 => n19379, A2 => n19381, ZN => n4007);
   U28 : OR2_X1 port map( A1 => n19381, A2 => n19380, ZN => n19204);
   U30 : NAND2_X1 port map( A1 => n19039, A2 => n24582, ZN => n194);
   U36 : INV_X1 port map( A => n16037, ZN => n18516);
   U40 : INV_X1 port map( A => n365, ZN => n46);
   U41 : INV_X1 port map( A => n17043, ZN => n17373);
   U49 : INV_X1 port map( A => n3544, ZN => n41);
   U50 : OR2_X1 port map( A1 => n14926, A2 => n16028, ZN => n161);
   U51 : OR2_X1 port map( A1 => n15694, A2 => n16062, ZN => n15600);
   U52 : INV_X1 port map( A => n16428, ZN => n15958);
   U54 : XNOR2_X1 port map( A => n15096, B => n12, ZN => n15100);
   U56 : INV_X1 port map( A => n15358, ZN => n75);
   U57 : INV_X1 port map( A => n15422, ZN => n14442);
   U59 : OR2_X1 port map( A1 => n14340, A2 => n25197, ZN => n76);
   U60 : OR2_X1 port map( A1 => n13921, A2 => n13653, ZN => n96);
   U61 : OR2_X1 port map( A1 => n13956, A2 => n13733, ZN => n813);
   U62 : AND2_X1 port map( A1 => n12704, A2 => n14078, ZN => n13628);
   U63 : AND3_X1 port map( A1 => n25435, A2 => n14235, A3 => n24402, ZN => n182
                           );
   U66 : INV_X1 port map( A => n14209, ZN => n13811);
   U67 : OR2_X1 port map( A1 => n13953, A2 => n24999, ZN => n507);
   U69 : OR2_X1 port map( A1 => n13209, A2 => n13208, ZN => n136);
   U70 : NAND2_X1 port map( A1 => n10395, A2 => n10394, ZN => n508);
   U74 : AND2_X1 port map( A1 => n13222, A2 => n13227, ZN => n29);
   U76 : AND2_X1 port map( A1 => n12454, A2 => n13061, ZN => n4320);
   U78 : INV_X1 port map( A => n11892, ZN => n12257);
   U85 : INV_X1 port map( A => n10630, ZN => n44);
   U86 : OAI21_X1 port map( B1 => n11338, B2 => n24082, A => n10491, ZN => 
                           n11935);
   U90 : OAI211_X1 port map( C1 => n25, C2 => n9817, A => n25046, B => n24, ZN 
                           => n655);
   U93 : AND2_X1 port map( A1 => n25069, A2 => n9886, ZN => n52);
   U94 : INV_X1 port map( A => n10148, ZN => n10120);
   U96 : XNOR2_X1 port map( A => n8505, B => n8504, ZN => n8521);
   U98 : CLKBUF_X1 port map( A => Key(174), Z => n187);
   U104 : NAND2_X1 port map( A1 => n7815, A2 => n9070, ZN => n8507);
   U106 : OR2_X1 port map( A1 => n248, A2 => n7232, ZN => n3192);
   U107 : OR2_X1 port map( A1 => n7099, A2 => n127, ZN => n126);
   U108 : OR2_X1 port map( A1 => n7522, A2 => n23, ZN => n2949);
   U110 : BUF_X1 port map( A => n7057, Z => n9068);
   U111 : INV_X1 port map( A => n7526, ZN => n23);
   U115 : MUX2_X1 port map( A => n6107, B => n6108, S => n7033, Z => n7526);
   U116 : AND2_X1 port map( A1 => n4672, A2 => n7947, ZN => n13);
   U118 : OR2_X1 port map( A1 => n6945, A2 => n6944, ZN => n70);
   U123 : AND2_X1 port map( A1 => n23252, A2 => n3720, ZN => n23254);
   U124 : NOR2_X1 port map( A1 => n7284, A2 => n7776, ZN => n7522);
   U127 : NAND2_X1 port map( A1 => n17691, A2 => n17690, ZN => n18004);
   U129 : OR2_X1 port map( A1 => n13345, A2 => n12859, ZN => n13349);
   U130 : INV_X1 port map( A => n22982, ZN => n22530);
   U133 : AND2_X1 port map( A1 => n16449, A2 => n223, ZN => n131);
   U135 : OR2_X1 port map( A1 => n7781, A2 => n7787, ZN => n5266);
   U137 : NOR2_X1 port map( A1 => n22987, A2 => n23379, ZN => n22988);
   U139 : OR2_X1 port map( A1 => n18994, A2 => n20319, ZN => n615);
   U142 : AND2_X1 port map( A1 => n23505, A2 => n3978, ZN => n23513);
   U145 : NOR2_X1 port map( A1 => n23937, A2 => n24948, ZN => n104);
   U147 : OR2_X1 port map( A1 => n22729, A2 => n22093, ZN => n20893);
   U148 : OR2_X1 port map( A1 => n23479, A2 => n23478, ZN => n22736);
   U156 : NAND2_X1 port map( A1 => n17620, A2 => n17623, ZN => n16901);
   U158 : MUX2_X2 port map( A => n20254, B => n20253, S => n21844, Z => n23860)
                           ;
   U162 : INV_X1 port map( A => n10168, ZN => n25);
   U163 : OR2_X1 port map( A1 => n10168, A2 => n10169, ZN => n24);
   U164 : BUF_X1 port map( A => n13453, Z => n14302);
   U166 : XNOR2_X2 port map( A => n2633, B => n2634, ZN => n23014);
   U167 : AND2_X2 port map( A1 => n2568, A2 => n2567, ZN => n2569);
   U170 : OAI21_X1 port map( B1 => n10028, B2 => n4787, A => n9023, ZN => 
                           n10941);
   U171 : OR2_X1 port map( A1 => n20183, A2 => n20042, ZN => n113);
   U172 : XNOR2_X1 port map( A => n11440, B => n11640, ZN => n12073);
   U174 : INV_X1 port map( A => n20913, ZN => n347);
   U178 : OAI22_X1 port map( A1 => n10793, A2 => n11196, B1 => n11199, B2 => 
                           n10789, ZN => n10628);
   U180 : OR2_X1 port map( A1 => n6819, A2 => n6895, ZN => n190);
   U181 : NAND2_X1 port map( A1 => n23393, A2 => n22026, ZN => n23386);
   U183 : NAND3_X1 port map( A1 => n24585, A2 => n16932, A3 => n17054, ZN => 
                           n3593);
   U187 : NAND2_X1 port map( A1 => n24589, A2 => n13386, ZN => n1);
   U188 : NAND2_X1 port map( A1 => n13644, A2 => n25011, ZN => n3);
   U190 : NAND2_X1 port map( A1 => n2801, A2 => n4, ZN => n7829);
   U193 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n20088);
   U194 : NAND2_X1 port map( A1 => n20084, A2 => n24338, ZN => n5);
   U195 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n6);
   U196 : NAND2_X1 port map( A1 => n20570, A2 => n20616, ZN => n8);
   U198 : NOR2_X1 port map( A1 => n25469, A2 => n9, ZN => n1988);
   U199 : NOR2_X1 port map( A1 => n19170, A2 => n19173, ZN => n9);
   U202 : XNOR2_X1 port map( A => n18044, B => n17590, ZN => n10);
   U205 : BUF_X1 port map( A => n6849, Z => n249);
   U208 : XNOR2_X2 port map( A => n14884, B => n11, ZN => n16595);
   U209 : XNOR2_X1 port map( A => n15176, B => n12451, ZN => n11);
   U210 : OAI21_X1 port map( B1 => n24397, B2 => n23595, A => n21944, ZN => 
                           n21945);
   U214 : NAND3_X1 port map( A1 => n5296, A2 => n10930, A3 => n10596, ZN => 
                           n4213);
   U215 : AOI22_X1 port map( A1 => n13813, A2 => n14209, B1 => n3340, B2 => 
                           n13422, ZN => n12982);
   U216 : NAND2_X1 port map( A1 => n13421, A2 => n1314, ZN => n14209);
   U218 : NAND2_X1 port map( A1 => n4259, A2 => n13, ZN => n7949);
   U220 : OR2_X2 port map( A1 => n2773, A2 => n7951, ZN => n9149);
   U221 : NAND2_X1 port map( A1 => n7035, A2 => n25424, ZN => n6105);
   U223 : NOR2_X1 port map( A1 => n3333, A2 => n3334, ZN => n14);
   U226 : AOI22_X1 port map( A1 => n8841, A2 => n15, B1 => n8842, B2 => n9729, 
                           ZN => n10523);
   U227 : OAI21_X1 port map( B1 => n9493, B2 => n426, A => n9731, ZN => n15);
   U239 : NAND2_X1 port map( A1 => n9558, A2 => n4454, ZN => n777);
   U240 : NAND3_X1 port map( A1 => n13964, A2 => n13962, A3 => n13963, ZN => 
                           n3801);
   U244 : NOR2_X1 port map( A1 => n25246, A2 => n17419, ZN => n17226);
   U247 : NAND2_X1 port map( A1 => n3356, A2 => n25292, ZN => n20);
   U248 : OR2_X1 port map( A1 => n13010, A2 => n12919, ZN => n21);
   U249 : NAND3_X1 port map( A1 => n20519, A2 => n351, A3 => n22, ZN => n73);
   U252 : NAND2_X2 port map( A1 => n660, A2 => n9616, ZN => n11205);
   U257 : AOI22_X2 port map( A1 => n20222, A2 => n20272, B1 => n20515, B2 => 
                           n20221, ZN => n21568);
   U259 : NAND2_X1 port map( A1 => n17267, A2 => n15673, ZN => n26);
   U260 : NAND2_X1 port map( A1 => n16710, A2 => n17326, ZN => n27);
   U261 : NAND3_X1 port map( A1 => n10001, A2 => n10002, A3 => n10000, ZN => 
                           n10004);
   U263 : AOI21_X1 port map( B1 => n6782, B2 => n6781, A => n6780, ZN => n28);
   U265 : NAND2_X1 port map( A1 => n12924, A2 => n29, ZN => n12571);
   U267 : NAND2_X2 port map( A1 => n608, A2 => n9204, ZN => n10585);
   U269 : XNOR2_X2 port map( A => n5952, B => Key(169), ZN => n6488);
   U270 : NAND2_X1 port map( A1 => n12984, A2 => n780, ZN => n779);
   U272 : NAND3_X1 port map( A1 => n4296, A2 => n8026, A3 => n8025, ZN => n9040
                           );
   U280 : INV_X1 port map( A => n11598, ZN => n31);
   U281 : OR3_X1 port map( A1 => n7909, A2 => n7155, A3 => n7908, ZN => n7156);
   U284 : XNOR2_X1 port map( A => n15443, B => n15442, ZN => n15545);
   U285 : NOR2_X1 port map( A1 => n13028, A2 => n13023, ZN => n11406);
   U286 : NAND2_X1 port map( A1 => n34, A2 => n32, ZN => n13854);
   U287 : NAND2_X1 port map( A1 => n12549, A2 => n24220, ZN => n32);
   U291 : NAND3_X2 port map( A1 => n2424, A2 => n12575, A3 => n2423, ZN => 
                           n13845);
   U294 : AND2_X1 port map( A1 => n18902, A2 => n18772, ZN => n762);
   U295 : BUF_X1 port map( A => n9269, Z => n9947);
   U296 : NAND2_X1 port map( A1 => n38, A2 => n24527, ZN => n14044);
   U298 : NAND2_X1 port map( A1 => n3559, A2 => n3558, ZN => n38);
   U301 : INV_X1 port map( A => n18465, ZN => n39);
   U302 : AND3_X2 port map( A1 => n3251, A2 => n3250, A3 => n3252, ZN => n11564
                           );
   U304 : NAND2_X1 port map( A1 => n42, A2 => n41, ZN => n40);
   U306 : NAND3_X2 port map( A1 => n2750, A2 => n6219, A3 => n2749, ZN => n8341
                           );
   U312 : NAND2_X1 port map( A1 => n9064, A2 => n10050, ZN => n9539);
   U313 : OR2_X1 port map( A1 => n10751, A2 => n10904, ZN => n10900);
   U316 : OR2_X2 port map( A1 => n7244, A2 => n7243, ZN => n8501);
   U325 : OAI21_X1 port map( B1 => n2119, B2 => n6734, A => n2118, ZN => n6064)
                           ;
   U329 : OAI21_X1 port map( B1 => n16539, B2 => n17633, A => n45, ZN => n16792
                           );
   U331 : MUX2_X2 port map( A => n22971, B => n22970, S => n22969, Z => n23350)
                           ;
   U332 : XNOR2_X1 port map( A => n47, B => n2735, ZN => Ciphertext(74));
   U333 : NAND3_X1 port map( A1 => n4605, A2 => n21955, A3 => n4607, ZN => n47)
                           ;
   U335 : NAND2_X2 port map( A1 => n9415, A2 => n4655, ZN => n10767);
   U338 : NAND2_X1 port map( A1 => n2821, A2 => n13438, ZN => n48);
   U346 : OAI21_X1 port map( B1 => n52, B2 => n9887, A => n51, ZN => n9890);
   U347 : NAND2_X1 port map( A1 => n9887, A2 => n9888, ZN => n51);
   U356 : INV_X1 port map( A => n20291, ZN => n55);
   U357 : NAND2_X1 port map( A1 => n6301, A2 => n6488, ZN => n6430);
   U361 : NAND2_X1 port map( A1 => n17572, A2 => n17042, ZN => n17043);
   U363 : NAND2_X1 port map( A1 => n1148, A2 => n6977, ZN => n6691);
   U364 : NAND2_X1 port map( A1 => n1649, A2 => n10141, ZN => n1648);
   U368 : XNOR2_X2 port map( A => n5913, B => Key(18), ZN => n5916);
   U369 : NAND2_X1 port map( A1 => n13236, A2 => n4499, ZN => n12937);
   U375 : NAND2_X1 port map( A1 => n2922, A2 => n9486, ZN => n9487);
   U376 : NAND3_X1 port map( A1 => n10181, A2 => n58, A3 => n10182, ZN => 
                           n10183);
   U377 : NAND2_X1 port map( A1 => n10179, A2 => n10178, ZN => n58);
   U380 : NAND3_X1 port map( A1 => n4846, A2 => n2259, A3 => n16355, ZN => 
                           n2258);
   U382 : NAND2_X1 port map( A1 => n13550, A2 => n14210, ZN => n59);
   U383 : NAND2_X1 port map( A1 => n6881, A2 => n6076, ZN => n6643);
   U384 : NAND2_X1 port map( A1 => n60, A2 => n942, ZN => n941);
   U385 : NAND2_X1 port map( A1 => n767, A2 => n6154, ZN => n60);
   U391 : NOR2_X2 port map( A1 => n13087, A2 => n13086, ZN => n13712);
   U392 : NAND2_X1 port map( A1 => n2938, A2 => n2941, ZN => n13087);
   U393 : OAI21_X1 port map( B1 => n3016, B2 => n20498, A => n61, ZN => n20270)
                           ;
   U398 : OAI21_X1 port map( B1 => n7228, B2 => n4812, A => n7947, ZN => n4811)
                           ;
   U400 : OR2_X1 port map( A1 => n15557, A2 => n25410, ZN => n15750);
   U404 : AOI22_X2 port map( A1 => n1570, A2 => n11038, B1 => n11040, B2 => 
                           n11039, ZN => n11983);
   U411 : NOR2_X1 port map( A1 => n23462, A2 => n22733, ZN => n23020);
   U412 : NAND2_X1 port map( A1 => n6052, A2 => n6051, ZN => n6054);
   U413 : NAND3_X1 port map( A1 => n16021, A2 => n287, A3 => n16846, ZN => 
                           n16027);
   U415 : NAND3_X1 port map( A1 => n7977, A2 => n3567, A3 => n3618, ZN => n7516
                           );
   U418 : AND3_X2 port map( A1 => n1873, A2 => n3613, A3 => n3612, ZN => n8807)
                           ;
   U419 : AOI22_X2 port map( A1 => n14025, A2 => n13877, B1 => n14334, B2 => 
                           n14333, ZN => n13595);
   U420 : NAND2_X1 port map( A1 => n66, A2 => n19032, ZN => n4245);
   U421 : NAND2_X1 port map( A1 => n19030, A2 => n19031, ZN => n66);
   U422 : INV_X1 port map( A => n25215, ZN => n370);
   U423 : NAND2_X1 port map( A1 => n24569, A2 => n25215, ZN => n5763);
   U431 : AOI21_X2 port map( B1 => n7488, B2 => n7487, A => n7486, ZN => n9081)
                           ;
   U432 : XNOR2_X1 port map( A => n68, B => n2319, ZN => Ciphertext(11));
   U433 : OAI211_X1 port map( C1 => n23082, C2 => n22578, A => n23081, B => 
                           n23080, ZN => n68);
   U436 : NAND2_X1 port map( A1 => n730, A2 => n3320, ZN => n7758);
   U438 : NAND2_X1 port map( A1 => n2387, A2 => n10884, ZN => n3416);
   U439 : NAND2_X1 port map( A1 => n2597, A2 => n22373, ZN => n2596);
   U442 : NAND2_X1 port map( A1 => n16717, A2 => n69, ZN => n2823);
   U443 : NAND3_X1 port map( A1 => n16715, A2 => n17598, A3 => n17596, ZN => 
                           n69);
   U445 : NAND2_X1 port map( A1 => n2996, A2 => n24458, ZN => n14382);
   U451 : NAND2_X1 port map( A1 => n1614, A2 => n1590, ZN => n71);
   U452 : NAND3_X1 port map( A1 => n73, A2 => n1438, A3 => n72, ZN => n21675);
   U453 : NAND2_X1 port map( A1 => n200, A2 => n20272, ZN => n72);
   U455 : AND2_X1 port map( A1 => n22889, A2 => n22093, ZN => n21774);
   U458 : NAND2_X1 port map( A1 => n13501, A2 => n13878, ZN => n13511);
   U459 : XNOR2_X1 port map( A => n15506, B => n75, ZN => n15361);
   U462 : NAND2_X1 port map( A1 => n17077, A2 => n17478, ZN => n16897);
   U466 : NAND3_X2 port map( A1 => n16374, A2 => n3775, A3 => n3774, ZN => 
                           n18532);
   U468 : NAND3_X1 port map( A1 => n616, A2 => n9071, A3 => n7430, ZN => n775);
   U469 : NAND2_X1 port map( A1 => n16210, A2 => n1496, ZN => n17387);
   U471 : NAND3_X1 port map( A1 => n6171, A2 => n6350, A3 => n6169, ZN => n77);
   U475 : NAND2_X1 port map( A1 => n22678, A2 => n23997, ZN => n2618);
   U478 : NAND2_X1 port map( A1 => n5208, A2 => n20193, ZN => n5207);
   U481 : NAND3_X1 port map( A1 => n10927, A2 => n10924, A3 => n10327, ZN => 
                           n10328);
   U483 : NAND3_X1 port map( A1 => n20388, A2 => n19345, A3 => n240, ZN => 
                           n19023);
   U484 : NAND2_X1 port map( A1 => n992, A2 => n78, ZN => n15757);
   U485 : NAND2_X1 port map( A1 => n16002, A2 => n16267, ZN => n78);
   U487 : BUF_X1 port map( A => n5902, Z => n6950);
   U489 : AOI21_X2 port map( B1 => n17410, B2 => n15026, A => n79, ZN => n18326
                           );
   U490 : OAI21_X1 port map( B1 => n17410, B2 => n17257, A => n15025, ZN => n79
                           );
   U493 : XNOR2_X2 port map( A => Key(61), B => Plaintext(61), ZN => n6963);
   U496 : NAND2_X1 port map( A1 => n2767, A2 => n17013, ZN => n4005);
   U499 : NAND2_X1 port map( A1 => n131, A2 => n16236, ZN => n16237);
   U500 : MUX2_X1 port map( A => n13073, B => n12532, S => n13067, Z => n12475)
                           ;
   U503 : BUF_X1 port map( A => n7147, Z => n7699);
   U508 : AND2_X2 port map( A1 => n6837, A2 => n467, ZN => n7989);
   U520 : NAND2_X1 port map( A1 => n81, A2 => n6540, ZN => n6167);
   U521 : NAND2_X1 port map( A1 => n5916, A2 => n6162, ZN => n81);
   U524 : NAND3_X2 port map( A1 => n13772, A2 => n82, A3 => n13771, ZN => 
                           n14775);
   U527 : INV_X1 port map( A => n22736, ZN => n23469);
   U528 : NAND2_X1 port map( A1 => n25191, A2 => n12928, ZN => n1971);
   U529 : NAND3_X2 port map( A1 => n3039, A2 => n136, A3 => n13214, ZN => 
                           n13988);
   U531 : NAND3_X2 port map( A1 => n7493, A2 => n7491, A3 => n7492, ZN => n3715
                           );
   U535 : BUF_X1 port map( A => n22575, Z => n23194);
   U538 : XNOR2_X1 port map( A => n85, B => n1875, ZN => Ciphertext(33));
   U539 : NOR2_X1 port map( A1 => n462, A2 => n22576, ZN => n85);
   U541 : INV_X1 port map( A => n20572, ZN => n87);
   U542 : XNOR2_X2 port map( A => n14681, B => n14680, ZN => n16109);
   U545 : NAND2_X1 port map( A1 => n88, A2 => n16124, ZN => n16127);
   U546 : NAND2_X1 port map( A1 => n578, A2 => n381, ZN => n88);
   U548 : NAND3_X1 port map( A1 => n24103, A2 => n7897, A3 => n24861, ZN => 
                           n5235);
   U549 : AOI21_X2 port map( B1 => n89, B2 => n10852, A => n2959, ZN => n11703)
                           ;
   U550 : NAND2_X1 port map( A1 => n1167, A2 => n10847, ZN => n89);
   U551 : NAND2_X1 port map( A1 => n14028, A2 => n13877, ZN => n13880);
   U559 : NAND3_X2 port map( A1 => n5388, A2 => n1749, A3 => n1405, ZN => n9188
                           );
   U560 : INV_X1 port map( A => n17099, ZN => n15869);
   U561 : NAND2_X1 port map( A1 => n17120, A2 => n17119, ZN => n17099);
   U564 : NAND2_X1 port map( A1 => n24378, A2 => n20102, ZN => n21035);
   U573 : INV_X1 port map( A => n11092, ZN => n11090);
   U574 : NAND2_X1 port map( A1 => n95, A2 => n11092, ZN => n10764);
   U575 : NAND3_X2 port map( A1 => n5362, A2 => n9535, A3 => n9534, ZN => 
                           n11092);
   U577 : XNOR2_X1 port map( A => n8541, B => n8540, ZN => n9495);
   U587 : OAI211_X2 port map( C1 => n15809, C2 => n15808, A => n15807, B => 
                           n15806, ZN => n18289);
   U588 : NAND3_X2 port map( A1 => n13381, A2 => n97, A3 => n96, ZN => n14620);
   U589 : NAND2_X1 port map( A1 => n13985, A2 => n13918, ZN => n97);
   U592 : NAND2_X1 port map( A1 => n25347, A2 => n20216, ZN => n101);
   U594 : NAND3_X2 port map( A1 => n15264, A2 => n3121, A3 => n15265, ZN => 
                           n17342);
   U596 : NAND2_X1 port map( A1 => n9487, A2 => n9488, ZN => n102);
   U599 : XNOR2_X2 port map( A => n5779, B => Key(91), ZN => n6712);
   U600 : NAND2_X1 port map( A1 => n3407, A2 => n6277, ZN => n791);
   U601 : NAND2_X1 port map( A1 => n6517, A2 => n315, ZN => n6277);
   U602 : OAI21_X1 port map( B1 => n15783, B2 => n4678, A => n2478, ZN => n2891
                           );
   U604 : OAI21_X2 port map( B1 => n6387, B2 => n6386, A => n6385, ZN => n3979)
                           ;
   U610 : BUF_X1 port map( A => n19250, Z => n1551);
   U612 : NAND3_X1 port map( A1 => n7718, A2 => n7715, A3 => n24577, ZN => 
                           n7560);
   U613 : NAND2_X1 port map( A1 => n23859, A2 => n23843, ZN => n22982);
   U616 : AOI22_X2 port map( A1 => n3191, A2 => n103, B1 => n10077, B2 => 
                           n10078, ZN => n12053);
   U617 : INV_X1 port map( A => n11002, ZN => n103);
   U618 : NAND2_X1 port map( A1 => n5342, A2 => n5119, ZN => n11002);
   U619 : NAND2_X1 port map( A1 => n23924, A2 => n104, ZN => n23915);
   U631 : NAND2_X1 port map( A1 => n1015, A2 => n1016, ZN => n1014);
   U634 : OAI211_X2 port map( C1 => n6750, C2 => n6749, A => n6748, B => n6747,
                           ZN => n7674);
   U640 : INV_X1 port map( A => n457, ZN => n19325);
   U641 : NAND2_X1 port map( A1 => n3748, A2 => n17872, ZN => n457);
   U646 : NAND2_X1 port map( A1 => n3302, A2 => n108, ZN => n3301);
   U647 : OR2_X1 port map( A1 => n14156, A2 => n5080, ZN => n108);
   U649 : XNOR2_X2 port map( A => Key(63), B => Plaintext(63), ZN => n5800);
   U651 : NAND2_X1 port map( A1 => n19244, A2 => n19615, ZN => n109);
   U654 : NAND3_X1 port map( A1 => n12652, A2 => n10360, A3 => n13177, ZN => 
                           n10394);
   U656 : NAND2_X1 port map( A1 => n15639, A2 => n16187, ZN => n2051);
   U659 : BUF_X2 port map( A => n17845, Z => n19464);
   U660 : NAND3_X1 port map( A1 => n3549, A2 => n7500, A3 => n7991, ZN => n2748
                           );
   U663 : AOI21_X2 port map( B1 => n15761, B2 => n3406, A => n15760, ZN => 
                           n17478);
   U666 : NAND2_X1 port map( A1 => n11199, A2 => n10630, ZN => n4047);
   U668 : XNOR2_X1 port map( A => n15072, B => n15073, ZN => n112);
   U670 : NOR2_X1 port map( A1 => n16350, A2 => n24467, ZN => n3333);
   U671 : NAND2_X1 port map( A1 => n16597, A2 => n15822, ZN => n16350);
   U677 : NAND2_X1 port map( A1 => n5462, A2 => n16732, ZN => n3306);
   U679 : NAND2_X1 port map( A1 => n19398, A2 => n24326, ZN => n114);
   U680 : NAND2_X1 port map( A1 => n19399, A2 => n18899, ZN => n115);
   U685 : OAI21_X1 port map( B1 => n3655, B2 => n16876, A => n17356, ZN => n119
                           );
   U687 : NAND2_X1 port map( A1 => n16546, A2 => n17068, ZN => n16733);
   U689 : AND2_X1 port map( A1 => n14124, A2 => n3341, ZN => n13815);
   U690 : NAND2_X1 port map( A1 => n371, A2 => n16578, ZN => n15538);
   U693 : XNOR2_X1 port map( A => n18466, B => n16037, ZN => n18401);
   U694 : NAND3_X2 port map( A1 => n10920, A2 => n10921, A3 => n3182, ZN => 
                           n12388);
   U699 : NAND2_X1 port map( A1 => n122, A2 => n121, ZN => n120);
   U700 : INV_X1 port map( A => n6802, ZN => n121);
   U701 : INV_X1 port map( A => n24772, ZN => n122);
   U702 : OAI21_X1 port map( B1 => n12537, B2 => n14271, A => n123, ZN => n2774
                           );
   U703 : INV_X1 port map( A => n13839, ZN => n123);
   U704 : NAND2_X1 port map( A1 => n9633, A2 => n9635, ZN => n10039);
   U705 : XNOR2_X2 port map( A => n8870, B => n8871, ZN => n9635);
   U706 : NOR2_X2 port map( A1 => n13007, A2 => n13008, ZN => n13830);
   U711 : INV_X1 port map( A => n6826, ZN => n6100);
   U712 : NAND2_X1 port map( A1 => n6602, A2 => n7013, ZN => n6826);
   U714 : NAND3_X2 port map( A1 => n6227, A2 => n6228, A3 => n6229, ZN => n7733
                           );
   U716 : NAND2_X1 port map( A1 => n14308, A2 => n14307, ZN => n13956);
   U718 : NAND2_X1 port map( A1 => n4249, A2 => n16002, ZN => n994);
   U719 : NAND2_X1 port map( A1 => n16004, A2 => n25009, ZN => n4249);
   U723 : OR2_X1 port map( A1 => n24470, A2 => n10935, ZN => n10509);
   U724 : BUF_X1 port map( A => n16431, Z => n17174);
   U725 : OAI21_X1 port map( B1 => n7100, B2 => n126, A => n125, ZN => n7105);
   U726 : NAND2_X1 port map( A1 => n7103, A2 => n127, ZN => n125);
   U727 : INV_X1 port map( A => n7101, ZN => n127);
   U729 : OR2_X2 port map( A1 => n6131, A2 => n128, ZN => n7615);
   U730 : AOI21_X1 port map( B1 => n6129, B2 => n6260, A => n6259, ZN => n128);
   U733 : NAND2_X1 port map( A1 => n6608, A2 => n6712, ZN => n1925);
   U735 : AND2_X2 port map( A1 => n727, A2 => n728, ZN => n20319);
   U737 : NAND2_X1 port map( A1 => n16126, A2 => n24458, ZN => n129);
   U743 : NAND2_X1 port map( A1 => n133, A2 => n24429, ZN => n17156);
   U745 : NAND2_X1 port map( A1 => n16046, A2 => n16045, ZN => n133);
   U747 : NAND2_X1 port map( A1 => n135, A2 => n24093, ZN => n10375);
   U751 : NAND3_X1 port map( A1 => n431, A2 => n7476, A3 => n7477, ZN => n7425)
                           ;
   U756 : OR2_X1 port map( A1 => n1147, A2 => n6976, ZN => n6388);
   U757 : XNOR2_X2 port map( A => n5829, B => Key(134), ZN => n6358);
   U759 : NAND2_X1 port map( A1 => n7185, A2 => n1862, ZN => n7246);
   U760 : NAND3_X2 port map( A1 => n2308, A2 => n2310, A3 => n2307, ZN => 
                           n11749);
   U763 : NAND2_X2 port map( A1 => n12732, A2 => n137, ZN => n14510);
   U765 : OR2_X2 port map( A1 => n16541, A2 => n16542, ZN => n18659);
   U767 : AOI22_X1 port map( A1 => n15945, A2 => n15943, B1 => n16443, B2 => 
                           n16440, ZN => n138);
   U768 : MUX2_X2 port map( A => n9768, B => n9767, S => n11163, Z => n12002);
   U770 : OAI21_X1 port map( B1 => n17443, B2 => n17444, A => n139, ZN => 
                           n17448);
   U772 : NAND2_X1 port map( A1 => n6904, A2 => n6902, ZN => n6903);
   U774 : NAND2_X2 port map( A1 => n4813, A2 => n4811, ZN => n8867);
   U777 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => n23414);
   U778 : OAI21_X1 port map( B1 => n23411, B2 => n24426, A => n23420, ZN => 
                           n140);
   U779 : NAND2_X1 port map( A1 => n23413, A2 => n142, ZN => n141);
   U781 : NAND2_X1 port map( A1 => n7103, A2 => n6165, ZN => n7098);
   U782 : NAND2_X1 port map( A1 => n1611, A2 => n4819, ZN => n2144);
   U784 : NAND3_X1 port map( A1 => n4326, A2 => n11499, A3 => n11058, ZN => 
                           n2152);
   U790 : NAND2_X1 port map( A1 => n19380, A2 => n24335, ZN => n19379);
   U791 : OR2_X1 port map( A1 => n25035, A2 => n23411, ZN => n3157);
   U796 : XNOR2_X1 port map( A => n144, B => n4153, ZN => Ciphertext(88));
   U797 : NAND2_X1 port map( A1 => n3156, A2 => n23414, ZN => n144);
   U798 : NAND3_X1 port map( A1 => n145, A2 => n2435, A3 => n10301, ZN => n2433
                           );
   U799 : NAND2_X1 port map( A1 => n2386, A2 => n10302, ZN => n145);
   U800 : NAND2_X1 port map( A1 => n7133, A2 => n146, ZN => n1848);
   U801 : NAND2_X1 port map( A1 => n7132, A2 => n7598, ZN => n146);
   U802 : AOI21_X2 port map( B1 => n12590, B2 => n13350, A => n2481, ZN => 
                           n14064);
   U805 : NAND3_X1 port map( A1 => n17236, A2 => n17237, A3 => n3872, ZN => 
                           n17238);
   U806 : NAND2_X1 port map( A1 => n9858, A2 => n238, ZN => n9861);
   U810 : XNOR2_X1 port map( A => n147, B => n8539, ZN => n8540);
   U811 : XNOR2_X1 port map( A => n8891, B => n8538, ZN => n147);
   U813 : NOR2_X2 port map( A1 => n12812, A2 => n12813, ZN => n14325);
   U814 : NAND2_X1 port map( A1 => n4962, A2 => n4963, ZN => n12907);
   U817 : OR2_X1 port map( A1 => n5992, A2 => n25045, ZN => n7018);
   U818 : OAI22_X2 port map( A1 => n16436, A2 => n16863, B1 => n16435, B2 => 
                           n17171, ZN => n18335);
   U829 : NOR2_X2 port map( A1 => n9439, A2 => n9438, ZN => n12108);
   U830 : XNOR2_X1 port map( A => n149, B => n4873, ZN => n17606);
   U831 : XNOR2_X1 port map( A => n18183, B => n18579, ZN => n149);
   U832 : BUF_X1 port map( A => n9944, Z => n9897);
   U834 : BUF_X1 port map( A => n5794, Z => n6623);
   U837 : OR2_X2 port map( A1 => n12887, A2 => n12888, ZN => n14153);
   U838 : INV_X1 port map( A => n17027, ZN => n17023);
   U839 : NAND2_X1 port map( A1 => n17391, A2 => n17185, ZN => n17027);
   U848 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => n151);
   U849 : NAND2_X1 port map( A1 => n15828, A2 => n1846, ZN => n152);
   U850 : NAND2_X1 port map( A1 => n15829, A2 => n15638, ZN => n153);
   U855 : NAND2_X1 port map( A1 => n14130, A2 => n4844, ZN => n13896);
   U856 : NAND2_X2 port map( A1 => n1564, A2 => n3493, ZN => n14130);
   U861 : AND2_X2 port map( A1 => n10675, A2 => n10673, ZN => n10985);
   U862 : OAI211_X2 port map( C1 => n14058, C2 => n14057, A => n2756, B => n155
                           , ZN => n15119);
   U863 : NAND2_X1 port map( A1 => n14056, A2 => n14058, ZN => n155);
   U864 : NAND2_X1 port map( A1 => n5863, A2 => n24592, ZN => n6260);
   U867 : NAND2_X1 port map( A1 => n3529, A2 => n3530, ZN => n156);
   U868 : NAND3_X1 port map( A1 => n7209, A2 => n7210, A3 => n2875, ZN => n9769
                           );
   U869 : NAND2_X1 port map( A1 => n17181, A2 => n15907, ZN => n15645);
   U874 : XNOR2_X2 port map( A => n14095, B => n14094, ZN => n16368);
   U875 : NAND2_X1 port map( A1 => n158, A2 => n23058, ZN => n22644);
   U876 : INV_X1 port map( A => n1322, ZN => n158);
   U877 : NAND2_X1 port map( A1 => n322, A2 => n23040, ZN => n1322);
   U879 : OR2_X2 port map( A1 => n5611, A2 => n5610, ZN => n24012);
   U881 : NOR2_X1 port map( A1 => n159, A2 => n23985, ZN => n23986);
   U882 : NAND2_X1 port map( A1 => n4476, A2 => n23984, ZN => n159);
   U883 : OAI21_X1 port map( B1 => n17067, B2 => n17069, A => n369, ZN => n723)
                           ;
   U886 : NAND2_X1 port map( A1 => n19646, A2 => n20343, ZN => n19648);
   U887 : NAND3_X1 port map( A1 => n160, A2 => n19104, A3 => n1706, ZN => 
                           n20518);
   U889 : NAND2_X1 port map( A1 => n15771, A2 => n161, ZN => n15770);
   U890 : NAND2_X1 port map( A1 => n162, A2 => n6307, ZN => n7863);
   U891 : NAND2_X1 port map( A1 => n909, A2 => n908, ZN => n162);
   U893 : NAND3_X2 port map( A1 => n15732, A2 => n15731, A3 => n468, ZN => 
                           n18382);
   U896 : NAND2_X1 port map( A1 => n24570, A2 => n17052, ZN => n3434);
   U898 : OAI211_X2 port map( C1 => n3921, C2 => n24257, A => n3924, B => n3920
                           , ZN => n7380);
   U899 : NAND2_X2 port map( A1 => n4858, A2 => n3494, ZN => n17131);
   U900 : NAND2_X1 port map( A1 => n5162, A2 => n7237, ZN => n4020);
   U906 : AND2_X2 port map( A1 => n5197, A2 => n5199, ZN => n10935);
   U907 : XNOR2_X1 port map( A => n15404, B => n164, ZN => n15406);
   U908 : XNOR2_X1 port map( A => n15402, B => n15401, ZN => n164);
   U916 : NAND3_X1 port map( A1 => n3429, A2 => n1582, A3 => n1581, ZN => n1580
                           );
   U920 : INV_X1 port map( A => n22988, ZN => n22992);
   U929 : AND3_X2 port map( A1 => n1881, A2 => n2956, A3 => n20091, ZN => 
                           n21182);
   U932 : MUX2_X1 port map( A => n5427, B => n20498, S => n19824, Z => n19828);
   U933 : NAND2_X1 port map( A1 => n20268, A2 => n1155, ZN => n19824);
   U935 : NAND2_X1 port map( A1 => n17211, A2 => n24529, ZN => n16880);
   U942 : NAND2_X1 port map( A1 => n20227, A2 => n20498, ZN => n171);
   U943 : NAND2_X1 port map( A1 => n172, A2 => n19082, ZN => n20501);
   U944 : NAND2_X1 port map( A1 => n5006, A2 => n5007, ZN => n172);
   U945 : NAND2_X1 port map( A1 => n17068, A2 => n1139, ZN => n16732);
   U949 : INV_X1 port map( A => n20249, ZN => n174);
   U950 : NAND2_X1 port map( A1 => n19788, A2 => n20241, ZN => n20248);
   U953 : NAND2_X1 port map( A1 => n175, A2 => n5518, ZN => n5517);
   U954 : NAND2_X1 port map( A1 => n787, A2 => n1534, ZN => n175);
   U959 : NAND2_X1 port map( A1 => n13722, A2 => n391, ZN => n4650);
   U967 : AND2_X2 port map( A1 => n2147, A2 => n2146, ZN => n7908);
   U974 : NAND2_X1 port map( A1 => n20383, A2 => n20459, ZN => n20464);
   U977 : MUX2_X2 port map( A => n19716, B => n19715, S => n19714, Z => n21506)
                           ;
   U978 : OR2_X2 port map( A1 => n6626, A2 => n6627, ZN => n7789);
   U979 : NOR2_X2 port map( A1 => n11075, A2 => n11074, ZN => n12196);
   U981 : NAND2_X1 port map( A1 => n2682, A2 => n4765, ZN => n178);
   U982 : NAND2_X1 port map( A1 => n363, A2 => n19191, ZN => n19566);
   U983 : OAI21_X1 port map( B1 => n20312, B2 => n20125, A => n179, ZN => 
                           n19967);
   U984 : NAND2_X1 port map( A1 => n20125, A2 => n20309, ZN => n179);
   U989 : XNOR2_X1 port map( A => n180, B => n20935, ZN => Ciphertext(152));
   U990 : NAND4_X1 port map( A1 => n4954, A2 => n5732, A3 => n4953, A4 => 
                           n21833, ZN => n180);
   U991 : NAND3_X1 port map( A1 => n11148, A2 => n11147, A3 => n11143, ZN => 
                           n10962);
   U992 : XNOR2_X1 port map( A => n181, B => n8936, ZN => n8939);
   U993 : XNOR2_X1 port map( A => n8937, B => n9188, ZN => n181);
   U995 : NOR2_X2 port map( A1 => n19800, A2 => n19801, ZN => n4227);
   U996 : NAND2_X1 port map( A1 => n17729, A2 => n16888, ZN => n17690);
   U997 : NAND2_X1 port map( A1 => n9683, A2 => n4069, ZN => n9686);
   U998 : NOR2_X1 port map( A1 => n260, A2 => n10044, ZN => n9683);
   U999 : NAND2_X1 port map( A1 => n19519, A2 => n19522, ZN => n19525);
   U1000 : INV_X1 port map( A => n7330, ZN => n5704);
   U1001 : NAND2_X1 port map( A1 => n3469, A2 => n7896, ZN => n7330);
   U1003 : AND2_X2 port map( A1 => n4726, A2 => n6197, ZN => n2624);
   U1005 : AOI21_X1 port map( B1 => n14231, B2 => n4560, A => n182, ZN => n4558
                           );
   U1010 : NAND2_X1 port map( A1 => n12428, A2 => n14315, ZN => n183);
   U1011 : NAND2_X1 port map( A1 => n12427, A2 => n14307, ZN => n185);
   U1013 : OR2_X2 port map( A1 => n7265, A2 => n7264, ZN => n8899);
   U1015 : OR2_X1 port map( A1 => n16809, A2 => n17081, ZN => n16590);
   U1016 : OR2_X1 port map( A1 => n19596, A2 => n18830, ZN => n19254);
   U1022 : NAND2_X1 port map( A1 => n1588, A2 => n22132, ZN => n22343);
   U1024 : NAND2_X1 port map( A1 => n3712, A2 => n16490, ZN => n15761);
   U1027 : NAND2_X1 port map( A1 => n23254, A2 => n189, ZN => n188);
   U1028 : INV_X1 port map( A => n23256, ZN => n189);
   U1031 : XNOR2_X2 port map( A => n14610, B => n14609, ZN => n16043);
   U1032 : OR3_X1 port map( A1 => n9985, A2 => n9980, A3 => n9981, ZN => n9739)
                           ;
   U1034 : BUF_X1 port map( A => n6275, Z => n6517);
   U1039 : NAND2_X1 port map( A1 => n17284, A2 => n17293, ZN => n17540);
   U1040 : NAND2_X2 port map( A1 => n2934, A2 => n2935, ZN => n17284);
   U1041 : AND3_X2 port map( A1 => n2698, A2 => n2697, A3 => n2696, ZN => 
                           n21084);
   U1042 : NAND3_X2 port map( A1 => n4339, A2 => n22332, A3 => n22331, ZN => 
                           n23165);
   U1043 : NAND2_X1 port map( A1 => n12710, A2 => n12707, ZN => n13074);
   U1047 : OAI21_X2 port map( B1 => n1373, B2 => n1406, A => n4252, ZN => 
                           n11057);
   U1048 : NAND3_X1 port map( A1 => n190, A2 => n6893, A3 => n6357, ZN => n730)
                           ;
   U1054 : NAND2_X1 port map( A1 => n14075, A2 => n396, ZN => n13851);
   U1059 : OAI21_X1 port map( B1 => n19387, B2 => n24477, A => n191, ZN => 
                           n2706);
   U1061 : NAND2_X1 port map( A1 => n10621, A2 => n10620, ZN => n10622);
   U1062 : NAND2_X1 port map( A1 => n232, A2 => n11212, ZN => n10621);
   U1066 : NOR2_X2 port map( A1 => n17200, A2 => n17201, ZN => n18290);
   U1069 : NAND3_X1 port map( A1 => n17572, A2 => n17042, A3 => n17573, ZN => 
                           n15995);
   U1071 : NAND2_X2 port map( A1 => n7455, A2 => n5161, ZN => n9041);
   U1075 : NAND3_X1 port map( A1 => n1861, A2 => n25366, A3 => n13345, ZN => 
                           n12575);
   U1082 : MUX2_X2 port map( A => n10418, B => n10417, S => n10416, Z => n11771
                           );
   U1087 : NAND2_X1 port map( A1 => n19404, A2 => n24929, ZN => n19189);
   U1088 : NAND2_X1 port map( A1 => n196, A2 => n194, ZN => n19040);
   U1090 : OAI21_X1 port map( B1 => n5233, B2 => n19036, A => n19037, ZN => 
                           n196);
   U1091 : AOI21_X2 port map( B1 => n15998, B2 => n15997, A => n15996, ZN => 
                           n18312);
   U1104 : NAND3_X1 port map( A1 => n197, A2 => n20508, A3 => n25223, ZN => 
                           n4328);
   U1105 : NAND4_X2 port map( A1 => n6691, A2 => n4828, A3 => n6689, A4 => 
                           n4829, ZN => n7413);
   U1106 : XNOR2_X1 port map( A => Key(6), B => Plaintext(6), ZN => n6434);
   U1107 : OR2_X1 port map( A1 => n11089, A2 => n11297, ZN => n1058);
   U1108 : OR2_X1 port map( A1 => n10451, A2 => n1499, ZN => n3443);
   U1111 : OR2_X1 port map( A1 => n13693, A2 => n13975, ZN => n14508);
   U1114 : OR2_X1 port map( A1 => n17343, A2 => n17241, ZN => n1284);
   U1116 : INV_X1 port map( A => n19485, ZN => n5280);
   U1119 : AND2_X1 port map( A1 => n23748, A2 => n997, ZN => n23744);
   U1120 : OR2_X1 port map( A1 => n22633, A2 => n2040, ZN => n509);
   U1121 : OR2_X1 port map( A1 => n22634, A2 => n509, ZN => n22640);
   U1122 : AND2_X1 port map( A1 => n6426, A2 => n6467, ZN => n198);
   U1123 : BUF_X1 port map( A => n6805, Z => n8530);
   U1124 : AND2_X1 port map( A1 => n7128, A2 => n7322, ZN => n199);
   U1125 : AND2_X1 port map( A1 => n20515, A2 => n20517, ZN => n200);
   U1128 : OR2_X1 port map( A1 => n10833, A2 => n9291, ZN => n201);
   U1130 : OR2_X1 port map( A1 => n10296, A2 => n5101, ZN => n202);
   U1132 : OR2_X1 port map( A1 => n10240, A2 => n10496, ZN => n203);
   U1133 : AND3_X1 port map( A1 => n11147, A2 => n11151, A3 => n714, ZN => n204
                           );
   U1135 : AND2_X2 port map( A1 => n10569, A2 => n10568, ZN => n13954);
   U1137 : OR2_X1 port map( A1 => n14002, A2 => n14003, ZN => n205);
   U1140 : OR3_X1 port map( A1 => n17322, A2 => n17321, A3 => n17320, ZN => 
                           n206);
   U1141 : OR2_X1 port map( A1 => n17323, A2 => n17324, ZN => n207);
   U1142 : OR3_X1 port map( A1 => n17332, A2 => n17335, A3 => n376, ZN => n208)
                           ;
   U1145 : AND2_X1 port map( A1 => n18764, A2 => n1475, ZN => n209);
   U1149 : OR2_X1 port map( A1 => n22456, A2 => n22270, ZN => n211);
   U1151 : OR3_X1 port map( A1 => n23839, A2 => n23857, A3 => n24469, ZN => 
                           n212);
   U1153 : OR2_X2 port map( A1 => n21871, A2 => n2921, ZN => n23317);
   U1155 : XNOR2_X1 port map( A => n14561, B => n14560, ZN => n16149);
   U1166 : XNOR2_X2 port map( A => n13199, B => n13198, ZN => n16597);
   U1168 : XNOR2_X2 port map( A => n8496, B => n8495, ZN => n9798);
   U1169 : XNOR2_X2 port map( A => n14878, B => n14877, ZN => n15921);
   U1182 : XNOR2_X2 port map( A => n5896, B => Key(53), ZN => n6560);
   U1188 : NOR2_X1 port map( A1 => n15617, A2 => n15616, ZN => n17062);
   U1190 : NOR2_X2 port map( A1 => n14037, A2 => n3891, ZN => n14846);
   U1198 : XNOR2_X1 port map( A => n8136, B => n8135, ZN => n9893);
   U1199 : AND2_X2 port map( A1 => n3045, A2 => n3044, ZN => n21591);
   U1211 : BUF_X1 port map( A => n11217, Z => n232);
   U1212 : OAI21_X1 port map( B1 => n5448, B2 => n10093, A => n10092, ZN => 
                           n11217);
   U1216 : NOR2_X1 port map( A1 => n11928, A2 => n11927, ZN => n14304);
   U1227 : XNOR2_X2 port map( A => n9093, B => n9094, ZN => n10060);
   U1229 : AND2_X2 port map( A1 => n6092, A2 => n6093, ZN => n5202);
   U1233 : OAI21_X2 port map( B1 => n8384, B2 => n9327, A => n8383, ZN => 
                           n10931);
   U1236 : OAI211_X2 port map( C1 => n7378, C2 => n7641, A => n2787, B => n7377
                           , ZN => n8517);
   U1244 : XNOR2_X1 port map( A => n8037, B => n5157, ZN => n9859);
   U1248 : XNOR2_X1 port map( A => n4385, B => n17652, ZN => n19485);
   U1256 : XNOR2_X2 port map( A => n11533, B => n11532, ZN => n12471);
   U1262 : XNOR2_X1 port map( A => n14412, B => n14411, ZN => n16428);
   U1264 : OR2_X1 port map( A1 => n19596, A2 => n25001, ZN => n808);
   U1272 : XNOR2_X1 port map( A => n8482, B => n8481, ZN => n9997);
   U1273 : OAI211_X2 port map( C1 => n7645, C2 => n7736, A => n7644, B => n7643
                           , ZN => n8898);
   U1275 : XNOR2_X2 port map( A => Key(183), B => Plaintext(183), ZN => n6438);
   U1279 : AOI21_X2 port map( B1 => n5814, B2 => n6242, A => n5813, ZN => n7577
                           );
   U1281 : XNOR2_X1 port map( A => n6000, B => Key(116), ZN => n6849);
   U1289 : XNOR2_X2 port map( A => n8750, B => n8749, ZN => n9762);
   U1297 : XNOR2_X2 port map( A => n4610, B => n4611, ZN => n3461);
   U1304 : BUF_X1 port map( A => n9255, Z => n261);
   U1305 : OAI211_X1 port map( C1 => n1183, C2 => n9934, A => n1182, B => n9933
                           , ZN => n10245);
   U1310 : XNOR2_X2 port map( A => n5943, B => Key(182), ZN => n6174);
   U1314 : XNOR2_X1 port map( A => n21056, B => n21057, ZN => n22244);
   U1316 : NOR2_X1 port map( A1 => n19510, A2 => n1419, ZN => n20249);
   U1319 : INV_X1 port map( A => n19310, ZN => n264);
   U1322 : NOR3_X1 port map( A1 => n17576, A2 => n1638, A3 => n1637, ZN => 
                           n17772);
   U1327 : INV_X1 port map( A => n17352, ZN => n266);
   U1328 : INV_X1 port map( A => n16333, ZN => n267);
   U1332 : INV_X1 port map( A => n10552, ZN => n11160);
   U1334 : INV_X1 port map( A => n7591, ZN => n268);
   U1336 : INV_X1 port map( A => n7965, ZN => n270);
   U1337 : OR2_X1 port map( A1 => n6174, A2 => n4866, ZN => n6334);
   U1338 : INV_X1 port map( A => n5804, ZN => n271);
   U1340 : CLKBUF_X1 port map( A => Key(83), Z => n2120);
   U1341 : CLKBUF_X1 port map( A => Key(11), Z => n1856);
   U1343 : CLKBUF_X1 port map( A => Key(124), Z => n765);
   U1344 : CLKBUF_X1 port map( A => Key(18), Z => n1833);
   U1345 : CLKBUF_X1 port map( A => Key(92), Z => n3183);
   U1347 : CLKBUF_X1 port map( A => Key(108), Z => n2834);
   U1349 : CLKBUF_X1 port map( A => Key(24), Z => n1865);
   U1351 : CLKBUF_X1 port map( A => Key(59), Z => n22886);
   U1353 : CLKBUF_X1 port map( A => Key(56), Z => n23679);
   U1354 : CLKBUF_X1 port map( A => Key(144), Z => n1952);
   U1355 : CLKBUF_X1 port map( A => Key(154), Z => n2744);
   U1356 : NOR2_X1 port map( A1 => n24492, A2 => n23361, ZN => n937);
   U1357 : INV_X1 port map( A => n22395, ZN => n23292);
   U1359 : AND2_X1 port map( A1 => n5223, A2 => n5222, ZN => n23227);
   U1360 : OAI21_X1 port map( B1 => n22503, B2 => n22504, A => n22502, ZN => 
                           n23442);
   U1363 : OAI211_X1 port map( C1 => n22393, C2 => n22958, A => n2857, B => 
                           n1889, ZN => n22395);
   U1364 : OAI21_X1 port map( B1 => n22966, B2 => n334, A => n833, ZN => n22970
                           );
   U1365 : OAI21_X1 port map( B1 => n335, B2 => n810, A => n809, ZN => n21842);
   U1370 : OAI21_X1 port map( B1 => n330, B2 => n25414, A => n520, ZN => n3642)
                           ;
   U1371 : XNOR2_X1 port map( A => n20002, B => n21083, ZN => n22228);
   U1375 : XNOR2_X1 port map( A => n20731, B => n20730, ZN => n22323);
   U1377 : INV_X1 port map( A => n22449, ZN => n274);
   U1378 : XNOR2_X1 port map( A => n3871, B => n20252, ZN => n22354);
   U1386 : OAI21_X1 port map( B1 => n343, B2 => n20269, A => n1154, ZN => 
                           n19091);
   U1387 : OAI21_X1 port map( B1 => n1256, B2 => n345, A => n1255, ZN => n20876
                           );
   U1389 : OR2_X1 port map( A1 => n20051, A2 => n2168, ZN => n1072);
   U1390 : AND2_X1 port map( A1 => n20338, A2 => n20666, ZN => n19710);
   U1393 : INV_X1 port map( A => n19875, ZN => n275);
   U1397 : AND2_X1 port map( A1 => n348, A2 => n20479, ZN => n1023);
   U1398 : INV_X1 port map( A => n20370, ZN => n277);
   U1401 : OR2_X1 port map( A1 => n4075, A2 => n18927, ZN => n17942);
   U1403 : OR2_X1 port map( A1 => n19613, A2 => n355, ZN => n1805);
   U1404 : OR2_X1 port map( A1 => n19360, A2 => n18817, ZN => n1265);
   U1405 : AND2_X1 port map( A1 => n19565, A2 => n19191, ZN => n1051);
   U1406 : AND2_X1 port map( A1 => n363, A2 => n19570, ZN => n1049);
   U1408 : INV_X1 port map( A => n355, ZN => n278);
   U1409 : XNOR2_X1 port map( A => n18282, B => n3753, ZN => n3773);
   U1410 : XNOR2_X1 port map( A => n18479, B => n18480, ZN => n19575);
   U1412 : INV_X1 port map( A => n19543, ZN => n279);
   U1414 : XNOR2_X1 port map( A => n18321, B => n18322, ZN => n19568);
   U1417 : XNOR2_X1 port map( A => n17922, B => n17923, ZN => n4748);
   U1418 : XNOR2_X1 port map( A => n17819, B => n444, ZN => n17820);
   U1419 : XNOR2_X1 port map( A => n25390, B => n450, ZN => n17360);
   U1424 : AOI21_X1 port map( B1 => n17143, B2 => n368, A => n17146, ZN => n474
                           );
   U1425 : AOI22_X1 port map( A1 => n16560, A2 => n17408, B1 => n17613, B2 => 
                           n17409, ZN => n16563);
   U1426 : OAI211_X1 port map( C1 => n366, C2 => n17473, A => n17474, B => 
                           n17475, ZN => n515);
   U1428 : AND2_X1 port map( A1 => n17044, A2 => n373, ZN => n16767);
   U1429 : INV_X1 port map( A => n4004, ZN => n281);
   U1430 : CLKBUF_X1 port map( A => n16527, Z => n17453);
   U1431 : INV_X1 port map( A => n17173, ZN => n282);
   U1432 : BUF_X1 port map( A => n16660, Z => n17031);
   U1433 : INV_X1 port map( A => n1139, ZN => n283);
   U1435 : INV_X1 port map( A => n17053, ZN => n284);
   U1437 : INV_X1 port map( A => n17400, ZN => n285);
   U1440 : NAND2_X1 port map( A1 => n15835, A2 => n15836, ZN => n16888);
   U1442 : BUF_X1 port map( A => n17065, Z => n369);
   U1449 : INV_X1 port map( A => n17461, ZN => n287);
   U1451 : INV_X1 port map( A => n15560, ZN => n16023);
   U1455 : CLKBUF_X1 port map( A => n15710, Z => n16438);
   U1458 : INV_X1 port map( A => n16334, ZN => n290);
   U1459 : INV_X1 port map( A => n16042, ZN => n291);
   U1463 : XNOR2_X1 port map( A => n14723, B => n14722, ZN => n15584);
   U1464 : INV_X1 port map( A => n16149, ZN => n293);
   U1465 : XNOR2_X1 port map( A => n13499, B => n13498, ZN => n16332);
   U1466 : XNOR2_X1 port map( A => n14969, B => n14968, ZN => n16451);
   U1468 : XNOR2_X1 port map( A => n14979, B => n14919, ZN => n1091);
   U1471 : INV_X1 port map( A => n14997, ZN => n295);
   U1472 : OAI21_X1 port map( B1 => n14123, B2 => n14208, A => n2214, ZN => 
                           n14210);
   U1473 : AND2_X1 port map( A1 => n394, A2 => n13951, ZN => n749);
   U1474 : INV_X1 port map( A => n4844, ZN => n14132);
   U1475 : INV_X1 port map( A => n14034, ZN => n296);
   U1476 : INV_X1 port map( A => n14149, ZN => n297);
   U1477 : INV_X1 port map( A => n14044, ZN => n298);
   U1478 : INV_X1 port map( A => n13488, ZN => n299);
   U1480 : NAND3_X1 port map( A1 => n12422, A2 => n1086, A3 => n1087, ZN => 
                           n13900);
   U1483 : INV_X1 port map( A => n13847, ZN => n300);
   U1485 : OR2_X1 port map( A1 => n12483, A2 => n12715, ZN => n4057);
   U1487 : INV_X1 port map( A => n13328, ZN => n301);
   U1488 : XNOR2_X1 port map( A => n12044, B => n12043, ZN => n2295);
   U1489 : OR2_X1 port map( A1 => n13056, A2 => n13057, ZN => n11438);
   U1491 : INV_X1 port map( A => n12784, ZN => n302);
   U1492 : INV_X1 port map( A => n12796, ZN => n303);
   U1493 : XNOR2_X1 port map( A => n12290, B => n12289, ZN => n13114);
   U1496 : INV_X1 port map( A => n4766, ZN => n304);
   U1499 : XNOR2_X1 port map( A => n11977, B => n11295, ZN => n12114);
   U1504 : OR2_X1 port map( A1 => n11101, A2 => n10914, ZN => n10220);
   U1506 : NOR2_X1 port map( A1 => n11342, A2 => n10632, ZN => n10491);
   U1507 : AND2_X1 port map( A1 => n10891, A2 => n10889, ZN => n10438);
   U1511 : INV_X1 port map( A => n11122, ZN => n305);
   U1518 : XNOR2_X1 port map( A => n7550, B => n7549, ZN => n9281);
   U1519 : INV_X1 port map( A => n1595, ZN => n3292);
   U1523 : INV_X1 port map( A => n10061, ZN => n309);
   U1524 : XNOR2_X1 port map( A => n9105, B => n9104, ZN => n9127);
   U1526 : INV_X1 port map( A => n8818, ZN => n310);
   U1530 : OR2_X1 port map( A1 => n8008, A2 => n8007, ZN => n8970);
   U1531 : AND4_X1 port map( A1 => n1195, A2 => n1190, A3 => n1191, A4 => n1193
                           , ZN => n1110);
   U1532 : BUF_X1 port map( A => n7108, Z => n7532);
   U1534 : INV_X1 port map( A => n7609, ZN => n311);
   U1535 : BUF_X1 port map( A => n7589, Z => n7462);
   U1536 : CLKBUF_X1 port map( A => n7409, Z => n7982);
   U1540 : INV_X1 port map( A => n7917, ZN => n312);
   U1543 : INV_X1 port map( A => n1147, ZN => n6687);
   U1545 : CLKBUF_X1 port map( A => n6066, Z => n6688);
   U1548 : XNOR2_X1 port map( A => n5803, B => Key(67), ZN => n5804);
   U1549 : CLKBUF_X1 port map( A => n6400, Z => n6755);
   U1550 : CLKBUF_X1 port map( A => n6648, Z => n7011);
   U1552 : INV_X1 port map( A => n6358, ZN => n313);
   U1555 : CLKBUF_X1 port map( A => Key(109), Z => n925);
   U1556 : CLKBUF_X1 port map( A => Key(81), Z => n3062);
   U1557 : CLKBUF_X1 port map( A => Key(110), Z => n2049);
   U1558 : CLKBUF_X1 port map( A => Key(67), Z => n494);
   U1559 : CLKBUF_X1 port map( A => Key(126), Z => n1745);
   U1560 : CLKBUF_X1 port map( A => Key(123), Z => n21662);
   U1562 : CLKBUF_X1 port map( A => Key(177), Z => n20284);
   U1563 : CLKBUF_X1 port map( A => Key(170), Z => n1777);
   U1565 : CLKBUF_X1 port map( A => Key(31), Z => n2726);
   U1568 : CLKBUF_X1 port map( A => Key(128), Z => n2746);
   U1569 : CLKBUF_X1 port map( A => Key(125), Z => n2881);
   U1570 : CLKBUF_X1 port map( A => Key(88), Z => n891);
   U1572 : CLKBUF_X1 port map( A => Key(133), Z => n2826);
   U1573 : CLKBUF_X1 port map( A => Key(9), Z => n19392);
   U1574 : CLKBUF_X1 port map( A => Key(114), Z => n2211);
   U1575 : CLKBUF_X1 port map( A => Key(7), Z => n2222);
   U1576 : CLKBUF_X1 port map( A => Key(121), Z => n2145);
   U1577 : CLKBUF_X1 port map( A => Key(165), Z => n924);
   U1578 : CLKBUF_X1 port map( A => Key(21), Z => n17960);
   U1579 : CLKBUF_X1 port map( A => Key(160), Z => n1754);
   U1580 : CLKBUF_X1 port map( A => Key(135), Z => n3129);
   U1582 : CLKBUF_X1 port map( A => Key(129), Z => n876);
   U1584 : CLKBUF_X1 port map( A => Key(77), Z => n681);
   U1585 : CLKBUF_X1 port map( A => Key(118), Z => n3118);
   U1586 : CLKBUF_X1 port map( A => Key(104), Z => n3089);
   U1587 : CLKBUF_X1 port map( A => Key(130), Z => n2739);
   U1588 : CLKBUF_X1 port map( A => Key(70), Z => n663);
   U1589 : CLKBUF_X1 port map( A => Key(112), Z => n2126);
   U1590 : CLKBUF_X1 port map( A => Key(1), Z => n2805);
   U1591 : CLKBUF_X1 port map( A => Key(42), Z => n2761);
   U1592 : CLKBUF_X1 port map( A => Key(171), Z => n20690);
   U1593 : CLKBUF_X1 port map( A => Key(49), Z => n1827);
   U1594 : CLKBUF_X1 port map( A => Key(143), Z => n20609);
   U1596 : CLKBUF_X1 port map( A => Key(178), Z => n896);
   U1598 : CLKBUF_X1 port map( A => Key(39), Z => n2039);
   U1599 : CLKBUF_X1 port map( A => Key(17), Z => n1869);
   U1602 : CLKBUF_X1 port map( A => Key(52), Z => n1746);
   U1603 : CLKBUF_X1 port map( A => Key(22), Z => n1797);
   U1604 : CLKBUF_X1 port map( A => Key(95), Z => n14398);
   U1606 : CLKBUF_X1 port map( A => Key(147), Z => n1724);
   U1610 : CLKBUF_X1 port map( A => Key(16), Z => n853);
   U1611 : CLKBUF_X1 port map( A => Key(163), Z => n1757);
   U1613 : CLKBUF_X1 port map( A => Key(111), Z => n21204);
   U1615 : CLKBUF_X1 port map( A => Key(141), Z => n1804);
   U1616 : CLKBUF_X1 port map( A => Key(103), Z => n1951);
   U1617 : CLKBUF_X1 port map( A => Key(148), Z => n812);
   U1618 : CLKBUF_X1 port map( A => Key(120), Z => n3084);
   U1619 : CLKBUF_X1 port map( A => Key(127), Z => n1815);
   U1620 : CLKBUF_X1 port map( A => Key(76), Z => n2772);
   U1622 : CLKBUF_X1 port map( A => Key(71), Z => n2240);
   U1623 : CLKBUF_X1 port map( A => Key(85), Z => n2241);
   U1624 : CLKBUF_X1 port map( A => Key(69), Z => n860);
   U1625 : CLKBUF_X1 port map( A => Key(62), Z => n1863);
   U1626 : CLKBUF_X1 port map( A => Key(55), Z => n1739);
   U1627 : CLKBUF_X1 port map( A => Key(5), Z => n2991);
   U1628 : CLKBUF_X1 port map( A => Key(84), Z => n2193);
   U1629 : CLKBUF_X1 port map( A => Key(173), Z => n3158);
   U1630 : CLKBUF_X1 port map( A => Key(159), Z => n2044);
   U1631 : CLKBUF_X1 port map( A => Key(145), Z => n1792);
   U1632 : CLKBUF_X1 port map( A => Key(19), Z => n1835);
   U1634 : CLKBUF_X1 port map( A => Key(138), Z => n1801);
   U1635 : CLKBUF_X1 port map( A => Key(96), Z => n2717);
   U1636 : CLKBUF_X1 port map( A => Key(180), Z => n912);
   U1637 : CLKBUF_X1 port map( A => Key(47), Z => n889);
   U1639 : CLKBUF_X1 port map( A => Key(155), Z => n2989);
   U1640 : INV_X1 port map( A => n6521, ZN => n315);
   U1641 : CLKBUF_X1 port map( A => Key(75), Z => n2882);
   U1642 : CLKBUF_X1 port map( A => Key(169), Z => n899);
   U1644 : CLKBUF_X1 port map( A => Key(162), Z => n921);
   U1645 : CLKBUF_X1 port map( A => Key(153), Z => n1891);
   U1646 : CLKBUF_X1 port map( A => Key(139), Z => n1810);
   U1648 : CLKBUF_X1 port map( A => Key(191), Z => n2847);
   U1649 : INV_X1 port map( A => n6243, ZN => n316);
   U1650 : CLKBUF_X1 port map( A => Key(34), Z => n1789);
   U1651 : CLKBUF_X1 port map( A => Key(6), Z => n21623);
   U1652 : CLKBUF_X1 port map( A => Key(27), Z => n763);
   U1653 : CLKBUF_X1 port map( A => Key(188), Z => n3131);
   U1654 : CLKBUF_X1 port map( A => Key(10), Z => n20995);
   U1655 : CLKBUF_X1 port map( A => Key(181), Z => n1767);
   U1658 : CLKBUF_X1 port map( A => Key(80), Z => n2236);
   U1659 : CLKBUF_X1 port map( A => Key(86), Z => n3178);
   U1660 : CLKBUF_X1 port map( A => Key(72), Z => n1758);
   U1661 : CLKBUF_X1 port map( A => Key(73), Z => n881);
   U1663 : CLKBUF_X1 port map( A => Key(65), Z => n20046);
   U1665 : CLKBUF_X1 port map( A => Key(51), Z => n2087);
   U1666 : CLKBUF_X1 port map( A => Key(66), Z => n2990);
   U1667 : CLKBUF_X1 port map( A => Key(12), Z => n2208);
   U1668 : CLKBUF_X1 port map( A => Key(87), Z => n1826);
   U1669 : CLKBUF_X1 port map( A => Key(23), Z => n2190);
   U1670 : CLKBUF_X1 port map( A => Key(36), Z => n1364);
   U1671 : CLKBUF_X1 port map( A => Key(78), Z => n1924);
   U1672 : CLKBUF_X1 port map( A => Key(43), Z => n1768);
   U1673 : CLKBUF_X1 port map( A => Key(50), Z => n2005);
   U1674 : NOR2_X1 port map( A1 => n23511, A2 => n23512, ZN => n23522);
   U1675 : OAI211_X1 port map( C1 => n23965, C2 => n23964, A => n23963, B => 
                           n878, ZN => n3150);
   U1676 : OR2_X1 port map( A1 => n23728, A2 => n23727, ZN => n786);
   U1677 : OR2_X1 port map( A1 => n22531, A2 => n22532, ZN => n852);
   U1678 : OR2_X1 port map( A1 => n23692, A2 => n23689, ZN => n1145);
   U1679 : NOR2_X1 port map( A1 => n23619, A2 => n23634, ZN => n23652);
   U1680 : NOR2_X1 port map( A1 => n23292, A2 => n23303, ZN => n23298);
   U1682 : INV_X1 port map( A => n23311, ZN => n4108);
   U1683 : AND2_X1 port map( A1 => n23911, A2 => n23924, ZN => n23941);
   U1687 : AND2_X1 port map( A1 => n1683, A2 => n1686, ZN => n23327);
   U1694 : BUF_X1 port map( A => n24010, Z => n23982);
   U1696 : OAI21_X1 port map( B1 => n21378, B2 => n25543, A => n5048, ZN => 
                           n22442);
   U1699 : INV_X1 port map( A => n23227, ZN => n317);
   U1701 : INV_X1 port map( A => n23810, ZN => n318);
   U1702 : AND3_X1 port map( A1 => n5422, A2 => n5419, A3 => n1397, ZN => 
                           n23361);
   U1703 : INV_X1 port map( A => n21863, ZN => n23903);
   U1705 : OAI21_X1 port map( B1 => n22497, B2 => n4719, A => n2364, ZN => 
                           n23443);
   U1711 : INV_X1 port map( A => n23442, ZN => n321);
   U1713 : INV_X1 port map( A => n22698, ZN => n322);
   U1714 : INV_X1 port map( A => n23972, ZN => n878);
   U1716 : AND3_X1 port map( A1 => n4781, A2 => n1691, A3 => n22729, ZN => 
                           n23517);
   U1719 : OAI21_X1 port map( B1 => n4591, B2 => n22408, A => n24951, ZN => 
                           n22414);
   U1720 : INV_X1 port map( A => n23543, ZN => n323);
   U1723 : OAI21_X1 port map( B1 => n20980, B2 => n20979, A => n24902, ZN => 
                           n1007);
   U1725 : AND2_X1 port map( A1 => n22808, A2 => n4427, ZN => n23993);
   U1726 : INV_X1 port map( A => n24879, ZN => n324);
   U1728 : OR2_X1 port map( A1 => n24951, A2 => n22565, ZN => n650);
   U1729 : OR2_X1 port map( A1 => n22953, A2 => n21878, ZN => n1257);
   U1730 : OR2_X1 port map( A1 => n22034, A2 => n24884, ZN => n1258);
   U1731 : AND2_X1 port map( A1 => n22667, A2 => n22670, ZN => n919);
   U1732 : INV_X1 port map( A => n22219, ZN => n22217);
   U1733 : OR2_X1 port map( A1 => n4468, A2 => n4467, ZN => n481);
   U1734 : INV_X1 port map( A => n3781, ZN => n1686);
   U1736 : OR2_X1 port map( A1 => n22322, A2 => n22456, ZN => n22327);
   U1737 : NOR2_X1 port map( A1 => n21802, A2 => n22198, ZN => n23634);
   U1738 : INV_X1 port map( A => n22356, ZN => n21348);
   U1741 : AND2_X1 port map( A1 => n25082, A2 => n22361, ZN => n1249);
   U1742 : OR2_X1 port map( A1 => n21841, A2 => n22257, ZN => n810);
   U1744 : OR2_X1 port map( A1 => n22426, A2 => n2674, ZN => n776);
   U1745 : XNOR2_X1 port map( A => n20783, B => n20782, ZN => n5084);
   U1746 : XNOR2_X1 port map( A => n20746, B => n20745, ZN => n22454);
   U1747 : OR2_X1 port map( A1 => n21856, A2 => n22769, ZN => n534);
   U1749 : OR2_X1 port map( A1 => n21792, A2 => n3231, ZN => n1163);
   U1751 : OR2_X1 port map( A1 => n22261, A2 => n22398, ZN => n22262);
   U1752 : INV_X1 port map( A => n2601, ZN => n1146);
   U1753 : OR2_X1 port map( A1 => n22056, A2 => n21836, ZN => n1310);
   U1757 : CLKBUF_X1 port map( A => n21766, Z => n22206);
   U1758 : INV_X1 port map( A => n22953, ZN => n1293);
   U1759 : INV_X1 port map( A => n23574, ZN => n325);
   U1760 : INV_X1 port map( A => n24971, ZN => n326);
   U1761 : XNOR2_X1 port map( A => n21006, B => n21007, ZN => n22926);
   U1764 : AND2_X1 port map( A1 => n4273, A2 => n22655, ZN => n22811);
   U1766 : CLKBUF_X1 port map( A => n21265, Z => n22614);
   U1767 : INV_X1 port map( A => n22888, ZN => n327);
   U1769 : INV_X1 port map( A => n22228, ZN => n328);
   U1772 : CLKBUF_X1 port map( A => n21759, Z => n22197);
   U1773 : INV_X1 port map( A => n22323, ZN => n329);
   U1774 : XNOR2_X1 port map( A => n20083, B => n20082, ZN => n22355);
   U1777 : INV_X1 port map( A => n23999, ZN => n330);
   U1779 : XNOR2_X1 port map( A => n20988, B => n20987, ZN => n22715);
   U1780 : INV_X1 port map( A => n22657, ZN => n331);
   U1781 : INV_X1 port map( A => n22257, ZN => n332);
   U1782 : INV_X1 port map( A => n21934, ZN => n333);
   U1784 : INV_X1 port map( A => n22968, ZN => n334);
   U1785 : XNOR2_X1 port map( A => n21595, B => n21594, ZN => n22033);
   U1786 : XNOR2_X1 port map( A => n20642, B => n20643, ZN => n22333);
   U1790 : CLKBUF_X1 port map( A => n21209, Z => n20634);
   U1791 : INV_X1 port map( A => n22252, ZN => n335);
   U1792 : INV_X1 port map( A => n22222, ZN => n336);
   U1793 : XNOR2_X1 port map( A => n21180, B => n21179, ZN => n22448);
   U1794 : INV_X1 port map( A => n22832, ZN => n337);
   U1795 : INV_X1 port map( A => n22965, ZN => n338);
   U1796 : XNOR2_X1 port map( A => n21621, B => n21985, ZN => n20957);
   U1797 : XNOR2_X1 port map( A => n21176, B => n20594, ZN => n21562);
   U1798 : XNOR2_X1 port map( A => n1153, B => n20904, ZN => n21496);
   U1799 : XNOR2_X1 port map( A => n21569, B => n21402, ZN => n21246);
   U1800 : XNOR2_X1 port map( A => n21688, B => n596, ZN => n21690);
   U1802 : NAND3_X1 port map( A1 => n19048, A2 => n19050, A3 => n19049, ZN => 
                           n20870);
   U1803 : XNOR2_X1 port map( A => n21687, B => n21689, ZN => n596);
   U1814 : OAI21_X1 port map( B1 => n19706, B2 => n20614, A => n19705, ZN => 
                           n21975);
   U1815 : AND3_X1 port map( A1 => n4183, A2 => n20266, A3 => n20265, ZN => 
                           n4185);
   U1820 : MUX2_X1 port map( A => n21009, B => n24581, S => n20289, Z => n20295
                           );
   U1824 : OAI211_X1 port map( C1 => n19939, C2 => n24077, A => n3650, B => 
                           n19339, ZN => n21106);
   U1825 : OR2_X1 port map( A1 => n20592, A2 => n20593, ZN => n2362);
   U1826 : OAI21_X1 port map( B1 => n636, B2 => n20527, A => n20526, ZN => 
                           n21013);
   U1829 : NOR2_X1 port map( A1 => n20074, A2 => n19855, ZN => n588);
   U1831 : NAND2_X1 port map( A1 => n19938, A2 => n19939, ZN => n2946);
   U1832 : AND2_X1 port map( A1 => n20255, A2 => n19743, ZN => n1256);
   U1833 : INV_X1 port map( A => n19511, ZN => n754);
   U1834 : OR2_X1 port map( A1 => n24076, A2 => n20616, ZN => n19703);
   U1835 : AOI22_X1 port map( A1 => n20478, A2 => n1024, B1 => n1023, B2 => 
                           n20480, ZN => n1022);
   U1836 : INV_X1 port map( A => n20191, ZN => n1242);
   U1837 : INV_X1 port map( A => n19743, ZN => n2024);
   U1840 : INV_X1 port map( A => n19984, ZN => n885);
   U1842 : AND2_X1 port map( A1 => n20578, A2 => n20576, ZN => n1205);
   U1843 : OR2_X1 port map( A1 => n20165, A2 => n20395, ZN => n2426);
   U1844 : OR2_X1 port map( A1 => n1591, A2 => n17943, ZN => n21031);
   U1845 : INV_X1 port map( A => n17943, ZN => n21033);
   U1847 : INV_X1 port map( A => n20262, ZN => n20409);
   U1849 : INV_X1 port map( A => n19887, ZN => n339);
   U1850 : NAND2_X1 port map( A1 => n1716, A2 => n1421, ZN => n20094);
   U1851 : AND2_X1 port map( A1 => n20523, A2 => n20522, ZN => n21009);
   U1853 : NAND2_X1 port map( A1 => n1980, A2 => n18394, ZN => n20022);
   U1854 : OR2_X1 port map( A1 => n19619, A2 => n19618, ZN => n594);
   U1856 : INV_X1 port map( A => n20319, ZN => n340);
   U1857 : NOR2_X1 port map( A1 => n20142, A2 => n19975, ZN => n19680);
   U1858 : BUF_X1 port map( A => n19774, Z => n20384);
   U1859 : AND3_X1 port map( A1 => n4916, A2 => n2983, A3 => n4915, ZN => 
                           n17567);
   U1860 : NOR2_X1 port map( A1 => n20497, A2 => n20498, ZN => n20502);
   U1865 : NAND2_X1 port map( A1 => n18547, A2 => n3055, ZN => n20614);
   U1867 : INV_X1 port map( A => n20055, ZN => n19928);
   U1868 : INV_X1 port map( A => n20317, ZN => n341);
   U1869 : AOI21_X1 port map( B1 => n19529, B2 => n1013, A => n1011, ZN => 
                           n1010);
   U1871 : AND2_X1 port map( A1 => n3277, A2 => n3989, ZN => n818);
   U1873 : NAND2_X1 port map( A1 => n5646, A2 => n18827, ZN => n20476);
   U1876 : INV_X1 port map( A => n20498, ZN => n343);
   U1880 : INV_X1 port map( A => n20413, ZN => n345);
   U1883 : INV_X1 port map( A => n20214, ZN => n20199);
   U1886 : INV_X1 port map( A => n20909, ZN => n346);
   U1887 : OAI21_X1 port map( B1 => n1046, B2 => n1050, A => n1048, ZN => 
                           n20214);
   U1891 : INV_X1 port map( A => n20353, ZN => n348);
   U1892 : OR2_X1 port map( A1 => n17554, A2 => n19531, ZN => n1015);
   U1893 : NAND2_X1 port map( A1 => n19533, A2 => n19531, ZN => n1016);
   U1894 : INV_X1 port map( A => n20367, ZN => n349);
   U1895 : OR2_X1 port map( A1 => n18443, A2 => n19164, ZN => n1977);
   U1896 : AOI22_X1 port map( A1 => n1001, A2 => n280, B1 => n19576, B2 => 
                           n25072, ZN => n1000);
   U1897 : OAI21_X1 port map( B1 => n19629, B2 => n4543, A => n3379, ZN => 
                           n19840);
   U1898 : OR2_X1 port map( A1 => n1107, A2 => n264, ZN => n1160);
   U1899 : INV_X1 port map( A => n20460, ZN => n350);
   U1900 : INV_X1 port map( A => n20515, ZN => n351);
   U1901 : NOR2_X1 port map( A1 => n24982, A2 => n1002, ZN => n1001);
   U1902 : INV_X1 port map( A => n19007, ZN => n1005);
   U1903 : XNOR2_X1 port map( A => n4890, B => n18384, ZN => n18597);
   U1904 : AND2_X1 port map( A1 => n1052, A2 => n5634, ZN => n1050);
   U1905 : AND2_X1 port map( A1 => n1051, A2 => n1047, ZN => n1046);
   U1906 : AOI21_X1 port map( B1 => n19269, B2 => n19534, A => n4172, ZN => 
                           n1012);
   U1907 : NAND2_X1 port map( A1 => n1291, A2 => n19435, ZN => n1290);
   U1908 : OR2_X1 port map( A1 => n19435, A2 => n18833, ZN => n1287);
   U1909 : BUF_X1 port map( A => n18772, Z => n19125);
   U1912 : AND2_X1 port map( A1 => n18788, A2 => n19397, ZN => n18900);
   U1913 : NAND3_X1 port map( A1 => n19060, A2 => n19059, A3 => n19007, ZN => 
                           n19062);
   U1921 : AND2_X1 port map( A1 => n4436, A2 => n1300, ZN => n4435);
   U1922 : OR2_X1 port map( A1 => n19311, A2 => n19309, ZN => n696);
   U1923 : INV_X1 port map( A => n19186, ZN => n19404);
   U1924 : INV_X1 port map( A => n19421, ZN => n1306);
   U1925 : AND2_X1 port map( A1 => n19419, A2 => n19420, ZN => n1307);
   U1926 : AND2_X1 port map( A1 => n988, A2 => n24982, ZN => n1443);
   U1928 : XNOR2_X1 port map( A => n17647, B => n17646, ZN => n19490);
   U1931 : INV_X1 port map( A => n19487, ZN => n352);
   U1934 : INV_X1 port map( A => n3773, ZN => n353);
   U1935 : INV_X1 port map( A => n19575, ZN => n354);
   U1936 : INV_X1 port map( A => n19238, ZN => n355);
   U1938 : XNOR2_X1 port map( A => n17508, B => n17507, ZN => n19300);
   U1939 : INV_X1 port map( A => n19126, ZN => n19543);
   U1940 : INV_X1 port map( A => n19418, ZN => n19419);
   U1941 : INV_X1 port map( A => n19296, ZN => n356);
   U1942 : INV_X1 port map( A => n19502, ZN => n357);
   U1945 : XNOR2_X1 port map( A => n18427, B => n18426, ZN => n19162);
   U1947 : XNOR2_X1 port map( A => n16939, B => n16938, ZN => n19311);
   U1948 : INV_X1 port map( A => n19273, ZN => n1053);
   U1949 : XNOR2_X1 port map( A => n18625, B => n18624, ZN => n19441);
   U1950 : INV_X1 port map( A => n19500, ZN => n358);
   U1954 : INV_X1 port map( A => n19570, ZN => n960);
   U1955 : XNOR2_X1 port map( A => n18462, B => n18461, ZN => n988);
   U1957 : OR2_X1 port map( A1 => n19568, A2 => n19192, ZN => n1047);
   U1960 : XNOR2_X1 port map( A => n4274, B => n16626, ZN => n19559);
   U1962 : INV_X1 port map( A => n18832, ZN => n361);
   U1963 : XNOR2_X1 port map( A => n18273, B => n18274, ZN => n19126);
   U1964 : XNOR2_X1 port map( A => n18699, B => n18698, ZN => n19407);
   U1966 : XNOR2_X1 port map( A => n17308, B => n17307, ZN => n19329);
   U1969 : XNOR2_X1 port map( A => n18632, B => n18631, ZN => n19438);
   U1972 : XNOR2_X1 port map( A => n18379, B => n18378, ZN => n19428);
   U1973 : INV_X1 port map( A => n19568, ZN => n362);
   U1974 : INV_X1 port map( A => n19192, ZN => n363);
   U1975 : XNOR2_X1 port map( A => n17787, B => n17786, ZN => n19370);
   U1977 : XNOR2_X1 port map( A => n17874, B => n3725, ZN => n966);
   U1978 : XNOR2_X1 port map( A => n17638, B => n17637, ZN => n18051);
   U1980 : XNOR2_X1 port map( A => n18334, B => n18407, ZN => n17648);
   U1981 : XNOR2_X1 port map( A => n934, B => n25411, ZN => n18683);
   U1982 : AOI22_X1 port map( A1 => n4267, A2 => n4266, B1 => n16610, B2 => 
                           n17054, ZN => n17933);
   U1985 : XNOR2_X1 port map( A => n18674, B => n18295, ZN => n18387);
   U1992 : XNOR2_X1 port map( A => n17807, B => n17913, ZN => n18390);
   U1993 : OAI211_X1 port map( C1 => n17030, C2 => n16662, A => n4036, B => 
                           n4035, ZN => n17840);
   U1998 : OAI211_X1 port map( C1 => n3601, C2 => n3603, A => n3600, B => n3599
                           , ZN => n18541);
   U2001 : AND2_X1 port map( A1 => n3260, A2 => n16968, ZN => n17662);
   U2002 : NAND2_X1 port map( A1 => n15882, A2 => n935, ZN => n934);
   U2003 : INV_X1 port map( A => n15610, ZN => n1135);
   U2004 : AND2_X1 port map( A1 => n2133, A2 => n2134, ZN => n1253);
   U2008 : NAND2_X1 port map( A1 => n16679, A2 => n5521, ZN => n17807);
   U2009 : NAND3_X1 port map( A1 => n1269, A2 => n15635, A3 => n15636, ZN => 
                           n17875);
   U2010 : OAI211_X1 port map( C1 => n2429, C2 => n17483, A => n17480, B => 
                           n2428, ZN => n18365);
   U2012 : OAI21_X1 port map( B1 => n17027, B2 => n3598, A => n17026, ZN => 
                           n18096);
   U2014 : AND2_X1 port map( A1 => n17084, A2 => n16581, ZN => n575);
   U2015 : OR2_X1 port map( A1 => n17465, A2 => n25572, ZN => n1313);
   U2016 : INV_X1 port map( A => n18310, ZN => n364);
   U2017 : INV_X1 port map( A => n16615, ZN => n469);
   U2020 : AOI21_X1 port map( B1 => n16964, B2 => n16828, A => n17441, ZN => 
                           n16430);
   U2021 : AND2_X1 port map( A1 => n2508, A2 => n2509, ZN => n491);
   U2022 : NOR2_X1 port map( A1 => n282, A2 => n17175, ZN => n16523);
   U2023 : OAI211_X1 port map( C1 => n16726, C2 => n16974, A => n17335, B => 
                           n16915, ZN => n16605);
   U2026 : OAI21_X1 port map( B1 => n24585, B2 => n16932, A => n1270, ZN => 
                           n1269);
   U2027 : INV_X1 port map( A => n16746, ZN => n828);
   U2029 : OR2_X1 port map( A1 => n16973, A2 => n17335, ZN => n17337);
   U2030 : OR2_X1 port map( A1 => n17482, A2 => n17481, ZN => n2428);
   U2032 : OR2_X1 port map( A1 => n15884, A2 => n15883, ZN => n935);
   U2033 : OR2_X1 port map( A1 => n17242, A2 => n17240, ZN => n1283);
   U2034 : AND2_X1 port map( A1 => n17193, A2 => n17031, ZN => n572);
   U2035 : INV_X1 port map( A => n16731, ZN => n17067);
   U2038 : AOI21_X1 port map( B1 => n16929, B2 => n16932, A => n17059, ZN => 
                           n1270);
   U2040 : INV_X1 port map( A => n17284, ZN => n17230);
   U2041 : OR2_X1 port map( A1 => n17068, A2 => n1139, ZN => n1138);
   U2042 : INV_X1 port map( A => n17302, ZN => n470);
   U2043 : INV_X1 port map( A => n16539, ZN => n365);
   U2044 : MUX2_X1 port map( A => n15163, B => n15162, S => n5447, Z => n17379)
                           ;
   U2046 : INV_X1 port map( A => n17293, ZN => n16951);
   U2048 : INV_X1 port map( A => n16871, ZN => n3602);
   U2049 : INV_X1 port map( A => n17629, ZN => n366);
   U2050 : NOR2_X1 port map( A1 => n17368, A2 => n24471, ZN => n1546);
   U2051 : OR2_X1 port map( A1 => n16795, A2 => n16551, ZN => n16620);
   U2059 : NAND2_X1 port map( A1 => n16245, A2 => n2202, ZN => n17015);
   U2060 : AND3_X1 port map( A1 => n1965, A2 => n16006, A3 => n1964, ZN => 
                           n16846);
   U2061 : INV_X1 port map( A => n17413, ZN => n16957);
   U2062 : INV_X1 port map( A => n25246, ZN => n1230);
   U2064 : OAI21_X1 port map( B1 => n4675, B2 => n4677, A => n4676, ZN => 
                           n17175);
   U2065 : AND2_X1 port map( A1 => n25465, A2 => n17391, ZN => n875);
   U2066 : INV_X1 port map( A => n17227, ZN => n1231);
   U2067 : OR2_X1 port map( A1 => n17227, A2 => n17419, ZN => n1229);
   U2068 : INV_X1 port map( A => n15631, ZN => n17060);
   U2071 : NAND2_X1 port map( A1 => n16033, A2 => n1927, ZN => n17464);
   U2072 : AOI22_X1 port map( A1 => n16228, A2 => n16298, B1 => n16026, B2 => 
                           n16025, ZN => n17461);
   U2074 : INV_X1 port map( A => n17141, ZN => n368);
   U2075 : INV_X1 port map( A => n16261, ZN => n17166);
   U2080 : NOR2_X1 port map( A1 => n17622, A2 => n17624, ZN => n17472);
   U2083 : INV_X1 port map( A => n17088, ZN => n371);
   U2089 : AND2_X1 port map( A1 => n4646, A2 => n4645, ZN => n662);
   U2091 : OAI21_X1 port map( B1 => n4985, B2 => n4984, A => n4983, ZN => 
                           n17288);
   U2092 : AND2_X1 port map( A1 => n4197, A2 => n5212, ZN => n1232);
   U2093 : NOR2_X1 port map( A1 => n1382, A2 => n15866, ZN => n4985);
   U2094 : NAND4_X1 port map( A1 => n16088, A2 => n16104, A3 => n16087, A4 => 
                           n16086, ZN => n16261);
   U2095 : AND2_X1 port map( A1 => n15653, A2 => n16416, ZN => n4984);
   U2096 : INV_X1 port map( A => n17573, ZN => n373);
   U2098 : OAI211_X1 port map( C1 => n16199, C2 => n3143, A => n16201, B => 
                           n3542, ZN => n17386);
   U2099 : AND2_X1 port map( A1 => n3122, A2 => n2212, ZN => n16682);
   U2101 : INV_X1 port map( A => n16765, ZN => n374);
   U2103 : INV_X1 port map( A => n17336, ZN => n376);
   U2104 : OR2_X1 port map( A1 => n15653, A2 => n15868, ZN => n726);
   U2105 : OAI21_X1 port map( B1 => n5414, B2 => n16194, A => n3288, ZN => 
                           n17622);
   U2106 : NOR2_X1 port map( A1 => n1122, A2 => n16342, ZN => n16347);
   U2107 : OR2_X1 port map( A1 => n2251, A2 => n15537, ZN => n516);
   U2108 : OR2_X1 port map( A1 => n2607, A2 => n15564, ZN => n1097);
   U2109 : NOR2_X1 port map( A1 => n16404, A2 => n24062, ZN => n3143);
   U2110 : AND2_X1 port map( A1 => n15677, A2 => n15901, ZN => n521);
   U2112 : NOR2_X1 port map( A1 => n16392, A2 => n24537, ZN => n15850);
   U2114 : BUF_X1 port map( A => n15545, Z => n16475);
   U2115 : XNOR2_X1 port map( A => n2000, B => n14597, ZN => n16042);
   U2116 : INV_X1 port map( A => n15557, ZN => n16010);
   U2117 : XNOR2_X1 port map( A => n14527, B => n14526, ZN => n16389);
   U2118 : INV_X1 port map( A => n24981, ZN => n377);
   U2119 : XNOR2_X1 port map( A => n15140, B => n1105, ZN => n1103);
   U2121 : CLKBUF_X1 port map( A => n15640, Z => n15907);
   U2122 : INV_X1 port map( A => n16109, ZN => n379);
   U2124 : INV_X1 port map( A => n16423, ZN => n707);
   U2125 : XNOR2_X1 port map( A => n13476, B => n13475, ZN => n16333);
   U2126 : XNOR2_X1 port map( A => n13939, B => n13938, ZN => n15970);
   U2129 : XNOR2_X1 port map( A => n15116, B => n15115, ZN => n16360);
   U2130 : XNOR2_X1 port map( A => n15469, B => n15468, ZN => n16473);
   U2131 : INV_X1 port map( A => n16067, ZN => n380);
   U2132 : INV_X1 port map( A => n15646, ZN => n16401);
   U2133 : XNOR2_X1 port map( A => n5192, B => n14742, ZN => n15583);
   U2138 : OR2_X1 port map( A1 => n14926, A2 => n16029, ZN => n2651);
   U2145 : XNOR2_X1 port map( A => n4399, B => n15189, ZN => n15198);
   U2147 : INV_X1 port map( A => n16176, ZN => n15655);
   U2148 : INV_X1 port map( A => n16125, ZN => n381);
   U2149 : CLKBUF_X1 port map( A => n13940, Z => n15971);
   U2150 : XNOR2_X1 port map( A => n15014, B => n15013, ZN => n15560);
   U2153 : XNOR2_X1 port map( A => n14706, B => n14707, ZN => n16107);
   U2154 : INV_X1 port map( A => n15549, ZN => n382);
   U2156 : INV_X1 port map( A => n15715, ZN => n383);
   U2157 : XNOR2_X1 port map( A => n15086, B => n15085, ZN => n16290);
   U2158 : XNOR2_X1 port map( A => n15137, B => n15136, ZN => n16001);
   U2160 : XNOR2_X1 port map( A => n12909, B => n14840, ZN => n16349);
   U2165 : INV_X1 port map( A => n16449, ZN => n385);
   U2166 : INV_X1 port map( A => n16381, ZN => n386);
   U2167 : XNOR2_X1 port map( A => n14380, B => n14379, ZN => n16121);
   U2168 : INV_X1 port map( A => n15564, ZN => n387);
   U2169 : INV_X1 port map( A => n16332, ZN => n388);
   U2171 : XNOR2_X1 port map( A => n14657, B => n14656, ZN => n16129);
   U2172 : XNOR2_X1 port map( A => n14890, B => n14894, ZN => n796);
   U2174 : CLKBUF_X1 port map( A => n16219, Z => n16458);
   U2177 : XNOR2_X1 port map( A => n14904, B => n540, ZN => n14905);
   U2178 : INV_X1 port map( A => n16219, ZN => n389);
   U2179 : XNOR2_X1 port map( A => n12679, B => n14845, ZN => n15070);
   U2180 : XNOR2_X1 port map( A => n4859, B => n1907, ZN => n15405);
   U2181 : INV_X1 port map( A => n14788, ZN => n1111);
   U2182 : INV_X1 port map( A => n3787, ZN => n15188);
   U2183 : XNOR2_X1 port map( A => n15446, B => n15109, ZN => n540);
   U2184 : INV_X1 port map( A => n15177, ZN => n5215);
   U2185 : XNOR2_X1 port map( A => n15293, B => n1104, ZN => n1102);
   U2190 : XNOR2_X1 port map( A => n15138, B => n15483, ZN => n1105);
   U2191 : NAND2_X1 port map( A1 => n4558, A2 => n13690, ZN => n15003);
   U2194 : NAND2_X1 port map( A1 => n4330, A2 => n13483, ZN => n15190);
   U2195 : XNOR2_X1 port map( A => n15386, B => n1833, ZN => n1104);
   U2203 : NAND2_X1 port map( A1 => n2382, A2 => n2381, ZN => n15463);
   U2205 : NAND4_X1 port map( A1 => n14259, A2 => n14260, A3 => n14258, A4 => 
                           n14257, ZN => n14958);
   U2206 : INV_X1 port map( A => n14043, ZN => n985);
   U2207 : NAND3_X1 port map( A1 => n2911, A2 => n13934, A3 => n2910, ZN => 
                           n14997);
   U2209 : OR2_X1 port map( A1 => n13667, A2 => n5753, ZN => n13679);
   U2210 : NAND3_X1 port map( A1 => n5332, A2 => n13567, A3 => n3983, ZN => 
                           n15244);
   U2214 : NOR2_X1 port map( A1 => n13895, A2 => n14130, ZN => n620);
   U2215 : OAI21_X1 port map( B1 => n13655, B2 => n13379, A => n13989, ZN => 
                           n13381);
   U2216 : AND2_X1 port map( A1 => n14206, A2 => n14205, ZN => n13551);
   U2217 : NOR2_X1 port map( A1 => n14327, A2 => n13864, ZN => n5246);
   U2218 : NOR2_X1 port map( A1 => n13596, A2 => n13969, ZN => n5520);
   U2219 : OR2_X1 port map( A1 => n14328, A2 => n14041, ZN => n12803);
   U2221 : OR2_X1 port map( A1 => n10396, A2 => n508, ZN => n967);
   U2223 : OR2_X1 port map( A1 => n13995, A2 => n14235, ZN => n795);
   U2224 : INV_X1 port map( A => n14076, ZN => n13852);
   U2225 : OR2_X1 port map( A1 => n13921, A2 => n13922, ZN => n760);
   U2226 : AND2_X1 port map( A1 => n24949, A2 => n13796, ZN => n14180);
   U2228 : INV_X1 port map( A => n3959, ZN => n13534);
   U2229 : OR2_X1 port map( A1 => n14327, A2 => n14325, ZN => n13863);
   U2230 : NOR2_X1 port map( A1 => n14034, A2 => n14149, ZN => n14151);
   U2231 : OR2_X1 port map( A1 => n13851, A2 => n14078, ZN => n13631);
   U2232 : OR2_X1 port map( A1 => n13609, A2 => n14085, ZN => n1060);
   U2234 : INV_X1 port map( A => n4116, ZN => n14241);
   U2235 : NAND2_X1 port map( A1 => n2317, A2 => n2316, ZN => n14034);
   U2236 : INV_X1 port map( A => n13533, ZN => n14088);
   U2237 : OR2_X1 port map( A1 => n14022, A2 => n4510, ZN => n13607);
   U2238 : INV_X1 port map( A => n13951, ZN => n391);
   U2239 : NAND2_X1 port map( A1 => n1017, A2 => n12890, ZN => n14149);
   U2240 : OR2_X1 port map( A1 => n14089, A2 => n13533, ZN => n3959);
   U2241 : OAI21_X1 port map( B1 => n12778, B2 => n12777, A => n12776, ZN => 
                           n13796);
   U2243 : AND2_X1 port map( A1 => n612, A2 => n13502, ZN => n13506);
   U2244 : AND2_X1 port map( A1 => n13656, A2 => n13918, ZN => n755);
   U2245 : INV_X1 port map( A => n13818, ZN => n392);
   U2248 : NOR2_X1 port map( A1 => n623, A2 => n12913, ZN => n622);
   U2249 : NAND2_X1 port map( A1 => n1081, A2 => n5022, ZN => n4510);
   U2251 : AND4_X1 port map( A1 => n13334, A2 => n13333, A3 => n13332, A4 => 
                           n13331, ZN => n13682);
   U2252 : OAI211_X1 port map( C1 => n1632, C2 => n13134, A => n1631, B => 
                           n1630, ZN => n13552);
   U2254 : INV_X1 port map( A => n14049, ZN => n13518);
   U2255 : INV_X1 port map( A => n14035, ZN => n1028);
   U2256 : OR3_X1 port map( A1 => n12119, A2 => n12118, A3 => n12117, ZN => 
                           n1553);
   U2259 : AND2_X1 port map( A1 => n5470, A2 => n4923, ZN => n1127);
   U2260 : INV_X1 port map( A => n13503, ZN => n612);
   U2261 : AND3_X1 port map( A1 => n5310, A2 => n5309, A3 => n5314, ZN => 
                           n14143);
   U2262 : INV_X1 port map( A => n14324, ZN => n14041);
   U2263 : OR2_X1 port map( A1 => n13128, A2 => n13127, ZN => n14211);
   U2266 : OAI211_X2 port map( C1 => n24487, C2 => n12558, A => n12557, B => 
                           n12556, ZN => n14078);
   U2267 : OAI21_X1 port map( B1 => n13021, B2 => n13020, A => n13019, ZN => 
                           n14225);
   U2268 : AND2_X1 port map( A1 => n12828, A2 => n1508, ZN => n13502);
   U2270 : INV_X1 port map( A => n13907, ZN => n394);
   U2271 : AND3_X1 port map( A1 => n4596, A2 => n4595, A3 => n25053, ZN => 
                           n13681);
   U2272 : INV_X1 port map( A => n24999, ZN => n395);
   U2273 : INV_X1 port map( A => n13419, ZN => n1314);
   U2275 : OR2_X1 port map( A1 => n12463, A2 => n12464, ZN => n493);
   U2276 : AND2_X1 port map( A1 => n1082, A2 => n12504, ZN => n13537);
   U2278 : NAND3_X1 port map( A1 => n12456, A2 => n12458, A3 => n12457, ZN => 
                           n14049);
   U2279 : INV_X1 port map( A => n14269, ZN => n397);
   U2280 : OAI21_X1 port map( B1 => n3975, B2 => n3974, A => n3972, ZN => 
                           n14048);
   U2281 : AND2_X1 port map( A1 => n12661, A2 => n13115, ZN => n1267);
   U2282 : OR2_X1 port map( A1 => n4587, A2 => n12995, ZN => n1018);
   U2283 : OAI21_X1 port map( B1 => n12937, B2 => n4493, A => n1445, ZN => 
                           n4491);
   U2285 : OR2_X1 port map( A1 => n13220, A2 => n24513, ZN => n780);
   U2286 : NOR2_X1 port map( A1 => n12690, A2 => n12910, ZN => n12598);
   U2287 : INV_X1 port map( A => n10200, ZN => n499);
   U2288 : OR2_X1 port map( A1 => n12179, A2 => n13093, ZN => n597);
   U2289 : OR2_X1 port map( A1 => n11328, A2 => n12993, ZN => n1020);
   U2290 : BUF_X1 port map( A => n12868, Z => n13119);
   U2292 : NOR2_X1 port map( A1 => n12834, A2 => n13274, ZN => n1201);
   U2294 : AND2_X1 port map( A1 => n24346, A2 => n13272, ZN => n4446);
   U2295 : INV_X1 port map( A => n12695, ZN => n1200);
   U2296 : OR2_X1 port map( A1 => n12792, A2 => n12995, ZN => n12991);
   U2298 : AND2_X1 port map( A1 => n12859, A2 => n12860, ZN => n12863);
   U2299 : AOI21_X1 port map( B1 => n1069, B2 => n12178, A => n13092, ZN => 
                           n4333);
   U2300 : OR2_X1 port map( A1 => n12433, A2 => n13144, ZN => n1915);
   U2301 : OR2_X1 port map( A1 => n12738, A2 => n13162, ZN => n3710);
   U2302 : AND2_X1 port map( A1 => n12648, A2 => n12178, ZN => n10200);
   U2306 : XNOR2_X1 port map( A => n12026, B => n12027, ZN => n13325);
   U2307 : INV_X1 port map( A => n12859, ZN => n398);
   U2309 : CLKBUF_X1 port map( A => n12519, Z => n12523);
   U2310 : BUF_X1 port map( A => n12520, Z => n13040);
   U2311 : INV_X1 port map( A => n12454, ZN => n13063);
   U2314 : XNOR2_X1 port map( A => n12361, B => n12360, ZN => n12861);
   U2317 : INV_X1 port map( A => n1324, ZN => n10360);
   U2318 : INV_X1 port map( A => n12576, ZN => n399);
   U2320 : XNOR2_X1 port map( A => n9971, B => n9970, ZN => n12178);
   U2321 : INV_X1 port map( A => n13335, ZN => n400);
   U2322 : AND2_X1 port map( A1 => n13027, A2 => n13028, ZN => n563);
   U2324 : INV_X1 port map( A => n13050, ZN => n401);
   U2326 : INV_X1 port map( A => n12725, ZN => n403);
   U2328 : INV_X1 port map( A => n12600, ZN => n404);
   U2329 : XNOR2_X1 port map( A => n12238, B => n12237, ZN => n13110);
   U2333 : XNOR2_X1 port map( A => n11364, B => n11365, ZN => n13213);
   U2335 : XNOR2_X1 port map( A => n12071, B => n12070, ZN => n13329);
   U2336 : INV_X1 port map( A => n13301, ZN => n405);
   U2337 : XNOR2_X1 port map( A => n10708, B => n10709, ZN => n13130);
   U2339 : INV_X1 port map( A => n13124, ZN => n406);
   U2340 : XNOR2_X1 port map( A => n11379, B => n11378, ZN => n12784);
   U2342 : XNOR2_X1 port map( A => n11443, B => n11444, ZN => n12796);
   U2343 : INV_X1 port map( A => n13267, ZN => n407);
   U2345 : INV_X1 port map( A => n12795, ZN => n408);
   U2347 : INV_X1 port map( A => n13056, ZN => n409);
   U2352 : XNOR2_X1 port map( A => n4485, B => n11744, ZN => n13227);
   U2353 : XNOR2_X1 port map( A => n11810, B => n11811, ZN => n13235);
   U2354 : XNOR2_X1 port map( A => n12389, B => n11247, ZN => n11827);
   U2355 : INV_X1 port map( A => n11796, ZN => n3648);
   U2356 : XNOR2_X1 port map( A => n9407, B => n9406, ZN => n9408);
   U2357 : XNOR2_X1 port map( A => n11414, B => n12365, ZN => n11356);
   U2358 : XNOR2_X1 port map( A => n11743, B => n11745, ZN => n4485);
   U2361 : XNOR2_X1 port map( A => n11464, B => n2241, ZN => n11315);
   U2362 : INV_X1 port map( A => n11253, ZN => n11915);
   U2363 : XNOR2_X1 port map( A => n1177, B => n11983, ZN => n12088);
   U2366 : XNOR2_X1 port map( A => n4670, B => n4668, ZN => n11180);
   U2370 : MUX2_X1 port map( A => n11219, B => n11218, S => n233, Z => n11568);
   U2372 : INV_X1 port map( A => n11845, ZN => n12283);
   U2374 : AND3_X1 port map( A1 => n10503, A2 => n3511, A3 => n3510, ZN => 
                           n4670);
   U2375 : AOI22_X1 port map( A1 => n10319, A2 => n10590, B1 => n10583, B2 => 
                           n10318, ZN => n12248);
   U2378 : NAND3_X1 port map( A1 => n10294, A2 => n10295, A3 => n202, ZN => 
                           n11698);
   U2379 : AND3_X1 port map( A1 => n9571, A2 => n9572, A3 => n4040, ZN => 
                           n12402);
   U2380 : NAND4_X1 port map( A1 => n1226, A2 => n1223, A3 => n1227, A4 => 
                           n1225, ZN => n11253);
   U2381 : OAI211_X1 port map( C1 => n10743, C2 => n10858, A => n10742, B => 
                           n10741, ZN => n12066);
   U2382 : AND3_X1 port map( A1 => n527, A2 => n526, A3 => n11050, ZN => n12082
                           );
   U2383 : NAND4_X1 port map( A1 => n11174, A2 => n3384, A3 => n10383, A4 => 
                           n3385, ZN => n11959);
   U2384 : AND2_X1 port map( A1 => n531, A2 => n532, ZN => n530);
   U2389 : OR2_X1 port map( A1 => n11203, A2 => n11204, ZN => n3011);
   U2390 : INV_X1 port map( A => n3443, ZN => n10202);
   U2391 : NAND3_X1 port map( A1 => n10928, A2 => n10929, A3 => n4691, ZN => 
                           n12315);
   U2392 : AND2_X1 port map( A1 => n10804, A2 => n10798, ZN => n10806);
   U2393 : OAI21_X1 port map( B1 => n10642, B2 => n11046, A => n529, ZN => 
                           n5671);
   U2395 : NOR2_X1 port map( A1 => n10967, A2 => n10971, ZN => n10818);
   U2396 : MUX2_X1 port map( A => n9210, B => n9209, S => n10587, Z => n9216);
   U2397 : OR2_X1 port map( A1 => n10805, A2 => n10799, ZN => n735);
   U2398 : OR2_X1 port map( A1 => n11082, A2 => n5559, ZN => n1264);
   U2399 : OR2_X1 port map( A1 => n11205, A2 => n11338, ZN => n10821);
   U2400 : OR2_X1 port map( A1 => n10527, A2 => n11529, ZN => n525);
   U2402 : OR2_X1 port map( A1 => n11091, A2 => n1057, ZN => n1056);
   U2403 : INV_X1 port map( A => n10491, ZN => n10233);
   U2405 : INV_X1 port map( A => n11212, ZN => n3868);
   U2406 : NOR2_X1 port map( A1 => n11099, A2 => n939, ZN => n10782);
   U2408 : NOR2_X1 port map( A1 => n10617, A2 => n10411, ZN => n559);
   U2409 : INV_X1 port map( A => n11024, ZN => n895);
   U2410 : INV_X1 port map( A => n11302, ZN => n11300);
   U2412 : INV_X1 port map( A => n10887, ZN => n10301);
   U2413 : INV_X1 port map( A => n939, ZN => n10911);
   U2414 : CLKBUF_X1 port map( A => n11172, Z => n1338);
   U2415 : INV_X1 port map( A => n232, ZN => n10812);
   U2416 : INV_X1 port map( A => n10583, ZN => n9443);
   U2418 : INV_X1 port map( A => n10798, ZN => n10805);
   U2419 : INV_X1 port map( A => n4531, ZN => n528);
   U2420 : INV_X1 port map( A => n11059, ZN => n410);
   U2424 : NAND2_X1 port map( A1 => n5535, A2 => n5534, ZN => n10762);
   U2426 : INV_X1 port map( A => n9432, ZN => n412);
   U2427 : INV_X1 port map( A => n10523, ZN => n11024);
   U2428 : INV_X1 port map( A => n10277, ZN => n413);
   U2430 : OR2_X1 port map( A1 => n1181, A2 => n1963, ZN => n10798);
   U2431 : INV_X1 port map( A => n11342, ZN => n414);
   U2432 : OR2_X1 port map( A1 => n9618, A2 => n9617, ZN => n660);
   U2434 : INV_X1 port map( A => n11499, ZN => n1218);
   U2435 : AND2_X1 port map( A1 => n10778, A2 => n9502, ZN => n1552);
   U2436 : INV_X1 port map( A => n10886, ZN => n10541);
   U2438 : NAND2_X1 port map( A1 => n9502, A2 => n10778, ZN => n11099);
   U2439 : OAI21_X1 port map( B1 => n9840, B2 => n10099, A => n9839, ZN => 
                           n10703);
   U2440 : INV_X1 port map( A => n11032, ZN => n415);
   U2441 : AND2_X1 port map( A1 => n9250, A2 => n1816, ZN => n10855);
   U2444 : OR2_X1 port map( A1 => n9201, A2 => n627, ZN => n9582);
   U2446 : INV_X1 port map( A => n11039, ZN => n416);
   U2448 : INV_X1 port map( A => n11163, ZN => n417);
   U2449 : INV_X1 port map( A => n10889, ZN => n418);
   U2453 : OAI211_X1 port map( C1 => n3722, C2 => n5609, A => n5608, B => n3721
                           , ZN => n11121);
   U2454 : OR2_X1 port map( A1 => n9128, A2 => n9129, ZN => n11036);
   U2455 : OAI21_X1 port map( B1 => n9598, B2 => n9597, A => n9596, ZN => 
                           n10614);
   U2458 : AOI22_X1 port map( A1 => n2140, A2 => n1796, B1 => n9501, B2 => n246
                           , ZN => n10778);
   U2462 : INV_X1 port map( A => n11298, ZN => n419);
   U2464 : INV_X1 port map( A => n11130, ZN => n420);
   U2466 : OAI22_X1 port map( A1 => n5523, A2 => n24054, B1 => n9945, B2 => 
                           n1165, ZN => n1181);
   U2467 : OAI21_X1 port map( B1 => n10122, B2 => n9841, A => n24087, ZN => 
                           n2256);
   U2468 : OR2_X1 port map( A1 => n9225, A2 => n9740, ZN => n1168);
   U2469 : NOR2_X1 port map( A1 => n2294, A2 => n1021, ZN => n9693);
   U2470 : INV_X1 port map( A => n3305, ZN => n699);
   U2471 : INV_X1 port map( A => n24085, ZN => n2257);
   U2474 : OR2_X1 port map( A1 => n9808, A2 => n9807, ZN => n1318);
   U2475 : INV_X1 port map( A => n9417, ZN => n9758);
   U2477 : NOR2_X1 port map( A1 => n9872, A2 => n1021, ZN => n1519);
   U2479 : AND2_X1 port map( A1 => n9886, A2 => n9565, ZN => n956);
   U2480 : AOI21_X1 port map( B1 => n3292, B2 => n9281, A => n9468, ZN => n665)
                           ;
   U2482 : AND2_X1 port map( A1 => n8521, A2 => n9798, ZN => n9314);
   U2483 : BUF_X1 port map( A => n8483, Z => n9999);
   U2484 : OR2_X1 port map( A1 => n24446, A2 => n4096, ZN => n4097);
   U2485 : INV_X1 port map( A => n10108, ZN => n9524);
   U2487 : INV_X1 port map( A => n9237, ZN => n9697);
   U2488 : INV_X1 port map( A => n4254, ZN => n1275);
   U2489 : OR2_X1 port map( A1 => n9295, A2 => n9781, ZN => n5025);
   U2490 : AND2_X1 port map( A1 => n24535, A2 => n9990, ZN => n9425);
   U2491 : NOR2_X1 port map( A1 => n25005, A2 => n9418, ZN => n9615);
   U2492 : INV_X1 port map( A => n9027, ZN => n1021);
   U2493 : CLKBUF_X1 port map( A => n9297, Z => n9780);
   U2495 : INV_X1 port map( A => n3292, ZN => n1185);
   U2496 : BUF_X1 port map( A => n9398, Z => n10136);
   U2498 : INV_X1 port map( A => n10251, ZN => n10250);
   U2499 : NOR2_X1 port map( A1 => n24087, A2 => n9843, ZN => n2413);
   U2500 : OR2_X1 port map( A1 => n10058, A2 => n4096, ZN => n794);
   U2501 : CLKBUF_X1 port map( A => n9419, Z => n9754);
   U2505 : INV_X1 port map( A => n8359, ZN => n421);
   U2507 : INV_X1 port map( A => n24534, ZN => n422);
   U2509 : XNOR2_X1 port map( A => n7454, B => n7453, ZN => n9962);
   U2511 : INV_X1 port map( A => n24505, ZN => n424);
   U2514 : INV_X1 port map( A => n9779, ZN => n425);
   U2515 : XNOR2_X1 port map( A => n8785, B => n8784, ZN => n9418);
   U2516 : INV_X1 port map( A => n9491, ZN => n426);
   U2517 : INV_X1 port map( A => n9945, ZN => n9942);
   U2518 : BUF_X1 port map( A => n8523, Z => n9530);
   U2519 : BUF_X1 port map( A => n10071, Z => n1330);
   U2520 : BUF_X1 port map( A => n9218, Z => n10065);
   U2521 : XNOR2_X1 port map( A => n7042, B => n7041, ZN => n9918);
   U2522 : INV_X1 port map( A => n10109, ZN => n4254);
   U2524 : XNOR2_X1 port map( A => n8816, B => n8817, ZN => n10018);
   U2526 : INV_X1 port map( A => n10071, ZN => n427);
   U2528 : XNOR2_X1 port map( A => n8464, B => n8463, ZN => n9786);
   U2531 : XNOR2_X1 port map( A => n8944, B => n8943, ZN => n10046);
   U2532 : XNOR2_X1 port map( A => n8767, B => n8768, ZN => n9752);
   U2534 : XNOR2_X1 port map( A => n7497, B => n7496, ZN => n9964);
   U2536 : INV_X1 port map( A => n9837, ZN => n428);
   U2537 : XNOR2_X1 port map( A => n8626, B => n8625, ZN => n10109);
   U2540 : INV_X1 port map( A => n9127, ZN => n429);
   U2541 : XNOR2_X1 port map( A => n8559, B => n2274, ZN => n2276);
   U2542 : INV_X1 port map( A => n8951, ZN => n5184);
   U2543 : XNOR2_X1 port map( A => n5344, B => n8798, ZN => n8198);
   U2545 : XNOR2_X1 port map( A => n8613, B => n8280, ZN => n9089);
   U2546 : XNOR2_X1 port map( A => n8980, B => n1110, ZN => n8778);
   U2548 : XNOR2_X1 port map( A => n8787, B => n8450, ZN => n9012);
   U2557 : OAI21_X1 port map( B1 => n5116, B2 => n7952, A => n2490, ZN => n9159
                           );
   U2560 : OAI21_X1 port map( B1 => n3267, B2 => n7843, A => n3265, ZN => n8615
                           );
   U2561 : NAND3_X1 port map( A1 => n7745, A2 => n7746, A3 => n1972, ZN => 
                           n9002);
   U2562 : OR2_X1 port map( A1 => n4975, A2 => n7859, ZN => n8789);
   U2567 : NAND2_X1 port map( A1 => n7484, A2 => n4001, ZN => n8795);
   U2569 : NOR2_X1 port map( A1 => n7807, A2 => n7806, ZN => n8450);
   U2571 : NAND3_X1 port map( A1 => n7178, A2 => n7177, A3 => n7176, ZN => 
                           n8917);
   U2572 : MUX2_X1 port map( A => n7446, B => n7447, S => n5607, Z => n8492);
   U2574 : NAND3_X1 port map( A1 => n2263, A2 => n7509, A3 => n2261, ZN => 
                           n8769);
   U2575 : AND2_X1 port map( A1 => n7158, A2 => n5345, ZN => n7161);
   U2577 : NAND3_X1 port map( A1 => n1848, A2 => n7137, A3 => n7138, ZN => 
                           n8647);
   U2579 : NAND2_X1 port map( A1 => n7729, A2 => n7728, ZN => n8914);
   U2581 : AOI22_X1 port map( A1 => n8024, A2 => n3258, B1 => n3259, B2 => 
                           n7532, ZN => n3257);
   U2583 : OR2_X1 port map( A1 => n3236, A2 => n2640, ZN => n3235);
   U2584 : AND2_X1 port map( A1 => n4145, A2 => n7953, ZN => n842);
   U2585 : AND2_X1 port map( A1 => n7282, A2 => n7281, ZN => n533);
   U2586 : OAI21_X1 port map( B1 => n806, B2 => n1345, A => n2223, ZN => n7487)
                           ;
   U2588 : OAI21_X1 port map( B1 => n3500, B2 => n7580, A => n3498, ZN => n8981
                           );
   U2589 : AND2_X1 port map( A1 => n7533, A2 => n7747, ZN => n3258);
   U2591 : INV_X1 port map( A => n7349, ZN => n1279);
   U2592 : OR2_X1 port map( A1 => n7651, A2 => n7650, ZN => n989);
   U2593 : OAI21_X1 port map( B1 => n7322, B2 => n7890, A => n311, ZN => n1124)
                           ;
   U2594 : INV_X1 port map( A => n941, ZN => n7622);
   U2596 : OR2_X1 port map( A1 => n2522, A2 => n8003, ZN => n736);
   U2598 : AND2_X1 port map( A1 => n7537, A2 => n7748, ZN => n8011);
   U2599 : INV_X1 port map( A => n7444, ZN => n7163);
   U2600 : OR2_X1 port map( A1 => n7593, A2 => n7592, ZN => n1190);
   U2601 : INV_X1 port map( A => n7754, ZN => n7542);
   U2602 : OR2_X1 port map( A1 => n7760, A2 => n7646, ZN => n6194);
   U2603 : INV_X1 port map( A => n7683, ZN => n7235);
   U2605 : INV_X1 port map( A => n512, ZN => n7634);
   U2607 : INV_X1 port map( A => n1162, ZN => n7676);
   U2608 : INV_X1 port map( A => n7074, ZN => n7506);
   U2609 : OR3_X1 port map( A1 => n7350, A2 => n5468, A3 => n7346, ZN => n7253)
                           ;
   U2610 : INV_X1 port map( A => n7078, ZN => n3275);
   U2611 : NAND2_X1 port map( A1 => n6581, A2 => n5604, ZN => n7924);
   U2612 : INV_X1 port map( A => n7914, ZN => n430);
   U2614 : CLKBUF_X1 port map( A => n6806, Z => n7667);
   U2615 : CLKBUF_X1 port map( A => n7246, Z => n7855);
   U2616 : OAI21_X1 port map( B1 => n6443, B2 => n6296, A => n6213, ZN => n2640
                           );
   U2617 : OR2_X1 port map( A1 => n270, A2 => n7962, ZN => n584);
   U2618 : INV_X1 port map( A => n7533, ZN => n1975);
   U2619 : INV_X1 port map( A => n2624, ZN => n7748);
   U2620 : AND2_X1 port map( A1 => n2401, A2 => n2400, ZN => n2402);
   U2621 : NOR2_X1 port map( A1 => n1162, A2 => n1085, ZN => n1084);
   U2622 : NAND2_X1 port map( A1 => n3608, A2 => n6313, ZN => n7861);
   U2624 : NAND2_X1 port map( A1 => n764, A2 => n1174, ZN => n7683);
   U2626 : NAND2_X1 port map( A1 => n1433, A2 => n2899, ZN => n7732);
   U2627 : INV_X1 port map( A => n7423, ZN => n431);
   U2628 : NAND2_X1 port map( A1 => n943, A2 => n944, ZN => n942);
   U2633 : OAI211_X1 port map( C1 => n5729, C2 => n6049, A => n504, B => n502, 
                           ZN => n7108);
   U2636 : AND2_X1 port map( A1 => n5890, A2 => n5889, ZN => n7896);
   U2637 : INV_X1 port map( A => n7217, ZN => n433);
   U2638 : INV_X1 port map( A => n7983, ZN => n7827);
   U2640 : INV_X1 port map( A => n7224, ZN => n434);
   U2641 : OAI21_X1 port map( B1 => n5142, B2 => n5143, A => n6273, ZN => n7803
                           );
   U2646 : AND2_X1 port map( A1 => n5912, A2 => n5911, ZN => n7347);
   U2647 : INV_X1 port map( A => n7915, ZN => n435);
   U2648 : INV_X1 port map( A => n7664, ZN => n436);
   U2650 : NAND2_X1 port map( A1 => n6103, A2 => n6102, ZN => n7768);
   U2651 : NAND2_X1 port map( A1 => n1695, A2 => n568, ZN => n1162);
   U2653 : INV_X1 port map( A => n6323, ZN => n944);
   U2654 : OAI211_X1 port map( C1 => n6412, C2 => n6051, A => n6411, B => n6410
                           , ZN => n7853);
   U2658 : AOI21_X1 port map( B1 => n5088, B2 => n7024, A => n2738, ZN => n2737
                           );
   U2661 : INV_X1 port map( A => n7962, ZN => n437);
   U2663 : OAI21_X1 port map( B1 => n709, B2 => n6553, A => n708, ZN => n1750);
   U2664 : AOI22_X1 port map( A1 => n7005, A2 => n6835, B1 => n7004, B2 => 
                           n6836, ZN => n467);
   U2665 : OR2_X1 port map( A1 => n6177, A2 => n6178, ZN => n7646);
   U2667 : INV_X1 port map( A => n1379, ZN => n1085);
   U2668 : OR2_X1 port map( A1 => n6463, A2 => n6464, ZN => n773);
   U2669 : AND2_X1 port map( A1 => n6274, A2 => n6324, ZN => n6522);
   U2670 : OAI21_X1 port map( B1 => n6906, B2 => n6905, A => n6373, ZN => n6475
                           );
   U2671 : AND2_X1 port map( A1 => n6519, A2 => n6275, ZN => n6524);
   U2672 : AND2_X1 port map( A1 => n6957, A2 => n6705, ZN => n709);
   U2673 : AND2_X1 port map( A1 => n6641, A2 => n6642, ZN => n5635);
   U2674 : NAND2_X1 port map( A1 => n6328, A2 => n5451, ZN => n1079);
   U2676 : OAI21_X1 port map( B1 => n669, B2 => n6674, A => n668, ZN => n6676);
   U2677 : INV_X1 port map( A => n6570, ZN => n4754);
   U2678 : OR2_X1 port map( A1 => n6588, A2 => n625, ZN => n6226);
   U2682 : CLKBUF_X1 port map( A => n6187, Z => n6347);
   U2684 : INV_X1 port map( A => n6999, ZN => n947);
   U2687 : OR2_X1 port map( A1 => n7035, A2 => n625, ZN => n6591);
   U2688 : INV_X1 port map( A => n625, ZN => n7033);
   U2689 : INV_X1 port map( A => n4324, ZN => n708);
   U2690 : BUF_X1 port map( A => n6381, Z => n7025);
   U2691 : INV_X1 port map( A => n6453, ZN => n1106);
   U2693 : INV_X1 port map( A => n6683, ZN => n6939);
   U2696 : INV_X1 port map( A => n6174, ZN => n438);
   U2697 : INV_X1 port map( A => n6367, ZN => n439);
   U2700 : BUF_X1 port map( A => n5887, Z => n6679);
   U2702 : INV_X1 port map( A => n6324, ZN => n440);
   U2703 : NOR2_X1 port map( A1 => n6757, A2 => n6578, ZN => n669);
   U2705 : INV_X1 port map( A => n1804, ZN => n931);
   U2706 : INV_X1 port map( A => n5824, ZN => n6372);
   U2707 : INV_X1 port map( A => n6496, ZN => n441);
   U2709 : INV_X1 port map( A => n6578, ZN => n5805);
   U2710 : INV_X1 port map( A => n23868, ZN => n4189);
   U2711 : INV_X1 port map( A => n6381, ZN => n442);
   U2712 : AOI21_X1 port map( B1 => n6498, B2 => n6034, A => n6434, ZN => n2218
                           );
   U2714 : AND3_X1 port map( A1 => n6777, A2 => n6198, A3 => n6775, ZN => n1295
                           );
   U2715 : CLKBUF_X1 port map( A => Key(102), Z => n677);
   U2717 : CLKBUF_X1 port map( A => Key(140), Z => n3190);
   U2721 : CLKBUF_X1 port map( A => Key(64), Z => n2970);
   U2722 : CLKBUF_X1 port map( A => Key(53), Z => n2215);
   U2723 : INV_X1 port map( A => n2744, ZN => n444);
   U2725 : CLKBUF_X1 port map( A => Key(30), Z => n3133);
   U2726 : XNOR2_X1 port map( A => Key(44), B => Plaintext(44), ZN => n6955);
   U2727 : INV_X1 port map( A => n1952, ZN => n445);
   U2728 : CLKBUF_X1 port map( A => Key(57), Z => n887);
   U2729 : CLKBUF_X1 port map( A => Key(167), Z => n2743);
   U2730 : CLKBUF_X1 port map( A => Key(151), Z => n1874);
   U2731 : CLKBUF_X1 port map( A => Key(61), Z => n21046);
   U2732 : CLKBUF_X1 port map( A => Key(91), Z => n1935);
   U2733 : CLKBUF_X1 port map( A => Key(164), Z => n2137);
   U2734 : CLKBUF_X1 port map( A => Key(90), Z => n2034);
   U2737 : INV_X1 port map( A => n768, ZN => n447);
   U2740 : INV_X1 port map( A => n7008, ZN => n448);
   U2741 : CLKBUF_X1 port map( A => Key(187), Z => n888);
   U2743 : XNOR2_X1 port map( A => Plaintext(145), B => Key(145), ZN => n5824);
   U2744 : INV_X1 port map( A => n2834, ZN => n449);
   U2746 : INV_X1 port map( A => n1833, ZN => n450);
   U2749 : XNOR2_X1 port map( A => Key(187), B => Plaintext(187), ZN => n6195);
   U2750 : CLKBUF_X1 port map( A => Key(132), Z => n3155);
   U2751 : CLKBUF_X1 port map( A => Key(54), Z => n2795);
   U2753 : INV_X1 port map( A => n22886, ZN => n451);
   U2754 : INV_X1 port map( A => n1865, ZN => n452);
   U2756 : CLKBUF_X1 port map( A => Key(179), Z => n21964);
   U2757 : INV_X1 port map( A => n6050, ZN => n453);
   U2758 : CLKBUF_X1 port map( A => Key(122), Z => n23476);
   U2759 : CLKBUF_X1 port map( A => Key(186), Z => n1726);
   U2760 : XNOR2_X1 port map( A => Key(85), B => Plaintext(85), ZN => n6243);
   U2761 : CLKBUF_X1 port map( A => Key(134), Z => n729);
   U2762 : CLKBUF_X1 port map( A => Key(8), Z => n3152);
   U2763 : INV_X1 port map( A => n7029, ZN => n454);
   U2764 : CLKBUF_X1 port map( A => Key(26), Z => n3073);
   U2765 : INV_X1 port map( A => n765, ZN => n455);
   U2766 : CLKBUF_X1 port map( A => Key(13), Z => n3125);
   U2767 : NAND2_X1 port map( A1 => n19323, A2 => n456, ZN => n19936);
   U2768 : NAND2_X1 port map( A1 => n458, A2 => n457, ZN => n456);
   U2769 : OAI211_X2 port map( C1 => n13378, C2 => n13484, A => n205, B => n459
                           , ZN => n14805);
   U2770 : NAND2_X1 port map( A1 => n13485, A2 => n652, ZN => n459);
   U2772 : OR2_X1 port map( A1 => n18959, A2 => n19470, ZN => n18961);
   U2773 : NAND2_X1 port map( A1 => n12272, A2 => n12864, ZN => n13115);
   U2775 : AOI22_X1 port map( A1 => n21919, A2 => n329, B1 => n22451, B2 => 
                           n22323, ZN => n21920);
   U2777 : NAND2_X1 port map( A1 => n1192, A2 => n1196, ZN => n7237);
   U2779 : NOR2_X1 port map( A1 => n5415, A2 => n22824, ZN => n462);
   U2780 : OAI21_X1 port map( B1 => n23948, B2 => n22826, A => n463, ZN => 
                           n23949);
   U2782 : OAI211_X2 port map( C1 => n10894, C2 => n3119, A => n465, B => n464,
                           ZN => n12020);
   U2783 : NAND2_X1 port map( A1 => n10892, A2 => n3119, ZN => n464);
   U2784 : NAND2_X1 port map( A1 => n10893, A2 => n11085, ZN => n465);
   U2786 : NAND2_X1 port map( A1 => n470, A2 => n469, ZN => n468);
   U2790 : NAND2_X1 port map( A1 => n7192, A2 => n8371, ZN => n472);
   U2791 : NAND2_X1 port map( A1 => n17142, A2 => n17141, ZN => n473);
   U2793 : NAND2_X1 port map( A1 => n3306, A2 => n16611, ZN => n16614);
   U2794 : NAND3_X1 port map( A1 => n7828, A2 => n7829, A3 => n7827, ZN => 
                           n7830);
   U2795 : NAND2_X1 port map( A1 => n1694, A2 => n12965, ZN => n12968);
   U2796 : NAND2_X1 port map( A1 => n477, A2 => n475, ZN => n7717);
   U2797 : NAND2_X1 port map( A1 => n8371, A2 => n24577, ZN => n475);
   U2799 : NAND2_X1 port map( A1 => n7715, A2 => n24878, ZN => n477);
   U2800 : NAND3_X1 port map( A1 => n16509, A2 => n16508, A3 => n25376, ZN => 
                           n1812);
   U2802 : OAI211_X1 port map( C1 => n16235, C2 => n257, A => n478, B => n385, 
                           ZN => n14974);
   U2803 : NAND2_X1 port map( A1 => n16235, A2 => n16450, ZN => n478);
   U2804 : NAND2_X1 port map( A1 => n480, A2 => n479, ZN => n10769);
   U2805 : NAND3_X1 port map( A1 => n10767, A2 => n10890, A3 => n4422, ZN => 
                           n479);
   U2806 : NAND2_X1 port map( A1 => n10768, A2 => n412, ZN => n480);
   U2807 : MUX2_X1 port map( A => n23967, B => n25017, S => n23972, Z => n23959
                           );
   U2810 : OAI211_X2 port map( C1 => n1604, C2 => n20369, A => n484, B => n483,
                           ZN => n21750);
   U2811 : NAND2_X1 port map( A1 => n277, A2 => n24454, ZN => n483);
   U2812 : NAND2_X1 port map( A1 => n20370, A2 => n24531, ZN => n484);
   U2814 : NAND2_X1 port map( A1 => n17129, A2 => n17132, ZN => n486);
   U2815 : XNOR2_X1 port map( A => n488, B => n11348, ZN => n11349);
   U2816 : XNOR2_X1 port map( A => n11347, B => n11346, ZN => n488);
   U2817 : NAND3_X1 port map( A1 => n4013, A2 => n413, A3 => n10830, ZN => 
                           n9646);
   U2818 : NAND3_X1 port map( A1 => n4774, A2 => n17166, A3 => n25219, ZN => 
                           n514);
   U2822 : NAND3_X1 port map( A1 => n2485, A2 => n5624, A3 => n13353, ZN => 
                           n2484);
   U2823 : NAND2_X1 port map( A1 => n6718, A2 => n6712, ZN => n6713);
   U2824 : NAND2_X1 port map( A1 => n16193, A2 => n16191, ZN => n15677);
   U2829 : NAND3_X1 port map( A1 => n2728, A2 => n4554, A3 => n2727, ZN => n492
                           );
   U2831 : INV_X1 port map( A => Plaintext(65), ZN => n495);
   U2832 : NAND3_X1 port map( A1 => n9454, A2 => n9564, A3 => n9885, ZN => 
                           n2720);
   U2833 : OAI211_X1 port map( C1 => n5269, C2 => n15921, A => n496, B => n389,
                           ZN => n15779);
   U2834 : NAND2_X1 port map( A1 => n16464, A2 => n15921, ZN => n496);
   U2835 : NAND2_X1 port map( A1 => n13307, A2 => n11722, ZN => n13309);
   U2838 : OR2_X1 port map( A1 => n10201, A2 => n5323, ZN => n498);
   U2839 : NAND3_X1 port map( A1 => n1080, A2 => n4332, A3 => n499, ZN => n1081
                           );
   U2840 : AND2_X1 port map( A1 => n6622, A2 => n6114, ZN => n500);
   U2842 : NAND2_X1 port map( A1 => n1609, A2 => n6114, ZN => n505);
   U2843 : NAND2_X1 port map( A1 => n1609, A2 => n500, ZN => n504);
   U2844 : NAND2_X1 port map( A1 => n505, A2 => n501, ZN => n1610);
   U2845 : NAND2_X1 port map( A1 => n6619, A2 => n316, ZN => n501);
   U2846 : NAND3_X1 port map( A1 => n6619, A2 => n6622, A3 => n316, ZN => n502)
                           ;
   U2847 : INV_X1 port map( A => n507, ZN => n3302);
   U2848 : NOR2_X1 port map( A1 => n508, A2 => n14158, ZN => n13467);
   U2849 : NAND2_X1 port map( A1 => n508, A2 => n14158, ZN => n13776);
   U2851 : NOR2_X1 port map( A1 => n5080, A2 => n24999, ZN => n11022);
   U2852 : NAND2_X1 port map( A1 => n5079, A2 => n507, ZN => n13469);
   U2853 : OR2_X1 port map( A1 => n22634, A2 => n22633, ZN => n510);
   U2854 : NAND2_X1 port map( A1 => n22636, A2 => n510, ZN => n22641);
   U2856 : NAND2_X1 port map( A1 => n512, A2 => n25253, ZN => n7914);
   U2857 : NAND2_X1 port map( A1 => n512, A2 => n7449, ZN => n6486);
   U2858 : NAND2_X1 port map( A1 => n3347, A2 => n511, ZN => n7398);
   U2859 : AND2_X1 port map( A1 => n512, A2 => n7918, ZN => n511);
   U2860 : NAND2_X1 port map( A1 => n430, A2 => n312, ZN => n8075);
   U2861 : NAND3_X1 port map( A1 => n3348, A2 => n512, A3 => n435, ZN => n7159)
                           ;
   U2862 : NAND3_X1 port map( A1 => n2376, A2 => n2679, A3 => n22592, ZN => 
                           n710);
   U2863 : OR2_X1 port map( A1 => n25475, A2 => n8839, ZN => n5277);
   U2865 : AOI21_X1 port map( B1 => n20041, B2 => n20039, A => n19862, ZN => 
                           n513);
   U2868 : NAND2_X1 port map( A1 => n515, A2 => n1841, ZN => n18473);
   U2869 : NAND2_X1 port map( A1 => n517, A2 => n516, ZN => n17088);
   U2870 : OAI22_X1 port map( A1 => n15536, A2 => n15788, B1 => n15535, B2 => 
                           n2253, ZN => n517);
   U2871 : OR2_X1 port map( A1 => n16231, A2 => n16232, ZN => n15935);
   U2872 : OAI22_X1 port map( A1 => n2814, A2 => n16739, B1 => n371, B2 => 
                           n16649, ZN => n17090);
   U2873 : AOI22_X2 port map( A1 => n5471, A2 => n12206, B1 => n5472, B2 => 
                           n3876, ZN => n13460);
   U2874 : XNOR2_X1 port map( A => n12207, B => n455, ZN => n12208);
   U2877 : OAI21_X1 port map( B1 => n19400, B2 => n18900, A => n19163, ZN => 
                           n519);
   U2880 : NAND2_X1 port map( A1 => n23995, A2 => n25079, ZN => n520);
   U2881 : OR2_X1 port map( A1 => n10308, A2 => n4998, ZN => n758);
   U2882 : NAND2_X1 port map( A1 => n6341, A2 => n6187, ZN => n6448);
   U2883 : NOR2_X1 port map( A1 => n521, A2 => n15676, ZN => n15678);
   U2884 : NAND2_X1 port map( A1 => n523, A2 => n17449, ZN => n522);
   U2887 : NAND2_X1 port map( A1 => n2714, A2 => n10552, ZN => n3196);
   U2889 : NAND3_X2 port map( A1 => n10526, A2 => n525, A3 => n10525, ZN => 
                           n12277);
   U2890 : NAND2_X1 port map( A1 => n3556, A2 => n3555, ZN => n16112);
   U2892 : NAND2_X1 port map( A1 => n10013, A2 => n4531, ZN => n526);
   U2893 : NAND2_X1 port map( A1 => n10014, A2 => n528, ZN => n527);
   U2896 : NAND2_X1 port map( A1 => n11046, A2 => n11044, ZN => n529);
   U2897 : INV_X1 port map( A => n10158, ZN => n3305);
   U2898 : OR2_X1 port map( A1 => n1100, A2 => n22359, ZN => n972);
   U2899 : NOR2_X1 port map( A1 => n5475, A2 => n20257, ZN => n5473);
   U2900 : INV_X1 port map( A => n20255, ZN => n20412);
   U2901 : NAND2_X1 port map( A1 => n10242, A2 => n10497, ZN => n531);
   U2902 : NAND2_X1 port map( A1 => n10241, A2 => n2546, ZN => n532);
   U2903 : NAND2_X1 port map( A1 => n14075, A2 => n14076, ZN => n13629);
   U2905 : OR2_X1 port map( A1 => n25046, A2 => n8327, ZN => n9591);
   U2906 : OR2_X1 port map( A1 => n20422, A2 => n20419, ZN => n1660);
   U2907 : NAND2_X1 port map( A1 => n17160, A2 => n17163, ZN => n16264);
   U2910 : NAND2_X1 port map( A1 => n21293, A2 => n22771, ZN => n535);
   U2912 : OAI21_X1 port map( B1 => n23833, B2 => n23827, A => n318, ZN => n536
                           );
   U2913 : NAND2_X1 port map( A1 => n537, A2 => n11125, ZN => n9243);
   U2914 : OAI22_X1 port map( A1 => n305, A2 => n10460, B1 => n11124, B2 => 
                           n10850, ZN => n537);
   U2915 : NAND2_X1 port map( A1 => n16035, A2 => n16733, ZN => n2096);
   U2916 : OAI21_X1 port map( B1 => n13030, B2 => n302, A => n538, ZN => n12494
                           );
   U2917 : NAND2_X1 port map( A1 => n12786, A2 => n13023, ZN => n538);
   U2918 : AOI22_X1 port map( A1 => n3627, A2 => n3783, B1 => n3626, B2 => 
                           n17316, ZN => n539);
   U2919 : INV_X1 port map( A => n542, ZN => n541);
   U2920 : OAI21_X1 port map( B1 => n11175, B2 => n10940, A => n10939, ZN => 
                           n542);
   U2921 : NAND2_X1 port map( A1 => n543, A2 => n1375, ZN => n11242);
   U2923 : NAND2_X1 port map( A1 => n12624, A2 => n12878, ZN => n5191);
   U2924 : NAND2_X1 port map( A1 => n14182, A2 => n14178, ZN => n13797);
   U2925 : INV_X1 port map( A => n13234, ZN => n545);
   U2926 : NAND2_X1 port map( A1 => n12936, A2 => n13234, ZN => n546);
   U2929 : NAND2_X1 port map( A1 => n18903, A2 => n353, ZN => n548);
   U2930 : NAND2_X1 port map( A1 => n18904, A2 => n3773, ZN => n549);
   U2935 : OAI211_X1 port map( C1 => n22624, C2 => n23058, A => n553, B => n552
                           , ZN => n22626);
   U2936 : NAND2_X1 port map( A1 => n22643, A2 => n23059, ZN => n552);
   U2937 : NAND2_X1 port map( A1 => n23055, A2 => n22698, ZN => n553);
   U2938 : NAND2_X1 port map( A1 => n23301, A2 => n554, ZN => n664);
   U2939 : AOI22_X1 port map( A1 => n23298, A2 => n23297, B1 => n23300, B2 => 
                           n23299, ZN => n554);
   U2940 : INV_X1 port map( A => n19422, ZN => n1309);
   U2941 : NAND3_X1 port map( A1 => n555, A2 => n4475, A3 => n4474, ZN => 
                           n23977);
   U2942 : NAND2_X1 port map( A1 => n23975, A2 => n23987, ZN => n555);
   U2944 : INV_X1 port map( A => n557, ZN => n556);
   U2945 : OAI21_X1 port map( B1 => n9827, B2 => n10186, A => n9586, ZN => n557
                           );
   U2946 : NAND2_X1 port map( A1 => n561, A2 => n558, ZN => n10345);
   U2947 : NAND2_X1 port map( A1 => n560, A2 => n559, ZN => n558);
   U2948 : INV_X1 port map( A => n10341, ZN => n560);
   U2949 : NAND2_X1 port map( A1 => n10342, A2 => n10411, ZN => n561);
   U2951 : OR2_X1 port map( A1 => n16106, A2 => n16108, ZN => n15854);
   U2952 : INV_X1 port map( A => n13074, ZN => n12708);
   U2953 : NAND2_X1 port map( A1 => n4124, A2 => n562, ZN => n4123);
   U2954 : NAND2_X1 port map( A1 => n13029, A2 => n563, ZN => n562);
   U2955 : NAND3_X2 port map( A1 => n564, A2 => n15079, A3 => n15080, ZN => 
                           n17424);
   U2957 : NAND2_X1 port map( A1 => n13350, A2 => n12349, ZN => n12330);
   U2959 : NAND3_X1 port map( A1 => n424, A2 => n10089, A3 => n1348, ZN => 
                           n9784);
   U2960 : XNOR2_X1 port map( A => n565, B => n22875, ZN => Ciphertext(9));
   U2961 : OAI211_X1 port map( C1 => n24350, C2 => n22578, A => n1197, B => 
                           n22873, ZN => n565);
   U2962 : NAND2_X1 port map( A1 => n4165, A2 => n2815, ZN => n566);
   U2963 : NAND2_X1 port map( A1 => n17090, A2 => n17091, ZN => n567);
   U2964 : OR2_X1 port map( A1 => n6742, A2 => n6104, ZN => n568);
   U2965 : NAND2_X1 port map( A1 => n7280, A2 => n8512, ZN => n569);
   U2966 : OAI22_X1 port map( A1 => n21930, A2 => n22465, B1 => n22462, B2 => 
                           n22459, ZN => n570);
   U2967 : NAND2_X1 port map( A1 => n17032, A2 => n571, ZN => n18073);
   U2968 : NAND2_X1 port map( A1 => n2111, A2 => n572, ZN => n571);
   U2970 : NAND2_X1 port map( A1 => n574, A2 => n573, ZN => n2032);
   U2971 : INV_X1 port map( A => n24037, ZN => n573);
   U2972 : NAND2_X1 port map( A1 => n6921, A2 => n6920, ZN => n574);
   U2973 : NAND2_X1 port map( A1 => n25366, A2 => n25415, ZN => n2422);
   U2975 : OAI21_X2 port map( B1 => n16842, B2 => n17166, A => n16841, ZN => 
                           n18121);
   U2977 : NAND2_X1 port map( A1 => n10858, A2 => n10860, ZN => n10280);
   U2978 : NAND2_X1 port map( A1 => n5064, A2 => n9250, ZN => n10860);
   U2979 : OR2_X1 port map( A1 => n10099, A2 => n10100, ZN => n4302);
   U2981 : NAND2_X1 port map( A1 => n19599, A2 => n19598, ZN => n576);
   U2983 : NAND2_X1 port map( A1 => n579, A2 => n25449, ZN => n578);
   U2984 : INV_X1 port map( A => n16123, ZN => n579);
   U2985 : OAI211_X1 port map( C1 => n1231, C2 => n16957, A => n1230, B => 
                           n1229, ZN => n1228);
   U2986 : NAND3_X1 port map( A1 => n580, A2 => n1482, A3 => n2066, ZN => n1722
                           );
   U2988 : AND2_X1 port map( A1 => n339, A2 => n19883, ZN => n19916);
   U2989 : NAND2_X1 port map( A1 => n1551, A2 => n4842, ZN => n4841);
   U2990 : NAND2_X1 port map( A1 => n7666, A2 => n7665, ZN => n8534);
   U2991 : NAND2_X1 port map( A1 => n581, A2 => n2121, ZN => n16531);
   U2992 : NAND2_X1 port map( A1 => n16526, A2 => n17451, ZN => n581);
   U2993 : NAND2_X1 port map( A1 => n2223, A2 => n584, ZN => n7687);
   U2994 : NAND2_X1 port map( A1 => n9675, A2 => n9674, ZN => n1346);
   U2995 : AND2_X2 port map( A1 => n586, A2 => n585, ZN => n21985);
   U2996 : NAND2_X1 port map( A1 => n20302, A2 => n20301, ZN => n585);
   U2997 : NAND2_X1 port map( A1 => n20300, A2 => n20299, ZN => n586);
   U2998 : OAI21_X1 port map( B1 => n12526, B2 => n25337, A => n902, ZN => 
                           n11452);
   U3000 : AOI21_X1 port map( B1 => n20066, B2 => n20074, A => n588, ZN => n587
                           );
   U3002 : INV_X1 port map( A => n15584, ZN => n16105);
   U3003 : OR2_X1 port map( A1 => n6195, A2 => n6444, ZN => n640);
   U3004 : NAND2_X1 port map( A1 => n589, A2 => n4044, ZN => n15841);
   U3005 : NAND2_X1 port map( A1 => n692, A2 => n4045, ZN => n589);
   U3006 : OAI21_X1 port map( B1 => n429, B2 => n10060, A => n590, ZN => n10067
                           );
   U3007 : NAND2_X1 port map( A1 => n10060, A2 => n10061, ZN => n590);
   U3008 : OR2_X1 port map( A1 => n17093, A2 => n24410, ZN => n17687);
   U3009 : BUF_X2 port map( A => n6374, Z => n6904);
   U3010 : NAND3_X1 port map( A1 => n24468, A2 => n21840, A3 => n21822, ZN => 
                           n21296);
   U3014 : NAND2_X1 port map( A1 => n22403, A2 => n21885, ZN => n593);
   U3016 : NAND2_X1 port map( A1 => n6128, A2 => n6530, ZN => n6129);
   U3019 : AOI21_X1 port map( B1 => n907, B2 => n905, A => n142, ZN => n595);
   U3020 : NAND2_X1 port map( A1 => n6257, A2 => n6256, ZN => n2824);
   U3022 : NAND2_X1 port map( A1 => n4906, A2 => n13094, ZN => n598);
   U3024 : NAND2_X1 port map( A1 => n11410, A2 => n11409, ZN => n2117);
   U3025 : AND3_X2 port map( A1 => n599, A2 => n13649, A3 => n13650, ZN => 
                           n14104);
   U3027 : OAI211_X2 port map( C1 => n20567, C2 => n20566, A => n24530, B => 
                           n600, ZN => n21579);
   U3028 : NAND2_X1 port map( A1 => n20565, A2 => n20564, ZN => n600);
   U3029 : NAND2_X1 port map( A1 => n20502, A2 => n20501, ZN => n5424);
   U3030 : NAND2_X1 port map( A1 => n605, A2 => n602, ZN => n22854);
   U3032 : INV_X1 port map( A => n5421, ZN => n603);
   U3034 : NAND2_X1 port map( A1 => n22855, A2 => n24356, ZN => n605);
   U3035 : INV_X1 port map( A => n14382, ZN => n15620);
   U3036 : NAND3_X1 port map( A1 => n10253, A2 => n10730, A3 => n606, ZN => 
                           n10262);
   U3037 : OR2_X1 port map( A1 => n10255, A2 => n10254, ZN => n606);
   U3038 : NAND2_X1 port map( A1 => n10254, A2 => n10129, ZN => n10251);
   U3042 : AND2_X2 port map( A1 => n2048, A2 => n1471, ZN => n14327);
   U3046 : OAI21_X2 port map( B1 => n16653, B2 => n16652, A => n16651, ZN => 
                           n18239);
   U3047 : NAND2_X1 port map( A1 => n611, A2 => n610, ZN => n9839);
   U3048 : NAND2_X1 port map( A1 => n428, A2 => n8359, ZN => n610);
   U3049 : NAND2_X1 port map( A1 => n9838, A2 => n9837, ZN => n611);
   U3050 : NAND2_X1 port map( A1 => n10094, A2 => n9515, ZN => n9838);
   U3052 : XNOR2_X2 port map( A => n17511, B => n17512, ZN => n19297);
   U3053 : NAND2_X1 port map( A1 => n7887, A2 => n7883, ZN => n3130);
   U3054 : NAND2_X1 port map( A1 => n7882, A2 => n7585, ZN => n7887);
   U3057 : NAND2_X1 port map( A1 => n380, A2 => n16064, ZN => n613);
   U3058 : AND2_X1 port map( A1 => n22262, A2 => n1276, ZN => n22135);
   U3059 : NAND2_X1 port map( A1 => n615, A2 => n614, ZN => n19715);
   U3060 : NAND2_X1 port map( A1 => n20319, A2 => n19889, ZN => n614);
   U3061 : NOR2_X1 port map( A1 => n616, A2 => n7427, ZN => n7199);
   U3062 : NAND2_X1 port map( A1 => n7812, A2 => n9068, ZN => n616);
   U3063 : INV_X1 port map( A => n617, ZN => n16053);
   U3064 : NAND2_X1 port map( A1 => n24352, A2 => n15706, ZN => n617);
   U3066 : NOR2_X1 port map( A1 => n14131, A2 => n620, ZN => n14133);
   U3067 : NAND2_X1 port map( A1 => n619, A2 => n618, ZN => n12941);
   U3068 : NAND2_X1 port map( A1 => n5751, A2 => n14132, ZN => n618);
   U3070 : NOR2_X1 port map( A1 => n1508, A2 => n12597, ZN => n623);
   U3071 : NAND2_X1 port map( A1 => n12912, A2 => n1508, ZN => n624);
   U3073 : NAND2_X1 port map( A1 => n25424, A2 => n625, ZN => n7031);
   U3074 : NAND2_X1 port map( A1 => n625, A2 => n6104, ZN => n6005);
   U3075 : NAND3_X1 port map( A1 => n6593, A2 => n6592, A3 => n626, ZN => n6594
                           );
   U3076 : NAND2_X1 port map( A1 => n454, A2 => n7033, ZN => n626);
   U3077 : NOR2_X1 port map( A1 => n9398, A2 => n9365, ZN => n627);
   U3078 : AND2_X1 port map( A1 => n10136, A2 => n24026, ZN => n9201);
   U3079 : NAND2_X1 port map( A1 => n14853, A2 => n14852, ZN => n628);
   U3080 : NAND2_X1 port map( A1 => n21286, A2 => n629, ZN => n21288);
   U3081 : OAI211_X1 port map( C1 => n317, C2 => n23229, A => n23218, B => n630
                           , ZN => n629);
   U3082 : NAND2_X1 port map( A1 => n317, A2 => n23220, ZN => n630);
   U3083 : INV_X1 port map( A => n16311, ZN => n16012);
   U3084 : NAND2_X1 port map( A1 => n631, A2 => n16311, ZN => n633);
   U3085 : OAI21_X1 port map( B1 => n2173, B2 => n15198, A => n632, ZN => n631)
                           ;
   U3086 : NAND2_X1 port map( A1 => n15198, A2 => n16312, ZN => n632);
   U3089 : NAND2_X1 port map( A1 => n634, A2 => n633, ZN => n635);
   U3091 : OAI21_X1 port map( B1 => n17331, B2 => n635, A => n17335, ZN => 
                           n17339);
   U3092 : NOR2_X1 port map( A1 => n19972, A2 => n636, ZN => n19973);
   U3093 : OAI21_X1 port map( B1 => n20530, B2 => n636, A => n2852, ZN => 
                           n18886);
   U3094 : INV_X1 port map( A => n20289, ZN => n636);
   U3095 : NAND2_X1 port map( A1 => n637, A2 => n6196, ZN => n4726);
   U3096 : NAND2_X1 port map( A1 => n6448, A2 => n637, ZN => n4878);
   U3097 : NAND2_X1 port map( A1 => n640, A2 => n6188, ZN => n637);
   U3098 : XNOR2_X1 port map( A => n25390, B => n447, ZN => n18241);
   U3099 : XNOR2_X1 port map( A => n25390, B => n452, ZN => n16635);
   U3100 : XNOR2_X1 port map( A => n17873, B => n445, ZN => n17644);
   U3101 : XNOR2_X1 port map( A => n25390, B => n449, ZN => n18125);
   U3102 : NOR2_X1 port map( A1 => n372, A2 => n17053, ZN => n4298);
   U3104 : NAND2_X1 port map( A1 => n9358, A2 => n9357, ZN => n3324);
   U3106 : NAND2_X1 port map( A1 => n24398, A2 => n24585, ZN => n16609);
   U3109 : NAND2_X1 port map( A1 => n25408, A2 => n12490, ZN => n642);
   U3111 : NAND2_X1 port map( A1 => n12534, A2 => n12535, ZN => n12533);
   U3112 : NAND2_X1 port map( A1 => n645, A2 => n376, ZN => n644);
   U3115 : NAND2_X1 port map( A1 => n994, A2 => n16266, ZN => n646);
   U3117 : NAND2_X1 port map( A1 => n10594, A2 => n10505, ZN => n10930);
   U3120 : NAND3_X1 port map( A1 => n10688, A2 => n10687, A3 => n10686, ZN => 
                           n10689);
   U3121 : OR2_X1 port map( A1 => n17299, A2 => n17297, ZN => n16702);
   U3122 : OR2_X1 port map( A1 => n22782, A2 => n24406, ZN => n22365);
   U3123 : NAND3_X1 port map( A1 => n1198, A2 => n22872, A3 => n22578, ZN => 
                           n1197);
   U3127 : NAND3_X2 port map( A1 => n15608, A2 => n879, A3 => n880, ZN => 
                           n17068);
   U3130 : NAND2_X1 port map( A1 => n16069, A2 => n4105, ZN => n649);
   U3131 : NAND2_X1 port map( A1 => n651, A2 => n650, ZN => n21938);
   U3132 : NAND2_X1 port map( A1 => n21935, A2 => n326, ZN => n651);
   U3133 : XNOR2_X1 port map( A => n15222, B => n15221, ZN => n16192);
   U3134 : NOR2_X1 port map( A1 => n13486, A2 => n24462, ZN => n652);
   U3135 : NAND3_X1 port map( A1 => n10547, A2 => n10705, A3 => n10702, ZN => 
                           n10551);
   U3139 : AOI22_X1 port map( A1 => n12866, A2 => n12865, B1 => n1513, B2 => 
                           n13114, ZN => n4798);
   U3140 : NAND3_X1 port map( A1 => n9456, A2 => n9455, A3 => n9887, ZN => n957
                           );
   U3142 : NAND2_X1 port map( A1 => n657, A2 => n438, ZN => n656);
   U3143 : NAND2_X1 port map( A1 => n6439, A2 => n6438, ZN => n657);
   U3144 : NAND2_X1 port map( A1 => n6440, A2 => n6174, ZN => n658);
   U3145 : NAND3_X2 port map( A1 => n2943, A2 => n7649, A3 => n989, ZN => n9043
                           );
   U3146 : XNOR2_X1 port map( A => n659, B => n5598, ZN => Ciphertext(136));
   U3147 : OAI211_X1 port map( C1 => n23718, C2 => n3283, A => n3280, B => 
                           n23717, ZN => n659);
   U3148 : NOR2_X2 port map( A1 => n11252, A2 => n661, ZN => n14294);
   U3149 : OAI22_X1 port map( A1 => n12987, A2 => n13220, B1 => n4652, B2 => 
                           n12767, ZN => n661);
   U3150 : NAND2_X1 port map( A1 => n374, A2 => n662, ZN => n17044);
   U3151 : NAND2_X1 port map( A1 => n24903, A2 => n23303, ZN => n23295);
   U3152 : XNOR2_X1 port map( A => n664, B => n23302, ZN => Ciphertext(57));
   U3153 : NAND3_X1 port map( A1 => n13506, A2 => n13507, A3 => n13505, ZN => 
                           n13508);
   U3154 : NAND3_X1 port map( A1 => n4597, A2 => n4600, A3 => n13437, ZN => 
                           n2821);
   U3155 : XNOR2_X2 port map( A => n5822, B => Key(146), ZN => n6377);
   U3156 : OAI211_X2 port map( C1 => n17325, C2 => n17326, A => n207, B => n206
                           , ZN => n18447);
   U3157 : XNOR2_X1 port map( A => n11768, B => n11764, ZN => n667);
   U3159 : NAND2_X1 port map( A1 => n6674, A2 => n6675, ZN => n668);
   U3160 : NAND2_X1 port map( A1 => n14584, A2 => n213, ZN => n14585);
   U3162 : XNOR2_X1 port map( A => n18152, B => n18147, ZN => n670);
   U3163 : OAI211_X1 port map( C1 => n1771, C2 => n13962, A => n671, B => n4293
                           , ZN => n1770);
   U3164 : NAND2_X1 port map( A1 => n13962, A2 => n13963, ZN => n671);
   U3165 : AND2_X2 port map( A1 => n3744, A2 => n15768, ZN => n16809);
   U3166 : NAND3_X1 port map( A1 => n2003, A2 => n2002, A3 => n672, ZN => 
                           n14976);
   U3168 : NOR2_X1 port map( A1 => n16851, A2 => n1653, ZN => n16847);
   U3169 : NAND3_X1 port map( A1 => n674, A2 => n6494, A3 => n6489, ZN => n6492
                           );
   U3170 : NAND2_X1 port map( A1 => n6487, A2 => n6488, ZN => n674);
   U3171 : NAND3_X1 port map( A1 => n675, A2 => n9884, A3 => n9563, ZN => n9891
                           );
   U3172 : NAND2_X1 port map( A1 => n9883, A2 => n9882, ZN => n675);
   U3173 : OAI211_X1 port map( C1 => n7634, C2 => n7918, A => n312, B => n920, 
                           ZN => n1280);
   U3174 : NAND2_X1 port map( A1 => n7923, A2 => n5607, ZN => n1088);
   U3175 : NAND2_X1 port map( A1 => n12833, A2 => n5645, ZN => n12850);
   U3176 : NAND2_X1 port map( A1 => n9419, A2 => n9613, ZN => n9972);
   U3177 : NAND2_X1 port map( A1 => n1345, A2 => n270, ZN => n2223);
   U3179 : AND2_X1 port map( A1 => n2677, A2 => n710, ZN => n5259);
   U3180 : NAND2_X1 port map( A1 => n676, A2 => n13055, ZN => n13059);
   U3181 : NOR2_X1 port map( A1 => n409, A2 => n13057, ZN => n676);
   U3182 : OR2_X1 port map( A1 => n1248, A2 => n22359, ZN => n782);
   U3183 : NAND2_X1 port map( A1 => n2939, A2 => n401, ZN => n2938);
   U3184 : NAND2_X1 port map( A1 => n1962, A2 => n1961, ZN => n1959);
   U3185 : OAI21_X1 port map( B1 => n11085, B2 => n418, A => n678, ZN => n10894
                           );
   U3186 : NAND2_X1 port map( A1 => n11085, A2 => n10890, ZN => n678);
   U3187 : XNOR2_X1 port map( A => n14827, B => n15446, ZN => n14430);
   U3188 : INV_X1 port map( A => n16572, ZN => n17116);
   U3189 : OAI211_X1 port map( C1 => n19070, C2 => n19612, A => n19069, B => 
                           n19068, ZN => n1155);
   U3192 : NAND3_X1 port map( A1 => n7841, A2 => n8370, A3 => n7843, ZN => 
                           n7842);
   U3194 : NAND2_X1 port map( A1 => n680, A2 => n4753, ZN => n7578);
   U3195 : NAND2_X1 port map( A1 => n4751, A2 => n4752, ZN => n680);
   U3196 : NAND2_X1 port map( A1 => n10684, A2 => n10363, ZN => n3934);
   U3197 : NAND2_X1 port map( A1 => n6405, A2 => n6404, ZN => n1558);
   U3199 : NAND2_X1 port map( A1 => n4806, A2 => n4807, ZN => n693);
   U3200 : NAND2_X1 port map( A1 => n2090, A2 => n16109, ZN => n682);
   U3201 : NAND2_X1 port map( A1 => n4689, A2 => n379, ZN => n683);
   U3204 : OAI22_X1 port map( A1 => n442, A2 => n249, B1 => n7021, B2 => n7026,
                           ZN => n6638);
   U3205 : NAND2_X1 port map( A1 => n13548, A2 => n13551, ZN => n684);
   U3207 : OAI21_X1 port map( B1 => n707, B2 => n16170, A => n706, ZN => n15960
                           );
   U3208 : NAND3_X1 port map( A1 => n685, A2 => n12461, A3 => n12482, ZN => 
                           n3454);
   U3209 : INV_X1 port map( A => n12709, ZN => n685);
   U3210 : OAI22_X1 port map( A1 => n16031, A2 => n24403, B1 => n16276, B2 => 
                           n16274, ZN => n16032);
   U3212 : NAND2_X1 port map( A1 => n3050, A2 => n4369, ZN => n7421);
   U3213 : NAND2_X1 port map( A1 => n16534, A2 => n16533, ZN => n686);
   U3216 : NAND2_X1 port map( A1 => n6380, A2 => n6379, ZN => n4641);
   U3217 : XNOR2_X1 port map( A => n11796, B => n12138, ZN => n11469);
   U3220 : NAND2_X1 port map( A1 => n16973, A2 => n17336, ZN => n16726);
   U3221 : NAND2_X1 port map( A1 => n25462, A2 => n25022, ZN => n21146);
   U3224 : NAND2_X1 port map( A1 => n19611, A2 => n2764, ZN => n1590);
   U3225 : NAND2_X1 port map( A1 => n13417, A2 => n24503, ZN => n689);
   U3226 : NAND2_X1 port map( A1 => n25278, A2 => n14099, ZN => n690);
   U3229 : NAND3_X1 port map( A1 => n693, A2 => n16686, A3 => n3723, ZN => 
                           n17248);
   U3230 : NAND2_X1 port map( A1 => n24339, A2 => n324, ZN => n23389);
   U3232 : NAND2_X1 port map( A1 => n731, A2 => n800, ZN => n7214);
   U3233 : NAND3_X1 port map( A1 => n3169, A2 => n14748, A3 => n16762, ZN => 
                           n829);
   U3235 : AOI21_X1 port map( B1 => n22848, B2 => n21709, A => n22907, ZN => 
                           n695);
   U3236 : OR2_X2 port map( A1 => n722, A2 => n2449, ZN => n12414);
   U3238 : NAND2_X1 port map( A1 => n5633, A2 => n19191, ZN => n5632);
   U3239 : NAND2_X1 port map( A1 => n18923, A2 => n696, ZN => n17011);
   U3240 : NAND2_X1 port map( A1 => n14180, A2 => n14178, ZN => n13771);
   U3241 : INV_X1 port map( A => n697, ZN => n22269);
   U3242 : OAI22_X1 port map( A1 => n22268, A2 => n22267, B1 => n22266, B2 => 
                           n25381, ZN => n697);
   U3245 : NAND3_X1 port map( A1 => n822, A2 => n821, A3 => n699, ZN => n698);
   U3247 : NAND2_X1 port map( A1 => n15314, A2 => n17342, ZN => n16778);
   U3249 : NAND2_X1 port map( A1 => n6037, A2 => n6503, ZN => n703);
   U3250 : OAI21_X1 port map( B1 => n13840, B2 => n397, A => n704, ZN => n13842
                           );
   U3251 : NAND2_X1 port map( A1 => n13840, A2 => n13837, ZN => n704);
   U3252 : NAND3_X1 port map( A1 => n13189, A2 => n3957, A3 => n13190, ZN => 
                           n14108);
   U3253 : NAND3_X1 port map( A1 => n9657, A2 => n9996, A3 => n9658, ZN => n867
                           );
   U3254 : OR2_X1 port map( A1 => n16266, A2 => n16268, ZN => n992);
   U3255 : AND2_X1 port map( A1 => n14290, A2 => n13907, ZN => n11454);
   U3256 : OR3_X1 port map( A1 => n19393, A2 => n18788, A3 => n24407, ZN => 
                           n18789);
   U3257 : OAI21_X1 port map( B1 => n6329, B2 => n4621, A => n6471, ZN => n1078
                           );
   U3258 : OAI21_X1 port map( B1 => n406, B2 => n25430, A => n705, ZN => n12875
                           );
   U3259 : NAND2_X1 port map( A1 => n13352, A2 => n13353, ZN => n705);
   U3262 : NAND2_X1 port map( A1 => n6049, A2 => n6623, ZN => n6624);
   U3263 : NAND2_X1 port map( A1 => n1918, A2 => n11208, ZN => n11211);
   U3265 : NAND2_X1 port map( A1 => n6425, A2 => n198, ZN => n2542);
   U3267 : NAND2_X1 port map( A1 => n9979, A2 => n712, ZN => n711);
   U3268 : INV_X1 port map( A => n713, ZN => n712);
   U3269 : OAI21_X1 port map( B1 => n9429, B2 => n9981, A => n9980, ZN => n713)
                           ;
   U3271 : NAND3_X1 port map( A1 => n10156, A2 => n25206, A3 => n10120, ZN => 
                           n2254);
   U3272 : NAND3_X1 port map( A1 => n5277, A2 => n25007, A3 => n5278, ZN => 
                           n5272);
   U3273 : INV_X1 port map( A => n716, ZN => Ciphertext(116));
   U3274 : OAI211_X1 port map( C1 => n21952, C2 => n21951, A => n21949, B => 
                           n21950, ZN => n716);
   U3275 : NAND2_X1 port map( A1 => n7212, A2 => n8530, ZN => n800);
   U3276 : NAND3_X1 port map( A1 => n346, A2 => n20486, A3 => n19634, ZN => 
                           n19638);
   U3277 : NAND2_X1 port map( A1 => n17255, A2 => n16561, ZN => n17257);
   U3279 : NAND2_X1 port map( A1 => n7720, A2 => n7719, ZN => n8730);
   U3280 : NAND3_X1 port map( A1 => n719, A2 => n1465, A3 => n718, ZN => n23956
                           );
   U3281 : NAND2_X1 port map( A1 => n23953, A2 => n23969, ZN => n718);
   U3282 : NAND2_X1 port map( A1 => n23954, A2 => n23955, ZN => n719);
   U3283 : OAI211_X2 port map( C1 => n3971, C2 => n13162, A => n3970, B => 
                           n3969, ZN => n1355);
   U3284 : NAND2_X1 port map( A1 => n19190, A2 => n20511, ZN => n837);
   U3286 : OR2_X2 port map( A1 => n720, A2 => n4941, ZN => n3725);
   U3288 : NAND2_X1 port map( A1 => n721, A2 => n23011, ZN => n23493);
   U3289 : NAND2_X1 port map( A1 => n23480, A2 => n2710, ZN => n721);
   U3290 : AOI21_X1 port map( B1 => n10657, B2 => n10656, A => n10661, ZN => 
                           n722);
   U3291 : AOI21_X1 port map( B1 => n10727, B2 => n10726, A => n10868, ZN => 
                           n1900);
   U3292 : NAND2_X1 port map( A1 => n10286, A2 => n1658, ZN => n10727);
   U3295 : XNOR2_X1 port map( A => n14979, B => n14980, ZN => n14981);
   U3296 : OAI211_X2 port map( C1 => n13526, C2 => n13527, A => n3329, B => 
                           n3331, ZN => n14979);
   U3297 : NAND2_X1 port map( A1 => n12862, A2 => n725, ZN => n13871);
   U3298 : NAND2_X1 port map( A1 => n12858, A2 => n12863, ZN => n725);
   U3300 : NAND2_X1 port map( A1 => n13602, A2 => n14317, ZN => n13603);
   U3301 : NAND2_X1 port map( A1 => n17304, A2 => n17305, ZN => n1244);
   U3302 : NAND2_X1 port map( A1 => n14302, A2 => n14306, ZN => n13889);
   U3303 : OAI21_X1 port map( B1 => n6718, B2 => n24051, A => n24500, ZN => 
                           n6237);
   U3305 : NAND2_X1 port map( A1 => n313, A2 => n6893, ZN => n6816);
   U3306 : XNOR2_X2 port map( A => n5826, B => Key(137), ZN => n6893);
   U3307 : NAND2_X1 port map( A1 => n20317, A2 => n340, ZN => n4960);
   U3308 : NAND2_X1 port map( A1 => n17503, A2 => n17502, ZN => n727);
   U3309 : INV_X1 port map( A => n2229, ZN => n728);
   U3313 : NAND3_X1 port map( A1 => n2325, A2 => n17227, A3 => n16954, ZN => 
                           n4974);
   U3314 : NAND2_X1 port map( A1 => n798, A2 => n7665, ZN => n731);
   U3316 : NAND2_X1 port map( A1 => n732, A2 => n19162, ZN => n1979);
   U3317 : NAND2_X1 port map( A1 => n3726, A2 => n19163, ZN => n732);
   U3318 : NAND2_X1 port map( A1 => n13212, A2 => n13211, ZN => n13005);
   U3319 : NAND2_X1 port map( A1 => n733, A2 => n16734, ZN => n16735);
   U3320 : NAND2_X1 port map( A1 => n16733, A2 => n16732, ZN => n733);
   U3321 : NAND2_X1 port map( A1 => n6904, A2 => n6089, ZN => n6090);
   U3323 : NAND3_X1 port map( A1 => n1058, A2 => n2878, A3 => n11302, ZN => 
                           n734);
   U3324 : OAI21_X1 port map( B1 => n10650, B2 => n10651, A => n735, ZN => 
                           n10652);
   U3325 : NAND3_X2 port map( A1 => n737, A2 => n736, A3 => n8004, ZN => n8965)
                           ;
   U3326 : NAND2_X1 port map( A1 => n7756, A2 => n7755, ZN => n737);
   U3331 : NAND4_X1 port map( A1 => n741, A2 => n14367, A3 => n14366, A4 => 
                           n740, ZN => n14368);
   U3332 : NAND2_X1 port map( A1 => n14363, A2 => n5526, ZN => n740);
   U3333 : NAND2_X1 port map( A1 => n14365, A2 => n14364, ZN => n741);
   U3334 : NAND2_X1 port map( A1 => n19395, A2 => n19162, ZN => n18790);
   U3338 : NAND3_X1 port map( A1 => n4215, A2 => n21366, A3 => n21365, ZN => 
                           Ciphertext(160));
   U3339 : NAND2_X1 port map( A1 => n16347, A2 => n25441, ZN => n2702);
   U3340 : NAND2_X1 port map( A1 => n744, A2 => n743, ZN => n1832);
   U3341 : AOI21_X1 port map( B1 => n24080, B2 => n15822, A => n16597, ZN => 
                           n743);
   U3342 : NAND2_X1 port map( A1 => n16595, A2 => n24467, ZN => n744);
   U3343 : NAND3_X1 port map( A1 => n10134, A2 => n10141, A3 => n10138, ZN => 
                           n9370);
   U3346 : INV_X1 port map( A => n16398, ZN => n746);
   U3348 : NAND2_X1 port map( A1 => n3937, A2 => n22461, ZN => n747);
   U3349 : NAND2_X1 port map( A1 => n24253, A2 => n24592, ZN => n6015);
   U3352 : OR2_X1 port map( A1 => n16546, A2 => n17068, ZN => n1071);
   U3353 : NAND2_X1 port map( A1 => n24973, A2 => n749, ZN => n2303);
   U3355 : NAND3_X2 port map( A1 => n751, A2 => n16617, A3 => n752, ZN => 
                           n18431);
   U3356 : NAND2_X1 port map( A1 => n3377, A2 => n469, ZN => n752);
   U3357 : OAI21_X1 port map( B1 => n19817, B2 => n754, A => n753, ZN => n19512
                           );
   U3358 : NAND2_X1 port map( A1 => n19817, A2 => n1344, ZN => n753);
   U3360 : NAND2_X1 port map( A1 => n757, A2 => n756, ZN => n15718);
   U3361 : NAND2_X1 port map( A1 => n24981, A2 => n15951, ZN => n756);
   U3362 : NAND3_X1 port map( A1 => n10307, A2 => n759, A3 => n758, ZN => 
                           n11776);
   U3363 : OAI21_X1 port map( B1 => n10305, B2 => n10306, A => n4998, ZN => 
                           n759);
   U3366 : NAND2_X1 port map( A1 => n762, A2 => n19543, ZN => n3665);
   U3367 : NAND2_X1 port map( A1 => n2879, A2 => n7010, ZN => n764);
   U3369 : NAND2_X1 port map( A1 => n766, A2 => n437, ZN => n1192);
   U3370 : NAND2_X1 port map( A1 => n7235, A2 => n7961, ZN => n766);
   U3372 : NAND3_X1 port map( A1 => n6153, A2 => n6277, A3 => n440, ZN => n767)
                           ;
   U3374 : NAND2_X1 port map( A1 => n1160, A2 => n1161, ZN => n1159);
   U3375 : NAND2_X1 port map( A1 => n5744, A2 => n1689, ZN => n11133);
   U3376 : NOR2_X1 port map( A1 => n420, A2 => n10838, ZN => n5744);
   U3377 : NAND2_X1 port map( A1 => n12597, A2 => n12824, ZN => n12690);
   U3378 : NAND2_X1 port map( A1 => n770, A2 => n769, ZN => n14080);
   U3380 : NAND2_X1 port map( A1 => n14076, A2 => n396, ZN => n770);
   U3381 : NAND3_X1 port map( A1 => n771, A2 => n20370, A3 => n349, ZN => n3430
                           );
   U3382 : NAND2_X1 port map( A1 => n6556, A2 => n6697, ZN => n1961);
   U3383 : NAND2_X1 port map( A1 => n19581, A2 => n19579, ZN => n18880);
   U3385 : OAI22_X1 port map( A1 => n3211, A2 => n3212, B1 => n3210, B2 => 
                           n22972, ZN => n772);
   U3386 : AOI21_X2 port map( B1 => n19440, B2 => n3986, A => n19439, ZN => 
                           n20588);
   U3388 : NAND2_X1 port map( A1 => n3116, A2 => n3072, ZN => n9254);
   U3391 : AOI22_X1 port map( A1 => n4513, A2 => n23645, B1 => n24320, B2 => 
                           n23652, ZN => n22153);
   U3396 : NOR2_X1 port map( A1 => n1201, A2 => n1200, ZN => n4447);
   U3397 : NOR2_X1 port map( A1 => n5472, A2 => n4923, ZN => n898);
   U3398 : XNOR2_X1 port map( A => n15342, B => n15238, ZN => n15239);
   U3401 : NAND2_X1 port map( A1 => n7431, A2 => n775, ZN => n8339);
   U3404 : NAND2_X1 port map( A1 => n7057, A2 => n9067, ZN => n3249);
   U3405 : NAND3_X2 port map( A1 => n3171, A2 => n2078, A3 => n6340, ZN => 
                           n9067);
   U3406 : AOI21_X1 port map( B1 => n777, B2 => n9560, A => n9559, ZN => n9561)
                           ;
   U3407 : NAND2_X1 port map( A1 => n1365, A2 => n16073, ZN => n16074);
   U3408 : NAND2_X1 port map( A1 => n778, A2 => n14178, ZN => n4593);
   U3409 : NAND2_X1 port map( A1 => n14181, A2 => n13796, ZN => n778);
   U3412 : NAND4_X1 port map( A1 => n23872, A2 => n3077, A3 => n3078, A4 => 
                           n23871, ZN => n23874);
   U3413 : XNOR2_X1 port map( A => n781, B => n21080, ZN => n21082);
   U3414 : XNOR2_X1 port map( A => n21081, B => n21429, ZN => n781);
   U3415 : NAND2_X1 port map( A1 => n7211, A2 => n7662, ZN => n6548);
   U3416 : NAND2_X1 port map( A1 => n9589, A2 => n9588, ZN => n3551);
   U3419 : NAND2_X1 port map( A1 => n14320, A2 => n13871, ZN => n14459);
   U3421 : NAND2_X1 port map( A1 => n22671, A2 => n22784, ZN => n22672);
   U3428 : NAND3_X1 port map( A1 => n23587, A2 => n23588, A3 => n23586, ZN => 
                           n23590);
   U3429 : NAND2_X1 port map( A1 => n10117, A2 => n784, ZN => n9532);
   U3430 : NAND2_X1 port map( A1 => n9530, A2 => n9531, ZN => n784);
   U3432 : INV_X1 port map( A => n17734, ZN => n4934);
   U3433 : NAND2_X1 port map( A1 => n1086, A2 => n1087, ZN => n12423);
   U3434 : NAND2_X1 port map( A1 => n13177, A2 => n12506, ZN => n13174);
   U3435 : OAI211_X2 port map( C1 => n3656, C2 => n20165, A => n19950, B => 
                           n19949, ZN => n21713);
   U3438 : OR2_X1 port map( A1 => n10065, A2 => n10064, ZN => n787);
   U3439 : OAI21_X1 port map( B1 => n4083, B2 => n5158, A => n4082, ZN => n788)
                           ;
   U3440 : NOR2_X2 port map( A1 => n19020, A2 => n789, ZN => n21639);
   U3441 : OAI22_X1 port map( A1 => n20532, A2 => n20536, B1 => n19019, B2 => 
                           n20447, ZN => n789);
   U3443 : XNOR2_X1 port map( A => n4687, B => n4688, ZN => n801);
   U3444 : NAND4_X1 port map( A1 => n3425, A2 => n3426, A3 => n13964, A4 => 
                           n3427, ZN => n790);
   U3446 : NAND3_X1 port map( A1 => n6464, A2 => n6459, A3 => n6455, ZN => 
                           n2078);
   U3447 : NAND2_X1 port map( A1 => n3815, A2 => n16603, ZN => n3816);
   U3448 : NAND2_X1 port map( A1 => n2028, A2 => n2027, ZN => n4511);
   U3450 : XNOR2_X1 port map( A => n792, B => n23183, ZN => Ciphertext(29));
   U3451 : OAI22_X1 port map( A1 => n23180, A2 => n23179, B1 => n23182, B2 => 
                           n23181, ZN => n792);
   U3452 : NAND2_X1 port map( A1 => n1145, A2 => n23688, ZN => n1144);
   U3453 : INV_X1 port map( A => n933, ZN => n7710);
   U3454 : NAND2_X1 port map( A1 => n7865, A2 => n7862, ZN => n933);
   U3455 : NAND3_X1 port map( A1 => n10729, A2 => n10482, A3 => n10481, ZN => 
                           n1178);
   U3456 : NAND3_X1 port map( A1 => n6938, A2 => n6281, A3 => n793, ZN => n5911
                           );
   U3457 : OR2_X1 port map( A1 => n6944, A2 => n5910, ZN => n793);
   U3458 : NAND2_X1 port map( A1 => n5910, A2 => n5887, ZN => n6938);
   U3461 : XNOR2_X2 port map( A => n796, B => n838, ZN => n16274);
   U3462 : OR2_X1 port map( A1 => n16334, A2 => n25092, ZN => n981);
   U3463 : NAND2_X1 port map( A1 => n14021, A2 => n14022, ZN => n13540);
   U3464 : NAND2_X1 port map( A1 => n22762, A2 => n23294, ZN => n22761);
   U3467 : NAND2_X1 port map( A1 => n4336, A2 => n13067, ZN => n4340);
   U3471 : XNOR2_X1 port map( A => n17678, B => n17679, ZN => n797);
   U3473 : OAI21_X1 port map( B1 => n8528, B2 => n269, A => n799, ZN => n798);
   U3474 : NAND2_X1 port map( A1 => n7211, A2 => n8531, ZN => n799);
   U3476 : NAND2_X1 port map( A1 => n7933, A2 => n7932, ZN => n2165);
   U3477 : NAND2_X1 port map( A1 => n7163, A2 => n7923, ZN => n7933);
   U3478 : NAND3_X2 port map( A1 => n8352, A2 => n3708, A3 => n8351, ZN => 
                           n8952);
   U3480 : AOI21_X1 port map( B1 => n3764, B2 => n3765, A => n16406, ZN => n802
                           );
   U3481 : NAND2_X1 port map( A1 => n949, A2 => n6097, ZN => n8005);
   U3483 : INV_X1 port map( A => n16997, ZN => n17000);
   U3484 : NAND2_X1 port map( A1 => n17574, A2 => n17368, ZN => n16997);
   U3487 : XNOR2_X1 port map( A => n804, B => n14470, ZN => n14471);
   U3488 : XNOR2_X1 port map( A => n14469, B => n14675, ZN => n804);
   U3490 : INV_X1 port map( A => n7682, ZN => n806);
   U3495 : NOR2_X1 port map( A1 => n808, A2 => n19255, ZN => n19073);
   U3496 : NAND2_X1 port map( A1 => n21841, A2 => n22255, ZN => n809);
   U3497 : AOI22_X2 port map( A1 => n14007, A2 => n14006, B1 => n14005, B2 => 
                           n14004, ZN => n14980);
   U3500 : NAND2_X1 port map( A1 => n16902, A2 => n16539, ZN => n17473);
   U3501 : NAND2_X1 port map( A1 => n1116, A2 => n1118, ZN => n5906);
   U3502 : NAND3_X1 port map( A1 => n13462, A2 => n814, A3 => n813, ZN => 
                           n14676);
   U3503 : NAND2_X1 port map( A1 => n4921, A2 => n13959, ZN => n814);
   U3504 : NAND2_X1 port map( A1 => n17012, A2 => n4004, ZN => n3516);
   U3505 : INV_X1 port map( A => n7920, ZN => n1282);
   U3507 : NAND2_X1 port map( A1 => n20912, A2 => n815, ZN => n21736);
   U3508 : NAND3_X1 port map( A1 => n817, A2 => n347, A3 => n816, ZN => n815);
   U3509 : NAND2_X1 port map( A1 => n20911, A2 => n346, ZN => n816);
   U3510 : NAND2_X1 port map( A1 => n20910, A2 => n20909, ZN => n817);
   U3511 : NAND2_X1 port map( A1 => n21888, A2 => n22265, ZN => n22266);
   U3513 : NAND3_X1 port map( A1 => n819, A2 => n4188, A3 => n4187, ZN => 
                           Ciphertext(166));
   U3514 : OAI21_X1 port map( B1 => n4193, B2 => n4192, A => n23868, ZN => n819
                           );
   U3515 : XNOR2_X1 port map( A => n820, B => n19946, ZN => n19966);
   U3516 : XNOR2_X1 port map( A => n19955, B => n24899, ZN => n820);
   U3517 : NOR2_X2 port map( A1 => n1312, A2 => n20037, ZN => n23857);
   U3519 : NAND2_X1 port map( A1 => n14507, A2 => n24556, ZN => n13977);
   U3520 : NAND2_X1 port map( A1 => n9850, A2 => n9849, ZN => n821);
   U3521 : NAND2_X1 port map( A1 => n9384, A2 => n9592, ZN => n822);
   U3522 : INV_X1 port map( A => n17486, ZN => n17093);
   U3524 : NAND2_X1 port map( A1 => n14327, A2 => n14328, ZN => n14329);
   U3525 : NAND3_X1 port map( A1 => n1589, A2 => n4235, A3 => n4237, ZN => 
                           n4229);
   U3526 : NAND2_X1 port map( A1 => n4230, A2 => n23200, ZN => n1589);
   U3528 : INV_X1 port map( A => n2632, ZN => n12829);
   U3529 : NAND2_X1 port map( A1 => n13265, A2 => n2632, ZN => n2631);
   U3530 : NAND2_X1 port map( A1 => n4653, A2 => n17641, ZN => n19917);
   U3531 : XNOR2_X1 port map( A => n823, B => n18492, ZN => n18494);
   U3532 : XNOR2_X1 port map( A => n18490, B => n18491, ZN => n823);
   U3533 : OAI211_X1 port map( C1 => n22537, C2 => n23265, A => n825, B => n824
                           , ZN => n22538);
   U3534 : NAND2_X1 port map( A1 => n22535, A2 => n23265, ZN => n824);
   U3535 : NAND2_X1 port map( A1 => n22536, A2 => n23281, ZN => n825);
   U3536 : NAND2_X1 port map( A1 => n829, A2 => n826, ZN => n18251);
   U3537 : NAND2_X1 port map( A1 => n828, A2 => n827, ZN => n826);
   U3538 : INV_X1 port map( A => n17248, ZN => n827);
   U3539 : AOI22_X1 port map( A1 => n6558, A2 => n830, B1 => n6415, B2 => n6560
                           , ZN => n6417);
   U3540 : NAND2_X1 port map( A1 => n6693, A2 => n6695, ZN => n830);
   U3541 : XNOR2_X1 port map( A => n831, B => n20505, ZN => n20521);
   U3542 : XNOR2_X1 port map( A => n20504, B => n21600, ZN => n831);
   U3543 : NAND3_X1 port map( A1 => n212, A2 => n4903, A3 => n832, ZN => n2760)
                           ;
   U3544 : NAND2_X1 port map( A1 => n22530, A2 => n23860, ZN => n832);
   U3546 : NAND2_X1 port map( A1 => n22966, A2 => n24411, ZN => n833);
   U3547 : OAI22_X1 port map( A1 => n834, A2 => n14063, B1 => n13847, B2 => 
                           n13845, ZN => n13849);
   U3548 : NOR2_X1 port map( A1 => n13844, A2 => n13843, ZN => n834);
   U3549 : AOI22_X2 port map( A1 => n13310, A2 => n13309, B1 => n13312, B2 => 
                           n13311, ZN => n13924);
   U3552 : NAND3_X1 port map( A1 => n6051, A2 => n6746, A3 => n453, ZN => n6747
                           );
   U3553 : XNOR2_X2 port map( A => n5831, B => Key(142), ZN => n6795);
   U3554 : NAND2_X1 port map( A1 => n1774, A2 => n12665, ZN => n1773);
   U3555 : NOR2_X2 port map( A1 => n837, A2 => n19193, ZN => n21514);
   U3557 : XNOR2_X1 port map( A => n14891, B => n14893, ZN => n838);
   U3558 : NAND3_X1 port map( A1 => n22461, A2 => n22462, A3 => n3845, ZN => 
                           n4339);
   U3559 : NAND3_X1 port map( A1 => n13185, A2 => n24640, A3 => n12740, ZN => 
                           n13105);
   U3560 : NAND2_X1 port map( A1 => n5451, A2 => n4621, ZN => n4620);
   U3561 : NAND2_X1 port map( A1 => n1599, A2 => n1793, ZN => n20376);
   U3562 : NAND2_X1 port map( A1 => n6776, A2 => n6292, ZN => n6481);
   U3563 : AND2_X2 port map( A1 => n10674, A2 => n1453, ZN => n11163);
   U3565 : NOR2_X1 port map( A1 => n1294, A2 => n1295, ZN => n839);
   U3566 : NAND2_X1 port map( A1 => n19686, A2 => n20149, ZN => n19687);
   U3567 : NAND2_X1 port map( A1 => n23690, A2 => n2305, ZN => n22998);
   U3569 : NAND3_X2 port map( A1 => n4619, A2 => n6316, A3 => n6317, ZN => 
                           n7865);
   U3570 : OAI21_X1 port map( B1 => n22109, B2 => n22929, A => n22108, ZN => 
                           n840);
   U3571 : NAND2_X1 port map( A1 => n1530, A2 => n841, ZN => n8088);
   U3572 : NAND2_X1 port map( A1 => n3352, A2 => n842, ZN => n841);
   U3573 : XNOR2_X1 port map( A => n843, B => n23564, ZN => Ciphertext(112));
   U3574 : OAI211_X1 port map( C1 => n23563, C2 => n23562, A => n23560, B => 
                           n23561, ZN => n843);
   U3576 : NAND2_X1 port map( A1 => n12633, A2 => n12206, ZN => n5470);
   U3580 : OAI21_X2 port map( B1 => n25036, B2 => n14083, A => n12574, ZN => 
                           n14857);
   U3581 : NAND3_X1 port map( A1 => n13206, A2 => n1335, A3 => n13207, ZN => 
                           n1725);
   U3583 : OAI22_X1 port map( A1 => n845, A2 => n20186, B1 => n20043, B2 => 
                           n20191, ZN => n20044);
   U3584 : NAND2_X1 port map( A1 => n20041, A2 => n20042, ZN => n845);
   U3585 : NAND2_X1 port map( A1 => n2346, A2 => n19592, ZN => n19589);
   U3588 : NAND2_X1 port map( A1 => n9929, A2 => n9934, ZN => n847);
   U3589 : NAND2_X1 port map( A1 => n7838, A2 => n25217, ZN => n848);
   U3592 : NAND2_X1 port map( A1 => n16250, A2 => n16018, ZN => n849);
   U3595 : NOR2_X1 port map( A1 => n22533, A2 => n852, ZN => n22534);
   U3596 : AOI21_X1 port map( B1 => n18718, B2 => n19497, A => n19499, ZN => 
                           n18723);
   U3597 : XNOR2_X1 port map( A => n854, B => n20812, ZN => n20814);
   U3598 : XNOR2_X1 port map( A => n20811, B => n24896, ZN => n854);
   U3601 : NAND2_X1 port map( A1 => n14010, A2 => n14254, ZN => n855);
   U3602 : NAND2_X1 port map( A1 => n14255, A2 => n14252, ZN => n856);
   U3606 : NAND2_X1 port map( A1 => n10219, A2 => n857, ZN => n11616);
   U3607 : NAND2_X1 port map( A1 => n10220, A2 => n10782, ZN => n857);
   U3609 : INV_X1 port map( A => n8697, ZN => n5553);
   U3610 : XNOR2_X1 port map( A => n9106, B => n8959, ZN => n8697);
   U3611 : XNOR2_X1 port map( A => n11943, B => n11944, ZN => n3473);
   U3614 : NAND3_X1 port map( A1 => n5187, A2 => n5188, A3 => n20255, ZN => 
                           n5186);
   U3617 : NAND3_X1 port map( A1 => n5366, A2 => n281, A3 => n5367, ZN => n5599
                           );
   U3619 : NAND3_X1 port map( A1 => n22506, A2 => n23443, A3 => n321, ZN => 
                           n23444);
   U3621 : OAI211_X1 port map( C1 => n1175, C2 => n6776, A => n6290, B => n6775
                           , ZN => n6199);
   U3622 : OAI21_X1 port map( B1 => n20226, B2 => n3016, A => n862, ZN => 
                           n20271);
   U3623 : NAND2_X1 port map( A1 => n3016, A2 => n20268, ZN => n862);
   U3624 : NAND2_X1 port map( A1 => n6894, A2 => n313, ZN => n2914);
   U3625 : OAI21_X1 port map( B1 => n13013, B2 => n13245, A => n863, ZN => 
                           n12563);
   U3626 : NAND2_X1 port map( A1 => n13245, A2 => n25199, ZN => n863);
   U3627 : OR2_X1 port map( A1 => n19786, A2 => n19987, ZN => n19753);
   U3628 : NOR2_X1 port map( A1 => n21382, A2 => n22323, ZN => n22322);
   U3629 : OR2_X1 port map( A1 => n13132, A2 => n25033, ZN => n1844);
   U3630 : OAI21_X1 port map( B1 => n10570, B2 => n416, A => n864, ZN => n10576
                           );
   U3631 : NAND2_X1 port map( A1 => n10570, A2 => n10571, ZN => n864);
   U3632 : XNOR2_X2 port map( A => n1884, B => n14404, ZN => n16170);
   U3633 : INV_X1 port map( A => n21909, ZN => n22275);
   U3634 : NAND2_X1 port map( A1 => n21910, A2 => n22138, ZN => n21909);
   U3635 : INV_X1 port map( A => n1095, ZN => n15709);
   U3637 : XNOR2_X1 port map( A => n868, B => n14414, ZN => n14422);
   U3638 : XNOR2_X1 port map( A => n14960, B => n14413, ZN => n868);
   U3639 : NAND3_X1 port map( A1 => n6338, A2 => n6510, A3 => n6337, ZN => 
                           n3171);
   U3641 : NAND2_X1 port map( A1 => n4499, A2 => n13298, ZN => n1818);
   U3642 : NAND2_X1 port map( A1 => n3557, A2 => n13200, ZN => n870);
   U3643 : NAND2_X1 port map( A1 => n22952, A2 => n871, ZN => n1889);
   U3644 : NOR2_X1 port map( A1 => n24884, A2 => n22954, ZN => n871);
   U3646 : NAND2_X1 port map( A1 => n6359, A2 => n6360, ZN => n873);
   U3647 : NAND2_X1 port map( A1 => n25041, A2 => n22836, ZN => n22895);
   U3649 : NAND2_X2 port map( A1 => n874, A2 => n4796, ZN => n13868);
   U3650 : NAND2_X1 port map( A1 => n4333, A2 => n4332, ZN => n874);
   U3651 : NOR2_X1 port map( A1 => n5481, A2 => n19532, ZN => n5475);
   U3652 : AOI21_X1 port map( B1 => n17388, B2 => n17387, A => n875, ZN => 
                           n17393);
   U3654 : AOI22_X1 port map( A1 => n877, A2 => n23531, B1 => n23008, B2 => 
                           n23505, ZN => n22930);
   U3655 : NAND2_X1 port map( A1 => n23013, A2 => n24313, ZN => n877);
   U3656 : NAND2_X1 port map( A1 => n21356, A2 => n23828, ZN => n21357);
   U3657 : NAND2_X1 port map( A1 => n8528, A2 => n269, ZN => n4994);
   U3660 : NAND3_X1 port map( A1 => n24589, A2 => n13646, A3 => n13824, ZN => 
                           n13650);
   U3662 : NAND2_X1 port map( A1 => n16509, A2 => n15605, ZN => n880);
   U3664 : NAND2_X1 port map( A1 => n9601, A2 => n9602, ZN => n9607);
   U3665 : NAND2_X1 port map( A1 => n6916, A2 => n6912, ZN => n5845);
   U3666 : AND3_X1 port map( A1 => n3350, A2 => n13991, A3 => n3349, ZN => 
                           n1112);
   U3667 : INV_X1 port map( A => n17122, ZN => n2580);
   U3668 : OAI211_X1 port map( C1 => n10414, C2 => n10617, A => n10413, B => 
                           n977, ZN => n11237);
   U3669 : NAND2_X1 port map( A1 => n882, A2 => n1975, ZN => n8026);
   U3670 : NAND2_X1 port map( A1 => n1840, A2 => n8023, ZN => n882);
   U3671 : NAND2_X1 port map( A1 => n7882, A2 => n7883, ZN => n7885);
   U3672 : OR2_X2 port map( A1 => n5850, A2 => n5849, ZN => n7883);
   U3674 : NAND2_X1 port map( A1 => n19515, A2 => n19984, ZN => n883);
   U3675 : NAND2_X1 port map( A1 => n19516, A2 => n885, ZN => n884);
   U3677 : XNOR2_X1 port map( A => n1111, B => n1359, ZN => n14370);
   U3678 : NAND2_X1 port map( A1 => n7322, A2 => n7323, ZN => n2733);
   U3679 : AND2_X2 port map( A1 => n6009, A2 => n6008, ZN => n7322);
   U3680 : XNOR2_X2 port map( A => Key(74), B => Plaintext(74), ZN => n5774);
   U3681 : AND2_X1 port map( A1 => n16572, A2 => n890, ZN => n16802);
   U3682 : INV_X1 port map( A => n17122, ZN => n890);
   U3685 : NAND2_X1 port map( A1 => n2753, A2 => n22240, ZN => n22062);
   U3686 : NAND2_X1 port map( A1 => n1243, A2 => n1246, ZN => n892);
   U3687 : NAND2_X1 port map( A1 => n24480, A2 => n11143, ZN => n10304);
   U3691 : NAND2_X1 port map( A1 => n13322, A2 => n13318, ZN => n893);
   U3692 : OAI21_X1 port map( B1 => n11525, B2 => n895, A => n894, ZN => n10581
                           );
   U3693 : NAND2_X1 port map( A1 => n11525, A2 => n25060, ZN => n894);
   U3694 : AOI22_X1 port map( A1 => n17454, A2 => n17455, B1 => n17456, B2 => 
                           n17457, ZN => n17458);
   U3696 : OAI21_X1 port map( B1 => n6371, B2 => n6658, A => n6370, ZN => n897)
                           ;
   U3698 : NAND2_X1 port map( A1 => n19821, A2 => n19788, ZN => n19819);
   U3699 : NAND2_X1 port map( A1 => n1680, A2 => n2853, ZN => n23579);
   U3700 : OR2_X1 port map( A1 => n25401, A2 => n6488, ZN => n5953);
   U3701 : NOR2_X1 port map( A1 => n1127, A2 => n898, ZN => n14308);
   U3702 : NOR2_X1 port map( A1 => n900, A2 => n10788, ZN => n4051);
   U3703 : NOR2_X1 port map( A1 => n1824, A2 => n10793, ZN => n900);
   U3704 : XNOR2_X2 port map( A => n5817, B => Key(126), ZN => n6367);
   U3706 : OAI21_X1 port map( B1 => n16475, B2 => n16474, A => n901, ZN => 
                           n15460);
   U3707 : NAND2_X1 port map( A1 => n16475, A2 => n15546, ZN => n901);
   U3708 : XNOR2_X1 port map( A => n18308, B => n934, ZN => n17926);
   U3709 : NAND2_X1 port map( A1 => n11438, A2 => n25337, ZN => n902);
   U3710 : NAND2_X1 port map( A1 => n20560, A2 => n20094, ZN => n19727);
   U3711 : AOI21_X2 port map( B1 => n19726, B2 => n19719, A => n19725, ZN => 
                           n20560);
   U3712 : XNOR2_X1 port map( A => n903, B => n21696, ZN => n21698);
   U3713 : XNOR2_X1 port map( A => n21695, B => n21694, ZN => n903);
   U3714 : NAND3_X1 port map( A1 => n14416, A2 => n14278, A3 => n24958, ZN => 
                           n13444);
   U3715 : NAND3_X1 port map( A1 => n2514, A2 => n14946, A3 => n13801, ZN => 
                           n13802);
   U3716 : NAND2_X1 port map( A1 => n906, A2 => n23411, ZN => n905);
   U3717 : INV_X1 port map( A => n23410, ZN => n906);
   U3718 : NAND2_X1 port map( A1 => n23418, A2 => n24947, ZN => n907);
   U3719 : NAND3_X1 port map( A1 => n3544, A2 => n16406, A3 => n24062, ZN => 
                           n5212);
   U3720 : NAND2_X1 port map( A1 => n6488, A2 => n6781, ZN => n908);
   U3721 : NAND2_X1 port map( A1 => n6305, A2 => n6304, ZN => n909);
   U3722 : NAND2_X1 port map( A1 => n910, A2 => n24007, ZN => n3485);
   U3723 : NAND2_X1 port map( A1 => n3486, A2 => n24005, ZN => n910);
   U3724 : XNOR2_X1 port map( A => n911, B => n14903, ZN => n14906);
   U3725 : XNOR2_X1 port map( A => n14901, B => n15112, ZN => n911);
   U3728 : NAND3_X1 port map( A1 => n914, A2 => n5029, A3 => n5032, ZN => 
                           Ciphertext(14));
   U3729 : NAND2_X1 port map( A1 => n5028, A2 => n5031, ZN => n914);
   U3730 : NAND2_X1 port map( A1 => n915, A2 => n13988, ZN => n13990);
   U3731 : INV_X1 port map( A => n13987, ZN => n915);
   U3732 : NAND2_X1 port map( A1 => n5416, A2 => n13247, ZN => n13987);
   U3733 : NAND2_X1 port map( A1 => n7328, A2 => n7897, ZN => n7332);
   U3734 : NAND2_X1 port map( A1 => n24952, A2 => n23112, ZN => n5035);
   U3735 : XNOR2_X1 port map( A => n916, B => n449, ZN => Ciphertext(180));
   U3736 : NAND2_X1 port map( A1 => n23950, A2 => n23951, ZN => n916);
   U3737 : OR2_X1 port map( A1 => n6987, A2 => n6244, ZN => n6247);
   U3740 : OAI211_X2 port map( C1 => n5595, C2 => n7187, A => n918, B => n7645,
                           ZN => n8909);
   U3741 : NAND2_X1 port map( A1 => n5593, A2 => n5595, ZN => n918);
   U3742 : AOI21_X1 port map( B1 => n22468, B2 => n22675, A => n919, ZN => 
                           n22470);
   U3743 : NAND2_X1 port map( A1 => n7918, A2 => n435, ZN => n920);
   U3744 : OR3_X1 port map( A1 => n20290, A2 => n21008, A3 => n20523, ZN => 
                           n2852);
   U3746 : NAND3_X2 port map( A1 => n21933, A2 => n21932, A3 => n21931, ZN => 
                           n23201);
   U3747 : NAND2_X1 port map( A1 => n1299, A2 => n18914, ZN => n18916);
   U3748 : OR2_X1 port map( A1 => n19185, A2 => n19548, ZN => n1710);
   U3750 : OR2_X1 port map( A1 => n3822, A2 => n17613, ZN => n16562);
   U3751 : NAND2_X1 port map( A1 => n17408, A2 => n16561, ZN => n3822);
   U3752 : NAND4_X2 port map( A1 => n5984, A2 => n5985, A3 => n5983, A4 => 
                           n5982, ZN => n7604);
   U3753 : AND2_X1 port map( A1 => n17173, A2 => n927, ZN => n16435);
   U3754 : NAND2_X1 port map( A1 => n17175, A2 => n16434, ZN => n927);
   U3755 : AOI21_X1 port map( B1 => n17174, B2 => n282, A => n17175, ZN => 
                           n4413);
   U3756 : NAND2_X1 port map( A1 => n22961, A2 => n24343, ZN => n932);
   U3757 : XNOR2_X1 port map( A => n928, B => n931, ZN => Ciphertext(69));
   U3758 : NAND3_X1 port map( A1 => n929, A2 => n3014, A3 => n22995, ZN => n928
                           );
   U3759 : NAND3_X1 port map( A1 => n930, A2 => n932, A3 => n23340, ZN => n929)
                           ;
   U3760 : OR2_X1 port map( A1 => n23354, A2 => n23349, ZN => n930);
   U3761 : INV_X1 port map( A => n932, ZN => n22996);
   U3762 : AOI21_X1 port map( B1 => n933, B2 => n7868, A => n3570, ZN => n7711)
                           ;
   U3763 : XNOR2_X1 port map( A => n18310, B => n934, ZN => n16000);
   U3764 : XNOR2_X1 port map( A => n934, B => n1777, ZN => n17883);
   U3765 : XNOR2_X1 port map( A => n18285, B => n934, ZN => n18286);
   U3766 : NAND2_X1 port map( A1 => n936, A2 => n24585, ZN => n17056);
   U3767 : INV_X1 port map( A => n16932, ZN => n936);
   U3768 : NOR2_X1 port map( A1 => n24398, A2 => n16932, ZN => n16610);
   U3769 : NAND2_X1 port map( A1 => n23350, A2 => n23349, ZN => n938);
   U3770 : NAND2_X1 port map( A1 => n937, A2 => n23350, ZN => n3014);
   U3771 : OAI21_X1 port map( B1 => n24343, B2 => n24400, A => n938, ZN => 
                           n23037);
   U3772 : AOI22_X1 port map( A1 => n22979, A2 => n22996, B1 => n23363, B2 => 
                           n938, ZN => n22980);
   U3774 : NAND2_X1 port map( A1 => n24753, A2 => n939, ZN => n11096);
   U3776 : XNOR2_X1 port map( A => n13642, B => n13641, ZN => n940);
   U3777 : NAND2_X1 port map( A1 => n24960, A2 => n25500, ZN => n15811);
   U3778 : OAI21_X1 port map( B1 => n3544, B2 => n24960, A => n15646, ZN => 
                           n16199);
   U3779 : NAND2_X1 port map( A1 => n941, A2 => n7382, ZN => n7303);
   U3780 : NAND3_X1 port map( A1 => n7386, A2 => n7618, A3 => n941, ZN => n7203
                           );
   U3781 : NAND2_X1 port map( A1 => n7383, A2 => n941, ZN => n7389);
   U3782 : AOI21_X1 port map( B1 => n7616, B2 => n941, A => n7615, ZN => n7624)
                           ;
   U3783 : INV_X1 port map( A => n6156, ZN => n943);
   U3784 : NAND2_X1 port map( A1 => n8005, A2 => n7754, ZN => n8003);
   U3785 : NAND3_X1 port map( A1 => n945, A2 => n6074, A3 => n6073, ZN => n7754
                           );
   U3786 : NAND2_X1 port map( A1 => n6657, A2 => n946, ZN => n945);
   U3787 : NAND2_X1 port map( A1 => n6658, A2 => n947, ZN => n946);
   U3788 : NAND2_X1 port map( A1 => n950, A2 => n448, ZN => n949);
   U3789 : NAND2_X1 port map( A1 => n6834, A2 => n7009, ZN => n950);
   U3792 : NAND3_X1 port map( A1 => n18967, A2 => n19300, A3 => n3653, ZN => 
                           n951);
   U3793 : INV_X1 port map( A => n19297, ZN => n3653);
   U3794 : NAND3_X1 port map( A1 => n18856, A2 => n18970, A3 => n18928, ZN => 
                           n952);
   U3796 : NAND2_X1 port map( A1 => n9475, A2 => n9476, ZN => n953);
   U3797 : AOI21_X1 port map( B1 => n9473, B2 => n9864, A => n9860, ZN => n954)
                           ;
   U3798 : AND2_X1 port map( A1 => n10886, A2 => n10887, ZN => n9477);
   U3799 : NAND2_X1 port map( A1 => n9456, A2 => n956, ZN => n955);
   U3800 : NAND2_X1 port map( A1 => n961, A2 => n959, ZN => n958);
   U3801 : NAND3_X1 port map( A1 => n362, A2 => n19192, A3 => n960, ZN => n959)
                           ;
   U3802 : NAND2_X1 port map( A1 => n19571, A2 => n19570, ZN => n961);
   U3803 : AOI21_X1 port map( B1 => n19567, B2 => n19566, A => n19565, ZN => 
                           n962);
   U3804 : NAND3_X1 port map( A1 => n17230, A2 => n2285, A3 => n16951, ZN => 
                           n14589);
   U3805 : NAND3_X1 port map( A1 => n1656, A2 => n1655, A3 => n24537, ZN => 
                           n963);
   U3806 : OAI21_X1 port map( B1 => n16917, B2 => n17335, A => n16915, ZN => 
                           n16919);
   U3809 : XNOR2_X1 port map( A => n966, B => n18436, ZN => n18441);
   U3810 : INV_X1 port map( A => n966, ZN => n4808);
   U3811 : INV_X1 port map( A => n17874, ZN => n4942);
   U3812 : NAND2_X1 port map( A1 => n967, A2 => n4356, ZN => n4355);
   U3813 : NAND3_X1 port map( A1 => n967, A2 => n14159, A3 => n5080, ZN => 
                           n3085);
   U3814 : AOI22_X2 port map( A1 => n1235, A2 => n15868, B1 => n15867, B2 => 
                           n16141, ZN => n17119);
   U3815 : AND2_X2 port map( A1 => n969, A2 => n968, ZN => n17120);
   U3816 : NAND2_X1 port map( A1 => n15855, A2 => n24928, ZN => n968);
   U3818 : NAND3_X1 port map( A1 => n23828, A2 => n23827, A3 => n318, ZN => 
                           n21349);
   U3819 : AND2_X1 port map( A1 => n4219, A2 => n1099, ZN => n971);
   U3820 : NAND2_X1 port map( A1 => n303, A2 => n12795, ZN => n973);
   U3822 : OAI21_X1 port map( B1 => n12799, B2 => n12798, A => n12797, ZN => 
                           n974);
   U3823 : INV_X1 port map( A => n1646, ZN => n975);
   U3824 : AOI21_X2 port map( B1 => n976, B2 => n12802, A => n12801, ZN => 
                           n14328);
   U3826 : NAND2_X1 port map( A1 => n978, A2 => n10611, ZN => n977);
   U3827 : NAND2_X1 port map( A1 => n10614, A2 => n10486, ZN => n10611);
   U3828 : NAND2_X1 port map( A1 => n979, A2 => n980, ZN => n978);
   U3829 : NAND2_X1 port map( A1 => n10412, A2 => n10411, ZN => n979);
   U3830 : NAND2_X1 port map( A1 => n10486, A2 => n10411, ZN => n980);
   U3831 : OAI211_X1 port map( C1 => n388, C2 => n16334, A => n981, B => n15755
                           , ZN => n5317);
   U3833 : NAND2_X1 port map( A1 => n21031, A2 => n21038, ZN => n2248);
   U3835 : OR2_X1 port map( A1 => n298, A2 => n13863, ZN => n984);
   U3836 : NAND2_X1 port map( A1 => n986, A2 => n16342, ZN => n17620);
   U3837 : NAND2_X1 port map( A1 => n987, A2 => n4926, ZN => n986);
   U3839 : NOR2_X1 port map( A1 => n19575, A2 => n988, ZN => n1098);
   U3840 : MUX2_X1 port map( A => n988, B => n24982, S => n19575, Z => n1004);
   U3841 : NAND2_X1 port map( A1 => n7390, A2 => n7647, ZN => n7649);
   U3842 : INV_X1 port map( A => n7646, ZN => n7390);
   U3843 : AND2_X1 port map( A1 => n12817, A2 => n14088, ZN => n990);
   U3844 : NAND2_X1 port map( A1 => n4510, A2 => n14085, ZN => n12817);
   U3845 : NAND2_X1 port map( A1 => n13537, A2 => n13536, ZN => n14085);
   U3848 : NAND2_X1 port map( A1 => n15757, A2 => n16001, ZN => n995);
   U3849 : XNOR2_X2 port map( A => n15144, B => n15145, ZN => n16266);
   U3852 : AOI21_X1 port map( B1 => n3856, B2 => n22253, A => n332, ZN => n996)
                           ;
   U3854 : AOI21_X1 port map( B1 => n22254, B2 => n24468, A => n24362, ZN => 
                           n998);
   U3856 : NAND2_X1 port map( A1 => n20354, A2 => n20352, ZN => n999);
   U3857 : NAND2_X1 port map( A1 => n20003, A2 => n20479, ZN => n20352);
   U3858 : INV_X1 port map( A => n19057, ZN => n19060);
   U3859 : INV_X1 port map( A => n19578, ZN => n1002);
   U3861 : NAND2_X1 port map( A1 => n1005, A2 => n1004, ZN => n1003);
   U3862 : AND2_X1 port map( A1 => n23645, A2 => n23640, ZN => n23653);
   U3863 : OAI211_X1 port map( C1 => n22116, C2 => n22072, A => n22169, B => 
                           n22115, ZN => n1006);
   U3864 : OAI211_X1 port map( C1 => n20353, C2 => n20480, A => n1008, B => 
                           n20003, ZN => n1992);
   U3866 : NAND4_X2 port map( A1 => n4717, A2 => n4716, A3 => n3388, A4 => 
                           n3389, ZN => n20479);
   U3867 : INV_X1 port map( A => n20479, ZN => n2168);
   U3868 : INV_X1 port map( A => n1012, ZN => n1011);
   U3869 : INV_X1 port map( A => n19269, ZN => n1013);
   U3870 : NAND3_X1 port map( A1 => n1019, A2 => n12991, A3 => n1018, ZN => 
                           n1017);
   U3871 : NAND2_X1 port map( A1 => n2608, A2 => n1020, ZN => n1019);
   U3873 : NAND2_X1 port map( A1 => n9872, A2 => n1021, ZN => n9879);
   U3874 : NAND3_X1 port map( A1 => n4993, A2 => n2294, A3 => n1021, ZN => 
                           n9032);
   U3875 : MUX2_X1 port map( A => n9872, B => n24549, S => n9027, Z => n9549);
   U3877 : INV_X1 port map( A => n20003, ZN => n20477);
   U3878 : NOR2_X1 port map( A1 => n20003, A2 => n20479, ZN => n1024);
   U3880 : NAND2_X1 port map( A1 => n1028, A2 => n1027, ZN => n1026);
   U3882 : AND2_X1 port map( A1 => n18834, A2 => n24478, ZN => n2695);
   U3883 : NAND2_X1 port map( A1 => n19438, A2 => n24478, ZN => n18835);
   U3884 : NAND2_X1 port map( A1 => n18642, A2 => n1029, ZN => n18643);
   U3885 : AND2_X1 port map( A1 => n24478, A2 => n25422, ZN => n1029);
   U3887 : INV_X1 port map( A => n18651, ZN => n1030);
   U3888 : NAND2_X1 port map( A1 => n19081, A2 => n24478, ZN => n18651);
   U3891 : NAND2_X1 port map( A1 => n17629, A2 => n16539, ZN => n1032);
   U3892 : INV_X1 port map( A => n2566, ZN => n1033);
   U3893 : XNOR2_X1 port map( A => n18633, B => n5120, ZN => n18634);
   U3895 : NAND3_X1 port map( A1 => n17629, A2 => n2561, A3 => n17633, ZN => 
                           n1036);
   U3896 : NAND2_X1 port map( A1 => n1038, A2 => n434, ZN => n1037);
   U3897 : NAND2_X1 port map( A1 => n1039, A2 => n7078, ZN => n1038);
   U3898 : NAND2_X1 port map( A1 => n7674, A2 => n25251, ZN => n1039);
   U3899 : NAND2_X1 port map( A1 => n1041, A2 => n6869, ZN => n1040);
   U3900 : NAND2_X1 port map( A1 => n7506, A2 => n1379, ZN => n6869);
   U3901 : NAND2_X1 port map( A1 => n7510, A2 => n7509, ZN => n1041);
   U3902 : NAND2_X1 port map( A1 => n1162, A2 => n7224, ZN => n7509);
   U3903 : OR2_X2 port map( A1 => n6868, A2 => n6867, ZN => n7224);
   U3904 : NAND2_X1 port map( A1 => n7078, A2 => n7674, ZN => n7510);
   U3905 : NAND2_X1 port map( A1 => n3274, A2 => n3273, ZN => n7078);
   U3906 : NAND2_X1 port map( A1 => n1043, A2 => n1042, ZN => n1045);
   U3907 : NAND2_X1 port map( A1 => n297, A2 => n14153, ZN => n1042);
   U3908 : NAND2_X1 port map( A1 => n14154, A2 => n13805, ZN => n1043);
   U3909 : NAND3_X2 port map( A1 => n1045, A2 => n14152, A3 => n1044, ZN => 
                           n15055);
   U3910 : NAND2_X1 port map( A1 => n14151, A2 => n14150, ZN => n1044);
   U3911 : NAND2_X1 port map( A1 => n1049, A2 => n19568, ZN => n1048);
   U3912 : INV_X1 port map( A => n19191, ZN => n5634);
   U3913 : XNOR2_X2 port map( A => n18307, B => n18306, ZN => n19191);
   U3914 : NAND2_X1 port map( A1 => n19568, A2 => n1053, ZN => n1052);
   U3915 : INV_X1 port map( A => n11297, ZN => n11091);
   U3916 : NAND2_X1 port map( A1 => n9528, A2 => n2855, ZN => n11297);
   U3918 : NAND2_X1 port map( A1 => n1055, A2 => n11302, ZN => n1054);
   U3919 : INV_X1 port map( A => n11297, ZN => n1055);
   U3920 : NAND2_X1 port map( A1 => n10762, A2 => n11298, ZN => n1057);
   U3921 : AOI22_X2 port map( A1 => n10896, A2 => n1059, B1 => n10898, B2 => 
                           n10897, ZN => n11627);
   U3922 : INV_X1 port map( A => n1055, ZN => n1059);
   U3923 : NAND2_X1 port map( A1 => n391, A2 => n11454, ZN => n2301);
   U3924 : NAND2_X1 port map( A1 => n14088, A2 => n4510, ZN => n1062);
   U3925 : INV_X1 port map( A => n25372, ZN => n21648);
   U3926 : XNOR2_X1 port map( A => n21650, B => n1063, ZN => n21651);
   U3927 : XNOR2_X1 port map( A => n25372, B => n24319, ZN => n1063);
   U3929 : OAI22_X1 port map( A1 => n22941, A2 => n337, B1 => n22832, B2 => 
                           n22940, ZN => n1066);
   U3931 : NAND2_X1 port map( A1 => n25063, A2 => n1066, ZN => n1065);
   U3932 : NAND2_X1 port map( A1 => n22830, A2 => n22832, ZN => n1068);
   U3933 : NOR2_X1 port map( A1 => n23398, A2 => n23420, ZN => n22868);
   U3934 : NAND2_X1 port map( A1 => n13097, A2 => n1069, ZN => n1080);
   U3936 : NAND2_X1 port map( A1 => n13094, A2 => n3492, ZN => n1069);
   U3937 : NAND3_X1 port map( A1 => n16612, A2 => n16730, A3 => n283, ZN => 
                           n1070);
   U3938 : NAND2_X1 port map( A1 => n5761, A2 => n1071, ZN => n16613);
   U3939 : NAND2_X1 port map( A1 => n1073, A2 => n1072, ZN => n20053);
   U3940 : NAND2_X1 port map( A1 => n20480, A2 => n20476, ZN => n20051);
   U3941 : NAND2_X1 port map( A1 => n20048, A2 => n2168, ZN => n1073);
   U3942 : NAND2_X1 port map( A1 => n1075, A2 => n23311, ZN => n5660);
   U3943 : NAND2_X1 port map( A1 => n5662, A2 => n5664, ZN => n1074);
   U3946 : OAI22_X1 port map( A1 => n21891, A2 => n24881, B1 => n4109, B2 => 
                           n22974, ZN => n1076);
   U3947 : NOR2_X1 port map( A1 => n7590, A2 => n7591, ZN => n1194);
   U3948 : OAI21_X2 port map( B1 => n5452, B2 => n1079, A => n1077, ZN => n7591
                           );
   U3949 : NAND2_X1 port map( A1 => n1078, A2 => n1698, ZN => n1077);
   U3950 : NAND2_X1 port map( A1 => n6315, A2 => n6467, ZN => n6328);
   U3951 : NAND3_X1 port map( A1 => n13119, A2 => n13113, A3 => n12503, ZN => 
                           n1082);
   U3952 : NAND2_X1 port map( A1 => n7508, A2 => n1083, ZN => n2263);
   U3953 : NAND2_X1 port map( A1 => n1084, A2 => n7506, ZN => n1083);
   U3954 : INV_X1 port map( A => n13900, ZN => n13958);
   U3955 : NAND2_X1 port map( A1 => n12659, A2 => n12503, ZN => n1087);
   U3956 : NAND2_X1 port map( A1 => n12291, A2 => n3328, ZN => n1086);
   U3957 : NAND2_X1 port map( A1 => n13958, A2 => n13903, ZN => n13459);
   U3958 : AOI21_X1 port map( B1 => n7262, B2 => n1088, A => n7261, ZN => n7265
                           );
   U3959 : XNOR2_X1 port map( A => n1089, B => n8263, ZN => n8267);
   U3960 : INV_X1 port map( A => n8851, ZN => n1089);
   U3961 : XNOR2_X1 port map( A => n1090, B => n8851, ZN => n8838);
   U3962 : INV_X1 port map( A => n8835, ZN => n1090);
   U3963 : XNOR2_X1 port map( A => n1091, B => n15338, ZN => n14652);
   U3964 : XNOR2_X1 port map( A => n1091, B => n15485, ZN => n15492);
   U3965 : XNOR2_X1 port map( A => n1091, B => n15239, ZN => n15243);
   U3968 : OAI21_X1 port map( B1 => n9953, B2 => n9955, A => n9949, ZN => n1093
                           );
   U3970 : NAND2_X1 port map( A1 => n16439, A2 => n1095, ZN => n16446);
   U3971 : OAI22_X1 port map( A1 => n1097, A2 => n16492, B1 => n16490, B2 => 
                           n387, ZN => n1096);
   U3973 : NAND3_X1 port map( A1 => n21839, A2 => n22361, A3 => n245, ZN => 
                           n1099);
   U3974 : NAND2_X1 port map( A1 => n24608, A2 => n22356, ZN => n1100);
   U3977 : NAND2_X1 port map( A1 => n6189, A2 => n1106, ZN => n4881);
   U3978 : NAND2_X1 port map( A1 => n6195, A2 => n6445, ZN => n6453);
   U3979 : NAND2_X1 port map( A1 => n19315, A2 => n19312, ZN => n1107);
   U3980 : NAND2_X1 port map( A1 => n17563, A2 => n1107, ZN => n17565);
   U3981 : NOR2_X1 port map( A1 => n1109, A2 => n19984, ZN => n1108);
   U3982 : NOR2_X2 port map( A1 => n1159, A2 => n18926, ZN => n19984);
   U3983 : INV_X1 port map( A => n24464, ZN => n1109);
   U3984 : XNOR2_X1 port map( A => n1110, B => n8615, ZN => n8071);
   U3985 : XNOR2_X1 port map( A => n9034, B => n1110, ZN => n9037);
   U3986 : XNOR2_X1 port map( A => n8491, B => n1110, ZN => n7980);
   U3987 : XNOR2_X1 port map( A => n8537, B => n1110, ZN => n7594);
   U3988 : NAND2_X1 port map( A1 => n16474, A2 => n16473, ZN => n15688);
   U3989 : NAND3_X1 port map( A1 => n16469, A2 => n15546, A3 => n16471, ZN => 
                           n1113);
   U3990 : NAND3_X1 port map( A1 => n16472, A2 => n16473, A3 => n16474, ZN => 
                           n1114);
   U3991 : MUX2_X1 port map( A => n16578, B => n17086, S => n16649, Z => n15875
                           );
   U3992 : NAND2_X1 port map( A1 => n15795, A2 => n16069, ZN => n1115);
   U3994 : NAND2_X1 port map( A1 => n1119, A2 => n6255, ZN => n1116);
   U3995 : NAND2_X1 port map( A1 => n5905, A2 => n25437, ZN => n1118);
   U3996 : AOI21_X1 port map( B1 => n6254, B2 => n1119, A => n6528, ZN => n6258
                           );
   U3997 : NAND2_X1 port map( A1 => n6948, A2 => n6529, ZN => n1119);
   U3998 : OAI22_X1 port map( A1 => n19565, A2 => n19273, B1 => n19192, B2 => 
                           n19570, ZN => n19274);
   U3999 : XNOR2_X2 port map( A => n18330, B => n18329, ZN => n19570);
   U4000 : NAND2_X1 port map( A1 => n19274, A2 => n18907, ZN => n1120);
   U4001 : NAND2_X1 port map( A1 => n363, A2 => n19570, ZN => n18907);
   U4002 : NAND2_X1 port map( A1 => n18794, A2 => n18793, ZN => n1121);
   U4004 : INV_X1 port map( A => n15667, ZN => n1123);
   U4005 : NOR2_X1 port map( A1 => n3947, A2 => n25092, ZN => n16335);
   U4006 : AND2_X1 port map( A1 => n267, A2 => n16332, ZN => n16339);
   U4008 : OAI21_X2 port map( B1 => n12426, B2 => n13150, A => n1125, ZN => 
                           n14307);
   U4009 : NAND2_X1 port map( A1 => n1126, A2 => n13129, ZN => n1125);
   U4010 : OAI21_X1 port map( B1 => n13148, B2 => n13130, A => n13131, ZN => 
                           n1126);
   U4011 : NAND3_X1 port map( A1 => n1128, A2 => n7139, A3 => n7896, ZN => 
                           n7143);
   U4012 : NAND2_X1 port map( A1 => n1130, A2 => n3469, ZN => n1128);
   U4013 : INV_X1 port map( A => n3469, ZN => n7902);
   U4014 : NAND2_X2 port map( A1 => n1129, A2 => n1398, ZN => n3469);
   U4015 : NAND2_X1 port map( A1 => n5876, A2 => n5875, ZN => n1129);
   U4016 : INV_X1 port map( A => n7327, ZN => n1130);
   U4018 : NAND3_X1 port map( A1 => n1138, A2 => n17067, A3 => n17066, ZN => 
                           n1133);
   U4019 : NAND2_X1 port map( A1 => n17069, A2 => n1139, ZN => n16734);
   U4020 : NAND3_X1 port map( A1 => n15609, A2 => n1136, A3 => n1134, ZN => 
                           n18262);
   U4021 : NAND2_X1 port map( A1 => n1135, A2 => n283, ZN => n1134);
   U4022 : NAND2_X1 port map( A1 => n16730, A2 => n1137, ZN => n1136);
   U4023 : AND2_X1 port map( A1 => n1139, A2 => n16546, ZN => n1137);
   U4024 : XNOR2_X1 port map( A => n1140, B => n23693, ZN => Ciphertext(129));
   U4025 : NAND3_X1 port map( A1 => n1143, A2 => n1142, A3 => n1141, ZN => 
                           n1140);
   U4026 : NAND2_X1 port map( A1 => n23691, A2 => n25026, ZN => n1141);
   U4027 : NAND2_X1 port map( A1 => n25405, A2 => n23686, ZN => n1142);
   U4028 : NOR2_X1 port map( A1 => n23670, A2 => n25026, ZN => n23686);
   U4029 : NAND2_X1 port map( A1 => n1144, A2 => n23670, ZN => n1143);
   U4030 : NAND3_X1 port map( A1 => n4702, A2 => n4703, A3 => n4700, ZN => 
                           Ciphertext(130));
   U4031 : NAND2_X1 port map( A1 => n22200, A2 => n1146, ZN => n22179);
   U4032 : NAND2_X1 port map( A1 => n325, A2 => n1146, ZN => n4362);
   U4033 : OAI21_X1 port map( B1 => n325, B2 => n1146, A => n22200, ZN => 
                           n21804);
   U4035 : NAND2_X1 port map( A1 => n6976, A2 => n1147, ZN => n6692);
   U4037 : NAND2_X1 port map( A1 => n6686, A2 => n1147, ZN => n6390);
   U4039 : INV_X1 port map( A => n6690, ZN => n1149);
   U4040 : NAND2_X1 port map( A1 => n1150, A2 => n4110, ZN => n1613);
   U4042 : NAND2_X1 port map( A1 => n4175, A2 => n20384, ZN => n1152);
   U4043 : NAND2_X1 port map( A1 => n1613, A2 => n4176, ZN => n21743);
   U4044 : OAI21_X2 port map( B1 => n19882, B2 => n20554, A => n19881, ZN => 
                           n1153);
   U4045 : XNOR2_X1 port map( A => n1153, B => n21985, ZN => n20818);
   U4046 : XNOR2_X1 port map( A => n1153, B => n452, ZN => n20991);
   U4047 : XNOR2_X1 port map( A => n1153, B => n1758, ZN => n21462);
   U4049 : NOR2_X1 port map( A1 => n23652, A2 => n23649, ZN => n22151);
   U4050 : NAND2_X1 port map( A1 => n20856, A2 => n2601, ZN => n1156);
   U4051 : NAND2_X1 port map( A1 => n21802, A2 => n22200, ZN => n1158);
   U4052 : NAND2_X1 port map( A1 => n18922, A2 => n264, ZN => n1161);
   U4053 : NAND2_X1 port map( A1 => n14044, A2 => n5246, ZN => n1930);
   U4054 : NAND2_X1 port map( A1 => n20111, A2 => n19916, ZN => n5123);
   U4055 : NOR2_X2 port map( A1 => n17714, A2 => n17713, ZN => n19883);
   U4056 : NAND3_X1 port map( A1 => n1162, A2 => n7078, A3 => n25251, ZN => 
                           n7075);
   U4057 : MUX2_X2 port map( A => n7226, B => n7227, S => n7676, Z => n8491);
   U4059 : NAND2_X1 port map( A1 => n24083, A2 => n9944, ZN => n1165);
   U4061 : MUX2_X1 port map( A => n10848, B => n10850, S => n11122, Z => n1166)
                           ;
   U4063 : NAND2_X1 port map( A1 => n3546, A2 => n1479, ZN => n10848);
   U4064 : INV_X1 port map( A => n11124, ZN => n1167);
   U4066 : NAND2_X1 port map( A1 => n10721, A2 => n11124, ZN => n1170);
   U4067 : OAI211_X1 port map( C1 => n7008, C2 => n7009, A => n1173, B => n7006
                           , ZN => n1174);
   U4068 : NAND2_X1 port map( A1 => n7009, A2 => n7004, ZN => n1173);
   U4069 : NAND2_X1 port map( A1 => n283, A2 => n17068, ZN => n16611);
   U4070 : NAND3_X1 port map( A1 => n283, A2 => n17068, A3 => n16612, ZN => 
                           n5307);
   U4071 : INV_X1 port map( A => n6198, ZN => n1175);
   U4073 : NOR2_X1 port map( A1 => n25480, A2 => n1176, ZN => n5964);
   U4074 : AOI21_X1 port map( B1 => n6923, B2 => n6922, A => n1176, ZN => n6928
                           );
   U4075 : INV_X1 port map( A => n6776, ZN => n1176);
   U4076 : XNOR2_X1 port map( A => n1177, B => n21662, ZN => n10431);
   U4077 : XNOR2_X1 port map( A => n1177, B => n21553, ZN => n9406);
   U4078 : XNOR2_X1 port map( A => n11735, B => n1177, ZN => n10638);
   U4079 : XNOR2_X1 port map( A => n11564, B => n1177, ZN => n11537);
   U4080 : NAND3_X2 port map( A1 => n9404, A2 => n9405, A3 => n1178, ZN => 
                           n1177);
   U4081 : NOR2_X2 port map( A1 => n19840, A2 => n1179, ZN => n3198);
   U4082 : OAI22_X1 port map( A1 => n3203, A2 => n19390, B1 => n24909, B2 => 
                           n3202, ZN => n1179);
   U4083 : AND2_X1 port map( A1 => n3198, A2 => n19839, ZN => n19842);
   U4085 : NAND2_X1 port map( A1 => n411, A2 => n10798, ZN => n1180);
   U4086 : NAND2_X1 port map( A1 => n10651, A2 => n10245, ZN => n10243);
   U4087 : NAND2_X1 port map( A1 => n9932, A2 => n25217, ZN => n1182);
   U4088 : AOI22_X1 port map( A1 => n9345, A2 => n9928, B1 => n9926, B2 => 
                           n9925, ZN => n1183);
   U4089 : AOI21_X2 port map( B1 => n1186, B2 => n1185, A => n1184, ZN => 
                           n10651);
   U4090 : NAND2_X1 port map( A1 => n1602, A2 => n4166, ZN => n1184);
   U4091 : OAI21_X2 port map( B1 => n17730, B2 => n1189, A => n1187, ZN => 
                           n18370);
   U4092 : MUX2_X1 port map( A => n17731, B => n1188, S => n25472, Z => n1187);
   U4093 : NAND2_X1 port map( A1 => n17733, A2 => n17486, ZN => n1188);
   U4094 : MUX2_X1 port map( A => n17728, B => n17729, S => n17486, Z => n1189)
                           ;
   U4095 : NOR2_X2 port map( A1 => n15841, A2 => n15840, ZN => n17486);
   U4096 : NAND2_X1 port map( A1 => n1194, A2 => n7588, ZN => n1191);
   U4097 : NAND3_X1 port map( A1 => n1839, A2 => n7590, A3 => n7462, ZN => 
                           n1193);
   U4098 : NAND2_X1 port map( A1 => n7588, A2 => n7590, ZN => n7593);
   U4099 : NAND3_X1 port map( A1 => n2035, A2 => n7591, A3 => n7464, ZN => 
                           n1195);
   U4100 : NAND2_X1 port map( A1 => n7236, A2 => n7962, ZN => n1196);
   U4101 : NAND2_X1 port map( A1 => n25024, A2 => n23064, ZN => n1198);
   U4102 : NAND2_X1 port map( A1 => n1199, A2 => n10951, ZN => n10957);
   U4103 : NAND2_X1 port map( A1 => n2754, A2 => n10950, ZN => n1199);
   U4104 : NAND2_X1 port map( A1 => n10698, A2 => n25074, ZN => n10950);
   U4105 : NAND2_X1 port map( A1 => n13275, A2 => n1201, ZN => n13276);
   U4107 : NOR2_X1 port map( A1 => n367, A2 => n4004, ZN => n3655);
   U4109 : OR2_X1 port map( A1 => n16272, A2 => n4516, ZN => n1202);
   U4110 : NAND2_X1 port map( A1 => n296, A2 => n1028, ZN => n1204);
   U4111 : NAND3_X1 port map( A1 => n296, A2 => n1028, A3 => n14153, ZN => 
                           n14152);
   U4113 : NOR2_X1 port map( A1 => n13512, A2 => n14031, ZN => n1203);
   U4114 : AND2_X1 port map( A1 => n20193, A2 => n20576, ZN => n1206);
   U4116 : NAND2_X1 port map( A1 => n3198, A2 => n20576, ZN => n20438);
   U4118 : NAND2_X1 port map( A1 => n1208, A2 => n15811, ZN => n15812);
   U4119 : NAND2_X1 port map( A1 => n16404, A2 => n16401, ZN => n1208);
   U4121 : OR2_X1 port map( A1 => n9523, A2 => n1210, ZN => n3028);
   U4122 : INV_X1 port map( A => n9843, ZN => n1210);
   U4123 : OR2_X1 port map( A1 => n1211, A2 => n19103, ZN => n18021);
   U4124 : NOR2_X1 port map( A1 => n19360, A2 => n24312, ZN => n1211);
   U4126 : INV_X1 port map( A => n18817, ZN => n1212);
   U4127 : NAND2_X1 port map( A1 => n16404, A2 => n15646, ZN => n1214);
   U4129 : NAND2_X1 port map( A1 => n9803, A2 => n11053, ZN => n1216);
   U4130 : NAND2_X1 port map( A1 => n1218, A2 => n11058, ZN => n1217);
   U4131 : NAND2_X1 port map( A1 => n1523, A2 => n11499, ZN => n1219);
   U4132 : NAND2_X1 port map( A1 => n9802, A2 => n11499, ZN => n1220);
   U4133 : NAND2_X1 port map( A1 => n24499, A2 => n12459, ZN => n12653);
   U4135 : OAI21_X1 port map( B1 => n13177, B2 => n13176, A => n12506, ZN => 
                           n10362);
   U4137 : INV_X1 port map( A => n11205, ZN => n1224);
   U4138 : NAND2_X1 port map( A1 => n4152, A2 => n10819, ZN => n1226);
   U4140 : NAND3_X1 port map( A1 => n25025, A2 => n11342, A3 => n1224, ZN => 
                           n1223);
   U4141 : NAND2_X1 port map( A1 => n10232, A2 => n414, ZN => n1227);
   U4143 : NAND2_X1 port map( A1 => n1233, A2 => n1228, ZN => n18146);
   U4144 : NAND2_X1 port map( A1 => n14353, A2 => n25246, ZN => n1233);
   U4145 : NAND2_X1 port map( A1 => n15865, A2 => n15866, ZN => n1235);
   U4147 : XNOR2_X2 port map( A => n21315, B => n21314, ZN => n22222);
   U4148 : INV_X1 port map( A => n22221, ZN => n1238);
   U4149 : XNOR2_X2 port map( A => n21330, B => n21329, ZN => n22221);
   U4150 : NAND2_X1 port map( A1 => n1239, A2 => n10558, ZN => n10337);
   U4151 : INV_X1 port map( A => n25250, ZN => n1239);
   U4152 : NAND3_X1 port map( A1 => n1239, A2 => n10559, A3 => n10655, ZN => 
                           n4540);
   U4153 : NAND2_X1 port map( A1 => n1240, A2 => n10314, ZN => n10316);
   U4154 : NAND2_X1 port map( A1 => n10558, A2 => n25250, ZN => n1240);
   U4155 : NOR2_X1 port map( A1 => n19862, A2 => n1242, ZN => n19865);
   U4156 : OAI21_X1 port map( B1 => n20038, B2 => n20191, A => n1241, ZN => 
                           n20040);
   U4157 : NAND2_X1 port map( A1 => n20038, A2 => n20039, ZN => n1241);
   U4158 : NOR2_X1 port map( A1 => n20185, A2 => n1242, ZN => n20187);
   U4159 : NAND2_X1 port map( A1 => n1244, A2 => n17598, ZN => n1243);
   U4160 : NAND3_X1 port map( A1 => n3316, A2 => n4574, A3 => n1483, ZN => 
                           n1245);
   U4161 : NAND2_X1 port map( A1 => n17596, A2 => n24543, ZN => n1246);
   U4162 : NOR2_X1 port map( A1 => n14180, A2 => n1247, ZN => n14183);
   U4163 : INV_X1 port map( A => n14181, ZN => n1247);
   U4164 : INV_X1 port map( A => n21839, ZN => n22358);
   U4165 : NOR2_X1 port map( A1 => n22361, A2 => n22358, ZN => n1248);
   U4166 : AND2_X1 port map( A1 => n21782, A2 => n22361, ZN => n22359);
   U4167 : INV_X1 port map( A => n21838, ZN => n21782);
   U4170 : NAND2_X1 port map( A1 => n24172, A2 => n19459, ZN => n1251);
   U4171 : NAND2_X1 port map( A1 => n15938, A2 => n16247, ZN => n2359);
   U4172 : NAND2_X1 port map( A1 => n16018, A2 => n15938, ZN => n15568);
   U4173 : NAND2_X1 port map( A1 => n17058, A2 => n17057, ZN => n1252);
   U4174 : NAND2_X1 port map( A1 => n1254, A2 => n7893, ZN => n7455);
   U4175 : NAND2_X1 port map( A1 => n1254, A2 => n7889, ZN => n7325);
   U4176 : OAI21_X1 port map( B1 => n20410, B2 => n20411, A => n345, ZN => 
                           n1255);
   U4177 : NAND2_X1 port map( A1 => n20872, A2 => n20412, ZN => n20873);
   U4178 : MUX2_X1 port map( A => n25421, B => n20411, S => n20262, Z => n20872
                           );
   U4179 : MUX2_X1 port map( A => n22952, B => n22033, S => n22954, Z => n1259)
                           ;
   U4180 : XNOR2_X2 port map( A => n21605, B => n21604, ZN => n22954);
   U4182 : AND2_X1 port map( A1 => n15804, A2 => n1261, ZN => n4337);
   U4183 : NOR2_X1 port map( A1 => n15856, A2 => n1261, ZN => n15858);
   U4185 : MUX2_X1 port map( A => n15856, B => n16117, S => n1261, Z => n4338);
   U4186 : MUX2_X1 port map( A => n15614, B => n15613, S => n1261, Z => n15617)
                           ;
   U4188 : XNOR2_X2 port map( A => n14481, B => n14480, ZN => n1261);
   U4190 : INV_X1 port map( A => n1263, ZN => n1262);
   U4193 : NAND2_X1 port map( A1 => n3119, A2 => n10767, ZN => n11082);
   U4194 : NAND2_X1 port map( A1 => n1503, A2 => n1504, ZN => n20383);
   U4195 : NAND2_X1 port map( A1 => n3943, A2 => n1506, ZN => n1503);
   U4196 : NAND2_X1 port map( A1 => n1266, A2 => n1265, ZN => n3943);
   U4197 : NAND2_X1 port map( A1 => n1268, A2 => n12503, ZN => n5402);
   U4200 : XNOR2_X1 port map( A => n18258, B => n25000, ZN => n18619);
   U4202 : NAND2_X1 port map( A1 => n9524, A2 => n9774, ZN => n1272);
   U4203 : NAND2_X1 port map( A1 => n25393, A2 => n9772, ZN => n1273);
   U4206 : INV_X1 port map( A => n22268, ZN => n1276);
   U4209 : NAND2_X1 port map( A1 => n7914, A2 => n7917, ZN => n1281);
   U4210 : NAND2_X1 port map( A1 => n7634, A2 => n7449, ZN => n7920);
   U4211 : INV_X1 port map( A => n17237, ZN => n1285);
   U4212 : OAI211_X1 port map( C1 => n16859, C2 => n17236, A => n1284, B => 
                           n1283, ZN => n16860);
   U4213 : NAND2_X1 port map( A1 => n17341, A2 => n3872, ZN => n1286);
   U4214 : INV_X1 port map( A => n17346, ZN => n17236);
   U4215 : NAND2_X2 port map( A1 => n1763, A2 => n15365, ZN => n17346);
   U4216 : AND3_X2 port map( A1 => n15309, A2 => n1812, A3 => n15310, ZN => 
                           n17241);
   U4217 : INV_X1 port map( A => n1289, ZN => n1288);
   U4218 : AOI21_X1 port map( B1 => n18835, B2 => n19437, A => n25422, ZN => 
                           n1289);
   U4219 : NAND2_X1 port map( A1 => n361, A2 => n18834, ZN => n19437);
   U4220 : AND2_X1 port map( A1 => n19441, A2 => n25422, ZN => n1291);
   U4221 : INV_X1 port map( A => n19441, ZN => n19245);
   U4222 : AND2_X1 port map( A1 => n24922, A2 => n24885, ZN => n22956);
   U4223 : NOR2_X1 port map( A1 => n22958, A2 => n1292, ZN => n21879);
   U4224 : NAND2_X1 port map( A1 => n24884, A2 => n1293, ZN => n1292);
   U4225 : NOR2_X1 port map( A1 => n6481, A2 => n6198, ZN => n1294);
   U4227 : INV_X1 port map( A => n9418, ZN => n9973);
   U4228 : NAND2_X1 port map( A1 => n25005, A2 => n9418, ZN => n9417);
   U4229 : NAND2_X1 port map( A1 => n1296, A2 => n1712, ZN => n19726);
   U4230 : NAND2_X1 port map( A1 => n1714, A2 => n19404, ZN => n1296);
   U4232 : OR2_X1 port map( A1 => n6244, A2 => n1297, ZN => n6641);
   U4233 : NAND2_X1 port map( A1 => n6987, A2 => n6640, ZN => n1297);
   U4235 : INV_X1 port map( A => n19261, ZN => n1299);
   U4236 : NOR2_X1 port map( A1 => n19264, A2 => n1300, ZN => n17558);
   U4237 : AOI21_X1 port map( B1 => n1299, B2 => n19264, A => n1300, ZN => 
                           n18918);
   U4238 : INV_X1 port map( A => n18914, ZN => n1300);
   U4239 : NAND2_X1 port map( A1 => n1304, A2 => n1301, ZN => n21282);
   U4240 : NAND2_X1 port map( A1 => n22578, A2 => n1302, ZN => n1301);
   U4241 : NAND2_X1 port map( A1 => n23064, A2 => n23077, ZN => n1302);
   U4244 : NAND2_X1 port map( A1 => n1309, A2 => n18586, ZN => n1308);
   U4245 : AOI21_X1 port map( B1 => n1311, B2 => n1310, A => n328, ZN => n1312)
                           ;
   U4246 : INV_X1 port map( A => n21794, ZN => n1311);
   U4247 : NAND3_X2 port map( A1 => n2811, A2 => n16501, A3 => n1313, ZN => 
                           n18331);
   U4250 : NAND2_X1 port map( A1 => n12979, A2 => n25053, ZN => n1315);
   U4252 : INV_X1 port map( A => n9808, ZN => n9339);
   U4253 : AND2_X1 port map( A1 => n10284, A2 => n11113, ZN => n10285);
   U4254 : NAND2_X1 port map( A1 => n10870, A2 => n10873, ZN => n10284);
   U4255 : NAND2_X1 port map( A1 => n9337, A2 => n9529, ZN => n1317);
   U4256 : NAND3_X1 port map( A1 => n6274, A2 => n6324, A3 => n315, ZN => n1320
                           );
   U4258 : NAND2_X1 port map( A1 => n6518, A2 => n6517, ZN => n1321);
   U4259 : NAND3_X1 port map( A1 => n1322, A2 => n23053, A3 => n23052, ZN => 
                           n23054);
   U4260 : INV_X1 port map( A => n23571, ZN => n1323);
   U4261 : INV_X2 port map( A => n18596, ZN => n19760);
   U4262 : XNOR2_X1 port map( A => n11237, B => n11568, ZN => n11880);
   U4263 : AND2_X1 port map( A1 => n5440, A2 => n13868, ZN => n13600);
   U4264 : XNOR2_X1 port map( A => n10320, B => n1325, ZN => n1324);
   U4265 : XOR2_X1 port map( A => n11536, B => n10310, Z => n1325);
   U4266 : OR2_X1 port map( A1 => n10772, A2 => n415, ZN => n11033);
   U4269 : INV_X1 port map( A => n24397, ZN => n1328);
   U4270 : OAI211_X1 port map( C1 => n12931, C2 => n12930, A => n4457, B => 
                           n12929, ZN => n1331);
   U4271 : OR2_X1 port map( A1 => n8752, A2 => n2159, ZN => n1332);
   U4272 : XNOR2_X1 port map( A => n14426, B => n14425, ZN => n16423);
   U4273 : XNOR2_X1 port map( A => n8717, B => n8718, ZN => n10071);
   U4274 : OAI211_X1 port map( C1 => n12931, C2 => n12930, A => n4457, B => 
                           n12929, ZN => n14129);
   U4276 : XOR2_X1 port map( A => n18266, B => n18265, Z => n1334);
   U4277 : XOR2_X1 port map( A => n11364, B => n11365, Z => n1335);
   U4278 : XNOR2_X1 port map( A => n3141, B => n21748, ZN => n1336);
   U4279 : XOR2_X1 port map( A => n8088, B => n9169, Z => n1337);
   U4280 : OR2_X1 port map( A1 => n17293, A2 => n17233, ZN => n1339);
   U4282 : XNOR2_X1 port map( A => n3141, B => n21748, ZN => n22245);
   U4287 : NAND2_X1 port map( A1 => n14236, A2 => n14235, ZN => n1342);
   U4288 : NAND2_X1 port map( A1 => n14234, A2 => n14233, ZN => n1343);
   U4292 : XOR2_X1 port map( A => n11243, B => n11741, Z => n12322);
   U4293 : INV_X1 port map( A => n15715, ZN => n16474);
   U4294 : OAI21_X1 port map( B1 => n15820, B2 => n15819, A => n16426, ZN => 
                           n15835);
   U4295 : OAI211_X2 port map( C1 => n11008, C2 => n4088, A => n4495, B => 
                           n1921, ZN => n12295);
   U4296 : AND2_X1 port map( A1 => n19320, A2 => n19319, ZN => n1344);
   U4297 : NAND2_X1 port map( A1 => n10093, A2 => n9676, ZN => n1347);
   U4298 : XNOR2_X1 port map( A => n2276, B => n1903, ZN => n1348);
   U4299 : XNOR2_X1 port map( A => n1903, B => n2276, ZN => n9779);
   U4300 : NAND3_X1 port map( A1 => n1727, A2 => n2926, A3 => n5231, ZN => 
                           n1349);
   U4302 : NOR2_X1 port map( A1 => n13523, A2 => n13522, ZN => n1351);
   U4303 : XNOR2_X1 port map( A => n20750, B => n20749, ZN => n1352);
   U4304 : XNOR2_X1 port map( A => n11650, B => n11649, ZN => n1353);
   U4306 : NAND3_X1 port map( A1 => n1727, A2 => n2926, A3 => n5231, ZN => 
                           n23157);
   U4307 : NOR2_X1 port map( A1 => n13523, A2 => n13522, ZN => n15005);
   U4308 : XNOR2_X1 port map( A => n18527, B => n18526, ZN => n19238);
   U4309 : XNOR2_X1 port map( A => n20750, B => n20749, ZN => n22270);
   U4310 : XNOR2_X1 port map( A => n11650, B => n11649, ZN => n13159);
   U4311 : XOR2_X1 port map( A => n14763, B => n15106, Z => n14767);
   U4312 : XOR2_X1 port map( A => n14858, B => n14857, Z => n15160);
   U4314 : AOI21_X2 port map( B1 => n15759, B2 => n5666, A => n5668, ZN => 
                           n16539);
   U4315 : OAI21_X1 port map( B1 => n1871, B2 => n9691, A => n9690, ZN => 
                           n10961);
   U4316 : INV_X1 port map( A => n11158, ZN => n1358);
   U4320 : NOR2_X1 port map( A1 => n13799, A2 => n13798, ZN => n1359);
   U4322 : XOR2_X1 port map( A => n18379, B => n18378, Z => n1361);
   U4323 : NOR2_X1 port map( A1 => n13799, A2 => n13798, ZN => n14982);
   U4324 : XNOR2_X1 port map( A => n8939, B => n2276, ZN => n9255);
   U4325 : MUX2_X1 port map( A => n22706, B => n23278, S => n23265, Z => n22707
                           );
   U4326 : INV_X1 port map( A => n23265, ZN => n23274);
   U4327 : AND2_X1 port map( A1 => n13035, A2 => n13036, ZN => n1362);
   U4329 : OAI21_X2 port map( B1 => n12923, B2 => n12924, A => n12922, ZN => 
                           n14127);
   U4330 : XOR2_X1 port map( A => n8427, B => n8846, Z => n8628);
   U4332 : XNOR2_X2 port map( A => n5894, B => Key(50), ZN => n6699);
   U4333 : AOI22_X1 port map( A1 => n16015, A2 => n16345, B1 => n16014, B2 => 
                           n24539, ZN => n17463);
   U4335 : INV_X1 port map( A => n16106, ZN => n4689);
   U4336 : AOI21_X1 port map( B1 => n15592, B2 => n15591, A => n15590, ZN => 
                           n17065);
   U4337 : OAI21_X2 port map( B1 => n6711, B2 => n7998, A => n6710, ZN => n8846
                           );
   U4342 : INV_X1 port map( A => n7628, ZN => n7913);
   U4343 : OR2_X1 port map( A1 => n9433, A2 => n10037, ZN => n9714);
   U4344 : XNOR2_X1 port map( A => n310, B => n8506, ZN => n8084);
   U4345 : INV_X1 port map( A => n10169, ZN => n2207);
   U4347 : INV_X1 port map( A => n12040, ZN => n12213);
   U4348 : INV_X1 port map( A => n10934, ZN => n2311);
   U4349 : XNOR2_X1 port map( A => n3899, B => n12355, ZN => n11194);
   U4350 : INV_X1 port map( A => n11268, ZN => n3899);
   U4351 : OR2_X1 port map( A1 => n10811, A2 => n10812, ZN => n5629);
   U4352 : OR2_X1 port map( A1 => n11298, A2 => n10762, ZN => n10763);
   U4353 : INV_X1 port map( A => n25027, ZN => n3512);
   U4354 : OR2_X1 port map( A1 => n12773, A2 => n12774, ZN => n13069);
   U4355 : NOR2_X1 port map( A1 => n13071, A2 => n12470, ZN => n1544);
   U4356 : INV_X1 port map( A => n12856, ZN => n4196);
   U4357 : INV_X1 port map( A => n13347, ZN => n3766);
   U4358 : XNOR2_X1 port map( A => n11076, B => n11582, ZN => n12046);
   U4360 : XNOR2_X1 port map( A => n12131, B => n3206, ZN => n3204);
   U4361 : XNOR2_X1 port map( A => n12127, B => n2834, ZN => n3206);
   U4362 : XNOR2_X1 port map( A => n4996, B => n4995, ZN => n11328);
   U4363 : XNOR2_X1 port map( A => n11321, B => n11320, ZN => n4995);
   U4364 : NOR2_X1 port map( A1 => n12951, A2 => n2295, ZN => n12604);
   U4365 : AND2_X1 port map( A1 => n24346, A2 => n404, ZN => n3813);
   U4367 : XNOR2_X1 port map( A => n3862, B => n3861, ZN => n11722);
   U4368 : XNOR2_X1 port map( A => n11880, B => n11700, ZN => n3861);
   U4369 : XNOR2_X1 port map( A => n11699, B => n11702, ZN => n3862);
   U4371 : INV_X1 port map( A => n3341, ZN => n14206);
   U4372 : INV_X1 port map( A => n13386, ZN => n13646);
   U4373 : OR2_X1 port map( A1 => n13277, A2 => n24346, ZN => n4387);
   U4374 : INV_X1 port map( A => n13864, ZN => n5230);
   U4375 : MUX2_X1 port map( A => n13401, B => n13400, S => n14225, Z => n13402
                           );
   U4376 : INV_X1 port map( A => n15802, ZN => n16075);
   U4377 : INV_X1 port map( A => n16394, ZN => n16167);
   U4378 : AND2_X1 port map( A1 => n15198, A2 => n3554, ZN => n3553);
   U4379 : XNOR2_X1 port map( A => n2862, B => n14555, ZN => n16151);
   U4380 : INV_X1 port map( A => n16312, ZN => n16309);
   U4381 : OR2_X1 port map( A1 => n4869, A2 => n15647, ZN => n4575);
   U4382 : INV_X1 port map( A => n15640, ZN => n3380);
   U4383 : INV_X1 port map( A => n17183, ZN => n16204);
   U4384 : XNOR2_X1 port map( A => n4967, B => n4965, ZN => n16422);
   U4385 : XNOR2_X1 port map( A => n14428, B => n4966, ZN => n4965);
   U4386 : NOR2_X1 port map( A1 => n24981, A2 => n5039, ZN => n5038);
   U4387 : AND2_X1 port map( A1 => n16481, A2 => n16480, ZN => n5039);
   U4388 : AOI22_X1 port map( A1 => n16495, A2 => n16494, B1 => n16493, B2 => 
                           n16492, ZN => n16516);
   U4389 : OAI211_X1 port map( C1 => n16104, C2 => n16105, A => n3409, B => 
                           n3408, ZN => n17524);
   U4390 : OR2_X1 port map( A1 => n16103, A2 => n3410, ZN => n3409);
   U4391 : INV_X1 port map( A => n17524, ZN => n16863);
   U4392 : OR2_X1 port map( A1 => n16798, A2 => n5375, ZN => n5240);
   U4393 : XNOR2_X1 port map( A => n17814, B => n18562, ZN => n17815);
   U4394 : INV_X1 port map( A => n1653, ZN => n17144);
   U4395 : NAND3_X1 port map( A1 => n16468, A2 => n4725, A3 => n4724, ZN => 
                           n16984);
   U4397 : OR2_X1 port map( A1 => n15796, A2 => n382, ZN => n4858);
   U4398 : INV_X1 port map( A => n17515, ZN => n18258);
   U4399 : OR2_X1 port map( A1 => n19520, A2 => n19284, ZN => n4433);
   U4401 : XNOR2_X1 port map( A => n1386, B => n17092, ZN => n4214);
   U4403 : NAND2_X1 port map( A1 => n18840, A2 => n19322, ZN => n3584);
   U4404 : OR2_X1 port map( A1 => n18961, A2 => n19467, ZN => n3579);
   U4405 : INV_X1 port map( A => n17567, ZN => n19714);
   U4406 : OR2_X1 port map( A1 => n20203, A2 => n20204, ZN => n1664);
   U4407 : XNOR2_X1 port map( A => n3823, B => n21043, ZN => n21229);
   U4408 : XNOR2_X1 port map( A => n21266, B => n24485, ZN => n3746);
   U4410 : OR2_X1 port map( A1 => n20368, A2 => n24454, ZN => n20303);
   U4411 : XNOR2_X1 port map( A => n19161, B => n19160, ZN => n22255);
   U4412 : OR2_X1 port map( A1 => n6034, A2 => n441, ZN => n6171);
   U4414 : INV_X1 port map( A => n7782, ZN => n7174);
   U4415 : AND2_X1 port map( A1 => n2974, A2 => n2973, ZN => n6613);
   U4416 : INV_X1 port map( A => n7991, ZN => n7357);
   U4418 : INV_X1 port map( A => n8132, ZN => n8845);
   U4419 : INV_X1 port map( A => n8428, ZN => n4335);
   U4420 : XNOR2_X1 port map( A => n8476, B => n2191, ZN => n4395);
   U4422 : NAND2_X1 port map( A1 => n1693, A2 => n1692, ZN => n7234);
   U4423 : AND2_X1 port map( A1 => n7004, A2 => n448, ZN => n5148);
   U4424 : OR2_X1 port map( A1 => n7892, A2 => n7322, ZN => n3082);
   U4425 : XNOR2_X1 port map( A => n8730, B => n8468, ZN => n8797);
   U4427 : OR2_X1 port map( A1 => n9220, A2 => n9705, ZN => n3721);
   U4428 : NAND2_X1 port map( A1 => n7532, A2 => n7533, ZN => n1972);
   U4429 : INV_X1 port map( A => n8476, ZN => n4401);
   U4430 : OR2_X1 port map( A1 => n9127, A2 => n10063, ZN => n9220);
   U4431 : NOR2_X1 port map( A1 => n1517, A2 => n24549, ZN => n9876);
   U4432 : INV_X1 port map( A => n10138, ZN => n1649);
   U4433 : OR2_X1 port map( A1 => n10099, A2 => n9515, ZN => n10097);
   U4434 : OAI21_X1 port map( B1 => n2267, B2 => n9615, A => n1412, ZN => n3546
                           );
   U4435 : OR2_X1 port map( A1 => n9754, A2 => n9613, ZN => n1412);
   U4436 : AND2_X1 port map( A1 => n10161, A2 => n24984, ZN => n9382);
   U4437 : BUF_X1 port map( A => n9515, Z => n10098);
   U4440 : XNOR2_X1 port map( A => n8806, B => n1831, ZN => n2491);
   U4441 : NOR2_X1 port map( A1 => n4254, A2 => n25393, ZN => n3865);
   U4443 : AND2_X1 port map( A1 => n13049, A2 => n13048, ZN => n1545);
   U4444 : AND2_X1 port map( A1 => n2524, A2 => n2523, ZN => n10312);
   U4445 : INV_X1 port map( A => n3375, ZN => n11307);
   U4446 : AND2_X1 port map( A1 => n11012, A2 => n11045, ZN => n10415);
   U4447 : INV_X1 port map( A => n2295, ZN => n13327);
   U4448 : OR2_X1 port map( A1 => n13076, A2 => n3704, ZN => n13080);
   U4449 : INV_X1 port map( A => n3492, ZN => n4405);
   U4450 : OR2_X1 port map( A1 => n10711, A2 => n13132, ZN => n13158);
   U4451 : XNOR2_X1 port map( A => n11546, B => n11547, ZN => n12773);
   U4452 : INV_X1 port map( A => n11981, ZN => n4931);
   U4453 : INV_X1 port map( A => n12934, ZN => n5361);
   U4456 : OAI211_X1 port map( C1 => n13104, C2 => n13103, A => n12658, B => 
                           n12657, ZN => n12668);
   U4457 : INV_X1 port map( A => n3958, ZN => n12654);
   U4458 : XNOR2_X1 port map( A => n11760, B => n4134, ZN => n13223);
   U4459 : OR2_X1 port map( A1 => n3460, A2 => n3492, ZN => n5325);
   U4460 : XNOR2_X1 port map( A => n11268, B => n3900, ZN => n11626);
   U4461 : NOR2_X1 port map( A1 => n12583, A2 => n24554, ZN => n12624);
   U4462 : OR2_X1 port map( A1 => n13122, A2 => n5626, ZN => n2516);
   U4463 : OR2_X1 port map( A1 => n12873, A2 => n13123, ZN => n2515);
   U4465 : OR2_X1 port map( A1 => n12452, A2 => n304, ZN => n3523);
   U4466 : OR2_X1 port map( A1 => n12453, A2 => n4766, ZN => n3524);
   U4467 : OR2_X1 port map( A1 => n13025, A2 => n13030, ZN => n1634);
   U4469 : NOR2_X1 port map( A1 => n4790, A2 => n4789, ZN => n4788);
   U4470 : AND2_X1 port map( A1 => n4791, A2 => n3858, ZN => n3860);
   U4472 : OR2_X1 port map( A1 => n5359, A2 => n4499, ZN => n2715);
   U4473 : AND2_X1 port map( A1 => n12610, A2 => n1971, ZN => n1970);
   U4474 : OR2_X1 port map( A1 => n12606, A2 => n12683, ZN => n2840);
   U4475 : OAI21_X1 port map( B1 => n12965, B2 => n3813, A => n13273, ZN => 
                           n2158);
   U4476 : INV_X1 port map( A => n14167, ZN => n14164);
   U4478 : OR2_X1 port map( A1 => n4529, A2 => n12634, ZN => n2721);
   U4479 : AOI21_X1 port map( B1 => n14067, B2 => n13845, A => n13627, ZN => 
                           n12592);
   U4480 : INV_X1 port map( A => n15556, ZN => n2173);
   U4481 : AND3_X1 port map( A1 => n14327, A2 => n14044, A3 => n13864, ZN => 
                           n2225);
   U4482 : NOR2_X1 port map( A1 => n4870, A2 => n24062, ZN => n4869);
   U4484 : OR2_X1 port map( A1 => n16206, A2 => n15640, ZN => n16207);
   U4485 : AND2_X1 port map( A1 => n16324, A2 => n2610, ZN => n16194);
   U4486 : AOI22_X1 port map( A1 => n388, A2 => n290, B1 => n1123, B2 => n16331
                           , ZN => n16185);
   U4487 : XNOR2_X1 port map( A => n15237, B => n15236, ZN => n15674);
   U4488 : OAI21_X1 port map( B1 => n386, B2 => n15992, A => n15991, ZN => 
                           n4646);
   U4489 : INV_X1 port map( A => n15839, ZN => n16175);
   U4490 : XNOR2_X1 port map( A => n5757, B => n13424, ZN => n15915);
   U4491 : XNOR2_X1 port map( A => n4712, B => n3694, ZN => n16418);
   U4492 : INV_X1 port map( A => n16246, ZN => n16253);
   U4493 : AND2_X1 port map( A1 => n25484, A2 => n15764, ZN => n15940);
   U4496 : INV_X1 port map( A => n16418, ZN => n16413);
   U4497 : INV_X1 port map( A => n15842, ZN => n2996);
   U4499 : XNOR2_X1 port map( A => n14592, B => n1383, ZN => n4205);
   U4500 : XNOR2_X1 port map( A => n4095, B => n14593, ZN => n4204);
   U4501 : INV_X1 port map( A => n2253, ZN => n2251);
   U4503 : OAI21_X1 port map( B1 => n16274, B2 => n16029, A => n2280, ZN => 
                           n16034);
   U4504 : AOI22_X1 port map( A1 => n16133, A2 => n16075, B1 => n16132, B2 => 
                           n16131, ZN => n16431);
   U4505 : OR2_X1 port map( A1 => n15983, A2 => n16163, ZN => n3008);
   U4507 : NAND3_X1 port map( A1 => n16146, A2 => n2541, A3 => n16098, ZN => 
                           n16434);
   U4508 : AOI22_X1 port map( A1 => n16838, A2 => n16261, B1 => n16533, B2 => 
                           n17165, ZN => n16378);
   U4509 : XNOR2_X1 port map( A => n17811, B => n17969, ZN => n18248);
   U4511 : INV_X1 port map( A => n17815, ZN => n18287);
   U4512 : INV_X1 port map( A => n19278, ZN => n5573);
   U4513 : XNOR2_X1 port map( A => n17639, B => n18051, ZN => n18734);
   U4514 : XNOR2_X1 port map( A => n18578, B => n18577, ZN => n18998);
   U4515 : AND2_X1 port map( A1 => n18998, A2 => n19418, ZN => n19002);
   U4516 : INV_X1 port map( A => n19488, ZN => n19346);
   U4517 : AND2_X1 port map( A1 => n18734, A2 => n19476, ZN => n5685);
   U4518 : XNOR2_X1 port map( A => n18354, B => n18353, ZN => n18385);
   U4519 : INV_X1 port map( A => n18998, ZN => n19421);
   U4520 : OR2_X1 port map( A1 => n19413, A2 => n25469, ZN => n19409);
   U4521 : XNOR2_X1 port map( A => n2692, B => n17777, ZN => n2029);
   U4522 : XNOR2_X1 port map( A => n18681, B => n18682, ZN => n19408);
   U4524 : XNOR2_X1 port map( A => n18123, B => n23191, ZN => n18438);
   U4526 : OR2_X1 port map( A1 => n18907, A2 => n19568, ZN => n2512);
   U4527 : XNOR2_X1 port map( A => n4268, B => n18363, ZN => n4274);
   U4528 : INV_X1 port map( A => n18520, ZN => n16600);
   U4529 : XNOR2_X1 port map( A => n4808, B => n17375, ZN => n17376);
   U4530 : OR2_X1 port map( A1 => n25423, A2 => n19436, ZN => n5007);
   U4531 : AND2_X1 port map( A1 => n357, A2 => n19500, ZN => n18986);
   U4532 : XNOR2_X1 port map( A => n18175, B => n18174, ZN => n19520);
   U4533 : AND2_X1 port map( A1 => n5572, A2 => n2626, ZN => n20258);
   U4534 : AND2_X1 port map( A1 => n19540, A2 => n19126, ZN => n2626);
   U4535 : OR2_X1 port map( A1 => n2132, A2 => n24477, ZN => n4542);
   U4536 : XNOR2_X1 port map( A => n21164, B => n21165, ZN => n1605);
   U4537 : XNOR2_X1 port map( A => n4908, B => n21532, ZN => n17951);
   U4538 : INV_X1 port map( A => n21481, ZN => n4908);
   U4539 : AOI21_X1 port map( B1 => n22609, B2 => n22813, A => n4272, ZN => 
                           n22610);
   U4540 : NOR2_X1 port map( A1 => n22495, A2 => n22494, ZN => n4719);
   U4541 : OR2_X1 port map( A1 => n21822, A2 => n22257, ZN => n2987);
   U4542 : INV_X1 port map( A => n22255, ZN => n4373);
   U4543 : OAI21_X1 port map( B1 => n3741, B2 => n22811, A => n22813, ZN => 
                           n3740);
   U4544 : XNOR2_X1 port map( A => n20697, B => n5286, ZN => n20465);
   U4546 : OR2_X1 port map( A1 => n6688, A2 => n4830, ZN => n4829);
   U4547 : INV_X1 port map( A => n6648, ZN => n7006);
   U4548 : XNOR2_X1 port map( A => Plaintext(122), B => Key(122), ZN => n6648);
   U4549 : OR2_X1 port map( A1 => n6396, A2 => n6732, ZN => n4178);
   U4550 : NAND2_X1 port map( A1 => n6607, A2 => n6606, ZN => n1926);
   U4552 : OR2_X1 port map( A1 => n6528, A2 => n6529, ZN => n4681);
   U4553 : OR2_X1 port map( A1 => n6165, A2 => n7101, ZN => n6545);
   U4554 : OR2_X1 port map( A1 => n8022, A2 => n8021, ZN => n1840);
   U4555 : OAI21_X1 port map( B1 => n6094, B2 => n7006, A => n7005, ZN => n2879
                           );
   U4556 : AND2_X1 port map( A1 => n442, A2 => n7026, ZN => n5089);
   U4558 : INV_X1 port map( A => n5924, ZN => n3922);
   U4559 : AND2_X1 port map( A1 => n7776, A2 => n7767, ZN => n1786);
   U4561 : INV_X1 port map( A => n6805, ZN => n7665);
   U4562 : INV_X1 port map( A => n8782, ZN => n8537);
   U4563 : OR2_X1 port map( A1 => n7456, A2 => n311, ZN => n5161);
   U4564 : INV_X1 port map( A => n7257, ZN => n7341);
   U4565 : NAND2_X1 port map( A1 => n6537, A2 => n4744, ZN => n7664);
   U4566 : INV_X1 port map( A => n8336, ZN => n8172);
   U4567 : OR2_X1 port map( A1 => n4136, A2 => n4002, ZN => n4001);
   U4568 : NAND2_X1 port map( A1 => n4883, A2 => n7068, ZN => n2560);
   U4569 : OAI21_X1 port map( B1 => n7221, B2 => n7064, A => n431, ZN => n4883)
                           ;
   U4570 : NAND2_X1 port map( A1 => n5636, A2 => n5635, ZN => n7629);
   U4571 : NAND3_X1 port map( A1 => n4377, A2 => n7538, A3 => n7539, ZN => 
                           n9007);
   U4572 : XNOR2_X1 port map( A => n8150, B => n5504, ZN => n8157);
   U4573 : XNOR2_X1 port map( A => n4395, B => n8342, ZN => n8343);
   U4574 : XNOR2_X1 port map( A => n8612, B => n8981, ZN => n8889);
   U4575 : XNOR2_X1 port map( A => n7119, B => n7120, ZN => n9955);
   U4576 : INV_X1 port map( A => n9012, ZN => n8665);
   U4577 : XNOR2_X1 port map( A => n8451, B => n8454, ZN => n1906);
   U4578 : INV_X1 port map( A => n9335, ZN => n9334);
   U4579 : XNOR2_X1 port map( A => n8183, B => n3507, ZN => n3506);
   U4581 : AND2_X1 port map( A1 => n25207, A2 => n10149, ZN => n2740);
   U4582 : XNOR2_X1 port map( A => n8336, B => n1528, ZN => n8070);
   U4584 : INV_X1 port map( A => n9829, ZN => n10178);
   U4585 : INV_X1 port map( A => n10614, ZN => n10488);
   U4586 : INV_X1 port map( A => n9244, ZN => n9866);
   U4587 : XNOR2_X1 port map( A => n9079, B => n9078, ZN => n10050);
   U4588 : XNOR2_X1 port map( A => n2446, B => n8087, ZN => n9692);
   U4589 : OR2_X1 port map( A1 => n9454, A2 => n8157, ZN => n9566);
   U4590 : OR2_X1 port map( A1 => n9219, A2 => n10060, ZN => n5608);
   U4591 : INV_X1 port map( A => n9515, ZN => n4300);
   U4592 : AND2_X1 port map( A1 => n10100, A2 => n9837, ZN => n9327);
   U4593 : NOR2_X1 port map( A1 => n10406, A2 => n10405, ZN => n10992);
   U4594 : INV_X1 port map( A => n11036, ZN => n5392);
   U4596 : INV_X1 port map( A => n10935, ZN => n10508);
   U4597 : NAND3_X1 port map( A1 => n1671, A2 => n1670, A3 => n1668, ZN => 
                           n4422);
   U4598 : OR2_X1 port map( A1 => n9436, A2 => n9435, ZN => n1670);
   U4599 : NAND2_X1 port map( A1 => n1669, A2 => n9434, ZN => n1668);
   U4600 : INV_X1 port map( A => n9382, ZN => n5105);
   U4601 : OR2_X1 port map( A1 => n10172, A2 => n25, ZN => n4212);
   U4602 : OR2_X1 port map( A1 => n9815, A2 => n2207, ZN => n2548);
   U4603 : AND3_X1 port map( A1 => n10753, A2 => n2866, A3 => n2865, ZN => 
                           n10760);
   U4604 : NAND2_X1 port map( A1 => n2268, A2 => n9976, ZN => n10416);
   U4605 : AND2_X1 port map( A1 => n25499, A2 => n12942, ZN => n2918);
   U4606 : OR2_X1 port map( A1 => n3387, A2 => n10590, ZN => n10591);
   U4607 : INV_X1 port map( A => n11704, ZN => n3812);
   U4608 : XNOR2_X1 port map( A => n1388, B => n12340, ZN => n13353);
   U4609 : OAI21_X1 port map( B1 => n4462, B2 => n420, A => n4464, ZN => n4461)
                           ;
   U4610 : INV_X1 port map( A => n12613, ZN => n3859);
   U4611 : OR2_X1 port map( A1 => n10623, A2 => n11212, ZN => n10624);
   U4612 : XNOR2_X1 port map( A => n11820, B => n11819, ZN => n13301);
   U4613 : INV_X1 port map( A => n405, ZN => n4493);
   U4614 : AND2_X1 port map( A1 => n13245, A2 => n13014, ZN => n13018);
   U4615 : NOR2_X1 port map( A1 => n25198, A2 => n13014, ZN => n13016);
   U4616 : XNOR2_X1 port map( A => n11661, B => n3208, ZN => n11248);
   U4617 : AND2_X1 port map( A1 => n13228, A2 => n11328, ZN => n2291);
   U4618 : AND3_X1 port map( A1 => n12612, A2 => n3859, A3 => n13303, ZN => 
                           n4790);
   U4619 : OR2_X1 port map( A1 => n13018, A2 => n13017, ZN => n3558);
   U4620 : BUF_X1 port map( A => n13037, Z => n13044);
   U4621 : OR2_X1 port map( A1 => n13076, A2 => n12713, ZN => n2192);
   U4622 : INV_X1 port map( A => n24573, ZN => n3590);
   U4624 : AND3_X1 port map( A1 => n25494, A2 => n13051, A3 => n4094, ZN => 
                           n13086);
   U4625 : INV_X1 port map( A => n13998, ZN => n13993);
   U4626 : INV_X1 port map( A => n12897, ZN => n4861);
   U4627 : INV_X1 port map( A => n25248, ZN => n2437);
   U4628 : XNOR2_X1 port map( A => n10198, B => n10197, ZN => n3492);
   U4629 : OAI21_X1 port map( B1 => n12483, B2 => n12711, A => n4060, ZN => 
                           n4059);
   U4630 : AND2_X1 port map( A1 => n13989, A2 => n13918, ZN => n13984);
   U4631 : OR2_X1 port map( A1 => n4729, A2 => n3766, ZN => n2423);
   U4632 : OR2_X1 port map( A1 => n12899, A2 => n13279, ZN => n11867);
   U4633 : INV_X1 port map( A => n4241, ZN => n12946);
   U4634 : XNOR2_X1 port map( A => n11835, B => n11834, ZN => n12902);
   U4635 : OR3_X1 port map( A1 => n13222, A2 => n24965, A3 => n13227, ZN => 
                           n4484);
   U4636 : INV_X1 port map( A => n14150, ZN => n5102);
   U4637 : INV_X1 port map( A => n12767, ZN => n2493);
   U4638 : INV_X1 port map( A => n13216, ZN => n12986);
   U4639 : AOI22_X1 port map( A1 => n13009, A2 => n11754, B1 => n13221, B2 => 
                           n12885, ZN => n13010);
   U4642 : OR2_X1 port map( A1 => n2608, A2 => n2837, ZN => n12567);
   U4643 : AND2_X1 port map( A1 => n13796, A2 => n13792, ZN => n13579);
   U4644 : AND2_X1 port map( A1 => n3788, A2 => n3786, ZN => n3787);
   U4645 : OAI211_X1 port map( C1 => n14268, C2 => n123, A => n14267, B => 
                           n3789, ZN => n3788);
   U4646 : AND2_X1 port map( A1 => n13884, A2 => n13597, ZN => n13596);
   U4647 : OR2_X1 port map( A1 => n12918, A2 => n24490, ZN => n12570);
   U4648 : INV_X1 port map( A => n14048, ZN => n14050);
   U4649 : OAI21_X1 port map( B1 => n12426, B2 => n12666, A => n10787, ZN => 
                           n13953);
   U4650 : OR2_X1 port map( A1 => n12437, A2 => n13138, ZN => n2929);
   U4651 : OAI21_X1 port map( B1 => n5013, B2 => n25061, A => n13162, ZN => 
                           n5012);
   U4652 : OR2_X1 port map( A1 => n13164, A2 => n13163, ZN => n4867);
   U4653 : AND2_X1 port map( A1 => n4868, A2 => n14112, ZN => n13581);
   U4654 : AND2_X1 port map( A1 => n13485, A2 => n12669, ZN => n13262);
   U4655 : OR2_X1 port map( A1 => n14944, A2 => n25458, ZN => n14144);
   U4656 : INV_X1 port map( A => n14826, ZN => n15111);
   U4657 : INV_X1 port map( A => n13597, ZN => n13724);
   U4658 : OR2_X1 port map( A1 => n1578, A2 => n12555, ZN => n12556);
   U4659 : AND2_X1 port map( A1 => n5140, A2 => n4634, ZN => n12072);
   U4660 : AND2_X1 port map( A1 => n13325, A2 => n13323, ZN => n5140);
   U4661 : INV_X1 port map( A => n14325, ZN => n14330);
   U4663 : INV_X1 port map( A => n14221, ZN => n4019);
   U4664 : INV_X1 port map( A => n13829, ZN => n14119);
   U4665 : INV_X1 port map( A => n13966, ZN => n13883);
   U4666 : INV_X1 port map( A => n13997, ZN => n14235);
   U4667 : INV_X1 port map( A => n13682, ZN => n14233);
   U4668 : AND2_X1 port map( A1 => n14204, A2 => n3341, ZN => n13814);
   U4669 : AND2_X1 port map( A1 => n13446, A2 => n13445, ZN => n2863);
   U4670 : OAI21_X1 port map( B1 => n13819, B2 => n13385, A => n13646, ZN => 
                           n2658);
   U4671 : AND2_X1 port map( A1 => n1790, A2 => n16051, ZN => n15540);
   U4672 : OR2_X1 port map( A1 => n13440, A2 => n14101, ZN => n4598);
   U4673 : XNOR2_X1 port map( A => n14391, B => n15452, ZN => n15093);
   U4674 : XNOR2_X1 port map( A => n14358, B => n14357, ZN => n15842);
   U4675 : XNOR2_X1 port map( A => n13450, B => n3787, ZN => n3471);
   U4676 : XNOR2_X1 port map( A => n15177, B => n5216, ZN => n14964);
   U4677 : OR2_X1 port map( A1 => n13676, A2 => n5221, ZN => n13489);
   U4678 : OAI21_X1 port map( B1 => n13484, B2 => n13487, A => n3071, ZN => 
                           n4415);
   U4679 : INV_X1 port map( A => n16368, ZN => n15814);
   U4680 : OR2_X1 port map( A1 => n15940, A2 => n2605, ZN => n2604);
   U4681 : INV_X1 port map( A => n4765, ZN => n14201);
   U4683 : AOI22_X1 port map( A1 => n1621, A2 => n16285, B1 => n15747, B2 => 
                           n24539, ZN => n17623);
   U4684 : INV_X1 port map( A => n5376, ZN => n16622);
   U4685 : OAI21_X1 port map( B1 => n16481, B2 => n15953, A => n15696, ZN => 
                           n5495);
   U4686 : OAI21_X1 port map( B1 => n25238, B2 => n15695, A => n16483, ZN => 
                           n5493);
   U4687 : AND2_X1 port map( A1 => n17276, A2 => n17254, ZN => n17247);
   U4688 : AND2_X1 port map( A1 => n16368, A2 => n17183, ZN => n17181);
   U4690 : OR2_X1 port map( A1 => n2549, A2 => n17442, ZN => n16961);
   U4691 : OR2_X1 port map( A1 => n17356, A2 => n17351, ZN => n5366);
   U4692 : AND2_X1 port map( A1 => n24942, A2 => n17450, ZN => n17152);
   U4693 : INV_X1 port map( A => n3604, ZN => n3598);
   U4694 : OAI21_X1 port map( B1 => n16411, B2 => n3061, A => n3060, ZN => 
                           n16421);
   U4695 : INV_X1 port map( A => n17050, ZN => n2613);
   U4697 : AND2_X1 port map( A1 => n16323, A2 => n25447, ZN => n15258);
   U4698 : AND2_X1 port map( A1 => n4541, A2 => n15604, ZN => n15693);
   U4699 : OAI22_X1 port map( A1 => n4482, A2 => n17356, B1 => n16316, B2 => 
                           n367, ZN => n16318);
   U4700 : NAND3_X1 port map( A1 => n16758, A2 => n16757, A3 => n2324, ZN => 
                           n17931);
   U4701 : OR2_X1 port map( A1 => n15602, A2 => n16060, ZN => n1673);
   U4702 : INV_X1 port map( A => n18646, ZN => n18552);
   U4703 : NOR2_X1 port map( A1 => n16671, A2 => n2530, ZN => n2937);
   U4705 : OR2_X1 port map( A1 => n16978, A2 => n17336, ZN => n4246);
   U4706 : OR2_X1 port map( A1 => n16431, A2 => n16434, ZN => n16522);
   U4707 : NOR2_X1 port map( A1 => n5522, A2 => n17572, ZN => n3004);
   U4708 : AND2_X1 port map( A1 => n1616, A2 => n1615, ZN => n16719);
   U4709 : OR2_X1 port map( A1 => n17025, A2 => n17389, ZN => n1852);
   U4710 : OR2_X1 port map( A1 => n4566, A2 => n17602, ZN => n4565);
   U4711 : AOI21_X1 port map( B1 => n4564, B2 => n4563, A => n2968, ZN => n4562
                           );
   U4712 : OAI21_X1 port map( B1 => n3956, B2 => n25215, A => n3948, ZN => 
                           n18254);
   U4714 : AOI21_X1 port map( B1 => n3458, B2 => n3457, A => n3391, ZN => n3390
                           );
   U4715 : AND2_X1 port map( A1 => n25226, A2 => n25245, ZN => n3391);
   U4717 : INV_X1 port map( A => n18123, ZN => n18437);
   U4718 : INV_X1 port map( A => n19077, ZN => n18862);
   U4719 : OR3_X1 port map( A1 => n25245, A2 => n17131, A3 => n25226, ZN => 
                           n15806);
   U4720 : OR2_X1 port map( A1 => n17418, A2 => n17419, ZN => n2054);
   U4721 : NAND2_X1 port map( A1 => n2183, A2 => n2110, ZN => n17811);
   U4722 : AND2_X1 port map( A1 => n17198, A2 => n17395, ZN => n2112);
   U4723 : XNOR2_X1 port map( A => n18397, B => n17520, ZN => n18627);
   U4724 : OAI21_X1 port map( B1 => n17461, B2 => n288, A => n17464, ZN => 
                           n5158);
   U4725 : XNOR2_X1 port map( A => n3703, B => n18187, ZN => n18291);
   U4726 : AOI22_X1 port map( A1 => n3930, A2 => n16985, B1 => n3929, B2 => 
                           n17144, ZN => n3928);
   U4727 : OR2_X1 port map( A1 => n3432, A2 => n17053, ZN => n3431);
   U4728 : OR2_X1 port map( A1 => n16895, A2 => n2372, ZN => n2373);
   U4729 : AOI21_X1 port map( B1 => n5386, B2 => n17479, A => n2181, ZN => 
                           n2374);
   U4730 : INV_X1 port map( A => n16513, ZN => n16618);
   U4731 : OR2_X1 port map( A1 => n16703, A2 => n16705, ZN => n16617);
   U4732 : XNOR2_X1 port map( A => n24536, B => n17757, ZN => n18363);
   U4733 : NAND2_X1 port map( A1 => n4304, A2 => n16908, ZN => n2583);
   U4734 : NAND3_X1 port map( A1 => n16182, A2 => n16181, A3 => n5017, ZN => 
                           n17863);
   U4735 : AND2_X1 port map( A1 => n16984, A2 => n16985, ZN => n2161);
   U4736 : AND2_X1 port map( A1 => n17122, A2 => n17114, ZN => n16801);
   U4737 : AND2_X1 port map( A1 => n25422, A2 => n19436, ZN => n3985);
   U4738 : NOR2_X1 port map( A1 => n1427, A2 => n5573, ZN => n5569);
   U4739 : INV_X1 port map( A => n20192, ZN => n5208);
   U4740 : XNOR2_X1 port map( A => n21160, B => n21750, ZN => n21163);
   U4741 : XNOR2_X1 port map( A => n21266, B => n21160, ZN => n21611);
   U4742 : OAI211_X1 port map( C1 => n20220, C2 => n20510, A => n1809, B => 
                           n1808, ZN => n21495);
   U4743 : INV_X1 port map( A => n19710, ZN => n4713);
   U4748 : OAI22_X1 port map( A1 => n5499, A2 => n25345, B1 => n2606, B2 => 
                           n20214, ZN => n20513);
   U4750 : NAND2_X1 port map( A1 => n20207, A2 => n4264, ZN => n4263);
   U4751 : AND2_X1 port map( A1 => n20206, A2 => n4265, ZN => n4264);
   U4753 : OR2_X1 port map( A1 => n20548, A2 => n20124, ZN => n4569);
   U4754 : INV_X1 port map( A => n22721, ZN => n2711);
   U4755 : INV_X1 port map( A => n20336, ZN => n19708);
   U4756 : INV_X1 port map( A => n20459, ZN => n4489);
   U4757 : OAI22_X1 port map( A1 => n20128, A2 => n20130, B1 => n20130, B2 => 
                           n20129, ZN => n5491);
   U4758 : AND2_X1 port map( A1 => n21523, A2 => n2563, ZN => n20926);
   U4759 : INV_X1 port map( A => n3115, ZN => n2563);
   U4761 : NOR2_X1 port map( A1 => n19984, A2 => n19983, ZN => n2098);
   U4762 : OR2_X1 port map( A1 => n20117, A2 => n20116, ZN => n2873);
   U4763 : OR2_X1 port map( A1 => n20114, A2 => n20111, ZN => n2874);
   U4764 : XNOR2_X1 port map( A => n21599, B => n21520, ZN => n21192);
   U4765 : XNOR2_X1 port map( A => n21550, B => n21981, ZN => n21209);
   U4766 : NOR2_X1 port map( A1 => n25383, A2 => n2431, ZN => n20375);
   U4767 : OR2_X1 port map( A1 => n20374, A2 => n2432, ZN => n2431);
   U4768 : OR2_X1 port map( A1 => n19682, A2 => n20302, ZN => n2135);
   U4770 : NAND3_X1 port map( A1 => n19986, A2 => n19987, A3 => n21068, ZN => 
                           n3963);
   U4772 : XNOR2_X1 port map( A => n22006, B => n25400, ZN => n4396);
   U4773 : XNOR2_X1 port map( A => n2465, B => n25483, ZN => n20745);
   U4774 : XNOR2_X1 port map( A => n21699, B => n23183, ZN => n2465);
   U4775 : INV_X1 port map( A => n329, ZN => n5224);
   U4776 : XNOR2_X1 port map( A => n20972, B => n20678, ZN => n4100);
   U4777 : NOR2_X1 port map( A1 => n22209, A2 => n22064, ZN => n22092);
   U4778 : XNOR2_X1 port map( A => n21724, B => n21723, ZN => n2633);
   U4781 : XNOR2_X1 port map( A => n21737, B => n21734, ZN => n4687);
   U4782 : OR2_X1 port map( A1 => n23016, A2 => n23014, ZN => n22914);
   U4783 : XNOR2_X1 port map( A => n20918, B => n1628, ZN => n2315);
   U4784 : INV_X1 port map( A => n21538, ZN => n1628);
   U4785 : INV_X1 port map( A => n22227, ZN => n3231);
   U4786 : OR2_X1 port map( A1 => n22228, A2 => n22231, ZN => n3230);
   U4787 : XNOR2_X1 port map( A => n20324, B => n3746, ZN => n4169);
   U4788 : OR2_X1 port map( A1 => n22770, A2 => n5378, ZN => n5377);
   U4789 : INV_X1 port map( A => n22812, ZN => n4469);
   U4790 : OR2_X1 port map( A1 => n5712, A2 => n21856, ZN => n22772);
   U4794 : NAND4_X1 port map( A1 => n23202, A2 => n22569, A3 => n24889, A4 => 
                           n22561, ZN => n4237);
   U4795 : AND2_X1 port map( A1 => n23805, A2 => n24895, ZN => n2591);
   U4797 : INV_X1 port map( A => n3856, ZN => n19625);
   U4798 : INV_X1 port map( A => n23843, ZN => n23862);
   U4799 : INV_X1 port map( A => n6733, ZN => n2119);
   U4800 : XNOR2_X1 port map( A => n5847, B => Key(161), ZN => n6770);
   U4801 : OR2_X1 port map( A1 => n6297, A2 => n6438, ZN => n5946);
   U4802 : AOI21_X1 port map( B1 => n6703, B2 => n24405, A => n6959, ZN => 
                           n4324);
   U4803 : INV_X1 port map( A => n8021, ZN => n7531);
   U4804 : OR2_X1 port map( A1 => n6162, A2 => n6265, ZN => n2534);
   U4805 : OR2_X1 port map( A1 => n5910, A2 => n5887, ZN => n4503);
   U4807 : OAI21_X1 port map( B1 => n6771, B2 => n24037, A => n6770, ZN => 
                           n6772);
   U4808 : INV_X1 port map( A => n4672, ZN => n7945);
   U4809 : OR2_X1 port map( A1 => n7858, A2 => n7857, ZN => n4976);
   U4810 : INV_X1 port map( A => n7413, ZN => n4827);
   U4811 : NOR2_X1 port map( A1 => n5824, A2 => n6473, ZN => n6899);
   U4812 : OAI21_X1 port map( B1 => n5975, B2 => n6987, A => n5974, ZN => n5978
                           );
   U4813 : AND2_X1 port map( A1 => n5798, A2 => n5799, ZN => n7481);
   U4814 : OR2_X1 port map( A1 => n7861, A2 => n7862, ZN => n3571);
   U4815 : INV_X1 port map( A => n7781, ZN => n7419);
   U4816 : AND3_X1 port map( A1 => n3588, A2 => n3344, A3 => n7531, ZN => n3587
                           );
   U4817 : AND2_X1 port map( A1 => n4708, A2 => n4711, ZN => n4707);
   U4818 : AND3_X1 port map( A1 => n7930, A2 => n7931, A3 => n7929, ZN => n4545
                           );
   U4819 : INV_X1 port map( A => n2402, ZN => n8024);
   U4820 : OR2_X1 port map( A1 => n6768, A2 => n6767, ZN => n2976);
   U4821 : INV_X1 port map( A => n7335, ZN => n7592);
   U4823 : OR2_X1 port map( A1 => n6494, A2 => n6493, ZN => n1575);
   U4825 : OAI211_X1 port map( C1 => n1468, C2 => n4376, A => n7079, B => n4375
                           , ZN => n8452);
   U4826 : OR2_X1 port map( A1 => n6040, A2 => n6165, ZN => n6041);
   U4827 : INV_X1 port map( A => n8960, ZN => n8908);
   U4828 : OAI211_X1 port map( C1 => n6752, C2 => n6674, A => n6578, B => n1807
                           , ZN => n2495);
   U4829 : OR2_X1 port map( A1 => n6400, A2 => n6757, ZN => n1807);
   U4830 : INV_X1 port map( A => n6572, ZN => n6058);
   U4831 : OR2_X1 port map( A1 => n6059, A2 => n6967, ZN => n3838);
   U4832 : AND2_X1 port map( A1 => n2355, A2 => n1175, ZN => n2349);
   U4833 : INV_X1 port map( A => n6314, ZN => n5452);
   U4834 : OR2_X1 port map( A1 => n6233, A2 => n6715, ZN => n6110);
   U4835 : XNOR2_X1 port map( A => n8721, B => n2272, ZN => n8756);
   U4836 : INV_X1 port map( A => n8755, ZN => n2272);
   U4837 : OAI21_X1 port map( B1 => n7045, B2 => n7174, A => n3496, ZN => n8812
                           );
   U4838 : OAI21_X1 port map( B1 => n5606, B2 => n5605, A => n5607, ZN => n5603
                           );
   U4839 : AND2_X1 port map( A1 => n7157, A2 => n7156, ZN => n5345);
   U4840 : INV_X1 port map( A => n7364, ZN => n7911);
   U4841 : INV_X1 port map( A => n7629, ZN => n7910);
   U4842 : INV_X1 port map( A => n3979, ZN => n8371);
   U4843 : OR2_X1 port map( A1 => n6413, A2 => n7721, ZN => n1879);
   U4844 : OR2_X1 port map( A1 => n7115, A2 => n7761, ZN => n5691);
   U4845 : INV_X1 port map( A => n2145, ZN => n5690);
   U4847 : INV_X1 port map( A => n6549, ZN => n7671);
   U4848 : AND2_X1 port map( A1 => n3680, A2 => n7541, ZN => n3679);
   U4849 : XNOR2_X1 port map( A => n8796, B => n8795, ZN => n9137);
   U4850 : XNOR2_X1 port map( A => n9007, B => n2560, ZN => n9115);
   U4851 : INV_X1 port map( A => n7553, ZN => n2323);
   U4852 : OAI22_X1 port map( A1 => n7043, A2 => n3730, B1 => n9355, B2 => 
                           n7044, ZN => n4481);
   U4854 : OR2_X1 port map( A1 => n7073, A2 => n437, ZN => n3814);
   U4855 : XNOR2_X1 port map( A => n4802, B => n8691, ZN => n8994);
   U4856 : OR2_X1 port map( A1 => n7909, A2 => n7364, ZN => n4825);
   U4857 : XNOR2_X1 port map( A => n8237, B => n3715, ZN => n4913);
   U4858 : XNOR2_X1 port map( A => n4378, B => n8639, ZN => n9111);
   U4859 : INV_X1 port map( A => n10186, ZN => n9520);
   U4860 : OAI21_X1 port map( B1 => n9717, B2 => n9716, A => n9715, ZN => 
                           n10533);
   U4861 : AND2_X1 port map( A1 => n9713, A2 => n10037, ZN => n1669);
   U4863 : INV_X1 port map( A => n9702, ZN => n4656);
   U4864 : AND2_X1 port map( A1 => n3762, A2 => n10571, ZN => n3758);
   U4865 : AND2_X1 port map( A1 => n10942, A2 => n5392, ZN => n3761);
   U4866 : INV_X1 port map( A => n9355, ZN => n3730);
   U4867 : AND2_X1 port map( A1 => n10848, A2 => n10850, ZN => n5077);
   U4868 : INV_X1 port map( A => n11121, ZN => n10460);
   U4869 : AND2_X1 port map( A1 => n10682, A2 => n11004, ZN => n11006);
   U4870 : AND2_X1 port map( A1 => n9673, A2 => n5279, ZN => n1532);
   U4871 : INV_X1 port map( A => n9795, ZN => n5279);
   U4873 : INV_X1 port map( A => n11190, ZN => n10480);
   U4874 : OAI21_X1 port map( B1 => n1519, B2 => n2294, A => n4993, ZN => n1518
                           );
   U4875 : OAI21_X1 port map( B1 => n9693, B2 => n9876, A => n9692, ZN => n1520
                           );
   U4876 : OR2_X1 port map( A1 => n9664, A2 => n9985, ZN => n2011);
   U4877 : INV_X1 port map( A => n9737, ZN => n9982);
   U4880 : OR2_X1 port map( A1 => n8526, A2 => n9334, ZN => n2046);
   U4881 : AND2_X1 port map( A1 => n9838, A2 => n428, ZN => n9517);
   U4882 : INV_X1 port map( A => n10482, ZN => n10457);
   U4883 : INV_X1 port map( A => n12147, ZN => n12282);
   U4885 : OR2_X1 port map( A1 => n10489, A2 => n10617, ZN => n5062);
   U4887 : OR2_X1 port map( A1 => n2148, A2 => n10985, ZN => n11164);
   U4889 : OR2_X1 port map( A1 => n10283, A2 => n10190, ZN => n2226);
   U4890 : AND2_X1 port map( A1 => n5393, A2 => n5392, ZN => n5391);
   U4891 : OR2_X1 port map( A1 => n10620, A2 => n233, ZN => n3724);
   U4892 : AND2_X1 port map( A1 => n2849, A2 => n10218, ZN => n10219);
   U4893 : XNOR2_X1 port map( A => n2917, B => n12023, ZN => n12181);
   U4894 : AND2_X1 port map( A1 => n11122, A2 => n10722, ZN => n10723);
   U4895 : OR2_X1 port map( A1 => n10936, A2 => n10935, ZN => n2307);
   U4896 : OR2_X1 port map( A1 => n5296, A2 => n2311, ZN => n2310);
   U4897 : OR2_X1 port map( A1 => n10549, A2 => n10699, ZN => n4758);
   U4899 : OR2_X1 port map( A1 => n2584, A2 => n10596, ZN => n10600);
   U4900 : OR2_X1 port map( A1 => n301, A2 => n2295, ZN => n5312);
   U4901 : XNOR2_X1 port map( A => n11567, B => n11566, ZN => n12520);
   U4902 : INV_X1 port map( A => n12396, ZN => n3269);
   U4903 : OR2_X1 port map( A1 => n3573, A2 => n11069, ZN => n10348);
   U4904 : INV_X1 port map( A => n11295, ZN => n3448);
   U4905 : XNOR2_X1 port map( A => n11385, B => n11653, ZN => n11848);
   U4906 : NAND2_X1 port map( A1 => n10659, A2 => n10660, ZN => n2450);
   U4907 : INV_X1 port map( A => n12167, ZN => n11486);
   U4908 : XNOR2_X1 port map( A => n12381, B => n12048, ZN => n11812);
   U4909 : OR2_X1 port map( A1 => n11050, A2 => n11051, ZN => n3144);
   U4910 : INV_X1 port map( A => n11787, ZN => n12081);
   U4911 : OR2_X1 port map( A1 => n10293, A2 => n11129, ZN => n10295);
   U4912 : XNOR2_X1 port map( A => n4670, B => n23476, ZN => n11225);
   U4913 : AND2_X1 port map( A1 => n14141, A2 => n14143, ZN => n2178);
   U4914 : INV_X1 port map( A => n403, ZN => n3974);
   U4915 : AOI21_X1 port map( B1 => n13178, B2 => n24499, A => n3968, ZN => 
                           n3975);
   U4916 : OR2_X1 port map( A1 => n12469, A2 => n12470, ZN => n4336);
   U4917 : INV_X1 port map( A => n12470, ZN => n13066);
   U4918 : OR2_X1 port map( A1 => n13234, A2 => n13298, ZN => n2544);
   U4919 : AND2_X1 port map( A1 => n14124, A2 => n14208, ZN => n13813);
   U4920 : INV_X1 port map( A => n13843, ZN => n14067);
   U4921 : OR2_X1 port map( A1 => n14294, A2 => n13907, ZN => n11369);
   U4922 : OR2_X1 port map( A1 => n13568, A2 => n13569, ZN => n2603);
   U4923 : NOR2_X1 port map( A1 => n14017, A2 => n2573, ZN => n14020);
   U4924 : AND2_X1 port map( A1 => n14089, A2 => n13533, ZN => n2573);
   U4925 : INV_X1 port map( A => n13901, ZN => n13959);
   U4927 : INV_X1 port map( A => n14301, ZN => n3966);
   U4928 : OAI211_X1 port map( C1 => n13591, C2 => n13864, A => n2417, B => 
                           n5150, ZN => n14698);
   U4929 : OR2_X1 port map( A1 => n12803, A2 => n298, ZN => n2417);
   U4931 : AND2_X1 port map( A1 => n14321, A2 => n3401, ZN => n13500);
   U4932 : XNOR2_X1 port map( A => n15005, B => n1907, ZN => n13524);
   U4933 : INV_X1 port map( A => n15476, ZN => n1907);
   U4934 : OR2_X1 port map( A1 => n13807, A2 => n3717, ZN => n13515);
   U4935 : OR2_X1 port map( A1 => n4452, A2 => n14165, ZN => n4451);
   U4936 : OAI211_X1 port map( C1 => n4763, C2 => n14166, A => n14170, B => 
                           n4762, ZN => n14697);
   U4937 : OR2_X1 port map( A1 => n14171, A2 => n14172, ZN => n4762);
   U4938 : AND2_X1 port map( A1 => n14268, A2 => n14269, ZN => n12542);
   U4939 : OR2_X1 port map( A1 => n14226, A2 => n14225, ZN => n1747);
   U4941 : NOR2_X1 port map( A1 => n14000, A2 => n12669, ZN => n14004);
   U4943 : AND2_X1 port map( A1 => n14102, A2 => n14216, ZN => n4876);
   U4944 : INV_X1 port map( A => n14102, ZN => n4877);
   U4945 : AND2_X1 port map( A1 => n2570, A2 => n3888, ZN => n14202);
   U4946 : OR2_X1 port map( A1 => n3338, A2 => n12639, ZN => n4765);
   U4947 : OR2_X1 port map( A1 => n13701, A2 => n13923, ZN => n13707);
   U4948 : AND2_X1 port map( A1 => n13995, A2 => n25435, ZN => n14236);
   U4949 : OAI21_X1 port map( B1 => n3808, B2 => n3807, A => n13712, ZN => 
                           n11681);
   U4952 : INV_X1 port map( A => n2242, ZN => n3233);
   U4954 : OR2_X1 port map( A1 => n14334, A2 => n14336, ZN => n3059);
   U4955 : XNOR2_X1 port map( A => n13906, B => n5251, ZN => n15411);
   U4956 : INV_X1 port map( A => n14940, ZN => n4557);
   U4957 : OAI21_X1 port map( B1 => n24152, B2 => n14306, A => n12120, ZN => 
                           n12176);
   U4958 : NAND2_X1 port map( A1 => n13525, A2 => n13864, ZN => n2507);
   U4959 : AND2_X1 port map( A1 => n3777, A2 => n3776, ZN => n14437);
   U4960 : XNOR2_X1 port map( A => n15111, B => n15112, ZN => n15114);
   U4961 : AND2_X1 port map( A1 => n4382, A2 => n4383, ZN => n13263);
   U4963 : OR2_X1 port map( A1 => n4016, A2 => n2457, ZN => n4015);
   U4964 : XNOR2_X1 port map( A => n4637, B => n4635, ZN => n4897);
   U4965 : INV_X1 port map( A => n2375, ZN => n16050);
   U4966 : INV_X1 port map( A => n14915, ZN => n4095);
   U4967 : NOR2_X1 port map( A1 => n11806, A2 => n13966, ZN => n13470);
   U4968 : OR2_X1 port map( A1 => n13968, A2 => n13969, ZN => n3802);
   U4969 : OR2_X1 port map( A1 => n4019, A2 => n14219, ZN => n13831);
   U4970 : AOI21_X1 port map( B1 => n2170, B2 => n2172, A => n1868, ZN => n1867
                           );
   U4971 : OAI211_X1 port map( C1 => n14107, C2 => n14112, A => n14109, B => 
                           n13582, ZN => n3983);
   U4972 : XNOR2_X1 port map( A => n15071, B => n14594, ZN => n14389);
   U4973 : OR2_X1 port map( A1 => n14144, A2 => n3887, ZN => n3678);
   U4974 : XNOR2_X1 port map( A => n14902, B => n14936, ZN => n4966);
   U4975 : OAI21_X1 port map( B1 => n3756, B2 => n13843, A => n300, ZN => n3755
                           );
   U4976 : AOI22_X1 port map( A1 => n13597, A2 => n13966, B1 => n11806, B2 => 
                           n13969, ZN => n13598);
   U4977 : OAI211_X1 port map( C1 => n14123, C2 => n13814, A => n13548, B => 
                           n14122, ZN => n2382);
   U4978 : XNOR2_X1 port map( A => n15062, B => n15133, ZN => n15462);
   U4979 : XNOR2_X1 port map( A => n15119, B => n14775, ZN => n15461);
   U4980 : AOI21_X1 port map( B1 => n13477, B2 => n14141, A => n14140, ZN => 
                           n5297);
   U4981 : INV_X1 port map( A => n14141, ZN => n5299);
   U4982 : INV_X1 port map( A => n16095, ZN => n1762);
   U4984 : XNOR2_X1 port map( A => n13441, B => n4582, ZN => n4581);
   U4985 : OR2_X1 port map( A1 => n16410, A2 => n16414, ZN => n3061);
   U4986 : OR2_X1 port map( A1 => n15583, A2 => n16100, ZN => n5245);
   U4987 : AND2_X1 port map( A1 => n17275, A2 => n17273, ZN => n2511);
   U4989 : OR2_X1 port map( A1 => n16225, A2 => n24506, ZN => n5383);
   U4990 : OR2_X1 port map( A1 => n2587, A2 => n16796, ZN => n5243);
   U4991 : AND2_X1 port map( A1 => n15953, A2 => n16480, ZN => n4773);
   U4993 : AND2_X1 port map( A1 => n17326, A2 => n17265, ZN => n17266);
   U4994 : OR2_X1 port map( A1 => n16324, A2 => n16323, ZN => n15899);
   U4995 : INV_X1 port map( A => n17015, ZN => n17214);
   U4996 : OR2_X1 port map( A1 => n17324, A2 => n17326, ZN => n3991);
   U4997 : INV_X1 port map( A => n16892, ZN => n16893);
   U5000 : INV_X1 port map( A => n15612, ZN => n15856);
   U5001 : INV_X1 port map( A => n15611, ZN => n16117);
   U5002 : OR2_X1 port map( A1 => n16118, A2 => n15804, ZN => n2518);
   U5003 : AND2_X1 port map( A1 => n17435, A2 => n17434, ZN => n16429);
   U5004 : AND2_X1 port map( A1 => n17421, A2 => n17381, ZN => n17426);
   U5005 : OR2_X1 port map( A1 => n17185, A2 => n25465, ZN => n17025);
   U5006 : OR2_X1 port map( A1 => n17123, A2 => n4664, ZN => n4663);
   U5007 : INV_X1 port map( A => n1896, ZN => n4664);
   U5009 : NOR2_X1 port map( A1 => n17282, A2 => n17254, ZN => n4941);
   U5010 : INV_X1 port map( A => n5018, ZN => n16662);
   U5012 : OR2_X1 port map( A1 => n3955, A2 => n370, ZN => n3953);
   U5013 : NAND3_X1 port map( A1 => n2265, A2 => n16953, A3 => n2264, ZN => 
                           n17791);
   U5014 : INV_X1 port map( A => n17532, ZN => n18293);
   U5015 : AND2_X1 port map( A1 => n17618, A2 => n17617, ZN => n18018);
   U5016 : OR2_X1 port map( A1 => n17457, A2 => n5073, ZN => n17459);
   U5017 : XNOR2_X1 port map( A => n17724, B => n17725, ZN => n18812);
   U5018 : OAI21_X1 port map( B1 => n3602, B2 => n17391, A => n17388, ZN => 
                           n3601);
   U5019 : NOR2_X1 port map( A1 => n17186, A2 => n3317, ZN => n3603);
   U5020 : XNOR2_X1 port map( A => n24888, B => n18275, ZN => n18475);
   U5021 : INV_X1 port map( A => n19445, ZN => n19449);
   U5022 : OR2_X1 port map( A1 => n16740, A2 => n17084, ZN => n4614);
   U5024 : OR2_X1 port map( A1 => n16557, A2 => n17211, ZN => n16259);
   U5026 : XNOR2_X1 port map( A => n17709, B => n18466, ZN => n17882);
   U5027 : AND2_X1 port map( A1 => n17312, A2 => n17305, ZN => n3626);
   U5028 : INV_X1 port map( A => n18812, ZN => n19390);
   U5029 : AND2_X1 port map( A1 => n17524, A2 => n17171, ZN => n16823);
   U5030 : XNOR2_X1 port map( A => n3706, B => n18660, ZN => n2692);
   U5031 : AND2_X1 port map( A1 => n17575, A2 => n17574, ZN => n1637);
   U5032 : AOI21_X1 port map( B1 => n1640, B2 => n1639, A => n17574, ZN => 
                           n1638);
   U5033 : XNOR2_X1 port map( A => n17970, B => n17811, ZN => n18463);
   U5035 : INV_X1 port map( A => n18128, ZN => n18371);
   U5037 : INV_X1 port map( A => n18448, ZN => n3197);
   U5038 : OR2_X1 port map( A1 => n19088, A2 => n19419, ZN => n19089);
   U5039 : OR2_X1 port map( A1 => n16630, A2 => n16629, ZN => n16631);
   U5040 : XNOR2_X1 port map( A => n18257, B => n18256, ZN => n19278);
   U5041 : INV_X1 port map( A => n19470, ZN => n3748);
   U5042 : XNOR2_X1 port map( A => n2283, B => n18388, ZN => n18458);
   U5043 : OR2_X1 port map( A1 => n16734, A2 => n17067, ZN => n5674);
   U5044 : XNOR2_X1 port map( A => n18227, B => n18293, ZN => n17679);
   U5045 : XNOR2_X1 port map( A => n17112, B => n17113, ZN => n17496);
   U5046 : OR2_X1 port map( A1 => n16845, A2 => n2064, ZN => n5136);
   U5047 : XNOR2_X1 port map( A => n18559, B => n23151, ZN => n2334);
   U5048 : XNOR2_X1 port map( A => n17673, B => n2332, ZN => n19488);
   U5049 : INV_X1 port map( A => n20386, ZN => n19345);
   U5051 : NOR2_X1 port map( A1 => n19361, A2 => n19210, ZN => n4853);
   U5052 : OR2_X1 port map( A1 => n18998, A2 => n19420, ZN => n19088);
   U5053 : OAI21_X1 port map( B1 => n19426, B2 => n19760, A => n2663, ZN => 
                           n19761);
   U5054 : INV_X1 port map( A => n19302, ZN => n18766);
   U5055 : AND2_X1 port map( A1 => n19413, A2 => n19408, ZN => n1890);
   U5056 : AND2_X1 port map( A1 => n2216, A2 => n19376, ZN => n2410);
   U5057 : BUF_X1 port map( A => n19021, Z => n17762);
   U5058 : OR2_X1 port map( A1 => n19460, A2 => n18976, ZN => n18978);
   U5059 : OR2_X1 port map( A1 => n20536, A2 => n20145, ZN => n20146);
   U5060 : OR2_X1 port map( A1 => n18851, A2 => n19479, ZN => n4403);
   U5061 : OR2_X1 port map( A1 => n17554, A2 => n19272, ZN => n4916);
   U5062 : OR2_X1 port map( A1 => n19539, A2 => n3773, ZN => n3751);
   U5063 : OR2_X1 port map( A1 => n19520, A2 => n19522, ZN => n18206);
   U5064 : AND2_X1 port map( A1 => n19568, A2 => n19570, ZN => n3995);
   U5065 : OAI21_X1 port map( B1 => n19570, B2 => n19191, A => n19192, ZN => 
                           n3996);
   U5066 : OAI21_X1 port map( B1 => n19106, B2 => n19105, A => n2464, ZN => 
                           n2462);
   U5067 : INV_X1 port map( A => n19799, ZN => n1522);
   U5068 : INV_X1 port map( A => n19128, ZN => n18767);
   U5069 : INV_X1 port map( A => n18790, ZN => n19400);
   U5070 : INV_X1 port map( A => n19522, ZN => n18895);
   U5072 : INV_X1 port map( A => n19304, ZN => n18947);
   U5074 : AND2_X1 port map( A1 => n19531, A2 => n24329, ZN => n19535);
   U5075 : AND2_X1 port map( A1 => n19579, A2 => n19580, ZN => n2069);
   U5076 : XNOR2_X1 port map( A => n18066, B => n18065, ZN => n19077);
   U5077 : INV_X1 port map( A => n19311, ZN => n5371);
   U5078 : XNOR2_X1 port map( A => n17008, B => n17007, ZN => n19312);
   U5079 : XNOR2_X1 port map( A => n5302, B => n5305, ZN => n5301);
   U5080 : XNOR2_X1 port map( A => n17033, B => n3534, ZN => n17034);
   U5081 : AND2_X1 port map( A1 => n20598, A2 => n20599, ZN => n19740);
   U5082 : OR2_X1 port map( A1 => n25223, A2 => n20215, ZN => n2606);
   U5083 : XNOR2_X1 port map( A => n2569, B => n25222, ZN => n21494);
   U5084 : XNOR2_X1 port map( A => n21501, B => n21500, ZN => n21502);
   U5085 : INV_X1 port map( A => n20533, ZN => n20539);
   U5088 : INV_X1 port map( A => n18729, ZN => n19228);
   U5089 : AND2_X1 port map( A1 => n20111, A2 => n20109, ZN => n3326);
   U5091 : AND2_X1 port map( A1 => n19658, A2 => n3240, ZN => n3241);
   U5093 : OR2_X1 port map( A1 => n18783, A2 => n19407, ZN => n5670);
   U5094 : OR2_X1 port map( A1 => n20016, A2 => n20137, ZN => n19994);
   U5095 : INV_X1 port map( A => n19917, ZN => n20117);
   U5096 : AND2_X1 port map( A1 => n18994, A2 => n20319, ZN => n19691);
   U5098 : OR2_X1 port map( A1 => n5189, A2 => n2024, ZN => n5185);
   U5099 : AND2_X1 port map( A1 => n20960, A2 => n20451, ZN => n1614);
   U5100 : XNOR2_X1 port map( A => n21573, B => n21721, ZN => n21217);
   U5101 : OAI21_X1 port map( B1 => n22465, B2 => n22462, A => n22464, ZN => 
                           n3906);
   U5102 : INV_X1 port map( A => n24042, ZN => n2679);
   U5103 : OR2_X1 port map( A1 => n20446, A2 => n20447, ZN => n3075);
   U5105 : OR2_X1 port map( A1 => n22421, A2 => n2674, ZN => n2671);
   U5106 : OR2_X1 port map( A1 => n22887, A2 => n22728, ZN => n3836);
   U5107 : XNOR2_X1 port map( A => n21608, B => n20826, ZN => n20881);
   U5108 : OR2_X1 port map( A1 => n22241, A2 => n22242, ZN => n2753);
   U5109 : AOI21_X2 port map( B1 => n2356, B2 => n19156, A => n2358, ZN => 
                           n21266);
   U5110 : INV_X1 port map( A => n20697, ZN => n21325);
   U5111 : NOR2_X1 port map( A1 => n22656, A2 => n25241, ZN => n3741);
   U5112 : INV_X1 port map( A => n1605, ZN => n2393);
   U5113 : NOR2_X1 port map( A1 => n22592, A2 => n1605, ZN => n22590);
   U5114 : AND2_X1 port map( A1 => n25066, A2 => n2393, ZN => n21188);
   U5116 : OAI21_X1 port map( B1 => n2828, B2 => n21368, A => n5539, ZN => 
                           n22511);
   U5117 : AND2_X1 port map( A1 => n25471, A2 => n22590, ZN => n22318);
   U5118 : OR2_X1 port map( A1 => n24971, A2 => n1593, ZN => n21936);
   U5119 : NOR2_X1 port map( A1 => n21883, A2 => n22401, ZN => n22263);
   U5120 : AND2_X1 port map( A1 => n22335, A2 => n22338, ZN => n4442);
   U5121 : AND2_X1 port map( A1 => n22268, A2 => n22396, ZN => n3781);
   U5122 : NOR2_X1 port map( A1 => n4098, A2 => n22975, ZN => n4372);
   U5124 : NOR2_X1 port map( A1 => n22198, A2 => n23574, ZN => n23573);
   U5125 : OR2_X1 port map( A1 => n22166, A2 => n22072, ZN => n1679);
   U5126 : AND2_X1 port map( A1 => n22911, A2 => n23464, ZN => n2691);
   U5127 : INV_X1 port map( A => n22072, ZN => n4064);
   U5128 : OR2_X1 port map( A1 => n22092, A2 => n22156, ZN => n22067);
   U5129 : XNOR2_X1 port map( A => n20835, B => n20834, ZN => n23575);
   U5132 : INV_X1 port map( A => n21903, ZN => n2477);
   U5133 : OR2_X1 port map( A1 => n24895, A2 => n23002, ZN => n21902);
   U5134 : INV_X1 port map( A => n24895, ZN => n4533);
   U5135 : OAI21_X1 port map( B1 => n4473, B2 => n22812, A => n4471, ZN => 
                           n22826);
   U5136 : OR2_X1 port map( A1 => n22658, A2 => n4469, ZN => n4471);
   U5137 : OR2_X1 port map( A1 => n23480, A2 => n23481, ZN => n2539);
   U5138 : OR2_X1 port map( A1 => n23053, A2 => n23048, ZN => n3909);
   U5139 : NAND2_X1 port map( A1 => n23042, A2 => n3913, ZN => n3912);
   U5140 : AND2_X1 port map( A1 => n23049, A2 => n23048, ZN => n3913);
   U5141 : OR2_X1 port map( A1 => n21930, A2 => n22464, ZN => n21931);
   U5142 : AND2_X1 port map( A1 => n5084, A2 => n22400, ZN => n21915);
   U5143 : INV_X1 port map( A => n4236, ZN => n4233);
   U5144 : INV_X1 port map( A => Key(58), ZN => n4236);
   U5145 : NOR2_X1 port map( A1 => n21924, A2 => n2376, ZN => n21925);
   U5146 : AOI22_X1 port map( A1 => n1440, A2 => n22326, B1 => n21918, B2 => 
                           n5224, ZN => n5223);
   U5147 : OAI22_X1 port map( A1 => n22284, A2 => n2904, B1 => n22563, B2 => 
                           n22285, ZN => n22287);
   U5148 : INV_X1 port map( A => n22563, ZN => n2904);
   U5149 : NOR2_X1 port map( A1 => n25550, A2 => n23277, ZN => n22536);
   U5150 : INV_X1 port map( A => n23317, ZN => n23318);
   U5151 : OAI21_X1 port map( B1 => n22863, B2 => n22862, A => n23462, ZN => 
                           n1799);
   U5152 : OR2_X1 port map( A1 => n22858, A2 => n22857, ZN => n3264);
   U5153 : OAI21_X1 port map( B1 => n23443, B2 => n22527, A => n5348, ZN => 
                           n22529);
   U5154 : OR2_X1 port map( A1 => n23443, A2 => n1370, ZN => n4033);
   U5155 : INV_X1 port map( A => n2710, ZN => n23491);
   U5156 : AOI21_X1 port map( B1 => n2313, B2 => n22206, A => n22209, ZN => 
                           n5226);
   U5157 : AOI21_X1 port map( B1 => n22156, B2 => n22159, A => n22092, ZN => 
                           n5227);
   U5158 : INV_X1 port map( A => n22208, ZN => n2313);
   U5159 : NOR2_X1 port map( A1 => n22058, A2 => n22228, ZN => n4398);
   U5160 : INV_X1 port map( A => n3227, ZN => n3226);
   U5161 : AND2_X1 port map( A1 => n23853, A2 => n24469, ZN => n3737);
   U5162 : OR2_X1 port map( A1 => n3641, A2 => n23998, ZN => n3640);
   U5164 : NOR2_X1 port map( A1 => n22810, A2 => n22813, ZN => n4468);
   U5165 : OR2_X1 port map( A1 => n24012, A2 => n24006, ZN => n3486);
   U5166 : OR2_X1 port map( A1 => n6752, A2 => n6675, ZN => n6753);
   U5167 : OR2_X1 port map( A1 => n6758, A2 => n6757, ZN => n3276);
   U5169 : AND2_X1 port map( A1 => n6776, A2 => n6198, ZN => n4078);
   U5170 : OR2_X1 port map( A1 => n6679, A2 => n6944, ZN => n2843);
   U5171 : INV_X1 port map( A => n4866, ZN => n6335);
   U5172 : OR2_X1 port map( A1 => n6530, A2 => n6531, ZN => n4746);
   U5173 : AOI21_X1 port map( B1 => n6516, B2 => n6515, A => n6514, ZN => n6806
                           );
   U5175 : NOR2_X1 port map( A1 => n7952, A2 => n7423, ZN => n4483);
   U5176 : AND2_X1 port map( A1 => n1698, A2 => n4621, ZN => n2160);
   U5177 : INV_X1 port map( A => n4621, ZN => n6425);
   U5179 : AND2_X1 port map( A1 => n6712, A2 => n24501, ZN => n3445);
   U5180 : OR2_X1 port map( A1 => n7255, A2 => n7600, ZN => n1902);
   U5181 : AND2_X1 port map( A1 => n6682, A2 => n6685, ZN => n4826);
   U5182 : NAND2_X1 port map( A1 => n2279, A2 => n2278, ZN => n7864);
   U5183 : NAND3_X1 port map( A1 => n6293, A2 => n6481, A3 => n6198, ZN => 
                           n2278);
   U5184 : OR2_X1 port map( A1 => n6489, A2 => n6493, ZN => n6781);
   U5185 : INV_X1 port map( A => n7732, ZN => n7640);
   U5186 : OR2_X1 port map( A1 => n4621, A2 => n6470, ZN => n6203);
   U5187 : OAI21_X1 port map( B1 => n25404, B2 => n1698, A => n5966, ZN => 
                           n1696);
   U5188 : AOI21_X1 port map( B1 => n2351, B2 => n2350, A => n5964, ZN => n7461
                           );
   U5189 : INV_X1 port map( A => n2352, ZN => n2351);
   U5190 : OR2_X1 port map( A1 => n6692, A2 => n6977, ZN => n4828);
   U5191 : AND2_X1 port map( A1 => n7532, A2 => n5738, ZN => n2196);
   U5192 : INV_X1 port map( A => n2534, ZN => n7100);
   U5193 : OAI211_X1 port map( C1 => n7103, C2 => n6539, A => n2532, B => n6543
                           , ZN => n7104);
   U5195 : OR2_X1 port map( A1 => n7975, A2 => n7976, ZN => n7517);
   U5197 : INV_X1 port map( A => n7234, ZN => n7682);
   U5198 : AND2_X1 port map( A1 => n6733, A2 => n6395, ZN => n2900);
   U5200 : INV_X1 port map( A => n7525, ZN => n1677);
   U5201 : OR2_X1 port map( A1 => n7768, A2 => n7526, ZN => n4247);
   U5202 : AND2_X1 port map( A1 => n5574, A2 => n3444, ZN => n1641);
   U5203 : INV_X1 port map( A => n1558, ZN => n1559);
   U5204 : OR2_X1 port map( A1 => n25253, A2 => n7449, ZN => n7636);
   U5206 : AND2_X1 port map( A1 => n6301, A2 => n6784, ZN => n1561);
   U5207 : INV_X1 port map( A => n9066, ZN => n7427);
   U5208 : NOR2_X1 port map( A1 => n7217, A2 => n8316, ZN => n7698);
   U5209 : INV_X1 port map( A => n7595, ZN => n7135);
   U5210 : OR2_X1 port map( A1 => n6805, A2 => n8527, ZN => n6549);
   U5212 : INV_X1 port map( A => n7860, ZN => n4537);
   U5214 : OR2_X1 port map( A1 => n6403, A2 => n6752, ZN => n1735);
   U5215 : OR2_X1 port map( A1 => n6630, A2 => n6407, ZN => n6412);
   U5216 : INV_X1 port map( A => n7474, ZN => n5413);
   U5217 : INV_X1 port map( A => n7615, ZN => n7385);
   U5218 : OR2_X1 port map( A1 => n7896, A2 => n3469, ZN => n2846);
   U5220 : INV_X1 port map( A => n8457, ZN => n8764);
   U5221 : INV_X1 port map( A => n4400, ZN => n7971);
   U5222 : INV_X1 port map( A => n7349, ZN => n8508);
   U5223 : AND2_X1 port map( A1 => n4259, A2 => n7657, ZN => n7228);
   U5224 : AND2_X1 port map( A1 => n5651, A2 => n6772, ZN => n2836);
   U5225 : AND2_X1 port map( A1 => n6312, A2 => n6311, ZN => n3608);
   U5226 : AND2_X1 port map( A1 => n7862, A2 => n7864, ZN => n7553);
   U5227 : INV_X1 port map( A => n8005, ZN => n7543);
   U5228 : AOI21_X1 port map( B1 => n6171, B2 => n6170, A => n6350, ZN => n5068
                           );
   U5229 : AND2_X1 port map( A1 => n6191, A2 => n7761, ZN => n7391);
   U5230 : INV_X1 port map( A => n5202, ZN => n3268);
   U5231 : NOR2_X1 port map( A1 => n8005, A2 => n7292, ZN => n2520);
   U5232 : OR2_X1 port map( A1 => n9066, A2 => n9067, ZN => n7428);
   U5233 : NOR2_X1 port map( A1 => n7588, A2 => n7335, ZN => n7338);
   U5234 : INV_X1 port map( A => n7943, ZN => n6931);
   U5235 : OR2_X1 port map( A1 => n7489, A2 => n7943, ZN => n6929);
   U5236 : INV_X1 port map( A => n8316, ZN => n8314);
   U5237 : INV_X1 port map( A => n7255, ZN => n7598);
   U5238 : INV_X1 port map( A => n7537, ZN => n8013);
   U5239 : OR2_X1 port map( A1 => n6582, A2 => n6755, ZN => n5604);
   U5240 : INV_X1 port map( A => n5607, ZN => n5460);
   U5241 : OR2_X1 port map( A1 => n6243, A2 => n6114, ZN => n6720);
   U5242 : OR2_X1 port map( A1 => n6824, A2 => n6829, ZN => n4122);
   U5243 : AND2_X1 port map( A1 => n7475, A2 => n7474, ZN => n7221);
   U5244 : INV_X1 port map( A => n1345, ZN => n3488);
   U5245 : OR2_X1 port map( A1 => n7961, A2 => n7683, ZN => n7485);
   U5246 : OR2_X1 port map( A1 => n7942, A2 => n4672, ZN => n3677);
   U5247 : AND2_X1 port map( A1 => n7861, A2 => n7707, ZN => n7271);
   U5248 : INV_X1 port map( A => n7861, ZN => n7868);
   U5250 : NAND2_X1 port map( A1 => n1839, A2 => n7462, ZN => n5552);
   U5251 : AND2_X1 port map( A1 => n268, A2 => n5970, ZN => n5549);
   U5252 : OR2_X1 port map( A1 => n7908, A2 => n7364, ZN => n5390);
   U5254 : AND2_X1 port map( A1 => n25252, A2 => n7768, ZN => n7525);
   U5255 : INV_X1 port map( A => n7322, ZN => n7891);
   U5256 : OR2_X1 port map( A1 => n4839, A2 => n442, ZN => n3142);
   U5257 : INV_X1 port map( A => n7578, ZN => n7576);
   U5259 : AND2_X1 port map( A1 => n7141, A2 => n7902, ZN => n2780);
   U5260 : NAND3_X1 port map( A1 => n5265, A2 => n5268, A3 => n5263, ZN => 
                           n8477);
   U5261 : AND2_X1 port map( A1 => n7734, A2 => n7642, ZN => n7730);
   U5262 : OR2_X1 port map( A1 => n6950, A2 => n25437, ZN => n4757);
   U5263 : AOI21_X1 port map( B1 => n3923, B2 => n6553, A => n3922, ZN => n3921
                           );
   U5264 : OR2_X1 port map( A1 => n6137, A2 => n6705, ZN => n3924);
   U5265 : OR2_X1 port map( A1 => n440, A2 => n6524, ZN => n6154);
   U5266 : OR2_X1 port map( A1 => n6963, A2 => n6570, ZN => n6571);
   U5267 : OR2_X1 port map( A1 => n6688, A2 => n6686, ZN => n6567);
   U5268 : OR2_X1 port map( A1 => n1985, A2 => n7965, ZN => n7236);
   U5269 : OR2_X1 port map( A1 => n7070, A2 => n7962, ZN => n1984);
   U5270 : AND2_X1 port map( A1 => n5713, A2 => n7433, ZN => n2858);
   U5271 : OR2_X1 port map( A1 => n7175, A2 => n7782, ZN => n7176);
   U5272 : AOI21_X1 port map( B1 => n4705, B2 => n3344, A => n3587, ZN => n4710
                           );
   U5274 : OR2_X1 port map( A1 => n3979, A2 => n8367, ZN => n7558);
   U5275 : INV_X1 port map( A => n8616, ZN => n8400);
   U5276 : AND2_X1 port map( A1 => n7740, A2 => n7811, ZN => n4803);
   U5277 : OR2_X1 port map( A1 => n9469, A2 => n1595, ZN => n1594);
   U5278 : INV_X1 port map( A => n9959, ZN => n2876);
   U5279 : AND2_X2 port map( A1 => n2275, A2 => n4785, ZN => n8721);
   U5280 : OR2_X1 port map( A1 => n4784, A2 => n7661, ZN => n2275);
   U5281 : XNOR2_X1 port map( A => n8806, B => n8492, ZN => n8714);
   U5282 : OR2_X1 port map( A1 => n7345, A2 => n7600, ZN => n1999);
   U5283 : INV_X1 port map( A => n8501, ZN => n8973);
   U5284 : INV_X1 port map( A => n2058, ZN => n5328);
   U5285 : INV_X1 port map( A => n8798, ZN => n5343);
   U5286 : XNOR2_X1 port map( A => n2560, B => n8923, ZN => n7083);
   U5287 : XNOR2_X1 port map( A => n8416, B => n8415, ZN => n10157);
   U5288 : AND2_X1 port map( A1 => n9843, A2 => n10149, ZN => n9844);
   U5289 : INV_X1 port map( A => n9211, ZN => n7437);
   U5291 : INV_X1 port map( A => n25232, ZN => n5621);
   U5292 : AND2_X1 port map( A1 => n10951, A2 => n25074, ZN => n5106);
   U5293 : INV_X1 port map( A => n10703, ZN => n5107);
   U5294 : AND2_X1 port map( A1 => n9435, A2 => n9635, ZN => n1939);
   U5295 : XNOR2_X1 port map( A => n8130, B => n8129, ZN => n9944);
   U5296 : AND2_X1 port map( A1 => n24083, A2 => n9899, ZN => n9289);
   U5297 : OR2_X1 port map( A1 => n10168, A2 => n10166, ZN => n2091);
   U5298 : INV_X1 port map( A => n10811, ZN => n5628);
   U5299 : INV_X1 port map( A => n10314, ZN => n10165);
   U5300 : AND2_X1 port map( A1 => n11215, A2 => n10669, ZN => n5085);
   U5301 : AND2_X1 port map( A1 => n10942, A2 => n11039, ZN => n2870);
   U5302 : AND2_X1 port map( A1 => n9872, A2 => n2294, ZN => n2293);
   U5303 : AOI21_X1 port map( B1 => n9883, B2 => n25069, A => n9563, ZN => 
                           n5066);
   U5305 : INV_X1 port map( A => n11046, ZN => n10641);
   U5306 : INV_X1 port map( A => n10757, ZN => n2867);
   U5307 : NAND2_X1 port map( A1 => n9342, A2 => n1464, ZN => n1658);
   U5308 : OR2_X1 port map( A1 => n9668, A2 => n9999, ZN => n9311);
   U5309 : OR2_X1 port map( A1 => n10054, A2 => n10052, ZN => n1871);
   U5311 : AND2_X1 port map( A1 => n10989, A2 => n10406, ZN => n10996);
   U5312 : OR2_X1 port map( A1 => n25229, A2 => n10737, ZN => n10283);
   U5313 : INV_X1 port map( A => n10858, ZN => n10859);
   U5314 : NOR2_X1 port map( A1 => n8178, A2 => n8179, ZN => n10994);
   U5315 : AND2_X1 port map( A1 => n10406, A2 => n10990, ZN => n8146);
   U5316 : OR2_X1 port map( A1 => n3467, A2 => n11101, ZN => n2849);
   U5317 : INV_X1 port map( A => n10891, ZN => n2185);
   U5318 : OR3_X1 port map( A1 => n10830, A2 => n10831, A3 => n10836, ZN => 
                           n4778);
   U5319 : OR2_X1 port map( A1 => n25217, A2 => n9603, ZN => n2928);
   U5320 : INV_X1 port map( A => n12261, ZN => n12218);
   U5321 : NOR2_X1 port map( A1 => n4251, A2 => n11059, ZN => n4392);
   U5322 : AND2_X1 port map( A1 => n11052, A2 => n11058, ZN => n4391);
   U5323 : INV_X1 port map( A => n10627, ZN => n11563);
   U5324 : OR2_X1 port map( A1 => n10924, A2 => n10993, ZN => n4929);
   U5325 : OR2_X1 port map( A1 => n10185, A2 => n9520, ZN => n5534);
   U5326 : INV_X1 port map( A => n10558, ZN => n10556);
   U5327 : INV_X1 port map( A => n4521, ZN => n9810);
   U5328 : NAND4_X1 port map( A1 => n2152, A2 => n11056, A3 => n3163, A4 => 
                           n1389, ZN => n4759);
   U5329 : INV_X1 port map( A => n10504, ZN => n4671);
   U5330 : INV_X1 port map( A => n10951, ZN => n10955);
   U5331 : INV_X1 port map( A => n11152, ZN => n11147);
   U5332 : AND3_X1 port map( A1 => n10447, A2 => n10448, A3 => n10446, ZN => 
                           n11412);
   U5333 : AOI21_X1 port map( B1 => n11300, B2 => n419, A => n11299, ZN => 
                           n11306);
   U5334 : INV_X1 port map( A => n11146, ZN => n2060);
   U5335 : NOR2_X1 port map( A1 => n25249, A2 => n10714, ZN => n11131);
   U5337 : INV_X1 port map( A => n10398, ZN => n10661);
   U5338 : INV_X1 port map( A => n2243, ZN => n10830);
   U5339 : INV_X1 port map( A => n10941, ZN => n10944);
   U5340 : OAI21_X1 port map( B1 => n9919, B2 => n9355, A => n3967, ZN => n9136
                           );
   U5341 : AND2_X1 port map( A1 => n9135, A2 => n9912, ZN => n2810);
   U5342 : AND2_X1 port map( A1 => n9461, A2 => n9463, ZN => n3967);
   U5343 : INV_X1 port map( A => n11113, ZN => n11110);
   U5345 : INV_X1 port map( A => n12221, ZN => n5180);
   U5346 : INV_X1 port map( A => n11044, ZN => n4532);
   U5347 : INV_X1 port map( A => n11012, ZN => n2681);
   U5348 : NOR2_X1 port map( A1 => n11024, A2 => n8934, ZN => n3771);
   U5349 : AND2_X1 port map( A1 => n10858, A2 => n25230, ZN => n5727);
   U5350 : INV_X1 port map( A => n12134, ZN => n12109);
   U5351 : INV_X1 port map( A => n11628, ZN => n12356);
   U5352 : INV_X1 port map( A => n5340, ZN => n10261);
   U5353 : OAI21_X1 port map( B1 => n10148, B2 => n5357, A => n5355, ZN => 
                           n10867);
   U5354 : INV_X1 port map( A => n1658, ZN => n10875);
   U5356 : INV_X1 port map( A => n5448, ZN => n2498);
   U5357 : OR2_X1 port map( A1 => n11070, A2 => n25203, ZN => n3573);
   U5358 : INV_X1 port map( A => n11412, ZN => n12168);
   U5359 : INV_X1 port map( A => n1499, ZN => n10759);
   U5360 : NOR2_X1 port map( A1 => n10753, A2 => n1499, ZN => n3750);
   U5361 : INV_X1 port map( A => n3324, ZN => n10291);
   U5362 : XNOR2_X1 port map( A => n12261, B => n3158, ZN => n12220);
   U5363 : OR2_X1 port map( A1 => n4937, A2 => n10734, ZN => n2830);
   U5364 : XNOR2_X1 port map( A => n3418, B => n12180, ZN => n12182);
   U5365 : XNOR2_X1 port map( A => n12306, B => n3133, ZN => n3418);
   U5366 : XNOR2_X1 port map( A => n11913, B => n11914, ZN => n2271);
   U5367 : XNOR2_X1 port map( A => n12128, B => n12355, ZN => n3207);
   U5368 : INV_X1 port map( A => n2739, ZN => n4107);
   U5369 : XNOR2_X1 port map( A => n11268, B => n3901, ZN => n12266);
   U5370 : INV_X1 port map( A => n12315, ZN => n5181);
   U5371 : OR2_X1 port map( A1 => n10940, A2 => n24591, ZN => n3252);
   U5372 : XNOR2_X1 port map( A => n25396, B => n5514, ZN => n11571);
   U5373 : INV_X1 port map( A => n11542, ZN => n1699);
   U5374 : INV_X1 port map( A => n4759, ZN => n11706);
   U5376 : NAND2_X1 port map( A1 => n11081, A2 => n4421, ZN => n10222);
   U5377 : OR2_X1 port map( A1 => n10767, A2 => n4422, ZN => n4421);
   U5378 : INV_X1 port map( A => n13153, ZN => n1632);
   U5379 : INV_X1 port map( A => n11424, ZN => n10490);
   U5380 : AND2_X1 port map( A1 => n2628, A2 => n11342, ZN => n10493);
   U5381 : OR2_X1 port map( A1 => n10425, A2 => n10596, ZN => n4211);
   U5382 : INV_X1 port map( A => n1543, ZN => n1538);
   U5383 : INV_X1 port map( A => n1544, ZN => n1537);
   U5385 : INV_X1 port map( A => n11199, ZN => n10229);
   U5386 : XNOR2_X1 port map( A => n11401, B => n2602, ZN => n11665);
   U5388 : AND2_X1 port map( A1 => n24930, A2 => n3688, ZN => n11596);
   U5389 : NOR2_X1 port map( A1 => n414, A2 => n4711, ZN => n11934);
   U5391 : INV_X1 port map( A => n12219, ZN => n5182);
   U5392 : AOI22_X1 port map( A1 => n9241, A2 => n11124, B1 => n10846, B2 => 
                           n305, ZN => n9242);
   U5393 : AND2_X1 port map( A1 => n2680, A2 => n11012, ZN => n10013);
   U5394 : OR2_X1 port map( A1 => n13347, A2 => n12636, ZN => n12858);
   U5395 : AND2_X1 port map( A1 => n13169, A2 => n13167, ZN => n12721);
   U5397 : INV_X1 port map( A => n302, ZN => n1636);
   U5402 : INV_X1 port map( A => n24512, ZN => n13215);
   U5403 : OR2_X1 port map( A1 => n13040, A2 => n12800, ZN => n4639);
   U5405 : OR2_X1 port map( A1 => n12685, A2 => n5311, ZN => n5314);
   U5406 : OR2_X1 port map( A1 => n12684, A2 => n24422, ZN => n5309);
   U5407 : NOR2_X1 port map( A1 => n3689, A2 => n24373, ZN => n13172);
   U5408 : INV_X1 port map( A => n12669, ZN => n3563);
   U5409 : AND2_X1 port map( A1 => n14333, A2 => n14339, ZN => n13878);
   U5410 : OR2_X1 port map( A1 => n13146, A2 => n13145, ZN => n5543);
   U5411 : OR2_X1 port map( A1 => n5412, A2 => n12858, ZN => n3339);
   U5412 : INV_X1 port map( A => n13109, ZN => n4529);
   U5413 : INV_X1 port map( A => n13485, ZN => n14005);
   U5414 : INV_X1 port map( A => n14362, ZN => n3698);
   U5415 : AND2_X1 port map( A1 => n13569, A2 => n13394, ZN => n3808);
   U5416 : NOR2_X1 port map( A1 => n11601, A2 => n11600, ZN => n3807);
   U5417 : AND2_X1 port map( A1 => n13323, A2 => n2295, ZN => n12848);
   U5419 : INV_X1 port map( A => n14107, ZN => n13566);
   U5420 : INV_X1 port map( A => n13265, ZN => n5644);
   U5421 : INV_X1 port map( A => n14129, ZN => n13893);
   U5422 : AND2_X1 port map( A1 => n13868, A2 => n14317, ZN => n3501);
   U5423 : INV_X1 port map( A => n13647, ZN => n13819);
   U5424 : INV_X1 port map( A => n14328, ZN => n2505);
   U5425 : AND2_X1 port map( A1 => n12633, A2 => n4923, ZN => n5471);
   U5426 : OR2_X1 port map( A1 => n13953, A2 => n14158, ZN => n4356);
   U5427 : INV_X1 port map( A => n14211, ZN => n13437);
   U5429 : AOI22_X1 port map( A1 => n12876, A2 => n13357, B1 => n13359, B2 => 
                           n24554, ZN => n2889);
   U5431 : AND2_X1 port map( A1 => n14035, A2 => n14034, ZN => n13806);
   U5433 : OAI21_X1 port map( B1 => n12507, B2 => n12506, A => n3633, ZN => 
                           n3632);
   U5434 : OR2_X1 port map( A1 => n14022, A2 => n13533, ZN => n13609);
   U5435 : AND2_X1 port map( A1 => n12018, A2 => n1527, ZN => n1526);
   U5437 : NOR2_X1 port map( A1 => n14172, A2 => n14165, ZN => n3383);
   U5439 : NOR2_X1 port map( A1 => n14000, A2 => n12668, ZN => n13676);
   U5440 : INV_X1 port map( A => n14165, ZN => n13741);
   U5442 : INV_X1 port map( A => n14190, ZN => n14142);
   U5443 : INV_X1 port map( A => n12536, ZN => n13759);
   U5444 : AND2_X1 port map( A1 => n14274, A2 => n14268, ZN => n13764);
   U5445 : AOI21_X1 port map( B1 => n13733, B2 => n13732, A => n13731, ZN => 
                           n14594);
   U5446 : AND2_X1 port map( A1 => n14106, A2 => n14108, ZN => n1933);
   U5447 : AND3_X1 port map( A1 => n13792, A2 => n13796, A3 => n13578, ZN => 
                           n4331);
   U5448 : OR2_X1 port map( A1 => n14302, A2 => n14301, ZN => n13454);
   U5449 : AND2_X1 port map( A1 => n14153, A2 => n3717, ZN => n3716);
   U5450 : INV_X1 port map( A => n14089, ZN => n14018);
   U5451 : OR2_X1 port map( A1 => n13824, A2 => n13560, ZN => n13389);
   U5453 : INV_X1 port map( A => n13048, ZN => n12489);
   U5454 : INV_X1 port map( A => n4059, ZN => n4058);
   U5456 : OR2_X1 port map( A1 => n12843, A2 => n12946, ZN => n2770);
   U5457 : OR2_X1 port map( A1 => n12844, A2 => n12845, ZN => n2769);
   U5458 : AND2_X1 port map( A1 => n14294, A2 => n14290, ZN => n13722);
   U5459 : NOR2_X1 port map( A1 => n13895, A2 => n4844, ZN => n4043);
   U5460 : AND2_X1 port map( A1 => n399, A2 => n13338, ZN => n12959);
   U5461 : INV_X1 port map( A => n14124, ZN => n14123);
   U5462 : INV_X1 port map( A => n13422, ZN => n2378);
   U5463 : INV_X1 port map( A => n14205, ZN => n2379);
   U5465 : OR2_X1 port map( A1 => n14219, A2 => n14222, ZN => n13022);
   U5466 : OR2_X1 port map( A1 => n13863, A2 => n13864, ZN => n12814);
   U5468 : OAI211_X1 port map( C1 => n5485, C2 => n5487, A => n5483, B => n5482
                           , ZN => n14966);
   U5469 : OAI21_X1 port map( B1 => n15216, B2 => n15215, A => n16641, ZN => 
                           n16945);
   U5473 : OR2_X1 port map( A1 => n16422, A2 => n16427, ZN => n16171);
   U5474 : OAI21_X1 port map( B1 => n13724, B2 => n11806, A => n1771, ZN => 
                           n13727);
   U5475 : AND2_X1 port map( A1 => n14078, A2 => n14077, ZN => n2122);
   U5476 : AND2_X1 port map( A1 => n16443, A2 => n16442, ZN => n2809);
   U5477 : OR2_X1 port map( A1 => n16038, A2 => n16043, ZN => n3578);
   U5478 : XNOR2_X1 port map( A => n14830, B => n1371, ZN => n15564);
   U5479 : INV_X1 port map( A => n14500, ZN => n14806);
   U5480 : OR2_X1 port map( A1 => n386, A2 => n25210, ZN => n4026);
   U5481 : XNOR2_X1 port map( A => n15435, B => n15434, ZN => n15470);
   U5482 : OR2_X1 port map( A1 => n15714, A2 => n16470, ZN => n4972);
   U5483 : INV_X1 port map( A => n24539, ZN => n4927);
   U5484 : OR2_X1 port map( A1 => n15977, A2 => n16394, ZN => n1656);
   U5485 : INV_X1 port map( A => n16225, ZN => n16301);
   U5486 : OR2_X1 port map( A1 => n15686, A2 => n16437, ZN => n2637);
   U5487 : OR2_X1 port map( A1 => n16076, A2 => n14664, ZN => n3636);
   U5488 : INV_X1 port map( A => n16207, ZN => n4914);
   U5490 : AND2_X1 port map( A1 => n17421, A2 => n16945, ZN => n2234);
   U5491 : NOR2_X1 port map( A1 => n2375, A2 => n4897, ZN => n15691);
   U5492 : NOR2_X1 port map( A1 => n16048, A2 => n15605, ZN => n15604);
   U5493 : XNOR2_X1 port map( A => n3471, B => n14962, ZN => n2407);
   U5494 : INV_X1 port map( A => n15953, ZN => n15717);
   U5495 : XNOR2_X1 port map( A => n5009, B => n15352, ZN => n15353);
   U5496 : OR2_X1 port map( A1 => n17085, A2 => n17088, ZN => n3103);
   U5497 : INV_X1 port map( A => n4985, ZN => n4981);
   U5498 : INV_X1 port map( A => n15314, ZN => n17343);
   U5501 : XNOR2_X1 port map( A => n2969, B => n1907, ZN => n14693);
   U5502 : AND2_X1 port map( A1 => n16595, A2 => n24587, ZN => n15824);
   U5503 : AND2_X1 port map( A1 => n5447, A2 => n5667, ZN => n5668);
   U5504 : OAI211_X1 port map( C1 => n5447, C2 => n16001, A => n15758, B => 
                           n3658, ZN => n5666);
   U5505 : OAI21_X1 port map( B1 => n16185, B2 => n15915, A => n5317, ZN => 
                           n1516);
   U5506 : OR2_X1 port map( A1 => n16355, A2 => n16360, ZN => n4496);
   U5507 : OR2_X1 port map( A1 => n16770, A2 => n17039, ZN => n17363);
   U5509 : INV_X1 port map( A => n15937, ZN => n5168);
   U5510 : NOR2_X1 port map( A1 => n15695, A2 => n15953, ZN => n16482);
   U5511 : XNOR2_X1 port map( A => n14262, B => n14263, ZN => n15837);
   U5512 : AND2_X1 port map( A1 => n4046, A2 => n15837, ZN => n15839);
   U5514 : AND2_X1 port map( A1 => n16551, A2 => n5376, ZN => n15739);
   U5516 : OR2_X1 port map( A1 => n14787, A2 => n24163, ZN => n3067);
   U5517 : XNOR2_X1 port map( A => n14822, B => n14821, ZN => n16230);
   U5518 : INV_X1 port map( A => n17320, ZN => n2287);
   U5519 : AND2_X1 port map( A1 => n16769, A2 => n17364, ZN => n2530);
   U5520 : OAI21_X1 port map( B1 => n24586, B2 => n4807, A => n4806, ZN => 
                           n16687);
   U5521 : OR2_X1 port map( A1 => n4353, A2 => n15594, ZN => n4938);
   U5522 : OR2_X1 port map( A1 => n3702, A2 => n16438, ZN => n2202);
   U5523 : AND2_X1 port map( A1 => n16241, A2 => n16437, ZN => n3702);
   U5524 : INV_X1 port map( A => n17212, ZN => n5512);
   U5525 : INV_X1 port map( A => n15470, ZN => n16472);
   U5528 : INV_X1 port map( A => n17728, ZN => n1704);
   U5529 : OR2_X1 port map( A1 => n17690, A2 => n17485, ZN => n1701);
   U5531 : AND2_X1 port map( A1 => n14585, A2 => n1676, ZN => n1675);
   U5532 : INV_X1 port map( A => n17433, ZN => n3000);
   U5533 : AND2_X1 port map( A1 => n17312, A2 => n17316, ZN => n16716);
   U5534 : OR2_X1 port map( A1 => n17596, A2 => n24543, ZN => n4564);
   U5535 : OR2_X1 port map( A1 => n17364, A2 => n25058, ZN => n3951);
   U5536 : OR2_X1 port map( A1 => n16064, A2 => n16067, ZN => n4105);
   U5537 : NOR2_X1 port map( A1 => n25245, A2 => n17132, ZN => n3457);
   U5538 : OR2_X1 port map( A1 => n15668, A2 => n290, ZN => n2286);
   U5539 : OR2_X1 port map( A1 => n17319, A2 => n16607, ZN => n16923);
   U5540 : OAI21_X1 port map( B1 => n13547, B2 => n267, A => n13546, ZN => 
                           n17225);
   U5541 : INV_X1 port map( A => n17225, ZN => n16956);
   U5542 : INV_X1 port map( A => n17387, ZN => n3604);
   U5543 : NAND3_X1 port map( A1 => n382, A2 => n25446, A3 => n15550, ZN => 
                           n5596);
   U5544 : AOI22_X1 port map( A1 => n16828, A2 => n16962, B1 => n1612, B2 => 
                           n24444, ZN => n17128);
   U5545 : OR2_X1 port map( A1 => n15266, A2 => n24429, ZN => n3121);
   U5547 : OAI21_X1 port map( B1 => n15940, B2 => n24163, A => n24162, ZN => 
                           n2344);
   U5548 : INV_X1 port map( A => n16927, ZN => n17322);
   U5549 : INV_X1 port map( A => n16971, ZN => n17332);
   U5550 : OR2_X1 port map( A1 => n25409, A2 => n15584, ZN => n3503);
   U5551 : AND2_X1 port map( A1 => n17316, A2 => n24543, ZN => n3627);
   U5552 : AND2_X1 port map( A1 => n17320, A2 => n16927, ZN => n17267);
   U5553 : AND2_X1 port map( A1 => n17371, A2 => n17042, ZN => n16766);
   U5554 : OR2_X1 port map( A1 => n17414, A2 => n17225, ZN => n5705);
   U5555 : INV_X1 port map( A => n16486, ZN => n16518);
   U5556 : AND2_X1 port map( A1 => n16851, A2 => n17138, ZN => n3930);
   U5557 : AND2_X1 port map( A1 => n17145, A2 => n16984, ZN => n3929);
   U5558 : INV_X1 port map( A => n3778, ZN => n14864);
   U5559 : OR2_X1 port map( A1 => n17608, A2 => n17409, ZN => n16743);
   U5560 : OR2_X1 port map( A1 => n16311, A2 => n16312, ZN => n1817);
   U5561 : OR2_X1 port map( A1 => n16298, A2 => n4957, ZN => n4956);
   U5562 : INV_X1 port map( A => n17131, ZN => n16655);
   U5563 : AND3_X1 port map( A1 => n17081, A2 => n17078, A3 => n17478, ZN => 
                           n2181);
   U5566 : NOR2_X1 port map( A1 => n16353, A2 => n16595, ZN => n3334);
   U5567 : INV_X1 port map( A => n17114, ZN => n4304);
   U5568 : INV_X1 port map( A => n17520, ZN => n18311);
   U5569 : INV_X1 port map( A => n16921, ZN => n17596);
   U5570 : AND2_X1 port map( A1 => n17068, A2 => n16731, ZN => n4286);
   U5571 : INV_X1 port map( A => n16769, ZN => n3685);
   U5572 : NOR2_X1 port map( A1 => n1451, A2 => n1498, ZN => n1497);
   U5573 : AND2_X1 port map( A1 => n15970, A2 => n16186, ZN => n3223);
   U5574 : INV_X1 port map( A => n17624, ZN => n4284);
   U5575 : INV_X1 port map( A => n17622, ZN => n4285);
   U5576 : AND2_X1 port map( A1 => n16112, A2 => n17524, ZN => n17527);
   U5578 : AOI21_X1 port map( B1 => n17314, B2 => n16921, A => n2968, ZN => 
                           n3782);
   U5580 : OR2_X1 port map( A1 => n16440, A2 => n16442, ZN => n15947);
   U5581 : XNOR2_X1 port map( A => n18375, B => n16866, ZN => n16867);
   U5582 : INV_X1 port map( A => n16846, ZN => n16499);
   U5583 : OR2_X1 port map( A1 => n16034, A2 => n15573, ZN => n1927);
   U5584 : INV_X1 port map( A => n17410, ZN => n17609);
   U5585 : INV_X1 port map( A => n16561, ZN => n17407);
   U5586 : OR2_X1 port map( A1 => n16961, A2 => n17445, ZN => n3260);
   U5587 : NAND2_X1 port map( A1 => n15845, A2 => n2992, ZN => n17122);
   U5589 : XNOR2_X1 port map( A => n18157, B => n24886, ZN => n18159);
   U5590 : INV_X1 port map( A => n4114, ZN => n2216);
   U5591 : OR2_X1 port map( A1 => n19312, A2 => n19310, ZN => n18843);
   U5592 : XNOR2_X1 port map( A => n4269, B => n18429, ZN => n4268);
   U5593 : INV_X1 port map( A => n18694, ZN => n4269);
   U5594 : INV_X1 port map( A => n19413, ZN => n3491);
   U5595 : BUF_X1 port map( A => n16910, Z => n17907);
   U5596 : XNOR2_X1 port map( A => n2001, B => n18128, ZN => n18464);
   U5597 : INV_X1 port map( A => n18129, ZN => n2001);
   U5598 : INV_X1 port map( A => n18172, ZN => n4971);
   U5599 : INV_X1 port map( A => n19255, ZN => n18870);
   U5600 : XNOR2_X1 port map( A => n18520, B => n18519, ZN => n19064);
   U5601 : AND2_X1 port map( A1 => n19238, A2 => n18883, ZN => n19067);
   U5602 : AND2_X1 port map( A1 => n19331, A2 => n4291, ZN => n5213);
   U5603 : INV_X1 port map( A => n20586, ZN => n19951);
   U5604 : AND2_X1 port map( A1 => n280, A2 => n19575, ZN => n5155);
   U5606 : INV_X1 port map( A => n19064, ZN => n2298);
   U5607 : AND2_X1 port map( A1 => n19065, A2 => n25012, ZN => n2328);
   U5608 : AND2_X1 port map( A1 => n25012, A2 => n19064, ZN => n19616);
   U5611 : AND2_X1 port map( A1 => n17945, A2 => n4291, ZN => n4288);
   U5612 : OR2_X1 port map( A1 => n19202, A2 => n3412, ZN => n19839);
   U5613 : NAND2_X1 port map( A1 => n276, A2 => n24463, ZN => n5132);
   U5615 : OR2_X1 port map( A1 => n17872, A2 => n18959, ZN => n3583);
   U5616 : AOI21_X1 port map( B1 => n20554, B2 => n20555, A => n2594, ZN => 
                           n20559);
   U5617 : INV_X1 port map( A => n1590, ZN => n2688);
   U5618 : OAI211_X1 port map( C1 => n19080, C2 => n5134, A => n19251, B => 
                           n1501, ZN => n5427);
   U5619 : AOI22_X1 port map( A1 => n19079, A2 => n19592, B1 => n2346, B2 => 
                           n1502, ZN => n1501);
   U5620 : AND2_X1 port map( A1 => n18808, A2 => n19078, ZN => n1502);
   U5621 : OR2_X1 port map( A1 => n19532, A2 => n19272, ZN => n5652);
   U5622 : NAND2_X1 port map( A1 => n4857, A2 => n1505, ZN => n1504);
   U5624 : OR2_X1 port map( A1 => n19009, A2 => n19170, ZN => n3820);
   U5625 : INV_X1 port map( A => n20149, ZN => n20147);
   U5626 : OR2_X1 port map( A1 => n19087, A2 => n24584, ZN => n3668);
   U5627 : INV_X1 port map( A => n5427, ZN => n20497);
   U5628 : AND2_X1 port map( A1 => n20268, A2 => n20501, ZN => n20225);
   U5629 : OAI21_X1 port map( B1 => n18720, B2 => n18721, A => n357, ZN => 
                           n18722);
   U5630 : INV_X1 port map( A => n5475, ZN => n5474);
   U5631 : INV_X1 port map( A => n5569, ZN => n5568);
   U5632 : INV_X1 port map( A => n20576, ZN => n19841);
   U5633 : OR2_X1 port map( A1 => n24583, A2 => n4291, ZN => n4287);
   U5634 : INV_X1 port map( A => n20345, ZN => n1557);
   U5636 : OR2_X1 port map( A1 => n100, A2 => n20507, ZN => n5499);
   U5637 : INV_X1 port map( A => n20614, ZN => n2330);
   U5638 : INV_X1 port map( A => n20617, ZN => n20570);
   U5639 : INV_X1 port map( A => n20616, ZN => n20569);
   U5640 : NOR2_X1 port map( A1 => n5590, A2 => n20414, ZN => n5733);
   U5641 : INV_X1 port map( A => n21533, ZN => n4164);
   U5643 : OAI21_X1 port map( B1 => n18828, B2 => n19002, A => n4195, ZN => 
                           n4194);
   U5644 : OR2_X1 port map( A1 => n19777, A2 => n20173, ZN => n20234);
   U5645 : OR2_X1 port map( A1 => n19255, A2 => n25001, ZN => n3388);
   U5646 : INV_X1 port map( A => n20269, ZN => n20224);
   U5647 : INV_X1 port map( A => n20414, ZN => n5591);
   U5648 : OR2_X1 port map( A1 => n19112, A2 => n2642, ZN => n18867);
   U5649 : OR2_X1 port map( A1 => n19252, A2 => n19078, ZN => n2804);
   U5650 : AND2_X1 port map( A1 => n7, A2 => n20614, ZN => n20572);
   U5652 : INV_X1 port map( A => n20145, ZN => n20447);
   U5653 : OR2_X1 port map( A1 => n20149, A2 => n19018, ZN => n20532);
   U5654 : OR2_X1 port map( A1 => n19168, A2 => n19002, ZN => n2927);
   U5655 : OR2_X1 port map( A1 => n25422, A2 => n19246, ZN => n3987);
   U5656 : INV_X1 port map( A => n20335, ZN => n20666);
   U5657 : OR2_X1 port map( A1 => n20142, A2 => n19979, ZN => n2074);
   U5658 : OR2_X1 port map( A1 => n5007, A2 => n19441, ZN => n2693);
   U5659 : OAI211_X1 port map( C1 => n20114, C2 => n19887, A => n19886, B => 
                           n19885, ZN => n20904);
   U5660 : INV_X1 port map( A => n18978, ZN => n17892);
   U5661 : INV_X1 port map( A => n1591, ZN => n19893);
   U5662 : INV_X1 port map( A => n20518, ZN => n20276);
   U5663 : INV_X1 port map( A => n20437, ZN => n20583);
   U5664 : INV_X1 port map( A => n20193, ZN => n20577);
   U5665 : OR2_X1 port map( A1 => n25205, A2 => n20231, ZN => n19803);
   U5666 : AND2_X1 port map( A1 => n2594, A2 => n20557, ZN => n19880);
   U5667 : AOI21_X1 port map( B1 => n352, B2 => n19345, A => n19344, ZN => 
                           n19348);
   U5668 : INV_X1 port map( A => n19383, ZN => n4008);
   U5669 : OR2_X1 port map( A1 => n19168, A2 => n19421, ZN => n4578);
   U5670 : INV_X1 port map( A => n19423, ZN => n4579);
   U5671 : OR2_X1 port map( A1 => n18818, A2 => n19211, ZN => n4851);
   U5672 : NOR2_X1 port map( A1 => n24275, A2 => n20913, ZN => n20362);
   U5673 : AND2_X1 port map( A1 => n5132, A2 => n5131, ZN => n5130);
   U5674 : INV_X1 port map( A => n20019, ZN => n4728);
   U5675 : INV_X1 port map( A => n19703, ZN => n20623);
   U5676 : INV_X1 port map( A => n19849, ZN => n19852);
   U5677 : INV_X1 port map( A => n19661, ZN => n19657);
   U5678 : NOR2_X1 port map( A1 => n20555, A2 => n20554, ZN => n2369);
   U5679 : INV_X1 port map( A => n20089, ZN => n2370);
   U5680 : AND2_X1 port map( A1 => n20330, A2 => n3480, ZN => n20090);
   U5681 : AND2_X1 port map( A1 => n4616, A2 => n4066, ZN => n20009);
   U5682 : AND2_X1 port map( A1 => n5686, A2 => n5685, ZN => n17895);
   U5683 : OR2_X1 port map( A1 => n20071, A2 => n3240, ZN => n19661);
   U5684 : AND2_X1 port map( A1 => n20518, A2 => n20516, ZN => n19799);
   U5685 : INV_X1 port map( A => n19979, ZN => n20296);
   U5686 : INV_X1 port map( A => n20142, ZN => n20297);
   U5687 : NAND2_X1 port map( A1 => n3239, A2 => n18846, ZN => n19658);
   U5688 : OR2_X1 port map( A1 => n19406, A2 => n19407, ZN => n18782);
   U5689 : OR2_X1 port map( A1 => n25489, A2 => n19397, ZN => n4809);
   U5690 : NOR2_X1 port map( A1 => n19510, A2 => n1419, ZN => n3195);
   U5691 : INV_X1 port map( A => n20419, ZN => n4509);
   U5692 : INV_X1 port map( A => n20174, ZN => n20589);
   U5693 : NOR2_X1 port map( A1 => n20576, A2 => n20578, ZN => n20432);
   U5694 : NAND2_X1 port map( A1 => n19843, A2 => n19839, ZN => n20437);
   U5695 : OR2_X1 port map( A1 => n5207, A2 => n20194, ZN => n5206);
   U5696 : INV_X1 port map( A => n20411, ZN => n20263);
   U5698 : NAND2_X1 port map( A1 => n18974, A2 => n19478, ZN => n4402);
   U5699 : INV_X1 port map( A => n19658, ZN => n20069);
   U5700 : INV_X1 port map( A => n3428, ZN => n2432);
   U5701 : OAI21_X1 port map( B1 => n1601, B2 => n1600, A => n24454, ZN => 
                           n1599);
   U5702 : AND2_X1 port map( A1 => n20370, A2 => n20374, ZN => n1601);
   U5703 : OR2_X1 port map( A1 => n19173, A2 => n19407, ZN => n18826);
   U5704 : OAI22_X1 port map( A1 => n20280, A2 => n20279, B1 => n20343, B2 => 
                           n20345, ZN => n2699);
   U5705 : OAI21_X1 port map( B1 => n20298, B2 => n19979, A => n4615, ZN => 
                           n20302);
   U5706 : OR2_X1 port map( A1 => n19785, A2 => n24464, ZN => n19750);
   U5708 : OR2_X1 port map( A1 => n20022, A2 => n18395, ZN => n19729);
   U5709 : OR2_X1 port map( A1 => n18728, A2 => n2578, ZN => n2854);
   U5710 : AND2_X1 port map( A1 => n19490, A2 => n240, ZN => n2578);
   U5711 : OR2_X1 port map( A1 => n18717, A2 => n18990, ZN => n2304);
   U5712 : AOI21_X1 port map( B1 => n20562, B2 => n20094, A => n25221, ZN => 
                           n2469);
   U5713 : OR2_X1 port map( A1 => n20560, A2 => n20094, ZN => n2470);
   U5714 : INV_X1 port map( A => n20126, ZN => n20312);
   U5715 : AND2_X1 port map( A1 => n20345, A2 => n3671, ZN => n4460);
   U5717 : OR2_X1 port map( A1 => n20230, A2 => n343, ZN => n5425);
   U5718 : INV_X1 port map( A => n19586, ZN => n2068);
   U5719 : NOR2_X1 port map( A1 => n4480, A2 => n19592, ZN => n4479);
   U5720 : NOR2_X2 port map( A1 => n19604, A2 => n19603, ZN => n20960);
   U5723 : OR2_X1 port map( A1 => n20411, A2 => n4184, ZN => n4183);
   U5724 : OR2_X1 port map( A1 => n20591, A2 => n20588, ZN => n2724);
   U5726 : XNOR2_X1 port map( A => n21967, B => n21735, ZN => n4688);
   U5727 : AOI22_X1 port map( A1 => n17849, A2 => n20117, B1 => n3326, B2 => 
                           n25388, ZN => n3325);
   U5729 : NOR2_X1 port map( A1 => n22355, A2 => n22356, ZN => n4221);
   U5730 : INV_X1 port map( A => n19888, ZN => n4174);
   U5731 : XNOR2_X1 port map( A => n21640, B => n21596, ZN => n20831);
   U5733 : INV_X1 port map( A => n22803, ZN => n22585);
   U5735 : AND2_X1 port map( A1 => n22452, A2 => n21918, ZN => n5584);
   U5736 : NOR2_X1 port map( A1 => n22779, A2 => n22782, ZN => n22780);
   U5737 : INV_X1 port map( A => n23196, ZN => n4113);
   U5738 : INV_X1 port map( A => n22333, ZN => n21368);
   U5739 : OR2_X1 port map( A1 => n22977, A2 => n22389, ZN => n3210);
   U5740 : AOI21_X1 port map( B1 => n1766, B2 => n1765, A => n22941, ZN => 
                           n22942);
   U5741 : NAND2_X1 port map( A1 => n24932, A2 => n22829, ZN => n4608);
   U5742 : INV_X1 port map( A => n4633, ZN => n22436);
   U5743 : NOR2_X1 port map( A1 => n22959, A2 => n24885, ZN => n22858);
   U5744 : AND2_X1 port map( A1 => n24397, A2 => n23592, ZN => n21946);
   U5745 : INV_X1 port map( A => n22159, ZN => n2312);
   U5746 : INV_X1 port map( A => n21829, ZN => n1728);
   U5747 : NOR2_X1 port map( A1 => n21825, A2 => n22252, ZN => n22521);
   U5751 : NOR2_X1 port map( A1 => n331, A2 => n25241, ZN => n22609);
   U5752 : INV_X1 port map( A => n4273, ZN => n4168);
   U5753 : NAND2_X1 port map( A1 => n22363, A2 => n25241, ZN => n2528);
   U5754 : OAI21_X1 port map( B1 => n22806, B2 => n22807, A => n24992, ZN => 
                           n4427);
   U5755 : INV_X1 port map( A => n24325, ZN => n4630);
   U5756 : AND2_X1 port map( A1 => n24381, A2 => n23714, ZN => n3282);
   U5760 : OR2_X1 port map( A1 => n22450, A2 => n274, ZN => n5260);
   U5761 : INV_X1 port map( A => n23104, ZN => n23123);
   U5763 : OR2_X1 port map( A1 => n21379, A2 => n274, ZN => n5048);
   U5764 : OR2_X1 port map( A1 => n23165, A2 => n23178, ZN => n22553);
   U5765 : AOI22_X1 port map( A1 => n22324, A2 => n22325, B1 => n22452, B2 => 
                           n22456, ZN => n3682);
   U5766 : OR2_X1 port map( A1 => n23190, A2 => n23200, ZN => n3037);
   U5768 : INV_X1 port map( A => n22561, ZN => n22573);
   U5769 : INV_X1 port map( A => n3720, ZN => n2869);
   U5770 : OR2_X1 port map( A1 => n3720, A2 => n23252, ZN => n3719);
   U5771 : NAND2_X1 port map( A1 => n23252, A2 => n23253, ZN => n4243);
   U5773 : AND2_X1 port map( A1 => n3623, A2 => n22508, ZN => n2861);
   U5775 : AOI21_X1 port map( B1 => n25081, B2 => n1500, A => n24309, ZN => 
                           n2921);
   U5776 : OR2_X1 port map( A1 => n21886, A2 => n3781, ZN => n1684);
   U5777 : OR2_X1 port map( A1 => n1685, A2 => n3781, ZN => n1682);
   U5778 : OR2_X1 port map( A1 => n4372, A2 => n22972, ZN => n22978);
   U5779 : OR2_X1 port map( A1 => n22744, A2 => n4606, ZN => n4605);
   U5781 : OR2_X1 port map( A1 => n22430, A2 => n23368, ZN => n3528);
   U5782 : INV_X1 port map( A => n22026, ZN => n23392);
   U5783 : AND2_X1 port map( A1 => n23449, A2 => n22528, ZN => n4311);
   U5784 : INV_X1 port map( A => n23480, ZN => n23492);
   U5785 : OR2_X1 port map( A1 => n23480, A2 => n2710, ZN => n23485);
   U5787 : INV_X1 port map( A => n4949, ZN => n23516);
   U5788 : INV_X1 port map( A => n23531, ZN => n5701);
   U5789 : AND2_X1 port map( A1 => n23592, A2 => n23596, ZN => n5437);
   U5791 : AND3_X1 port map( A1 => n22727, A2 => n20893, A3 => n20892, ZN => 
                           n20895);
   U5792 : NOR2_X1 port map( A1 => n23645, A2 => n23634, ZN => n23629);
   U5793 : NOR2_X1 port map( A1 => n23665, A2 => n5507, ZN => n23669);
   U5794 : INV_X1 port map( A => n23727, ZN => n3283);
   U5796 : AND2_X1 port map( A1 => n24362, A2 => n4374, ZN => n23752);
   U5797 : AND2_X1 port map( A1 => n23767, A2 => n25051, ZN => n2982);
   U5798 : AND2_X1 port map( A1 => n23769, A2 => n25051, ZN => n2783);
   U5799 : OR2_X1 port map( A1 => n23789, A2 => n24307, ZN => n4954);
   U5800 : AND2_X1 port map( A1 => n22043, A2 => n23805, ZN => n3495);
   U5801 : OR2_X1 port map( A1 => n24392, A2 => n3201, ZN => n23789);
   U5802 : AND2_X1 port map( A1 => n3456, A2 => n3070, ZN => n21346);
   U5803 : OR2_X1 port map( A1 => n22214, A2 => n21341, ZN => n3070);
   U5804 : OR2_X1 port map( A1 => n21352, A2 => n21362, ZN => n4216);
   U5805 : INV_X1 port map( A => n25391, ZN => n23831);
   U5806 : AND2_X1 port map( A1 => n24428, A2 => n4186, ZN => n4192);
   U5807 : AND2_X1 port map( A1 => n25399, A2 => n23860, ZN => n4186);
   U5808 : OR2_X1 port map( A1 => n23861, A2 => n23860, ZN => n4190);
   U5810 : INV_X1 port map( A => n24006, ZN => n4478);
   U5811 : OR2_X1 port map( A1 => n4478, A2 => n24440, ZN => n4475);
   U5812 : OR2_X1 port map( A1 => n23988, A2 => n23983, ZN => n23989);
   U5813 : OR2_X1 port map( A1 => n23993, A2 => n24006, ZN => n23979);
   U5814 : INV_X1 port map( A => n24019, ZN => n24008);
   U5815 : NOR2_X1 port map( A1 => n22775, A2 => n22774, ZN => n5610);
   U5816 : AOI21_X1 port map( B1 => n2538, B2 => n23499, A => n2535, ZN => 
                           n23012);
   U5817 : OR2_X1 port map( A1 => n23058, A2 => n22699, ZN => n3914);
   U5818 : NOR2_X1 port map( A1 => n1422, A2 => n23200, ZN => n4234);
   U5819 : OAI21_X1 port map( B1 => n23218, B2 => n23219, A => n2084, ZN => 
                           n22652);
   U5820 : AND2_X1 port map( A1 => n22296, A2 => n23245, ZN => n3586);
   U5821 : OAI21_X1 port map( B1 => n22851, B2 => n2961, A => n2960, ZN => 
                           n22867);
   U5822 : OR2_X1 port map( A1 => n4032, A2 => n924, ZN => n4029);
   U5823 : AND4_X1 port map( A1 => n3441, A2 => n22085, A3 => n22084, A4 => 
                           n22083, ZN => Ciphertext(133));
   U5824 : INV_X1 port map( A => n1815, ZN => n2588);
   U5825 : NOR2_X1 port map( A1 => n24895, A2 => n22043, ZN => n2590);
   U5826 : AND2_X1 port map( A1 => n2475, A2 => n2473, ZN => n21905);
   U5827 : OR2_X1 port map( A1 => n23866, A2 => n24428, ZN => n4816);
   U5828 : AOI21_X1 port map( B1 => n22828, B2 => n25076, A => n3840, ZN => 
                           n3843);
   U5829 : INV_X1 port map( A => n20975, ZN => n5131);
   U5830 : INV_X1 port map( A => n17107, ZN => n4684);
   U5831 : XOR2_X1 port map( A => n14828, B => n14829, Z => n1371);
   U5832 : INV_X1 port map( A => n23723, ZN => n5284);
   U5833 : INV_X1 port map( A => n22354, ZN => n21844);
   U5834 : INV_X1 port map( A => n16578, ZN => n2814);
   U5835 : INV_X1 port map( A => n6560, ZN => n6934);
   U5836 : NAND3_X1 port map( A1 => n24474, A2 => n7657, A3 => n7947, ZN => 
                           n1372);
   U5837 : INV_X1 port map( A => n7589, ZN => n7588);
   U5838 : AND3_X1 port map( A1 => n5948, A2 => n5947, A3 => n5949, ZN => n7589
                           );
   U5839 : OR2_X1 port map( A1 => n9805, A2 => n9804, ZN => n1373);
   U5840 : OR2_X1 port map( A1 => n12546, A2 => n12903, ZN => n1374);
   U5841 : INV_X1 port map( A => n4897, ZN => n4541);
   U5842 : INV_X1 port map( A => n10746, ZN => n4341);
   U5843 : AND2_X1 port map( A1 => n10811, A2 => n1448, ZN => n1375);
   U5845 : XNOR2_X1 port map( A => n17992, B => n17991, ZN => n2540);
   U5846 : XNOR2_X1 port map( A => n9573, B => n3360, ZN => n13092);
   U5847 : INV_X1 port map( A => n13092, ZN => n12871);
   U5848 : AND2_X1 port map( A1 => n12767, A2 => n13216, ZN => n1376);
   U5849 : OR2_X1 port map( A1 => n25198, A2 => n13011, ZN => n1377);
   U5850 : INV_X1 port map( A => n7382, ZN => n1895);
   U5851 : OR3_X1 port map( A1 => n22941, A2 => n22829, A3 => n22832, ZN => 
                           n1378);
   U5852 : INV_X1 port map( A => n7573, ZN => n3366);
   U5853 : INV_X1 port map( A => n4880, ZN => n7651);
   U5854 : OR2_X1 port map( A1 => n6719, A2 => n6718, ZN => n1379);
   U5856 : INV_X1 port map( A => n7580, ZN => n4136);
   U5857 : INV_X1 port map( A => n23120, ZN => n5036);
   U5858 : INV_X1 port map( A => n20395, ZN => n3656);
   U5859 : AND2_X1 port map( A1 => n4136, A2 => n7575, ZN => n1380);
   U5860 : INV_X1 port map( A => n13969, ZN => n4293);
   U5861 : INV_X1 port map( A => n1535, ZN => n16615);
   U5862 : BUF_X1 port map( A => n12178, Z => n13097);
   U5863 : INV_X1 port map( A => n22809, ZN => n22812);
   U5864 : AND2_X1 port map( A1 => n16409, A2 => n14472, ZN => n1382);
   U5865 : INV_X1 port map( A => n23799, ZN => n23002);
   U5866 : XOR2_X1 port map( A => n15120, B => n1951, Z => n1383);
   U5867 : XOR2_X1 port map( A => n11847, B => n11846, Z => n1384);
   U5868 : XOR2_X1 port map( A => n9084, B => n9083, Z => n1385);
   U5869 : INV_X1 port map( A => n19613, ZN => n1806);
   U5870 : INV_X1 port map( A => n13996, ZN => n13995);
   U5871 : INV_X1 port map( A => n17391, ZN => n3317);
   U5872 : XOR2_X1 port map( A => n18269, B => n1835, Z => n1386);
   U5874 : XOR2_X1 port map( A => n12337, B => n12336, Z => n1388);
   U5875 : INV_X1 port map( A => n20588, ZN => n5093);
   U5877 : INV_X1 port map( A => n22464, ZN => n3908);
   U5879 : INV_X1 port map( A => n7767, ZN => n3013);
   U5880 : INV_X1 port map( A => n22387, ZN => n4109);
   U5881 : INV_X1 port map( A => n8934, ZN => n10922);
   U5882 : INV_X1 port map( A => n14112, ZN => n5333);
   U5883 : INV_X1 port map( A => n14850, ZN => n14416);
   U5884 : INV_X1 port map( A => n17351, ZN => n17013);
   U5885 : OR3_X1 port map( A1 => n11059, A2 => n11058, A3 => n11057, ZN => 
                           n1389);
   U5888 : INV_X1 port map( A => n3671, ZN => n20279);
   U5889 : INV_X1 port map( A => n22317, ZN => n2376);
   U5892 : INV_X1 port map( A => n12737, ZN => n5112);
   U5893 : OR3_X1 port map( A1 => n22926, A2 => n25070, A3 => n22188, ZN => 
                           n1390);
   U5894 : INV_X1 port map( A => n6498, ZN => n6271);
   U5895 : INV_X1 port map( A => n16991, ZN => n2064);
   U5896 : OR2_X1 port map( A1 => n25445, A2 => n13437, ZN => n1391);
   U5898 : AND2_X1 port map( A1 => n16002, A2 => n24366, ZN => n1392);
   U5899 : INV_X1 port map( A => n19490, ZN => n5454);
   U5900 : OR3_X1 port map( A1 => n405, A2 => n545, A3 => n4499, ZN => n1393);
   U5901 : OR2_X1 port map( A1 => n16817, A2 => n24410, ZN => n1394);
   U5903 : OR2_X1 port map( A1 => n14330, A2 => n14329, ZN => n1395);
   U5904 : OR3_X1 port map( A1 => n22107, A2 => n25070, A3 => n22927, ZN => 
                           n1396);
   U5905 : OR3_X1 port map( A1 => n22933, A2 => n22932, A3 => n25004, ZN => 
                           n1397);
   U5906 : INV_X1 port map( A => n22973, ZN => n3213);
   U5907 : INV_X1 port map( A => n13329, ZN => n4634);
   U5908 : NAND3_X1 port map( A1 => n6690, A2 => n24579, A3 => n6976, ZN => 
                           n1398);
   U5909 : OR2_X1 port map( A1 => n9625, A2 => n9681, ZN => n1399);
   U5910 : INV_X1 port map( A => n22838, ZN => n2326);
   U5911 : INV_X1 port map( A => n20549, ZN => n20124);
   U5912 : XNOR2_X1 port map( A => n8201, B => n8202, ZN => n10149);
   U5913 : INV_X1 port map( A => n10149, ZN => n9841);
   U5914 : OAI21_X1 port map( B1 => n3709, B2 => n1392, A => n4515, ZN => 
                           n16607);
   U5916 : INV_X1 port map( A => n13871, ZN => n3401);
   U5917 : INV_X1 port map( A => n16221, ZN => n16461);
   U5918 : OR2_X1 port map( A1 => n10680, A2 => n4737, ZN => n1401);
   U5919 : OR2_X1 port map( A1 => n7081, A2 => n7943, ZN => n1402);
   U5920 : XNOR2_X1 port map( A => n18145, B => n4214, ZN => n2464);
   U5921 : INV_X1 port map( A => n2464, ZN => n3412);
   U5922 : OR2_X1 port map( A1 => n4069, A2 => n10047, ZN => n1403);
   U5923 : INV_X1 port map( A => n8477, ZN => n2191);
   U5924 : INV_X1 port map( A => n12607, ZN => n13266);
   U5925 : XNOR2_X1 port map( A => n12001, B => n12000, ZN => n12607);
   U5926 : INV_X1 port map( A => n7733, ZN => n5432);
   U5927 : XNOR2_X1 port map( A => n8438, B => n8437, ZN => n10079);
   U5928 : INV_X1 port map( A => n16096, ZN => n4418);
   U5929 : OAI211_X1 port map( C1 => n19376, C2 => n19222, A => n5441, B => 
                           n5442, ZN => n20140);
   U5930 : OAI211_X1 port map( C1 => n4543, C2 => n19022, A => n4542, B => 
                           n19629, ZN => n19975);
   U5931 : INV_X1 port map( A => n19975, ZN => n20298);
   U5932 : INV_X1 port map( A => n17572, ZN => n3371);
   U5933 : INV_X1 port map( A => n9281, ZN => n9963);
   U5934 : XNOR2_X1 port map( A => n4182, B => n12271, ZN => n12865);
   U5935 : XNOR2_X1 port map( A => n18712, B => n18711, ZN => n22257);
   U5937 : AND3_X1 port map( A1 => n19112, A2 => n19233, A3 => n19608, ZN => 
                           n1404);
   U5938 : OR2_X1 port map( A1 => n7912, A2 => n7364, ZN => n1405);
   U5939 : INV_X1 port map( A => n9964, ZN => n3290);
   U5940 : INV_X1 port map( A => n20422, ZN => n1662);
   U5941 : AND2_X1 port map( A1 => n9806, A2 => n9807, ZN => n1406);
   U5942 : OR3_X1 port map( A1 => n14003, A2 => n13486, A3 => n14000, ZN => 
                           n1407);
   U5943 : INV_X1 port map( A => n12861, ZN => n5412);
   U5944 : INV_X1 port map( A => n6848, ZN => n4643);
   U5945 : XOR2_X1 port map( A => n18557, B => n18043, Z => n1408);
   U5946 : XNOR2_X1 port map( A => n8248, B => n8247, ZN => n10177);
   U5947 : XNOR2_X1 port map( A => n21518, B => n21519, ZN => n22946);
   U5948 : XNOR2_X1 port map( A => n14673, B => n14674, ZN => n16108);
   U5949 : INV_X1 port map( A => n16108, ZN => n2090);
   U5951 : XNOR2_X1 port map( A => n10530, B => n10529, ZN => n13165);
   U5952 : XOR2_X1 port map( A => n18489, B => n5286, Z => n1410);
   U5953 : XOR2_X1 port map( A => n14897, B => n21944, Z => n1411);
   U5955 : INV_X1 port map( A => n6955, ZN => n3926);
   U5957 : XNOR2_X1 port map( A => n17793, B => n17794, ZN => n19365);
   U5958 : INV_X1 port map( A => n20517, ZN => n3522);
   U5959 : INV_X1 port map( A => n17276, ZN => n17274);
   U5960 : INV_X1 port map( A => n18597, ZN => n19179);
   U5961 : AND3_X1 port map( A1 => n7855, A2 => n24072, A3 => n7721, ZN => 
                           n1413);
   U5962 : NAND3_X1 port map( A1 => n4838, A2 => n3142, A3 => n6003, ZN => 
                           n7893);
   U5963 : XOR2_X1 port map( A => n8588, B => n1776, Z => n1414);
   U5964 : OR2_X1 port map( A1 => n15625, A2 => n16147, ZN => n1415);
   U5965 : INV_X1 port map( A => n11529, ZN => n11026);
   U5966 : INV_X1 port map( A => n7862, ZN => n4536);
   U5967 : OR3_X1 port map( A1 => n17421, A2 => n17425, A3 => n17424, ZN => 
                           n1416);
   U5968 : OR2_X1 port map( A1 => n21852, A2 => n22656, ZN => n1417);
   U5969 : INV_X1 port map( A => n24572, ZN => n4225);
   U5971 : INV_X1 port map( A => n20042, ZN => n19862);
   U5972 : AND2_X1 port map( A1 => n10993, A2 => n10990, ZN => n1418);
   U5973 : XNOR2_X1 port map( A => n20709, B => n20710, ZN => n22562);
   U5974 : XNOR2_X1 port map( A => n18084, B => n5135, ZN => n18808);
   U5975 : AND2_X1 port map( A1 => n19301, A2 => n19300, ZN => n1419);
   U5976 : INV_X1 port map( A => n20597, ZN => n5044);
   U5977 : OR2_X1 port map( A1 => n20480, A2 => n20478, ZN => n1420);
   U5978 : XNOR2_X1 port map( A => n14648, B => n14647, ZN => n16073);
   U5979 : OR2_X1 port map( A1 => n5572, A2 => n19277, ZN => n1421);
   U5980 : OR2_X1 port map( A1 => n24889, A2 => n23201, ZN => n1422);
   U5981 : OR2_X1 port map( A1 => n19587, A2 => n24483, ZN => n1423);
   U5982 : INV_X1 port map( A => n16434, ZN => n17170);
   U5983 : AND2_X1 port map( A1 => n20593, A2 => n20590, ZN => n1424);
   U5984 : OR2_X1 port map( A1 => n19013, A2 => n19436, ZN => n1425);
   U5985 : OR2_X1 port map( A1 => n19584, A2 => n19105, ZN => n1426);
   U5986 : OR2_X1 port map( A1 => n19277, A2 => n19126, ZN => n1427);
   U5987 : NAND2_X1 port map( A1 => n1642, A2 => n5574, ZN => n7731);
   U5988 : INV_X1 port map( A => n7731, ZN => n5595);
   U5989 : AND2_X1 port map( A1 => n22656, A2 => n22606, ZN => n1428);
   U5990 : OR2_X1 port map( A1 => n19408, A2 => n19413, ZN => n1429);
   U5991 : AND2_X1 port map( A1 => n10596, A2 => n10935, ZN => n1430);
   U5992 : AND2_X1 port map( A1 => n22901, A2 => n22847, ZN => n1431);
   U5993 : AND2_X1 port map( A1 => n20019, A2 => n18985, ZN => n1432);
   U5994 : INV_X1 port map( A => n2321, ZN => n14090);
   U5995 : OAI211_X1 port map( C1 => n12501, C2 => n13148, A => n2575, B => 
                           n2574, ZN => n2321);
   U5996 : AND3_X1 port map( A1 => n6241, A2 => n6242, A3 => n6240, ZN => n1433
                           );
   U5997 : AND2_X1 port map( A1 => n16359, A2 => n16355, ZN => n1434);
   U5998 : OR3_X1 port map( A1 => n22505, A2 => n25063, A3 => n22722, ZN => 
                           n1435);
   U5999 : OR2_X1 port map( A1 => n19396, A2 => n19397, ZN => n1436);
   U6000 : OR3_X1 port map( A1 => n25572, A2 => n16846, A3 => n5052, ZN => 
                           n1437);
   U6001 : OR3_X1 port map( A1 => n20518, A2 => n20517, A3 => n20516, ZN => 
                           n1438);
   U6002 : INV_X1 port map( A => n10571, ZN => n3760);
   U6003 : INV_X1 port map( A => n22528, ZN => n3242);
   U6004 : AND2_X1 port map( A1 => n12471, A2 => n12773, ZN => n1439);
   U6005 : INV_X1 port map( A => n7890, ZN => n7606);
   U6006 : OR2_X1 port map( A1 => n24311, A2 => n22323, ZN => n1440);
   U6007 : INV_X1 port map( A => n13235, ZN => n12546);
   U6008 : AND2_X1 port map( A1 => n6729, A2 => n6732, ZN => n1441);
   U6009 : OR2_X1 port map( A1 => n23690, A2 => n23689, ZN => n1442);
   U6010 : INV_X1 port map( A => n20136, ZN => n1954);
   U6011 : INV_X1 port map( A => n23595, ZN => n23591);
   U6012 : OR2_X1 port map( A1 => n15670, A2 => n15915, ZN => n1444);
   U6013 : BUF_X1 port map( A => n5888, Z => n6940);
   U6015 : INV_X1 port map( A => n11116, ZN => n11111);
   U6016 : OR2_X1 port map( A1 => n14509, A2 => n14440, ZN => n1446);
   U6017 : AND2_X1 port map( A1 => n11159, A2 => n11158, ZN => n1447);
   U6018 : OR2_X1 port map( A1 => n10670, A2 => n11214, ZN => n1448);
   U6019 : AND2_X1 port map( A1 => n20126, A2 => n20124, ZN => n1449);
   U6020 : NOR2_X1 port map( A1 => n24588, A2 => n14303, ZN => n1450);
   U6021 : AND2_X1 port map( A1 => n17180, A2 => n17181, ZN => n1451);
   U6022 : OR2_X1 port map( A1 => n20437, A2 => n24940, ZN => n1452);
   U6024 : AND2_X1 port map( A1 => n9765, A2 => n9766, ZN => n1453);
   U6025 : INV_X1 port map( A => n17305, ZN => n3783);
   U6026 : INV_X1 port map( A => n21828, ZN => n3201);
   U6027 : AND2_X1 port map( A1 => n7588, A2 => n5971, ZN => n1454);
   U6028 : OR2_X1 port map( A1 => n3480, A2 => n20328, ZN => n1455);
   U6029 : OR2_X1 port map( A1 => n13316, A2 => n12945, ZN => n1456);
   U6030 : AND2_X1 port map( A1 => n331, A2 => n22656, ZN => n1457);
   U6032 : INV_X1 port map( A => n12928, ZN => n5672);
   U6033 : INV_X1 port map( A => n23714, ZN => n23716);
   U6034 : OR2_X1 port map( A1 => n13552, A2 => n24376, ZN => n1459);
   U6036 : XNOR2_X1 port map( A => n7356, B => n7355, ZN => n10125);
   U6037 : INV_X1 port map( A => n10125, ZN => n5057);
   U6038 : AND2_X1 port map( A1 => n9695, A2 => n9699, ZN => n1460);
   U6039 : XOR2_X1 port map( A => n21743, B => n860, Z => n1461);
   U6040 : NOR2_X1 port map( A1 => n23730, A2 => n24991, ZN => n1462);
   U6041 : INV_X1 port map( A => n11178, ZN => n3386);
   U6042 : AND2_X1 port map( A1 => n8318, A2 => n8319, ZN => n1463);
   U6043 : OR2_X1 port map( A1 => n25064, A2 => n1577, ZN => n1464);
   U6044 : INV_X1 port map( A => n14306, ZN => n1527);
   U6045 : INV_X1 port map( A => n20272, ZN => n20520);
   U6047 : OR2_X1 port map( A1 => n23969, A2 => n23972, ZN => n1465);
   U6049 : NOR2_X1 port map( A1 => n22159, A2 => n22158, ZN => n1467);
   U6050 : INV_X1 port map( A => n19381, ZN => n19377);
   U6051 : AND2_X1 port map( A1 => n13088, A2 => n13394, ZN => n14359);
   U6052 : AND2_X1 port map( A1 => n7506, A2 => n1379, ZN => n1468);
   U6053 : OR2_X1 port map( A1 => n20073, A2 => n20072, ZN => n1469);
   U6055 : INV_X1 port map( A => n17379, ZN => n5406);
   U6056 : OR2_X1 port map( A1 => n12793, A2 => n12792, ZN => n1471);
   U6057 : OR2_X1 port map( A1 => n15937, A2 => n24387, ZN => n1472);
   U6058 : AND2_X1 port map( A1 => n17298, A2 => n1535, ZN => n1473);
   U6059 : INV_X1 port map( A => n12540, ZN => n13220);
   U6060 : INV_X1 port map( A => n11755, ZN => n12885);
   U6061 : INV_X1 port map( A => n7590, ZN => n2035);
   U6062 : AND2_X1 port map( A1 => n14462, A2 => n3501, ZN => n1474);
   U6063 : INV_X1 port map( A => n7211, ZN => n7666);
   U6064 : NAND2_X1 port map( A1 => n4179, A2 => n13173, ZN => n14107);
   U6065 : NAND3_X1 port map( A1 => n19272, A2 => n19530, A3 => n1013, ZN => 
                           n1475);
   U6066 : INV_X1 port map( A => n4754, ZN => n4752);
   U6067 : INV_X1 port map( A => n17872, ZN => n18945);
   U6068 : BUF_X1 port map( A => n17872, Z => n19471);
   U6069 : INV_X1 port map( A => n22459, ZN => n22463);
   U6070 : OR2_X1 port map( A1 => n25058, A2 => n17362, ZN => n1476);
   U6071 : NOR2_X1 port map( A1 => n25075, A2 => n22655, ZN => n1477);
   U6072 : OR2_X1 port map( A1 => n22928, A2 => n24379, ZN => n1478);
   U6073 : INV_X1 port map( A => n17970, ZN => n5300);
   U6074 : INV_X1 port map( A => n2556, ZN => n5487);
   U6075 : OR2_X1 port map( A1 => n9236, A2 => n9416, ZN => n1479);
   U6076 : NAND2_X1 port map( A1 => n22490, A2 => n25055, ZN => n1480);
   U6077 : OR2_X1 port map( A1 => n11121, A2 => n11123, ZN => n1481);
   U6078 : NAND2_X1 port map( A1 => n22254, A2 => n21822, ZN => n1482);
   U6079 : OR2_X1 port map( A1 => n15646, A2 => n25500, ZN => n1483);
   U6080 : OR2_X1 port map( A1 => n20343, A2 => n20277, ZN => n1484);
   U6081 : OR2_X1 port map( A1 => n7782, A2 => n7418, ZN => n1485);
   U6083 : OR2_X1 port map( A1 => n20190, A2 => n20191, ZN => n1487);
   U6084 : BUF_X1 port map( A => n15674, Z => n16328);
   U6085 : AND2_X1 port map( A1 => n24954, A2 => n23993, ZN => n1488);
   U6086 : INV_X1 port map( A => n14143, ZN => n5641);
   U6087 : INV_X1 port map( A => n8527, ZN => n7087);
   U6088 : INV_X1 port map( A => n13549, ZN => n14204);
   U6089 : INV_X1 port map( A => n13569, ZN => n13589);
   U6091 : AND2_X1 port map( A1 => n19964, A2 => n349, ZN => n1489);
   U6092 : INV_X1 port map( A => n10548, ZN => n10702);
   U6093 : BUF_X1 port map( A => n12663, Z => n13152);
   U6094 : INV_X1 port map( A => n13968, ZN => n1771);
   U6095 : INV_X1 port map( A => n23327, ZN => n5659);
   U6096 : INV_X1 port map( A => n20400, ZN => n20417);
   U6097 : AND2_X1 port map( A1 => n7693, A2 => n7694, ZN => n1490);
   U6098 : OR2_X1 port map( A1 => n24498, A2 => n5131, ZN => n1491);
   U6099 : INV_X1 port map( A => n20091, ZN => n2368);
   U6100 : NAND2_X1 port map( A1 => n16990, A2 => n17039, ZN => n1492);
   U6101 : AND2_X1 port map( A1 => n20368, A2 => n20373, ZN => n3767);
   U6102 : INV_X1 port map( A => n14319, ZN => n4794);
   U6103 : OR2_X1 port map( A1 => n18912, A2 => n19138, ZN => n1493);
   U6104 : INV_X1 port map( A => n924, ZN => n4034);
   U6105 : AND2_X1 port map( A1 => n5353, A2 => n5354, ZN => n1494);
   U6106 : OR2_X1 port map( A1 => n11342, A2 => n3344, ZN => n1495);
   U6107 : INV_X1 port map( A => n21964, ZN => n2319);
   U6108 : INV_X1 port map( A => n21046, ZN => n4023);
   U6109 : INV_X1 port map( A => n2137, ZN => n4668);
   U6110 : INV_X1 port map( A => n925, ZN => n5433);
   U6111 : INV_X1 port map( A => n3155, ZN => n3901);
   U6112 : INV_X1 port map( A => n888, ZN => n1528);
   U6113 : INV_X1 port map( A => n4711, ZN => n3344);
   U6114 : INV_X1 port map( A => n22089, ZN => n5286);
   U6115 : INV_X1 port map( A => n853, ZN => n4153);
   U6116 : INV_X1 port map( A => n1831, ZN => n4761);
   U6117 : INV_X1 port map( A => n677, ZN => n5514);
   U6118 : INV_X1 port map( A => n2034, ZN => n3900);
   U6119 : INV_X1 port map( A => n763, ZN => n2964);
   U6120 : INV_X1 port map( A => n3152, ZN => n5251);
   U6121 : INV_X1 port map( A => n1935, ZN => n4589);
   U6122 : INV_X1 port map( A => n2970, ZN => n5598);
   U6123 : INV_X1 port map( A => n2743, ZN => n3208);
   U6124 : INV_X1 port map( A => Key(41), ZN => n3696);
   U6125 : NAND2_X1 port map( A1 => n1497, A2 => n1496, ZN => n17184);
   U6126 : OAI21_X1 port map( B1 => n16208, B2 => n16209, A => n16207, ZN => 
                           n1496);
   U6127 : NOR2_X1 port map( A1 => n17182, A2 => n17183, ZN => n1498);
   U6128 : NAND2_X1 port map( A1 => n10753, A2 => n1499, ZN => n4506);
   U6129 : NAND2_X1 port map( A1 => n4505, A2 => n1499, ZN => n4507);
   U6130 : NAND2_X1 port map( A1 => n10452, A2 => n1499, ZN => n10290);
   U6131 : AND2_X1 port map( A1 => n10455, A2 => n1499, ZN => n2385);
   U6132 : NAND2_X1 port map( A1 => n23334, A2 => n24341, ZN => n1500);
   U6133 : XNOR2_X2 port map( A => n21396, B => n21397, ZN => n23334);
   U6135 : NAND2_X1 port map( A1 => n4052, A2 => n18862, ZN => n19080);
   U6137 : NAND2_X1 port map( A1 => n19361, A2 => n24447, ZN => n1506);
   U6138 : AND2_X1 port map( A1 => n25392, A2 => n24312, ZN => n1505);
   U6140 : INV_X1 port map( A => n4442, ZN => n1507);
   U6141 : NAND2_X1 port map( A1 => n12827, A2 => n25466, ZN => n1508);
   U6142 : NAND2_X1 port map( A1 => n14457, A2 => n4794, ZN => n14460);
   U6143 : OR2_X1 port map( A1 => n1509, A2 => n25398, ZN => n5698);
   U6144 : INV_X1 port map( A => n6523, ZN => n1509);
   U6145 : AND2_X1 port map( A1 => n16350, A2 => n1511, ZN => n16598);
   U6146 : OAI21_X1 port map( B1 => n24890, B2 => n16595, A => n24080, ZN => 
                           n1510);
   U6147 : NAND3_X1 port map( A1 => n15885, A2 => n15890, A3 => n24587, ZN => 
                           n1511);
   U6148 : NOR2_X1 port map( A1 => n24587, A2 => n16597, ZN => n1512);
   U6149 : NAND2_X1 port map( A1 => n1513, A2 => n13116, ZN => n2097);
   U6150 : NOR2_X1 port map( A1 => n3328, A2 => n12272, ZN => n1513);
   U6151 : NOR2_X1 port map( A1 => n22800, A2 => n1514, ZN => n22659);
   U6152 : NOR2_X1 port map( A1 => n12942, A2 => n1515, ZN => n11921);
   U6153 : NAND2_X1 port map( A1 => n1515, A2 => n13317, ZN => n13321);
   U6154 : INV_X1 port map( A => n4241, ZN => n1515);
   U6156 : NAND2_X1 port map( A1 => n1516, A2 => n2562, ZN => n5316);
   U6157 : NAND2_X1 port map( A1 => n1516, A2 => n16901, ZN => n17474);
   U6158 : INV_X1 port map( A => n9694, ZN => n1517);
   U6159 : INV_X1 port map( A => n2294, ZN => n9875);
   U6160 : NAND2_X1 port map( A1 => n1520, A2 => n1518, ZN => n10534);
   U6162 : NAND2_X1 port map( A1 => n19117, A2 => n1522, ZN => n1521);
   U6163 : INV_X1 port map( A => n11057, ZN => n1523);
   U6164 : NAND2_X1 port map( A1 => n1524, A2 => n11059, ZN => n10697);
   U6165 : NOR2_X1 port map( A1 => n1218, A2 => n11057, ZN => n1524);
   U6167 : AND2_X1 port map( A1 => n24588, A2 => n14301, ZN => n12018);
   U6169 : NAND2_X1 port map( A1 => n3352, A2 => n4144, ZN => n1530);
   U6170 : NAND2_X1 port map( A1 => n1531, A2 => n431, ZN => n3352);
   U6172 : NAND4_X1 port map( A1 => n5273, A2 => n1532, A3 => n5274, A4 => 
                           n5271, ZN => n10477);
   U6173 : NAND2_X1 port map( A1 => n9127, A2 => n10064, ZN => n1534);
   U6174 : OR2_X1 port map( A1 => n1535, A2 => n17296, ZN => n16513);
   U6175 : NOR2_X1 port map( A1 => n1535, A2 => n17299, ZN => n16706);
   U6176 : OR2_X1 port map( A1 => n4508, A2 => n1535, ZN => n16703);
   U6177 : NAND3_X1 port map( A1 => n1541, A2 => n13643, A3 => n1536, ZN => 
                           n13648);
   U6178 : NAND3_X1 port map( A1 => n1538, A2 => n13079, A3 => n1537, ZN => 
                           n1536);
   U6179 : NAND3_X1 port map( A1 => n1540, A2 => n13079, A3 => n1539, ZN => 
                           n13818);
   U6180 : NAND2_X1 port map( A1 => n1543, A2 => n4340, ZN => n1540);
   U6181 : NAND2_X1 port map( A1 => n1542, A2 => n13079, ZN => n1541);
   U6182 : INV_X1 port map( A => n4340, ZN => n1542);
   U6183 : NAND2_X1 port map( A1 => n13069, A2 => n13070, ZN => n1543);
   U6184 : NOR2_X1 port map( A1 => n3423, A2 => n1545, ZN => n3422);
   U6185 : XNOR2_X2 port map( A => n4316, B => n11617, ZN => n13048);
   U6186 : XNOR2_X2 port map( A => n11605, B => n11606, ZN => n13049);
   U6187 : NAND2_X1 port map( A1 => n1546, A2 => n17042, ZN => n3372);
   U6188 : AOI21_X1 port map( B1 => n17572, B2 => n1546, A => n3004, ZN => 
                           n3003);
   U6189 : XNOR2_X2 port map( A => Plaintext(29), B => Key(29), ZN => n6531);
   U6190 : MUX2_X1 port map( A => n18881, B => n18880, S => n2464, Z => n1547);
   U6192 : NAND2_X1 port map( A1 => n2069, A2 => n3412, ZN => n1548);
   U6193 : NAND2_X1 port map( A1 => n17224, A2 => n1549, ZN => n2324);
   U6194 : AND2_X1 port map( A1 => n25433, A2 => n17225, ZN => n1549);
   U6197 : NAND2_X1 port map( A1 => n6434, A2 => n6498, ZN => n6168);
   U6198 : AND2_X1 port map( A1 => n20909, A2 => n20491, ZN => n1550);
   U6199 : XNOR2_X2 port map( A => n7654, B => n7655, ZN => n9599);
   U6200 : OR2_X1 port map( A1 => n3353, A2 => n13829, ZN => n13556);
   U6201 : OR2_X1 port map( A1 => n4545, A2 => n7932, ZN => n2164);
   U6202 : AND2_X1 port map( A1 => n7924, A2 => n7932, ZN => n5606);
   U6203 : AND2_X1 port map( A1 => n4380, A2 => n4379, ZN => n1554);
   U6204 : OR2_X1 port map( A1 => n6789, A2 => n6905, ZN => n5247);
   U6205 : INV_X1 port map( A => n7007, ZN => n7005);
   U6206 : INV_X1 port map( A => n14242, ZN => n13633);
   U6208 : INV_X1 port map( A => n4436, ZN => n19265);
   U6209 : INV_X1 port map( A => n16397, ZN => n3630);
   U6210 : INV_X1 port map( A => n7803, ZN => n7795);
   U6211 : NOR2_X1 port map( A1 => n441, A2 => n6271, ZN => n5143);
   U6212 : OR2_X1 port map( A1 => n5707, A2 => n25433, ZN => n4572);
   U6213 : AND2_X1 port map( A1 => n25450, A2 => n1363, ZN => n21928);
   U6215 : INV_X1 port map( A => n16220, ZN => n5269);
   U6217 : OR2_X1 port map( A1 => n16901, A2 => n16902, ZN => n2247);
   U6218 : XNOR2_X1 port map( A => n18285, B => n18685, ZN => n18372);
   U6219 : INV_X1 port map( A => n15746, ZN => n1654);
   U6220 : OR2_X1 port map( A1 => n24540, A2 => n25441, ZN => n4926);
   U6221 : OAI211_X1 port map( C1 => n9857, C2 => n9864, A => n25464, B => 
                           n4622, ZN => n10517);
   U6223 : INV_X1 port map( A => n2404, ZN => n7085);
   U6224 : AND2_X1 port map( A1 => n7013, A2 => n6827, ZN => n1876);
   U6225 : OR2_X1 port map( A1 => n23281, A2 => n24349, ZN => n5529);
   U6226 : OR2_X1 port map( A1 => n24411, A2 => n22962, ZN => n22964);
   U6227 : INV_X1 port map( A => n22967, ZN => n21476);
   U6228 : OR2_X1 port map( A1 => n2587, A2 => n16550, ZN => n2508);
   U6229 : INV_X1 port map( A => n16550, ZN => n16794);
   U6230 : OR2_X1 port map( A1 => n16550, A2 => n16796, ZN => n16619);
   U6231 : OR2_X1 port map( A1 => n12648, A2 => n12178, ZN => n5321);
   U6232 : AND2_X1 port map( A1 => n24549, A2 => n9692, ZN => n9028);
   U6233 : OR2_X1 port map( A1 => n24549, A2 => n9027, ZN => n3117);
   U6234 : XNOR2_X1 port map( A => n1813, B => n8789, ZN => n8549);
   U6235 : INV_X1 port map( A => n8366, ZN => n1813);
   U6236 : XNOR2_X1 port map( A => n21215, B => n20223, ZN => n3871);
   U6238 : INV_X1 port map( A => n24547, ZN => n4334);
   U6239 : OR2_X1 port map( A1 => n6444, A2 => n6445, ZN => n6021);
   U6240 : OR2_X1 port map( A1 => n23069, A2 => n23064, ZN => n4990);
   U6241 : OR2_X1 port map( A1 => n12652, A2 => n403, ZN => n3935);
   U6243 : OR2_X1 port map( A1 => n25477, A2 => n20597, ZN => n5365);
   U6244 : XNOR2_X1 port map( A => n11309, B => n3647, ZN => n12792);
   U6245 : OAI21_X1 port map( B1 => n7893, B2 => n7604, A => n7606, ZN => n7326
                           );
   U6246 : NOR2_X1 port map( A1 => n9782, A2 => n9781, ZN => n9676);
   U6247 : AND2_X1 port map( A1 => n2718, A2 => n15811, ZN => n3316);
   U6248 : INV_X1 port map( A => n13888, ZN => n13945);
   U6249 : OAI21_X1 port map( B1 => n9064, B2 => n10050, A => n9866, ZN => 
                           n9869);
   U6250 : AOI21_X1 port map( B1 => n9064, B2 => n9244, A => n24446, ZN => 
                           n3489);
   U6251 : AND2_X1 port map( A1 => n9064, A2 => n24092, ZN => n10054);
   U6253 : AND2_X1 port map( A1 => n3195, A2 => n19939, ZN => n19817);
   U6254 : AND2_X1 port map( A1 => n19302, A2 => n19133, ZN => n3568);
   U6255 : NOR2_X1 port map( A1 => n388, A2 => n15667, ZN => n15917);
   U6256 : OR2_X1 port map( A1 => n14510, A2 => n13974, ZN => n3777);
   U6257 : INV_X1 port map( A => n13974, ZN => n14436);
   U6258 : NOR2_X1 port map( A1 => n13161, A2 => n12454, ZN => n5013);
   U6259 : AND2_X1 port map( A1 => n23869, A2 => n23905, ZN => n23888);
   U6260 : NOR2_X1 port map( A1 => n25414, A2 => n25079, ZN => n2616);
   U6262 : AND2_X1 port map( A1 => n25001, A2 => n19598, ZN => n4715);
   U6264 : OR2_X1 port map( A1 => n6775, A2 => n6292, ZN => n6293);
   U6265 : OR2_X1 port map( A1 => n6775, A2 => n6777, ZN => n2353);
   U6266 : NOR2_X1 port map( A1 => n10464, A2 => n10720, ZN => n4500);
   U6267 : AOI22_X1 port map( A1 => n7827, A2 => n7985, B1 => n7984, B2 => 
                           n7046, ZN => n7513);
   U6268 : AND2_X1 port map( A1 => n7985, A2 => n7983, ZN => n1690);
   U6269 : OR2_X1 port map( A1 => n7827, A2 => n7985, ZN => n2082);
   U6270 : INV_X1 port map( A => n21140, ZN => n22779);
   U6271 : INV_X1 port map( A => n18290, ZN => n17637);
   U6272 : OR2_X1 port map( A1 => n3472, A2 => n10125, ZN => n9379);
   U6273 : XNOR2_X1 port map( A => n15267, B => n15160, ZN => n3669);
   U6275 : AND2_X1 port map( A1 => n24321, A2 => n23303, ZN => n23300);
   U6276 : OR2_X1 port map( A1 => n24321, A2 => n23303, ZN => n3623);
   U6277 : OR2_X1 port map( A1 => n20255, A2 => n25421, ZN => n5189);
   U6278 : NOR2_X1 port map( A1 => n18895, A2 => n19526, ZN => n19720);
   U6279 : OAI22_X1 port map( A1 => n5003, A2 => n18795, B1 => n19526, B2 => 
                           n5496, ZN => n19528);
   U6280 : INV_X1 port map( A => n19526, ZN => n19283);
   U6282 : OR2_X1 port map( A1 => n22868, A2 => n23411, ZN => n2961);
   U6283 : AND2_X1 port map( A1 => n24421, A2 => n19290, ZN => n3094);
   U6284 : INV_X1 port map( A => n12792, ZN => n4680);
   U6285 : AND2_X1 port map( A1 => n13228, A2 => n12792, ZN => n13229);
   U6286 : AND2_X1 port map( A1 => n12792, A2 => n12995, ZN => n2837);
   U6287 : OR2_X1 port map( A1 => n7008, A2 => n7004, ZN => n6833);
   U6288 : XNOR2_X1 port map( A => n24413, B => n8981, ZN => n8183);
   U6289 : OR2_X1 port map( A1 => n22162, A2 => n22221, ZN => n21830);
   U6290 : OAI21_X1 port map( B1 => n18994, B2 => n20316, A => n20319, ZN => 
                           n2179);
   U6291 : AND2_X1 port map( A1 => n12993, A2 => n4587, ZN => n13230);
   U6292 : OR2_X1 port map( A1 => n12791, A2 => n12993, ZN => n5041);
   U6293 : OR2_X1 port map( A1 => n9449, A2 => n9907, ZN => n9936);
   U6294 : AND2_X1 port map( A1 => n23273, A2 => n25550, ZN => n22535);
   U6296 : AND2_X1 port map( A1 => n22409, A2 => n22407, ZN => n22133);
   U6297 : OR2_X1 port map( A1 => n22562, A2 => n22407, ZN => n1588);
   U6298 : OR2_X1 port map( A1 => n16109, A2 => n16108, ZN => n2020);
   U6299 : INV_X1 port map( A => n12272, ZN => n13113);
   U6300 : OR2_X1 port map( A1 => n6795, A2 => n6076, ZN => n3894);
   U6301 : OR2_X1 port map( A1 => n23555, A2 => n23546, ZN => n5397);
   U6302 : INV_X1 port map( A => n16452, ZN => n16235);
   U6303 : NOR2_X1 port map( A1 => n12785, A2 => n13027, ZN => n1635);
   U6304 : INV_X1 port map( A => n12785, ZN => n13029);
   U6305 : OAI21_X1 port map( B1 => n20963, B2 => n24354, A => n20962, ZN => 
                           n21452);
   U6306 : INV_X1 port map( A => n16192, ZN => n16196);
   U6307 : XNOR2_X1 port map( A => n15218, B => n14955, ZN => n2862);
   U6312 : AND2_X1 port map( A1 => n16266, A2 => n25009, ZN => n5667);
   U6313 : OAI22_X1 port map( A1 => n3287, A2 => n12824, B1 => n13288, B2 => 
                           n13289, ZN => n13297);
   U6314 : XNOR2_X1 port map( A => n15430, B => n15523, ZN => n15106);
   U6315 : OR2_X1 port map( A1 => n16356, A2 => n16290, ZN => n4846);
   U6316 : OAI21_X1 port map( B1 => n3517, B2 => n367, A => n3514, ZN => n3706)
                           ;
   U6317 : AOI22_X1 port map( A1 => n17356, A2 => n17351, B1 => n17012, B2 => 
                           n25491, ZN => n3517);
   U6318 : XNOR2_X1 port map( A => n21601, B => n21675, ZN => n21023);
   U6319 : AND2_X1 port map( A1 => n19366, A2 => n19370, ZN => n19098);
   U6321 : NOR2_X1 port map( A1 => n12459, A2 => n12724, ZN => n3968);
   U6323 : NOR2_X1 port map( A1 => n8021, A2 => n7278, ZN => n3259);
   U6324 : INV_X1 port map( A => n24415, ZN => n4350);
   U6326 : OAI211_X1 port map( C1 => n13119, C2 => n12660, A => n2571, B => 
                           n12865, ZN => n12422);
   U6327 : INV_X1 port map( A => n9989, ZN => n9747);
   U6329 : INV_X1 port map( A => n18982, ZN => n20137);
   U6330 : OR2_X1 port map( A1 => n3822, A2 => n17607, ZN => n16941);
   U6332 : OR2_X1 port map( A1 => n22099, A2 => n22729, ZN => n2981);
   U6333 : INV_X1 port map( A => n22729, ZN => n3837);
   U6334 : INV_X1 port map( A => n19300, ZN => n18970);
   U6335 : INV_X1 port map( A => n2607, ZN => n16229);
   U6336 : AND2_X1 port map( A1 => n16492, A2 => n24387, ZN => n5169);
   U6337 : OR2_X1 port map( A1 => n10007, A2 => n9484, ZN => n9722);
   U6338 : OR2_X1 port map( A1 => n6814, A2 => n6815, ZN => n2800);
   U6339 : NAND2_X1 port map( A1 => n18763, A2 => n4172, ZN => n1556);
   U6340 : NAND3_X1 port map( A1 => n1733, A2 => n20343, A3 => n1557, ZN => 
                           n19650);
   U6341 : NAND2_X1 port map( A1 => n1558, A2 => n4752, ZN => n1862);
   U6342 : NAND2_X1 port map( A1 => n4752, A2 => n1559, ZN => n6406);
   U6344 : OAI21_X1 port map( B1 => n8146, B2 => n10927, A => n1562, ZN => 
                           n10408);
   U6345 : NAND2_X1 port map( A1 => n10407, A2 => n10927, ZN => n1562);
   U6346 : NAND3_X1 port map( A1 => n13349, A2 => n13346, A3 => n12861, ZN => 
                           n2023);
   U6347 : NAND2_X1 port map( A1 => n6937, A2 => n1563, ZN => n6562);
   U6348 : NAND2_X1 port map( A1 => n6559, A2 => n6934, ZN => n1563);
   U6349 : INV_X1 port map( A => n12611, ZN => n13304);
   U6352 : NAND2_X1 port map( A1 => n13304, A2 => n12555, ZN => n1566);
   U6354 : INV_X1 port map( A => n12555, ZN => n13303);
   U6355 : XNOR2_X1 port map( A => n1568, B => n3093, ZN => n11336);
   U6356 : XNOR2_X1 port map( A => n1568, B => n2881, ZN => n12010);
   U6357 : XNOR2_X1 port map( A => n1568, B => n14398, ZN => n10706);
   U6358 : XNOR2_X1 port map( A => n1568, B => n2782, ZN => n11483);
   U6359 : XNOR2_X1 port map( A => n1568, B => n12314, ZN => n11614);
   U6360 : XNOR2_X1 port map( A => n1568, B => n12391, ZN => n12392);
   U6361 : OAI21_X1 port map( B1 => n11038, B2 => n10942, A => n1569, ZN => 
                           n11040);
   U6362 : NAND2_X1 port map( A1 => n10941, A2 => n11036, ZN => n1569);
   U6363 : NAND2_X1 port map( A1 => n11037, A2 => n11036, ZN => n1570);
   U6364 : NAND2_X1 port map( A1 => n10571, A2 => n10941, ZN => n11037);
   U6366 : NAND2_X1 port map( A1 => n12689, A2 => n12946, ZN => n1572);
   U6367 : NAND2_X1 port map( A1 => n7634, A2 => n1573, ZN => n7160);
   U6368 : NAND2_X1 port map( A1 => n1574, A2 => n25253, ZN => n1573);
   U6369 : NAND2_X1 port map( A1 => n7915, A2 => n7917, ZN => n1574);
   U6370 : NAND3_X1 port map( A1 => n1575, A2 => n6491, A3 => n6492, ZN => 
                           n7915);
   U6371 : INV_X1 port map( A => Plaintext(59), ZN => n1576);
   U6373 : INV_X1 port map( A => n10166, ZN => n1577);
   U6374 : NOR2_X1 port map( A1 => n12555, A2 => n25248, ZN => n13306);
   U6375 : NAND2_X1 port map( A1 => n12914, A2 => n12613, ZN => n1578);
   U6376 : NAND2_X1 port map( A1 => n1579, A2 => n14264, ZN => n5693);
   U6377 : AND2_X2 port map( A1 => n1583, A2 => n1580, ZN => n21115);
   U6378 : NAND2_X1 port map( A1 => n25383, A2 => n2432, ZN => n1581);
   U6379 : NAND2_X1 port map( A1 => n19963, A2 => n20369, ZN => n1582);
   U6380 : AOI21_X1 port map( B1 => n3767, B2 => n24558, A => n1489, ZN => 
                           n1583);
   U6381 : AND2_X1 port map( A1 => n17472, A2 => n17629, ZN => n1842);
   U6383 : NAND2_X1 port map( A1 => n22133, A2 => n1586, ZN => n1585);
   U6384 : NAND2_X1 port map( A1 => n22566, A2 => n22563, ZN => n1586);
   U6385 : NAND2_X1 port map( A1 => n22343, A2 => n22406, ZN => n1587);
   U6386 : NAND4_X1 port map( A1 => n4235, A2 => n1589, A3 => n4233, A4 => 
                           n4237, ZN => n4232);
   U6387 : NAND2_X1 port map( A1 => n1590, A2 => n20448, ZN => n20449);
   U6388 : NOR2_X1 port map( A1 => n1590, A2 => n20451, ZN => n20158);
   U6390 : NAND2_X1 port map( A1 => n1591, A2 => n20100, ZN => n17946);
   U6391 : AND2_X1 port map( A1 => n1591, A2 => n20103, ZN => n2358);
   U6392 : NOR2_X1 port map( A1 => n1591, A2 => n20101, ZN => n19915);
   U6393 : NAND2_X1 port map( A1 => n21033, A2 => n1591, ZN => n20105);
   U6394 : OAI21_X1 port map( B1 => n21033, B2 => n1591, A => n20101, ZN => 
                           n19156);
   U6395 : OAI21_X1 port map( B1 => n7645, B2 => n5595, A => n1592, ZN => n7569
                           );
   U6396 : NAND3_X1 port map( A1 => n25151, A2 => n24578, A3 => n7640, ZN => 
                           n1592);
   U6397 : NAND2_X1 port map( A1 => n4018, A2 => n6237, ZN => n1643);
   U6398 : INV_X1 port map( A => n22409, ZN => n1593);
   U6399 : OR2_X1 port map( A1 => n22341, A2 => n24971, ZN => n22568);
   U6400 : AOI22_X2 port map( A1 => n22343, A2 => n22412, B1 => n22342, B2 => 
                           n326, ZN => n23166);
   U6401 : NOR2_X1 port map( A1 => n9964, A2 => n1595, ZN => n9965);
   U6403 : AOI21_X1 port map( B1 => n9469, B2 => n1595, A => n9964, ZN => n8142
                           );
   U6405 : MUX2_X1 port map( A => n9964, B => n9203, S => n3292, Z => n9204);
   U6406 : AOI21_X1 port map( B1 => n1597, B2 => n7854, A => n1596, ZN => n1598
                           );
   U6407 : OR2_X1 port map( A1 => n7722, A2 => n7721, ZN => n1597);
   U6408 : OAI21_X2 port map( B1 => n1598, B2 => n1413, A => n7724, ZN => n8478
                           );
   U6409 : NOR2_X1 port map( A1 => n20370, A2 => n20369, ZN => n1600);
   U6412 : MUX2_X1 port map( A => n20368, B => n20370, S => n3428, Z => n1604);
   U6414 : AND2_X1 port map( A1 => n22592, A2 => n1605, ZN => n21189);
   U6415 : NAND2_X1 port map( A1 => n25066, A2 => n1605, ZN => n22450);
   U6416 : NOR2_X1 port map( A1 => n25066, A2 => n1605, ZN => n21923);
   U6417 : INV_X1 port map( A => n7735, ZN => n7641);
   U6418 : NAND2_X1 port map( A1 => n1607, A2 => n7735, ZN => n7644);
   U6419 : NAND2_X1 port map( A1 => n1608, A2 => n7732, ZN => n1607);
   U6420 : NAND2_X1 port map( A1 => n7731, A2 => n7733, ZN => n1608);
   U6421 : INV_X1 port map( A => n5796, ZN => n6049);
   U6422 : INV_X1 port map( A => n5796, ZN => n1609);
   U6423 : NAND2_X1 port map( A1 => n1610, A2 => n6728, ZN => n1642);
   U6424 : INV_X1 port map( A => n16830, ZN => n1611);
   U6426 : NAND2_X1 port map( A1 => n2688, A2 => n1614, ZN => n2687);
   U6427 : NOR2_X1 port map( A1 => n16714, A2 => n17312, ZN => n1616);
   U6428 : NAND2_X1 port map( A1 => n16715, A2 => n17304, ZN => n1615);
   U6429 : INV_X1 port map( A => n17304, ZN => n17597);
   U6430 : OAI211_X2 port map( C1 => n18815, C2 => n19384, A => n18814, B => 
                           n1617, ZN => n20491);
   U6431 : NAND2_X1 port map( A1 => n19633, A2 => n1617, ZN => n19636);
   U6432 : NAND2_X1 port map( A1 => n18813, A2 => n24909, ZN => n1617);
   U6433 : AND2_X1 port map( A1 => n1619, A2 => n23649, ZN => n23606);
   U6434 : NAND2_X1 port map( A1 => n23638, A2 => n1618, ZN => n23641);
   U6435 : AND3_X1 port map( A1 => n23640, A2 => n23639, A3 => n1619, ZN => 
                           n1618);
   U6436 : NAND3_X1 port map( A1 => n23638, A2 => n23640, A3 => n1619, ZN => 
                           n23631);
   U6437 : NAND2_X1 port map( A1 => n1622, A2 => n1620, ZN => n16348);
   U6438 : NAND2_X1 port map( A1 => n1621, A2 => n16345, ZN => n1620);
   U6439 : NOR2_X1 port map( A1 => n1654, A2 => n16342, ZN => n1621);
   U6440 : NAND2_X1 port map( A1 => n16346, A2 => n16281, ZN => n1622);
   U6442 : AOI21_X1 port map( B1 => n1624, B2 => n16764, A => n17274, ZN => 
                           n1623);
   U6443 : NAND2_X1 port map( A1 => n17248, A2 => n17273, ZN => n16764);
   U6445 : AOI21_X1 port map( B1 => n16762, B2 => n17252, A => n1626, ZN => 
                           n1625);
   U6446 : INV_X1 port map( A => n17275, ZN => n1626);
   U6447 : NAND2_X1 port map( A1 => n24300, A2 => n17272, ZN => n16762);
   U6448 : AND2_X1 port map( A1 => n22158, A2 => n2315, ZN => n22211);
   U6449 : OR2_X1 port map( A1 => n2315, A2 => n22158, ZN => n22065);
   U6450 : NAND2_X1 port map( A1 => n1467, A2 => n2315, ZN => n22161);
   U6451 : OAI22_X2 port map( A1 => n21771, A2 => n21770, B1 => n21769, B2 => 
                           n1627, ZN => n23596);
   U6452 : INV_X1 port map( A => n2315, ZN => n1627);
   U6453 : AND2_X1 port map( A1 => n18982, A2 => n1629, ZN => n5566);
   U6454 : NAND2_X1 port map( A1 => n19992, A2 => n25378, ZN => n19993);
   U6456 : NAND2_X1 port map( A1 => n1432, A2 => n25378, ZN => n5563);
   U6457 : NAND2_X1 port map( A1 => n13131, A2 => n13151, ZN => n13153);
   U6458 : NAND3_X1 port map( A1 => n13131, A2 => n1774, A3 => n13152, ZN => 
                           n1630);
   U6459 : NAND2_X1 port map( A1 => n13133, A2 => n13132, ZN => n1631);
   U6460 : NAND2_X1 port map( A1 => n24376, A2 => n13552, ZN => n4600);
   U6461 : NAND2_X1 port map( A1 => n14268, A2 => n14267, ZN => n13623);
   U6462 : NAND2_X1 port map( A1 => n1636, A2 => n1635, ZN => n1633);
   U6463 : NAND2_X1 port map( A1 => n3371, A2 => n17571, ZN => n1639);
   U6464 : NAND2_X1 port map( A1 => n3374, A2 => n17572, ZN => n1640);
   U6465 : NAND4_X1 port map( A1 => n1641, A2 => n1643, A3 => n7733, A4 => 
                           n1642, ZN => n7567);
   U6466 : NAND2_X1 port map( A1 => n1645, A2 => n1644, ZN => n22522);
   U6467 : OR2_X1 port map( A1 => n24362, A2 => n21841, ZN => n1644);
   U6468 : NAND2_X1 port map( A1 => n21822, A2 => n21841, ZN => n1645);
   U6469 : XNOR2_X2 port map( A => n19054, B => n19053, ZN => n21841);
   U6470 : NAND3_X1 port map( A1 => n21798, A2 => n21796, A3 => n21797, ZN => 
                           n23772);
   U6471 : NAND2_X1 port map( A1 => n1646, A2 => n12800, ZN => n12481);
   U6472 : NAND2_X1 port map( A1 => n1646, A2 => n12797, ZN => n4618);
   U6473 : NAND2_X1 port map( A1 => n1648, A2 => n1647, ZN => n9583);
   U6474 : NAND2_X1 port map( A1 => n10136, A2 => n10138, ZN => n1647);
   U6475 : NAND3_X1 port map( A1 => n9367, A2 => n9366, A3 => n1649, ZN => 
                           n9371);
   U6476 : MUX2_X1 port map( A => n5742, B => n9400, S => n10138, Z => n9401);
   U6477 : OAI21_X1 port map( B1 => n9201, B2 => n10146, A => n1649, ZN => 
                           n9202);
   U6478 : NAND2_X1 port map( A1 => n17145, A2 => n1653, ZN => n16848);
   U6480 : AOI21_X1 port map( B1 => n16496, B2 => n1653, A => n16847, ZN => 
                           n16497);
   U6482 : NAND2_X1 port map( A1 => n15977, A2 => n15849, ZN => n1655);
   U6483 : NAND2_X1 port map( A1 => n10284, A2 => n1658, ZN => n3532);
   U6485 : NAND2_X1 port map( A1 => n1658, A2 => n11113, ZN => n11114);
   U6487 : INV_X1 port map( A => n20430, ZN => n20209);
   U6488 : NAND2_X1 port map( A1 => n20400, A2 => n1663, ZN => n1661);
   U6489 : NOR2_X1 port map( A1 => n20415, A2 => n20419, ZN => n1663);
   U6490 : NAND2_X1 port map( A1 => n1666, A2 => n20597, ZN => n1665);
   U6491 : NAND2_X1 port map( A1 => n19846, A2 => n20599, ZN => n1666);
   U6492 : INV_X1 port map( A => n25477, ZN => n1667);
   U6493 : NAND2_X1 port map( A1 => n9718, A2 => n9635, ZN => n9436);
   U6494 : NAND2_X1 port map( A1 => n1672, A2 => n9634, ZN => n1671);
   U6495 : OAI21_X1 port map( B1 => n9434, B2 => n9710, A => n9714, ZN => n1672
                           );
   U6497 : NAND3_X1 port map( A1 => n16095, A2 => n15625, A3 => n16147, ZN => 
                           n1676);
   U6498 : XNOR2_X2 port map( A => n14567, B => n14566, ZN => n16095);
   U6499 : NAND2_X1 port map( A1 => n1677, A2 => n4247, ZN => n7528);
   U6500 : NAND2_X1 port map( A1 => n22113, A2 => n1678, ZN => n1680);
   U6501 : NOR2_X1 port map( A1 => n22072, A2 => n22917, ZN => n1678);
   U6504 : NOR2_X1 port map( A1 => n1681, A2 => n12768, ZN => n12769);
   U6505 : OAI21_X1 port map( B1 => n1681, B2 => n4651, A => n13218, ZN => 
                           n4547);
   U6506 : NAND2_X1 port map( A1 => n13215, A2 => n12767, ZN => n1681);
   U6508 : OR2_X1 port map( A1 => n21887, A2 => n22263, ZN => n1685);
   U6509 : NAND2_X1 port map( A1 => n1685, A2 => n21886, ZN => n1683);
   U6510 : AND2_X1 port map( A1 => n382, A2 => n16067, ZN => n16065);
   U6511 : AOI21_X1 port map( B1 => n380, B2 => n16064, A => n16060, ZN => 
                           n15796);
   U6512 : INV_X1 port map( A => n11128, ZN => n1689);
   U6516 : NAND3_X1 port map( A1 => n10839, A2 => n11129, A3 => n1689, ZN => 
                           n10716);
   U6517 : NAND3_X1 port map( A1 => n10840, A2 => n420, A3 => n1689, ZN => 
                           n10843);
   U6518 : NAND2_X1 port map( A1 => n1690, A2 => n7048, ZN => n6852);
   U6519 : OR2_X1 port map( A1 => n21774, A2 => n1691, ZN => n2513);
   U6520 : NAND2_X1 port map( A1 => n327, A2 => n22728, ZN => n1691);
   U6521 : NAND2_X1 port map( A1 => n7034, A2 => n454, ZN => n1692);
   U6522 : NAND2_X1 port map( A1 => n2270, A2 => n7035, ZN => n1693);
   U6523 : MUX2_X1 port map( A => n1345, B => n270, S => n7682, Z => n7071);
   U6524 : INV_X1 port map( A => n12964, ZN => n1694);
   U6525 : NAND2_X1 port map( A1 => n6740, A2 => n6739, ZN => n1695);
   U6526 : OAI21_X1 port map( B1 => n434, B2 => n7674, A => n7676, ZN => n7673)
                           ;
   U6527 : INV_X1 port map( A => n1696, ZN => n1697);
   U6528 : XNOR2_X2 port map( A => n5969, B => Key(179), ZN => n1698);
   U6529 : NAND2_X1 port map( A1 => n5966, A2 => n1698, ZN => n6468);
   U6530 : NAND2_X1 port map( A1 => n1697, A2 => n5449, ZN => n5450);
   U6531 : NOR2_X1 port map( A1 => n6469, A2 => n1698, ZN => n7692);
   U6532 : XNOR2_X1 port map( A => n11661, B => n1699, ZN => n10707);
   U6533 : XNOR2_X1 port map( A => n11750, B => n1700, ZN => n11752);
   U6534 : INV_X1 port map( A => n11661, ZN => n1700);
   U6535 : XNOR2_X1 port map( A => n25493, B => n18157, ZN => n18305);
   U6536 : NAND2_X1 port map( A1 => n15834, A2 => n25472, ZN => n1702);
   U6537 : NAND3_X1 port map( A1 => n1704, A2 => n17729, A3 => n17485, ZN => 
                           n1703);
   U6538 : NAND3_X1 port map( A1 => n17735, A2 => n24410, A3 => n17093, ZN => 
                           n1705);
   U6539 : OAI211_X1 port map( C1 => n19361, C2 => n25392, A => n1707, B => 
                           n19211, ZN => n1706);
   U6540 : NAND2_X1 port map( A1 => n25392, A2 => n19359, ZN => n1707);
   U6541 : NAND3_X1 port map( A1 => n15779, A2 => n15778, A3 => n15777, ZN => 
                           n17075);
   U6542 : INV_X1 port map( A => n17075, ZN => n17077);
   U6543 : OR2_X1 port map( A1 => n7460, A2 => n268, ZN => n1904);
   U6547 : OAI21_X1 port map( B1 => n19549, B2 => n1710, A => n19403, ZN => 
                           n2722);
   U6548 : INV_X1 port map( A => n19548, ZN => n1711);
   U6549 : NAND2_X1 port map( A1 => n19552, A2 => n1713, ZN => n1712);
   U6550 : AND2_X1 port map( A1 => n19185, A2 => n25057, ZN => n1713);
   U6551 : NAND2_X1 port map( A1 => n19552, A2 => n19185, ZN => n1714);
   U6552 : NOR2_X1 port map( A1 => n25057, A2 => n1715, ZN => n19725);
   U6553 : NAND2_X1 port map( A1 => n19546, A2 => n19186, ZN => n1715);
   U6557 : NAND2_X1 port map( A1 => n16038, A2 => n2253, ZN => n1718);
   U6560 : NAND2_X1 port map( A1 => n10573, A2 => n11037, ZN => n10575);
   U6561 : NAND2_X1 port map( A1 => n1721, A2 => n1720, ZN => n18941);
   U6562 : NAND2_X1 port map( A1 => n18937, A2 => n19327, ZN => n1720);
   U6563 : NAND2_X1 port map( A1 => n18936, A2 => n19328, ZN => n1721);
   U6564 : NAND2_X2 port map( A1 => n1722, A2 => n21296, ZN => n23828);
   U6565 : XNOR2_X2 port map( A => n1723, B => n7436, ZN => n3472);
   U6566 : XNOR2_X1 port map( A => n7552, B => n7435, ZN => n1723);
   U6567 : XNOR2_X1 port map( A => n11517, B => n11516, ZN => n11533);
   U6568 : OAI21_X1 port map( B1 => n12550, B2 => n13001, A => n1725, ZN => 
                           n12553);
   U6571 : XNOR2_X1 port map( A => n4386, B => n8702, ZN => n9737);
   U6572 : NOR2_X1 port map( A1 => n20264, A2 => n20262, ZN => n19741);
   U6573 : INV_X1 port map( A => n7863, ZN => n3570);
   U6574 : XNOR2_X1 port map( A => n25436, B => n14952, ZN => n14915);
   U6576 : NOR2_X1 port map( A1 => n18756, A2 => n5239, ZN => n5238);
   U6577 : OR2_X1 port map( A1 => n21385, A2 => n21918, ZN => n1727);
   U6578 : NAND3_X2 port map( A1 => n5288, A2 => n9373, A3 => n5740, ZN => 
                           n10756);
   U6579 : MUX2_X1 port map( A => n20515, B => n20514, S => n20517, Z => n20275
                           );
   U6580 : NAND2_X1 port map( A1 => n19267, A2 => n19266, ZN => n1729);
   U6581 : NAND2_X1 port map( A1 => n19268, A2 => n18917, ZN => n1730);
   U6582 : OAI21_X1 port map( B1 => n24399, B2 => n17559, A => n1731, ZN => 
                           n18759);
   U6583 : NAND2_X1 port map( A1 => n19264, A2 => n19261, ZN => n1731);
   U6585 : OAI21_X1 port map( B1 => n20343, B2 => n24414, A => n1732, ZN => 
                           n20278);
   U6586 : NAND2_X1 port map( A1 => n1733, A2 => n20346, ZN => n1732);
   U6587 : INV_X1 port map( A => n20277, ZN => n1733);
   U6588 : NAND3_X1 port map( A1 => n6403, A2 => n6401, A3 => n5805, ZN => 
                           n1734);
   U6589 : OAI21_X1 port map( B1 => n7563, B2 => n7853, A => n24072, ZN => 
                           n1737);
   U6590 : NAND3_X1 port map( A1 => n24977, A2 => n23416, A3 => n25035, ZN => 
                           n1738);
   U6591 : NAND3_X1 port map( A1 => n22563, A2 => n22562, A3 => n22409, ZN => 
                           n20714);
   U6592 : NAND3_X2 port map( A1 => n16816, A2 => n16815, A3 => n1394, ZN => 
                           n18149);
   U6593 : AOI21_X1 port map( B1 => n16112, B2 => n17170, A => n17171, ZN => 
                           n16134);
   U6595 : NOR2_X2 port map( A1 => n20283, A2 => n2138, ZN => n20475);
   U6596 : NOR2_X1 port map( A1 => n17437, A2 => n1782, ZN => n1781);
   U6599 : NAND2_X1 port map( A1 => n1741, A2 => n7826, ZN => n6855);
   U6600 : OAI21_X1 port map( B1 => n7828, B2 => n7048, A => n7825, ZN => n1741
                           );
   U6601 : NAND2_X1 port map( A1 => n14508, A2 => n14509, ZN => n14512);
   U6602 : NAND2_X1 port map( A1 => n13693, A2 => n24556, ZN => n14509);
   U6604 : NAND3_X1 port map( A1 => n14124, A2 => n14206, A3 => n14204, ZN => 
                           n3850);
   U6605 : NAND2_X1 port map( A1 => n24574, A2 => n10284, ZN => n9580);
   U6606 : NAND2_X1 port map( A1 => n2930, A2 => n2931, ZN => n5912);
   U6608 : NAND3_X1 port map( A1 => n4116, A2 => n14240, A3 => n13200, ZN => 
                           n4117);
   U6609 : NAND2_X1 port map( A1 => n7216, A2 => n1743, ZN => n1742);
   U6610 : INV_X1 port map( A => n2404, ZN => n1743);
   U6611 : NAND2_X1 port map( A1 => n7215, A2 => n2404, ZN => n1744);
   U6612 : NAND2_X1 port map( A1 => n6504, A2 => n6501, ZN => n6437);
   U6614 : AOI22_X1 port map( A1 => n3366, A2 => n7575, B1 => n7573, B2 => 
                           n7574, ZN => n3500);
   U6615 : NAND2_X1 port map( A1 => n14220, A2 => n14225, ZN => n1748);
   U6616 : AND2_X1 port map( A1 => n4884, A2 => n19237, ZN => n19610);
   U6617 : NAND2_X1 port map( A1 => n5387, A2 => n7913, ZN => n1749);
   U6618 : OAI21_X1 port map( B1 => n9187, B2 => n9397, A => n10141, ZN => 
                           n1751);
   U6619 : XNOR2_X1 port map( A => n1752, B => n23063, ZN => Ciphertext(5));
   U6620 : NAND2_X1 port map( A1 => n1834, A2 => n23061, ZN => n1752);
   U6621 : NAND2_X1 port map( A1 => n1753, A2 => n24043, ZN => n22594);
   U6622 : NAND2_X1 port map( A1 => n5046, A2 => n2393, ZN => n1753);
   U6624 : OR2_X1 port map( A1 => n13211, A2 => n13207, ZN => n13006);
   U6625 : NAND2_X1 port map( A1 => n5651, A2 => n6772, ZN => n5650);
   U6626 : NOR2_X1 port map( A1 => n19910, A2 => n19911, ZN => n1755);
   U6627 : XNOR2_X2 port map( A => n6035, B => Key(7), ZN => n6351);
   U6628 : XNOR2_X1 port map( A => n17813, B => n17812, ZN => n1759);
   U6629 : NAND2_X1 port map( A1 => n1761, A2 => n1760, ZN => n4420);
   U6630 : NAND2_X1 port map( A1 => n15864, A2 => n16095, ZN => n1760);
   U6631 : NAND2_X1 port map( A1 => n16151, A2 => n16149, ZN => n15864);
   U6632 : NAND2_X1 port map( A1 => n1415, A2 => n1762, ZN => n1761);
   U6633 : NAND3_X1 port map( A1 => n6752, A2 => n6578, A3 => n6751, ZN => 
                           n6402);
   U6634 : OAI21_X1 port map( B1 => n4772, B2 => n4773, A => n15952, ZN => 
                           n1763);
   U6635 : NAND2_X1 port map( A1 => n3413, A2 => n3414, ZN => n1764);
   U6636 : NAND2_X1 port map( A1 => n22939, A2 => n24932, ZN => n1765);
   U6637 : NAND2_X1 port map( A1 => n22027, A2 => n22938, ZN => n1766);
   U6639 : INV_X1 port map( A => n23869, ZN => n23889);
   U6641 : NAND3_X1 port map( A1 => n3268, A2 => n2522, A3 => n7758, ZN => 
                           n1769);
   U6642 : NAND3_X1 port map( A1 => n13157, A2 => n13151, A3 => n25033, ZN => 
                           n13154);
   U6644 : OR2_X2 port map( A1 => n13659, A2 => n13660, ZN => n12669);
   U6645 : NAND2_X1 port map( A1 => n1773, A2 => n1772, ZN => n13659);
   U6646 : NAND2_X1 port map( A1 => n12664, A2 => n13148, ZN => n1772);
   U6647 : INV_X1 port map( A => n13148, ZN => n1774);
   U6648 : XNOR2_X2 port map( A => n5879, B => Key(32), ZN => n5903);
   U6649 : NAND2_X1 port map( A1 => n1941, A2 => n10763, ZN => n10896);
   U6650 : NAND2_X1 port map( A1 => n18739, A2 => n18977, ZN => n17888);
   U6651 : NAND2_X2 port map( A1 => n20106, A2 => n2010, ZN => n21469);
   U6652 : INV_X1 port map( A => n10713, ZN => n10840);
   U6653 : OAI211_X1 port map( C1 => n13217, C2 => n12986, A => n4945, B => 
                           n13218, ZN => n12765);
   U6654 : NAND2_X1 port map( A1 => n13902, A2 => n4524, ZN => n13957);
   U6655 : NAND2_X1 port map( A1 => n6474, A2 => n6789, ZN => n6476);
   U6656 : XNOR2_X2 port map( A => n5979, B => Key(121), ZN => n7004);
   U6657 : OR2_X1 port map( A1 => n9064, A2 => n10050, ZN => n3998);
   U6658 : XNOR2_X2 port map( A => n5965, B => Key(177), ZN => n4621);
   U6660 : OR2_X1 port map( A1 => n15637, A2 => n16397, ZN => n2420);
   U6661 : NAND2_X1 port map( A1 => n1779, A2 => n1778, ZN => n7888);
   U6662 : NAND2_X1 port map( A1 => n7885, A2 => n7884, ZN => n1778);
   U6664 : NAND2_X1 port map( A1 => n1612, A2 => n1780, ZN => n17444);
   U6665 : NAND2_X1 port map( A1 => n17436, A2 => n1781, ZN => n1780);
   U6666 : NAND3_X1 port map( A1 => n17434, A2 => n17435, A3 => n17433, ZN => 
                           n1782);
   U6669 : NAND2_X1 port map( A1 => n1784, A2 => n13067, ZN => n1783);
   U6670 : NAND2_X1 port map( A1 => n12472, A2 => n12471, ZN => n1784);
   U6671 : XNOR2_X2 port map( A => Key(99), B => Plaintext(99), ZN => n7029);
   U6673 : OAI21_X1 port map( B1 => n1460, B2 => n9697, A => n1785, ZN => n9701
                           );
   U6674 : NAND2_X1 port map( A1 => n9698, A2 => n9697, ZN => n1785);
   U6675 : NAND2_X1 port map( A1 => n7288, A2 => n1786, ZN => n7287);
   U6676 : INV_X1 port map( A => n7510, ZN => n2262);
   U6677 : OAI21_X1 port map( B1 => n1788, B2 => n13096, A => n1787, ZN => 
                           n13100);
   U6678 : NAND2_X1 port map( A1 => n13096, A2 => n13095, ZN => n1787);
   U6679 : NAND2_X1 port map( A1 => n13097, A2 => n12871, ZN => n1788);
   U6680 : INV_X1 port map( A => n8221, ZN => n7811);
   U6681 : MUX2_X1 port map( A => n8220, B => n7812, S => n8221, Z => n7815);
   U6682 : NOR2_X1 port map( A1 => n15706, A2 => n4897, ZN => n1790);
   U6683 : OAI21_X1 port map( B1 => n15824, B2 => n24080, A => n2336, ZN => 
                           n1791);
   U6684 : INV_X1 port map( A => n9884, ZN => n5739);
   U6685 : INV_X1 port map( A => n19774, ZN => n20461);
   U6686 : OR2_X1 port map( A1 => n15803, A2 => n17134, ZN => n15807);
   U6687 : NAND2_X1 port map( A1 => n20372, A2 => n19962, ZN => n1793);
   U6688 : XNOR2_X1 port map( A => n15021, B => n15020, ZN => n4957);
   U6689 : NAND2_X1 port map( A1 => n19760, A2 => n18385, ZN => n1982);
   U6691 : INV_X1 port map( A => n16095, ZN => n16097);
   U6692 : INV_X1 port map( A => n9769, ZN => n10681);
   U6693 : XNOR2_X1 port map( A => n12167, B => n12295, ZN => n11946);
   U6694 : XNOR2_X1 port map( A => n3471, B => n14598, ZN => n2000);
   U6695 : OR3_X1 port map( A1 => n11169, A2 => n11171, A3 => n8660, ZN => 
                           n3384);
   U6696 : NAND2_X1 port map( A1 => n3982, A2 => n16528, ZN => n16529);
   U6697 : NAND2_X1 port map( A1 => n1795, A2 => n1794, ZN => n10001);
   U6698 : NAND2_X1 port map( A1 => n246, A2 => n9998, ZN => n1794);
   U6699 : NAND2_X1 port map( A1 => n25453, A2 => n1796, ZN => n1795);
   U6700 : INV_X1 port map( A => n9997, ZN => n1796);
   U6702 : AOI21_X1 port map( B1 => n6134, B2 => n6164, A => n6162, ZN => n1798
                           );
   U6703 : NAND2_X1 port map( A1 => n16219, A2 => n16220, ZN => n16216);
   U6704 : OR2_X1 port map( A1 => n9832, A2 => n9829, ZN => n9827);
   U6705 : NAND2_X1 port map( A1 => n6156, A2 => n6523, ZN => n6278);
   U6707 : NAND2_X1 port map( A1 => n9564, A2 => n9565, ZN => n9884);
   U6709 : XNOR2_X1 port map( A => n4670, B => n3512, ZN => n11690);
   U6710 : NAND2_X1 port map( A1 => n350, A2 => n3657, ZN => n20462);
   U6712 : NAND3_X1 port map( A1 => n2326, A2 => n22893, A3 => n22835, ZN => 
                           n1802);
   U6713 : NAND2_X1 port map( A1 => n5766, A2 => n25438, ZN => n1803);
   U6714 : INV_X1 port map( A => n6997, ZN => n3109);
   U6716 : OAI211_X1 port map( C1 => n19239, C2 => n278, A => n3919, B => n1805
                           , ZN => n3918);
   U6718 : INV_X1 port map( A => n20218, ZN => n1809);
   U6719 : OAI21_X1 port map( B1 => n4684, B2 => n17130, A => n1811, ZN => 
                           n16789);
   U6720 : NAND2_X1 port map( A1 => n4684, A2 => n25227, ZN => n1811);
   U6721 : XNOR2_X2 port map( A => n5871, B => Key(42), ZN => n5924);
   U6722 : NAND2_X1 port map( A1 => n2892, A2 => n5105, ZN => n10934);
   U6723 : AND2_X1 port map( A1 => n7604, A2 => n7323, ZN => n2552);
   U6724 : NAND2_X1 port map( A1 => n13216, A2 => n13217, ZN => n12539);
   U6725 : AND2_X2 port map( A1 => n5297, A2 => n5298, ZN => n15446);
   U6726 : INV_X1 port map( A => n16171, ZN => n15820);
   U6727 : NAND2_X1 port map( A1 => n6487, A2 => n6301, ZN => n6302);
   U6729 : NAND2_X1 port map( A1 => n3064, A2 => n3066, ZN => n12529);
   U6730 : AND3_X2 port map( A1 => n14887, A2 => n14888, A3 => n15925, ZN => 
                           n17608);
   U6731 : OAI21_X1 port map( B1 => n348, B2 => n4065, A => n20476, ZN => n5244
                           );
   U6732 : NOR2_X1 port map( A1 => n16539, A2 => n2247, ZN => n2246);
   U6733 : XNOR2_X2 port map( A => n11318, B => n11317, ZN => n12993);
   U6734 : NAND2_X1 port map( A1 => n25246, A2 => n17413, ZN => n17418);
   U6735 : NAND2_X1 port map( A1 => n7792, A2 => n7793, ZN => n8366);
   U6736 : NAND2_X1 port map( A1 => n2160, A2 => n6326, ZN => n6327);
   U6738 : NAND2_X1 port map( A1 => n9753, A2 => n9613, ZN => n1814);
   U6739 : NAND2_X1 port map( A1 => n10855, A2 => n25230, ZN => n10282);
   U6740 : NAND2_X1 port map( A1 => n5065, A2 => n5066, ZN => n1816);
   U6741 : NAND2_X1 port map( A1 => n16310, A2 => n1817, ZN => n16313);
   U6742 : AND3_X1 port map( A1 => n250, A2 => n6848, A3 => n7025, ZN => n2738)
                           ;
   U6743 : OR2_X1 port map( A1 => n15846, A2 => n16154, ZN => n2992);
   U6744 : NAND2_X1 port map( A1 => n1818, A2 => n2544, ZN => n2543);
   U6745 : XNOR2_X1 port map( A => n3931, B => n5513, ZN => n16440);
   U6746 : INV_X1 port map( A => n17130, ZN => n3458);
   U6747 : NAND2_X1 port map( A1 => n13891, A2 => n1819, ZN => n15523);
   U6748 : NAND2_X1 port map( A1 => n1820, A2 => n13728, ZN => n1819);
   U6749 : NAND2_X1 port map( A1 => n13889, A2 => n13944, ZN => n1820);
   U6751 : OR2_X1 port map( A1 => n15929, A2 => n15725, ZN => n15730);
   U6752 : INV_X1 port map( A => n13394, ZN => n2629);
   U6753 : OR2_X1 port map( A1 => n6556, A2 => n6414, ZN => n6935);
   U6754 : INV_X1 port map( A => n13807, ZN => n14035);
   U6755 : INV_X1 port map( A => n9681, ZN => n4069);
   U6756 : INV_X1 port map( A => n15583, ZN => n5100);
   U6757 : XNOR2_X1 port map( A => n2077, B => n11906, ZN => n5749);
   U6758 : INV_X1 port map( A => n24542, ZN => n17598);
   U6759 : XNOR2_X1 port map( A => n3233, B => n15191, ZN => n15155);
   U6761 : XNOR2_X1 port map( A => n12214, B => n11990, ZN => n1821);
   U6762 : NAND3_X2 port map( A1 => n5527, A2 => n5525, A3 => n13588, ZN => 
                           n15230);
   U6763 : NAND2_X1 port map( A1 => n1823, A2 => n1436, ZN => n1822);
   U6764 : INV_X1 port map( A => n18901, ZN => n1823);
   U6765 : NAND2_X1 port map( A1 => n11201, A2 => n10630, ZN => n1824);
   U6766 : NAND3_X1 port map( A1 => n6949, A2 => n6255, A3 => n5903, ZN => 
                           n5528);
   U6767 : NAND2_X1 port map( A1 => n1825, A2 => n377, ZN => n5546);
   U6768 : NOR2_X1 port map( A1 => n15695, A2 => n25238, ZN => n1825);
   U6769 : NAND2_X1 port map( A1 => n1441, A2 => n6731, ZN => n1922);
   U6770 : NAND2_X1 port map( A1 => n6734, A2 => n6238, ZN => n6731);
   U6772 : NAND2_X1 port map( A1 => n20909, A2 => n20491, ZN => n20483);
   U6773 : NAND3_X1 port map( A1 => n16262, A2 => n16261, A3 => n25219, ZN => 
                           n16263);
   U6774 : NAND2_X1 port map( A1 => n353, A2 => n19125, ZN => n5571);
   U6775 : XOR2_X1 port map( A => n18281, B => n18280, Z => n3753);
   U6776 : INV_X1 port map( A => n13302, ZN => n1828);
   U6777 : NAND2_X1 port map( A1 => n9664, A2 => n9985, ZN => n9742);
   U6778 : NAND2_X1 port map( A1 => n2668, A2 => n2669, ZN => n2238);
   U6779 : NAND3_X2 port map( A1 => n4889, A2 => n1402, A3 => n1372, ZN => 
                           n8787);
   U6780 : OAI21_X1 port map( B1 => n25223, B2 => n25347, A => n1996, ZN => 
                           n19816);
   U6781 : AOI22_X1 port map( A1 => n1830, A2 => n6468, B1 => n5451, B2 => 
                           n6467, ZN => n7690);
   U6782 : NAND2_X1 port map( A1 => n25404, A2 => n6425, ZN => n1830);
   U6783 : OR2_X1 port map( A1 => n23062, A2 => n322, ZN => n1834);
   U6784 : INV_X1 port map( A => n10100, ZN => n9836);
   U6785 : OAI21_X1 port map( B1 => n17003, B2 => n17051, A => n3643, ZN => 
                           n3646);
   U6789 : XNOR2_X1 port map( A => n10601, B => n3565, ZN => n10602);
   U6790 : INV_X1 port map( A => n5971, ZN => n1839);
   U6791 : NAND2_X1 port map( A1 => n1842, A2 => n17473, ZN => n1841);
   U6792 : INV_X1 port map( A => n4503, ZN => n5884);
   U6793 : NAND2_X1 port map( A1 => n1844, A2 => n1843, ZN => n12501);
   U6794 : NAND2_X1 port map( A1 => n25033, A2 => n13130, ZN => n1843);
   U6795 : OAI21_X1 port map( B1 => n10254, B2 => n5057, A => n9379, ZN => 
                           n5289);
   U6796 : OAI211_X1 port map( C1 => n15972, C2 => n15971, A => n3630, B => 
                           n1845, ZN => n3629);
   U6797 : NAND2_X1 port map( A1 => n15971, A2 => n1846, ZN => n1845);
   U6798 : INV_X1 port map( A => n15638, ZN => n1846);
   U6799 : NAND2_X1 port map( A1 => n1847, A2 => n1275, ZN => n4255);
   U6800 : NAND2_X1 port map( A1 => n10110, A2 => n10107, ZN => n1847);
   U6801 : INV_X1 port map( A => n9121, ZN => n7895);
   U6802 : NAND2_X1 port map( A1 => n7888, A2 => n7887, ZN => n9121);
   U6803 : NAND2_X1 port map( A1 => n4676, A2 => n4675, ZN => n3555);
   U6804 : NAND2_X1 port map( A1 => n1850, A2 => n1849, ZN => n4676);
   U6805 : NAND2_X1 port map( A1 => n2479, A2 => n25030, ZN => n1849);
   U6806 : NAND2_X1 port map( A1 => n2480, A2 => n24586, ZN => n1850);
   U6807 : NAND2_X1 port map( A1 => n6455, A2 => n25428, ZN => n6507);
   U6808 : NAND3_X1 port map( A1 => n17024, A2 => n2230, A3 => n1852, ZN => 
                           n17026);
   U6811 : NAND2_X1 port map( A1 => n17015, A2 => n17208, ZN => n16557);
   U6812 : NAND2_X1 port map( A1 => n19888, A2 => n20316, ZN => n3541);
   U6813 : NAND2_X1 port map( A1 => n2251, A2 => n15263, ZN => n15264);
   U6814 : INV_X1 port map( A => n15319, ZN => n15126);
   U6815 : INV_X1 port map( A => n13583, ZN => n14105);
   U6816 : NAND2_X1 port map( A1 => n9993, A2 => n24534, ZN => n1857);
   U6817 : NAND2_X1 port map( A1 => n9994, A2 => n422, ZN => n1858);
   U6820 : NAND2_X1 port map( A1 => n12637, A2 => n398, ZN => n1859);
   U6821 : NAND2_X1 port map( A1 => n12638, A2 => n1861, ZN => n1860);
   U6822 : INV_X1 port map( A => n398, ZN => n1861);
   U6824 : XNOR2_X1 port map( A => n24472, B => n1381, ZN => n20839);
   U6827 : NAND2_X1 port map( A1 => n3324, A2 => n10757, ZN => n9364);
   U6828 : NAND2_X1 port map( A1 => n14008, A2 => n14252, ZN => n13701);
   U6829 : NAND2_X1 port map( A1 => n15925, A2 => n3778, ZN => n1872);
   U6830 : NAND2_X1 port map( A1 => n3380, A2 => n15904, ZN => n14138);
   U6831 : OAI21_X1 port map( B1 => n5246, B2 => n14042, A => n298, ZN => n2155
                           );
   U6832 : NAND2_X1 port map( A1 => n6755, A2 => n6673, ZN => n6579);
   U6833 : OR3_X1 port map( A1 => n7350, A2 => n7349, A3 => n7346, ZN => n7352)
                           ;
   U6834 : NAND3_X1 port map( A1 => n19530, A2 => n19270, A3 => n24329, ZN => 
                           n5654);
   U6835 : OAI22_X1 port map( A1 => n13773, A2 => n14179, B1 => n13774, B2 => 
                           n24949, ZN => n1866);
   U6836 : NOR2_X1 port map( A1 => n14088, A2 => n14092, ZN => n1868);
   U6838 : NAND2_X1 port map( A1 => n12845, A2 => n1456, ZN => n12846);
   U6839 : NAND2_X1 port map( A1 => n12947, A2 => n12945, ZN => n12845);
   U6840 : OAI211_X1 port map( C1 => n16724, C2 => n2666, A => n2665, B => 
                           n2664, ZN => n17676);
   U6841 : NAND3_X1 port map( A1 => n312, A2 => n7636, A3 => n435, ZN => n6495)
                           ;
   U6842 : XNOR2_X1 port map( A => n15150, B => n14414, ZN => n3308);
   U6843 : XNOR2_X1 port map( A => n15159, B => n15161, ZN => n3670);
   U6844 : OAI21_X1 port map( B1 => n15314, B2 => n17240, A => n17346, ZN => 
                           n15473);
   U6845 : NAND2_X1 port map( A1 => n7580, A2 => n7573, ZN => n3548);
   U6847 : INV_X1 port map( A => n16029, ZN => n16273);
   U6848 : NOR2_X1 port map( A1 => n6818, A2 => n6895, ZN => n3414);
   U6849 : NAND2_X1 port map( A1 => n2290, A2 => n12794, ZN => n2048);
   U6850 : NAND2_X1 port map( A1 => n12991, A2 => n4587, ZN => n12794);
   U6851 : NAND2_X1 port map( A1 => n1872, A2 => n16459, ZN => n15704);
   U6853 : OR3_X1 port map( A1 => n14130, A2 => n14127, A3 => n14126, ZN => 
                           n13407);
   U6854 : NAND2_X1 port map( A1 => n22771, A2 => n22774, ZN => n22773);
   U6855 : NAND2_X1 port map( A1 => n5498, A2 => n14256, ZN => n14259);
   U6856 : XNOR2_X1 port map( A => n4590, B => n12196, ZN => n12095);
   U6857 : OR2_X1 port map( A1 => n1971, A2 => n4861, ZN => n4860);
   U6858 : NAND2_X1 port map( A1 => n3616, A2 => n7747, ZN => n1873);
   U6859 : INV_X1 port map( A => n11806, ZN => n13963);
   U6861 : OAI21_X1 port map( B1 => n271, B2 => n6752, A => n2494, ZN => n2496)
                           ;
   U6862 : AOI21_X1 port map( B1 => n16851, B2 => n16850, A => n2105, ZN => 
                           n16853);
   U6863 : INV_X1 port map( A => n5255, ZN => n8671);
   U6864 : INV_X1 port map( A => n12636, ZN => n13348);
   U6865 : INV_X1 port map( A => n10613, ZN => n10412);
   U6866 : INV_X1 port map( A => n13305, ZN => n12917);
   U6867 : INV_X1 port map( A => n10596, ZN => n10936);
   U6868 : INV_X1 port map( A => n11070, ZN => n11068);
   U6869 : INV_X1 port map( A => n13906, ZN => n15410);
   U6870 : INV_X1 port map( A => n13868, ZN => n14458);
   U6871 : OAI21_X1 port map( B1 => n7313, B2 => n7582, A => n7314, ZN => n7470
                           );
   U6872 : INV_X1 port map( A => n8667, ZN => n8039);
   U6873 : INV_X1 port map( A => n12003, ZN => n2917);
   U6874 : INV_X1 port map( A => n8203, ZN => n9052);
   U6875 : INV_X1 port map( A => n223, ZN => n15726);
   U6876 : INV_X1 port map( A => n24012, ZN => n4477);
   U6877 : XNOR2_X1 port map( A => n14486, B => n14485, ZN => n15612);
   U6878 : OAI211_X1 port map( C1 => n15573, C2 => n15572, A => n2651, B => 
                           n16274, ZN => n2648);
   U6879 : XNOR2_X1 port map( A => n15153, B => n1920, ZN => n14841);
   U6880 : NAND2_X1 port map( A1 => n7015, A2 => n1876, ZN => n6828);
   U6885 : NAND2_X1 port map( A1 => n7564, A2 => n6413, ZN => n1880);
   U6886 : NAND2_X1 port map( A1 => n6925, A2 => n6480, ZN => n6923);
   U6887 : NAND2_X1 port map( A1 => n20559, A2 => n20092, ZN => n1881);
   U6888 : NAND2_X1 port map( A1 => n405, A2 => n13235, ZN => n5359);
   U6889 : NAND2_X1 port map( A1 => n4617, A2 => n16461, ZN => n14887);
   U6890 : AND3_X2 port map( A1 => n12572, A2 => n12571, A3 => n12570, ZN => 
                           n14075);
   U6891 : NAND2_X1 port map( A1 => n1883, A2 => n1882, ZN => n16669);
   U6892 : OR3_X1 port map( A1 => n17347, A2 => n17241, A3 => n17342, ZN => 
                           n1882);
   U6894 : XNOR2_X1 port map( A => n14403, B => n14891, ZN => n1884);
   U6896 : NAND2_X1 port map( A1 => n1885, A2 => n5361, ZN => n5360);
   U6897 : NAND2_X1 port map( A1 => n407, A2 => n13264, ZN => n1885);
   U6898 : AOI21_X1 port map( B1 => n9329, B2 => n9503, A => n1886, ZN => n9333
                           );
   U6899 : NAND2_X1 port map( A1 => n2011, A2 => n9736, ZN => n9430);
   U6902 : OAI21_X1 port map( B1 => n10536, B2 => n4998, A => n10535, ZN => 
                           n1887);
   U6905 : AOI22_X1 port map( A1 => n9845, A2 => n10151, B1 => n10152, B2 => 
                           n9843, ZN => n10154);
   U6906 : OAI21_X1 port map( B1 => n10669, B2 => n24340, A => n1910, ZN => 
                           n11218);
   U6908 : MUX2_X1 port map( A => n6878, B => n6877, S => n6876, Z => n1888);
   U6910 : NAND3_X1 port map( A1 => n385, A2 => n16448, A3 => n223, ZN => 
                           n15728);
   U6911 : OAI21_X1 port map( B1 => n7943, B2 => n4259, A => n1892, ZN => n7229
                           );
   U6912 : NAND2_X1 port map( A1 => n7943, A2 => n7942, ZN => n1892);
   U6913 : NAND2_X1 port map( A1 => n13460, A2 => n14307, ZN => n13902);
   U6917 : INV_X1 port map( A => n15861, ZN => n16116);
   U6918 : OR2_X1 port map( A1 => n10303, A2 => n10302, ZN => n5678);
   U6919 : NAND2_X1 port map( A1 => n16535, A2 => n4774, ZN => n16536);
   U6920 : XNOR2_X2 port map( A => n21628, B => n21629, ZN => n22832);
   U6921 : NAND2_X1 port map( A1 => n13171, A2 => n11597, ZN => n1893);
   U6922 : NAND2_X1 port map( A1 => n11596, A2 => n13165, ZN => n1894);
   U6923 : NAND3_X1 port map( A1 => n7617, A2 => n7384, A3 => n1895, ZN => 
                           n7202);
   U6924 : XNOR2_X1 port map( A => n8190, B => n8189, ZN => n9842);
   U6926 : NOR2_X1 port map( A1 => n3817, A2 => n16974, ZN => n3815);
   U6927 : OAI21_X1 port map( B1 => n3578, B2 => n15790, A => n1897, ZN => 
                           n3576);
   U6932 : NAND2_X1 port map( A1 => n1902, A2 => n1901, ZN => n7603);
   U6933 : NAND2_X1 port map( A1 => n7600, A2 => n7595, ZN => n1901);
   U6934 : INV_X1 port map( A => n12541, ZN => n4651);
   U6935 : XNOR2_X1 port map( A => n8558, B => n3048, ZN => n1903);
   U6936 : NAND2_X1 port map( A1 => n22831, A2 => n337, ZN => n1905);
   U6937 : XNOR2_X2 port map( A => n5937, B => Key(1), ZN => n6456);
   U6938 : NAND2_X1 port map( A1 => n9306, A2 => n9788, ZN => n8455);
   U6939 : INV_X1 port map( A => n16048, ZN => n15606);
   U6940 : NAND2_X1 port map( A1 => n294, A2 => n16048, ZN => n4624);
   U6941 : AND2_X1 port map( A1 => n7749, A2 => n8012, ZN => n7535);
   U6944 : NAND2_X1 port map( A1 => n24570, A2 => n372, ZN => n1909);
   U6945 : NAND2_X1 port map( A1 => n24340, A2 => n11216, ZN => n1910);
   U6946 : NAND2_X1 port map( A1 => n16389, A2 => n1912, ZN => n1911);
   U6947 : NOR2_X1 port map( A1 => n15977, A2 => n16394, ZN => n1912);
   U6948 : NAND2_X1 port map( A1 => n14546, A2 => n15977, ZN => n1913);
   U6949 : OAI21_X1 port map( B1 => n17069, B2 => n369, A => n1914, ZN => 
                           n15610);
   U6950 : NAND2_X1 port map( A1 => n17065, A2 => n16731, ZN => n1914);
   U6952 : NAND2_X1 port map( A1 => n1916, A2 => n1915, ZN => n12733);
   U6953 : NAND2_X1 port map( A1 => n11109, A2 => n13144, ZN => n1916);
   U6954 : OR2_X1 port map( A1 => n11210, A2 => n11209, ZN => n1918);
   U6956 : NOR2_X1 port map( A1 => n19791, A2 => n174, ZN => n5338);
   U6957 : NOR2_X1 port map( A1 => n9760, A2 => n9764, ZN => n10076);
   U6958 : AOI22_X2 port map( A1 => n10609, A2 => n10966, B1 => n10608, B2 => 
                           n1919, ZN => n12031);
   U6959 : AOI21_X1 port map( B1 => n10607, B2 => n10970, A => n10606, ZN => 
                           n1919);
   U6961 : OR2_X1 port map( A1 => n10444, A2 => n10751, ZN => n10447);
   U6962 : NAND2_X1 port map( A1 => n260, A2 => n10044, ZN => n10047);
   U6963 : OR2_X1 port map( A1 => n2576, A2 => n6658, ZN => n3110);
   U6964 : NAND2_X1 port map( A1 => n24998, A2 => n23689, ZN => n23688);
   U6965 : INV_X1 port map( A => n16962, ZN => n17441);
   U6966 : NOR2_X1 port map( A1 => n23464, A2 => n23014, ZN => n22863);
   U6967 : OAI21_X1 port map( B1 => n3422, B2 => n13051, A => n3420, ZN => 
                           n13386);
   U6968 : INV_X1 port map( A => n8928, ZN => n8557);
   U6969 : INV_X1 port map( A => n17321, ZN => n15673);
   U6970 : XNOR2_X1 port map( A => n15175, B => n15003, ZN => n5210);
   U6971 : NAND2_X1 port map( A1 => n12526, A2 => n12796, ZN => n3066);
   U6972 : OR2_X1 port map( A1 => n10907, A2 => n10901, ZN => n4342);
   U6973 : INV_X1 port map( A => n17386, ZN => n17179);
   U6974 : OR2_X1 port map( A1 => n11067, A2 => n11062, ZN => n10059);
   U6975 : INV_X1 port map( A => n10128, ZN => n10254);
   U6976 : INV_X1 port map( A => n4422, ZN => n5559);
   U6977 : INV_X1 port map( A => n13279, ZN => n13283);
   U6978 : INV_X1 port map( A => n8157, ZN => n9567);
   U6979 : INV_X1 port map( A => n8119, ZN => n9190);
   U6980 : INV_X1 port map( A => n17410, ZN => n4487);
   U6981 : INV_X1 port map( A => n23326, ZN => n3564);
   U6982 : NOR2_X1 port map( A1 => n3544, A2 => n16202, ZN => n3543);
   U6983 : INV_X1 port map( A => n2674, ZN => n22420);
   U6984 : INV_X1 port map( A => n9140, ZN => n5346);
   U6985 : AOI21_X1 port map( B1 => n22948, B2 => n22947, A => n2673, ZN => 
                           n22949);
   U6986 : NOR2_X1 port map( A1 => n17616, A2 => n17609, ZN => n17610);
   U6987 : XNOR2_X1 port map( A => n13710, B => n13709, ZN => n3779);
   U6988 : XNOR2_X1 port map( A => n8615, B => n8616, ZN => n9090);
   U6989 : XNOR2_X1 port map( A => Plaintext(185), B => Key(185), ZN => n4866);
   U6990 : OAI22_X1 port map( A1 => n24492, A2 => n23350, B1 => n23354, B2 => 
                           n23359, ZN => n23363);
   U6991 : XNOR2_X1 port map( A => n12219, B => n11542, ZN => n11787);
   U6992 : OAI21_X2 port map( B1 => n2008, B2 => n5900, A => n5899, ZN => n7897
                           );
   U6993 : NAND2_X1 port map( A1 => n2459, A2 => n7911, ZN => n2458);
   U6994 : OAI22_X1 port map( A1 => n25432, A2 => n16349, B1 => n16595, B2 => 
                           n24467, ZN => n15671);
   U6995 : NAND2_X1 port map( A1 => n16225, A2 => n15774, ZN => n16024);
   U6996 : NAND3_X1 port map( A1 => n2306, A2 => n24420, A3 => n10369, ZN => 
                           n1921);
   U6997 : NAND2_X1 port map( A1 => n2461, A2 => n7628, ZN => n2460);
   U6998 : NAND2_X1 port map( A1 => n6617, A2 => n1922, ZN => n7787);
   U6999 : INV_X1 port map( A => n17463, ZN => n5052);
   U7000 : NAND3_X1 port map( A1 => n2721, A2 => n12635, A3 => n1923, ZN => 
                           n14200);
   U7001 : NAND3_X1 port map( A1 => n12633, A2 => n4529, A3 => n12632, ZN => 
                           n1923);
   U7003 : NAND3_X1 port map( A1 => n1459, A2 => n25445, A3 => n13417, ZN => 
                           n13553);
   U7004 : OAI21_X2 port map( B1 => n7639, B2 => n7638, A => n1928, ZN => n8760
                           );
   U7005 : NAND2_X1 port map( A1 => n7637, A2 => n7915, ZN => n1928);
   U7006 : XNOR2_X1 port map( A => n1929, B => n11991, ZN => n10672);
   U7007 : XNOR2_X1 port map( A => n10647, B => n10646, ZN => n1929);
   U7008 : NAND2_X1 port map( A1 => n24082, A2 => n11338, ZN => n2675);
   U7010 : XNOR2_X1 port map( A => n1931, B => n23401, ZN => Ciphertext(84));
   U7011 : NAND3_X1 port map( A1 => n2630, A2 => n23400, A3 => n23399, ZN => 
                           n1931);
   U7013 : AOI22_X1 port map( A1 => n1933, A2 => n1932, B1 => n13584, B2 => 
                           n1932, ZN => n5708);
   U7014 : INV_X1 port map( A => n4868, ZN => n1932);
   U7015 : OR2_X1 port map( A1 => n7358, A2 => n7412, ZN => n7360);
   U7016 : INV_X1 port map( A => n25201, ZN => n17211);
   U7017 : NAND2_X1 port map( A1 => n4491, A2 => n4492, ZN => n14126);
   U7018 : OAI21_X1 port map( B1 => n21362, B2 => n21363, A => n1934, ZN => 
                           n21364);
   U7019 : INV_X1 port map( A => n16691, ZN => n16496);
   U7020 : NOR2_X1 port map( A1 => n19659, A2 => n3241, ZN => n1936);
   U7021 : XNOR2_X1 port map( A => n17829, B => n17830, ZN => n19459);
   U7023 : OAI21_X1 port map( B1 => n16965, B2 => n17127, A => n17445, ZN => 
                           n17661);
   U7025 : NAND2_X1 port map( A1 => n1938, A2 => n24599, ZN => n2398);
   U7026 : NAND2_X1 port map( A1 => n25064, A2 => n10168, ZN => n1938);
   U7027 : NAND2_X1 port map( A1 => n9710, A2 => n1939, ZN => n8886);
   U7028 : INV_X1 port map( A => n18432, ZN => n17862);
   U7029 : OAI21_X2 port map( B1 => n2653, B2 => n16744, A => n2652, ZN => 
                           n18432);
   U7030 : OAI211_X1 port map( C1 => n10384, C2 => n11524, A => n1940, B => 
                           n11529, ZN => n2124);
   U7031 : NAND2_X1 port map( A1 => n11089, A2 => n11298, ZN => n1941);
   U7032 : XNOR2_X1 port map( A => n15251, B => n3787, ZN => n4399);
   U7033 : INV_X1 port map( A => n13264, ZN => n12932);
   U7034 : NAND3_X1 port map( A1 => n2506, A2 => n2504, A3 => n5151, ZN => 
                           n2503);
   U7036 : NAND3_X1 port map( A1 => n14171, A2 => n14165, A3 => n14164, ZN => 
                           n13734);
   U7039 : NAND2_X1 port map( A1 => n3266, A2 => n7841, ZN => n3265);
   U7040 : NAND3_X1 port map( A1 => n3058, A2 => n1945, A3 => n1944, ZN => 
                           n12276);
   U7041 : NAND2_X1 port map( A1 => n10572, A2 => n11038, ZN => n1944);
   U7042 : NAND2_X1 port map( A1 => n10513, A2 => n10571, ZN => n1945);
   U7044 : OR2_X1 port map( A1 => n13048, A2 => n12490, ZN => n2792);
   U7045 : NAND2_X1 port map( A1 => n15687, A2 => n257, ZN => n1946);
   U7046 : NAND2_X1 port map( A1 => n1948, A2 => n16235, ZN => n1947);
   U7047 : OAI21_X1 port map( B1 => n15726, B2 => n16447, A => n16239, ZN => 
                           n1948);
   U7048 : INV_X1 port map( A => n14389, ZN => n15504);
   U7049 : NAND2_X1 port map( A1 => n1950, A2 => n1949, ZN => n19801);
   U7050 : NAND2_X1 port map( A1 => n19799, A2 => n20517, ZN => n1949);
   U7051 : NAND2_X1 port map( A1 => n19797, A2 => n3522, ZN => n1950);
   U7053 : OAI211_X1 port map( C1 => n22628, C2 => n21895, A => n21897, B => 
                           n21896, ZN => n21899);
   U7054 : XOR2_X1 port map( A => n8867, B => n8446, Z => n3507);
   U7055 : AOI22_X2 port map( A1 => n9026, A2 => n9564, B1 => n9025, B2 => 
                           n9565, ZN => n10942);
   U7056 : INV_X1 port map( A => n22462, ZN => n3938);
   U7057 : NAND2_X1 port map( A1 => n1955, A2 => n1953, ZN => n20139);
   U7058 : NAND2_X1 port map( A1 => n1954, A2 => n20134, ZN => n1953);
   U7059 : NAND2_X1 port map( A1 => n4728, A2 => n20136, ZN => n1955);
   U7060 : NOR2_X2 port map( A1 => n10344, A2 => n10345, ZN => n11951);
   U7061 : NAND3_X1 port map( A1 => n1957, A2 => n1472, A3 => n1956, ZN => 
                           n16971);
   U7062 : NAND2_X1 port map( A1 => n15932, A2 => n16494, ZN => n1956);
   U7063 : NAND2_X1 port map( A1 => n15566, A2 => n16231, ZN => n1957);
   U7064 : NAND2_X1 port map( A1 => n6595, A2 => n6594, ZN => n7782);
   U7065 : NAND3_X1 port map( A1 => n21889, A2 => n5665, A3 => n22966, ZN => 
                           n5664);
   U7066 : XNOR2_X1 port map( A => n5200, B => n15033, ZN => n4723);
   U7068 : NAND2_X1 port map( A1 => n1959, A2 => n5893, ZN => n1958);
   U7069 : NAND2_X1 port map( A1 => n2007, A2 => n2006, ZN => n1960);
   U7070 : NAND3_X1 port map( A1 => n7350, A2 => n8508, A3 => n7347, ZN => 
                           n6219);
   U7071 : NAND2_X1 port map( A1 => n6695, A2 => n6699, ZN => n1962);
   U7072 : OAI22_X1 port map( A1 => n5616, A2 => n9897, B1 => n227, B2 => n9945
                           , ZN => n1963);
   U7073 : NAND3_X1 port map( A1 => n3186, A2 => n3187, A3 => n16005, ZN => 
                           n1965);
   U7074 : NAND2_X1 port map( A1 => n17463, A2 => n16846, ZN => n4198);
   U7075 : OR2_X1 port map( A1 => n16007, A2 => n16266, ZN => n1964);
   U7077 : NAND2_X1 port map( A1 => n14231, A2 => n14230, ZN => n13994);
   U7078 : NAND2_X1 port map( A1 => n13680, A2 => n24402, ZN => n1968);
   U7079 : NAND3_X1 port map( A1 => n14231, A2 => n24402, A3 => n13682, ZN => 
                           n1967);
   U7080 : NOR2_X2 port map( A1 => n13683, A2 => n13681, ZN => n14231);
   U7081 : NAND2_X1 port map( A1 => n14232, A2 => n25434, ZN => n1969);
   U7083 : NOR2_X1 port map( A1 => n7531, A2 => n1975, ZN => n3616);
   U7084 : NAND2_X1 port map( A1 => n7277, A2 => n1975, ZN => n8351);
   U7085 : AOI21_X1 port map( B1 => n3611, B2 => n1975, A => n2196, ZN => n3613
                           );
   U7086 : NAND2_X1 port map( A1 => n7747, A2 => n5738, ZN => n1973);
   U7087 : NAND2_X1 port map( A1 => n3588, A2 => n1975, ZN => n1974);
   U7088 : OAI21_X1 port map( B1 => n6672, B2 => n4754, A => n1976, ZN => n6670
                           );
   U7089 : NAND2_X1 port map( A1 => n6669, A2 => n4754, ZN => n1976);
   U7092 : OAI21_X1 port map( B1 => n18901, B2 => n18442, A => n1979, ZN => 
                           n1978);
   U7093 : NAND2_X1 port map( A1 => n18428, A2 => n25489, ZN => n18901);
   U7094 : NAND2_X1 port map( A1 => n1981, A2 => n19179, ZN => n1980);
   U7095 : NAND2_X1 port map( A1 => n1982, A2 => n19003, ZN => n1981);
   U7096 : NAND2_X1 port map( A1 => n18777, A2 => n19428, ZN => n19003);
   U7097 : NAND2_X1 port map( A1 => n16465, A2 => n16221, ZN => n3778);
   U7098 : INV_X1 port map( A => n15922, ZN => n1983);
   U7099 : NAND2_X1 port map( A1 => n1985, A2 => n7682, ZN => n7685);
   U7100 : NAND2_X1 port map( A1 => n1345, A2 => n7683, ZN => n7966);
   U7101 : NAND2_X1 port map( A1 => n270, A2 => n1985, ZN => n5684);
   U7102 : OAI21_X1 port map( B1 => n270, B2 => n1985, A => n7234, ZN => n7036)
                           ;
   U7104 : NAND2_X1 port map( A1 => n1988, A2 => n19171, ZN => n1987);
   U7105 : NAND2_X1 port map( A1 => n25469, A2 => n19412, ZN => n1990);
   U7107 : NAND2_X1 port map( A1 => n19627, A2 => n20479, ZN => n1991);
   U7108 : NAND2_X1 port map( A1 => n19628, A2 => n2168, ZN => n1993);
   U7111 : NAND2_X1 port map( A1 => n25347, A2 => n20507, ZN => n1996);
   U7112 : OAI21_X1 port map( B1 => n23320, B2 => n23311, A => n23313, ZN => 
                           n2920);
   U7113 : NAND2_X1 port map( A1 => n6274, A2 => n1509, ZN => n6028);
   U7116 : NAND2_X1 port map( A1 => n13724, A2 => n13965, ZN => n13725);
   U7117 : NAND2_X1 port map( A1 => n7771, A2 => n6126, ZN => n2004);
   U7118 : OAI21_X1 port map( B1 => n16109, B2 => n2090, A => n2089, ZN => 
                           n15592);
   U7119 : NAND3_X1 port map( A1 => n19427, A2 => n19760, A3 => n19176, ZN => 
                           n2663);
   U7120 : OR2_X1 port map( A1 => n22734, A2 => n23014, ZN => n2709);
   U7122 : INV_X1 port map( A => n14697, ZN => n14809);
   U7123 : INV_X1 port map( A => n6952, ZN => n6949);
   U7124 : OR2_X1 port map( A1 => n12447, A2 => n13165, ZN => n3442);
   U7125 : AND2_X1 port map( A1 => n7953, A2 => n7952, ZN => n7956);
   U7126 : AOI21_X1 port map( B1 => n14169, B2 => n14165, A => n14164, ZN => 
                           n4763);
   U7127 : OAI211_X1 port map( C1 => n2529, C2 => n1477, A => n2528, B => n2527
                           , ZN => n23911);
   U7128 : INV_X1 port map( A => n19163, ZN => n3727);
   U7130 : XNOR2_X1 port map( A => n21343, B => n21344, ZN => n2415);
   U7131 : INV_X1 port map( A => n17195, ZN => n4039);
   U7132 : OR2_X1 port map( A1 => n6699, A2 => n6697, ZN => n6415);
   U7133 : NAND2_X1 port map( A1 => n6699, A2 => n6556, ZN => n2006);
   U7135 : AOI21_X1 port map( B1 => n13482, B2 => n13769, A => n4331, ZN => 
                           n4330);
   U7136 : NAND2_X1 port map( A1 => n293, A2 => n16095, ZN => n16146);
   U7138 : NAND2_X1 port map( A1 => n2009, A2 => n22487, ZN => n22489);
   U7139 : NAND3_X1 port map( A1 => n22895, A2 => n2326, A3 => n2327, ZN => 
                           n2009);
   U7140 : NAND3_X1 port map( A1 => n23314, A2 => n2919, A3 => n23319, ZN => 
                           n23316);
   U7141 : OAI211_X2 port map( C1 => n20000, C2 => n20539, A => n19999, B => 
                           n2012, ZN => n3819);
   U7142 : OAI21_X1 port map( B1 => n19998, B2 => n20150, A => n20145, ZN => 
                           n2012);
   U7143 : NAND2_X1 port map( A1 => n2015, A2 => n2013, ZN => n11551);
   U7144 : NAND2_X1 port map( A1 => n12470, A2 => n11541, ZN => n2013);
   U7145 : NAND2_X1 port map( A1 => n11549, A2 => n13066, ZN => n2015);
   U7146 : NOR2_X1 port map( A1 => n13072, A2 => n12774, ZN => n11549);
   U7148 : NAND2_X1 port map( A1 => n19572, A2 => n20369, ZN => n2017);
   U7150 : OAI211_X1 port map( C1 => n2090, C2 => n16106, A => n24928, B => 
                           n2020, ZN => n15629);
   U7153 : OAI21_X1 port map( B1 => n7993, B2 => n7499, A => n7501, ZN => n7505
                           );
   U7154 : NOR2_X1 port map( A1 => n5573, A2 => n19275, ZN => n19542);
   U7157 : NAND2_X1 port map( A1 => n7457, A2 => n2022, ZN => n8498);
   U7158 : OR2_X1 port map( A1 => n7458, A2 => n7573, ZN => n2022);
   U7159 : XNOR2_X1 port map( A => n25481, B => n364, ZN => n17590);
   U7160 : NAND2_X1 port map( A1 => n10595, A2 => n1430, ZN => n10597);
   U7161 : NAND3_X1 port map( A1 => n2023, A2 => n2284, A3 => n5411, ZN => 
                           n13997);
   U7162 : OR2_X1 port map( A1 => n19908, A2 => n2024, ZN => n2568);
   U7163 : AOI21_X1 port map( B1 => n20412, B2 => n25420, A => n19741, ZN => 
                           n19908);
   U7164 : OR2_X1 port map( A1 => n413, A2 => n10518, ZN => n9291);
   U7165 : INV_X1 port map( A => n19530, ZN => n5480);
   U7168 : NAND2_X1 port map( A1 => n3407, A2 => n6324, ZN => n2025);
   U7169 : OR2_X2 port map( A1 => n6330, A2 => n6331, ZN => n9066);
   U7172 : OAI21_X1 port map( B1 => n7568, B2 => n7641, A => n7567, ZN => n2026
                           );
   U7173 : NAND2_X1 port map( A1 => n6936, A2 => n6560, ZN => n2027);
   U7174 : NAND2_X1 port map( A1 => n6697, A2 => n6699, ZN => n6936);
   U7175 : NAND2_X1 port map( A1 => n6935, A2 => n6934, ZN => n2028);
   U7178 : XNOR2_X2 port map( A => n9163, B => n9162, ZN => n10138);
   U7179 : OR2_X1 port map( A1 => n10176, A2 => n9829, ZN => n9584);
   U7180 : INV_X1 port map( A => n20039, ZN => n20185);
   U7181 : XNOR2_X1 port map( A => n9199, B => n9200, ZN => n9398);
   U7182 : NAND2_X1 port map( A1 => n2030, A2 => n9703, ZN => n9708);
   U7183 : NAND2_X1 port map( A1 => n9702, A2 => n9705, ZN => n2030);
   U7184 : NAND2_X1 port map( A1 => n3677, A2 => n4259, ZN => n3676);
   U7186 : NAND3_X1 port map( A1 => n11885, A2 => n11149, A3 => n24480, ZN => 
                           n5000);
   U7187 : AND2_X1 port map( A1 => n17048, A2 => n17050, ZN => n15956);
   U7188 : OR3_X1 port map( A1 => n25081, A2 => n22932, A3 => n24342, ZN => 
                           n21427);
   U7189 : NAND3_X1 port map( A1 => n6439, A2 => n6296, A3 => n6438, ZN => 
                           n5947);
   U7190 : NAND3_X1 port map( A1 => n3763, A2 => n6147, A3 => n6940, ZN => 
                           n5889);
   U7193 : INV_X1 port map( A => n16604, ZN => n3817);
   U7196 : NAND2_X1 port map( A1 => n2184, A2 => n10890, ZN => n2766);
   U7197 : NAND2_X1 port map( A1 => n4308, A2 => n278, ZN => n4307);
   U7198 : OAI21_X1 port map( B1 => n4442, B2 => n4441, A => n22274, ZN => 
                           n2038);
   U7199 : AOI22_X1 port map( A1 => n9498, A2 => n10090, B1 => n1348, B2 => 
                           n9497, ZN => n3088);
   U7200 : NOR2_X1 port map( A1 => n5102, A2 => n14153, ZN => n2775);
   U7202 : OAI21_X1 port map( B1 => n6088, B2 => n6372, A => n6900, ZN => n6087
                           );
   U7203 : NAND2_X1 port map( A1 => n6088, A2 => n6473, ZN => n6900);
   U7204 : NAND3_X1 port map( A1 => n6196, A2 => n6019, A3 => n6347, ZN => 
                           n6020);
   U7205 : XNOR2_X1 port map( A => n18580, B => n18581, ZN => n2041);
   U7207 : NOR2_X1 port map( A1 => n20089, A2 => n20557, ZN => n3482);
   U7208 : OAI211_X1 port map( C1 => n7292, C2 => n5202, A => n2522, B => n2043
                           , ZN => n3681);
   U7209 : NAND2_X1 port map( A1 => n5202, A2 => n432, ZN => n2043);
   U7210 : NAND2_X1 port map( A1 => n6478, A2 => n6873, ZN => n2045);
   U7211 : MUX2_X1 port map( A => n12820, B => n12821, S => n14054, Z => n12823
                           );
   U7212 : NAND2_X1 port map( A1 => n8525, A2 => n2046, ZN => n11168);
   U7213 : XNOR2_X1 port map( A => n21582, B => n20777, ZN => n3038);
   U7214 : AOI22_X2 port map( A1 => n19690, A2 => n19689, B1 => n2322, B2 => 
                           n20534, ZN => n21582);
   U7215 : NAND2_X1 port map( A1 => n19503, A2 => n358, ZN => n19504);
   U7216 : OR2_X1 port map( A1 => n1355, A2 => n14049, ZN => n12821);
   U7217 : OAI21_X1 port map( B1 => n9500, B2 => n10000, A => n9499, ZN => 
                           n10775);
   U7218 : NAND2_X1 port map( A1 => n9671, A2 => n9798, ZN => n10000);
   U7219 : AND2_X2 port map( A1 => n15969, A2 => n15968, ZN => n17572);
   U7220 : NOR2_X1 port map( A1 => n13159, A2 => n12440, ZN => n13062);
   U7221 : INV_X1 port map( A => n13837, ZN => n14271);
   U7222 : OR2_X1 port map( A1 => n24974, A2 => n13907, ZN => n13949);
   U7223 : NAND2_X1 port map( A1 => n3214, A2 => n19787, ZN => n3962);
   U7224 : INV_X1 port map( A => n9787, ZN => n4256);
   U7225 : OR2_X1 port map( A1 => n7414, A2 => n3549, ZN => n5329);
   U7226 : XNOR2_X1 port map( A => n11658, B => n2047, ZN => n10949);
   U7227 : XNOR2_X1 port map( A => n10923, B => n11942, ZN => n2047);
   U7228 : OR2_X1 port map( A1 => n13323, A2 => n2295, ZN => n12684);
   U7229 : NAND2_X1 port map( A1 => n2051, A2 => n16397, ZN => n3628);
   U7231 : INV_X1 port map( A => n25198, ZN => n13244);
   U7232 : XNOR2_X1 port map( A => n2052, B => n18176, ZN => n18180);
   U7233 : INV_X1 port map( A => n18588, ZN => n2052);
   U7234 : OAI21_X1 port map( B1 => n5704, B2 => n7329, A => n7897, ZN => n5703
                           );
   U7235 : INV_X1 port map( A => n4291, ZN => n18934);
   U7236 : XNOR2_X1 port map( A => n15219, B => n14724, ZN => n15319);
   U7237 : XNOR2_X1 port map( A => n24976, B => n2242, ZN => n14715);
   U7238 : INV_X1 port map( A => n7477, ZN => n4144);
   U7239 : INV_X1 port map( A => n20401, ZN => n5590);
   U7240 : INV_X1 port map( A => n21751, ZN => n21231);
   U7241 : OAI22_X1 port map( A1 => n3503, A2 => n3410, B1 => n5459, B2 => 
                           n16105, ZN => n15798);
   U7242 : NOR2_X1 port map( A1 => n13325, A2 => n13323, ZN => n12955);
   U7243 : INV_X1 port map( A => n14667, ZN => n3232);
   U7244 : INV_X1 port map( A => n17312, ZN => n17599);
   U7245 : XNOR2_X1 port map( A => n8119, B => n5328, ZN => n8439);
   U7246 : XNOR2_X1 port map( A => n21591, B => n4263, ZN => n20212);
   U7247 : XNOR2_X1 port map( A => n2053, B => n3901, ZN => Ciphertext(12));
   U7248 : OAI21_X1 port map( B1 => n22480, B2 => n23112, A => n22479, ZN => 
                           n2053);
   U7249 : NAND2_X1 port map( A1 => n17180, A2 => n16368, ZN => n16205);
   U7251 : OAI21_X1 port map( B1 => n17416, B2 => n17415, A => n17419, ZN => 
                           n2055);
   U7253 : OAI21_X1 port map( B1 => n7261, B2 => n7923, A => n2056, ZN => n7446
                           );
   U7254 : NAND2_X1 port map( A1 => n7923, A2 => n7932, ZN => n2056);
   U7256 : NAND2_X1 port map( A1 => n16704, A2 => n16708, ZN => n2057);
   U7257 : NAND3_X1 port map( A1 => n11884, A2 => n11145, A3 => n2059, ZN => 
                           n10535);
   U7258 : NOR2_X1 port map( A1 => n11152, A2 => n2060, ZN => n2059);
   U7264 : NAND2_X1 port map( A1 => n6522, A2 => n25398, ZN => n2061);
   U7266 : NAND2_X1 port map( A1 => n16844, A2 => n16991, ZN => n2062);
   U7267 : INV_X1 port map( A => n13260, ZN => n3791);
   U7269 : OR2_X1 port map( A1 => n25046, A2 => n10170, ZN => n9816);
   U7270 : NAND2_X1 port map( A1 => n21840, A2 => n24362, ZN => n2066);
   U7271 : NAND2_X2 port map( A1 => n19585, A2 => n2067, ZN => n20451);
   U7272 : NAND2_X1 port map( A1 => n2069, A2 => n2068, ZN => n2067);
   U7274 : INV_X1 port map( A => n14075, ZN => n14079);
   U7275 : NOR2_X1 port map( A1 => n24586, A2 => n16109, ZN => n5464);
   U7277 : NOR2_X1 port map( A1 => n15783, A2 => n379, ZN => n15590);
   U7278 : XNOR2_X1 port map( A => n2070, B => n14452, ZN => n14453);
   U7279 : XNOR2_X1 port map( A => n14451, B => n15188, ZN => n2070);
   U7281 : NAND3_X2 port map( A1 => n10002, A2 => n9800, A3 => n9801, ZN => 
                           n11499);
   U7282 : NAND3_X1 port map( A1 => n20299, A2 => n2074, A3 => n2073, ZN => 
                           n4932);
   U7283 : NAND2_X1 port map( A1 => n19979, A2 => n20298, ZN => n2073);
   U7284 : INV_X1 port map( A => n12717, ZN => n10532);
   U7285 : NAND2_X1 port map( A1 => n13169, A2 => n4766, ZN => n12717);
   U7286 : NAND2_X1 port map( A1 => n16683, A2 => n16681, ZN => n17272);
   U7287 : NAND2_X1 port map( A1 => n2076, A2 => n2075, ZN => n16683);
   U7288 : NAND2_X1 port map( A1 => n16082, A2 => n16102, ZN => n2075);
   U7289 : NAND2_X1 port map( A1 => n6122, A2 => n6245, ZN => n6989);
   U7290 : XNOR2_X1 port map( A => n25234, B => n25371, ZN => n12372);
   U7291 : NAND3_X1 port map( A1 => n10140, A2 => n10142, A3 => n10141, ZN => 
                           n10143);
   U7292 : INV_X1 port map( A => n11905, ZN => n2077);
   U7294 : NOR2_X1 port map( A1 => n10048, A2 => n10046, ZN => n2079);
   U7296 : NAND2_X1 port map( A1 => n7982, A2 => n7985, ZN => n2081);
   U7297 : NAND2_X1 port map( A1 => n4071, A2 => n23256, ZN => n2083);
   U7298 : NAND2_X1 port map( A1 => n23218, A2 => n23217, ZN => n2084);
   U7299 : NAND2_X1 port map( A1 => n21368, A2 => n20649, ZN => n4352);
   U7300 : OAI21_X1 port map( B1 => n341, B2 => n20316, A => n2913, ZN => 
                           n20323);
   U7304 : NOR2_X2 port map( A1 => n12589, A2 => n12588, ZN => n14063);
   U7305 : XNOR2_X1 port map( A => n2085, B => n8050, ZN => n8053);
   U7306 : XNOR2_X1 port map( A => n8049, B => n25407, ZN => n2085);
   U7308 : OR2_X1 port map( A1 => n7279, A2 => n7250, ZN => n2749);
   U7309 : INV_X1 port map( A => n11369, ZN => n14298);
   U7310 : INV_X1 port map( A => n23772, ZN => n23782);
   U7311 : XNOR2_X1 port map( A => n14689, B => n14815, ZN => n2969);
   U7312 : MUX2_X2 port map( A => n6701, B => n6700, S => n6934, Z => n7992);
   U7313 : XNOR2_X1 port map( A => n2088, B => n22986, ZN => Ciphertext(165));
   U7314 : NOR2_X1 port map( A1 => n22984, A2 => n22985, ZN => n2088);
   U7315 : OR2_X1 port map( A1 => n6146, A2 => n5887, ZN => n6682);
   U7316 : XNOR2_X1 port map( A => n12212, B => n12213, ZN => n12215);
   U7317 : NAND2_X1 port map( A1 => n6601, A2 => n6827, ZN => n6230);
   U7318 : NAND2_X1 port map( A1 => n16106, A2 => n16109, ZN => n2089);
   U7319 : OAI21_X1 port map( B1 => n22634, B2 => n24389, A => n21943, ZN => 
                           n21951);
   U7321 : OAI211_X1 port map( C1 => n25064, C2 => n1577, A => n24599, B => 
                           n2091, ZN => n2999);
   U7322 : NAND2_X1 port map( A1 => n4933, A2 => n4932, ZN => n19978);
   U7323 : XNOR2_X1 port map( A => n8557, B => n8826, ZN => n8441);
   U7324 : OR2_X1 port map( A1 => n5051, A2 => n7889, ZN => n2092);
   U7327 : NAND2_X1 port map( A1 => n20143, A2 => n5445, ZN => n5444);
   U7329 : NAND3_X1 port map( A1 => n3189, A2 => n4488, A3 => n17256, ZN => 
                           n17259);
   U7330 : NOR2_X1 port map( A1 => n19446, A2 => n19449, ZN => n5233);
   U7332 : INV_X1 port map( A => n6533, ZN => n4199);
   U7333 : OR2_X1 port map( A1 => n25046, A2 => n10166, ZN => n9588);
   U7334 : NAND3_X1 port map( A1 => n16813, A2 => n16814, A3 => n24410, ZN => 
                           n16816);
   U7335 : NAND2_X1 port map( A1 => n6755, A2 => n6757, ZN => n6756);
   U7336 : NOR2_X1 port map( A1 => n16186, A2 => n16397, ZN => n15828);
   U7337 : NAND3_X1 port map( A1 => n25061, A2 => n1353, A3 => n12454, ZN => 
                           n3969);
   U7338 : NAND2_X1 port map( A1 => n2625, A2 => n5570, ZN => n19743);
   U7339 : NAND2_X1 port map( A1 => n2095, A2 => n2094, ZN => n13523);
   U7340 : NAND2_X1 port map( A1 => n13520, A2 => n25247, ZN => n2094);
   U7341 : NAND2_X1 port map( A1 => n13519, A2 => n14054, ZN => n2095);
   U7343 : NAND3_X1 port map( A1 => n6753, A2 => n6754, A3 => n3276, ZN => 
                           n3274);
   U7345 : NAND2_X1 port map( A1 => n10648, A2 => n10649, ZN => n10650);
   U7346 : NAND3_X1 port map( A1 => n6408, A2 => n6412, A3 => n6409, ZN => 
                           n6411);
   U7347 : NAND2_X1 port map( A1 => n2096, A2 => n16036, ZN => n5308);
   U7349 : INV_X1 port map( A => n8436, ZN => n9001);
   U7350 : AND2_X1 port map( A1 => n13940, A2 => n16397, ZN => n16400);
   U7351 : NOR2_X1 port map( A1 => n10790, A2 => n11199, ZN => n4625);
   U7352 : OAI21_X1 port map( B1 => n24092, B2 => n10053, A => n4097, ZN => 
                           n9870);
   U7354 : NAND3_X1 port map( A1 => n15542, A2 => n15543, A3 => n15544, ZN => 
                           n15873);
   U7355 : INV_X1 port map( A => n13418, ZN => n4895);
   U7356 : NAND3_X1 port map( A1 => n2099, A2 => n13105, A3 => n12743, ZN => 
                           n12746);
   U7357 : NAND2_X1 port map( A1 => n12741, A2 => n13183, ZN => n2099);
   U7358 : NAND2_X1 port map( A1 => n3701, A2 => n13569, ZN => n3700);
   U7359 : OAI21_X1 port map( B1 => n13713, B2 => n3699, A => n3697, ZN => 
                           n13396);
   U7360 : NAND3_X1 port map( A1 => n5025, A2 => n5026, A3 => n425, ZN => n4561
                           );
   U7361 : XNOR2_X1 port map( A => n8542, B => n9044, ZN => n8543);
   U7362 : NAND2_X1 port map( A1 => n6952, A2 => n5903, ZN => n5905);
   U7363 : XNOR2_X2 port map( A => n5791, B => Key(89), ZN => n6114);
   U7364 : INV_X1 port map( A => n2546, ZN => n10497);
   U7365 : INV_X1 port map( A => n23342, ZN => n22961);
   U7366 : OR2_X1 port map( A1 => n15594, A2 => n24826, ZN => n15598);
   U7367 : INV_X1 port map( A => n16901, ZN => n2566);
   U7369 : INV_X1 port map( A => n10772, ZN => n4281);
   U7370 : NAND2_X1 port map( A1 => n2102, A2 => n2101, ZN => n6582);
   U7371 : NAND2_X1 port map( A1 => n6758, A2 => n6675, ZN => n2101);
   U7372 : NAND2_X1 port map( A1 => n5804, A2 => n6751, ZN => n2102);
   U7374 : XNOR2_X2 port map( A => n19738, B => n19737, ZN => n21848);
   U7377 : INV_X1 port map( A => n19854, ZN => n2104);
   U7379 : AND3_X2 port map( A1 => n2515, A2 => n2516, A3 => n2517, ZN => 
                           n14945);
   U7381 : NOR2_X1 port map( A1 => n16848, A2 => n17140, ZN => n2105);
   U7382 : NAND3_X1 port map( A1 => n1377, A2 => n3691, A3 => n13013, ZN => 
                           n3690);
   U7383 : NAND2_X1 port map( A1 => n4177, A2 => n6616, ZN => n6617);
   U7385 : NAND2_X1 port map( A1 => n7364, A2 => n7628, ZN => n7627);
   U7387 : OR2_X1 port map( A1 => n13124, A2 => n13350, ZN => n12873);
   U7388 : NAND3_X1 port map( A1 => n10943, A2 => n3760, A3 => n10944, ZN => 
                           n10945);
   U7389 : XNOR2_X2 port map( A => n18036, B => n18035, ZN => n19598);
   U7390 : XNOR2_X1 port map( A => n2106, B => n23657, ZN => Ciphertext(124));
   U7391 : NAND3_X1 port map( A1 => n23656, A2 => n23654, A3 => n23655, ZN => 
                           n2106);
   U7392 : NAND3_X1 port map( A1 => n11876, A2 => n11874, A3 => n11875, ZN => 
                           n13597);
   U7393 : NAND2_X1 port map( A1 => n16135, A2 => n2107, ZN => n18277);
   U7394 : NAND2_X1 port map( A1 => n17527, A2 => n17170, ZN => n2107);
   U7395 : NAND2_X1 port map( A1 => n4678, A2 => n24532, ZN => n4677);
   U7396 : OAI21_X1 port map( B1 => n8522, B2 => n9999, A => n2108, ZN => n3261
                           );
   U7397 : NAND3_X1 port map( A1 => n9310, A2 => n4137, A3 => n8521, ZN => 
                           n2108);
   U7398 : NAND2_X1 port map( A1 => n14002, A2 => n14003, ZN => n14006);
   U7400 : AOI21_X1 port map( B1 => n2109, B2 => n6030, A => n6512, ZN => n5941
                           );
   U7401 : NAND2_X1 port map( A1 => n6454, A2 => n6456, ZN => n2109);
   U7402 : NAND3_X1 port map( A1 => n3100, A2 => n10801, A3 => n10648, ZN => 
                           n10246);
   U7403 : NAND3_X1 port map( A1 => n4342, A2 => n10899, A3 => n4341, ZN => 
                           n4343);
   U7404 : OAI21_X1 port map( B1 => n2112, B2 => n285, A => n2111, ZN => n2110)
                           ;
   U7405 : INV_X1 port map( A => n4039, ZN => n2111);
   U7406 : INV_X1 port map( A => n4869, ZN => n4574);
   U7407 : XNOR2_X1 port map( A => n15398, B => n15495, ZN => n2113);
   U7408 : NAND2_X1 port map( A1 => n24532, A2 => n25030, ZN => n2478);
   U7410 : NAND2_X1 port map( A1 => n11407, A2 => n11408, ZN => n2116);
   U7411 : NAND2_X1 port map( A1 => n6734, A2 => n6730, ZN => n2118);
   U7412 : INV_X1 port map( A => n16526, ZN => n16832);
   U7413 : OR2_X1 port map( A1 => n523, A2 => n17450, ZN => n2121);
   U7414 : NAND2_X1 port map( A1 => n16979, A2 => n17450, ZN => n16526);
   U7415 : NAND3_X1 port map( A1 => n3575, A2 => n4358, A3 => n10902, ZN => 
                           n4357);
   U7417 : NOR2_X1 port map( A1 => n5315, A2 => n2246, ZN => n16904);
   U7420 : NAND3_X1 port map( A1 => n25323, A2 => n16197, A3 => n24482, ZN => 
                           n5165);
   U7421 : MUX2_X2 port map( A => n19718, B => n19717, S => n20117, Z => n21297
                           );
   U7422 : XNOR2_X2 port map( A => n8229, B => n8228, ZN => n9832);
   U7423 : AOI22_X1 port map( A1 => n17323, A2 => n4426, B1 => n15673, B2 => 
                           n17320, ZN => n17269);
   U7424 : NOR2_X1 port map( A1 => n7013, A2 => n25045, ZN => n6600);
   U7425 : AND2_X1 port map( A1 => n3358, A2 => n7948, ZN => n4812);
   U7426 : NOR2_X2 port map( A1 => n19527, A2 => n19528, ZN => n20370);
   U7427 : XNOR2_X1 port map( A => n24508, B => n14805, ZN => n3940);
   U7428 : INV_X1 port map( A => n22575, ZN => n23202);
   U7429 : OR2_X1 port map( A1 => n14205, A2 => n13549, ZN => n2214);
   U7430 : XNOR2_X1 port map( A => n14972, B => n14971, ZN => n4115);
   U7431 : OAI211_X1 port map( C1 => n24310, C2 => n19606, A => n4141, B => 
                           n19608, ZN => n2764);
   U7433 : INV_X1 port map( A => n13978, ZN => n13391);
   U7435 : NAND2_X1 port map( A1 => n2128, A2 => n2127, ZN => n7226);
   U7436 : NAND2_X1 port map( A1 => n7225, A2 => n25251, ZN => n2127);
   U7437 : NAND2_X1 port map( A1 => n3275, A2 => n7677, ZN => n2128);
   U7438 : INV_X1 port map( A => n13583, ZN => n4868);
   U7439 : MUX2_X2 port map( A => n6251, B => n6250, S => n7734, Z => n8806);
   U7440 : NAND2_X1 port map( A1 => n2130, A2 => n2129, ZN => n10546);
   U7441 : NAND2_X1 port map( A1 => n10540, A2 => n10302, ZN => n2129);
   U7442 : NAND2_X1 port map( A1 => n10539, A2 => n2389, ZN => n2130);
   U7443 : NAND3_X1 port map( A1 => n3791, A2 => n3792, A3 => n2131, ZN => 
                           n13450);
   U7444 : NAND2_X1 port map( A1 => n13257, A2 => n13974, ZN => n2131);
   U7449 : NAND4_X2 port map( A1 => n7202, A2 => n7201, A3 => n7203, A4 => 
                           n7620, ZN => n4378);
   U7450 : NOR2_X1 port map( A1 => n4812, A2 => n4093, ZN => n3359);
   U7451 : NAND2_X1 port map( A1 => n19391, A2 => n19389, ZN => n2132);
   U7452 : NAND2_X1 port map( A1 => n5710, A2 => n20474, ZN => n5711);
   U7453 : NAND2_X1 port map( A1 => n5556, A2 => n5557, ZN => n5555);
   U7454 : OR2_X1 port map( A1 => n7384, A2 => n7619, ZN => n7621);
   U7455 : NAND2_X1 port map( A1 => n17063, A2 => n24385, ZN => n2133);
   U7456 : NAND2_X1 port map( A1 => n17064, A2 => n17054, ZN => n2134);
   U7457 : NAND2_X1 port map( A1 => n4692, A2 => n19681, ZN => n2136);
   U7460 : NOR2_X1 port map( A1 => n20278, A2 => n20345, ZN => n2138);
   U7461 : NAND2_X1 port map( A1 => n6810, A2 => n2139, ZN => n8353);
   U7462 : OR2_X1 port map( A1 => n436, A2 => n8530, ZN => n2139);
   U7463 : NAND2_X1 port map( A1 => n6547, A2 => n6546, ZN => n6805);
   U7464 : NOR2_X1 port map( A1 => n9796, A2 => n9798, ZN => n2140);
   U7465 : XNOR2_X1 port map( A => n14443, B => n3695, ZN => n3694);
   U7466 : NAND2_X1 port map( A1 => n7101, A2 => n6133, ZN => n6134);
   U7467 : NAND2_X1 port map( A1 => n2388, A2 => n10302, ZN => n4327);
   U7468 : NAND3_X1 port map( A1 => n10541, A2 => n24345, A3 => n10301, ZN => 
                           n10213);
   U7469 : NAND2_X1 port map( A1 => n2142, A2 => n2141, ZN => n22386);
   U7470 : NAND2_X1 port map( A1 => n22384, A2 => n23318, ZN => n2141);
   U7471 : NAND2_X1 port map( A1 => n2143, A2 => n23317, ZN => n2142);
   U7473 : NAND3_X1 port map( A1 => n9474, A2 => n9857, A3 => n239, ZN => n9476
                           );
   U7474 : NAND3_X1 port map( A1 => n5402, A2 => n3339, A3 => n12631, ZN => 
                           n3338);
   U7475 : OAI21_X1 port map( B1 => n3404, B2 => n3401, A => n14320, ZN => 
                           n13602);
   U7476 : AOI22_X1 port map( A1 => n16354, A2 => n16980, B1 => n17453, B2 => 
                           n16979, ZN => n16370);
   U7477 : NAND2_X1 port map( A1 => n7450, A2 => n7155, ZN => n7630);
   U7478 : NAND2_X1 port map( A1 => n4439, A2 => n19597, ZN => n4438);
   U7480 : INV_X1 port map( A => n5649, ZN => n5648);
   U7481 : NAND3_X1 port map( A1 => n6636, A2 => n7021, A3 => n7027, ZN => 
                           n2146);
   U7482 : NAND2_X1 port map( A1 => n6638, A2 => n6637, ZN => n2147);
   U7483 : AND2_X1 port map( A1 => n7008, A2 => n7004, ZN => n6095);
   U7484 : NAND3_X1 port map( A1 => n15814, A2 => n16206, A3 => n3380, ZN => 
                           n15643);
   U7485 : NAND2_X1 port map( A1 => n11163, A2 => n10552, ZN => n2148);
   U7486 : NAND3_X1 port map( A1 => n9721, A2 => n9725, A3 => n10005, ZN => 
                           n9654);
   U7487 : MUX2_X1 port map( A => n15673, B => n17319, S => n17320, Z => n17325
                           );
   U7488 : NAND2_X2 port map( A1 => n2288, A2 => n2163, ZN => n17320);
   U7489 : OR2_X1 port map( A1 => n6325, A2 => n25398, ZN => n2149);
   U7490 : INV_X1 port map( A => n15893, ZN => n13374);
   U7491 : NAND2_X1 port map( A1 => n24080, A2 => n16595, ZN => n15893);
   U7493 : NAND2_X1 port map( A1 => n12467, A2 => n13521, ZN => n2150);
   U7494 : NAND2_X1 port map( A1 => n13611, A2 => n14058, ZN => n2151);
   U7495 : INV_X1 port map( A => n17686, ZN => n17689);
   U7496 : NAND2_X1 port map( A1 => n17484, A2 => n17730, ZN => n17686);
   U7497 : INV_X1 port map( A => n17414, ZN => n17224);
   U7498 : INV_X1 port map( A => n10064, ZN => n9704);
   U7499 : XNOR2_X1 port map( A => n12020, B => n12183, ZN => n11699);
   U7500 : XNOR2_X1 port map( A => n18004, B => n2964, ZN => n18005);
   U7502 : NAND3_X1 port map( A1 => n16235, A2 => n16449, A3 => n15725, ZN => 
                           n15729);
   U7503 : NAND3_X1 port map( A1 => n4198, A2 => n17461, A3 => n16021, ZN => 
                           n16993);
   U7506 : OAI21_X1 port map( B1 => n13026, B2 => n13029, A => n13025, ZN => 
                           n2153);
   U7507 : XNOR2_X1 port map( A => n18680, B => n2154, ZN => n18681);
   U7508 : XNOR2_X1 port map( A => n3703, B => n18679, ZN => n2154);
   U7509 : AND2_X1 port map( A1 => n12541, A2 => n12540, ZN => n12810);
   U7510 : NAND2_X1 port map( A1 => n2157, A2 => n2156, ZN => n10580);
   U7511 : NAND2_X1 port map( A1 => n11525, A2 => n11529, ZN => n2156);
   U7512 : NAND2_X1 port map( A1 => n1332, A2 => n11026, ZN => n2157);
   U7514 : NAND2_X1 port map( A1 => n23820, A2 => n23810, ZN => n23821);
   U7516 : NAND2_X1 port map( A1 => n6697, A2 => n6560, ZN => n5907);
   U7517 : NAND2_X1 port map( A1 => n24958, A2 => n24572, ZN => n13619);
   U7519 : NOR2_X2 port map( A1 => n8752, A2 => n2159, ZN => n11520);
   U7520 : OAI21_X1 port map( B1 => n9766, B2 => n9763, A => n8751, ZN => n2159
                           );
   U7521 : XNOR2_X1 port map( A => n9073, B => n5614, ZN => n8125);
   U7522 : XNOR2_X1 port map( A => n4025, B => n8981, ZN => n4024);
   U7523 : OR2_X1 port map( A1 => n10886, A2 => n10887, ZN => n3221);
   U7527 : XNOR2_X1 port map( A => n17660, B => n18626, ZN => n2335);
   U7528 : AND3_X2 port map( A1 => n4522, A2 => n4521, A3 => n4523, ZN => 
                           n11059);
   U7529 : OAI211_X1 port map( C1 => n9507, C2 => n9786, A => n2486, B => 
                           n24575, ZN => n4522);
   U7530 : AOI21_X2 port map( B1 => n16987, B2 => n16986, A => n2161, ZN => 
                           n18513);
   U7531 : NOR2_X1 port map( A1 => n4392, A2 => n4391, ZN => n4390);
   U7532 : XNOR2_X1 port map( A => n2162, B => n21448, ZN => n19161);
   U7533 : XNOR2_X1 port map( A => n19124, B => n21541, ZN => n2162);
   U7534 : OR2_X1 port map( A1 => n14522, A2 => n16116, ZN => n2935);
   U7535 : INV_X1 port map( A => n16246, ZN => n2605);
   U7536 : OR2_X1 port map( A1 => n15672, A2 => n15887, ZN => n2163);
   U7537 : OAI22_X1 port map( A1 => n7126, A2 => n7581, B1 => n7879, B2 => 
                           n7582, ZN => n7124);
   U7538 : NAND2_X1 port map( A1 => n10054, A2 => n10053, ZN => n10055);
   U7539 : NAND2_X1 port map( A1 => n2165, A2 => n2164, ZN => n7934);
   U7540 : OR2_X1 port map( A1 => n11023, A2 => n8934, ZN => n10920);
   U7541 : NAND2_X1 port map( A1 => n6020, A2 => n6021, ZN => n2166);
   U7542 : NAND2_X1 port map( A1 => n2167, A2 => n414, ZN => n5516);
   U7543 : NAND2_X1 port map( A1 => n2675, A2 => n11206, ZN => n2167);
   U7544 : OR2_X2 port map( A1 => n3166, A2 => n10022, ZN => n11044);
   U7545 : OAI21_X1 port map( B1 => n12534, B2 => n13048, A => n25494, ZN => 
                           n2639);
   U7547 : NAND2_X1 port map( A1 => n20194, A2 => n19744, ZN => n2169);
   U7548 : NAND2_X1 port map( A1 => n2171, A2 => n14090, ZN => n2170);
   U7549 : NAND2_X1 port map( A1 => n14088, A2 => n14089, ZN => n2171);
   U7550 : NAND2_X1 port map( A1 => n14091, A2 => n2321, ZN => n2172);
   U7551 : XNOR2_X1 port map( A => n2174, B => n22697, ZN => Ciphertext(185));
   U7552 : OAI21_X1 port map( B1 => n22696, B2 => n25076, A => n22695, ZN => 
                           n2174);
   U7554 : INV_X1 port map( A => n13228, ZN => n4587);
   U7555 : NAND3_X1 port map( A1 => n7540, A2 => n2522, A3 => n8006, ZN => 
                           n5203);
   U7556 : NAND2_X1 port map( A1 => n17252, A2 => n17272, ZN => n17282);
   U7557 : NOR2_X2 port map( A1 => n6127, A2 => n2175, ZN => n8824);
   U7559 : OR2_X2 port map( A1 => n5141, A2 => n12072, ZN => n14306);
   U7561 : INV_X1 port map( A => n13490, ZN => n3071);
   U7562 : INV_X1 port map( A => n7972, ZN => n7514);
   U7563 : INV_X1 port map( A => n18080, ZN => n3990);
   U7564 : AND3_X2 port map( A1 => n4352, A2 => n3476, A3 => n4349, ZN => 
                           n23218);
   U7565 : NAND2_X1 port map( A1 => n2177, A2 => n2176, ZN => n4801);
   U7566 : NAND2_X1 port map( A1 => n4400, A2 => n7972, ZN => n2176);
   U7568 : NAND2_X1 port map( A1 => n25360, A2 => n2178, ZN => n12702);
   U7569 : NAND2_X1 port map( A1 => n2180, A2 => n2179, ZN => n20321);
   U7571 : OAI21_X1 port map( B1 => n16869, B2 => n16870, A => n17196, ZN => 
                           n2183);
   U7572 : NOR2_X1 port map( A1 => n2185, A2 => n11084, ZN => n2184);
   U7573 : NAND3_X1 port map( A1 => n3984, A2 => n1425, A3 => n3987, ZN => 
                           n20533);
   U7574 : XNOR2_X1 port map( A => n2186, B => n21696, ZN => n18861);
   U7575 : XNOR2_X1 port map( A => n18746, B => n21247, ZN => n2186);
   U7576 : NAND2_X1 port map( A1 => n2188, A2 => n2187, ZN => n22458);
   U7577 : NAND2_X1 port map( A1 => n22456, A2 => n22455, ZN => n2187);
   U7580 : NAND2_X1 port map( A1 => n14945, A2 => n14944, ZN => n13801);
   U7581 : MUX2_X1 port map( A => n17346, B => n17345, S => n17344, Z => n17350
                           );
   U7582 : NAND2_X1 port map( A1 => n17240, A2 => n15314, ZN => n17344);
   U7583 : NAND2_X1 port map( A1 => n20039, A2 => n25478, ZN => n18729);
   U7584 : OR2_X1 port map( A1 => n16145, A2 => n16095, ZN => n2541);
   U7586 : INV_X1 port map( A => n12850, ZN => n14025);
   U7587 : NAND2_X1 port map( A1 => n6623, A2 => n316, ZN => n6621);
   U7588 : NAND4_X1 port map( A1 => n3708, A2 => n4707, A3 => n8351, A4 => 
                           n4706, ZN => n4709);
   U7589 : XNOR2_X1 port map( A => n2194, B => n21613, ZN => n22027);
   U7590 : XNOR2_X1 port map( A => n21612, B => n21611, ZN => n2194);
   U7591 : NAND3_X1 port map( A1 => n6684, A2 => n6944, A3 => n6683, ZN => 
                           n6685);
   U7592 : NAND2_X1 port map( A1 => n7582, A2 => n7313, ZN => n7583);
   U7593 : NAND2_X1 port map( A1 => n5138, A2 => n5139, ZN => n5137);
   U7594 : NAND2_X1 port map( A1 => n2195, A2 => n7598, ZN => n7259);
   U7595 : NAND2_X1 port map( A1 => n7258, A2 => n7595, ZN => n2195);
   U7596 : NAND2_X1 port map( A1 => n16122, A2 => n16123, ZN => n15846);
   U7600 : NAND3_X1 port map( A1 => n22742, A2 => n22743, A3 => n2199, ZN => 
                           n22746);
   U7604 : XNOR2_X2 port map( A => n2203, B => n3107, ZN => n10128);
   U7605 : XNOR2_X1 port map( A => n7471, B => n8703, ZN => n2203);
   U7606 : INV_X1 port map( A => n12951, ZN => n3256);
   U7607 : OAI21_X1 port map( B1 => n19084, B2 => n24584, A => n2204, ZN => 
                           n19000);
   U7608 : NAND2_X1 port map( A1 => n19084, A2 => n19418, ZN => n2204);
   U7609 : NAND3_X1 port map( A1 => n4159, A2 => n4163, A3 => n4162, ZN => 
                           n4158);
   U7610 : INV_X1 port map( A => n13167, ZN => n3688);
   U7611 : XNOR2_X1 port map( A => n2206, B => n20628, ZN => n20083);
   U7612 : XNOR2_X1 port map( A => n25202, B => n20047, ZN => n2206);
   U7613 : XNOR2_X2 port map( A => n15243, B => n15242, ZN => n16324);
   U7614 : NAND2_X1 port map( A1 => n6588, A2 => n7029, ZN => n6225);
   U7615 : NAND2_X1 port map( A1 => n6615, A2 => n6063, ZN => n2400);
   U7616 : INV_X1 port map( A => n14104, ZN => n14816);
   U7617 : OAI21_X1 port map( B1 => n22812, B2 => n22606, A => n22810, ZN => 
                           n2529);
   U7619 : OR2_X1 port map( A1 => n6296, A2 => n6297, ZN => n4865);
   U7620 : NAND3_X1 port map( A1 => n2493, A2 => n13216, A3 => n4651, ZN => 
                           n4546);
   U7621 : NAND2_X1 port map( A1 => n6722, A2 => n6243, ZN => n6721);
   U7622 : NAND2_X1 port map( A1 => n16382, A2 => n15837, ZN => n15990);
   U7623 : NAND2_X1 port map( A1 => n7107, A2 => n7250, ZN => n5928);
   U7624 : NAND2_X1 port map( A1 => n24576, A2 => n7862, ZN => n7708);
   U7625 : NAND3_X1 port map( A1 => n22330, A2 => n22329, A3 => n22464, ZN => 
                           n22331);
   U7626 : NAND2_X1 port map( A1 => n6969, A2 => n6570, ZN => n6057);
   U7627 : MUX2_X2 port map( A => n14114, B => n14113, S => n14112, Z => n15082
                           );
   U7628 : XNOR2_X2 port map( A => n8976, B => n4070, ZN => n9681);
   U7629 : OAI21_X1 port map( B1 => n5368, B2 => n2209, A => n2639, ZN => 
                           n12536);
   U7630 : NAND2_X1 port map( A1 => n4094, A2 => n13049, ZN => n2209);
   U7631 : INV_X1 port map( A => n14265, ZN => n5694);
   U7632 : INV_X1 port map( A => n8296, ZN => n2273);
   U7634 : OAI22_X1 port map( A1 => n12584, A2 => n12625, B1 => n12981, B2 => 
                           n13363, ZN => n12585);
   U7636 : XNOR2_X1 port map( A => n2210, B => n20794, ZN => n20796);
   U7637 : XNOR2_X1 port map( A => n20793, B => n21115, ZN => n2210);
   U7638 : INV_X1 port map( A => n7348, ZN => n5468);
   U7639 : OAI21_X1 port map( B1 => n20823, B2 => n23217, A => n20824, ZN => 
                           n3086);
   U7640 : OAI21_X1 port map( B1 => n4017, B2 => n20093, A => n20023, ZN => 
                           n20025);
   U7641 : INV_X1 port map( A => n14943, ZN => n2684);
   U7643 : NAND2_X1 port map( A1 => n3588, A2 => n7533, ZN => n4296);
   U7644 : OAI22_X1 port map( A1 => n21834, A2 => n3231, B1 => n21835, B2 => 
                           n21836, ZN => n3227);
   U7645 : OAI211_X1 port map( C1 => n16021, C2 => n17461, A => n3114, B => 
                           n5052, ZN => n3112);
   U7647 : NAND3_X1 port map( A1 => n15611, A2 => n15612, A3 => n16120, ZN => 
                           n2212);
   U7648 : XNOR2_X1 port map( A => n2213, B => n12025, ZN => n12026);
   U7649 : XNOR2_X1 port map( A => n12184, B => n12024, ZN => n2213);
   U7650 : NAND2_X1 port map( A1 => n2309, A2 => n10933, ZN => n2308);
   U7651 : OR2_X1 port map( A1 => n12911, A2 => n13288, ZN => n12694);
   U7652 : NAND2_X1 port map( A1 => n7961, A2 => n7683, ZN => n7684);
   U7654 : OR2_X1 port map( A1 => n16129, A2 => n16076, ZN => n14662);
   U7655 : NAND3_X2 port map( A1 => n10591, A2 => n10593, A3 => n10592, ZN => 
                           n12127);
   U7657 : XOR2_X1 port map( A => n18149, B => n3118, Z => n5327);
   U7658 : NOR2_X1 port map( A1 => n1353, A2 => n13162, ZN => n5011);
   U7659 : NAND2_X1 port map( A1 => n19098, A2 => n19367, ZN => n17801);
   U7660 : NAND2_X1 port map( A1 => n2219, A2 => n2218, ZN => n2217);
   U7661 : NAND2_X1 port map( A1 => n6350, A2 => n6271, ZN => n2219);
   U7663 : NAND2_X1 port map( A1 => n2221, A2 => n6346, ZN => n6348);
   U7664 : NAND2_X1 port map( A1 => n6345, A2 => n6445, ZN => n2221);
   U7666 : NAND2_X1 port map( A1 => n7124, A2 => n7123, ZN => n2224);
   U7667 : INV_X1 port map( A => n18796, ZN => n19281);
   U7669 : XNOR2_X1 port map( A => n14724, B => n2145, ZN => n13867);
   U7670 : NAND2_X1 port map( A1 => n2227, A2 => n2226, ZN => n12128);
   U7671 : OAI211_X1 port map( C1 => n10282, C2 => n10856, A => n10281, B => 
                           n10280, ZN => n2227);
   U7672 : NAND3_X2 port map( A1 => n20007, A2 => n5193, A3 => n20006, ZN => 
                           n22006);
   U7673 : OAI22_X1 port map( A1 => n4968, A2 => n3218, B1 => n17501, B2 => 
                           n24441, ZN => n2229);
   U7674 : NAND2_X1 port map( A1 => n10274, A2 => n10273, ZN => n11492);
   U7675 : NAND2_X1 port map( A1 => n17186, A2 => n17389, ZN => n2230);
   U7676 : NAND3_X1 port map( A1 => n2231, A2 => n18911, A3 => n1493, ZN => 
                           n20127);
   U7677 : OAI21_X1 port map( B1 => n19140, B2 => n19560, A => n25448, ZN => 
                           n2231);
   U7678 : XNOR2_X1 port map( A => n2232, B => n23489, ZN => Ciphertext(99));
   U7679 : NAND2_X1 port map( A1 => n23487, A2 => n23488, ZN => n2232);
   U7680 : NAND2_X1 port map( A1 => n12826, A2 => n12824, ZN => n12828);
   U7681 : NAND2_X1 port map( A1 => n2566, A2 => n16539, ZN => n16540);
   U7683 : NOR2_X1 port map( A1 => n5409, A2 => n16945, ZN => n2233);
   U7684 : NAND2_X1 port map( A1 => n6828, A2 => n6829, ZN => n6830);
   U7685 : NAND2_X1 port map( A1 => n18784, A2 => n18785, ZN => n18786);
   U7686 : NAND2_X1 port map( A1 => n2235, A2 => n6265, ZN => n6270);
   U7687 : NAND2_X1 port map( A1 => n6542, A2 => n7101, ZN => n2235);
   U7690 : NAND2_X1 port map( A1 => n2238, A2 => n23321, ZN => n23323);
   U7693 : NAND2_X1 port map( A1 => n6601, A2 => n5992, ZN => n6099);
   U7699 : INV_X1 port map( A => n18749, ZN => n3284);
   U7700 : NAND2_X1 port map( A1 => n6949, A2 => n25437, ZN => n5881);
   U7701 : OAI21_X1 port map( B1 => n12834, B2 => n4389, A => n13278, ZN => 
                           n4388);
   U7702 : NAND3_X1 port map( A1 => n4840, A2 => n17351, A3 => n17014, ZN => 
                           n4888);
   U7703 : OAI21_X1 port map( B1 => n10553, B2 => n1447, A => n2592, ZN => 
                           n2762);
   U7704 : XNOR2_X1 port map( A => n2242, B => n15347, ZN => n15349);
   U7705 : XNOR2_X1 port map( A => n25417, B => n2242, ZN => n14769);
   U7706 : XNOR2_X1 port map( A => n2242, B => n15514, ZN => n15517);
   U7707 : NOR2_X1 port map( A1 => n2243, A2 => n10831, ZN => n10832);
   U7708 : NAND2_X1 port map( A1 => n10275, A2 => n2243, ZN => n10515);
   U7709 : NAND2_X1 port map( A1 => n4779, A2 => n2243, ZN => n10276);
   U7710 : NAND2_X1 port map( A1 => n10834, A2 => n2243, ZN => n9647);
   U7711 : NOR2_X1 port map( A1 => n10850, A2 => n10720, ZN => n10722);
   U7712 : INV_X1 port map( A => n11123, ZN => n2244);
   U7713 : OAI211_X1 port map( C1 => n17134, C2 => n25245, A => n25226, B => 
                           n2245, ZN => n16656);
   U7714 : NAND2_X1 port map( A1 => n16655, A2 => n25245, ZN => n2245);
   U7716 : NAND2_X1 port map( A1 => n21035, A2 => n20101, ZN => n2249);
   U7720 : OAI21_X1 port map( B1 => n15588, B2 => n2253, A => n15587, ZN => 
                           n15589);
   U7721 : NAND3_X1 port map( A1 => n2255, A2 => n2256, A3 => n2254, ZN => 
                           n10623);
   U7722 : NAND3_X1 port map( A1 => n10156, A2 => n2257, A3 => n9843, ZN => 
                           n2255);
   U7724 : NAND2_X1 port map( A1 => n19370, A2 => n24968, ZN => n5461);
   U7725 : NAND2_X1 port map( A1 => n16359, A2 => n24456, ZN => n2259);
   U7726 : NAND2_X1 port map( A1 => n2262, A2 => n7676, ZN => n2261);
   U7727 : NAND3_X1 port map( A1 => n2933, A2 => n17284, A3 => n2266, ZN => 
                           n2265);
   U7728 : NAND2_X1 port map( A1 => n16950, A2 => n17293, ZN => n2266);
   U7729 : OR2_X1 port map( A1 => n2266, A2 => n17289, ZN => n2264);
   U7730 : INV_X1 port map( A => n9236, ZN => n2267);
   U7732 : NAND2_X1 port map( A1 => n9418, A2 => n9752, ZN => n2269);
   U7733 : OAI21_X1 port map( B1 => n454, B2 => n6588, A => n7031, ZN => n2270)
                           ;
   U7734 : INV_X1 port map( A => n6588, ZN => n7030);
   U7735 : XNOR2_X1 port map( A => n12240, B => n2271, ZN => n12245);
   U7736 : XNOR2_X1 port map( A => n11917, B => n2271, ZN => n11919);
   U7737 : XNOR2_X1 port map( A => n8721, B => n729, ZN => n3797);
   U7738 : XNOR2_X1 port map( A => n8721, B => n2273, ZN => n8036);
   U7739 : INV_X1 port map( A => n8721, ZN => n2274);
   U7740 : NAND2_X1 port map( A1 => n13466, A2 => n13744, ZN => n3381);
   U7741 : XNOR2_X1 port map( A => n11433, B => n12048, ZN => n2277);
   U7742 : XNOR2_X1 port map( A => n2277, B => n12342, ZN => n12348);
   U7743 : INV_X1 port map( A => n2277, ZN => n12341);
   U7744 : NAND3_X1 port map( A1 => n6926, A2 => n1175, A3 => n6291, ZN => 
                           n2279);
   U7746 : NAND2_X1 port map( A1 => n16029, A2 => n16028, ZN => n2280);
   U7747 : NAND2_X1 port map( A1 => n14927, A2 => n2281, ZN => n5336);
   U7748 : INV_X1 port map( A => n16274, ZN => n2281);
   U7749 : NAND2_X1 port map( A1 => n17467, A2 => n2064, ZN => n2282);
   U7750 : INV_X1 port map( A => n18633, ZN => n2283);
   U7751 : OR2_X1 port map( A1 => n13349, A2 => n25366, ZN => n2284);
   U7752 : AND2_X1 port map( A1 => n14231, A2 => n14235, ZN => n2977);
   U7753 : NAND3_X1 port map( A1 => n17284, A2 => n2285, A3 => n17283, ZN => 
                           n17285);
   U7754 : AOI21_X2 port map( B1 => n16755, B2 => n2285, A => n16544, ZN => 
                           n17993);
   U7755 : INV_X1 port map( A => n2285, ZN => n17287);
   U7756 : NAND2_X1 port map( A1 => n17293, A2 => n2285, ZN => n17231);
   U7757 : AND2_X1 port map( A1 => n2285, A2 => n16950, ZN => n4986);
   U7758 : NAND3_X1 port map( A1 => n2287, A2 => n16927, A3 => n17321, ZN => 
                           n3992);
   U7759 : NAND2_X1 port map( A1 => n15671, A2 => n24890, ZN => n2288);
   U7760 : NAND2_X1 port map( A1 => n2289, A2 => n12791, ZN => n2292);
   U7761 : INV_X1 port map( A => n12993, ZN => n2289);
   U7762 : NAND2_X1 port map( A1 => n2292, A2 => n2291, ZN => n2290);
   U7763 : OR2_X1 port map( A1 => n2294, A2 => n9872, ZN => n2444);
   U7764 : NAND3_X1 port map( A1 => n9872, A2 => n24549, A3 => n2294, ZN => 
                           n9547);
   U7765 : NAND2_X1 port map( A1 => n307, A2 => n2293, ZN => n9253);
   U7766 : NAND2_X1 port map( A1 => n13330, A2 => n2295, ZN => n5313);
   U7767 : AOI21_X1 port map( B1 => n13330, B2 => n25425, A => n2295, ZN => 
                           n12606);
   U7768 : NAND2_X1 port map( A1 => n21077, A2 => n22180, ZN => n2297);
   U7769 : NAND2_X1 port map( A1 => n2298, A2 => n25012, ZN => n4308);
   U7770 : NOR2_X1 port map( A1 => n19241, A2 => n2298, ZN => n18836);
   U7771 : OAI21_X1 port map( B1 => n2328, B2 => n2298, A => n278, ZN => n3055)
                           ;
   U7772 : OAI21_X1 port map( B1 => n3919, B2 => n1806, A => n2298, ZN => 
                           n18884);
   U7773 : INV_X1 port map( A => n13450, ZN => n14911);
   U7774 : XNOR2_X1 port map( A => n15093, B => n2299, ZN => n14392);
   U7775 : XNOR2_X1 port map( A => n13450, B => n2300, ZN => n2299);
   U7776 : INV_X1 port map( A => n14737, ZN => n2300);
   U7777 : NAND2_X1 port map( A1 => n13722, A2 => n13951, ZN => n2302);
   U7778 : INV_X1 port map( A => n20184, ZN => n20188);
   U7779 : NAND2_X1 port map( A1 => n19862, A2 => n25211, ZN => n20184);
   U7780 : INV_X1 port map( A => n2305, ZN => n23665);
   U7781 : NOR2_X1 port map( A1 => n24998, A2 => n23666, ZN => n5506);
   U7782 : NOR2_X1 port map( A1 => n23689, A2 => n24998, ZN => n22186);
   U7783 : NOR2_X1 port map( A1 => n23690, A2 => n24998, ZN => n23691);
   U7784 : OAI21_X1 port map( B1 => n23677, B2 => n24998, A => n23676, ZN => 
                           n23681);
   U7785 : NAND2_X1 port map( A1 => n22747, A2 => n2305, ZN => n23676);
   U7786 : NAND3_X1 port map( A1 => n25405, A2 => n23678, A3 => n24998, ZN => 
                           n22193);
   U7788 : NAND2_X1 port map( A1 => n2306, A2 => n11005, ZN => n10363);
   U7789 : NAND2_X1 port map( A1 => n10365, A2 => n2306, ZN => n10368);
   U7790 : INV_X1 port map( A => n10930, ZN => n2309);
   U7791 : NAND2_X1 port map( A1 => n5198, A2 => n10935, ZN => n5296);
   U7792 : AND2_X1 port map( A1 => n25018, A2 => n2312, ZN => n21765);
   U7793 : NAND2_X1 port map( A1 => n2315, A2 => n25018, ZN => n2314);
   U7795 : NAND2_X1 port map( A1 => n12893, A2 => n12894, ZN => n2316);
   U7796 : NAND2_X1 port map( A1 => n12895, A2 => n12896, ZN => n2317);
   U7797 : NAND2_X1 port map( A1 => n14685, A2 => n14686, ZN => n2320);
   U7798 : XNOR2_X1 port map( A => n14493, B => n2320, ZN => n11682);
   U7799 : XNOR2_X1 port map( A => n24966, B => n2318, ZN => n3695);
   U7800 : INV_X1 port map( A => n3696, ZN => n2318);
   U7801 : XNOR2_X1 port map( A => n24966, B => n2319, ZN => n14528);
   U7802 : AND2_X1 port map( A1 => n13533, A2 => n2321, ZN => n14017);
   U7805 : NAND4_X2 port map( A1 => n7190, A2 => n7189, A3 => n7188, A4 => 
                           n2323, ZN => n9059);
   U7806 : NAND2_X1 port map( A1 => n17224, A2 => n25433, ZN => n2325);
   U7807 : NAND2_X1 port map( A1 => n22893, A2 => n22717, ZN => n2327);
   U7808 : INV_X1 port map( A => n22836, ZN => n22717);
   U7809 : NAND2_X1 port map( A1 => n2330, A2 => n20571, ZN => n20619);
   U7810 : NAND2_X1 port map( A1 => n3795, A2 => n2330, ZN => n3794);
   U7811 : XNOR2_X1 port map( A => n2331, B => n2335, ZN => n2333);
   U7812 : XNOR2_X1 port map( A => n17528, B => n2334, ZN => n2331);
   U7813 : XNOR2_X1 port map( A => n17963, B => n17672, ZN => n2332);
   U7814 : NAND2_X1 port map( A1 => n2333, A2 => n19488, ZN => n18727);
   U7815 : NAND2_X1 port map( A1 => n16211, A2 => n24080, ZN => n2336);
   U7818 : NAND2_X1 port map( A1 => n5375, A2 => n2587, ZN => n2338);
   U7821 : NAND2_X1 port map( A1 => n2341, A2 => n23443, ZN => n4309);
   U7822 : NAND2_X1 port map( A1 => n2342, A2 => n22527, ZN => n2341);
   U7823 : NAND2_X1 port map( A1 => n24989, A2 => n1370, ZN => n2342);
   U7824 : INV_X1 port map( A => n23441, ZN => n22506);
   U7826 : INV_X1 port map( A => n19590, ZN => n2346);
   U7827 : NAND2_X1 port map( A1 => n18806, A2 => n2347, ZN => n18091);
   U7828 : NAND2_X1 port map( A1 => n5134, A2 => n24483, ZN => n2347);
   U7829 : INV_X1 port map( A => n5964, ZN => n2348);
   U7830 : NAND2_X1 port map( A1 => n2353, A2 => n2354, ZN => n2352);
   U7831 : NAND2_X1 port map( A1 => n2355, A2 => n1175, ZN => n2350);
   U7832 : NAND2_X1 port map( A1 => n6480, A2 => n6775, ZN => n2354);
   U7833 : NAND2_X1 port map( A1 => n2357, A2 => n20099, ZN => n2356);
   U7834 : NAND2_X1 port map( A1 => n20104, A2 => n24378, ZN => n2357);
   U7835 : NAND3_X1 port map( A1 => n15941, A2 => n25389, A3 => n2359, ZN => 
                           n15765);
   U7836 : AOI21_X1 port map( B1 => n16254, B2 => n2359, A => n16253, ZN => 
                           n16255);
   U7837 : NAND3_X1 port map( A1 => n277, A2 => n20374, A3 => n24558, ZN => 
                           n20305);
   U7839 : NOR2_X1 port map( A1 => n20591, A2 => n5093, ZN => n2361);
   U7840 : NAND2_X1 port map( A1 => n20589, A2 => n2361, ZN => n2360);
   U7841 : NAND2_X1 port map( A1 => n20591, A2 => n1424, ZN => n2363);
   U7843 : NAND2_X1 port map( A1 => n4719, A2 => n2364, ZN => n4718);
   U7844 : NAND2_X1 port map( A1 => n22497, A2 => n2364, ZN => n4720);
   U7847 : OAI21_X1 port map( B1 => n2368, B2 => n20092, A => n2367, ZN => 
                           n2365);
   U7848 : NAND2_X1 port map( A1 => n2369, A2 => n2370, ZN => n2366);
   U7849 : NAND2_X1 port map( A1 => n1455, A2 => n20092, ZN => n2367);
   U7850 : NAND2_X1 port map( A1 => n20090, A2 => n20555, ZN => n2371);
   U7852 : NAND3_X2 port map( A1 => n15776, A2 => n4956, A3 => n15775, ZN => 
                           n17078);
   U7856 : NAND2_X1 port map( A1 => n18998, A2 => n24584, ZN => n18586);
   U7857 : OAI21_X1 port map( B1 => n16509, B2 => n25376, A => n16508, ZN => 
                           n4896);
   U7858 : OAI211_X1 port map( C1 => n16509, C2 => n25376, A => n16508, B => 
                           n4899, ZN => n16510);
   U7859 : NAND2_X1 port map( A1 => n294, A2 => n25376, ZN => n4899);
   U7860 : OAI21_X1 port map( B1 => n25259, B2 => n15604, A => n25376, ZN => 
                           n15608);
   U7861 : NAND2_X1 port map( A1 => n4300, A2 => n10094, ZN => n8381);
   U7862 : NAND2_X1 port map( A1 => n9327, A2 => n4300, ZN => n5334);
   U7863 : NAND3_X1 port map( A1 => n421, A2 => n10095, A3 => n4300, ZN => 
                           n9516);
   U7865 : NOR2_X1 port map( A1 => n24043, A2 => n25471, ZN => n22591);
   U7866 : NAND2_X1 port map( A1 => n22448, A2 => n24043, ZN => n2395);
   U7867 : NAND3_X1 port map( A1 => n22448, A2 => n274, A3 => n24043, ZN => 
                           n2677);
   U7869 : NAND3_X1 port map( A1 => n2378, A2 => n2380, A3 => n2377, ZN => 
                           n2381);
   U7870 : NAND2_X1 port map( A1 => n2379, A2 => n13549, ZN => n2377);
   U7871 : NAND2_X1 port map( A1 => n14204, A2 => n3341, ZN => n2380);
   U7872 : OAI211_X1 port map( C1 => n4145, C2 => n4144, A => n2383, B => n3352
                           , ZN => n8406);
   U7873 : NAND2_X1 port map( A1 => n7477, A2 => n2384, ZN => n2383);
   U7874 : INV_X1 port map( A => n7953, ZN => n2384);
   U7876 : MUX2_X1 port map( A => n10754, B => n10755, S => n10759, Z => n10761
                           );
   U7877 : INV_X1 port map( A => n10885, ZN => n2386);
   U7878 : NOR2_X1 port map( A1 => n2388, A2 => n10302, ZN => n2387);
   U7879 : NAND2_X1 port map( A1 => n9477, A2 => n2389, ZN => n9478);
   U7880 : INV_X1 port map( A => n10302, ZN => n2389);
   U7881 : NAND2_X1 port map( A1 => n9448, A2 => n24083, ZN => n2390);
   U7883 : NAND2_X1 port map( A1 => n9447, A2 => n24054, ZN => n2392);
   U7885 : INV_X1 port map( A => n2397, ZN => n21371);
   U7886 : AOI21_X1 port map( B1 => n2397, B2 => n22792, A => n22791, ZN => 
                           n22794);
   U7887 : AND2_X1 port map( A1 => n22617, A2 => n2397, ZN => n22789);
   U7888 : NOR2_X1 port map( A1 => n2397, A2 => n22617, ZN => n22618);
   U7890 : MUX2_X1 port map( A => n22617, B => n2397, S => n22792, Z => n22474)
                           ;
   U7892 : NOR2_X1 port map( A1 => n21371, A2 => n22790, ZN => n2396);
   U7893 : NAND2_X1 port map( A1 => n22612, A2 => n2397, ZN => n4081);
   U7894 : NAND2_X1 port map( A1 => n2398, A2 => n10169, ZN => n2399);
   U7895 : NAND2_X1 port map( A1 => n2207, A2 => n10166, ZN => n2908);
   U7896 : MUX2_X1 port map( A => n9816, B => n9815, S => n2207, Z => n9819);
   U7898 : NAND2_X1 port map( A1 => n7747, A2 => n2402, ZN => n3174);
   U7900 : AND2_X1 port map( A1 => n2402, A2 => n7532, ZN => n7277);
   U7901 : NAND3_X1 port map( A1 => n3615, A2 => n2402, A3 => n8021, ZN => 
                           n4706);
   U7902 : NAND2_X1 port map( A1 => n433, A2 => n2404, ZN => n4365);
   U7903 : OAI211_X1 port map( C1 => n7697, C2 => n2404, A => n7696, B => n2403
                           , ZN => n7702);
   U7904 : NAND3_X1 port map( A1 => n7695, A2 => n1490, A3 => n2404, ZN => 
                           n2403);
   U7905 : MUX2_X1 port map( A => n2404, B => n7699, S => n7148, Z => n7152);
   U7906 : NAND3_X1 port map( A1 => n2404, A2 => n7148, A3 => n7217, ZN => 
                           n8319);
   U7908 : XNOR2_X1 port map( A => n2405, B => n11781, ZN => n11786);
   U7909 : XNOR2_X1 port map( A => n11242, B => n2406, ZN => n2405);
   U7910 : INV_X1 port map( A => n12214, ZN => n2406);
   U7911 : XNOR2_X1 port map( A => n15296, B => n14961, ZN => n2408);
   U7912 : NAND2_X1 port map( A1 => n4433, A2 => n2409, ZN => n4431);
   U7913 : INV_X1 port map( A => n19522, ZN => n2409);
   U7914 : NAND2_X1 port map( A1 => n2410, A2 => n19371, ZN => n5441);
   U7915 : OAI21_X1 port map( B1 => n19223, B2 => n2410, A => n19222, ZN => 
                           n19224);
   U7917 : OAI22_X1 port map( A1 => n23787, A2 => n2590, B1 => n2591, B2 => 
                           n2411, ZN => n2589);
   U7918 : AND2_X1 port map( A1 => n23786, A2 => n3201, ZN => n2411);
   U7919 : NAND2_X1 port map( A1 => n2412, A2 => n15198, ZN => n15767);
   U7920 : NAND2_X1 port map( A1 => n16010, A2 => n2173, ZN => n15751);
   U7921 : INV_X1 port map( A => n15556, ZN => n2412);
   U7922 : NAND2_X1 port map( A1 => n2413, A2 => n24085, ZN => n3029);
   U7923 : NAND2_X1 port map( A1 => n24802, A2 => n19480, ZN => n17894);
   U7925 : XNOR2_X1 port map( A => n21342, B => n21345, ZN => n2416);
   U7926 : NAND2_X1 port map( A1 => n2419, A2 => n2418, ZN => n17437);
   U7927 : NAND3_X1 port map( A1 => n2420, A2 => n25502, A3 => n15973, ZN => 
                           n2418);
   U7928 : NOR3_X1 port map( A1 => n21863, A2 => n23892, A3 => n23893, ZN => 
                           n23894);
   U7929 : OR2_X2 port map( A1 => n23891, A2 => n2421, ZN => n21863);
   U7930 : OAI22_X1 port map( A1 => n22772, A2 => n22370, B1 => n22682, B2 => 
                           n22679, ZN => n2421);
   U7931 : OAI211_X1 port map( C1 => n25415, C2 => n398, A => n2422, B => n5412
                           , ZN => n2424);
   U7932 : NAND2_X1 port map( A1 => n12861, A2 => n12636, ZN => n4729);
   U7933 : NAND2_X1 port map( A1 => n20460, A2 => n24460, ZN => n20165);
   U7935 : NAND2_X1 port map( A1 => n20385, A2 => n20395, ZN => n2427);
   U7937 : NAND2_X1 port map( A1 => n11302, A2 => n11297, ZN => n10434);
   U7938 : NAND2_X1 port map( A1 => n17479, A2 => n17478, ZN => n2429);
   U7939 : INV_X1 port map( A => n17078, ZN => n17479);
   U7940 : NAND2_X1 port map( A1 => n2430, A2 => n17160, ZN => n5225);
   U7941 : NAND2_X1 port map( A1 => n10538, A2 => n10885, ZN => n2435);
   U7942 : NAND2_X1 port map( A1 => n10541, A2 => n2388, ZN => n10544);
   U7943 : NAND2_X1 port map( A1 => n10888, A2 => n2388, ZN => n3417);
   U7944 : INV_X1 port map( A => n11722, ZN => n12915);
   U7945 : NAND3_X1 port map( A1 => n2437, A2 => n13304, A3 => n13307, ZN => 
                           n2436);
   U7946 : NAND2_X1 port map( A1 => n12904, A2 => n12915, ZN => n2438);
   U7947 : INV_X1 port map( A => n9872, ZN => n9251);
   U7948 : XNOR2_X2 port map( A => n8083, B => n8082, ZN => n9872);
   U7949 : NAND3_X1 port map( A1 => n2445, A2 => n2444, A3 => n2440, ZN => 
                           n10924);
   U7950 : NAND3_X1 port map( A1 => n2442, A2 => n2441, A3 => n307, ZN => n2440
                           );
   U7951 : NAND2_X1 port map( A1 => n2443, A2 => n9694, ZN => n2441);
   U7952 : NAND2_X1 port map( A1 => n9872, A2 => n9692, ZN => n2442);
   U7953 : NAND3_X1 port map( A1 => n9027, A2 => n9872, A3 => n2443, ZN => 
                           n2445);
   U7954 : INV_X1 port map( A => n9692, ZN => n2443);
   U7955 : XNOR2_X1 port map( A => n8862, B => n8086, ZN => n2446);
   U7956 : NAND3_X1 port map( A1 => n6143, A2 => n2447, A3 => n7615, ZN => 
                           n6151);
   U7957 : AND2_X1 port map( A1 => n2448, A2 => n6142, ZN => n2447);
   U7958 : OAI21_X1 port map( B1 => n10658, B2 => n10398, A => n2450, ZN => 
                           n2449);
   U7959 : NAND2_X1 port map( A1 => n25250, A2 => n10660, ZN => n10658);
   U7961 : AND2_X1 port map( A1 => n355, A2 => n19613, ZN => n18837);
   U7962 : XNOR2_X1 port map( A => n18666, B => n18491, ZN => n18538);
   U7963 : NOR2_X2 port map( A1 => n2451, A2 => n17367, ZN => n18491);
   U7964 : NAND2_X1 port map( A1 => n2452, A2 => n2453, ZN => n2451);
   U7966 : NAND2_X1 port map( A1 => n17365, A2 => n24569, ZN => n2453);
   U7970 : NAND3_X2 port map( A1 => n1390, A2 => n2887, A3 => n2456, ZN => 
                           n23592);
   U7971 : AND2_X1 port map( A1 => n24974, A2 => n14289, ZN => n2457);
   U7972 : NAND3_X1 port map( A1 => n24974, A2 => n14289, A3 => n13909, ZN => 
                           n3069);
   U7973 : OAI21_X1 port map( B1 => n13948, B2 => n2457, A => n391, ZN => 
                           n13910);
   U7974 : OAI21_X2 port map( B1 => n5622, B2 => n7911, A => n2458, ZN => n9034
                           );
   U7975 : OAI21_X1 port map( B1 => n7628, B2 => n7909, A => n2460, ZN => n2459
                           );
   U7976 : INV_X1 port map( A => n7155, ZN => n2461);
   U7978 : NAND2_X1 port map( A1 => n19107, A2 => n2464, ZN => n19584);
   U7979 : NAND2_X1 port map( A1 => n18445, A2 => n19875, ZN => n2466);
   U7980 : NAND2_X1 port map( A1 => n18444, A2 => n20023, ZN => n2467);
   U7982 : NAND2_X1 port map( A1 => n5051, A2 => n2471, ZN => n3083);
   U7983 : NOR2_X1 port map( A1 => n311, A2 => n7604, ZN => n2471);
   U7984 : INV_X1 port map( A => n12955, ZN => n2472);
   U7985 : NOR2_X1 port map( A1 => n23805, A2 => n2477, ZN => n2476);
   U7986 : NAND3_X1 port map( A1 => n4533, A2 => n21837, A3 => n2474, ZN => 
                           n2473);
   U7987 : AND2_X1 port map( A1 => n24983, A2 => n21903, ZN => n2474);
   U7989 : NAND2_X1 port map( A1 => n21837, A2 => n23002, ZN => n23787);
   U7990 : NOR2_X1 port map( A1 => n25030, A2 => n16106, ZN => n4675);
   U7991 : NAND2_X1 port map( A1 => n24928, A2 => n16107, ZN => n2479);
   U7992 : NAND2_X1 port map( A1 => n16109, A2 => n16108, ZN => n2480);
   U7993 : NAND2_X1 port map( A1 => n2484, A2 => n2482, ZN => n2481);
   U7994 : NAND2_X1 port map( A1 => n25430, A2 => n2483, ZN => n2482);
   U7995 : NOR2_X1 port map( A1 => n12349, A2 => n13350, ZN => n2483);
   U7996 : INV_X1 port map( A => n13123, ZN => n5624);
   U7997 : INV_X1 port map( A => n25430, ZN => n2485);
   U7998 : NAND2_X1 port map( A1 => n4256, A2 => n9507, ZN => n2486);
   U7999 : NAND2_X1 port map( A1 => n21954, A2 => n24911, ZN => n2488);
   U8000 : OAI22_X1 port map( A1 => n4171, A2 => n23370, B1 => n22430, B2 => 
                           n24404, ZN => n2487);
   U8001 : AOI21_X1 port map( B1 => n4606, B2 => n2488, A => n2487, ZN => n2489
                           );
   U8002 : XNOR2_X1 port map( A => n2489, B => n21711, ZN => Ciphertext(77));
   U8003 : XNOR2_X1 port map( A => n2491, B => n24413, ZN => n8445);
   U8004 : NAND2_X1 port map( A1 => n7223, A2 => n7952, ZN => n2490);
   U8005 : NAND3_X1 port map( A1 => n7953, A2 => n7952, A3 => n4144, ZN => 
                           n2880);
   U8006 : OAI21_X1 port map( B1 => n12767, B2 => n13216, A => n2492, ZN => 
                           n12811);
   U8007 : NAND2_X1 port map( A1 => n24513, A2 => n13216, ZN => n2492);
   U8008 : NAND3_X1 port map( A1 => n12987, A2 => n12986, A3 => n2493, ZN => 
                           n12988);
   U8009 : NAND2_X1 port map( A1 => n6752, A2 => n6675, ZN => n2494);
   U8010 : NAND2_X1 port map( A1 => n2497, A2 => n2501, ZN => n5101);
   U8011 : NAND2_X1 port map( A1 => n2498, A2 => n2499, ZN => n2497);
   U8012 : NAND2_X1 port map( A1 => n2500, A2 => n2499, ZN => n10838);
   U8013 : NAND2_X1 port map( A1 => n9298, A2 => n9676, ZN => n2499);
   U8014 : NAND2_X1 port map( A1 => n2501, A2 => n5448, ZN => n2500);
   U8015 : NAND3_X1 port map( A1 => n298, A2 => n14327, A3 => n5230, ZN => 
                           n2502);
   U8016 : NAND2_X1 port map( A1 => n14325, A2 => n2505, ZN => n2504);
   U8017 : INV_X1 port map( A => n13590, ZN => n2506);
   U8018 : NAND2_X1 port map( A1 => n2587, A2 => n4760, ZN => n2509);
   U8019 : NAND2_X1 port map( A1 => n2511, A2 => n17274, ZN => n2510);
   U8021 : OR2_X1 port map( A1 => n3888, A2 => n14944, ZN => n2514);
   U8023 : NAND2_X1 port map( A1 => n12621, A2 => n12622, ZN => n2517);
   U8024 : NOR2_X2 port map( A1 => n12628, A2 => n12627, ZN => n14944);
   U8025 : NAND2_X1 port map( A1 => n15857, A2 => n2518, ZN => n15805);
   U8026 : NAND2_X1 port map( A1 => n16116, A2 => n15857, ZN => n5176);
   U8028 : NAND2_X1 port map( A1 => n2520, A2 => n7757, ZN => n2521);
   U8029 : NAND2_X1 port map( A1 => n23285, A2 => n23292, ZN => n22508);
   U8030 : NAND3_X1 port map( A1 => n10698, A2 => n10952, A3 => n25232, ZN => 
                           n2523);
   U8031 : NAND3_X1 port map( A1 => n10951, A2 => n25232, A3 => n10548, ZN => 
                           n2524);
   U8032 : NAND2_X1 port map( A1 => n25038, A2 => n17330, ZN => n17331);
   U8033 : NAND2_X1 port map( A1 => n12916, A2 => n2526, ZN => n3493);
   U8034 : NAND2_X1 port map( A1 => n13311, A2 => n11722, ZN => n2526);
   U8035 : OR2_X1 port map( A1 => n13305, A2 => n12613, ZN => n13311);
   U8037 : NAND3_X1 port map( A1 => n2531, A2 => n6266, A3 => n7101, ZN => 
                           n2533);
   U8038 : INV_X1 port map( A => n7098, ZN => n2531);
   U8039 : NAND2_X1 port map( A1 => n5916, A2 => n7103, ZN => n2532);
   U8040 : NAND2_X1 port map( A1 => n6267, A2 => n6165, ZN => n6265);
   U8041 : NAND2_X1 port map( A1 => n2536, A2 => n3181, ZN => n2535);
   U8042 : NAND2_X1 port map( A1 => n2537, A2 => n23478, ZN => n2536);
   U8043 : NOR2_X1 port map( A1 => n23479, A2 => n23499, ZN => n2537);
   U8045 : INV_X1 port map( A => n2540, ZN => n19211);
   U8046 : NAND2_X1 port map( A1 => n24447, A2 => n19359, ZN => n4315);
   U8047 : NAND2_X1 port map( A1 => n19210, A2 => n24447, ZN => n19215);
   U8048 : AOI22_X1 port map( A1 => n3943, A2 => n4135, B1 => n18021, B2 => 
                           n24447, ZN => n19878);
   U8049 : OAI21_X1 port map( B1 => n6329, B2 => n6425, A => n2542, ZN => n6330
                           );
   U8051 : NAND2_X1 port map( A1 => n14036, A2 => n14035, ZN => n3893);
   U8052 : NAND2_X1 port map( A1 => n10971, A2 => n2546, ZN => n10816);
   U8053 : AND2_X2 port map( A1 => n3597, A2 => n3596, ZN => n2546);
   U8054 : NAND2_X1 port map( A1 => n2546, A2 => n10969, ZN => n10495);
   U8055 : NAND2_X1 port map( A1 => n10815, A2 => n2546, ZN => n3595);
   U8056 : XNOR2_X1 port map( A => n25483, B => n21478, ZN => n21479);
   U8059 : INV_X1 port map( A => n17438, ZN => n2549);
   U8060 : OAI21_X1 port map( B1 => n17442, B2 => n17441, A => n2550, ZN => 
                           n16829);
   U8062 : NAND2_X1 port map( A1 => n18808, A2 => n19590, ZN => n19252);
   U8064 : NAND2_X1 port map( A1 => n4286, A2 => n369, ZN => n15609);
   U8065 : NOR2_X1 port map( A1 => n7609, A2 => n7604, ZN => n7608);
   U8066 : NAND2_X1 port map( A1 => n7890, A2 => n7323, ZN => n6010);
   U8067 : NAND2_X1 port map( A1 => n7890, A2 => n2552, ZN => n2551);
   U8068 : NAND2_X1 port map( A1 => n7608, A2 => n7893, ZN => n2553);
   U8070 : NAND2_X1 port map( A1 => n7322, A2 => n7605, ZN => n2555);
   U8071 : NAND3_X1 port map( A1 => n4293, A2 => n13963, A3 => n13968, ZN => 
                           n2557);
   U8072 : INV_X1 port map( A => n14732, ZN => n15285);
   U8073 : NAND3_X1 port map( A1 => n2558, A2 => n2556, A3 => n2557, ZN => 
                           n14732);
   U8074 : NAND3_X1 port map( A1 => n2559, A2 => n1771, A3 => n4305, ZN => 
                           n2558);
   U8075 : OR2_X1 port map( A1 => n13883, A2 => n11806, ZN => n2559);
   U8076 : NAND3_X1 port map( A1 => n13968, A2 => n13724, A3 => n13969, ZN => 
                           n2556);
   U8077 : NAND2_X1 port map( A1 => n11805, A2 => n13724, ZN => n13964);
   U8078 : NAND2_X1 port map( A1 => n2558, A2 => n2557, ZN => n14397);
   U8079 : XNOR2_X1 port map( A => n8450, B => n2560, ZN => n8252);
   U8080 : XNOR2_X1 port map( A => n2560, B => n8517, ZN => n8292);
   U8081 : INV_X2 port map( A => n2562, ZN => n17633);
   U8082 : INV_X1 port map( A => n24959, ZN => n9372);
   U8083 : AOI21_X1 port map( B1 => n10252, B2 => n9378, A => n9211, ZN => 
                           n2564);
   U8084 : INV_X1 port map( A => n3472, ZN => n2565);
   U8085 : NAND3_X1 port map( A1 => n17633, A2 => n16902, A3 => n2566, ZN => 
                           n16903);
   U8086 : OR2_X1 port map( A1 => n46, A2 => n2566, ZN => n17632);
   U8087 : NAND2_X1 port map( A1 => n19742, A2 => n20255, ZN => n2567);
   U8088 : XNOR2_X1 port map( A => n2569, B => n21084, ZN => n20223);
   U8089 : XNOR2_X1 port map( A => n2569, B => n21985, ZN => n21987);
   U8090 : XNOR2_X1 port map( A => n2569, B => n21622, ZN => n19748);
   U8091 : XNOR2_X1 port map( A => n20815, B => n2569, ZN => n20817);
   U8093 : INV_X1 port map( A => n3888, ZN => n14199);
   U8094 : INV_X1 port map( A => n14949, ZN => n14950);
   U8095 : NAND2_X1 port map( A1 => n2684, A2 => n14202, ZN => n14949);
   U8096 : INV_X1 port map( A => n14945, ZN => n2570);
   U8098 : NAND2_X1 port map( A1 => n12660, A2 => n12272, ZN => n2571);
   U8099 : INV_X1 port map( A => n2572, ZN => n4921);
   U8100 : NAND2_X1 port map( A1 => n13460, A2 => n13900, ZN => n2572);
   U8101 : OAI21_X1 port map( B1 => n13733, B2 => n13460, A => n2572, ZN => 
                           n12428);
   U8102 : NAND2_X1 port map( A1 => n12499, A2 => n25033, ZN => n2574);
   U8103 : NAND2_X1 port map( A1 => n12500, A2 => n10711, ZN => n2575);
   U8104 : AND2_X1 port map( A1 => n439, A2 => n6996, ZN => n6811);
   U8105 : NAND2_X1 port map( A1 => n2576, A2 => n6658, ZN => n4149);
   U8106 : NAND3_X1 port map( A1 => n2576, A2 => n6367, A3 => n6999, ZN => 
                           n7000);
   U8107 : NAND3_X1 port map( A1 => n2576, A2 => n6658, A3 => n6367, ZN => 
                           n6074);
   U8108 : NAND2_X1 port map( A1 => n6997, A2 => n2576, ZN => n5818);
   U8109 : INV_X1 port map( A => n6996, ZN => n2576);
   U8110 : AOI21_X1 port map( B1 => n22364, B2 => n22365, A => n22675, ZN => 
                           n22368);
   U8111 : XNOR2_X1 port map( A => n4978, B => n21134, ZN => n2577);
   U8112 : INV_X1 port map( A => n18582, ZN => n17643);
   U8116 : INV_X1 port map( A => n17115, ZN => n2581);
   U8117 : OAI22_X1 port map( A1 => n10509, A2 => n2311, B1 => n10936, B2 => 
                           n2584, ZN => n10510);
   U8118 : NAND2_X1 port map( A1 => n10931, A2 => n10935, ZN => n2584);
   U8119 : NAND2_X1 port map( A1 => n10128, A2 => n2585, ZN => n10127);
   U8120 : NAND2_X1 port map( A1 => n5057, A2 => n24959, ZN => n9212);
   U8121 : NAND2_X1 port map( A1 => n10132, A2 => n24959, ZN => n9377);
   U8122 : NAND2_X1 port map( A1 => n7438, A2 => n24959, ZN => n7439);
   U8123 : MUX2_X1 port map( A => n10251, B => n10252, S => n9372, Z => n10253)
                           ;
   U8125 : AND2_X1 port map( A1 => n16796, A2 => n2587, ZN => n5762);
   U8126 : NAND2_X1 port map( A1 => n2586, A2 => n5375, ZN => n16797);
   U8127 : AND2_X1 port map( A1 => n2587, A2 => n16795, ZN => n2586);
   U8128 : MUX2_X1 port map( A => n16795, B => n2587, S => n16796, Z => n15737)
                           ;
   U8129 : NAND2_X1 port map( A1 => n5376, A2 => n2587, ZN => n2728);
   U8130 : NAND2_X1 port map( A1 => n16794, A2 => n2587, ZN => n5242);
   U8131 : INV_X1 port map( A => n22043, ZN => n23790);
   U8132 : XNOR2_X1 port map( A => n2589, B => n2588, ZN => Ciphertext(151));
   U8133 : INV_X1 port map( A => n10985, ZN => n2592);
   U8134 : AND2_X1 port map( A1 => n6713, A2 => n2593, ZN => n6717);
   U8135 : NAND2_X1 port map( A1 => n24050, A2 => n6235, ZN => n2593);
   U8136 : INV_X1 port map( A => n3480, ZN => n2594);
   U8137 : AOI21_X1 port map( B1 => n20555, B2 => n2594, A => n20330, ZN => 
                           n3478);
   U8138 : NAND2_X1 port map( A1 => n20331, A2 => n2594, ZN => n20332);
   U8139 : NAND2_X1 port map( A1 => n2596, A2 => n330, ZN => n2595);
   U8140 : NAND2_X1 port map( A1 => n22677, A2 => n23997, ZN => n2597);
   U8141 : NAND2_X1 port map( A1 => n6971, A2 => n6690, ZN => n2600);
   U8144 : NAND2_X1 port map( A1 => n6974, A2 => n2600, ZN => n4544);
   U8145 : XNOR2_X2 port map( A => n20855, B => n20854, ZN => n2601);
   U8146 : NAND2_X1 port map( A1 => n22175, A2 => n2601, ZN => n22198);
   U8147 : NOR2_X1 port map( A1 => n23571, A2 => n2601, ZN => n23572);
   U8148 : MUX2_X1 port map( A => n2601, B => n23576, S => n22175, Z => n22080)
                           ;
   U8149 : NAND2_X1 port map( A1 => n22174, A2 => n2601, ZN => n22178);
   U8150 : OAI22_X1 port map( A1 => n4360, A2 => n2601, B1 => n24369, B2 => 
                           n1323, ZN => n23577);
   U8151 : OAI22_X1 port map( A1 => n21760, A2 => n2601, B1 => n23574, B2 => 
                           n22201, ZN => n21761);
   U8152 : XNOR2_X1 port map( A => n2602, B => n2222, ZN => n11813);
   U8153 : XNOR2_X1 port map( A => n12096, B => n2602, ZN => n12098);
   U8154 : XNOR2_X1 port map( A => n12381, B => n2602, ZN => n11999);
   U8155 : XNOR2_X1 port map( A => n12241, B => n2602, ZN => n11432);
   U8156 : INV_X1 port map( A => n2603, ZN => n13587);
   U8157 : NAND2_X1 port map( A1 => n2629, A2 => n2603, ZN => n13570);
   U8160 : NAND2_X1 port map( A1 => n2607, A2 => n15564, ZN => n15565);
   U8161 : NOR2_X1 port map( A1 => n15933, A2 => n24387, ZN => n15932);
   U8162 : NAND2_X1 port map( A1 => n387, A2 => n24387, ZN => n3712);
   U8163 : NAND2_X1 port map( A1 => n5097, A2 => n24387, ZN => n5096);
   U8164 : AOI21_X1 port map( B1 => n387, B2 => n16232, A => n24387, ZN => 
                           n5024);
   U8165 : OAI21_X1 port map( B1 => n387, B2 => n2607, A => n16491, ZN => 
                           n16493);
   U8166 : OAI211_X1 port map( C1 => n24750, C2 => n25049, A => n4587, B => 
                           n2608, ZN => n12999);
   U8167 : NAND2_X1 port map( A1 => n25049, A2 => n12993, ZN => n2608);
   U8168 : OAI21_X1 port map( B1 => n15742, B2 => n16193, A => n2610, ZN => 
                           n15259);
   U8169 : NOR2_X1 port map( A1 => n16324, A2 => n25447, ZN => n15675);
   U8170 : NAND3_X1 port map( A1 => n16328, A2 => n16323, A3 => n2610, ZN => 
                           n15900);
   U8172 : MUX2_X1 port map( A => n25447, B => n16323, S => n16324, Z => n16330
                           );
   U8173 : INV_X1 port map( A => n8874, ZN => n2612);
   U8174 : XNOR2_X1 port map( A => n2611, B => n8874, ZN => n8301);
   U8175 : INV_X1 port map( A => n8457, ZN => n2611);
   U8176 : XNOR2_X1 port map( A => n2612, B => n8897, ZN => n8622);
   U8177 : NAND2_X1 port map( A1 => n372, A2 => n17053, ZN => n2615);
   U8178 : NAND3_X1 port map( A1 => n372, A2 => n17053, A3 => n2613, ZN => 
                           n2614);
   U8179 : NAND2_X1 port map( A1 => n2615, A2 => n17051, ZN => n3435);
   U8180 : NAND2_X1 port map( A1 => n330, A2 => n23998, ZN => n22376);
   U8181 : OR2_X1 port map( A1 => n2616, A2 => n24439, ZN => n24002);
   U8182 : NAND2_X1 port map( A1 => n330, A2 => n25439, ZN => n2617);
   U8184 : INV_X1 port map( A => n2621, ZN => n7791);
   U8185 : OR2_X1 port map( A1 => n2620, A2 => n7781, ZN => n2621);
   U8186 : INV_X1 port map( A => n7788, ZN => n2620);
   U8187 : NAND2_X1 port map( A1 => n7441, A2 => n2621, ZN => n7443);
   U8188 : NAND2_X1 port map( A1 => n21762, A2 => n22929, ZN => n5687);
   U8189 : NOR2_X1 port map( A1 => n22188, A2 => n22715, ZN => n21762);
   U8190 : NAND2_X1 port map( A1 => n8011, A2 => n8015, ZN => n2622);
   U8191 : INV_X1 port map( A => n8011, ZN => n2623);
   U8192 : NAND2_X1 port map( A1 => n8012, A2 => n2624, ZN => n6207);
   U8193 : NOR2_X1 port map( A1 => n2624, A2 => n7537, ZN => n7293);
   U8194 : NAND3_X1 port map( A1 => n2640, A2 => n2624, A3 => n7537, ZN => 
                           n7538);
   U8195 : NAND2_X1 port map( A1 => n8013, A2 => n2624, ZN => n3236);
   U8196 : MUX2_X1 port map( A => n8016, B => n8013, S => n2624, Z => n3238);
   U8197 : NOR2_X1 port map( A1 => n20258, A2 => n5569, ZN => n2625);
   U8198 : NAND2_X1 port map( A1 => n2627, A2 => n25054, ZN => n5570);
   U8199 : OAI21_X1 port map( B1 => n5572, B2 => n19125, A => n5571, ZN => 
                           n2627);
   U8200 : AND2_X1 port map( A1 => n15706, A2 => n16048, ZN => n15539);
   U8201 : NAND2_X1 port map( A1 => n11205, A2 => n11338, ZN => n2628);
   U8202 : NAND2_X1 port map( A1 => n2629, A2 => n14361, ZN => n13572);
   U8203 : NOR2_X1 port map( A1 => n2629, A2 => n14361, ZN => n14363);
   U8204 : NAND2_X1 port map( A1 => n13397, A2 => n1486, ZN => n15019);
   U8205 : NAND2_X1 port map( A1 => n24426, A2 => n23406, ZN => n2630);
   U8206 : NOR2_X1 port map( A1 => n24074, A2 => n23420, ZN => n23406);
   U8209 : NOR2_X1 port map( A1 => n24877, A2 => n23461, ZN => n22491);
   U8210 : XNOR2_X1 port map( A => n21725, B => n21722, ZN => n2634);
   U8211 : NAND2_X1 port map( A1 => n16441, A2 => n24293, ZN => n2635);
   U8212 : INV_X1 port map( A => n16440, ZN => n2636);
   U8214 : NAND2_X1 port map( A1 => n12536, A2 => n13757, ZN => n13837);
   U8215 : NAND3_X1 port map( A1 => n25451, A2 => n8014, A3 => n2640, ZN => 
                           n7299);
   U8216 : NAND2_X1 port map( A1 => n7293, A2 => n2640, ZN => n6214);
   U8217 : NAND3_X1 port map( A1 => n8016, A2 => n8015, A3 => n2640, ZN => 
                           n8017);
   U8218 : NAND2_X1 port map( A1 => n8011, A2 => n2640, ZN => n8020);
   U8219 : AOI21_X1 port map( B1 => n7296, B2 => n7297, A => n2640, ZN => n7301
                           );
   U8221 : NAND2_X1 port map( A1 => n17411, A2 => n17612, ZN => n2641);
   U8222 : NAND2_X1 port map( A1 => n2645, A2 => n19233, ZN => n2642);
   U8224 : INV_X1 port map( A => n19607, ZN => n2644);
   U8225 : INV_X1 port map( A => n19608, ZN => n2645);
   U8227 : NAND2_X1 port map( A1 => n6838, A2 => n6991, ZN => n2646);
   U8228 : NAND2_X1 port map( A1 => n6841, A2 => n6640, ZN => n6639);
   U8231 : NAND2_X1 port map( A1 => n15574, A2 => n16273, ZN => n2649);
   U8232 : NAND3_X1 port map( A1 => n2281, A2 => n16030, A3 => n16029, ZN => 
                           n2650);
   U8233 : NAND2_X2 port map( A1 => n14786, A2 => n3067, ZN => n17410);
   U8234 : MUX2_X1 port map( A => n17613, B => n16743, S => n17407, Z => n2652)
                           ;
   U8235 : INV_X1 port map( A => n17607, ZN => n17613);
   U8236 : NAND2_X1 port map( A1 => n17609, A2 => n17608, ZN => n2653);
   U8243 : NAND3_X1 port map( A1 => n24876, A2 => n24507, A3 => n24589, ZN => 
                           n2657);
   U8245 : NAND3_X1 port map( A1 => n5509, A2 => n5511, A3 => n2659, ZN => 
                           n17515);
   U8246 : NAND2_X1 port map( A1 => n16878, A2 => n17015, ZN => n2659);
   U8247 : INV_X1 port map( A => n22901, ZN => n5463);
   U8249 : AOI21_X1 port map( B1 => n2711, B2 => n1431, A => n2661, ZN => n2660
                           );
   U8250 : INV_X1 port map( A => n22848, ZN => n2661);
   U8251 : NAND2_X1 port map( A1 => n22904, A2 => n22842, ZN => n22848);
   U8253 : INV_X1 port map( A => n19762, ZN => n19427);
   U8254 : NOR2_X2 port map( A1 => n19761, A2 => n2662, ZN => n19953);
   U8256 : INV_X1 port map( A => n18385, ZN => n19183);
   U8258 : NAND2_X1 port map( A1 => n16724, A2 => n5484, ZN => n2664);
   U8259 : NAND2_X1 port map( A1 => n16723, A2 => n5484, ZN => n2665);
   U8260 : OR2_X1 port map( A1 => n16723, A2 => n5484, ZN => n2666);
   U8261 : XNOR2_X1 port map( A => n18456, B => n2667, ZN => n18457);
   U8262 : XNOR2_X1 port map( A => n2667, B => n18637, ZN => n18226);
   U8263 : XNOR2_X1 port map( A => n2667, B => n17663, ZN => n17533);
   U8264 : XNOR2_X1 port map( A => n2667, B => n18291, ZN => n17804);
   U8266 : NAND2_X1 port map( A1 => n2670, A2 => n23318, ZN => n2669);
   U8267 : NAND2_X1 port map( A1 => n3564, A2 => n24316, ZN => n2670);
   U8270 : XNOR2_X2 port map( A => n21529, B => n21528, ZN => n2674);
   U8271 : NAND2_X1 port map( A1 => n22421, A2 => n2674, ZN => n21547);
   U8272 : NAND2_X1 port map( A1 => n22422, A2 => n2674, ZN => n21548);
   U8274 : NOR2_X1 port map( A1 => n21530, A2 => n2674, ZN => n21531);
   U8277 : INV_X1 port map( A => n10416, ZN => n2680);
   U8278 : NAND2_X1 port map( A1 => n11012, A2 => n4531, ZN => n11010);
   U8279 : NAND2_X1 port map( A1 => n4530, A2 => n2681, ZN => n10353);
   U8280 : NAND3_X1 port map( A1 => n11045, A2 => n2680, A3 => n2681, ZN => 
                           n11049);
   U8282 : NAND2_X1 port map( A1 => n2683, A2 => n14945, ZN => n2682);
   U8286 : INV_X1 port map( A => n17192, ZN => n17028);
   U8287 : NAND2_X1 port map( A1 => n2689, A2 => n17399, ZN => n17401);
   U8288 : NAND2_X1 port map( A1 => n17398, A2 => n285, ZN => n2689);
   U8289 : AOI22_X1 port map( A1 => n3176, A2 => n23460, B1 => n2691, B2 => 
                           n23461, ZN => n2690);
   U8290 : NAND2_X1 port map( A1 => n21797, A2 => n21796, ZN => n4000);
   U8291 : OAI211_X2 port map( C1 => n24570, C2 => n4299, A => n16776, B => 
                           n4297, ZN => n18660);
   U8292 : NAND4_X2 port map( A1 => n19247, A2 => n2694, A3 => n2693, A4 => 
                           n19246, ZN => n20599);
   U8293 : NAND2_X1 port map( A1 => n2695, A2 => n19245, ZN => n2694);
   U8294 : NAND2_X1 port map( A1 => n20027, A2 => n20343, ZN => n2696);
   U8295 : NAND2_X1 port map( A1 => n19645, A2 => n20279, ZN => n2697);
   U8296 : NAND2_X1 port map( A1 => n2699, A2 => n20277, ZN => n2698);
   U8297 : AND2_X1 port map( A1 => n20346, A2 => n19809, ZN => n20027);
   U8299 : INV_X1 port map( A => n19809, ZN => n20280);
   U8300 : NAND2_X1 port map( A1 => n2702, A2 => n2703, ZN => n2701);
   U8301 : NAND2_X1 port map( A1 => n16283, A2 => n1654, ZN => n2703);
   U8302 : XNOR2_X1 port map( A => n17592, B => n16574, ZN => n2704);
   U8303 : INV_X1 port map( A => n17592, ZN => n18374);
   U8304 : XNOR2_X1 port map( A => n18284, B => n2704, ZN => n16582);
   U8307 : OAI21_X1 port map( B1 => n16185, B2 => n16337, A => n16184, ZN => 
                           n16871);
   U8308 : MUX2_X1 port map( A => n17179, B => n3602, S => n17389, Z => n17190)
                           ;
   U8311 : NAND3_X1 port map( A1 => n25382, A2 => n22900, A3 => n25569, ZN => 
                           n2708);
   U8312 : OAI21_X2 port map( B1 => n2709, B2 => n23020, A => n22735, ZN => 
                           n23480);
   U8315 : NAND2_X1 port map( A1 => n22896, A2 => n22835, ZN => n2713);
   U8316 : NOR2_X1 port map( A1 => n4737, A2 => n11163, ZN => n2714);
   U8317 : NAND3_X1 port map( A1 => n10053, A2 => n9244, A3 => n4096, ZN => 
                           n3049);
   U8319 : AOI22_X2 port map( A1 => n10437, A2 => n11092, B1 => n10436, B2 => 
                           n11300, ZN => n11646);
   U8320 : INV_X1 port map( A => n3698, ZN => n5526);
   U8321 : NOR2_X1 port map( A1 => n17031, A2 => n4039, ZN => n4038);
   U8323 : OR2_X1 port map( A1 => n6560, A2 => n6694, ZN => n6933);
   U8324 : INV_X1 port map( A => n19452, ZN => n19352);
   U8325 : INV_X1 port map( A => n23505, ZN => n23525);
   U8326 : INV_X1 port map( A => n20134, ZN => n19755);
   U8327 : INV_X1 port map( A => n3362, ZN => n7475);
   U8328 : XNOR2_X1 port map( A => n8591, B => n8590, ZN => n10006);
   U8329 : XNOR2_X1 port map( A => n8427, B => n8238, ZN => n8731);
   U8330 : OAI21_X2 port map( B1 => n16653, B2 => n16647, A => n15552, ZN => 
                           n18351);
   U8332 : OAI21_X1 port map( B1 => n9024, B2 => n9886, A => n2720, ZN => n8179
                           );
   U8333 : OAI21_X1 port map( B1 => n1376, B2 => n12768, A => n4945, ZN => 
                           n4943);
   U8334 : AOI21_X2 port map( B1 => n19405, B2 => n19404, A => n2722, ZN => 
                           n20593);
   U8335 : NAND2_X1 port map( A1 => n25064, A2 => n9814, ZN => n9512);
   U8337 : NAND3_X1 port map( A1 => n3734, A2 => n20176, A3 => n20588, ZN => 
                           n2725);
   U8338 : OAI22_X1 port map( A1 => n4270, A2 => n16268, B1 => n16004, B2 => 
                           n15758, ZN => n3709);
   U8340 : NAND2_X1 port map( A1 => n3452, A2 => n3455, ZN => n12748);
   U8341 : NAND2_X1 port map( A1 => n16146, A2 => n16145, ZN => n16152);
   U8342 : NAND2_X1 port map( A1 => n5375, A2 => n16622, ZN => n2727);
   U8344 : NAND2_X1 port map( A1 => n2732, A2 => n2731, ZN => n2730);
   U8345 : NAND2_X1 port map( A1 => n10122, A2 => n9843, ZN => n2731);
   U8346 : NAND2_X1 port map( A1 => n2868, A2 => n23236, ZN => n3124);
   U8347 : NAND2_X1 port map( A1 => n2816, A2 => n2819, ZN => n2734);
   U8349 : NAND2_X1 port map( A1 => n5087, A2 => n7022, ZN => n2736);
   U8352 : NAND2_X1 port map( A1 => n5015, A2 => n8005, ZN => n7540);
   U8353 : OAI211_X1 port map( C1 => n12582, C2 => n12844, A => n12581, B => 
                           n12845, ZN => n13427);
   U8354 : NAND2_X1 port map( A1 => n24085, A2 => n2740, ZN => n3742);
   U8355 : AND2_X1 port map( A1 => n9529, A2 => n9806, ZN => n10114);
   U8358 : NAND3_X1 port map( A1 => n7307, A2 => n7114, A3 => n6190, ZN => 
                           n6193);
   U8359 : XOR2_X1 port map( A => n12121, B => n12378, Z => n3881);
   U8360 : XNOR2_X1 port map( A => n9012, B => n8940, ZN => n2785);
   U8361 : INV_X1 port map( A => n19952, ZN => n3933);
   U8362 : NAND2_X1 port map( A1 => n2748, A2 => n3550, ZN => n7362);
   U8363 : NAND2_X1 port map( A1 => n15688, A2 => n15471, ZN => n3872);
   U8364 : NAND2_X1 port map( A1 => n6218, A2 => n7250, ZN => n2750);
   U8365 : XNOR2_X1 port map( A => n18675, B => n4711, ZN => n17716);
   U8367 : NAND3_X1 port map( A1 => n12629, A2 => n3889, A3 => n14945, ZN => 
                           n3884);
   U8368 : OAI21_X1 port map( B1 => n10369, B2 => n10365, A => n2751, ZN => 
                           n9770);
   U8370 : INV_X1 port map( A => n7043, ZN => n3729);
   U8371 : NAND2_X1 port map( A1 => n2752, A2 => n3532, ZN => n4577);
   U8373 : NAND2_X1 port map( A1 => n15790, A2 => n16042, ZN => n15266);
   U8374 : NAND3_X1 port map( A1 => n4256, A2 => n10080, A3 => n10088, ZN => 
                           n4521);
   U8377 : XNOR2_X1 port map( A => n17932, B => n17756, ZN => n17761);
   U8378 : XNOR2_X1 port map( A => n18195, B => n18276, ZN => n17756);
   U8379 : NAND2_X1 port map( A1 => n9531, A2 => n9806, ZN => n9335);
   U8381 : NAND3_X1 port map( A1 => n3192, A2 => n24861, A3 => n7899, ZN => 
                           n2759);
   U8382 : XNOR2_X1 port map( A => n17973, B => n17972, ZN => n19094);
   U8383 : INV_X1 port map( A => n13427, ZN => n13627);
   U8384 : OR2_X1 port map( A1 => n11522, A2 => n10922, ZN => n10525);
   U8385 : OAI21_X1 port map( B1 => n23138, B2 => n23143, A => n23145, ZN => 
                           n4631);
   U8386 : NAND2_X1 port map( A1 => n23138, A2 => n23154, ZN => n23145);
   U8388 : NAND2_X1 port map( A1 => n2807, A2 => n7284, ZN => n2806);
   U8389 : XNOR2_X1 port map( A => n2760, B => n20625, ZN => Ciphertext(167));
   U8390 : OR2_X1 port map( A1 => n6426, A2 => n4621, ZN => n5449);
   U8392 : NOR2_X1 port map( A1 => n16220, A2 => n16219, ZN => n16466);
   U8393 : INV_X1 port map( A => n13317, ZN => n12844);
   U8394 : OR2_X1 port map( A1 => n5434, A2 => n17069, ZN => n5462);
   U8396 : OR2_X1 port map( A1 => n13703, A2 => n14250, ZN => n13704);
   U8397 : OR2_X1 port map( A1 => n25200, A2 => n17212, ZN => n16556);
   U8398 : INV_X1 port map( A => n10846, ZN => n11124);
   U8399 : XNOR2_X1 port map( A => n18448, B => n18254, ZN => n17990);
   U8400 : AND2_X1 port map( A1 => n7268, A2 => n7843, ZN => n3266);
   U8401 : NOR2_X1 port map( A1 => n3717, A2 => n14150, ZN => n13513);
   U8402 : INV_X1 port map( A => n17012, ZN => n17353);
   U8403 : NOR2_X1 port map( A1 => n3027, A2 => n23357, ZN => n23358);
   U8404 : XNOR2_X1 port map( A => n18090, B => n18089, ZN => n19591);
   U8405 : INV_X1 port map( A => n7278, ZN => n8023);
   U8406 : INV_X1 port map( A => n16431, ZN => n17522);
   U8407 : INV_X1 port map( A => n12648, ZN => n13096);
   U8408 : NOR2_X1 port map( A1 => n23860, A2 => n24675, ZN => n4904);
   U8409 : XNOR2_X1 port map( A => n21168, B => n4455, ZN => n22449);
   U8410 : XNOR2_X1 port map( A => n8410, B => n8409, ZN => n9348);
   U8412 : NAND2_X1 port map( A1 => n10309, A2 => n11160, ZN => n2763);
   U8413 : INV_X1 port map( A => n7347, ZN => n8512);
   U8414 : NAND2_X1 port map( A1 => n13063, A2 => n24601, ZN => n13065);
   U8415 : AOI22_X2 port map( A1 => n6790, A2 => n6789, B1 => n6787, B2 => 
                           n6788, ZN => n7975);
   U8416 : NAND2_X1 port map( A1 => n11521, A2 => n3771, ZN => n3770);
   U8417 : XNOR2_X1 port map( A => n13906, B => n2765, ZN => n15167);
   U8421 : NOR2_X1 port map( A1 => n367, A2 => n17356, ZN => n2767);
   U8422 : OAI22_X1 port map( A1 => n12716, A2 => n13165, B1 => n12717, B2 => 
                           n13167, ZN => n12723);
   U8423 : NAND2_X1 port map( A1 => n12718, A2 => n4766, ZN => n12716);
   U8424 : NAND2_X1 port map( A1 => n338, A2 => n22967, ZN => n22129);
   U8425 : NAND2_X1 port map( A1 => n7319, A2 => n3300, ZN => n2768);
   U8426 : NAND2_X1 port map( A1 => n14031, A2 => n14151, ZN => n4963);
   U8428 : NAND2_X1 port map( A1 => n284, A2 => n16628, ZN => n16630);
   U8429 : NOR2_X1 port map( A1 => n24487, A2 => n5175, ZN => n5174);
   U8430 : NAND2_X1 port map( A1 => n14146, A2 => n14198, ZN => n14147);
   U8431 : NAND2_X1 port map( A1 => n15940, A2 => n16253, ZN => n2771);
   U8432 : NAND2_X1 port map( A1 => n7950, A2 => n7949, ZN => n2773);
   U8433 : NAND3_X1 port map( A1 => n10075, A2 => n10068, A3 => n10070, ZN => 
                           n2778);
   U8434 : OAI21_X1 port map( B1 => n17712, B2 => n19352, A => n2779, ZN => 
                           n17713);
   U8435 : NAND3_X1 port map( A1 => n17711, A2 => n19444, A3 => n25002, ZN => 
                           n2779);
   U8436 : NAND2_X1 port map( A1 => n16161, A2 => n16391, ZN => n15621);
   U8437 : NAND2_X1 port map( A1 => n15977, A2 => n16389, ZN => n16161);
   U8438 : XNOR2_X1 port map( A => n17816, B => n17900, ZN => n18348);
   U8439 : NAND2_X1 port map( A1 => n15792, A2 => n15791, ZN => n16575);
   U8441 : OR2_X1 port map( A1 => n12763, A2 => n11580, ZN => n11595);
   U8442 : OR2_X1 port map( A1 => n16961, A2 => n16828, ZN => n4817);
   U8443 : AND2_X1 port map( A1 => n10851, A2 => n305, ZN => n2959);
   U8444 : OR2_X1 port map( A1 => n9885, A2 => n8157, ZN => n9024);
   U8445 : AND2_X1 port map( A1 => n7023, A2 => n7021, ZN => n5087);
   U8448 : XNOR2_X1 port map( A => n17882, B => n18463, ZN => n5159);
   U8449 : XNOR2_X1 port map( A => n4024, B => n8982, ZN => n8984);
   U8450 : NAND2_X1 port map( A1 => n10524, A2 => n11529, ZN => n10526);
   U8451 : OAI21_X1 port map( B1 => n21188, B2 => n21189, A => n24043, ZN => 
                           n2781);
   U8452 : NAND2_X1 port map( A1 => n6722, A2 => n316, ZN => n6115);
   U8453 : BUF_X1 port map( A => n6208, Z => n6296);
   U8456 : OAI22_X1 port map( A1 => n9949, A2 => n9955, B1 => n9388, B2 => 
                           n9269, ZN => n9360);
   U8457 : NAND3_X1 port map( A1 => n6838, A2 => n6987, A3 => n6244, ZN => 
                           n6839);
   U8458 : NAND2_X1 port map( A1 => n4976, A2 => n7856, ZN => n4975);
   U8461 : AOI22_X1 port map( A1 => n23771, A2 => n23772, B1 => n23777, B2 => 
                           n2783, ZN => n23773);
   U8464 : INV_X1 port map( A => n17312, ZN => n2968);
   U8466 : NAND2_X1 port map( A1 => n3255, A2 => n12847, ZN => n13503);
   U8467 : NAND2_X1 port map( A1 => n5910, A2 => n6146, ZN => n6145);
   U8468 : NAND2_X1 port map( A1 => n4901, A2 => n7732, ZN => n2787);
   U8470 : OR2_X1 port map( A1 => n6970, A2 => n6969, ZN => n2788);
   U8471 : NAND2_X1 port map( A1 => n11529, A2 => n11524, ZN => n3182);
   U8473 : NAND2_X1 port map( A1 => n16240, A2 => n17216, ZN => n2789);
   U8474 : NAND2_X1 port map( A1 => n3117, A2 => n9251, ZN => n3116);
   U8475 : OAI21_X2 port map( B1 => n13749, B2 => n13748, A => n13747, ZN => 
                           n15219);
   U8476 : XNOR2_X1 port map( A => n8674, B => n8673, ZN => n8677);
   U8478 : NAND2_X1 port map( A1 => n2792, A2 => n2791, ZN => n12444);
   U8479 : NAND2_X1 port map( A1 => n13049, A2 => n12490, ZN => n2791);
   U8480 : NAND2_X1 port map( A1 => n13024, A2 => n12786, ZN => n12787);
   U8481 : NAND2_X1 port map( A1 => n2794, A2 => n2793, ZN => n12790);
   U8482 : NAND2_X1 port map( A1 => n12785, A2 => n302, ZN => n2793);
   U8485 : NOR2_X1 port map( A1 => n19558, A2 => n19555, ZN => n19140);
   U8486 : NAND2_X1 port map( A1 => n21476, A2 => n22965, ZN => n21959);
   U8489 : XNOR2_X1 port map( A => n8911, B => n8912, ZN => n9989);
   U8490 : OR2_X1 port map( A1 => n11045, A2 => n11051, ZN => n11013);
   U8491 : AND2_X1 port map( A1 => n4351, A2 => n4348, ZN => n3476);
   U8492 : INV_X1 port map( A => n19598, ZN => n19601);
   U8494 : XNOR2_X1 port map( A => n2797, B => n8570, ZN => n8571);
   U8495 : XNOR2_X1 port map( A => n8566, B => n8567, ZN => n2797);
   U8496 : NAND2_X1 port map( A1 => n10812, A2 => n5085, ZN => n3870);
   U8497 : NAND2_X1 port map( A1 => n2799, A2 => n2798, ZN => n23223);
   U8498 : NAND2_X1 port map( A1 => n23221, A2 => n24967, ZN => n2798);
   U8499 : NAND2_X1 port map( A1 => n23222, A2 => n23218, ZN => n2799);
   U8500 : OAI21_X1 port map( B1 => n6811, B2 => n6371, A => n7002, ZN => n2801
                           );
   U8501 : INV_X1 port map( A => n2803, ZN => n2802);
   U8502 : OAI22_X1 port map( A1 => n18918, A2 => n18919, B1 => n18917, B2 => 
                           n18916, ZN => n2803);
   U8503 : AOI22_X1 port map( A1 => n9761, A2 => n427, B1 => n9760, B2 => n1330
                           , ZN => n10674);
   U8504 : OAI211_X2 port map( C1 => n1551, C2 => n1423, A => n2804, B => n4841
                           , ZN => n20289);
   U8506 : OR2_X1 port map( A1 => n22945, A2 => n21531, ZN => n4170);
   U8507 : INV_X1 port map( A => n20688, ZN => n3087);
   U8508 : NOR2_X1 port map( A1 => n3615, A2 => n8021, ZN => n3614);
   U8511 : NAND2_X1 port map( A1 => n2636, A2 => n2809, ZN => n16444);
   U8513 : NAND3_X1 port map( A1 => n24103, A2 => n7896, A3 => n7897, ZN => 
                           n5901);
   U8514 : NAND2_X1 port map( A1 => n9136, A2 => n2810, ZN => n10371);
   U8517 : NAND2_X1 port map( A1 => n16500, A2 => n25572, ZN => n2811);
   U8518 : NAND3_X1 port map( A1 => n11045, A2 => n4531, A3 => n11046, ZN => 
                           n10643);
   U8520 : XNOR2_X1 port map( A => n13524, B => n15281, ZN => n2812);
   U8521 : OAI211_X1 port map( C1 => n2814, C2 => n17085, A => n17086, B => 
                           n2813, ZN => n15552);
   U8523 : INV_X1 port map( A => n17087, ZN => n2815);
   U8524 : NAND2_X1 port map( A1 => n2818, A2 => n2817, ZN => n2816);
   U8525 : INV_X1 port map( A => n22221, ZN => n2817);
   U8526 : NAND2_X1 port map( A1 => n22214, A2 => n25461, ZN => n2818);
   U8527 : NAND2_X1 port map( A1 => n21789, A2 => n22221, ZN => n2819);
   U8530 : NAND2_X1 port map( A1 => n10907, A2 => n10901, ZN => n10444);
   U8531 : INV_X1 port map( A => n13158, ZN => n12666);
   U8532 : NAND2_X1 port map( A1 => n13338, A2 => n13335, ZN => n12838);
   U8533 : NOR2_X2 port map( A1 => n16719, A2 => n2823, ZN => n18637);
   U8535 : NAND2_X1 port map( A1 => n13949, A2 => n13463, ZN => n13464);
   U8536 : NAND3_X1 port map( A1 => n2827, A2 => n22555, A3 => n22554, ZN => 
                           n22557);
   U8537 : NAND3_X1 port map( A1 => n22552, A2 => n22553, A3 => n22551, ZN => 
                           n2827);
   U8538 : AOI22_X1 port map( A1 => n15472, A2 => n17341, B1 => n17235, B2 => 
                           n16780, ZN => n2829);
   U8539 : OR2_X1 port map( A1 => n19233, A2 => n19112, ZN => n4141);
   U8541 : NAND2_X1 port map( A1 => n3985, A2 => n3986, ZN => n3984);
   U8544 : OAI21_X1 port map( B1 => n22263, B2 => n22264, A => n22262, ZN => 
                           n2833);
   U8545 : NAND3_X1 port map( A1 => n3295, A2 => n3293, A3 => n3405, ZN => 
                           n10482);
   U8546 : OAI22_X1 port map( A1 => n23660, A2 => n23686, B1 => n23662, B2 => 
                           n23661, ZN => n23664);
   U8547 : AOI21_X1 port map( B1 => n10462, B2 => n10463, A => n5077, ZN => 
                           n4501);
   U8549 : OR2_X1 port map( A1 => n10087, A2 => n10088, ZN => n2835);
   U8550 : NAND2_X1 port map( A1 => n11195, A2 => n11199, ZN => n10479);
   U8551 : INV_X1 port map( A => n7155, ZN => n7365);
   U8552 : OR2_X1 port map( A1 => n9723, A2 => n9484, ZN => n9655);
   U8553 : XNOR2_X1 port map( A => n14741, B => n14740, ZN => n5192);
   U8554 : INV_X1 port map( A => n4114, ZN => n19367);
   U8555 : INV_X1 port map( A => n14944, ZN => n12629);
   U8556 : XNOR2_X2 port map( A => n2839, B => n2838, ZN => n16106);
   U8557 : XNOR2_X1 port map( A => n15195, B => n15447, ZN => n2838);
   U8558 : XNOR2_X1 port map( A => n15156, B => n14668, ZN => n2839);
   U8560 : NAND3_X1 port map( A1 => n3515, A2 => n3516, A3 => n17013, ZN => 
                           n3514);
   U8561 : XNOR2_X1 port map( A => n3605, B => n18541, ZN => n18039);
   U8562 : INV_X1 port map( A => n15899, ZN => n15676);
   U8564 : XNOR2_X1 port map( A => n8960, B => n8244, ZN => n8436);
   U8565 : AOI21_X1 port map( B1 => n4729, B2 => n12407, A => n13347, ZN => 
                           n12421);
   U8566 : NAND2_X1 port map( A1 => n13957, A2 => n14311, ZN => n13904);
   U8569 : NAND3_X1 port map( A1 => n12935, A2 => n13235, A3 => n2842, ZN => 
                           n13238);
   U8571 : NOR2_X1 port map( A1 => n16302, A2 => n16022, ZN => n16299);
   U8572 : AOI21_X1 port map( B1 => n15917, B2 => n25092, A => n15916, ZN => 
                           n15918);
   U8573 : INV_X1 port map( A => n13903, ZN => n4525);
   U8574 : NAND3_X1 port map( A1 => n6147, A2 => n6678, A3 => n2843, ZN => 
                           n6148);
   U8575 : NAND2_X1 port map( A1 => n6679, A2 => n6281, ZN => n6147);
   U8579 : OAI21_X1 port map( B1 => n18897, B2 => n18896, A => n18895, ZN => 
                           n2844);
   U8581 : NAND2_X1 port map( A1 => n2846, A2 => n2845, ZN => n7233);
   U8582 : NAND2_X1 port map( A1 => n3469, A2 => n248, ZN => n2845);
   U8584 : OR2_X1 port map( A1 => n9753, A2 => n9613, ZN => n9750);
   U8585 : OR2_X1 port map( A1 => n4980, A2 => n14165, ZN => n4979);
   U8586 : OR2_X1 port map( A1 => n16311, A2 => n25410, ZN => n3743);
   U8588 : OAI21_X1 port map( B1 => n7648, B2 => n7651, A => n7305, ZN => n2848
                           );
   U8589 : NAND4_X2 port map( A1 => n7830, A2 => n7831, A3 => n7832, A4 => 
                           n7833, ZN => n8667);
   U8590 : NAND2_X1 port map( A1 => n16450, A2 => n223, ZN => n15929);
   U8591 : NAND3_X1 port map( A1 => n9706, A2 => n10062, A3 => n10064, ZN => 
                           n9707);
   U8592 : NAND4_X2 port map( A1 => n8017, A2 => n8020, A3 => n8018, A4 => 
                           n8019, ZN => n9169);
   U8593 : NAND2_X1 port map( A1 => n2850, A2 => n7005, ZN => n5145);
   U8594 : OAI21_X1 port map( B1 => n7011, B2 => n6650, A => n6649, ZN => n2850
                           );
   U8595 : INV_X1 port map( A => n12017, ZN => n4448);
   U8596 : XNOR2_X1 port map( A => n11753, B => n12395, ZN => n13224);
   U8597 : MUX2_X2 port map( A => n22720, B => n22719, S => n22893, Z => n23499
                           );
   U8599 : INV_X1 port map( A => n15657, ZN => n4046);
   U8601 : AOI21_X1 port map( B1 => n2851, B2 => n13313, A => n13923, ZN => 
                           n13314);
   U8602 : NAND2_X1 port map( A1 => n14253, A2 => n13924, ZN => n2851);
   U8603 : NAND2_X1 port map( A1 => n14118, A2 => n14221, ZN => n13403);
   U8604 : NAND2_X1 port map( A1 => n13399, A2 => n14219, ZN => n14118);
   U8605 : NAND3_X1 port map( A1 => n21712, A2 => n22072, A3 => n22916, ZN => 
                           n2853);
   U8606 : NOR2_X1 port map( A1 => n19973, A2 => n19974, ZN => n21534);
   U8608 : XOR2_X1 port map( A => n18666, B => n18239, Z => n4855);
   U8610 : OR2_X1 port map( A1 => n25486, A2 => n9845, ZN => n9523);
   U8611 : OR2_X1 port map( A1 => n9527, A2 => n9772, ZN => n2855);
   U8612 : OR2_X1 port map( A1 => n11806, A2 => n13968, ZN => n3425);
   U8613 : NAND2_X1 port map( A1 => n12630, A2 => n13117, ZN => n12631);
   U8614 : NAND2_X1 port map( A1 => n3607, A2 => n10325, ZN => n10330);
   U8615 : INV_X1 port map( A => n22394, ZN => n2857);
   U8616 : NAND2_X1 port map( A1 => n6121, A2 => n6642, ZN => n6124);
   U8620 : MUX2_X1 port map( A => n20353, B => n20476, S => n20480, Z => n2864)
                           ;
   U8621 : NAND2_X1 port map( A1 => n10759, A2 => n10757, ZN => n2865);
   U8622 : NAND2_X1 port map( A1 => n10758, A2 => n2867, ZN => n2866);
   U8623 : XNOR2_X1 port map( A => n11868, B => n3648, ZN => n3647);
   U8624 : NOR2_X1 port map( A1 => n23256, A2 => n2869, ZN => n2868);
   U8626 : AND2_X1 port map( A1 => n9281, A2 => n9468, ZN => n9471);
   U8628 : OAI22_X1 port map( A1 => n10512, A2 => n10570, B1 => n2870, B2 => 
                           n11038, ZN => n3058);
   U8629 : OR2_X1 port map( A1 => n9459, A2 => n9460, ZN => n9465);
   U8630 : NOR2_X1 port map( A1 => n20014, A2 => n20019, ZN => n5405);
   U8631 : NOR2_X1 port map( A1 => n9683, A2 => n9684, ZN => n8978);
   U8633 : XNOR2_X1 port map( A => n12325, B => n12144, ZN => n11388);
   U8634 : OAI21_X2 port map( B1 => n5671, B2 => n2680, A => n10645, ZN => 
                           n12144);
   U8635 : NAND3_X1 port map( A1 => n3615, A2 => n8023, A3 => n7747, ZN => 
                           n7745);
   U8637 : NAND2_X1 port map( A1 => n12670, A2 => n12671, ZN => n12677);
   U8638 : NAND2_X1 port map( A1 => n2871, A2 => n5341, ZN => n5340);
   U8639 : NAND2_X1 port map( A1 => n9391, A2 => n9953, ZN => n2871);
   U8640 : AOI22_X2 port map( A1 => n19274, A2 => n362, B1 => n2872, B2 => 
                           n19570, ZN => n20414);
   U8641 : NAND2_X1 port map( A1 => n5632, A2 => n19569, ZN => n2872);
   U8642 : NAND2_X1 port map( A1 => n7918, A2 => n7917, ZN => n8076);
   U8644 : NAND2_X1 port map( A1 => n9325, A2 => n9788, ZN => n5353);
   U8645 : INV_X1 port map( A => n14104, ZN => n4875);
   U8649 : XOR2_X1 port map( A => n21324, B => n23045, Z => n4456);
   U8650 : XNOR2_X1 port map( A => n21455, B => n21039, ZN => n21041);
   U8653 : NAND2_X1 port map( A1 => n11089, A2 => n419, ZN => n2878);
   U8654 : NAND2_X1 port map( A1 => n7957, A2 => n2880, ZN => n8770);
   U8655 : AND3_X2 port map( A1 => n5679, A2 => n11027, A3 => n11028, ZN => 
                           n12234);
   U8656 : OR2_X1 port map( A1 => n5673, A2 => n12928, ZN => n4457);
   U8657 : INV_X1 port map( A => n4899, ZN => n4898);
   U8658 : INV_X1 port map( A => n16616, ZN => n16705);
   U8659 : INV_X1 port map( A => n13224, ZN => n13009);
   U8660 : NAND2_X1 port map( A1 => n2884, A2 => n18807, ZN => n4550);
   U8661 : NAND2_X1 port map( A1 => n4551, A2 => n19250, ZN => n2884);
   U8662 : INV_X1 port map( A => n23748, ZN => n22308);
   U8664 : MUX2_X2 port map( A => n14121, B => n14120, S => n14119, Z => n15284
                           );
   U8665 : NAND2_X1 port map( A1 => n10411, A2 => n10612, ZN => n10616);
   U8666 : NAND2_X1 port map( A1 => n16285, A2 => n16342, ZN => n15679);
   U8667 : NAND2_X1 port map( A1 => n21762, A2 => n22926, ZN => n2887);
   U8668 : NAND2_X1 port map( A1 => n7769, A2 => n7771, ZN => n7770);
   U8669 : NAND2_X1 port map( A1 => n7767, A2 => n7527, ZN => n7769);
   U8670 : OAI21_X1 port map( B1 => n16923, B2 => n17320, A => n16924, ZN => 
                           n2890);
   U8672 : OAI21_X1 port map( B1 => n19335, B2 => n19496, A => n19334, ZN => 
                           n19338);
   U8673 : NAND2_X1 port map( A1 => n19335, A2 => n25459, ZN => n19334);
   U8674 : NAND2_X1 port map( A1 => n4520, A2 => n4929, ZN => n4928);
   U8675 : OR2_X1 port map( A1 => n12483, A2 => n12707, ZN => n13076);
   U8676 : INV_X1 port map( A => n2891, ZN => n3424);
   U8677 : OAI22_X1 port map( A1 => n4922, A2 => n6871, B1 => n6876, B2 => 
                           n6874, ZN => n5856);
   U8679 : NAND2_X1 port map( A1 => n23941, A2 => n23937, ZN => n23913);
   U8680 : OAI21_X1 port map( B1 => n8419, B2 => n8420, A => n8418, ZN => n2892
                           );
   U8681 : NAND3_X1 port map( A1 => n4281, A2 => n10911, A3 => n415, ZN => 
                           n9509);
   U8682 : INV_X1 port map( A => n6703, ZN => n3923);
   U8683 : NAND2_X1 port map( A1 => n2894, A2 => n7651, ZN => n2893);
   U8684 : INV_X1 port map( A => n7649, ZN => n2894);
   U8685 : NAND2_X1 port map( A1 => n2895, A2 => n10370, ZN => n10217);
   U8686 : NAND2_X1 port map( A1 => n10317, A2 => n10582, ZN => n2895);
   U8688 : NAND3_X1 port map( A1 => n4825, A2 => n7908, A3 => n7365, ZN => 
                           n2896);
   U8689 : INV_X1 port map( A => n2898, ZN => n2897);
   U8690 : OAI21_X1 port map( B1 => n7626, B2 => n7364, A => n7627, ZN => n2898
                           );
   U8691 : NAND2_X1 port map( A1 => n6393, A2 => n2900, ZN => n2899);
   U8692 : OAI211_X2 port map( C1 => n12444, C2 => n401, A => n12442, B => 
                           n12443, ZN => n14168);
   U8693 : INV_X1 port map( A => n9844, ZN => n3988);
   U8696 : XNOR2_X1 port map( A => n5304, B => n16037, ZN => n18002);
   U8697 : NAND2_X1 port map( A1 => n2902, A2 => n9064, ZN => n9689);
   U8698 : XNOR2_X2 port map( A => n9039, B => n9038, ZN => n9064);
   U8699 : INV_X1 port map( A => n10053, ZN => n2902);
   U8700 : OAI21_X1 port map( B1 => n5115, B2 => n19121, A => n5467, ZN => 
                           n5466);
   U8701 : NOR2_X1 port map( A1 => n12811, A2 => n4945, ZN => n12812);
   U8702 : AND2_X1 port map( A1 => n13839, A2 => n14267, ZN => n14276);
   U8704 : NAND2_X1 port map( A1 => n12521, A2 => n13040, ZN => n2905);
   U8705 : NAND2_X1 port map( A1 => n12522, A2 => n12478, ZN => n2906);
   U8706 : NOR2_X1 port map( A1 => n19130, A2 => n3568, ZN => n16505);
   U8707 : NAND2_X1 port map( A1 => n2908, A2 => n25, ZN => n2907);
   U8708 : NAND2_X1 port map( A1 => n9512, A2 => n10168, ZN => n2909);
   U8709 : NAND2_X1 port map( A1 => n14240, A2 => n4116, ZN => n2910);
   U8710 : NAND2_X1 port map( A1 => n13932, A2 => n13933, ZN => n2911);
   U8711 : NAND2_X1 port map( A1 => n2912, A2 => n3341, ZN => n14125);
   U8712 : NAND2_X1 port map( A1 => n14124, A2 => n14205, ZN => n2912);
   U8713 : OAI22_X1 port map( A1 => n12860, A2 => n13345, B1 => n13348, B2 => 
                           n12861, ZN => n5436);
   U8714 : XNOR2_X1 port map( A => n12410, B => n12409, ZN => n12411);
   U8715 : INV_X1 port map( A => n6072, ZN => n7002);
   U8716 : NAND2_X1 port map( A1 => n20316, A2 => n20319, ZN => n2913);
   U8718 : OR2_X1 port map( A1 => n5445, A2 => n20301, ZN => n5443);
   U8719 : INV_X1 port map( A => n4066, ZN => n19976);
   U8720 : XNOR2_X1 port map( A => n15040, B => n3462, ZN => n15332);
   U8721 : INV_X1 port map( A => n13289, ZN => n12692);
   U8722 : NAND2_X1 port map( A1 => n2914, A2 => n6893, ZN => n6897);
   U8723 : XNOR2_X2 port map( A => Key(111), B => Plaintext(111), ZN => n6987);
   U8724 : AOI21_X1 port map( B1 => n2915, B2 => n25466, A => n12910, ZN => 
                           n11803);
   U8725 : OR2_X1 port map( A1 => n13966, A2 => n13968, ZN => n3426);
   U8727 : AOI22_X1 port map( A1 => n5497, A2 => n14009, B1 => n14251, B2 => 
                           n13923, ZN => n13927);
   U8728 : NAND2_X1 port map( A1 => n17179, A2 => n17185, ZN => n16873);
   U8730 : OAI21_X1 port map( B1 => n6746, B2 => n6630, A => n6750, ZN => n6633
                           );
   U8733 : NAND2_X1 port map( A1 => n23312, A2 => n2920, ZN => n2919);
   U8734 : OR2_X1 port map( A1 => n16706, A2 => n16708, ZN => n5556);
   U8735 : XNOR2_X1 port map( A => n17899, B => n4155, ZN => n17771);
   U8736 : AOI22_X1 port map( A1 => n2923, A2 => n2922, B1 => n10012, B2 => 
                           n9724, ZN => n11172);
   U8737 : INV_X1 port map( A => n9652, ZN => n2922);
   U8738 : NAND2_X1 port map( A1 => n8609, A2 => n9725, ZN => n2923);
   U8739 : NAND3_X1 port map( A1 => n3513, A2 => n10548, A3 => n10504, ZN => 
                           n3510);
   U8740 : NOR2_X1 port map( A1 => n19499, A2 => n19498, ZN => n18721);
   U8741 : OAI21_X1 port map( B1 => n5144, B2 => n25325, A => n6503, ZN => 
                           n5142);
   U8742 : NAND3_X1 port map( A1 => n16942, A2 => n17408, A3 => n17407, ZN => 
                           n15025);
   U8743 : NAND2_X1 port map( A1 => n3690, A2 => n2924, ZN => n13907);
   U8744 : AOI22_X1 port map( A1 => n13248, A2 => n13245, B1 => n11288, B2 => 
                           n12808, ZN => n2924);
   U8745 : OAI21_X2 port map( B1 => n3041, B2 => n2925, A => n20020, ZN => 
                           n3823);
   U8746 : NAND2_X1 port map( A1 => n20015, A2 => n20016, ZN => n2925);
   U8747 : NAND2_X1 port map( A1 => n5190, A2 => n21384, ZN => n2926);
   U8748 : OAI211_X1 port map( C1 => n9928, C2 => n9600, A => n9599, B => n2928
                           , ZN => n4731);
   U8750 : XNOR2_X2 port map( A => n17586, B => n17585, ZN => n19477);
   U8751 : NAND2_X1 port map( A1 => n6944, A2 => n5909, ZN => n2930);
   U8752 : NAND2_X1 port map( A1 => n2932, A2 => n6940, ZN => n2931);
   U8753 : NAND2_X1 port map( A1 => n6679, A2 => n6146, ZN => n2932);
   U8754 : NAND2_X1 port map( A1 => n16951, A2 => n17287, ZN => n2933);
   U8755 : NAND2_X1 port map( A1 => n14521, A2 => n15804, ZN => n2934);
   U8756 : NAND2_X1 port map( A1 => n2936, A2 => n12763, ZN => n4638);
   U8757 : NAND2_X1 port map( A1 => n4640, A2 => n4639, ZN => n2936);
   U8758 : OAI21_X1 port map( B1 => n13048, B2 => n13051, A => n2940, ZN => 
                           n2939);
   U8759 : NAND2_X1 port map( A1 => n13049, A2 => n13048, ZN => n2940);
   U8760 : NAND2_X1 port map( A1 => n5368, A2 => n25408, ZN => n2941);
   U8761 : NAND2_X1 port map( A1 => n16621, A2 => n16795, ZN => n2942);
   U8762 : NAND2_X1 port map( A1 => n20225, A2 => n20269, ZN => n20229);
   U8763 : NAND2_X1 port map( A1 => n7766, A2 => n7648, ZN => n2943);
   U8764 : XNOR2_X1 port map( A => n2944, B => n8218, ZN => n9845);
   U8765 : XNOR2_X1 port map( A => n8793, B => n8217, ZN => n2944);
   U8766 : XNOR2_X1 port map( A => n5339, B => n21141, ZN => n20197);
   U8767 : XNOR2_X1 port map( A => n2945, B => n18057, ZN => n18059);
   U8768 : XNOR2_X1 port map( A => n18056, B => n25194, ZN => n2945);
   U8769 : NAND3_X1 port map( A1 => n19952, A2 => n19951, A3 => n20593, ZN => 
                           n19783);
   U8770 : AOI21_X1 port map( B1 => n19437, B2 => n19438, A => n19436, ZN => 
                           n19439);
   U8773 : NAND3_X1 port map( A1 => n6499, A2 => n6500, A3 => n6498, ZN => 
                           n6502);
   U8775 : NAND2_X1 port map( A1 => n2947, A2 => n9939, ZN => n3597);
   U8777 : NOR2_X1 port map( A1 => n12770, A2 => n12769, ZN => n12772);
   U8778 : OAI21_X2 port map( B1 => n19005, B2 => n19180, A => n19004, ZN => 
                           n20537);
   U8779 : OAI21_X1 port map( B1 => n18956, B2 => n18945, A => n3583, ZN => 
                           n3581);
   U8781 : INV_X1 port map( A => n7771, ZN => n7284);
   U8782 : OAI21_X2 port map( B1 => n10975, B2 => n10976, A => n10974, ZN => 
                           n12325);
   U8783 : NAND2_X1 port map( A1 => n9946, A2 => n9945, ZN => n9895);
   U8784 : NAND2_X1 port map( A1 => n2949, A2 => n2948, ZN => n7530);
   U8785 : NAND2_X1 port map( A1 => n7524, A2 => n23, ZN => n2948);
   U8786 : NAND2_X1 port map( A1 => n16962, A2 => n24444, ZN => n16826);
   U8788 : NAND2_X1 port map( A1 => n2952, A2 => n2951, ZN => n10209);
   U8789 : NAND2_X1 port map( A1 => n9470, A2 => n262, ZN => n2951);
   U8790 : NAND2_X1 port map( A1 => n9471, A2 => n2953, ZN => n2952);
   U8791 : INV_X1 port map( A => n9962, ZN => n2953);
   U8792 : NAND2_X1 port map( A1 => n3754, A2 => n13844, ZN => n2955);
   U8793 : NAND2_X1 port map( A1 => n24340, A2 => n10623, ZN => n10811);
   U8794 : NAND2_X1 port map( A1 => n20558, A2 => n20557, ZN => n2956);
   U8796 : OAI21_X1 port map( B1 => n13568, B2 => n13394, A => n3698, ZN => 
                           n13089);
   U8797 : XNOR2_X1 port map( A => n2957, B => n14763, ZN => n13606);
   U8798 : XNOR2_X1 port map( A => n13585, B => n14500, ZN => n2957);
   U8800 : AND2_X1 port map( A1 => n17442, A2 => n16826, ZN => n4819);
   U8802 : NAND3_X1 port map( A1 => n6216, A2 => n8511, A3 => n7351, ZN => 
                           n7251);
   U8804 : NAND2_X1 port map( A1 => n9781, A2 => n9295, ZN => n5082);
   U8805 : NAND2_X1 port map( A1 => n9222, A2 => n9223, ZN => n9224);
   U8806 : NAND2_X1 port map( A1 => n22866, A2 => n23411, ZN => n2960);
   U8807 : NAND2_X1 port map( A1 => n8370, A2 => n3979, ZN => n7266);
   U8808 : AND3_X1 port map( A1 => n6298, A2 => n4865, A3 => n6174, ZN => n6299
                           );
   U8810 : OAI22_X1 port map( A1 => n9430, A2 => n9737, B1 => n9978, B2 => 
                           n9429, ZN => n2962);
   U8811 : NOR2_X1 port map( A1 => n9431, A2 => n9982, ZN => n2963);
   U8812 : NAND2_X1 port map( A1 => n13035, A2 => n13036, ZN => n14675);
   U8813 : XNOR2_X2 port map( A => n14899, B => n5331, ZN => n16029);
   U8814 : NAND2_X1 port map( A1 => n24310, A2 => n4884, ZN => n4140);
   U8815 : NAND2_X1 port map( A1 => n9563, A2 => n9564, ZN => n9570);
   U8817 : INV_X1 port map( A => n17339, ZN => n5104);
   U8818 : OR2_X1 port map( A1 => n5910, A2 => n6146, ZN => n6945);
   U8819 : XNOR2_X2 port map( A => Key(189), B => Plaintext(189), ZN => n6445);
   U8820 : NAND2_X1 port map( A1 => n16404, A2 => n16403, ZN => n3765);
   U8822 : NAND2_X2 port map( A1 => n6865, A2 => n2965, ZN => n8987);
   U8823 : MUX2_X1 port map( A => n4951, B => n10729, S => n10728, Z => n11189)
                           ;
   U8825 : NAND2_X1 port map( A1 => n2966, A2 => n13284, ZN => n13286);
   U8826 : NAND2_X1 port map( A1 => n13283, A2 => n13282, ZN => n2966);
   U8828 : NAND3_X1 port map( A1 => n19942, A2 => n20450, A3 => n20377, ZN => 
                           n19943);
   U8829 : OAI21_X1 port map( B1 => n2613, B2 => n17048, A => n17049, ZN => 
                           n16774);
   U8830 : AOI21_X2 port map( B1 => n15954, B2 => n15955, A => n16482, ZN => 
                           n17049);
   U8832 : NAND2_X1 port map( A1 => n24506, A2 => n16226, ZN => n16298);
   U8833 : INV_X1 port map( A => n10839, ZN => n4464);
   U8835 : NAND2_X1 port map( A1 => n3499, A2 => n7580, ZN => n3498);
   U8836 : NAND2_X1 port map( A1 => n4631, A2 => n4630, ZN => n4628);
   U8838 : INV_X1 port map( A => n7992, ZN => n3549);
   U8839 : NOR2_X1 port map( A1 => n5594, A2 => n7733, ZN => n5593);
   U8840 : NAND2_X1 port map( A1 => n15533, A2 => n15534, ZN => n16742);
   U8841 : INV_X1 port map( A => n10518, ZN => n4013);
   U8842 : NAND2_X1 port map( A1 => n9938, A2 => n9905, ZN => n2971);
   U8843 : NAND3_X1 port map( A1 => n1485, A2 => n6618, A3 => n7419, ZN => 
                           n2972);
   U8844 : INV_X1 port map( A => n5349, ZN => n23449);
   U8845 : XNOR2_X2 port map( A => n20287, B => n20288, ZN => n22656);
   U8847 : OAI21_X2 port map( B1 => n12837, B2 => n12966, A => n12836, ZN => 
                           n14333);
   U8848 : NAND2_X1 port map( A1 => n6612, A2 => n24501, ZN => n2973);
   U8849 : NAND3_X1 port map( A1 => n6611, A2 => n6718, A3 => n6610, ZN => 
                           n2974);
   U8850 : OR2_X1 port map( A1 => n11867, A2 => n11873, ZN => n11876);
   U8852 : NAND3_X2 port map( A1 => n17097, A2 => n17095, A3 => n17096, ZN => 
                           n18356);
   U8853 : OR2_X1 port map( A1 => n13210, A2 => n5418, ZN => n3039);
   U8854 : INV_X1 port map( A => n18902, ZN => n19539);
   U8855 : XOR2_X1 port map( A => n18671, B => n18083, Z => n5135);
   U8857 : INV_X1 port map( A => n3720, ZN => n23245);
   U8858 : NOR2_X1 port map( A1 => n22279, A2 => n22280, ZN => n22944);
   U8859 : INV_X1 port map( A => n20094, ZN => n4017);
   U8860 : INV_X1 port map( A => n11101, ZN => n4143);
   U8861 : INV_X1 port map( A => n20519, ZN => n19925);
   U8862 : XNOR2_X1 port map( A => n5343, B => n7161, ZN => n8997);
   U8863 : NAND2_X1 port map( A1 => n19372, A2 => n19376, ZN => n19373);
   U8864 : AOI22_X1 port map( A1 => n14232, A2 => n14234, B1 => n2977, B2 => 
                           n13680, ZN => n14238);
   U8865 : MUX2_X1 port map( A => n4418, B => n24249, S => n15625, Z => n14745)
                           ;
   U8866 : XNOR2_X2 port map( A => n14572, B => n14573, ZN => n15625);
   U8868 : NAND2_X1 port map( A1 => n18889, A2 => n25057, ZN => n19403);
   U8869 : NAND2_X1 port map( A1 => n22661, A2 => n25160, ZN => n2978);
   U8871 : INV_X1 port map( A => n13929, ZN => n4837);
   U8872 : NAND2_X1 port map( A1 => n3926, A2 => n6956, ZN => n4323);
   U8873 : NAND2_X1 port map( A1 => n25078, A2 => n25375, ZN => n22095);
   U8874 : NAND2_X1 port map( A1 => n4322, A2 => n6960, ZN => n4321);
   U8875 : XNOR2_X1 port map( A => n2979, B => n14978, ZN => n14985);
   U8876 : XNOR2_X1 port map( A => n14981, B => n15342, ZN => n2979);
   U8877 : NAND2_X1 port map( A1 => n13118, A2 => n13117, ZN => n2980);
   U8879 : OR2_X1 port map( A1 => n1355, A2 => n14048, ZN => n13612);
   U8880 : AOI21_X2 port map( B1 => n16479, B2 => n16478, A => n16477, ZN => 
                           n16851);
   U8881 : NAND2_X1 port map( A1 => n23554, A2 => n24057, ZN => n23544);
   U8883 : INV_X1 port map( A => n18196, ZN => n4666);
   U8884 : INV_X1 port map( A => n12868, ZN => n3328);
   U8888 : NOR2_X1 port map( A1 => n23766, A2 => n2982, ZN => n23774);
   U8889 : NAND2_X1 port map( A1 => n4917, A2 => n19269, ZN => n2983);
   U8890 : INV_X1 port map( A => n4737, ZN => n2984);
   U8891 : NOR2_X1 port map( A1 => n25031, A2 => n17054, ZN => n16721);
   U8894 : NAND2_X1 port map( A1 => n2988, A2 => n2985, ZN => n19626);
   U8895 : NAND2_X1 port map( A1 => n2987, A2 => n2986, ZN => n2985);
   U8896 : NOR2_X1 port map( A1 => n22252, A2 => n21841, ZN => n2986);
   U8897 : NAND2_X1 port map( A1 => n19343, A2 => n22252, ZN => n2988);
   U8901 : INV_X1 port map( A => n13568, ZN => n3701);
   U8902 : NAND2_X1 port map( A1 => n19764, A2 => n20591, ZN => n19766);
   U8903 : OAI22_X1 port map( A1 => n11023, A2 => n11520, B1 => n11024, B2 => 
                           n11529, ZN => n11025);
   U8904 : NAND2_X1 port map( A1 => n11024, A2 => n11519, ZN => n11023);
   U8905 : INV_X1 port map( A => n7077, ZN => n4375);
   U8906 : XNOR2_X2 port map( A => n11774, B => n11775, ZN => n13291);
   U8907 : NAND2_X1 port map( A1 => n2993, A2 => n13790, ZN => n13791);
   U8908 : NAND2_X1 port map( A1 => n14140, A2 => n14141, ZN => n2993);
   U8909 : OAI22_X1 port map( A1 => n9229, A2 => n9709, B1 => n9711, B2 => 
                           n10039, ZN => n2994);
   U8910 : INV_X1 port map( A => n5249, ZN => n6788);
   U8911 : OAI21_X1 port map( B1 => n2996, B2 => n24459, A => n2995, ZN => 
                           n15844);
   U8912 : NAND2_X1 port map( A1 => n24459, A2 => n16125, ZN => n2995);
   U8913 : NAND3_X1 port map( A1 => n127, A2 => n6165, A3 => n6543, ZN => n6042
                           );
   U8914 : NOR2_X1 port map( A1 => n10502, A2 => n13167, ZN => n10531);
   U8916 : INV_X1 port map( A => n8012, ZN => n8016);
   U8917 : NAND2_X1 port map( A1 => n7002, A2 => n6815, ZN => n5819);
   U8919 : NAND2_X1 port map( A1 => n2999, A2 => n2998, ZN => n10174);
   U8920 : NAND2_X1 port map( A1 => n10171, A2 => n25046, ZN => n2998);
   U8923 : NAND2_X1 port map( A1 => n10702, A2 => n25074, ZN => n10704);
   U8924 : OR2_X1 port map( A1 => n24446, A2 => n9244, ZN => n9688);
   U8927 : NAND2_X1 port map( A1 => n16781, A2 => n17347, ZN => n3002);
   U8928 : NAND2_X1 port map( A1 => n17000, A2 => n16999, ZN => n3005);
   U8929 : NAND3_X1 port map( A1 => n4863, A2 => n22149, A3 => n4864, ZN => 
                           n4862);
   U8931 : NAND2_X1 port map( A1 => n7599, A2 => n7598, ZN => n3006);
   U8934 : NAND2_X1 port map( A1 => n15981, A2 => n16167, ZN => n3009);
   U8935 : NAND3_X1 port map( A1 => n24576, A2 => n7861, A3 => n3570, ZN => 
                           n7872);
   U8936 : XNOR2_X1 port map( A => n18687, B => n5304, ZN => n5303);
   U8937 : NAND2_X1 port map( A1 => n17179, A2 => n16871, ZN => n16872);
   U8938 : NAND2_X1 port map( A1 => n1324, A2 => n12725, ZN => n12460);
   U8939 : NAND2_X1 port map( A1 => n3543, A2 => n3545, ZN => n3542);
   U8940 : NAND2_X1 port map( A1 => n24386, A2 => n4435, ZN => n16885);
   U8941 : OAI21_X2 port map( B1 => n22944, B2 => n4632, A => n3718, ZN => 
                           n3720);
   U8942 : AND2_X1 port map( A1 => n21863, A2 => n23902, ZN => n22547);
   U8943 : NAND2_X1 port map( A1 => n5290, A2 => n18765, ZN => n19308);
   U8944 : AOI22_X2 port map( A1 => n3010, A2 => n12842, B1 => n12841, B2 => 
                           n12958, ZN => n14339);
   U8945 : OAI21_X1 port map( B1 => n3013, B2 => n7773, A => n3012, ZN => n6127
                           );
   U8946 : NAND2_X1 port map( A1 => n6113, A2 => n3013, ZN => n3012);
   U8947 : NAND2_X1 port map( A1 => n25252, A2 => n7526, ZN => n7773);
   U8948 : NAND3_X1 port map( A1 => n11214, A2 => n11212, A3 => n10812, ZN => 
                           n5627);
   U8949 : MUX2_X1 port map( A => n10555, B => n4736, S => n417, Z => n4740);
   U8951 : NAND2_X1 port map( A1 => n15656, A2 => n16381, ZN => n4835);
   U8952 : AOI21_X1 port map( B1 => n22290, B2 => n22291, A => n3018, ZN => 
                           n22292);
   U8953 : AND2_X1 port map( A1 => n22289, A2 => n22387, ZN => n3018);
   U8954 : NAND3_X1 port map( A1 => n3124, A2 => n23238, A3 => n23237, ZN => 
                           n3123);
   U8955 : XNOR2_X1 port map( A => n17756, B => n24536, ZN => n18049);
   U8956 : INV_X1 port map( A => n14373, ZN => n4834);
   U8957 : NAND3_X1 port map( A1 => n23743, A2 => n23748, A3 => n23740, ZN => 
                           n3097);
   U8958 : NAND3_X1 port map( A1 => n19951, A2 => n20587, A3 => n20590, ZN => 
                           n3466);
   U8962 : NAND2_X1 port map( A1 => n7514, A2 => n7977, ZN => n7405);
   U8963 : NOR2_X1 port map( A1 => n13995, A2 => n25435, ZN => n4560);
   U8964 : INV_X1 port map( A => n10799, ZN => n4527);
   U8965 : XNOR2_X1 port map( A => n3022, B => n12045, ZN => n11708);
   U8966 : XNOR2_X1 port map( A => n11705, B => n12121, ZN => n3022);
   U8970 : NAND2_X1 port map( A1 => n22391, A2 => n22974, ZN => n3024);
   U8971 : NAND2_X1 port map( A1 => n22868, A2 => n23411, ZN => n3025);
   U8973 : NOR2_X1 port map( A1 => n23356, A2 => n23355, ZN => n3027);
   U8974 : NOR2_X1 port map( A1 => n13712, A2 => n14361, ZN => n3030);
   U8975 : INV_X1 port map( A => n13711, ZN => n3031);
   U8976 : NOR2_X1 port map( A1 => n22415, A2 => n23300, ZN => n23309);
   U8977 : OAI211_X1 port map( C1 => n7582, C2 => n7581, A => n7583, B => n7882
                           , ZN => n5489);
   U8978 : NAND3_X1 port map( A1 => n3796, A2 => n20569, A3 => n20570, ZN => 
                           n3032);
   U8979 : OAI21_X1 port map( B1 => n3034, B2 => n24583, A => n3033, ZN => 
                           n18936);
   U8980 : NAND2_X1 port map( A1 => n24583, A2 => n19326, ZN => n3033);
   U8981 : INV_X1 port map( A => n18935, ZN => n3034);
   U8982 : OAI21_X1 port map( B1 => n21915, B2 => n22404, A => n22397, ZN => 
                           n3035);
   U8983 : XNOR2_X1 port map( A => n3036, B => n23191, ZN => Ciphertext(30));
   U8985 : XNOR2_X1 port map( A => n3038, B => n24100, ZN => n20779);
   U8986 : NAND2_X1 port map( A1 => n3040, A2 => n23418, ZN => n23400);
   U8987 : OAI21_X1 port map( B1 => n24978, B2 => n24426, A => n23416, ZN => 
                           n3040);
   U8990 : NAND3_X2 port map( A1 => n17303, A2 => n17302, A3 => n3376, ZN => 
                           n18465);
   U8991 : NAND2_X1 port map( A1 => n20210, A2 => n20597, ZN => n3044);
   U8993 : NAND2_X1 port map( A1 => n20209, A2 => n20208, ZN => n3046);
   U8994 : NAND2_X1 port map( A1 => n17029, A2 => n17030, ZN => n17032);
   U8995 : NAND2_X1 port map( A1 => n18968, A2 => n18967, ZN => n3844);
   U8997 : OAI22_X1 port map( A1 => n19251, A2 => n18862, B1 => n19252, B2 => 
                           n19592, ZN => n3047);
   U8999 : OR2_X1 port map( A1 => n6456, A2 => n6184, ZN => n6337);
   U9000 : NAND2_X1 port map( A1 => n12669, A2 => n24462, ZN => n3562);
   U9001 : XNOR2_X1 port map( A => n8556, B => n8557, ZN => n3048);
   U9002 : NAND2_X1 port map( A1 => n23364, A2 => n23365, ZN => n23367);
   U9004 : OAI21_X1 port map( B1 => n9867, B2 => n10053, A => n3049, ZN => 
                           n9245);
   U9005 : NAND2_X1 port map( A1 => n3052, A2 => n5512, ZN => n5511);
   U9006 : NOR2_X1 port map( A1 => n17211, A2 => n17016, ZN => n3052);
   U9007 : NAND2_X1 port map( A1 => n3589, A2 => n12713, ZN => n12430);
   U9008 : NAND2_X1 port map( A1 => n6940, A2 => n6683, ZN => n6144);
   U9009 : OAI21_X2 port map( B1 => n7322, B2 => n7326, A => n7325, ZN => n8771
                           );
   U9010 : OR2_X2 port map( A1 => n6157, A2 => n6158, ZN => n7382);
   U9011 : OAI21_X1 port map( B1 => n6953, B2 => n6949, A => n6141, ZN => n6157
                           );
   U9013 : OR2_X1 port map( A1 => n16655, A2 => n17134, ZN => n3053);
   U9014 : NAND2_X1 port map( A1 => n17129, A2 => n16655, ZN => n3054);
   U9015 : NAND2_X1 port map( A1 => n5714, A2 => n7800, ZN => n3056);
   U9016 : XNOR2_X1 port map( A => n3057, B => n15303, ZN => n14491);
   U9017 : XNOR2_X1 port map( A => n14490, B => n15446, ZN => n3057);
   U9020 : OAI211_X1 port map( C1 => n4341, C2 => n10445, A => n10751, B => 
                           n9553, ZN => n4040);
   U9021 : XNOR2_X1 port map( A => n18253, B => n5327, ZN => n5326);
   U9022 : OAI21_X1 port map( B1 => n24490, B2 => n12885, A => n3286, ZN => 
                           n12884);
   U9023 : XOR2_X1 port map( A => n12067, B => n3190, Z => n3361);
   U9024 : NAND2_X1 port map( A1 => n7675, A2 => n7672, ZN => n7227);
   U9026 : OAI21_X1 port map( B1 => n9403, B2 => n10734, A => n10731, ZN => 
                           n9404);
   U9029 : MUX2_X2 port map( A => n14134, B => n14133, S => n14132, Z => n15415
                           );
   U9031 : NAND2_X1 port map( A1 => n16415, A2 => n24231, ZN => n3060);
   U9033 : OAI21_X1 port map( B1 => n13793, B2 => n13579, A => n13769, ZN => 
                           n4592);
   U9034 : XNOR2_X1 port map( A => n17917, B => n17916, ZN => n18719);
   U9035 : NAND2_X1 port map( A1 => n3922, A2 => n6959, ZN => n6958);
   U9039 : INV_X1 port map( A => n12796, ZN => n3065);
   U9040 : NAND2_X1 port map( A1 => n25370, A2 => n24569, ZN => n3068);
   U9042 : MUX2_X2 port map( A => n17565, B => n17564, S => n5371, Z => n20317)
                           ;
   U9043 : NAND2_X1 port map( A1 => n20054, A2 => n25089, ZN => n20469);
   U9044 : NOR2_X1 port map( A1 => n13449, A2 => n13761, ZN => n3786);
   U9045 : INV_X1 port map( A => n7501, ZN => n7498);
   U9046 : NAND2_X1 port map( A1 => n9563, A2 => n8157, ZN => n9248);
   U9047 : AND2_X1 port map( A1 => n4117, A2 => n4118, ZN => n12495);
   U9048 : OAI21_X1 port map( B1 => n307, B2 => n4993, A => n9872, ZN => n3072)
                           ;
   U9049 : OR2_X1 port map( A1 => n13052, A2 => n13053, ZN => n4517);
   U9050 : INV_X1 port map( A => n3717, ZN => n14031);
   U9051 : XNOR2_X1 port map( A => n18100, B => n18099, ZN => n4139);
   U9052 : INV_X1 port map( A => n14245, ZN => n13200);
   U9053 : INV_X1 port map( A => n19275, ZN => n5572);
   U9056 : INV_X1 port map( A => n17165, ZN => n4774);
   U9057 : INV_X1 port map( A => n15191, ZN => n3234);
   U9058 : OAI22_X1 port map( A1 => n4885, A2 => n19609, B1 => n19610, B2 => 
                           n24310, ZN => n19611);
   U9059 : XNOR2_X1 port map( A => n14377, B => n15165, ZN => n14898);
   U9060 : NAND3_X1 port map( A1 => n10989, A2 => n10406, A3 => n3606, ZN => 
                           n3607);
   U9061 : NAND3_X1 port map( A1 => n3074, A2 => n6769, A3 => n6909, ZN => 
                           n6485);
   U9062 : NAND2_X1 port map( A1 => n6910, A2 => n6918, ZN => n3074);
   U9063 : NAND2_X1 port map( A1 => n23902, A2 => n25239, ZN => n3077);
   U9064 : NAND3_X1 port map( A1 => n23903, A2 => n23902, A3 => n23904, ZN => 
                           n3078);
   U9065 : NAND2_X1 port map( A1 => n10803, A2 => n10801, ZN => n3079);
   U9066 : NAND2_X1 port map( A1 => n21377, A2 => n3080, ZN => n23154);
   U9067 : OAI21_X1 port map( B1 => n21376, B2 => n22328, A => n22462, ZN => 
                           n3080);
   U9068 : NAND2_X1 port map( A1 => n3081, A2 => n14126, ZN => n13899);
   U9069 : OAI22_X1 port map( A1 => n13893, A2 => n14130, B1 => n13895, B2 => 
                           n4133, ZN => n3081);
   U9070 : NOR2_X1 port map( A1 => n16929, A2 => n24585, ZN => n16720);
   U9071 : OAI21_X1 port map( B1 => n13017, B2 => n13014, A => n12756, ZN => 
                           n13242);
   U9072 : XNOR2_X1 port map( A => n3086, B => n21398, ZN => Ciphertext(36));
   U9073 : NAND2_X1 port map( A1 => n14182, A2 => n13795, ZN => n13773);
   U9074 : NAND3_X1 port map( A1 => n6530, A2 => n6532, A3 => n6533, ZN => 
                           n5920);
   U9077 : NAND2_X1 port map( A1 => n3091, A2 => n3090, ZN => n22260);
   U9078 : NAND2_X1 port map( A1 => n25460, A2 => n22258, ZN => n3090);
   U9079 : NAND2_X1 port map( A1 => n22259, A2 => n997, ZN => n3091);
   U9081 : XNOR2_X2 port map( A => n5940, B => Key(5), ZN => n6510);
   U9082 : AOI21_X1 port map( B1 => n2953, B2 => n3292, A => n3289, ZN => 
                           n10208);
   U9083 : AND3_X1 port map( A1 => n5995, A2 => n5994, A3 => n6596, ZN => n3167
                           );
   U9084 : NAND2_X1 port map( A1 => n20192, A2 => n3198, ZN => n20434);
   U9085 : OAI21_X2 port map( B1 => n20327, B2 => n20571, A => n20326, ZN => 
                           n21606);
   U9086 : NAND2_X1 port map( A1 => n7602, A2 => n7257, ZN => n7258);
   U9088 : XNOR2_X1 port map( A => n14493, B => n21711, ZN => n14185);
   U9089 : XNOR2_X1 port map( A => n11915, B => n3812, ZN => n10239);
   U9090 : NAND3_X1 port map( A1 => n24286, A2 => n1357, A3 => n11151, ZN => 
                           n4999);
   U9091 : OR2_X1 port map( A1 => n6473, A2 => n6373, ZN => n6091);
   U9092 : NAND2_X1 port map( A1 => n12891, A2 => n13207, ZN => n13210);
   U9093 : XNOR2_X2 port map( A => n11358, B => n11359, ZN => n13207);
   U9095 : NAND2_X1 port map( A1 => n3094, A2 => n4262, ZN => n4260);
   U9096 : INV_X1 port map( A => n7108, ZN => n7747);
   U9100 : NAND2_X1 port map( A1 => n25460, A2 => n3096, ZN => n3095);
   U9101 : NOR2_X1 port map( A1 => n23748, A2 => n23730, ZN => n3096);
   U9103 : NAND3_X1 port map( A1 => n10799, A2 => n10649, A3 => n411, ZN => 
                           n3098);
   U9104 : INV_X1 port map( A => n10649, ZN => n3100);
   U9105 : NAND3_X2 port map( A1 => n3145, A2 => n11049, A3 => n3144, ZN => 
                           n12197);
   U9106 : NAND2_X1 port map( A1 => n3101, A2 => n22141, ZN => n3961);
   U9107 : NAND2_X1 port map( A1 => n21910, A2 => n22333, ZN => n3101);
   U9109 : OAI21_X2 port map( B1 => n3656, B2 => n20464, A => n3102, ZN => 
                           n21693);
   U9110 : NAND2_X1 port map( A1 => n20462, A2 => n20463, ZN => n3102);
   U9111 : OAI21_X1 port map( B1 => n6323, B2 => n6523, A => n6276, ZN => n3407
                           );
   U9112 : NAND2_X1 port map( A1 => n19304, A2 => n19132, ZN => n18765);
   U9114 : NAND2_X1 port map( A1 => n3104, A2 => n3103, ZN => n16650);
   U9115 : NAND2_X1 port map( A1 => n16648, A2 => n17088, ZN => n3104);
   U9116 : XNOR2_X1 port map( A => n3105, B => n9021, ZN => n9237);
   U9117 : XNOR2_X1 port map( A => n9019, B => n9020, ZN => n3105);
   U9118 : NAND2_X1 port map( A1 => n2008, A2 => n6697, ZN => n5897);
   U9119 : NAND2_X1 port map( A1 => n19207, A2 => n25474, ZN => n3106);
   U9120 : MUX2_X2 port map( A => n10289, B => n10288, S => n11111, Z => n12186
                           );
   U9121 : OR2_X1 port map( A1 => n10698, A2 => n25074, ZN => n10700);
   U9123 : INV_X1 port map( A => n18613, ZN => n18612);
   U9124 : XNOR2_X1 port map( A => n9015, B => n1864, ZN => n9018);
   U9125 : XNOR2_X1 port map( A => n7276, B => n8112, ZN => n3107);
   U9126 : NAND2_X1 port map( A1 => n7002, A2 => n6658, ZN => n3111);
   U9127 : OR2_X1 port map( A1 => n19105, A2 => n19107, ZN => n19202);
   U9128 : OR2_X1 port map( A1 => n10276, A2 => n10192, ZN => n4777);
   U9129 : INV_X1 port map( A => n15198, ZN => n3378);
   U9130 : INV_X1 port map( A => n13521, ZN => n14052);
   U9131 : NAND2_X1 port map( A1 => n16507, A2 => n3112, ZN => n17041);
   U9132 : NAND2_X1 port map( A1 => n16021, A2 => n16991, ZN => n3114);
   U9134 : NAND2_X1 port map( A1 => n10460, A2 => n10846, ZN => n10464);
   U9136 : INV_X1 port map( A => n16867, ZN => n18171);
   U9137 : NAND2_X1 port map( A1 => n9978, A2 => n9980, ZN => n9431);
   U9138 : NAND2_X1 port map( A1 => n3120, A2 => n12713, ZN => n12714);
   U9139 : OAI21_X1 port map( B1 => n12712, B2 => n12711, A => n12710, ZN => 
                           n3120);
   U9140 : NOR2_X2 port map( A1 => n4200, A2 => n13740, ZN => n15318);
   U9141 : XNOR2_X1 port map( A => n3123, B => n23239, ZN => Ciphertext(42));
   U9142 : INV_X1 port map( A => n11013, ZN => n11011);
   U9143 : NAND3_X1 port map( A1 => n6568, A2 => n6690, A3 => n6688, ZN => 
                           n6067);
   U9144 : INV_X1 port map( A => n19084, ZN => n19167);
   U9145 : OAI22_X1 port map( A1 => n13339, A2 => n231, B1 => n13337, B2 => 
                           n13338, ZN => n3126);
   U9146 : OAI21_X1 port map( B1 => n4672, B2 => n7947, A => n7656, ZN => n4784
                           );
   U9147 : NOR2_X1 port map( A1 => n22458, A2 => n5584, ZN => n5583);
   U9149 : NOR2_X1 port map( A1 => n275, A2 => n20094, ZN => n3127);
   U9150 : NOR2_X1 port map( A1 => n23683, A2 => n3128, ZN => Ciphertext(128));
   U9151 : AND2_X1 port map( A1 => n23684, A2 => n23685, ZN => n3128);
   U9154 : NAND2_X1 port map( A1 => n6906, A2 => n6372, ZN => n5250);
   U9155 : NAND3_X1 port map( A1 => n3130, A2 => n7583, A3 => n7312, ZN => 
                           n5859);
   U9156 : OR2_X1 port map( A1 => n10161, A2 => n10162, ZN => n10163);
   U9157 : MUX2_X2 port map( A => n16330, B => n16329, S => n16328, Z => n16979
                           );
   U9158 : NAND4_X2 port map( A1 => n15644, A2 => n15643, A3 => n15645, A4 => 
                           n15642, ZN => n16921);
   U9159 : NOR2_X1 port map( A1 => n404, A2 => n13274, ZN => n4389);
   U9160 : XOR2_X1 port map( A => n18283, B => n3073, Z => n5374);
   U9161 : INV_X1 port map( A => n14459, ZN => n13601);
   U9162 : OAI21_X1 port map( B1 => n18721, B2 => n19501, A => n4585, ZN => 
                           n18846);
   U9163 : XNOR2_X1 port map( A => n5373, B => n18286, ZN => n18288);
   U9165 : INV_X1 port map( A => n4590, ZN => n10771);
   U9166 : NAND2_X1 port map( A1 => n7307, A2 => n7647, ZN => n7765);
   U9167 : NAND2_X1 port map( A1 => n19962, A2 => n20370, ZN => n19963);
   U9168 : OAI21_X1 port map( B1 => n7576, B2 => n7318, A => n3548, ZN => n3300
                           );
   U9170 : AND2_X1 port map( A1 => n9212, A2 => n9211, ZN => n3134);
   U9171 : INV_X1 port map( A => n14360, ZN => n13568);
   U9172 : OAI21_X1 port map( B1 => n13587, B2 => n14359, A => n13586, ZN => 
                           n5527);
   U9173 : INV_X1 port map( A => n3461, ZN => n5323);
   U9174 : OAI22_X1 port map( A1 => n13627, A2 => n13843, B1 => n14063, B2 => 
                           n13847, ZN => n14265);
   U9175 : NOR2_X1 port map( A1 => n3324, A2 => n10756, ZN => n10755);
   U9176 : NAND2_X1 port map( A1 => n9301, A2 => n25043, ZN => n8609);
   U9177 : NAND2_X1 port map( A1 => n4140, A2 => n18120, ZN => n18135);
   U9178 : NAND2_X1 port map( A1 => n22583, A2 => n24559, ZN => n3135);
   U9179 : NAND2_X1 port map( A1 => n21238, A2 => n22803, ZN => n3136);
   U9180 : NAND2_X1 port map( A1 => n21237, A2 => n22799, ZN => n3137);
   U9181 : NAND3_X1 port map( A1 => n23507, A2 => n3139, A3 => n3138, ZN => 
                           n23509);
   U9182 : NAND2_X1 port map( A1 => n23504, A2 => n23531, ZN => n3138);
   U9183 : NAND2_X1 port map( A1 => n23513, A2 => n23503, ZN => n3139);
   U9184 : NAND2_X1 port map( A1 => n4950, A2 => n22919, ZN => n4949);
   U9185 : NAND2_X1 port map( A1 => n19657, A2 => n19850, ZN => n3140);
   U9186 : XOR2_X1 port map( A => n15409, B => n23620, Z => n4636);
   U9188 : NAND3_X1 port map( A1 => n5232, A2 => n9961, A3 => n3292, ZN => 
                           n3216);
   U9189 : OR2_X1 port map( A1 => n11174, A2 => n1338, ZN => n11176);
   U9190 : MUX2_X1 port map( A => n7405, B => n7406, S => n4400, Z => n7407);
   U9191 : NAND3_X1 port map( A1 => n10262, A2 => n10729, A3 => n10481, ZN => 
                           n10266);
   U9192 : XNOR2_X1 port map( A => n21029, B => n21030, ZN => n3141);
   U9193 : NAND2_X1 port map( A1 => n11047, A2 => n11048, ZN => n3145);
   U9194 : XNOR2_X2 port map( A => n8043, B => n8042, ZN => n9857);
   U9197 : AOI21_X1 port map( B1 => n3147, B2 => n3146, A => n23887, ZN => 
                           Ciphertext(170));
   U9198 : INV_X1 port map( A => n23877, ZN => n3146);
   U9199 : NAND2_X1 port map( A1 => n23878, A2 => n23879, ZN => n3147);
   U9200 : OAI21_X1 port map( B1 => n10095, B2 => n421, A => n3148, ZN => n9794
                           );
   U9201 : NAND2_X1 port map( A1 => n9790, A2 => n10095, ZN => n3148);
   U9202 : INV_X1 port map( A => n5009, ZN => n15351);
   U9205 : XNOR2_X1 port map( A => n3149, B => n23973, ZN => Ciphertext(183));
   U9206 : NAND2_X1 port map( A1 => n23971, A2 => n3150, ZN => n3149);
   U9207 : XNOR2_X1 port map( A => n14634, B => n15316, ZN => n14556);
   U9209 : NAND2_X1 port map( A1 => n7699, A2 => n7217, ZN => n7215);
   U9210 : NAND2_X1 port map( A1 => n6437, A2 => n5144, ZN => n3153);
   U9212 : NAND2_X1 port map( A1 => n24577, A2 => n7713, ZN => n7719);
   U9213 : NAND2_X1 port map( A1 => n5623, A2 => n7630, ZN => n5622);
   U9214 : NAND2_X1 port map( A1 => n23571, A2 => n23576, ZN => n22201);
   U9215 : INV_X1 port map( A => n7698, ZN => n7700);
   U9216 : OAI211_X1 port map( C1 => n23418, C2 => n142, A => n23402, B => 
                           n3157, ZN => n3156);
   U9218 : MUX2_X2 port map( A => n14177, B => n14176, S => n16204, Z => n17227
                           );
   U9220 : XNOR2_X1 port map( A => n3159, B => n21661, ZN => n21667);
   U9221 : XNOR2_X1 port map( A => n21663, B => n21660, ZN => n3159);
   U9222 : OAI21_X1 port map( B1 => n25299, B2 => n22243, A => n3160, ZN => 
                           n22183);
   U9223 : NAND2_X1 port map( A1 => n1336, A2 => n22243, ZN => n3160);
   U9224 : XNOR2_X1 port map( A => n3162, B => n21469, ZN => n4657);
   U9225 : XNOR2_X1 port map( A => n21306, B => n23798, ZN => n3162);
   U9226 : INV_X1 port map( A => n3811, ZN => n3810);
   U9227 : NAND2_X1 port map( A1 => n19592, A2 => n19587, ZN => n19251);
   U9228 : OR2_X2 port map( A1 => n11723, A2 => n5174, ZN => n11806);
   U9229 : NAND2_X1 port map( A1 => n9523, A2 => n25207, ZN => n4586);
   U9230 : OR3_X1 port map( A1 => n17464, A2 => n17463, A3 => n16499, ZN => 
                           n4970);
   U9232 : OR2_X1 port map( A1 => n7247, A2 => n7855, ZN => n7248);
   U9233 : OAI21_X1 port map( B1 => n16943, B2 => n17613, A => n16941, ZN => 
                           n16944);
   U9234 : NAND3_X1 port map( A1 => n16304, A2 => n16023, A3 => n15773, ZN => 
                           n15022);
   U9235 : XNOR2_X1 port map( A => n8268, B => n8269, ZN => n3307);
   U9237 : NAND2_X1 port map( A1 => n400, A2 => n13336, ZN => n5505);
   U9239 : NAND2_X1 port map( A1 => n6650, A2 => n7007, ZN => n6834);
   U9240 : NAND3_X1 port map( A1 => n11057, A2 => n11054, A3 => n11499, ZN => 
                           n3163);
   U9241 : OAI211_X2 port map( C1 => n13993, C2 => n14233, A => n13377, B => 
                           n13376, ZN => n15431);
   U9243 : OAI22_X1 port map( A1 => n10016, A2 => n25007, B1 => n10015, B2 => 
                           n25475, ZN => n3166);
   U9244 : NAND2_X1 port map( A1 => n7224, A2 => n7676, ZN => n4376);
   U9245 : NAND2_X1 port map( A1 => n10116, A2 => n10113, ZN => n9808);
   U9246 : XNOR2_X2 port map( A => n12204, B => n12205, ZN => n12856);
   U9247 : NAND2_X1 port map( A1 => n1149, A2 => n6975, ZN => n6979);
   U9248 : AND2_X2 port map( A1 => n20162, A2 => n20161, ZN => n21577);
   U9249 : NAND2_X1 port map( A1 => n3168, A2 => n13593, ZN => n13594);
   U9250 : OAI21_X1 port map( B1 => n14335, B2 => n25197, A => n13877, ZN => 
                           n3168);
   U9251 : NAND2_X1 port map( A1 => n3854, A2 => n17254, ZN => n3169);
   U9252 : XNOR2_X1 port map( A => n3170, B => n10917, ZN => n12510);
   U9253 : XNOR2_X1 port map( A => n12354, B => n11639, ZN => n3170);
   U9254 : NAND2_X1 port map( A1 => n24935, A2 => n16349, ZN => n15888);
   U9255 : INV_X1 port map( A => n7292, ZN => n5015);
   U9258 : OR2_X1 port map( A1 => n24512, A2 => n12540, ZN => n4946);
   U9260 : NAND2_X1 port map( A1 => n3172, A2 => n13103, ZN => n13106);
   U9261 : OAI22_X1 port map( A1 => n13185, A2 => n13102, B1 => n13101, B2 => 
                           n3958, ZN => n3172);
   U9265 : OAI211_X1 port map( C1 => n6528, C2 => n6255, A => n6947, B => n4757
                           , ZN => n4756);
   U9266 : OAI22_X2 port map( A1 => n12332, A2 => n12331, B1 => n5625, B2 => 
                           n12350, ZN => n13901);
   U9267 : XNOR2_X1 port map( A => n11564, B => n12297, ZN => n12028);
   U9269 : XNOR2_X1 port map( A => n14885, B => n14886, ZN => n15922);
   U9270 : XNOR2_X1 port map( A => n14880, B => n14879, ZN => n14881);
   U9271 : OR2_X1 port map( A1 => n6645, A2 => n6076, ZN => n3173);
   U9272 : INV_X1 port map( A => n9500, ZN => n4137);
   U9273 : NAND2_X1 port map( A1 => n16894, A2 => n16895, ZN => n4612);
   U9274 : INV_X1 port map( A => n18540, ZN => n17595);
   U9275 : XOR2_X1 port map( A => n8519, B => n8518, Z => n4138);
   U9276 : NAND3_X1 port map( A1 => n3174, A2 => n8022, A3 => n8021, ZN => 
                           n7746);
   U9277 : NAND2_X1 port map( A1 => n17085, A2 => n17086, ZN => n17089);
   U9278 : NAND2_X1 port map( A1 => n5280, A2 => n25473, ZN => n19024);
   U9279 : NAND2_X1 port map( A1 => n313, A2 => n6651, ZN => n6653);
   U9280 : NAND2_X1 port map( A1 => n3175, A2 => n23464, ZN => n22865);
   U9281 : OAI21_X1 port map( B1 => n24364, B2 => n23016, A => n23015, ZN => 
                           n3175);
   U9282 : INV_X1 port map( A => n22864, ZN => n3176);
   U9283 : OAI21_X1 port map( B1 => n3177, B2 => n15539, A => n16051, ZN => 
                           n15309);
   U9284 : NOR2_X1 port map( A1 => n4541, A2 => n16048, ZN => n3177);
   U9285 : NOR2_X1 port map( A1 => n14245, A2 => n13935, ZN => n14243);
   U9286 : XNOR2_X1 port map( A => n11915, B => n2145, ZN => n11799);
   U9288 : NAND3_X1 port map( A1 => n6985, A2 => n1130, A3 => n7898, ZN => 
                           n7900);
   U9289 : XNOR2_X1 port map( A => n3179, B => n21641, ZN => n21643);
   U9290 : XNOR2_X1 port map( A => n21675, B => n21638, ZN => n3179);
   U9291 : AOI21_X1 port map( B1 => n3180, B2 => n22724, A => n22938, ZN => 
                           n22726);
   U9292 : NAND2_X1 port map( A1 => n22723, A2 => n22722, ZN => n3180);
   U9293 : NAND3_X1 port map( A1 => n23011, A2 => n23479, A3 => n23480, ZN => 
                           n3181);
   U9294 : NOR2_X1 port map( A1 => n20598, A2 => n20427, ZN => n20425);
   U9295 : OAI211_X2 port map( C1 => n7716, C2 => n7561, A => n7560, B => n7559
                           , ZN => n8880);
   U9297 : NAND2_X1 port map( A1 => n9651, A2 => n9652, ZN => n9656);
   U9299 : NAND4_X2 port map( A1 => n9656, A2 => n9655, A3 => n3185, A4 => 
                           n9654, ZN => n11199);
   U9300 : NAND2_X1 port map( A1 => n9653, A2 => n10008, ZN => n3185);
   U9302 : MUX2_X1 port map( A => n12853, B => n12587, S => n12854, Z => n12589
                           );
   U9303 : XNOR2_X2 port map( A => n12188, B => n12187, ZN => n12854);
   U9304 : INV_X1 port map( A => n16269, ZN => n3186);
   U9305 : NAND2_X1 port map( A1 => n16004, A2 => n16268, ZN => n3187);
   U9306 : AOI21_X1 port map( B1 => n23386, B2 => n22032, A => n22031, ZN => 
                           n22041);
   U9307 : OAI22_X1 port map( A1 => n23033, A2 => n24972, B1 => n23034, B2 => 
                           n23830, ZN => n23035);
   U9308 : NAND2_X1 port map( A1 => n12758, A2 => n12784, ZN => n12761);
   U9309 : NAND2_X1 port map( A1 => n5832, A2 => n6885, ZN => n3188);
   U9311 : XNOR2_X1 port map( A => n17984, B => n17985, ZN => n19381);
   U9312 : NAND2_X1 port map( A1 => n10059, A2 => n10665, ZN => n3191);
   U9313 : OR2_X1 port map( A1 => n12928, A2 => n12897, ZN => n13281);
   U9314 : XNOR2_X1 port map( A => n8950, B => n8949, ZN => n9550);
   U9315 : NAND2_X1 port map( A1 => n6259, A2 => n24592, ZN => n5867);
   U9316 : XNOR2_X1 port map( A => n3193, B => n8249, ZN => n6048);
   U9317 : XNOR2_X1 port map( A => n9175, B => n5930, ZN => n3193);
   U9318 : NAND3_X2 port map( A1 => n16728, A2 => n3816, A3 => n16729, ZN => 
                           n4250);
   U9319 : XNOR2_X1 port map( A => n3194, B => n15183, ZN => n15186);
   U9320 : XNOR2_X1 port map( A => n15184, B => n21169, ZN => n3194);
   U9321 : INV_X1 port map( A => n11031, ZN => n11100);
   U9322 : NAND2_X1 port map( A1 => n3196, A2 => n4739, ZN => n4738);
   U9324 : XNOR2_X1 port map( A => n18451, B => n3197, ZN => n17701);
   U9325 : XNOR2_X2 port map( A => Key(123), B => Plaintext(123), ZN => n7008);
   U9326 : OAI21_X1 port map( B1 => n7891, B2 => n7890, A => n7889, ZN => n5054
                           );
   U9328 : NAND2_X1 port map( A1 => n9804, A2 => n9805, ZN => n10115);
   U9329 : NAND2_X1 port map( A1 => n3199, A2 => n10113, ZN => n5197);
   U9330 : NAND2_X1 port map( A1 => n10115, A2 => n9533, ZN => n3199);
   U9331 : NAND3_X1 port map( A1 => n3200, A2 => n13176, A3 => n10360, ZN => 
                           n12726);
   U9332 : NAND3_X1 port map( A1 => n13177, A2 => n13178, A3 => n3200, ZN => 
                           n13179);
   U9333 : INV_X1 port map( A => n12652, ZN => n3200);
   U9334 : NOR2_X1 port map( A1 => n22043, A2 => n3201, ZN => n22044);
   U9335 : NAND3_X1 port map( A1 => n21837, A2 => n24983, A3 => n4533, ZN => 
                           n21900);
   U9337 : OR2_X1 port map( A1 => n19389, A2 => n19386, ZN => n3202);
   U9339 : NAND2_X1 port map( A1 => n19388, A2 => n19389, ZN => n3203);
   U9340 : XNOR2_X2 port map( A => n17719, B => n17718, ZN => n19389);
   U9342 : XNOR2_X1 port map( A => n12133, B => n3207, ZN => n3205);
   U9346 : OAI21_X1 port map( B1 => n24881, B2 => n22973, A => n22387, ZN => 
                           n3211);
   U9347 : NOR2_X1 port map( A1 => n3213, A2 => n22977, ZN => n3212);
   U9349 : OR2_X1 port map( A1 => n18952, A2 => n24441, ZN => n3215);
   U9350 : NAND2_X1 port map( A1 => n3217, A2 => n3216, ZN => n11004);
   U9351 : NAND2_X1 port map( A1 => n7572, A2 => n8140, ZN => n3217);
   U9352 : MUX2_X1 port map( A => n17472, B => n17633, S => n16901, Z => n16793
                           );
   U9353 : INV_X1 port map( A => n19135, ZN => n18949);
   U9354 : NAND2_X1 port map( A1 => n3218, A2 => n19304, ZN => n19135);
   U9355 : INV_X1 port map( A => n19133, ZN => n3218);
   U9358 : NAND2_X1 port map( A1 => n4327, A2 => n3221, ZN => n3220);
   U9359 : NAND2_X1 port map( A1 => n399, A2 => n12956, ZN => n13339);
   U9361 : OAI21_X1 port map( B1 => n16400, B2 => n3223, A => n15972, ZN => 
                           n3222);
   U9362 : NOR2_X1 port map( A1 => n17453, A2 => n5072, ZN => n17454);
   U9363 : AOI22_X2 port map( A1 => n3225, A2 => n16368, B1 => n3224, B2 => 
                           n17180, ZN => n17450);
   U9364 : NAND2_X1 port map( A1 => n3299, A2 => n16367, ZN => n3224);
   U9365 : NAND2_X1 port map( A1 => n16365, A2 => n16366, ZN => n3225);
   U9366 : NAND2_X1 port map( A1 => n3229, A2 => n3231, ZN => n3228);
   U9367 : OAI21_X1 port map( B1 => n22233, B2 => n22234, A => n3230, ZN => 
                           n3229);
   U9368 : XNOR2_X1 port map( A => n3232, B => n15191, ZN => n13928);
   U9369 : XNOR2_X1 port map( A => n15374, B => n3234, ZN => n15377);
   U9370 : OAI211_X2 port map( C1 => n3238, C2 => n8014, A => n3237, B => n3235
                           , ZN => n9035);
   U9371 : NAND3_X1 port map( A1 => n7749, A2 => n8014, A3 => n25451, ZN => 
                           n3237);
   U9372 : INV_X1 port map( A => n19851, ZN => n3240);
   U9373 : OR2_X1 port map( A1 => n18847, A2 => n19334, ZN => n3239);
   U9374 : NAND2_X1 port map( A1 => n13486, A2 => n14000, ZN => n12678);
   U9375 : AOI21_X1 port map( B1 => n299, B2 => n13485, A => n14000, ZN => 
                           n13490);
   U9376 : NAND2_X1 port map( A1 => n13262, A2 => n14000, ZN => n4226);
   U9377 : XNOR2_X1 port map( A => n11644, B => n11643, ZN => n12440);
   U9378 : INV_X1 port map( A => n12440, ZN => n13162);
   U9381 : NAND3_X1 port map( A1 => n5347, A2 => n5350, A3 => n1480, ZN => 
                           n5349);
   U9383 : NAND2_X1 port map( A1 => n5106, A2 => n5621, ZN => n3243);
   U9386 : AND3_X2 port map( A1 => n3247, A2 => n3246, A3 => n4120, ZN => 
                           n10558);
   U9387 : NAND2_X1 port map( A1 => n9592, A2 => n10160, ZN => n3246);
   U9388 : NAND2_X1 port map( A1 => n10164, A2 => n10163, ZN => n3247);
   U9389 : NAND2_X1 port map( A1 => n3249, A2 => n9066, ZN => n3248);
   U9390 : INV_X1 port map( A => n12028, ZN => n12029);
   U9391 : OR2_X1 port map( A1 => n10939, A2 => n24591, ZN => n3250);
   U9392 : NAND2_X1 port map( A1 => n3253, A2 => n3386, ZN => n3251);
   U9393 : NAND2_X1 port map( A1 => n10313, A2 => n11168, ZN => n3253);
   U9394 : NAND2_X1 port map( A1 => n12955, A2 => n13330, ZN => n3255);
   U9395 : XNOR2_X2 port map( A => n12035, B => n12034, ZN => n13323);
   U9396 : XNOR2_X2 port map( A => n18107, B => n18108, ZN => n19112);
   U9397 : XNOR2_X1 port map( A => n4679, B => n18133, ZN => n19608);
   U9399 : AOI21_X1 port map( B1 => n3263, B2 => n8497, A => n9310, ZN => n3262
                           );
   U9400 : NAND2_X1 port map( A1 => n9998, A2 => n25453, ZN => n3263);
   U9401 : AOI21_X2 port map( B1 => n3264, B2 => n22958, A => n22861, ZN => 
                           n23416);
   U9403 : NAND3_X1 port map( A1 => n9658, A2 => n9747, A3 => n24535, ZN => 
                           n9663);
   U9404 : NAND2_X1 port map( A1 => n24577, A2 => n8370, ZN => n7841);
   U9405 : MUX2_X1 port map( A => n24878, B => n7713, S => n8368, Z => n3267);
   U9407 : XNOR2_X1 port map( A => n12275, B => n3269, ZN => n11167);
   U9408 : NAND2_X1 port map( A1 => n3271, A2 => n3270, ZN => n16222);
   U9409 : NAND3_X1 port map( A1 => n389, A2 => n16220, A3 => n16460, ZN => 
                           n3270);
   U9412 : XNOR2_X1 port map( A => n8731, B => n8421, ZN => n8425);
   U9414 : OAI21_X1 port map( B1 => n7479, B2 => n7954, A => n7478, ZN => n3272
                           );
   U9415 : NAND3_X1 port map( A1 => n6756, A2 => n3276, A3 => n5805, ZN => 
                           n3273);
   U9416 : NAND3_X1 port map( A1 => n19352, A2 => n19445, A3 => n25002, ZN => 
                           n3277);
   U9419 : NAND2_X1 port map( A1 => n3281, A2 => n23714, ZN => n22084);
   U9420 : NOR2_X1 port map( A1 => n23727, A2 => n22082, ZN => n3281);
   U9421 : NAND3_X1 port map( A1 => n23705, A2 => n23715, A3 => n3283, ZN => 
                           n23706);
   U9422 : AOI21_X1 port map( B1 => n23698, B2 => n3283, A => n3282, ZN => 
                           n23709);
   U9423 : NAND3_X1 port map( A1 => n22147, A2 => n22148, A3 => n3283, ZN => 
                           n4863);
   U9425 : NAND2_X1 port map( A1 => n12885, A2 => n13224, ZN => n3286);
   U9426 : NAND2_X1 port map( A1 => n13292, A2 => n13291, ZN => n3287);
   U9427 : MUX2_X1 port map( A => n12827, B => n13291, S => n12824, Z => n12825
                           );
   U9428 : NAND3_X1 port map( A1 => n24482, A2 => n16191, A3 => n16328, ZN => 
                           n3288);
   U9429 : NAND2_X1 port map( A1 => n3291, A2 => n3290, ZN => n3289);
   U9430 : OAI211_X1 port map( C1 => n9349, C2 => n9850, A => n3294, B => n3305
                           , ZN => n3293);
   U9431 : NAND2_X1 port map( A1 => n9349, A2 => n9384, ZN => n3294);
   U9432 : NAND2_X1 port map( A1 => n9383, A2 => n9592, ZN => n3295);
   U9433 : NAND2_X1 port map( A1 => n18987, A2 => n3296, ZN => n3297);
   U9434 : XNOR2_X2 port map( A => n17904, B => n17903, ZN => n19500);
   U9435 : NAND2_X1 port map( A1 => n13728, A2 => n24588, ZN => n3298);
   U9436 : NAND2_X1 port map( A1 => n15640, A2 => n16206, ZN => n3299);
   U9438 : NAND2_X1 port map( A1 => n3300, A2 => n7575, ZN => n7457);
   U9439 : NAND2_X1 port map( A1 => n3303, A2 => n3301, ZN => n14826);
   U9441 : NAND2_X1 port map( A1 => n3304, A2 => n13952, ZN => n14157);
   U9442 : NAND2_X1 port map( A1 => n5080, A2 => n13775, ZN => n3304);
   U9443 : AND2_X1 port map( A1 => n10728, A2 => n10482, ZN => n11184);
   U9444 : NAND2_X1 port map( A1 => n9385, A2 => n9520, ZN => n10257);
   U9445 : NAND2_X1 port map( A1 => n9386, A2 => n9832, ZN => n10259);
   U9446 : NAND3_X1 port map( A1 => n9522, A2 => n9521, A3 => n2257, ZN => 
                           n5492);
   U9447 : NAND2_X1 port map( A1 => n22390, A2 => n24881, ZN => n3309);
   U9448 : MUX2_X1 port map( A => n20960, B => n20961, S => n20451, Z => n20963
                           );
   U9449 : OAI21_X1 port map( B1 => n20451, B2 => n20159, A => n3310, ZN => 
                           n19945);
   U9450 : NAND2_X1 port map( A1 => n20159, A2 => n20377, ZN => n3310);
   U9451 : NAND2_X1 port map( A1 => n3313, A2 => n10595, ZN => n3312);
   U9452 : NAND2_X1 port map( A1 => n10425, A2 => n2311, ZN => n3313);
   U9453 : INV_X1 port map( A => n12530, ZN => n3314);
   U9455 : NAND3_X1 port map( A1 => n12773, A2 => n12471, A3 => n12470, ZN => 
                           n3315);
   U9457 : NAND2_X1 port map( A1 => n16327, A2 => n16197, ZN => n3318);
   U9458 : NAND2_X1 port map( A1 => n16196, A2 => n16195, ZN => n3319);
   U9459 : NAND2_X1 port map( A1 => n3321, A2 => n6652, ZN => n3320);
   U9460 : MUX2_X1 port map( A => n6895, B => n6651, S => n6358, Z => n3321);
   U9461 : NAND2_X1 port map( A1 => n6895, A2 => n6086, ZN => n6357);
   U9462 : XNOR2_X2 port map( A => n18593, B => n18592, ZN => n19418);
   U9463 : NAND2_X1 port map( A1 => n9374, A2 => n3324, ZN => n9375);
   U9464 : NAND2_X1 port map( A1 => n3325, A2 => n4909, ZN => n21481);
   U9465 : NAND2_X1 port map( A1 => n25388, A2 => n20109, ZN => n19885);
   U9466 : NAND2_X1 port map( A1 => n3327, A2 => n12865, ZN => n4181);
   U9467 : INV_X1 port map( A => n12272, ZN => n3327);
   U9468 : NAND2_X1 port map( A1 => n3330, A2 => n14166, ZN => n3329);
   U9469 : MUX2_X1 port map( A => n13744, B => n14165, S => n13742, Z => n3330)
                           ;
   U9470 : NOR2_X2 port map( A1 => n12449, A2 => n12448, ZN => n13742);
   U9472 : XNOR2_X1 port map( A => n12113, B => n12114, ZN => n12115);
   U9474 : XNOR2_X1 port map( A => n19832, B => n19833, ZN => n21847);
   U9475 : INV_X1 port map( A => n21847, ZN => n3336);
   U9476 : OAI21_X1 port map( B1 => n21848, B2 => n22686, A => n3335, ZN => 
                           n21850);
   U9477 : NAND2_X1 port map( A1 => n3336, A2 => n21848, ZN => n3335);
   U9478 : INV_X1 port map( A => n3339, ZN => n3337);
   U9479 : AND2_X1 port map( A1 => n14205, A2 => n3341, ZN => n3340);
   U9480 : OR2_X2 port map( A1 => n12962, A2 => n12961, ZN => n3341);
   U9481 : NAND2_X1 port map( A1 => n25209, A2 => n13931, ZN => n14247);
   U9482 : NAND2_X1 port map( A1 => n4059, A2 => n4057, ZN => n3342);
   U9483 : NAND2_X1 port map( A1 => n4057, A2 => n24573, ZN => n3343);
   U9484 : NAND2_X1 port map( A1 => n414, A2 => n11207, ZN => n10633);
   U9485 : INV_X1 port map( A => n7449, ZN => n3348);
   U9486 : INV_X1 port map( A => n25253, ZN => n3347);
   U9487 : NAND3_X1 port map( A1 => n3346, A2 => n7635, A3 => n6486, ZN => 
                           n3345);
   U9488 : NAND2_X1 port map( A1 => n13983, A2 => n13982, ZN => n3349);
   U9489 : NAND2_X1 port map( A1 => n13984, A2 => n13922, ZN => n3350);
   U9491 : MUX2_X1 port map( A => n13225, B => n13226, S => n24490, Z => n3351)
                           ;
   U9492 : NAND2_X1 port map( A1 => n14221, A2 => n14222, ZN => n3353);
   U9493 : NAND2_X1 port map( A1 => n3357, A2 => n11754, ZN => n3356);
   U9494 : NAND2_X1 port map( A1 => n13009, A2 => n24965, ZN => n3357);
   U9495 : NAND3_X1 port map( A1 => n19446, A2 => n19452, A3 => n19445, ZN => 
                           n19356);
   U9497 : INV_X1 port map( A => n4672, ZN => n3358);
   U9498 : OAI211_X2 port map( C1 => n3359, C2 => n6931, A => n6929, B => n6930
                           , ZN => n8897);
   U9499 : XNOR2_X1 port map( A => n11420, B => n3361, ZN => n3360);
   U9500 : NAND2_X1 port map( A1 => n3362, A2 => n7474, ZN => n7066);
   U9501 : NOR2_X1 port map( A1 => n3362, A2 => n7421, ZN => n7954);
   U9502 : NAND2_X1 port map( A1 => n7423, A2 => n3362, ZN => n7220);
   U9503 : NAND2_X1 port map( A1 => n7477, A2 => n7475, ZN => n3363);
   U9504 : NAND2_X1 port map( A1 => n1380, A2 => n7573, ZN => n3365);
   U9505 : NAND2_X1 port map( A1 => n3366, A2 => n7580, ZN => n7319);
   U9506 : NAND3_X1 port map( A1 => n3366, A2 => n7580, A3 => n7575, ZN => 
                           n4347);
   U9507 : NAND2_X1 port map( A1 => n5809, A2 => n3366, ZN => n5815);
   U9508 : NAND2_X1 port map( A1 => n10005, A2 => n10007, ZN => n9723);
   U9510 : INV_X1 port map( A => n9481, ZN => n10005);
   U9511 : NAND3_X1 port map( A1 => n14317, A2 => n14458, A3 => n14319, ZN => 
                           n3367);
   U9512 : NAND2_X1 port map( A1 => n13868, A2 => n13500, ZN => n3368);
   U9514 : XNOR2_X1 port map( A => n15177, B => n14815, ZN => n14402);
   U9515 : NAND2_X1 port map( A1 => n5522, A2 => n3371, ZN => n15998);
   U9516 : NOR2_X1 port map( A1 => n17043, A2 => n3374, ZN => n17576);
   U9517 : AOI22_X1 port map( A1 => n17372, A2 => n3371, B1 => n17373, B2 => 
                           n3374, ZN => n17374);
   U9518 : AOI22_X1 port map( A1 => n16678, A2 => n3374, B1 => n17572, B2 => 
                           n16677, ZN => n16679);
   U9519 : OAI211_X1 port map( C1 => n16767, C2 => n3374, A => n3373, B => 
                           n3372, ZN => n18233);
   U9520 : NAND2_X1 port map( A1 => n16766, A2 => n3374, ZN => n3373);
   U9521 : OR2_X2 port map( A1 => n15964, A2 => n15963, ZN => n5522);
   U9522 : NAND3_X1 port map( A1 => n1055, A2 => n11092, A3 => n11302, ZN => 
                           n3375);
   U9523 : OAI211_X1 port map( C1 => n11302, C2 => n9536, A => n3375, B => 
                           n1056, ZN => n9537);
   U9524 : INV_X1 port map( A => n16708, ZN => n3377);
   U9525 : NAND2_X1 port map( A1 => n1473, A2 => n16708, ZN => n3376);
   U9527 : NAND3_X1 port map( A1 => n16615, A2 => n17296, A3 => n3377, ZN => 
                           n15731);
   U9528 : NAND2_X1 port map( A1 => n3378, A2 => n25410, ZN => n16009);
   U9529 : OAI21_X1 port map( B1 => n16315, B2 => n3378, A => n16311, ZN => 
                           n15768);
   U9530 : OAI21_X1 port map( B1 => n16309, B2 => n3378, A => n3554, ZN => 
                           n16314);
   U9531 : AOI21_X1 port map( B1 => n15752, B2 => n3378, A => n16312, ZN => 
                           n15753);
   U9532 : NAND3_X1 port map( A1 => n19390, A2 => n19630, A3 => n24909, ZN => 
                           n3379);
   U9533 : OAI21_X1 port map( B1 => n16206, B2 => n3380, A => n17182, ZN => 
                           n14177);
   U9534 : OR2_X1 port map( A1 => n16367, A2 => n15640, ZN => n17182);
   U9535 : NAND3_X1 port map( A1 => n16367, A2 => n17180, A3 => n3380, ZN => 
                           n15910);
   U9537 : NAND3_X1 port map( A1 => n13529, A2 => n3382, A3 => n3381, ZN => 
                           n14892);
   U9538 : OAI21_X1 port map( B1 => n12445, B2 => n3383, A => n13526, ZN => 
                           n3382);
   U9539 : XNOR2_X1 port map( A => n11957, B => n11959, ZN => n12320);
   U9540 : NAND2_X1 port map( A1 => n11169, A2 => n11168, ZN => n11174);
   U9541 : NAND3_X1 port map( A1 => n3386, A2 => n11175, A3 => n24591, ZN => 
                           n3385);
   U9542 : NAND3_X1 port map( A1 => n3387, A2 => n10586, A3 => n10587, ZN => 
                           n10593);
   U9543 : NAND2_X1 port map( A1 => n10582, A2 => n10583, ZN => n3387);
   U9544 : NAND3_X1 port map( A1 => n18037, A2 => n19602, A3 => n19596, ZN => 
                           n3389);
   U9545 : NAND2_X1 port map( A1 => n16577, A2 => n17131, ZN => n3392);
   U9546 : NAND2_X1 port map( A1 => n5337, A2 => n3393, ZN => n19248);
   U9547 : NAND2_X1 port map( A1 => n3394, A2 => n19575, ZN => n3393);
   U9548 : INV_X1 port map( A => n19578, ZN => n3394);
   U9549 : NAND2_X1 port map( A1 => n25072, A2 => n19248, ZN => n4425);
   U9550 : XNOR2_X1 port map( A => n17592, B => n18283, ZN => n3397);
   U9551 : NAND3_X1 port map( A1 => n4774, A2 => n16375, A3 => n16262, ZN => 
                           n3395);
   U9552 : NAND2_X1 port map( A1 => n16089, A2 => n17165, ZN => n3396);
   U9553 : XNOR2_X1 port map( A => n3397, B => n18375, ZN => n18044);
   U9554 : XNOR2_X1 port map( A => n3398, B => n1466, ZN => n9365);
   U9555 : XNOR2_X1 port map( A => n9137, B => n9138, ZN => n3398);
   U9557 : INV_X1 port map( A => n14320, ZN => n3402);
   U9558 : INV_X1 port map( A => n14321, ZN => n3404);
   U9560 : NAND2_X1 port map( A1 => n3402, A2 => n3401, ZN => n3400);
   U9561 : NAND2_X1 port map( A1 => n3404, A2 => n14320, ZN => n3403);
   U9562 : NAND2_X1 port map( A1 => n9382, A2 => n10162, ZN => n3405);
   U9563 : NAND2_X1 port map( A1 => n15933, A2 => n16231, ZN => n3406);
   U9564 : NAND3_X1 port map( A1 => n17662, A2 => n3131, A3 => n17661, ZN => 
                           n16969);
   U9565 : NAND3_X1 port map( A1 => n16105, A2 => n25409, A3 => n3410, ZN => 
                           n3408);
   U9566 : INV_X1 port map( A => n16102, ZN => n3410);
   U9568 : NAND2_X1 port map( A1 => n22800, A2 => n22798, ZN => n3411);
   U9569 : XNOR2_X2 port map( A => n21197, B => n21196, ZN => n22803);
   U9571 : INV_X1 port map( A => n3414, ZN => n6892);
   U9572 : OR2_X1 port map( A1 => n6651, A2 => n6893, ZN => n3413);
   U9573 : NAND3_X1 port map( A1 => n24345, A2 => n10302, A3 => n2386, ZN => 
                           n3415);
   U9574 : NAND3_X1 port map( A1 => n3419, A2 => n19254, A3 => n25001, ZN => 
                           n5027);
   U9575 : NAND2_X1 port map( A1 => n25244, A2 => n19596, ZN => n3419);
   U9576 : NOR2_X1 port map( A1 => n3419, A2 => n18870, ZN => n18873);
   U9577 : OAI21_X1 port map( B1 => n5561, B2 => n3421, A => n13051, ZN => 
                           n3420);
   U9578 : NOR2_X1 port map( A1 => n25408, A2 => n13049, ZN => n3421);
   U9579 : AND2_X1 port map( A1 => n4850, A2 => n13050, ZN => n5561);
   U9580 : NOR2_X1 port map( A1 => n13049, A2 => n12490, ZN => n3423);
   U9581 : NAND2_X1 port map( A1 => n13968, A2 => n13969, ZN => n3427);
   U9582 : NAND2_X1 port map( A1 => n3767, A2 => n3428, ZN => n5764);
   U9583 : INV_X1 port map( A => n3767, ZN => n3429);
   U9585 : MUX2_X1 port map( A => n17050, B => n17049, S => n17048, Z => n3432)
                           ;
   U9586 : NAND2_X1 port map( A1 => n3435, A2 => n3434, ZN => n3433);
   U9587 : NAND2_X1 port map( A1 => n17053, A2 => n17048, ZN => n17052);
   U9588 : NAND2_X1 port map( A1 => n24162, A2 => n16016, ZN => n15941);
   U9589 : NAND2_X1 port map( A1 => n24162, A2 => n3436, ZN => n3437);
   U9590 : AND2_X1 port map( A1 => n16246, A2 => n16016, ZN => n3436);
   U9592 : NAND3_X1 port map( A1 => n392, A2 => n13080, A3 => n13081, ZN => 
                           n13559);
   U9593 : AOI21_X1 port map( B1 => n24984, B2 => n9384, A => n3438, ZN => 
                           n9854);
   U9594 : AND2_X1 port map( A1 => n9348, A2 => n10158, ZN => n3438);
   U9597 : NAND2_X1 port map( A1 => n12719, A2 => n13167, ZN => n12447);
   U9598 : NAND2_X1 port map( A1 => n3445, A2 => n24051, ZN => n3444);
   U9599 : NAND2_X1 port map( A1 => n24051, A2 => n24500, ZN => n6719);
   U9600 : NAND2_X1 port map( A1 => n9410, A2 => n10452, ZN => n3446);
   U9601 : NAND2_X1 port map( A1 => n9411, A2 => n10290, ZN => n3447);
   U9602 : XNOR2_X1 port map( A => n3448, B => n4670, ZN => n11504);
   U9603 : XNOR2_X1 port map( A => n11504, B => n11505, ZN => n11508);
   U9604 : OAI22_X1 port map( A1 => n4496, A2 => n24841, B1 => n16359, B2 => 
                           n3450, ZN => n3449);
   U9605 : NAND2_X1 port map( A1 => n3451, A2 => n16355, ZN => n3450);
   U9606 : INV_X1 port map( A => n16356, ZN => n3451);
   U9607 : INV_X1 port map( A => n1355, ZN => n3453);
   U9608 : OAI21_X1 port map( B1 => n13518, B2 => n13521, A => n3453, ZN => 
                           n3452);
   U9609 : NAND2_X1 port map( A1 => n14050, A2 => n1355, ZN => n3455);
   U9610 : INV_X1 port map( A => n3456, ZN => n22055);
   U9611 : NAND2_X1 port map( A1 => n336, A2 => n21829, ZN => n3456);
   U9613 : NOR2_X1 port map( A1 => n25244, A2 => n19071, ZN => n18831);
   U9614 : NOR2_X1 port map( A1 => n3461, A2 => n13094, ZN => n13095);
   U9615 : NOR2_X1 port map( A1 => n3461, A2 => n3492, ZN => n12505);
   U9616 : NOR2_X1 port map( A1 => n4405, A2 => n3461, ZN => n10199);
   U9617 : OAI21_X1 port map( B1 => n13093, B2 => n3461, A => n3460, ZN => 
                           n4906);
   U9618 : NAND2_X1 port map( A1 => n3461, A2 => n12648, ZN => n3460);
   U9619 : XNOR2_X1 port map( A => n25394, B => n14816, ZN => n14115);
   U9620 : XNOR2_X1 port map( A => n25394, B => n15002, ZN => n15004);
   U9621 : XNOR2_X1 port map( A => n14889, B => n25394, ZN => n15084);
   U9622 : NAND2_X1 port map( A1 => n3464, A2 => n13788, ZN => n3463);
   U9623 : NAND2_X1 port map( A1 => n14188, A2 => n14142, ZN => n3464);
   U9625 : INV_X1 port map( A => n19953, ZN => n20587);
   U9626 : NAND2_X1 port map( A1 => n4143, A2 => n10772, ZN => n10910);
   U9628 : NAND2_X1 port map( A1 => n7897, A2 => n3469, ZN => n7140);
   U9629 : NAND3_X1 port map( A1 => n7898, A2 => n7232, A3 => n3469, ZN => 
                           n5236);
   U9630 : INV_X1 port map( A => n3471, ZN => n14599);
   U9631 : NAND2_X1 port map( A1 => n9211, A2 => n3472, ZN => n9380);
   U9632 : NAND2_X1 port map( A1 => n10125, A2 => n3472, ZN => n10126);
   U9633 : NAND2_X1 port map( A1 => n5057, A2 => n3472, ZN => n9597);
   U9634 : AOI21_X1 port map( B1 => n10130, B2 => n9211, A => n3472, ZN => 
                           n10131);
   U9635 : OAI21_X1 port map( B1 => n5057, B2 => n3472, A => n7437, ZN => n7438
                           );
   U9636 : INV_X1 port map( A => n13274, ZN => n12963);
   U9637 : MUX2_X1 port map( A => n12695, B => n404, S => n13274, Z => n12697);
   U9638 : NOR2_X1 port map( A1 => n24967, A2 => n23220, ZN => n3475);
   U9639 : NOR2_X1 port map( A1 => n23212, A2 => n3475, ZN => n23232);
   U9640 : NAND2_X1 port map( A1 => n7991, A2 => n7993, ZN => n7414);
   U9641 : OAI21_X2 port map( B1 => n6677, B2 => n271, A => n6676, ZN => n7993)
                           ;
   U9642 : XNOR2_X1 port map( A => n21559, B => n2120, ZN => n21127);
   U9646 : NAND2_X1 port map( A1 => n20330, A2 => n3482, ZN => n3481);
   U9647 : NAND2_X1 port map( A1 => n18136, A2 => n20089, ZN => n3483);
   U9648 : XNOR2_X1 port map( A => n3484, B => n24009, ZN => Ciphertext(189));
   U9649 : OAI211_X1 port map( C1 => n24018, C2 => n24008, A => n3487, B => 
                           n3485, ZN => n3484);
   U9650 : NAND2_X1 port map( A1 => n24008, A2 => n5773, ZN => n3487);
   U9651 : NAND2_X1 port map( A1 => n806, A2 => n3488, ZN => n7073);
   U9652 : NAND2_X1 port map( A1 => n9247, A2 => n3489, ZN => n4594);
   U9653 : NAND2_X1 port map( A1 => n9326, A2 => n9787, ZN => n10087);
   U9654 : NAND2_X1 port map( A1 => n9507, A2 => n9787, ZN => n4208);
   U9655 : MUX2_X1 port map( A => n10080, B => n9507, S => n9787, Z => n8466);
   U9656 : NAND2_X1 port map( A1 => n9789, A2 => n9787, ZN => n9307);
   U9657 : NAND3_X1 port map( A1 => n3491, A2 => n19412, A3 => n19173, ZN => 
                           n19174);
   U9658 : MUX2_X1 port map( A => n5324, B => n5323, S => n4405, Z => n13098);
   U9659 : NAND2_X1 port map( A1 => n15795, A2 => n15794, ZN => n3494);
   U9661 : NAND2_X1 port map( A1 => n3495, A2 => n4533, ZN => n4953);
   U9662 : NAND2_X1 port map( A1 => n4533, A2 => n22043, ZN => n23792);
   U9663 : NAND2_X1 port map( A1 => n3497, A2 => n7789, ZN => n3496);
   U9664 : NAND2_X1 port map( A1 => n7441, A2 => n7788, ZN => n3497);
   U9665 : NAND2_X1 port map( A1 => n7781, A2 => n7787, ZN => n7441);
   U9666 : MUX2_X1 port map( A => n7579, B => n7578, S => n7577, Z => n3499);
   U9667 : OAI21_X1 port map( B1 => n14038, B2 => n3501, A => n14319, ZN => 
                           n5058);
   U9668 : AOI21_X1 port map( B1 => n14461, B2 => n14460, A => n1474, ZN => 
                           n14463);
   U9669 : XNOR2_X1 port map( A => n11660, B => n12391, ZN => n10196);
   U9671 : NAND3_X1 port map( A1 => n10283, A2 => n10859, A3 => n10855, ZN => 
                           n3502);
   U9672 : NOR2_X2 port map( A1 => n15798, A2 => n15787, ZN => n17134);
   U9674 : XNOR2_X1 port map( A => n8112, B => n8115, ZN => n3504);
   U9675 : XNOR2_X1 port map( A => n8114, B => n8113, ZN => n3505);
   U9677 : NAND2_X1 port map( A1 => n19206, A2 => n19381, ZN => n3508);
   U9679 : NAND2_X1 port map( A1 => n20131, A2 => n55, ZN => n19671);
   U9680 : NAND2_X1 port map( A1 => n3509, A2 => n4671, ZN => n3511);
   U9681 : INV_X1 port map( A => n10699, ZN => n3509);
   U9683 : NAND2_X1 port map( A1 => n2754, A2 => n25233, ZN => n3513);
   U9684 : NAND2_X1 port map( A1 => n266, A2 => n17012, ZN => n3515);
   U9685 : INV_X1 port map( A => n19094, ZN => n18877);
   U9686 : NOR2_X2 port map( A1 => n3518, A2 => n17986, ZN => n20554);
   U9687 : OAI21_X1 port map( B1 => n20518, B2 => n3519, A => n20517, ZN => 
                           n3520);
   U9688 : INV_X1 port map( A => n20516, ZN => n3519);
   U9690 : NAND2_X1 port map( A1 => n20273, A2 => n3522, ZN => n3521);
   U9691 : NAND2_X1 port map( A1 => n17078, A2 => n17075, ZN => n16892);
   U9692 : XNOR2_X1 port map( A => n15170, B => n14973, ZN => n3525);
   U9693 : XNOR2_X2 port map( A => n3525, B => n4115, ZN => n16449);
   U9694 : NAND2_X1 port map( A1 => n24911, A2 => n23375, ZN => n3527);
   U9695 : XNOR2_X1 port map( A => n3526, B => n22440, ZN => Ciphertext(76));
   U9696 : NAND3_X1 port map( A1 => n3528, A2 => n22439, A3 => n3527, ZN => 
                           n3526);
   U9697 : NAND3_X1 port map( A1 => n18944, A2 => n19472, A3 => n19322, ZN => 
                           n3529);
   U9698 : NAND3_X1 port map( A1 => n19471, A2 => n19322, A3 => n18956, ZN => 
                           n3530);
   U9699 : OAI22_X1 port map( A1 => n11116, A2 => n3532, B1 => n11111, B2 => 
                           n10725, ZN => n5335);
   U9700 : AOI21_X1 port map( B1 => n6235, B2 => n5784, A => n6232, ZN => n5785
                           );
   U9701 : MUX2_X1 port map( A => n6717, B => n6716, S => n6232, Z => n7074);
   U9702 : NAND2_X1 port map( A1 => n3533, A2 => n14064, ZN => n13430);
   U9703 : OAI21_X1 port map( B1 => n5694, B2 => n3533, A => n5693, ZN => n5692
                           );
   U9704 : INV_X1 port map( A => n18073, ZN => n17899);
   U9705 : XNOR2_X1 port map( A => n18073, B => n3535, ZN => n3534);
   U9706 : INV_X1 port map( A => n18523, ZN => n3535);
   U9709 : NAND2_X1 port map( A1 => n13806, A2 => n13805, ZN => n3539);
   U9710 : NAND2_X1 port map( A1 => n341, A2 => n20320, ZN => n3540);
   U9711 : INV_X1 port map( A => n24062, ZN => n3545);
   U9713 : NAND2_X1 port map( A1 => n16171, A2 => n244, ZN => n3547);
   U9714 : OAI21_X1 port map( B1 => n3366, B2 => n7579, A => n3548, ZN => n4345
                           );
   U9715 : NAND2_X1 port map( A1 => n7359, A2 => n7993, ZN => n3550);
   U9718 : OR2_X2 port map( A1 => n3552, A2 => n3551, ZN => n10411);
   U9719 : AOI21_X1 port map( B1 => n9591, B2 => n9590, A => n10168, ZN => 
                           n3552);
   U9721 : NAND2_X1 port map( A1 => n4677, A2 => n4676, ZN => n3556);
   U9722 : XNOR2_X1 port map( A => n14907, B => n23523, ZN => n14413);
   U9723 : AND2_X1 port map( A1 => n14240, A2 => n25209, ZN => n3557);
   U9724 : NAND2_X1 port map( A1 => n12805, A2 => n13017, ZN => n3559);
   U9727 : OR2_X1 port map( A1 => n12669, A2 => n3561, ZN => n12671);
   U9728 : NOR2_X1 port map( A1 => n12668, A2 => n13488, ZN => n3561);
   U9729 : AND2_X1 port map( A1 => n299, A2 => n12669, ZN => n13667);
   U9730 : OR2_X1 port map( A1 => n12669, A2 => n299, ZN => n5221);
   U9732 : NAND2_X1 port map( A1 => n14001, A2 => n3562, ZN => n14007);
   U9733 : OAI21_X1 port map( B1 => n23320, B2 => n23317, A => n3564, ZN => 
                           n21895);
   U9734 : MUX2_X1 port map( A => n23311, B => n24316, S => n23326, Z => n22384
                           );
   U9735 : OR2_X2 port map( A1 => n21877, A2 => n21876, ZN => n23326);
   U9736 : XNOR2_X1 port map( A => n11628, B => n445, ZN => n3565);
   U9737 : INV_X1 port map( A => n7516, ZN => n7404);
   U9741 : NAND2_X1 port map( A1 => n3571, A2 => n3570, ZN => n3569);
   U9742 : NAND2_X1 port map( A1 => n7554, A2 => n7863, ZN => n3572);
   U9743 : INV_X1 port map( A => n6922, ZN => n4042);
   U9744 : XNOR2_X2 port map( A => Key(167), B => Plaintext(167), ZN => n6198);
   U9745 : NAND2_X1 port map( A1 => n11000, A2 => n3573, ZN => n11001);
   U9746 : INV_X1 port map( A => n10907, ZN => n10747);
   U9747 : NAND2_X1 port map( A1 => n10902, A2 => n10907, ZN => n3574);
   U9748 : INV_X1 port map( A => n10751, ZN => n10902);
   U9749 : NAND2_X1 port map( A1 => n10747, A2 => n10746, ZN => n3575);
   U9750 : NAND3_X1 port map( A1 => n25409, A2 => n16101, A3 => n5100, ZN => 
                           n3592);
   U9753 : INV_X1 port map( A => n14625, ZN => n16038);
   U9754 : AND3_X2 port map( A1 => n3580, A2 => n3584, A3 => n3579, ZN => 
                           n20071);
   U9755 : NAND2_X1 port map( A1 => n3581, A2 => n19470, ZN => n3580);
   U9757 : NAND2_X1 port map( A1 => n22564, A2 => n21934, ZN => n22132);
   U9759 : AOI22_X1 port map( A1 => n22297, A2 => n25373, B1 => n3586, B2 => 
                           n3585, ZN => Ciphertext(44));
   U9760 : NAND2_X1 port map( A1 => n22294, A2 => n189, ZN => n3585);
   U9761 : NAND2_X1 port map( A1 => n3588, A2 => n7531, ZN => n3708);
   U9762 : NAND2_X1 port map( A1 => n3590, A2 => n12707, ZN => n12429);
   U9763 : NAND2_X1 port map( A1 => n13078, A2 => n24573, ZN => n3589);
   U9764 : NAND3_X1 port map( A1 => n12712, A2 => n12431, A3 => n3590, ZN => 
                           n12432);
   U9765 : NAND2_X1 port map( A1 => n11589, A2 => n3590, ZN => n11594);
   U9766 : NAND2_X1 port map( A1 => n24585, A2 => n17054, ZN => n17057);
   U9767 : OAI21_X1 port map( B1 => n16722, B2 => n24398, A => n3593, ZN => 
                           n16723);
   U9768 : NAND2_X1 port map( A1 => n10814, A2 => n10967, ZN => n3594);
   U9769 : NAND2_X1 port map( A1 => n9909, A2 => n9935, ZN => n3596);
   U9770 : NAND2_X1 port map( A1 => n17023, A2 => n3598, ZN => n3600);
   U9771 : NAND2_X1 port map( A1 => n16627, A2 => n17389, ZN => n3599);
   U9772 : XNOR2_X1 port map( A => n18261, B => n2717, ZN => n3605);
   U9773 : INV_X1 port map( A => n10326, ZN => n3606);
   U9775 : NAND3_X1 port map( A1 => n9814, A2 => n10169, A3 => n25046, ZN => 
                           n9589);
   U9776 : MUX2_X1 port map( A => n9814, B => n9817, S => n25046, Z => n8332);
   U9777 : NAND3_X1 port map( A1 => n16324, A2 => n24482, A3 => n16197, ZN => 
                           n16198);
   U9778 : NAND2_X1 port map( A1 => n15258, A2 => n24482, ZN => n5408);
   U9779 : INV_X1 port map( A => n8022, ZN => n3615);
   U9780 : NOR2_X1 port map( A1 => n7532, A2 => n8024, ZN => n3611);
   U9781 : NAND2_X1 port map( A1 => n3614, A2 => n7532, ZN => n3612);
   U9782 : XNOR2_X1 port map( A => n18467, B => n21335, ZN => n17430);
   U9783 : XNOR2_X1 port map( A => n18467, B => n729, ZN => n17797);
   U9784 : XNOR2_X1 port map( A => n18467, B => n2049, ZN => n18153);
   U9785 : INV_X1 port map( A => n19366, ZN => n19219);
   U9786 : OAI21_X1 port map( B1 => n24424, B2 => n24361, A => n3617, ZN => 
                           n5682);
   U9787 : NAND2_X1 port map( A1 => n24424, A2 => n19371, ZN => n3617);
   U9788 : OR2_X1 port map( A1 => n6878, A2 => n6768, ZN => n3618);
   U9789 : NAND3_X1 port map( A1 => n12917, A2 => n12612, A3 => n25248, ZN => 
                           n11714);
   U9791 : NOR2_X1 port map( A1 => n12612, A2 => n25248, ZN => n4789);
   U9792 : NAND2_X1 port map( A1 => n19060, A2 => n19059, ZN => n3620);
   U9794 : OR2_X1 port map( A1 => n22510, A2 => n23303, ZN => n3622);
   U9795 : NAND2_X1 port map( A1 => n22763, A2 => n22509, ZN => n3624);
   U9796 : INV_X1 port map( A => n23306, ZN => n3625);
   U9798 : NOR2_X1 port map( A1 => n12508, A2 => n12652, ZN => n3631);
   U9800 : OR2_X1 port map( A1 => n13614, A2 => n13610, ZN => n3634);
   U9802 : NAND2_X1 port map( A1 => n3635, A2 => n3634, ZN => n13616);
   U9803 : NAND2_X1 port map( A1 => n13611, A2 => n13614, ZN => n3635);
   U9804 : OAI211_X1 port map( C1 => n16130, C2 => n1365, A => n24826, B => 
                           n3636, ZN => n3639);
   U9807 : NAND2_X1 port map( A1 => n3638, A2 => n15800, ZN => n3637);
   U9808 : NOR2_X1 port map( A1 => n1365, A2 => n14664, ZN => n3638);
   U9809 : NAND2_X1 port map( A1 => n7663, A2 => n7662, ZN => n7670);
   U9810 : NAND2_X1 port map( A1 => n23999, A2 => n25079, ZN => n3641);
   U9811 : NOR2_X1 port map( A1 => n23994, A2 => n25079, ZN => n22676);
   U9814 : INV_X1 port map( A => n16670, ZN => n3645);
   U9817 : NAND3_X1 port map( A1 => n9899, A2 => n9286, A3 => n9287, ZN => 
                           n8139);
   U9819 : NAND2_X1 port map( A1 => n25021, A2 => n9898, ZN => n9286);
   U9820 : XNOR2_X1 port map( A => n21106, B => n23983, ZN => n21107);
   U9821 : NAND3_X1 port map( A1 => n19818, A2 => n20243, A3 => n20244, ZN => 
                           n3650);
   U9822 : NAND2_X1 port map( A1 => n3652, A2 => n3651, ZN => n19510);
   U9823 : NAND2_X1 port map( A1 => n19298, A2 => n19297, ZN => n3651);
   U9824 : NAND2_X1 port map( A1 => n19299, A2 => n3653, ZN => n3652);
   U9825 : NAND2_X1 port map( A1 => n1344, A2 => n19939, ZN => n19818);
   U9826 : NAND2_X1 port map( A1 => n9380, A2 => n9379, ZN => n10255);
   U9827 : OR2_X1 port map( A1 => n20462, A2 => n3656, ZN => n20396);
   U9828 : NAND2_X1 port map( A1 => n20393, A2 => n20394, ZN => n3657);
   U9829 : INV_X1 port map( A => n16004, ZN => n3658);
   U9830 : NAND2_X1 port map( A1 => n3658, A2 => n15758, ZN => n16270);
   U9834 : NOR2_X1 port map( A1 => n19275, A2 => n3773, ZN => n3661);
   U9835 : INV_X1 port map( A => n5573, ZN => n3662);
   U9837 : OAI21_X1 port map( B1 => n22358, B2 => n3664, A => n4203, ZN => 
                           n22045);
   U9838 : NAND2_X1 port map( A1 => n21348, A2 => n21782, ZN => n3664);
   U9839 : INV_X1 port map( A => n17300, ZN => n16704);
   U9840 : NAND2_X1 port map( A1 => n20422, A2 => n20399, ZN => n4265);
   U9841 : AOI21_X1 port map( B1 => n3667, B2 => n3666, A => n23860, ZN => 
                           n23855);
   U9842 : NAND3_X1 port map( A1 => n23851, A2 => n3183, A3 => n24428, ZN => 
                           n3666);
   U9843 : OR2_X1 port map( A1 => n23851, A2 => n3183, ZN => n3667);
   U9844 : NAND2_X1 port map( A1 => n23839, A2 => n23862, ZN => n23851);
   U9845 : OAI211_X1 port map( C1 => n5371, C2 => n4874, A => n3673, B => n3672
                           , ZN => n3671);
   U9846 : NAND2_X1 port map( A1 => n18747, A2 => n18923, ZN => n3672);
   U9847 : NAND2_X1 port map( A1 => n18748, A2 => n19315, ZN => n3673);
   U9848 : OAI21_X1 port map( B1 => n3674, B2 => n10064, A => n10060, ZN => 
                           n5609);
   U9850 : INV_X1 port map( A => n10063, ZN => n3674);
   U9851 : NAND2_X1 port map( A1 => n3676, A2 => n3675, ZN => n7493);
   U9852 : NAND2_X1 port map( A1 => n7489, A2 => n24475, ZN => n3675);
   U9853 : NAND2_X1 port map( A1 => n7947, A2 => n7942, ZN => n7489);
   U9855 : NAND2_X1 port map( A1 => n3681, A2 => n3679, ZN => n8132);
   U9856 : NAND3_X1 port map( A1 => n5015, A2 => n7754, A3 => n5202, ZN => 
                           n3680);
   U9857 : INV_X1 port map( A => n22270, ZN => n22324);
   U9860 : NAND4_X1 port map( A1 => n15920, A2 => n3685, A3 => n17366, A4 => 
                           n3684, ZN => n3683);
   U9861 : OR2_X1 port map( A1 => n17039, A2 => n25058, ZN => n3684);
   U9862 : NAND2_X1 port map( A1 => n25058, A2 => n16770, ZN => n17366);
   U9863 : AND2_X1 port map( A1 => n13164, A2 => n1353, ZN => n3686);
   U9864 : NAND2_X1 port map( A1 => n24601, A2 => n13061, ZN => n13164);
   U9866 : XNOR2_X2 port map( A => n20959, B => n20958, ZN => n22072);
   U9867 : NOR2_X1 port map( A1 => n22917, A2 => n22072, ZN => n4948);
   U9868 : INV_X1 port map( A => n12719, ZN => n3689);
   U9870 : NAND2_X1 port map( A1 => n13011, A2 => n13014, ZN => n3691);
   U9871 : NAND2_X1 port map( A1 => n19438, A2 => n361, ZN => n19246);
   U9872 : NAND2_X1 port map( A1 => n6076, A2 => n6795, ZN => n6362);
   U9875 : NAND2_X1 port map( A1 => n17370, A2 => n17369, ZN => n3693);
   U9876 : NAND2_X1 port map( A1 => n13395, A2 => n3698, ZN => n3697);
   U9877 : NAND2_X1 port map( A1 => n3700, A2 => n24995, ZN => n3699);
   U9878 : XNOR2_X1 port map( A => n12225, B => n20609, ZN => n11543);
   U9879 : XNOR2_X1 port map( A => n18301, B => n3703, ZN => n18567);
   U9880 : XNOR2_X1 port map( A => n3703, B => n18294, ZN => n16946);
   U9881 : NAND2_X1 port map( A1 => n13081, A2 => n13080, ZN => n13647);
   U9882 : NOR2_X1 port map( A1 => n13078, A2 => n24573, ZN => n3704);
   U9884 : XNOR2_X1 port map( A => n3706, B => n18233, ZN => n18613);
   U9885 : XNOR2_X1 port map( A => n14916, B => n14915, ZN => n3707);
   U9886 : INV_X1 port map( A => n16030, ZN => n4092);
   U9887 : MUX2_X1 port map( A => n16274, B => n24403, S => n16030, Z => n4091)
                           ;
   U9888 : NAND2_X1 port map( A1 => n21841, A2 => n22252, ZN => n22254);
   U9891 : NOR2_X1 port map( A1 => n17320, A2 => n4426, ZN => n16710);
   U9892 : NAND2_X1 port map( A1 => n17079, A2 => n17075, ZN => n17482);
   U9894 : NAND3_X1 port map( A1 => n22282, A2 => n3714, A3 => n2673, ZN => 
                           n3713);
   U9895 : NAND2_X1 port map( A1 => n22947, A2 => n22946, ZN => n3714);
   U9896 : XNOR2_X1 port map( A => n3715, B => n2847, ZN => n7494);
   U9897 : XNOR2_X1 port map( A => n3715, B => n889, ZN => n8996);
   U9898 : XNOR2_X1 port map( A => n3715, B => n22886, ZN => n8422);
   U9899 : XNOR2_X1 port map( A => n3715, B => n21533, ZN => n8629);
   U9900 : NAND3_X1 port map( A1 => n3717, A2 => n1028, A3 => n14150, ZN => 
                           n3892);
   U9901 : NAND2_X1 port map( A1 => n5102, A2 => n3716, ZN => n14032);
   U9902 : NAND2_X1 port map( A1 => n13805, A2 => n3717, ZN => n4962);
   U9903 : NAND2_X1 port map( A1 => n3720, A2 => n23250, ZN => n4072);
   U9904 : NOR2_X1 port map( A1 => n23236, A2 => n25373, ZN => n22648);
   U9905 : NAND3_X1 port map( A1 => n23241, A2 => n24914, A3 => n3719, ZN => 
                           n23244);
   U9906 : INV_X1 port map( A => n9220, ZN => n3722);
   U9907 : NAND2_X1 port map( A1 => n4806, A2 => n24586, ZN => n3723);
   U9908 : XNOR2_X1 port map( A => n3725, B => n921, ZN => n4873);
   U9909 : XNOR2_X1 port map( A => n18239, B => n3725, ZN => n17982);
   U9910 : XNOR2_X1 port map( A => n3725, B => n17840, ZN => n18537);
   U9911 : XNOR2_X1 port map( A => n3725, B => n18621, ZN => n17261);
   U9912 : INV_X1 port map( A => n24407, ZN => n3726);
   U9913 : AOI21_X1 port map( B1 => n3727, B2 => n3726, A => n19393, ZN => 
                           n19399);
   U9914 : NAND2_X1 port map( A1 => n25198, A2 => n13246, ZN => n12807);
   U9915 : NAND2_X1 port map( A1 => n13015, A2 => n25199, ZN => n12561);
   U9916 : NOR2_X1 port map( A1 => n10685, A2 => n4481, ZN => n11007);
   U9917 : NAND2_X1 port map( A1 => n11007, A2 => n11004, ZN => n3728);
   U9920 : NAND2_X1 port map( A1 => n3734, A2 => n3733, ZN => n3732);
   U9921 : NOR2_X1 port map( A1 => n19953, A2 => n20588, ZN => n3733);
   U9922 : INV_X1 port map( A => n20590, ZN => n3734);
   U9923 : INV_X1 port map( A => n16686, ZN => n3735);
   U9924 : NAND2_X1 port map( A1 => n16686, A2 => n25030, ZN => n3736);
   U9925 : NAND3_X1 port map( A1 => n17279, A2 => n17275, A3 => n17252, ZN => 
                           n17253);
   U9926 : OAI21_X1 port map( B1 => n16106, B2 => n16109, A => n2090, ZN => 
                           n15855);
   U9929 : XNOR2_X1 port map( A => n3738, B => n23841, ZN => Ciphertext(163));
   U9930 : NAND3_X1 port map( A1 => n3739, A2 => n4816, A3 => n23840, ZN => 
                           n3738);
   U9931 : XNOR2_X1 port map( A => n17913, B => n23602, ZN => n16947);
   U9932 : NAND2_X1 port map( A1 => n3740, A2 => n20444, ZN => n23843);
   U9933 : OAI21_X1 port map( B1 => n9340, B2 => n10148, A => n3742, ZN => 
                           n8225);
   U9934 : NOR2_X2 port map( A1 => n12578, A2 => n12579, ZN => n13843);
   U9935 : NAND3_X1 port map( A1 => n5099, A2 => n3749, A3 => n3747, ZN => 
                           n19697);
   U9936 : NAND2_X1 port map( A1 => n19325, A2 => n19472, ZN => n3747);
   U9937 : NOR2_X1 port map( A1 => n10202, A2 => n3750, ZN => n9411);
   U9938 : MUX2_X1 port map( A => n4733, B => n10752, S => n3750, Z => n4732);
   U9939 : NAND2_X1 port map( A1 => n19125, A2 => n19539, ZN => n3752);
   U9940 : INV_X1 port map( A => n14063, ZN => n3756);
   U9941 : AND2_X1 port map( A1 => n13627, A2 => n14063, ZN => n3754);
   U9942 : AOI21_X1 port map( B1 => n3760, B2 => n3761, A => n3758, ZN => n3757
                           );
   U9944 : NOR2_X1 port map( A1 => n10941, A2 => n11038, ZN => n3762);
   U9945 : NAND2_X1 port map( A1 => n6939, A2 => n5908, ZN => n3763);
   U9946 : NAND2_X1 port map( A1 => n3544, A2 => n24062, ZN => n3764);
   U9947 : NAND2_X1 port map( A1 => n11026, A2 => n3769, ZN => n3768);
   U9948 : NOR2_X1 port map( A1 => n11520, A2 => n10922, ZN => n3769);
   U9949 : NAND2_X1 port map( A1 => n3773, A2 => n19276, ZN => n3772);
   U9950 : AND2_X1 port map( A1 => n19278, A2 => n19126, ZN => n19276);
   U9952 : NAND2_X1 port map( A1 => n16371, A2 => n16616, ZN => n3774);
   U9953 : AOI21_X1 port map( B1 => n24556, B2 => n14510, A => n14439, ZN => 
                           n3776);
   U9954 : NAND2_X1 port map( A1 => n24062, A2 => n3779, ZN => n15647);
   U9955 : MUX2_X1 port map( A => n16404, B => n16202, S => n3544, Z => n15813)
                           ;
   U9956 : NAND2_X1 port map( A1 => n1130, A2 => n7230, ZN => n6982);
   U9957 : NOR2_X1 port map( A1 => n3780, A2 => n7327, ZN => n7329);
   U9958 : INV_X1 port map( A => n7232, ZN => n3780);
   U9959 : MUX2_X1 port map( A => n24543, B => n3783, S => n17312, Z => n17318)
                           ;
   U9960 : NAND2_X1 port map( A1 => n16716, A2 => n3783, ZN => n16717);
   U9961 : NAND2_X1 port map( A1 => n3785, A2 => n17410, ZN => n3784);
   U9962 : NAND2_X1 port map( A1 => n3822, A2 => n17409, ZN => n3785);
   U9963 : NOR2_X1 port map( A1 => n14165, A2 => n14167, ZN => n13466);
   U9964 : NAND2_X1 port map( A1 => n14268, A2 => n13840, ZN => n3789);
   U9966 : NAND2_X1 port map( A1 => n12739, A2 => n14436, ZN => n3792);
   U9967 : AND2_X1 port map( A1 => n20617, A2 => n20615, ZN => n3795);
   U9968 : OR2_X1 port map( A1 => n20614, A2 => n20571, ZN => n3796);
   U9969 : XNOR2_X1 port map( A => n3797, B => n8722, ZN => n8723);
   U9970 : INV_X1 port map( A => n729, ZN => n3798);
   U9971 : OAI21_X1 port map( B1 => n9978, B2 => n9986, A => n9665, ZN => n3800
                           );
   U9972 : NAND2_X1 port map( A1 => n3799, A2 => n9664, ZN => n9986);
   U9973 : INV_X1 port map( A => n9429, ZN => n3799);
   U9974 : INV_X1 port map( A => n9429, ZN => n9740);
   U9977 : NAND2_X1 port map( A1 => n21290, A2 => n21848, ZN => n3804);
   U9978 : NAND2_X1 port map( A1 => n21289, A2 => n25395, ZN => n3805);
   U9980 : NAND2_X2 port map( A1 => n11595, A2 => n11590, ZN => n13394);
   U9981 : NAND2_X1 port map( A1 => n20193, A2 => n20432, ZN => n5205);
   U9983 : NAND2_X1 port map( A1 => n19214, A2 => n19215, ZN => n3809);
   U9985 : NAND3_X1 port map( A1 => n404, A2 => n12695, A3 => n12834, ZN => 
                           n12696);
   U9986 : NAND3_X1 port map( A1 => n12964, A2 => n12963, A3 => n404, ZN => 
                           n12969);
   U9987 : NAND2_X1 port map( A1 => n7960, A2 => n437, ZN => n7964);
   U9988 : INV_X1 port map( A => n3818, ZN => n16976);
   U9990 : XNOR2_X1 port map( A => n3819, B => n21738, ZN => n20741);
   U9991 : XNOR2_X1 port map( A => n3819, B => n451, ZN => n20811);
   U9992 : XNOR2_X1 port map( A => n3819, B => n2215, ZN => n21431);
   U9993 : XNOR2_X1 port map( A => n3819, B => n21273, ZN => n20984);
   U9994 : XNOR2_X1 port map( A => n3819, B => n21633, ZN => n20679);
   U9995 : NAND3_X1 port map( A1 => n19171, A2 => n19169, A3 => n19170, ZN => 
                           n3821);
   U9996 : XNOR2_X1 port map( A => n3823, B => n20021, ZN => n20033);
   U9997 : XNOR2_X1 port map( A => n3823, B => n21160, ZN => n20551);
   U9998 : XNOR2_X1 port map( A => n3823, B => n23663, ZN => n21344);
   U9999 : XNOR2_X1 port map( A => n3823, B => n22525, ZN => n21424);
   U10001 : NAND2_X1 port map( A1 => n3828, A2 => n12854, ZN => n3826);
   U10002 : INV_X1 port map( A => n12854, ZN => n3827);
   U10003 : INV_X1 port map( A => n12853, ZN => n3828);
   U10006 : NAND2_X1 port map( A1 => n3832, A2 => n20131, ZN => n3831);
   U10007 : MUX2_X1 port map( A => n21008, B => n20522, S => n20289, Z => n3832
                           );
   U10009 : NOR2_X1 port map( A1 => n1449, A2 => n3835, ZN => n3834);
   U10010 : OAI21_X1 port map( B1 => n20126, B2 => n20125, A => n20130, ZN => 
                           n3835);
   U10011 : NAND3_X1 port map( A1 => n3837, A2 => n22727, A3 => n3836, ZN => 
                           n22730);
   U10013 : AND2_X1 port map( A1 => n6967, A2 => n6576, ZN => n3839);
   U10014 : OAI21_X1 port map( B1 => n23969, B2 => n3841, A => n3842, ZN => 
                           n3840);
   U10015 : NAND2_X1 port map( A1 => n23967, A2 => n23966, ZN => n3841);
   U10016 : NAND2_X1 port map( A1 => n22827, A2 => n23969, ZN => n3842);
   U10017 : XNOR2_X1 port map( A => n3843, B => n2126, ZN => Ciphertext(184));
   U10018 : NAND2_X1 port map( A1 => n16023, A2 => n4957, ZN => n16025);
   U10019 : OAI21_X1 port map( B1 => n18969, B2 => n18970, A => n3844, ZN => 
                           n18982);
   U10020 : OAI22_X1 port map( A1 => n19300, A2 => n19297, B1 => n18927, B2 => 
                           n19295, ZN => n18968);
   U10021 : INV_X1 port map( A => n1363, ZN => n3845);
   U10022 : NAND2_X1 port map( A1 => n13513, A2 => n14153, ZN => n13514);
   U10024 : NAND2_X1 port map( A1 => n13304, A2 => n12914, ZN => n3848);
   U10026 : INV_X1 port map( A => n14122, ZN => n3851);
   U10028 : XNOR2_X1 port map( A => n18704, B => n18701, ZN => n3852);
   U10029 : XNOR2_X1 port map( A => n18703, B => n18702, ZN => n3853);
   U10030 : NAND2_X1 port map( A1 => n3855, A2 => n17248, ZN => n3854);
   U10031 : INV_X1 port map( A => n17272, ZN => n3855);
   U10032 : OAI22_X1 port map( A1 => n335, A2 => n3856, B1 => n21826, B2 => 
                           n22252, ZN => n3890);
   U10033 : NOR2_X1 port map( A1 => n23744, A2 => n1462, ZN => n23731);
   U10034 : NAND2_X1 port map( A1 => n23735, A2 => n3857, ZN => n23737);
   U10035 : INV_X1 port map( A => n23744, ZN => n3857);
   U10036 : NAND3_X1 port map( A1 => n13311, A2 => n24487, A3 => n3859, ZN => 
                           n3858);
   U10037 : NOR2_X1 port map( A1 => n3866, A2 => n10111, ZN => n3863);
   U10038 : NAND2_X1 port map( A1 => n3865, A2 => n8644, ZN => n3864);
   U10039 : AOI21_X1 port map( B1 => n10107, B2 => n10106, A => n8644, ZN => 
                           n3866);
   U10041 : NAND3_X1 port map( A1 => n3868, A2 => n11214, A3 => n233, ZN => 
                           n3867);
   U10042 : NAND3_X1 port map( A1 => n24340, A2 => n10810, A3 => n11212, ZN => 
                           n3869);
   U10043 : NAND3_X1 port map( A1 => n25082, A2 => n245, A3 => n22356, ZN => 
                           n4203);
   U10044 : INV_X1 port map( A => n17341, ZN => n17347);
   U10045 : NAND3_X1 port map( A1 => n24307, A2 => n24895, A3 => n22043, ZN => 
                           n3878);
   U10046 : OAI21_X1 port map( B1 => n3876, B2 => n12673, A => n13661, ZN => 
                           n3873);
   U10048 : NAND2_X1 port map( A1 => n13111, A2 => n4923, ZN => n3874);
   U10049 : NAND2_X1 port map( A1 => n3876, A2 => n13107, ZN => n3875);
   U10050 : INV_X1 port map( A => n13110, ZN => n3876);
   U10051 : XNOR2_X1 port map( A => n3877, B => n22049, ZN => Ciphertext(150));
   U10052 : NAND3_X1 port map( A1 => n3879, A2 => n22048, A3 => n3878, ZN => 
                           n3877);
   U10053 : OAI21_X1 port map( B1 => n22047, B2 => n24307, A => n3880, ZN => 
                           n3879);
   U10054 : NAND2_X1 port map( A1 => n24307, A2 => n24983, ZN => n3880);
   U10055 : XNOR2_X1 port map( A => n11798, B => n3881, ZN => n12126);
   U10058 : INV_X1 port map( A => n14200, ZN => n3887);
   U10060 : NAND2_X1 port map( A1 => n3886, A2 => n3888, ZN => n3885);
   U10061 : NOR2_X1 port map( A1 => n14945, A2 => n3887, ZN => n3886);
   U10062 : INV_X1 port map( A => n14200, ZN => n3889);
   U10064 : NAND2_X1 port map( A1 => n3893, A2 => n3892, ZN => n3891);
   U10065 : INV_X1 port map( A => n3894, ZN => n5832);
   U10066 : NAND2_X1 port map( A1 => n3894, A2 => n6791, ZN => n6798);
   U10067 : NAND2_X1 port map( A1 => n24362, A2 => n332, ZN => n3895);
   U10068 : NAND2_X1 port map( A1 => n21840, A2 => n22257, ZN => n3896);
   U10071 : NAND2_X1 port map( A1 => n7881, A2 => n7884, ZN => n3898);
   U10073 : NAND2_X1 port map( A1 => n3904, A2 => n341, ZN => n3903);
   U10074 : MUX2_X1 port map( A => n18994, B => n20319, S => n19889, Z => n3904
                           );
   U10076 : INV_X1 port map( A => n22465, ZN => n21929);
   U10077 : XNOR2_X2 port map( A => n20814, B => n20813, ZN => n22465);
   U10078 : NAND2_X1 port map( A1 => n3907, A2 => n3906, ZN => n21377);
   U10080 : NAND2_X1 port map( A1 => n22463, A2 => n1363, ZN => n22329);
   U10083 : NAND2_X1 port map( A1 => n23042, A2 => n23048, ZN => n3910);
   U10084 : INV_X1 port map( A => n23048, ZN => n23059);
   U10087 : NOR2_X1 port map( A1 => n20602, A2 => n3916, ZN => n19848);
   U10088 : AND2_X1 port map( A1 => n25476, A2 => n20597, ZN => n3916);
   U10089 : INV_X1 port map( A => n19615, ZN => n3919);
   U10090 : INV_X1 port map( A => n7380, ZN => n7386);
   U10091 : NAND2_X1 port map( A1 => n5656, A2 => n3923, ZN => n3920);
   U10092 : XNOR2_X1 port map( A => n18605, B => n896, ZN => n17504);
   U10093 : AND2_X2 port map( A1 => n3928, A2 => n3927, ZN => n18605);
   U10094 : NAND2_X1 port map( A1 => n16519, A2 => n17139, ZN => n3927);
   U10095 : XNOR2_X1 port map( A => n15482, B => n15481, ZN => n3931);
   U10096 : NAND2_X1 port map( A1 => n3933, A2 => n20591, ZN => n3932);
   U10099 : NOR2_X1 port map( A1 => n22465, A2 => n3938, ZN => n3937);
   U10100 : INV_X1 port map( A => n22464, ZN => n22461);
   U10101 : NAND3_X1 port map( A1 => n22459, A2 => n3845, A3 => n22464, ZN => 
                           n3939);
   U10102 : XNOR2_X1 port map( A => n15431, B => n14805, ZN => n15268);
   U10103 : XNOR2_X1 port map( A => n3941, B => n3940, ZN => n3942);
   U10104 : XNOR2_X1 port map( A => n15410, B => n15431, ZN => n3941);
   U10105 : XNOR2_X2 port map( A => n3942, B => n13393, ZN => n15667);
   U10106 : OAI21_X1 port map( B1 => n12853, B2 => n3945, A => n3944, ZN => 
                           n13663);
   U10107 : NAND2_X1 port map( A1 => n12673, A2 => n12856, ZN => n3944);
   U10108 : OR2_X1 port map( A1 => n12672, A2 => n12856, ZN => n3945);
   U10109 : NAND2_X1 port map( A1 => n25455, A2 => n15667, ZN => n15670);
   U10111 : OAI21_X1 port map( B1 => n267, B2 => n3947, A => n3946, ZN => 
                           n15669);
   U10112 : NAND2_X1 port map( A1 => n267, A2 => n25455, ZN => n3946);
   U10113 : INV_X1 port map( A => n15667, ZN => n3947);
   U10114 : INV_X1 port map( A => n17039, ZN => n3950);
   U10115 : NAND2_X1 port map( A1 => n3955, A2 => n25215, ZN => n3948);
   U10116 : NAND2_X1 port map( A1 => n3950, A2 => n25058, ZN => n3949);
   U10117 : NAND2_X1 port map( A1 => n17037, A2 => n3951, ZN => n3956);
   U10118 : NAND2_X1 port map( A1 => n3953, A2 => n3952, ZN => n18023);
   U10119 : NAND2_X1 port map( A1 => n3956, A2 => n370, ZN => n3952);
   U10120 : XNOR2_X2 port map( A => n10988, B => n10987, ZN => n3958);
   U10121 : NAND2_X1 port map( A1 => n3958, A2 => n13102, ZN => n12511);
   U10122 : NAND2_X1 port map( A1 => n12742, A2 => n3958, ZN => n13104);
   U10123 : NAND2_X1 port map( A1 => n12744, A2 => n3958, ZN => n12741);
   U10124 : MUX2_X1 port map( A => n13187, B => n3958, S => n13102, Z => n11020
                           );
   U10125 : OR2_X1 port map( A1 => n13191, A2 => n3958, ZN => n3957);
   U10126 : OAI22_X1 port map( A1 => n2321, A2 => n13609, B1 => n14090, B2 => 
                           n3959, ZN => n13542);
   U10127 : OAI21_X2 port map( B1 => n22143, B2 => n22142, A => n3960, ZN => 
                           n23275);
   U10128 : NAND2_X1 port map( A1 => n3961, A2 => n22274, ZN => n3960);
   U10129 : INV_X1 port map( A => n19784, ZN => n21068);
   U10130 : OAI21_X1 port map( B1 => n24588, B2 => n3966, A => n3965, ZN => 
                           n3964);
   U10131 : NAND2_X1 port map( A1 => n24588, A2 => n13888, ZN => n3965);
   U10132 : NAND3_X1 port map( A1 => n9919, A2 => n9914, A3 => n9920, ZN => 
                           n9274);
   U10134 : NAND2_X1 port map( A1 => n13062, A2 => n12439, ZN => n3970);
   U10135 : MUX2_X1 port map( A => n12454, B => n1353, S => n13061, Z => n3971)
                           ;
   U10136 : NAND2_X1 port map( A1 => n3973, A2 => n12459, ZN => n3972);
   U10137 : NAND2_X1 port map( A1 => n12460, A2 => n12652, ZN => n3973);
   U10138 : NAND2_X1 port map( A1 => n16741, A2 => n16742, ZN => n3976);
   U10139 : NAND2_X1 port map( A1 => n17090, A2 => n16740, ZN => n3977);
   U10140 : INV_X1 port map( A => n16649, ZN => n17085);
   U10142 : NAND2_X1 port map( A1 => n4947, A2 => n4949, ZN => n3978);
   U10143 : NAND3_X1 port map( A1 => n3978, A2 => n22920, A3 => n23018, ZN => 
                           n5465);
   U10144 : NAND2_X1 port map( A1 => n3979, A2 => n24878, ZN => n7268);
   U10145 : MUX2_X1 port map( A => n3979, B => n24878, S => n8370, Z => n7840);
   U10148 : NAND2_X1 port map( A1 => n3982, A2 => n5072, ZN => n3981);
   U10149 : INV_X1 port map( A => n19245, ZN => n3986);
   U10151 : XNOR2_X1 port map( A => n3990, B => n18435, ZN => n18620);
   U10152 : NAND2_X1 port map( A1 => n10954, A2 => n10548, ZN => n10958);
   U10153 : OAI21_X1 port map( B1 => n3996, B2 => n3995, A => n3994, ZN => 
                           n19730);
   U10154 : NAND2_X1 port map( A1 => n363, A2 => n18340, ZN => n3994);
   U10155 : NAND2_X1 port map( A1 => n3997, A2 => n24446, ZN => n9086);
   U10156 : INV_X1 port map( A => n4096, ZN => n3997);
   U10157 : OAI21_X1 port map( B1 => n4096, B2 => n10058, A => n3998, ZN => 
                           n9691);
   U10158 : NOR3_X1 port map( A1 => n24921, A2 => n23752, A3 => n4000, ZN => 
                           n22524);
   U10159 : INV_X1 port map( A => n7481, ZN => n7575);
   U10160 : MUX2_X1 port map( A => n7577, B => n7573, S => n7481, Z => n4002);
   U10162 : NAND3_X1 port map( A1 => n17012, A2 => n17356, A3 => n4004, ZN => 
                           n4003);
   U10163 : NAND4_X2 port map( A1 => n4007, A2 => n19378, A3 => n4006, A4 => 
                           n4008, ZN => n20459);
   U10164 : NAND3_X1 port map( A1 => n19377, A2 => n25067, A3 => n18876, ZN => 
                           n4006);
   U10165 : NAND2_X1 port map( A1 => n4010, A2 => n20022, ZN => n4009);
   U10166 : NAND2_X1 port map( A1 => n19727, A2 => n19728, ZN => n4010);
   U10167 : NAND2_X1 port map( A1 => n4012, A2 => n4011, ZN => n10837);
   U10168 : NAND2_X1 port map( A1 => n10829, A2 => n4013, ZN => n4011);
   U10169 : NAND2_X1 port map( A1 => n10830, A2 => n10518, ZN => n4012);
   U10170 : NAND3_X1 port map( A1 => n10829, A2 => n10275, A3 => n4013, ZN => 
                           n10193);
   U10171 : NAND3_X1 port map( A1 => n13728, A2 => n24588, A3 => n13945, ZN => 
                           n4014);
   U10172 : NAND2_X1 port map( A1 => n13909, A2 => n13951, ZN => n4016);
   U10175 : NAND2_X1 port map( A1 => n14218, A2 => n4019, ZN => n13400);
   U10176 : MUX2_X1 port map( A => n14218, B => n4019, S => n14219, Z => n14121
                           );
   U10177 : NAND2_X1 port map( A1 => n4020, A2 => n21046, ZN => n4022);
   U10178 : NAND2_X1 port map( A1 => n4022, A2 => n4021, ZN => n4025);
   U10179 : NAND3_X1 port map( A1 => n5162, A2 => n7237, A3 => n4023, ZN => 
                           n4021);
   U10180 : NAND3_X1 port map( A1 => n16175, A2 => n4027, A3 => n4026, ZN => 
                           n16180);
   U10181 : NAND2_X1 port map( A1 => n15655, A2 => n15656, ZN => n4027);
   U10182 : OR2_X1 port map( A1 => n15993, A2 => n4027, ZN => n4645);
   U10183 : OR2_X1 port map( A1 => n22529, A2 => n4034, ZN => n4031);
   U10184 : OAI211_X1 port map( C1 => n4031, C2 => n4030, A => n4029, B => 
                           n4028, ZN => Ciphertext(93));
   U10185 : NAND2_X1 port map( A1 => n22529, A2 => n4034, ZN => n4028);
   U10186 : INV_X1 port map( A => n4032, ZN => n4030);
   U10187 : NAND3_X1 port map( A1 => n4033, A2 => n3242, A3 => n23437, ZN => 
                           n4032);
   U10188 : NAND2_X1 port map( A1 => n285, A2 => n25003, ZN => n4037);
   U10189 : INV_X1 port map( A => n17840, ZN => n17726);
   U10190 : NAND2_X1 port map( A1 => n4038, A2 => n285, ZN => n4035);
   U10191 : NAND3_X1 port map( A1 => n4037, A2 => n16661, A3 => n17399, ZN => 
                           n4036);
   U10192 : NAND2_X1 port map( A1 => n20437, A2 => n20194, ZN => n5209);
   U10193 : INV_X1 port map( A => n10445, ZN => n10905);
   U10194 : NAND2_X1 port map( A1 => n13266, A2 => n24443, ZN => n13268);
   U10195 : OAI21_X1 port map( B1 => n12932, B2 => n25015, A => n24443, ZN => 
                           n12933);
   U10198 : AOI22_X1 port map( A1 => n6480, A2 => n4042, B1 => n6479, B2 => 
                           n6924, ZN => n6482);
   U10199 : NAND2_X1 port map( A1 => n4043, A2 => n14130, ZN => n13410);
   U10200 : INV_X1 port map( A => n15656, ZN => n4045);
   U10201 : NAND2_X1 port map( A1 => n15839, A2 => n15655, ZN => n4044);
   U10202 : OAI21_X1 port map( B1 => n10630, B2 => n11201, A => n4047, ZN => 
                           n4050);
   U10204 : NAND2_X1 port map( A1 => n4050, A2 => n11195, ZN => n4048);
   U10205 : XNOR2_X1 port map( A => n8520, B => n4138, ZN => n9500);
   U10206 : NAND2_X1 port map( A1 => n10003, A2 => n9668, ZN => n9670);
   U10207 : OR2_X1 port map( A1 => n9500, A2 => n1796, ZN => n10003);
   U10208 : OAI22_X1 port map( A1 => n19252, A2 => n4052, B1 => n5134, B2 => 
                           n19250, ZN => n4549);
   U10209 : INV_X1 port map( A => n19587, ZN => n4052);
   U10210 : NAND2_X1 port map( A1 => n25480, A2 => n6198, ZN => n4053);
   U10212 : NAND3_X1 port map( A1 => n25446, A2 => n15694, A3 => n16063, ZN => 
                           n4054);
   U10213 : INV_X1 port map( A => n12482, ZN => n4061);
   U10214 : NAND2_X1 port map( A1 => n4055, A2 => n4057, ZN => n13636);
   U10215 : NAND2_X1 port map( A1 => n4058, A2 => n4056, ZN => n4055);
   U10216 : NAND2_X1 port map( A1 => n12482, A2 => n24573, ZN => n4056);
   U10217 : NAND2_X1 port map( A1 => n12483, A2 => n12710, ZN => n4060);
   U10218 : NAND2_X1 port map( A1 => n11024, A2 => n11518, ZN => n11522);
   U10219 : NAND2_X1 port map( A1 => n24902, A2 => n22166, ZN => n4062);
   U10221 : NOR2_X1 port map( A1 => n4064, A2 => n22166, ZN => n4063);
   U10222 : NAND3_X1 port map( A1 => n22117, A2 => n22170, A3 => n4064, ZN => 
                           n22118);
   U10223 : INV_X1 port map( A => n20480, ZN => n4065);
   U10226 : NOR2_X1 port map( A1 => n20296, A2 => n4066, ZN => n19047);
   U10227 : OAI21_X1 port map( B1 => n20298, B2 => n4066, A => n20140, ZN => 
                           n19035);
   U10228 : AOI21_X1 port map( B1 => n20296, B2 => n4066, A => n20142, ZN => 
                           n20143);
   U10229 : NAND3_X1 port map( A1 => n10048, A2 => n10046, A3 => n4069, ZN => 
                           n4068);
   U10230 : INV_X1 port map( A => n8977, ZN => n4070);
   U10231 : NAND2_X1 port map( A1 => n22298, A2 => n4072, ZN => n4071);
   U10232 : NAND2_X1 port map( A1 => n24914, A2 => n23251, ZN => n22298);
   U10234 : NAND2_X1 port map( A1 => n4075, A2 => n19296, ZN => n4077);
   U10236 : INV_X1 port map( A => n19295, ZN => n4075);
   U10237 : NAND2_X1 port map( A1 => n4077, A2 => n18970, ZN => n4076);
   U10238 : NAND2_X1 port map( A1 => n6924, A2 => n4078, ZN => n6779);
   U10240 : NAND3_X1 port map( A1 => n24953, A2 => n4081, A3 => n4080, ZN => 
                           n4079);
   U10241 : NAND2_X1 port map( A1 => n17465, A2 => n25572, ZN => n4082);
   U10242 : NOR2_X1 port map( A1 => n16021, A2 => n287, ZN => n4083);
   U10243 : XNOR2_X1 port map( A => n18197, B => n17959, ZN => n18692);
   U10244 : AND2_X2 port map( A1 => n4084, A2 => n1492, ZN => n18197);
   U10245 : OAI21_X1 port map( B1 => n16988, B2 => n4085, A => n5763, ZN => 
                           n4084);
   U10246 : INV_X1 port map( A => n17363, ZN => n4085);
   U10248 : XNOR2_X1 port map( A => n18044, B => n4087, ZN => n4086);
   U10249 : XNOR2_X1 port map( A => n18285, B => n18562, ZN => n4087);
   U10250 : INV_X1 port map( A => n11003, ZN => n4088);
   U10251 : NAND2_X1 port map( A1 => n10681, A2 => n10682, ZN => n11003);
   U10254 : NAND2_X1 port map( A1 => n10558, A2 => n10660, ZN => n10397);
   U10255 : NAND2_X1 port map( A1 => n13235, A2 => n12902, ZN => n4490);
   U10256 : NAND3_X1 port map( A1 => n24403, A2 => n15572, A3 => n4092, ZN => 
                           n4090);
   U10257 : INV_X1 port map( A => n7657, ZN => n4093);
   U10258 : INV_X1 port map( A => n12490, ZN => n4094);
   U10259 : XNOR2_X1 port map( A => n4095, B => n15016, ZN => n14387);
   U10260 : NAND2_X1 port map( A1 => n12649, A2 => n4405, ZN => n12179);
   U10261 : OAI21_X1 port map( B1 => n5323, B2 => n4405, A => n13094, ZN => 
                           n12870);
   U10262 : AND2_X1 port map( A1 => n10053, A2 => n4096, ZN => n10051);
   U10263 : NAND2_X1 port map( A1 => n2902, A2 => n9866, ZN => n9247);
   U10265 : XNOR2_X1 port map( A => n20677, B => n20679, ZN => n4101);
   U10266 : NAND2_X1 port map( A1 => n20684, A2 => n4109, ZN => n4102);
   U10268 : INV_X1 port map( A => n22389, ZN => n4098);
   U10269 : NAND2_X1 port map( A1 => n4372, A2 => n22387, ZN => n4099);
   U10271 : OAI211_X2 port map( C1 => n19426, C2 => n19177, A => n18598, B => 
                           n4103, ZN => n20615);
   U10272 : NAND2_X1 port map( A1 => n4104, A2 => n19427, ZN => n4103);
   U10273 : OAI21_X1 port map( B1 => n19177, B2 => n18597, A => n1361, ZN => 
                           n4104);
   U10274 : NAND2_X1 port map( A1 => n5495, A2 => n5493, ZN => n16549);
   U10275 : NAND2_X1 port map( A1 => n6924, A2 => n6775, ZN => n4106);
   U10276 : INV_X1 port map( A => n6292, ZN => n6924);
   U10277 : XNOR2_X1 port map( A => n24027, B => n8761, ZN => n11447);
   U10278 : XNOR2_X1 port map( A => n24027, B => n4107, ZN => n11321);
   U10279 : NAND2_X1 port map( A1 => n13935, A2 => n14245, ZN => n13932);
   U10281 : AND2_X1 port map( A1 => n23320, A2 => n4108, ZN => n22628);
   U10282 : NAND2_X1 port map( A1 => n19948, A2 => n20460, ZN => n4110);
   U10283 : INV_X1 port map( A => n20394, ZN => n19948);
   U10284 : NAND4_X1 port map( A1 => n4113, A2 => n23193, A3 => n23202, A4 => 
                           n2903, ZN => n4112);
   U10285 : NAND2_X1 port map( A1 => n19376, A2 => n25010, ZN => n17803);
   U10287 : NAND2_X1 port map( A1 => n25128, A2 => n14241, ZN => n4118);
   U10290 : NAND2_X1 port map( A1 => n10159, A2 => n10162, ZN => n4120);
   U10291 : NOR2_X1 port map( A1 => n7734, A2 => n7642, ZN => n5594);
   U10293 : NAND2_X1 port map( A1 => n6600, A2 => n6824, ZN => n4121);
   U10294 : OR2_X1 port map( A1 => n2793, A2 => n13030, ZN => n4124);
   U10295 : OR2_X2 port map( A1 => n5786, A2 => n5785, ZN => n7580);
   U10297 : NOR2_X1 port map( A1 => n23359, A2 => n22961, ZN => n23355);
   U10299 : NAND2_X1 port map( A1 => n22956, A2 => n4128, ZN => n4126);
   U10300 : NAND2_X1 port map( A1 => n22955, A2 => n22954, ZN => n4127);
   U10301 : INV_X1 port map( A => n22954, ZN => n4128);
   U10302 : NAND2_X1 port map( A1 => n4844, A2 => n4130, ZN => n4129);
   U10303 : NAND2_X1 port map( A1 => n14130, A2 => n13895, ZN => n4130);
   U10304 : NAND2_X1 port map( A1 => n13826, A2 => n4132, ZN => n4131);
   U10305 : NAND2_X1 port map( A1 => n4133, A2 => n1331, ZN => n4132);
   U10306 : INV_X1 port map( A => n14127, ZN => n4133);
   U10307 : NAND2_X1 port map( A1 => n12885, A2 => n13223, ZN => n12918);
   U10308 : XNOR2_X1 port map( A => n12400, B => n11757, ZN => n4134);
   U10309 : XNOR2_X1 port map( A => n11740, B => n11739, ZN => n11755);
   U10310 : INV_X1 port map( A => n19210, ZN => n4135);
   U10311 : NAND3_X1 port map( A1 => n9797, A2 => n9796, A3 => n4137, ZN => 
                           n9801);
   U10312 : NAND2_X1 port map( A1 => n9795, A2 => n4137, ZN => n10002);
   U10313 : NAND2_X1 port map( A1 => n9314, A2 => n4137, ZN => n9312);
   U10314 : NAND2_X1 port map( A1 => n19607, A2 => n4139, ZN => n18864);
   U10315 : NAND2_X1 port map( A1 => n4143, A2 => n11099, ZN => n4142);
   U10316 : XNOR2_X2 port map( A => n14813, B => n14812, ZN => n16232);
   U10317 : NAND2_X1 port map( A1 => n7476, A2 => n7423, ZN => n4145);
   U10318 : XNOR2_X1 port map( A => n4146, B => n8084, ZN => n8416);
   U10319 : INV_X1 port map( A => n8411, ZN => n4146);
   U10320 : XNOR2_X1 port map( A => n4147, B => n8084, ZN => n8750);
   U10321 : INV_X1 port map( A => n8745, ZN => n4147);
   U10322 : NAND2_X1 port map( A1 => n4148, A2 => n6659, ZN => n7155);
   U10323 : NAND3_X1 port map( A1 => n4150, A2 => n4151, A3 => n4149, ZN => 
                           n4148);
   U10324 : NAND2_X1 port map( A1 => n6657, A2 => n6072, ZN => n4151);
   U10325 : NOR2_X1 port map( A1 => n11338, A2 => n25025, ZN => n4152);
   U10328 : XNOR2_X1 port map( A => n16799, B => n4153, ZN => n17328);
   U10329 : XNOR2_X1 port map( A => n4154, B => n16799, ZN => n18076);
   U10330 : INV_X1 port map( A => n18096, ZN => n4154);
   U10331 : XNOR2_X1 port map( A => n18700, B => n4155, ZN => n18702);
   U10332 : INV_X1 port map( A => n16799, ZN => n4155);
   U10335 : OAI211_X1 port map( C1 => n11214, C2 => n233, A => n10810, B => 
                           n11215, ZN => n4156);
   U10336 : INV_X1 port map( A => n11216, ZN => n10810);
   U10337 : XNOR2_X1 port map( A => n4157, B => n21537, ZN => n21539);
   U10338 : XNOR2_X1 port map( A => n21535, B => n4158, ZN => n4157);
   U10339 : NAND2_X1 port map( A1 => n4161, A2 => n4160, ZN => n4159);
   U10340 : INV_X1 port map( A => n19973, ZN => n4160);
   U10341 : NOR2_X1 port map( A1 => n19974, A2 => n4164, ZN => n4161);
   U10342 : NAND2_X1 port map( A1 => n19973, A2 => n4164, ZN => n4162);
   U10343 : NAND2_X1 port map( A1 => n19974, A2 => n4164, ZN => n4163);
   U10344 : XNOR2_X1 port map( A => n18334, B => n4761, ZN => n18615);
   U10345 : NAND2_X1 port map( A1 => n17089, A2 => n17088, ZN => n4165);
   U10346 : NAND3_X1 port map( A1 => n262, A2 => n9468, A3 => n9281, ZN => 
                           n4166);
   U10349 : NAND2_X1 port map( A1 => n19235, A2 => n19237, ZN => n4167);
   U10350 : NAND2_X1 port map( A1 => n19235, A2 => n19112, ZN => n18869);
   U10351 : NAND2_X1 port map( A1 => n1428, A2 => n4168, ZN => n4282);
   U10352 : NAND2_X1 port map( A1 => n23372, A2 => n24412, ZN => n4171);
   U10353 : NAND2_X1 port map( A1 => n4170, A2 => n4632, ZN => n4633);
   U10354 : NAND2_X1 port map( A1 => n4171, A2 => n24404, ZN => n22993);
   U10355 : NAND2_X1 port map( A1 => n22610, A2 => n22611, ZN => n23048);
   U10356 : INV_X1 port map( A => n18761, ZN => n4172);
   U10357 : NAND2_X1 port map( A1 => n4172, A2 => n24329, ZN => n17554);
   U10358 : XNOR2_X1 port map( A => n21729, B => n1854, ZN => n20733);
   U10359 : NAND4_X2 port map( A1 => n4174, A2 => n19692, A3 => n19693, A4 => 
                           n4173, ZN => n21729);
   U10360 : NAND3_X1 port map( A1 => n20322, A2 => n24917, A3 => n19889, ZN => 
                           n4173);
   U10362 : NAND2_X1 port map( A1 => n1327, A2 => n24460, ZN => n4175);
   U10363 : NAND3_X1 port map( A1 => n19948, A2 => n20460, A3 => n20395, ZN => 
                           n4176);
   U10364 : NAND2_X1 port map( A1 => n4177, A2 => n6395, ZN => n6399);
   U10366 : OAI21_X1 port map( B1 => n13172, B2 => n13171, A => n13170, ZN => 
                           n4179);
   U10367 : XNOR2_X1 port map( A => n8988, B => n9041, ZN => n8621);
   U10368 : XNOR2_X1 port map( A => n4180, B => n9041, ZN => n8287);
   U10369 : INV_X1 port map( A => n8498, ZN => n4180);
   U10370 : XNOR2_X1 port map( A => n12269, B => n12270, ZN => n4182);
   U10371 : NAND2_X1 port map( A1 => n20413, A2 => n20264, ZN => n4184);
   U10372 : INV_X1 port map( A => n4190, ZN => n4193);
   U10373 : OR2_X1 port map( A1 => n23867, A2 => n4189, ZN => n4187);
   U10374 : NAND4_X1 port map( A1 => n4191, A2 => n23867, A3 => n4190, A4 => 
                           n4189, ZN => n4188);
   U10375 : INV_X1 port map( A => n4192, ZN => n4191);
   U10376 : NAND2_X1 port map( A1 => n20476, A2 => n20353, ZN => n20354);
   U10377 : OR2_X1 port map( A1 => n19420, A2 => n19418, ZN => n4195);
   U10378 : NAND2_X1 port map( A1 => n4196, A2 => n13110, ZN => n12632);
   U10379 : NAND2_X1 port map( A1 => n4196, A2 => n13108, ZN => n4924);
   U10380 : NAND2_X1 port map( A1 => n5211, A2 => n16404, ZN => n4197);
   U10381 : MUX2_X1 port map( A => n16956, B => n17414, S => n17413, Z => 
                           n14353);
   U10382 : NAND2_X1 port map( A1 => n4198, A2 => n25572, ZN => n16506);
   U10383 : INV_X1 port map( A => n13281, ZN => n12698);
   U10384 : NAND2_X1 port map( A1 => n4202, A2 => n4201, ZN => n4200);
   U10385 : NAND3_X1 port map( A1 => n14191, A2 => n14189, A3 => n14142, ZN => 
                           n4201);
   U10386 : NOR2_X1 port map( A1 => n8023, A2 => n8022, ZN => n4206);
   U10387 : NAND3_X1 port map( A1 => n4209, A2 => n9506, A3 => n4208, ZN => 
                           n4207);
   U10388 : NAND2_X1 port map( A1 => n10088, A2 => n9507, ZN => n4209);
   U10389 : NAND2_X1 port map( A1 => n24575, A2 => n9786, ZN => n4210);
   U10390 : NAND2_X1 port map( A1 => n10508, A2 => n10931, ZN => n10425);
   U10391 : NAND4_X1 port map( A1 => n4216, A2 => n4217, A3 => n4218, A4 => 
                           n21357, ZN => n4215);
   U10392 : NAND2_X1 port map( A1 => n21351, A2 => n21352, ZN => n4217);
   U10393 : AND2_X1 port map( A1 => n21350, A2 => n21349, ZN => n4218);
   U10394 : NAND2_X1 port map( A1 => n4221, A2 => n21844, ZN => n4219);
   U10396 : OAI211_X2 port map( C1 => n14060, C2 => n14415, A => n4224, B => 
                           n4222, ZN => n15133);
   U10398 : NAND3_X1 port map( A1 => n4225, A2 => n14849, A3 => n14415, ZN => 
                           n4224);
   U10399 : OAI211_X2 port map( C1 => n13263, C2 => n13484, A => n4226, B => 
                           n1407, ZN => n15062);
   U10400 : XNOR2_X1 port map( A => n4227, B => n20982, ZN => n21430);
   U10401 : XNOR2_X1 port map( A => n4227, B => n889, ZN => n20847);
   U10402 : XNOR2_X1 port map( A => n4227, B => n21630, ZN => n21631);
   U10403 : XNOR2_X1 port map( A => n4227, B => n4294, ZN => n20700);
   U10406 : NAND2_X1 port map( A1 => n4234, A2 => n4236, ZN => n4231);
   U10407 : NOR2_X1 port map( A1 => n20520, A2 => n20515, ZN => n19797);
   U10408 : NAND4_X2 port map( A1 => n4239, A2 => n19111, A3 => n4238, A4 => 
                           n4977, ZN => n20272);
   U10409 : NAND2_X1 port map( A1 => n19110, A2 => n24908, ZN => n4238);
   U10410 : NAND2_X1 port map( A1 => n19108, A2 => n19384, ZN => n4239);
   U10411 : NAND2_X1 port map( A1 => n12688, A2 => n13318, ZN => n4240);
   U10412 : OAI21_X1 port map( B1 => n12946, B2 => n13318, A => n4240, ZN => 
                           n12582);
   U10413 : NOR2_X1 port map( A1 => n4241, A2 => n13318, ZN => n12944);
   U10414 : NAND2_X1 port map( A1 => n13317, A2 => n4241, ZN => n12687);
   U10415 : XNOR2_X1 port map( A => n15504, B => n15503, ZN => n15511);
   U10416 : XNOR2_X1 port map( A => n4242, B => n23257, ZN => Ciphertext(47));
   U10417 : OAI211_X1 port map( C1 => n23256, C2 => n23255, A => n4244, B => 
                           n4243, ZN => n4242);
   U10418 : NAND2_X1 port map( A1 => n23256, A2 => n23254, ZN => n4244);
   U10419 : NOR2_X2 port map( A1 => n22287, A2 => n22286, ZN => n23256);
   U10421 : OAI21_X1 port map( B1 => n16269, B2 => n24366, A => n4249, ZN => 
                           n15162);
   U10422 : XNOR2_X1 port map( A => n4250, B => n18289, ZN => n18086);
   U10423 : XNOR2_X1 port map( A => n4250, B => n18190, ZN => n17788);
   U10424 : XNOR2_X1 port map( A => n4250, B => n20609, ZN => n18228);
   U10425 : XNOR2_X1 port map( A => n4250, B => n3158, ZN => n18638);
   U10426 : XNOR2_X1 port map( A => n4250, B => n21711, ZN => n18414);
   U10427 : XNOR2_X1 port map( A => n4250, B => n17851, ZN => n17852);
   U10428 : NAND2_X1 port map( A1 => n11058, A2 => n11057, ZN => n4251);
   U10429 : NAND2_X1 port map( A1 => n9808, A2 => n9809, ZN => n4252);
   U10430 : NAND2_X1 port map( A1 => n9776, A2 => n4254, ZN => n4253);
   U10431 : AOI21_X1 port map( B1 => n9836, B2 => n428, A => n4257, ZN => n9840
                           );
   U10432 : AND2_X1 port map( A1 => n8359, A2 => n10094, ZN => n4257);
   U10434 : NAND2_X1 port map( A1 => n9515, A2 => n9837, ZN => n4258);
   U10435 : OAI21_X1 port map( B1 => n9514, B2 => n428, A => n10097, ZN => 
                           n9518);
   U10436 : INV_X1 port map( A => n7948, ZN => n4259);
   U10437 : OAI211_X2 port map( C1 => n19289, C2 => n25448, A => n4261, B => 
                           n4260, ZN => n20419);
   U10438 : INV_X1 port map( A => n19559, ZN => n4262);
   U10439 : XNOR2_X1 port map( A => n21227, B => n4263, ZN => n22004);
   U10440 : XNOR2_X1 port map( A => n21231, B => n4263, ZN => n21233);
   U10441 : XNOR2_X1 port map( A => n24485, B => n4263, ZN => n21270);
   U10442 : XNOR2_X1 port map( A => n4263, B => n1935, ZN => n21544);
   U10443 : NAND2_X1 port map( A1 => n17054, A2 => n25031, ZN => n4266);
   U10444 : NAND2_X1 port map( A1 => n16609, A2 => n16722, ZN => n4267);
   U10445 : NOR2_X1 port map( A1 => n16001, A2 => n16266, ZN => n4270);
   U10446 : NAND2_X1 port map( A1 => n5447, A2 => n16266, ZN => n16272);
   U10447 : NAND2_X1 port map( A1 => n24385, A2 => n17059, ZN => n16722);
   U10450 : NOR2_X1 port map( A1 => n22657, A2 => n4273, ZN => n22363);
   U10452 : NAND2_X1 port map( A1 => n20442, A2 => n4273, ZN => n20443);
   U10453 : AND2_X1 port map( A1 => n22657, A2 => n4273, ZN => n4272);
   U10454 : OAI21_X1 port map( B1 => n1457, B2 => n22609, A => n4273, ZN => 
                           n4283);
   U10456 : NAND2_X1 port map( A1 => n4276, A2 => n20669, ZN => n20340);
   U10457 : OAI21_X1 port map( B1 => n20338, B2 => n20666, A => n20671, ZN => 
                           n4276);
   U10459 : INV_X1 port map( A => n7989, ZN => n7826);
   U10460 : NAND3_X1 port map( A1 => n7827, A2 => n7982, A3 => n7826, ZN => 
                           n4277);
   U10461 : NAND3_X1 port map( A1 => n7828, A2 => n7989, A3 => n7825, ZN => 
                           n4278);
   U10465 : OAI21_X2 port map( B1 => n22815, B2 => n22816, A => n22814, ZN => 
                           n24011);
   U10466 : NAND3_X1 port map( A1 => n4281, A2 => n24753, A3 => n11101, ZN => 
                           n11103);
   U10467 : NAND2_X1 port map( A1 => n4286, A2 => n17069, ZN => n17070);
   U10468 : NAND2_X1 port map( A1 => n17944, A2 => n4290, ZN => n4289);
   U10469 : OR2_X1 port map( A1 => n19327, A2 => n4291, ZN => n4290);
   U10470 : OAI21_X1 port map( B1 => n20666, B2 => n20670, A => n4292, ZN => 
                           n20351);
   U10471 : NAND2_X1 port map( A1 => n20336, A2 => n20668, ZN => n4292);
   U10472 : OAI21_X2 port map( B1 => n17310, B2 => n18933, A => n17309, ZN => 
                           n20668);
   U10473 : AOI22_X2 port map( A1 => n20351, A2 => n20341, B1 => n20670, B2 => 
                           n18745, ZN => n21247);
   U10474 : XNOR2_X1 port map( A => n4294, B => n22697, ZN => n20047);
   U10475 : XNOR2_X1 port map( A => n4294, B => n2036, ZN => n20983);
   U10476 : XNOR2_X1 port map( A => n4294, B => n21699, ZN => n21221);
   U10477 : XNOR2_X1 port map( A => n21054, B => n4294, ZN => n21564);
   U10479 : NAND2_X1 port map( A1 => n4295, A2 => n20302, ZN => n4692);
   U10480 : INV_X1 port map( A => n20009, ZN => n4295);
   U10481 : NAND2_X1 port map( A1 => n4298, A2 => n24570, ZN => n4297);
   U10482 : INV_X1 port map( A => n16774, ZN => n4299);
   U10484 : AND2_X1 port map( A1 => n4303, A2 => n17114, ZN => n5429);
   U10485 : NOR2_X1 port map( A1 => n17100, A2 => n17114, ZN => n5760);
   U10486 : INV_X1 port map( A => n17118, ZN => n4303);
   U10487 : OAI21_X1 port map( B1 => n16573, B2 => n25357, A => n4304, ZN => 
                           n4714);
   U10489 : MUX2_X1 port map( A => n13965, B => n11806, S => n13966, Z => 
                           n13885);
   U10490 : NAND2_X1 port map( A1 => n13965, A2 => n11806, ZN => n4305);
   U10491 : MUX2_X1 port map( A => n13725, B => n13883, S => n11806, Z => 
                           n13726);
   U10492 : NOR2_X1 port map( A1 => n20478, A2 => n20003, ZN => n19627);
   U10493 : NOR2_X2 port map( A1 => n18838, A2 => n4306, ZN => n20478);
   U10494 : AOI21_X1 port map( B1 => n19239, B2 => n19064, A => n4307, ZN => 
                           n4306);
   U10496 : NAND2_X1 port map( A1 => n19213, A2 => n4315, ZN => n4314);
   U10497 : XNOR2_X1 port map( A => n11615, B => n11614, ZN => n4316);
   U10498 : OAI21_X1 port map( B1 => n19363, B2 => n24424, A => n24968, ZN => 
                           n4317);
   U10499 : NAND3_X1 port map( A1 => n13065, A2 => n4319, A3 => n4318, ZN => 
                           n13385);
   U10500 : NAND3_X1 port map( A1 => n13064, A2 => n13063, A3 => n12737, ZN => 
                           n4318);
   U10501 : INV_X1 port map( A => n13159, ZN => n12737);
   U10502 : OAI21_X1 port map( B1 => n13062, B2 => n4320, A => n13163, ZN => 
                           n4319);
   U10503 : INV_X1 port map( A => n6956, ZN => n6702);
   U10504 : OAI21_X1 port map( B1 => n3926, B2 => n6703, A => n4323, ZN => 
                           n4322);
   U10505 : INV_X1 port map( A => n11009, ZN => n4326);
   U10506 : NOR2_X1 port map( A1 => n1218, A2 => n11009, ZN => n11055);
   U10507 : INV_X1 port map( A => n13796, ZN => n13774);
   U10508 : XNOR2_X1 port map( A => n4334, B => n8914, ZN => n8131);
   U10509 : XNOR2_X1 port map( A => n8914, B => n4335, ZN => n8197);
   U10510 : NAND2_X1 port map( A1 => n4336, A2 => n13072, ZN => n12775);
   U10511 : NAND3_X1 port map( A1 => n23179, A2 => n23167, A3 => n25488, ZN => 
                           n22555);
   U10512 : NAND3_X1 port map( A1 => n4344, A2 => n4347, A3 => n7130, ZN => 
                           n8826);
   U10513 : NAND2_X1 port map( A1 => n4345, A2 => n7320, ZN => n4344);
   U10514 : NAND2_X1 port map( A1 => n20650, A2 => n24415, ZN => n4348);
   U10516 : NAND2_X1 port map( A1 => n20648, A2 => n22141, ZN => n4351);
   U10518 : OR2_X1 port map( A1 => n15802, A2 => n1365, ZN => n15594);
   U10519 : INV_X1 port map( A => n24826, ZN => n4353);
   U10520 : NAND2_X1 port map( A1 => n4355, A2 => n14160, ZN => n4354);
   U10521 : XNOR2_X1 port map( A => n12048, B => n1792, ZN => n11916);
   U10522 : NAND2_X1 port map( A1 => n10899, A2 => n4341, ZN => n4358);
   U10523 : NAND2_X1 port map( A1 => n23722, A2 => n23727, ZN => n23726);
   U10525 : NAND2_X1 port map( A1 => n22081, A2 => n4360, ZN => n4359);
   U10526 : INV_X1 port map( A => n22079, ZN => n4360);
   U10527 : NAND2_X1 port map( A1 => n22080, A2 => n22079, ZN => n4361);
   U10528 : NAND2_X1 port map( A1 => n4364, A2 => n3726, ZN => n4363);
   U10529 : MUX2_X1 port map( A => n19163, B => n19393, S => n19162, Z => n4364
                           );
   U10531 : NAND2_X1 port map( A1 => n8316, A2 => n8315, ZN => n4366);
   U10534 : NAND3_X1 port map( A1 => n24532, A2 => n24586, A3 => n16107, ZN => 
                           n15628);
   U10535 : NAND2_X1 port map( A1 => n6942, A2 => n6941, ZN => n4369);
   U10536 : NAND2_X1 port map( A1 => n5560, A2 => n6947, ZN => n4370);
   U10537 : NOR3_X1 port map( A1 => n22974, A2 => n22975, A3 => n22387, ZN => 
                           n4371);
   U10538 : NOR2_X1 port map( A1 => n4373, A2 => n21822, ZN => n19343);
   U10539 : NOR2_X1 port map( A1 => n332, A2 => n21822, ZN => n4374);
   U10540 : XNOR2_X1 port map( A => n8039, B => n8452, ZN => n9114);
   U10541 : XNOR2_X1 port map( A => n9114, B => n9115, ZN => n9119);
   U10542 : OAI21_X1 port map( B1 => n7535, B2 => n7536, A => n8013, ZN => 
                           n4377);
   U10543 : XNOR2_X1 port map( A => n4378, B => n2034, ZN => n7204);
   U10544 : XNOR2_X1 port map( A => n4378, B => n2193, ZN => n8264);
   U10545 : XNOR2_X1 port map( A => n8485, B => n4378, ZN => n8246);
   U10546 : XNOR2_X1 port map( A => n8698, B => n4378, ZN => n7778);
   U10547 : NAND2_X1 port map( A1 => n12107, A2 => n400, ZN => n4379);
   U10548 : NAND2_X1 port map( A1 => n4381, A2 => n13335, ZN => n4380);
   U10549 : INV_X1 port map( A => n13337, ZN => n4381);
   U10550 : NAND2_X1 port map( A1 => n14005, A2 => n24462, ZN => n4383);
   U10551 : XNOR2_X1 port map( A => n17648, B => n4384, ZN => n4385);
   U10552 : INV_X1 port map( A => n17918, ZN => n4384);
   U10553 : XNOR2_X1 port map( A => n8697, B => n8696, ZN => n4386);
   U10554 : INV_X1 port map( A => n12834, ZN => n13273);
   U10555 : NAND3_X1 port map( A1 => n4394, A2 => n4393, A3 => n4390, ZN => 
                           n11736);
   U10556 : NAND3_X1 port map( A1 => n4326, A2 => n11057, A3 => n10694, ZN => 
                           n4393);
   U10557 : NOR2_X2 port map( A1 => n9794, A2 => n9793, ZN => n11052);
   U10558 : NAND2_X1 port map( A1 => n11055, A2 => n11054, ZN => n4394);
   U10559 : XNOR2_X1 port map( A => n21092, B => n24453, ZN => n21095);
   U10560 : XNOR2_X1 port map( A => n21542, B => n24453, ZN => n21546);
   U10561 : XNOR2_X1 port map( A => n21611, B => n4396, ZN => n20035);
   U10564 : NOR2_X1 port map( A1 => n4525, A2 => n13901, ZN => n14309);
   U10565 : OAI21_X1 port map( B1 => n7972, B2 => n7977, A => n4400, ZN => 
                           n7817);
   U10566 : MUX2_X1 port map( A => n7972, B => n7973, S => n4400, Z => n7979);
   U10567 : AOI21_X1 port map( B1 => n7049, B2 => n7819, A => n4400, ZN => 
                           n7050);
   U10568 : XNOR2_X1 port map( A => n8881, B => n4401, ZN => n8883);
   U10569 : OAI21_X1 port map( B1 => n20069, B2 => n20068, A => n20067, ZN => 
                           n20070);
   U10570 : NAND2_X1 port map( A1 => n20068, A2 => n19849, ZN => n20067);
   U10571 : NAND2_X1 port map( A1 => n18849, A2 => n18848, ZN => n4404);
   U10575 : NAND2_X1 port map( A1 => n23397, A2 => n23396, ZN => n4406);
   U10579 : NOR2_X1 port map( A1 => n23396, A2 => n23394, ZN => n4411);
   U10580 : AND2_X1 port map( A1 => n17172, A2 => n17175, ZN => n4414);
   U10583 : XNOR2_X1 port map( A => n15191, B => n15112, ZN => n14937);
   U10584 : XNOR2_X1 port map( A => n15246, B => n14937, ZN => n14583);
   U10585 : NAND2_X1 port map( A1 => n4419, A2 => n4417, ZN => n4416);
   U10586 : NAND2_X1 port map( A1 => n16148, A2 => n4418, ZN => n4417);
   U10587 : AOI21_X1 port map( B1 => n16097, B2 => n16096, A => n213, ZN => 
                           n4419);
   U10588 : AND2_X1 port map( A1 => n4422, A2 => n412, ZN => n10439);
   U10589 : NAND2_X1 port map( A1 => n10438, A2 => n4422, ZN => n10442);
   U10591 : NAND2_X1 port map( A1 => n14154, A2 => n14153, ZN => n4424);
   U10592 : NAND2_X1 port map( A1 => n4426, A2 => n17320, ZN => n17324);
   U10593 : INV_X1 port map( A => n16607, ZN => n4426);
   U10594 : NAND2_X2 port map( A1 => n4428, A2 => n6378, ZN => n7843);
   U10595 : NAND2_X1 port map( A1 => n6790, A2 => n6089, ZN => n4428);
   U10597 : OR2_X1 port map( A1 => n19283, A2 => n19127, ZN => n4429);
   U10598 : NAND3_X1 port map( A1 => n4432, A2 => n19518, A3 => n4431, ZN => 
                           n4430);
   U10599 : NAND2_X1 port map( A1 => n4433, A2 => n19526, ZN => n4432);
   U10601 : OAI211_X1 port map( C1 => n21814, C2 => n22063, A => n21813, B => 
                           n21812, ZN => n4434);
   U10603 : XNOR2_X2 port map( A => n16785, B => n16786, ZN => n4436);
   U10604 : AND2_X1 port map( A1 => n19266, A2 => n4436, ZN => n5239);
   U10605 : NAND2_X1 port map( A1 => n1299, A2 => n4436, ZN => n16822);
   U10607 : NAND2_X1 port map( A1 => n18916, A2 => n4436, ZN => n19149);
   U10608 : NAND3_X1 port map( A1 => n1336, A2 => n22244, A3 => n4437, ZN => 
                           n22246);
   U10609 : INV_X1 port map( A => n22059, ZN => n4437);
   U10610 : AOI21_X1 port map( B1 => n19601, B2 => n18037, A => n4438, ZN => 
                           n19603);
   U10611 : NAND2_X1 port map( A1 => n19255, A2 => n19598, ZN => n4439);
   U10613 : NAND3_X1 port map( A1 => n16075, A2 => n1365, A3 => n16077, ZN => 
                           n4440);
   U10614 : NOR2_X1 port map( A1 => n22334, A2 => n22333, ZN => n4441);
   U10616 : NAND2_X1 port map( A1 => n4449, A2 => n13266, ZN => n4443);
   U10617 : NAND2_X1 port map( A1 => n14301, A2 => n13888, ZN => n13944);
   U10620 : INV_X1 port map( A => n12835, ZN => n4445);
   U10621 : NAND2_X1 port map( A1 => n4930, A2 => n12680, ZN => n4449);
   U10622 : NAND2_X1 port map( A1 => n4450, A2 => n24391, ZN => n5295);
   U10624 : NAND2_X1 port map( A1 => n12819, A2 => n4451, ZN => n4721);
   U10625 : NAND2_X1 port map( A1 => n14168, A2 => n13742, ZN => n4452);
   U10627 : OAI211_X2 port map( C1 => n10185, C2 => n10186, A => n10184, B => 
                           n10183, ZN => n10660);
   U10628 : INV_X1 port map( A => n20434, ZN => n19225);
   U10629 : MUX2_X2 port map( A => n9583, B => n9582, S => n25463, Z => n10617)
                           ;
   U10630 : INV_X1 port map( A => n4882, ZN => n18028);
   U10633 : MUX2_X2 port map( A => n10067, B => n10066, S => n10065, Z => 
                           n11070);
   U10635 : OAI21_X1 port map( B1 => n239, B2 => n9864, A => n4453, ZN => n8064
                           );
   U10636 : NAND2_X1 port map( A1 => n9864, A2 => n9857, ZN => n4453);
   U10637 : INV_X1 port map( A => n9859, ZN => n4454);
   U10638 : MUX2_X1 port map( A => n9860, B => n9559, S => n239, Z => n9262);
   U10640 : XNOR2_X1 port map( A => n4456, B => n21167, ZN => n4455);
   U10641 : NAND2_X1 port map( A1 => n19276, A2 => n1334, ZN => n4458);
   U10643 : NAND2_X1 port map( A1 => n19125, A2 => n5573, ZN => n4459);
   U10644 : INV_X1 port map( A => n10713, ZN => n4463);
   U10645 : OAI21_X1 port map( B1 => n5744, B2 => n11131, A => n11129, ZN => 
                           n4465);
   U10646 : NOR2_X1 port map( A1 => n4463, A2 => n10838, ZN => n4462);
   U10647 : OAI21_X1 port map( B1 => n22656, B2 => n331, A => n4466, ZN => 
                           n4473);
   U10648 : NAND2_X1 port map( A1 => n22813, A2 => n22656, ZN => n4466);
   U10649 : OAI21_X1 port map( B1 => n22656, B2 => n22657, A => n25241, ZN => 
                           n4467);
   U10650 : INV_X1 port map( A => n22658, ZN => n4470);
   U10651 : XNOR2_X2 port map( A => n20408, B => n20407, ZN => n22813);
   U10652 : NAND2_X1 port map( A1 => n24015, A2 => n4478, ZN => n4474);
   U10653 : NAND2_X1 port map( A1 => n4478, A2 => n23993, ZN => n23987);
   U10654 : NAND2_X1 port map( A1 => n23982, A2 => n4478, ZN => n23981);
   U10655 : AOI21_X1 port map( B1 => n24954, B2 => n4477, A => n23983, ZN => 
                           n4476);
   U10656 : NAND4_X2 port map( A1 => n12436, A2 => n12437, A3 => n12438, A4 => 
                           n12435, ZN => n14167);
   U10657 : NOR2_X2 port map( A1 => n19593, A2 => n4479, ZN => n20377);
   U10658 : MUX2_X1 port map( A => n24483, B => n19591, S => n19077, Z => n4480
                           );
   U10659 : NOR2_X1 port map( A1 => n10365, A2 => n4481, ZN => n10321);
   U10660 : OAI21_X1 port map( B1 => n10684, B2 => n11004, A => n4481, ZN => 
                           n11008);
   U10661 : NAND2_X1 port map( A1 => n17012, A2 => n25491, ZN => n4482);
   U10662 : OAI21_X1 port map( B1 => n7956, B2 => n4483, A => n7955, ZN => 
                           n7957);
   U10663 : NAND2_X1 port map( A1 => n4486, A2 => n4484, ZN => n12887);
   U10665 : NAND3_X1 port map( A1 => n17613, A2 => n17409, A3 => n17608, ZN => 
                           n4488);
   U10666 : NAND3_X1 port map( A1 => n19948, A2 => n4489, A3 => n20461, ZN => 
                           n19949);
   U10667 : MUX2_X1 port map( A => n20383, B => n20384, S => n20459, Z => 
                           n20398);
   U10669 : NAND2_X1 port map( A1 => n12937, A2 => n4490, ZN => n4492);
   U10671 : NAND2_X1 port map( A1 => n11006, A2 => n24420, ZN => n4495);
   U10672 : NAND2_X1 port map( A1 => n11836, A2 => n12902, ZN => n4497);
   U10674 : NAND2_X1 port map( A1 => n17416, A2 => n16565, ZN => n4502);
   U10675 : AOI21_X1 port map( B1 => n4503, B2 => n6678, A => n6281, ZN => 
                           n6282);
   U10676 : XNOR2_X1 port map( A => n14843, B => n14842, ZN => n4504);
   U10677 : INV_X1 port map( A => n10753, ZN => n4505);
   U10678 : NAND2_X1 port map( A1 => n9364, A2 => n4506, ZN => n10204);
   U10679 : INV_X1 port map( A => n17297, ZN => n4508);
   U10680 : INV_X1 port map( A => n4510, ZN => n14021);
   U10681 : NAND2_X1 port map( A1 => n4510, A2 => n14022, ZN => n12513);
   U10682 : NAND2_X1 port map( A1 => n14086, A2 => n4510, ZN => n14087);
   U10683 : NAND2_X1 port map( A1 => n2008, A2 => n6933, ZN => n4512);
   U10684 : NAND2_X1 port map( A1 => n11113, A2 => n11116, ZN => n5351);
   U10685 : NAND2_X1 port map( A1 => n9789, A2 => n24575, ZN => n5354);
   U10686 : NAND2_X1 port map( A1 => n22151, A2 => n4513, ZN => n22152);
   U10687 : OR2_X1 port map( A1 => n23647, A2 => n23612, ZN => n4514);
   U10688 : OR2_X1 port map( A1 => n24366, A2 => n4516, ZN => n4515);
   U10689 : INV_X1 port map( A => n16001, ZN => n4516);
   U10690 : OAI21_X1 port map( B1 => n13055, B2 => n13054, A => n4517, ZN => 
                           n12484);
   U10691 : OR2_X1 port map( A1 => n13053, A2 => n13055, ZN => n12753);
   U10693 : NAND2_X1 port map( A1 => n4523, A2 => n4522, ZN => n9811);
   U10694 : NAND2_X1 port map( A1 => n9789, A2 => n9788, ZN => n4523);
   U10695 : NAND2_X1 port map( A1 => n13901, A2 => n4525, ZN => n4524);
   U10698 : NOR2_X1 port map( A1 => n10244, A2 => n10799, ZN => n10804);
   U10699 : NAND3_X1 port map( A1 => n10651, A2 => n10800, A3 => n4527, ZN => 
                           n10248);
   U10700 : NAND3_X1 port map( A1 => n10244, A2 => n10651, A3 => n4527, ZN => 
                           n9966);
   U10701 : AOI21_X1 port map( B1 => n411, B2 => n4527, A => n10805, ZN => 
                           n10428);
   U10702 : NAND2_X1 port map( A1 => n5427, A2 => n20269, ZN => n20230);
   U10703 : NOR2_X1 port map( A1 => n16845, A2 => n16846, ZN => n4528);
   U10704 : INV_X1 port map( A => n13353, ZN => n5626);
   U10705 : AND2_X1 port map( A1 => n5626, A2 => n5624, ZN => n5625);
   U10706 : NOR2_X1 port map( A1 => n4531, A2 => n11044, ZN => n4530);
   U10707 : INV_X1 port map( A => n11051, ZN => n4531);
   U10708 : OAI21_X1 port map( B1 => n11046, B2 => n2680, A => n4532, ZN => 
                           n11047);
   U10709 : MUX2_X1 port map( A => n11046, B => n11045, S => n11044, Z => 
                           n10418);
   U10711 : NAND2_X1 port map( A1 => n7867, A2 => n7862, ZN => n4534);
   U10713 : NAND2_X1 port map( A1 => n22832, A2 => n22936, ZN => n4609);
   U10714 : XNOR2_X1 port map( A => n12200, B => n12201, ZN => n12202);
   U10716 : INV_X1 port map( A => n19386, ZN => n4543);
   U10717 : NAND2_X2 port map( A1 => n4544, A2 => n6569, ZN => n7923);
   U10718 : OAI21_X1 port map( B1 => n13219, B2 => n13220, A => n4546, ZN => 
                           n4548);
   U10719 : NOR2_X1 port map( A1 => n4052, A2 => n18808, ZN => n4551);
   U10720 : INV_X1 port map( A => n18808, ZN => n5134);
   U10722 : INV_X1 port map( A => n16795, ZN => n4554);
   U10724 : NOR2_X1 port map( A1 => n4553, A2 => n16551, ZN => n4552);
   U10725 : XNOR2_X1 port map( A => n4556, B => n14430, ZN => n15308);
   U10726 : INV_X1 port map( A => n15303, ZN => n4556);
   U10727 : XNOR2_X1 port map( A => n4557, B => n14430, ZN => n13499);
   U10728 : XNOR2_X1 port map( A => n3990, B => n18579, ZN => n18581);
   U10729 : NAND2_X1 port map( A1 => n17596, A2 => n17597, ZN => n4563);
   U10730 : AND2_X1 port map( A1 => n17600, A2 => n2968, ZN => n4566);
   U10731 : NOR2_X1 port map( A1 => n4567, A2 => n13335, ZN => n4822);
   U10732 : XNOR2_X2 port map( A => n4820, B => n4568, ZN => n13335);
   U10733 : INV_X1 port map( A => n13341, ZN => n4567);
   U10734 : NAND3_X2 port map( A1 => n4570, A2 => n18913, A3 => n4569, ZN => 
                           n21678);
   U10736 : INV_X1 port map( A => n20125, ZN => n20545);
   U10738 : NAND2_X1 port map( A1 => n17226, A2 => n17227, ZN => n4573);
   U10739 : AOI21_X2 port map( B1 => n4576, B2 => n10459, A => n10458, ZN => 
                           n11653);
   U10740 : MUX2_X1 port map( A => n10730, B => n10734, S => n11190, Z => n4576
                           );
   U10741 : NAND2_X1 port map( A1 => n19420, A2 => n19418, ZN => n19168);
   U10742 : XNOR2_X1 port map( A => n14654, B => n14799, ZN => n4582);
   U10743 : XNOR2_X1 port map( A => n14599, B => n14909, ZN => n4583);
   U10744 : AOI21_X1 port map( B1 => n24499, B2 => n403, A => n1324, ZN => 
                           n13175);
   U10745 : NAND3_X1 port map( A1 => n12727, A2 => n12726, A3 => n4584, ZN => 
                           n13975);
   U10746 : NAND2_X1 port map( A1 => n13178, A2 => n12506, ZN => n4584);
   U10747 : MUX2_X1 port map( A => n12652, B => n12651, S => n12506, Z => 
                           n13668);
   U10748 : NAND2_X1 port map( A1 => n19501, A2 => n19500, ZN => n4585);
   U10749 : NAND2_X1 port map( A1 => n4586, A2 => n10148, ZN => n5355);
   U10750 : AOI21_X1 port map( B1 => n3317, B2 => n17390, A => n3604, ZN => 
                           n16875);
   U10751 : NAND2_X1 port map( A1 => n25465, A2 => n17185, ZN => n17390);
   U10752 : NAND2_X1 port map( A1 => n15880, A2 => n24385, ZN => n15635);
   U10753 : OR2_X1 port map( A1 => n7155, A2 => n4588, ZN => n7912);
   U10754 : NAND2_X1 port map( A1 => n5636, A2 => n5635, ZN => n4588);
   U10756 : XNOR2_X1 port map( A => n10771, B => n11913, ZN => n10564);
   U10757 : XNOR2_X1 port map( A => n10771, B => n4589, ZN => n9217);
   U10758 : XNOR2_X1 port map( A => n4590, B => n11582, ZN => n11512);
   U10759 : NAND2_X1 port map( A1 => n3653, A2 => n19300, ZN => n18932);
   U10760 : INV_X1 port map( A => n22406, ZN => n4591);
   U10761 : XNOR2_X1 port map( A => n15054, B => n14500, ZN => n15267);
   U10762 : NAND2_X1 port map( A1 => n13364, A2 => n13363, ZN => n4595);
   U10763 : NAND2_X1 port map( A1 => n12977, A2 => n13365, ZN => n4596);
   U10764 : INV_X1 port map( A => n24503, ZN => n4597);
   U10765 : NAND2_X1 port map( A1 => n4602, A2 => n19014, ZN => n4601);
   U10767 : NAND2_X1 port map( A1 => n25489, A2 => n24407, ZN => n4602);
   U10770 : NAND2_X1 port map( A1 => n23370, A2 => n24404, ZN => n22991);
   U10771 : NAND3_X1 port map( A1 => n23370, A2 => n24404, A3 => n4606, ZN => 
                           n4607);
   U10772 : INV_X1 port map( A => n23379, ZN => n4606);
   U10773 : NAND2_X1 port map( A1 => n4609, A2 => n4608, ZN => n21657);
   U10774 : XNOR2_X1 port map( A => n11435, B => n11665, ZN => n4610);
   U10775 : INV_X1 port map( A => n11665, ZN => n11764);
   U10776 : XNOR2_X1 port map( A => n9217, B => n11061, ZN => n4611);
   U10777 : XNOR2_X1 port map( A => n18540, B => n18080, ZN => n18183);
   U10779 : NAND2_X1 port map( A1 => n16893, A2 => n17481, ZN => n4613);
   U10780 : NAND2_X1 port map( A1 => n16739, A2 => n16578, ZN => n16740);
   U10781 : INV_X1 port map( A => n15873, ZN => n16739);
   U10782 : INV_X1 port map( A => n20140, ZN => n4616);
   U10783 : NOR2_X1 port map( A1 => n5269, A2 => n16217, ZN => n4617);
   U10784 : AND2_X1 port map( A1 => n16219, A2 => n15921, ZN => n16217);
   U10785 : NOR2_X1 port map( A1 => n10149, A2 => n25486, ZN => n5357);
   U10786 : NAND3_X1 port map( A1 => n6314, A2 => n4620, A3 => n6470, ZN => 
                           n4619);
   U10788 : NAND2_X1 port map( A1 => n9857, A2 => n239, ZN => n4622);
   U10790 : NAND2_X1 port map( A1 => n4625, A2 => n44, ZN => n10796);
   U10791 : AOI22_X1 port map( A1 => n24526, A2 => n11199, B1 => n4625, B2 => 
                           n11201, ZN => n11202);
   U10792 : NAND2_X1 port map( A1 => n23160, A2 => n24325, ZN => n4626);
   U10795 : INV_X1 port map( A => n22424, ZN => n4632);
   U10796 : XNOR2_X1 port map( A => n15269, B => n4636, ZN => n4635);
   U10797 : XNOR2_X1 port map( A => n14721, B => n15055, ZN => n15269);
   U10798 : XNOR2_X1 port map( A => n15268, B => n15267, ZN => n4637);
   U10799 : INV_X1 port map( A => n12797, ZN => n4640);
   U10800 : NAND2_X1 port map( A1 => n13792, A2 => n13795, ZN => n14181);
   U10801 : NAND2_X1 port map( A1 => n4644, A2 => n7022, ZN => n4642);
   U10802 : INV_X1 port map( A => n7266, ZN => n7193);
   U10803 : NOR2_X1 port map( A1 => n442, A2 => n4643, ZN => n4644);
   U10804 : NAND2_X1 port map( A1 => n4645, A2 => n4646, ZN => n17368);
   U10805 : NAND2_X1 port map( A1 => n19201, A2 => n4647, ZN => n19843);
   U10810 : XNOR2_X2 port map( A => n21682, B => n21683, ZN => n22901);
   U10811 : NAND2_X1 port map( A1 => n4651, A2 => n24513, ZN => n12987);
   U10813 : NAND2_X1 port map( A1 => n13220, A2 => n24513, ZN => n4652);
   U10814 : NAND2_X1 port map( A1 => n17896, A2 => n19479, ZN => n4653);
   U10815 : NAND2_X1 port map( A1 => n20117, A2 => n20109, ZN => n20113);
   U10816 : OAI22_X1 port map( A1 => n11081, A2 => n10766, B1 => n3119, B2 => 
                           n4654, ZN => n10770);
   U10817 : NAND2_X1 port map( A1 => n4656, A2 => n309, ZN => n4655);
   U10818 : XNOR2_X1 port map( A => n4657, B => n21023, ZN => n21026);
   U10819 : OAI21_X1 port map( B1 => n17124, B2 => n17123, A => n4664, ZN => 
                           n4658);
   U10820 : OAI21_X1 port map( B1 => n17124, B2 => n4663, A => n4658, ZN => 
                           n17587);
   U10821 : NAND2_X1 port map( A1 => n4661, A2 => n4659, ZN => n18430);
   U10822 : NAND3_X1 port map( A1 => n17117, A2 => n17824, A3 => n4660, ZN => 
                           n4659);
   U10823 : INV_X1 port map( A => n17123, ZN => n4660);
   U10824 : XNOR2_X1 port map( A => n4665, B => n18049, ZN => n4667);
   U10825 : XNOR2_X1 port map( A => n4666, B => n17588, ZN => n4665);
   U10827 : XNOR2_X1 port map( A => n4670, B => n4669, ZN => n12192);
   U10828 : INV_X1 port map( A => n2746, ZN => n4669);
   U10829 : NAND2_X1 port map( A1 => n7942, A2 => n4672, ZN => n7944);
   U10830 : NAND2_X1 port map( A1 => n6889, A2 => n6888, ZN => n4673);
   U10831 : NAND2_X1 port map( A1 => n6887, A2 => n6886, ZN => n4674);
   U10832 : NAND2_X1 port map( A1 => n16106, A2 => n16109, ZN => n4678);
   U10833 : XNOR2_X1 port map( A => n18560, B => n18464, ZN => n4679);
   U10834 : INV_X1 port map( A => n18560, ZN => n18130);
   U10835 : NAND2_X1 port map( A1 => n4680, A2 => n12993, ZN => n12890);
   U10836 : NAND2_X1 port map( A1 => n6526, A2 => n6952, ZN => n4682);
   U10837 : OAI211_X1 port map( C1 => n4684, C2 => n17130, A => n17134, B => 
                           n25226, ZN => n4683);
   U10839 : INV_X1 port map( A => n17134, ZN => n4686);
   U10841 : NAND2_X1 port map( A1 => n24407, A2 => n18788, ZN => n18443);
   U10843 : NAND2_X1 port map( A1 => n5149, A2 => n19395, ZN => n5501);
   U10844 : INV_X1 port map( A => n10992, ZN => n4691);
   U10846 : NAND2_X1 port map( A1 => n6053, A2 => n5775, ZN => n4694);
   U10847 : INV_X1 port map( A => n5774, ZN => n6409);
   U10848 : INV_X1 port map( A => n6744, ZN => n4696);
   U10849 : NAND2_X1 port map( A1 => n5777, A2 => n6628, ZN => n4697);
   U10850 : NAND4_X1 port map( A1 => n4699, A2 => n4698, A3 => n4704, A4 => 
                           n2744, ZN => n4702);
   U10851 : INV_X1 port map( A => n22999, ZN => n4698);
   U10852 : INV_X1 port map( A => n23000, ZN => n4699);
   U10853 : OAI21_X1 port map( B1 => n4701, B2 => n22999, A => n444, ZN => 
                           n4700);
   U10854 : INV_X1 port map( A => n4704, ZN => n4701);
   U10855 : NAND2_X1 port map( A1 => n23000, A2 => n444, ZN => n4703);
   U10856 : NAND3_X1 port map( A1 => n22749, A2 => n22998, A3 => n1442, ZN => 
                           n4704);
   U10857 : OAI21_X1 port map( B1 => n10095, B2 => n10098, A => n8359, ZN => 
                           n8384);
   U10858 : INV_X1 port map( A => n8351, ZN => n4705);
   U10860 : OAI211_X1 port map( C1 => n8352, C2 => n4711, A => n4710, B => 
                           n4709, ZN => n8354);
   U10861 : NAND2_X1 port map( A1 => n16418, A2 => n16408, ZN => n15866);
   U10862 : XNOR2_X1 port map( A => n14729, B => n14444, ZN => n4712);
   U10864 : NAND2_X1 port map( A1 => n5774, A2 => n6050, ZN => n6052);
   U10865 : NAND2_X1 port map( A1 => n5774, A2 => n6744, ZN => n6629);
   U10866 : NAND2_X1 port map( A1 => n5774, A2 => n6630, ZN => n5775);
   U10867 : NAND2_X1 port map( A1 => n6628, A2 => n5774, ZN => n6748);
   U10868 : NAND3_X1 port map( A1 => n6051, A2 => n5774, A3 => n4696, ZN => 
                           n6410);
   U10869 : AOI21_X1 port map( B1 => n6566, B2 => n6746, A => n5774, ZN => 
                           n7927);
   U10870 : NAND2_X1 port map( A1 => n20301, A2 => n20009, ZN => n19049);
   U10871 : MUX2_X1 port map( A => n14458, B => n3404, S => n3401, Z => n14318)
                           ;
   U10872 : NAND2_X1 port map( A1 => n24079, A2 => n4715, ZN => n4716);
   U10873 : NAND2_X1 port map( A1 => n5439, A2 => n24079, ZN => n4717);
   U10874 : XNOR2_X1 port map( A => n18041, B => n18040, ZN => n19071);
   U10875 : NAND2_X1 port map( A1 => n4720, A2 => n4718, ZN => n23425);
   U10876 : OAI22_X1 port map( A1 => n22528, A2 => n23425, B1 => n1370, B2 => 
                           n23442, ZN => n23453);
   U10877 : XNOR2_X1 port map( A => n4723, B => n14579, ZN => n14840);
   U10878 : NOR2_X2 port map( A1 => n4722, A2 => n4721, ZN => n14579);
   U10879 : AOI21_X1 port map( B1 => n12818, B2 => n14172, A => n13526, ZN => 
                           n4722);
   U10880 : NAND3_X1 port map( A1 => n16461, A2 => n16462, A3 => n16460, ZN => 
                           n4725);
   U10881 : OAI211_X2 port map( C1 => n9453, C2 => n9935, A => n9451, B => 
                           n9452, ZN => n10885);
   U10883 : NAND2_X1 port map( A1 => n6429, A2 => n6785, ZN => n4727);
   U10884 : NAND3_X1 port map( A1 => n25242, A2 => n20136, A3 => n4728, ZN => 
                           n19756);
   U10885 : NAND2_X1 port map( A1 => n5566, A2 => n4728, ZN => n5565);
   U10886 : AOI21_X1 port map( B1 => n20135, B2 => n4728, A => n19755, ZN => 
                           n19758);
   U10887 : NAND2_X1 port map( A1 => n5436, A2 => n4729, ZN => n12862);
   U10888 : OAI21_X1 port map( B1 => n10759, B2 => n10757, A => n10756, ZN => 
                           n4733);
   U10889 : XNOR2_X2 port map( A => n5981, B => Key(125), ZN => n7007);
   U10890 : NAND3_X1 port map( A1 => n15130, A2 => n4735, A3 => n4734, ZN => 
                           n17381);
   U10891 : NAND2_X1 port map( A1 => n15118, A2 => n24919, ZN => n4734);
   U10892 : OAI21_X1 port map( B1 => n1434, B2 => n15117, A => n24841, ZN => 
                           n4735);
   U10893 : NOR2_X1 port map( A1 => n10985, A2 => n10552, ZN => n4736);
   U10894 : NAND2_X1 port map( A1 => n10554, A2 => n4737, ZN => n4739);
   U10896 : NOR2_X1 port map( A1 => n11160, A2 => n11163, ZN => n10553);
   U10897 : NOR2_X2 port map( A1 => n4740, A2 => n4738, ZN => n11761);
   U10898 : MUX2_X1 port map( A => n24490, B => n13222, S => n24965, Z => n4741
                           );
   U10899 : NAND2_X1 port map( A1 => n17426, A2 => n17379, ZN => n4742);
   U10900 : NAND2_X1 port map( A1 => n4745, A2 => n25014, ZN => n4744);
   U10901 : NAND2_X1 port map( A1 => n4746, A2 => n4747, ZN => n4745);
   U10902 : NAND2_X1 port map( A1 => n6530, A2 => n24067, ZN => n4747);
   U10903 : XNOR2_X2 port map( A => Key(27), B => Plaintext(27), ZN => n6530);
   U10904 : NOR2_X1 port map( A1 => n19500, A2 => n4748, ZN => n18720);
   U10905 : NOR2_X1 port map( A1 => n19502, A2 => n3296, ZN => n18983);
   U10906 : NAND2_X1 port map( A1 => n19497, A2 => n3296, ZN => n19495);
   U10907 : OAI21_X1 port map( B1 => n19335, B2 => n19500, A => n3296, ZN => 
                           n17924);
   U10908 : AOI21_X1 port map( B1 => n18987, B2 => n17938, A => n4748, ZN => 
                           n17939);
   U10910 : NAND3_X1 port map( A1 => n20236, A2 => n20170, A3 => n20239, ZN => 
                           n4750);
   U10912 : NAND2_X1 port map( A1 => n5802, A2 => n5801, ZN => n4753);
   U10913 : NAND2_X1 port map( A1 => n14157, A2 => n14156, ZN => n14163);
   U10915 : XNOR2_X1 port map( A => n4759, B => n11838, ZN => n12239);
   U10916 : OAI211_X2 port map( C1 => n10550, C2 => n3509, A => n10551, B => 
                           n4758, ZN => n11838);
   U10918 : NOR2_X1 port map( A1 => n5376, A2 => n16796, ZN => n4760);
   U10919 : OAI21_X1 port map( B1 => n19597, B2 => n19598, A => n19255, ZN => 
                           n19075);
   U10920 : MUX2_X1 port map( A => n19255, B => n19596, S => n19597, Z => 
                           n18054);
   U10921 : NAND2_X1 port map( A1 => n4764, A2 => n24919, ZN => n15897);
   U10922 : NAND2_X1 port map( A1 => n15748, A2 => n16293, ZN => n4764);
   U10923 : NAND2_X1 port map( A1 => n16357, A2 => n16356, ZN => n15748);
   U10924 : NOR2_X1 port map( A1 => n4766, A2 => n13170, ZN => n12720);
   U10925 : NOR2_X1 port map( A1 => n4766, A2 => n13165, ZN => n13166);
   U10926 : XNOR2_X2 port map( A => n18180, B => n18179, ZN => n19522);
   U10927 : OR2_X1 port map( A1 => n14278, A2 => n24572, ZN => n4771);
   U10928 : NAND3_X1 port map( A1 => n4225, A2 => n14850, A3 => n4767, ZN => 
                           n4769);
   U10929 : XNOR2_X1 port map( A => n14980, B => n14789, ZN => n15338);
   U10932 : NAND2_X1 port map( A1 => n14416, A2 => n13617, ZN => n4770);
   U10933 : NAND2_X1 port map( A1 => n16484, A2 => n16481, ZN => n4772);
   U10934 : INV_X1 port map( A => n25218, ZN => n4775);
   U10937 : NAND2_X1 port map( A1 => n24927, A2 => n262, ZN => n7572);
   U10938 : INV_X1 port map( A => n10518, ZN => n4779);
   U10939 : OAI211_X1 port map( C1 => n10520, C2 => n10829, A => n4778, B => 
                           n4777, ZN => n10279);
   U10940 : NAND2_X1 port map( A1 => n10830, A2 => n10275, ZN => n10520);
   U10941 : NAND2_X1 port map( A1 => n19838, A2 => n20194, ZN => n4780);
   U10942 : NAND2_X1 port map( A1 => n25078, A2 => n22093, ZN => n4781);
   U10943 : INV_X1 port map( A => n4781, ZN => n21772);
   U10944 : OAI211_X1 port map( C1 => n22642, C2 => n22641, A => n22640, B => 
                           n4782, ZN => Ciphertext(118));
   U10946 : MUX2_X1 port map( A => n7660, B => n7659, S => n7947, Z => n4785);
   U10947 : AOI22_X1 port map( A1 => n9695, A2 => n10026, B1 => n9699, B2 => 
                           n9639, ZN => n4787);
   U10948 : OAI21_X2 port map( B1 => n4787, B2 => n9240, A => n9239, ZN => 
                           n11123);
   U10950 : NAND3_X1 port map( A1 => n4794, A2 => n14317, A3 => n13868, ZN => 
                           n4793);
   U10951 : NAND2_X1 port map( A1 => n14322, A2 => n14458, ZN => n4795);
   U10952 : NAND2_X2 port map( A1 => n5172, A2 => n5170, ZN => n14317);
   U10953 : NAND2_X1 port map( A1 => n12870, A2 => n13097, ZN => n4796);
   U10954 : NAND2_X1 port map( A1 => n12867, A2 => n13117, ZN => n4797);
   U10955 : NAND2_X1 port map( A1 => n4800, A2 => n7739, ZN => n4799);
   U10957 : INV_X1 port map( A => n8913, ZN => n4802);
   U10958 : OAI211_X2 port map( C1 => n4801, C2 => n7820, A => n6799, B => 
                           n7821, ZN => n8913);
   U10959 : NAND2_X1 port map( A1 => n8219, A2 => n7809, ZN => n4804);
   U10961 : NAND2_X1 port map( A1 => n14702, A2 => n24586, ZN => n4806);
   U10964 : OAI22_X1 port map( A1 => n19016, A2 => n19162, B1 => n19164, B2 => 
                           n4809, ZN => n18791);
   U10965 : XNOR2_X1 port map( A => n18434, B => n18478, ZN => n4810);
   U10967 : XNOR2_X1 port map( A => n18441, B => n18440, ZN => n19163);
   U10968 : NAND2_X1 port map( A1 => n7229, A2 => n7946, ZN => n4813);
   U10970 : INV_X1 port map( A => n10553, ZN => n4815);
   U10971 : NAND2_X1 port map( A1 => n16830, A2 => n17445, ZN => n4818);
   U10972 : NAND2_X1 port map( A1 => n12957, A2 => n13336, ZN => n4823);
   U10973 : XNOR2_X1 port map( A => n4821, B => n12105, ZN => n4820);
   U10974 : INV_X1 port map( A => n12106, ZN => n4821);
   U10975 : NAND2_X1 port map( A1 => n11022, A2 => n13775, ZN => n4824);
   U10976 : INV_X1 port map( A => n7358, ZN => n7415);
   U10977 : NAND2_X1 port map( A1 => n4827, A2 => n7358, ZN => n7994);
   U10978 : OR2_X1 port map( A1 => n6690, A2 => n6686, ZN => n4830);
   U10979 : INV_X1 port map( A => n9423, ZN => n9746);
   U10982 : NAND2_X1 port map( A1 => n4833, A2 => n9747, ZN => n4832);
   U10983 : AND2_X1 port map( A1 => n9991, A2 => n9990, ZN => n4833);
   U10985 : OAI21_X1 port map( B1 => n16383, B2 => n15656, A => n4835, ZN => 
                           n16387);
   U10987 : OAI22_X2 port map( A1 => n4837, A2 => n14236, B1 => n13994, B2 => 
                           n13930, ZN => n15112);
   U10988 : NAND2_X1 port map( A1 => n7022, A2 => n6846, ZN => n4839);
   U10989 : NAND3_X1 port map( A1 => n6001, A2 => n250, A3 => n4839, ZN => 
                           n4838);
   U10990 : AOI21_X1 port map( B1 => n16316, B2 => n17013, A => n4840, ZN => 
                           n16317);
   U10991 : INV_X1 port map( A => n17356, ZN => n4840);
   U10992 : OAI21_X1 port map( B1 => n19077, B2 => n24483, A => n4843, ZN => 
                           n4842);
   U10993 : NAND2_X1 port map( A1 => n24483, A2 => n19078, ZN => n4843);
   U10994 : INV_X1 port map( A => n21812, ZN => n4845);
   U10995 : NAND2_X1 port map( A1 => n22059, A2 => n22245, ZN => n21812);
   U10996 : NOR2_X1 port map( A1 => n21786, A2 => n4845, ZN => n21788);
   U10998 : NOR2_X1 port map( A1 => n7382, A2 => n7619, ZN => n4848);
   U10999 : OAI211_X2 port map( C1 => n4848, C2 => n7304, A => n7303, B => 
                           n7302, ZN => n8916);
   U11000 : INV_X1 port map( A => n12534, ZN => n4850);
   U11001 : NAND3_X1 port map( A1 => n401, A2 => n13051, A3 => n12534, ZN => 
                           n12443);
   U11002 : NAND2_X1 port map( A1 => n19211, A2 => n4853, ZN => n4852);
   U11004 : INV_X1 port map( A => n4854, ZN => n23762);
   U11005 : NAND2_X1 port map( A1 => n23767, A2 => n23769, ZN => n4854);
   U11006 : OAI22_X1 port map( A1 => n23783, A2 => n22523, B1 => n22524, B2 => 
                           n4854, ZN => n22526);
   U11007 : INV_X1 port map( A => n23769, ZN => n23778);
   U11008 : XNOR2_X1 port map( A => n18381, B => n4855, ZN => n16664);
   U11009 : XNOR2_X1 port map( A => n18381, B => n4856, ZN => n18013);
   U11010 : INV_X1 port map( A => n18183, ZN => n4856);
   U11011 : NAND2_X1 port map( A1 => n19210, A2 => n18816, ZN => n4857);
   U11012 : XNOR2_X1 port map( A => n15282, B => n15174, ZN => n4859);
   U11014 : NAND3_X1 port map( A1 => n23723, A2 => n23714, A3 => n23727, ZN => 
                           n4864);
   U11015 : NAND2_X1 port map( A1 => n23721, A2 => n23720, ZN => n22148);
   U11016 : XNOR2_X1 port map( A => n4862, B => n22150, ZN => Ciphertext(135));
   U11017 : NAND2_X1 port map( A1 => n438, A2 => n6295, ZN => n6211);
   U11018 : MUX2_X1 port map( A => n5946, B => n6173, S => n6174, Z => n5948);
   U11019 : NAND2_X1 port map( A1 => n16202, A2 => n16200, ZN => n4870);
   U11020 : MUX2_X1 port map( A => n11205, B => n11338, S => n11209, Z => n9645
                           );
   U11023 : NAND2_X1 port map( A1 => n264, A2 => n18841, ZN => n4874);
   U11024 : NAND2_X1 port map( A1 => n6174, A2 => n6335, ZN => n6176);
   U11026 : NAND2_X1 port map( A1 => n9880, A2 => n4993, ZN => n9252);
   U11028 : NAND2_X1 port map( A1 => n4878, A2 => n4881, ZN => n4880);
   U11029 : OAI21_X1 port map( B1 => n7647, B2 => n7761, A => n4879, ZN => 
                           n7766);
   U11030 : NAND2_X1 port map( A1 => n7646, A2 => n4880, ZN => n4879);
   U11031 : XNOR2_X1 port map( A => n18704, B => n4882, ZN => n17035);
   U11032 : XNOR2_X1 port map( A => n17900, B => n17817, ZN => n4882);
   U11033 : INV_X1 port map( A => n19237, ZN => n18863);
   U11034 : INV_X1 port map( A => n19112, ZN => n4884);
   U11035 : INV_X1 port map( A => n24310, ZN => n4885);
   U11036 : NAND2_X1 port map( A1 => n5446, A2 => n16269, ZN => n4886);
   U11037 : NAND2_X1 port map( A1 => n16270, A2 => n16271, ZN => n4887);
   U11038 : XNOR2_X1 port map( A => n18123, B => n18124, ZN => n18492);
   U11039 : XNOR2_X1 port map( A => n18184, B => n18492, ZN => n18127);
   U11040 : OAI21_X1 port map( B1 => n7228, B2 => n7080, A => n7943, ZN => 
                           n4889);
   U11041 : XNOR2_X1 port map( A => n18383, B => n1410, ZN => n4890);
   U11042 : OAI21_X1 port map( B1 => n25445, B2 => n4892, A => n4891, ZN => 
                           n4893);
   U11044 : NAND2_X1 port map( A1 => n14211, A2 => n24376, ZN => n4892);
   U11045 : AOI21_X2 port map( B1 => n4895, B2 => n1391, A => n4893, ZN => 
                           n14834);
   U11046 : INV_X1 port map( A => n24375, ZN => n4894);
   U11047 : NAND3_X1 port map( A1 => n16050, A2 => n294, A3 => n15606, ZN => 
                           n4900);
   U11048 : AOI21_X1 port map( B1 => n24574, B2 => n11111, A => n10868, ZN => 
                           n10877);
   U11049 : NAND2_X1 port map( A1 => n19704, A2 => n20615, ZN => n4991);
   U11050 : NAND2_X1 port map( A1 => n20616, A2 => n20617, ZN => n19704);
   U11051 : NAND2_X1 port map( A1 => n4902, A2 => n7376, ZN => n4901);
   U11052 : NAND2_X1 port map( A1 => n5432, A2 => n7735, ZN => n4902);
   U11053 : AOI22_X1 port map( A1 => n4904, A2 => n25240, B1 => n23866, B2 => 
                           n23857, ZN => n4903);
   U11054 : NAND3_X1 port map( A1 => n13093, A2 => n13096, A3 => n12871, ZN => 
                           n4907);
   U11055 : NAND2_X1 port map( A1 => n4910, A2 => n4912, ZN => n4909);
   U11056 : NAND2_X1 port map( A1 => n20117, A2 => n25034, ZN => n4910);
   U11057 : INV_X1 port map( A => n17951, ZN => n20848);
   U11058 : AOI21_X1 port map( B1 => n25262, B2 => n19883, A => n20109, ZN => 
                           n4912);
   U11059 : XNOR2_X1 port map( A => n9124, B => n4913, ZN => n9125);
   U11060 : XNOR2_X1 port map( A => n8236, B => n4913, ZN => n5504);
   U11061 : XNOR2_X1 port map( A => n8843, B => n4913, ZN => n8833);
   U11062 : NAND2_X1 port map( A1 => n15815, A2 => n4914, ZN => n15818);
   U11063 : NAND2_X1 port map( A1 => n4919, A2 => n19532, ZN => n4915);
   U11064 : INV_X1 port map( A => n19270, ZN => n19529);
   U11065 : NOR2_X1 port map( A1 => n24393, A2 => n4918, ZN => n4917);
   U11066 : INV_X1 port map( A => n19537, ZN => n4918);
   U11067 : OAI21_X1 port map( B1 => n19530, B2 => n19270, A => n19269, ZN => 
                           n4919);
   U11069 : INV_X1 port map( A => n6874, ZN => n4922);
   U11070 : NAND2_X1 port map( A1 => n314, A2 => n6767, ZN => n6878);
   U11071 : NAND2_X1 port map( A1 => n6876, A2 => n314, ZN => n6764);
   U11072 : NAND3_X1 port map( A1 => n6309, A2 => n6768, A3 => n314, ZN => 
                           n6312);
   U11073 : MUX2_X1 port map( A => n5855, B => n5854, S => n314, Z => n5858);
   U11075 : NOR2_X1 port map( A1 => n10942, A2 => n5392, ZN => n10513);
   U11076 : NOR2_X1 port map( A1 => n10571, A2 => n5392, ZN => n10572);
   U11077 : NAND2_X1 port map( A1 => n13109, A2 => n12856, ZN => n4925);
   U11078 : NAND2_X1 port map( A1 => n13265, A2 => n13267, ZN => n4930);
   U11079 : NOR2_X2 port map( A1 => n19046, A2 => n19045, ZN => n19979);
   U11080 : NAND2_X1 port map( A1 => n19977, A2 => n20140, ZN => n4933);
   U11081 : INV_X1 port map( A => n17485, ZN => n17733);
   U11082 : NOR2_X1 port map( A1 => n17485, A2 => n4934, ZN => n17484);
   U11083 : NAND2_X1 port map( A1 => n3978, A2 => n23531, ZN => n23009);
   U11084 : NAND3_X1 port map( A1 => n23013, A2 => n23533, A3 => n3978, ZN => 
                           n23024);
   U11085 : OR2_X2 port map( A1 => n9402, A2 => n9401, ZN => n11190);
   U11086 : NAND2_X1 port map( A1 => n10457, A2 => n10728, ZN => n4936);
   U11087 : NAND2_X1 port map( A1 => n4951, A2 => n10728, ZN => n4937);
   U11089 : NAND2_X1 port map( A1 => n4353, A2 => n14663, ZN => n4939);
   U11090 : INV_X1 port map( A => n14267, ZN => n14274);
   U11092 : NAND2_X1 port map( A1 => n12984, A2 => n12541, ZN => n4944);
   U11093 : INV_X1 port map( A => n13220, ZN => n4945);
   U11094 : INV_X1 port map( A => n23515, ZN => n4947);
   U11095 : MUX2_X1 port map( A => n22916, B => n4948, S => n22918, Z => n23515
                           );
   U11096 : OAI22_X1 port map( A1 => n21712, A2 => n22918, B1 => n22916, B2 => 
                           n22917, ZN => n4950);
   U11097 : AND2_X1 port map( A1 => n4951, A2 => n11190, ZN => n9403);
   U11098 : INV_X1 port map( A => n10730, ZN => n4951);
   U11099 : INV_X1 port map( A => n4957, ZN => n16304);
   U11101 : OAI22_X1 port map( A1 => n16300, A2 => n16299, B1 => n16303, B2 => 
                           n4957, ZN => n16308);
   U11102 : NAND2_X1 port map( A1 => n7666, A2 => n436, ZN => n6551);
   U11103 : NAND3_X1 port map( A1 => n7666, A2 => n436, A3 => n269, ZN => n8533
                           );
   U11104 : NAND2_X1 port map( A1 => n12925, A2 => n4958, ZN => n12609);
   U11105 : INV_X1 port map( A => n12899, ZN => n4958);
   U11107 : OAI21_X1 port map( B1 => n20317, B2 => n4961, A => n4960, ZN => 
                           n19716);
   U11108 : INV_X1 port map( A => n20316, ZN => n4961);
   U11109 : NAND2_X1 port map( A1 => n12898, A2 => n12897, ZN => n4964);
   U11110 : XNOR2_X1 port map( A => n14429, B => n14430, ZN => n4967);
   U11111 : OR2_X1 port map( A1 => n19128, A2 => n19304, ZN => n4968);
   U11113 : XNOR2_X1 port map( A => n4971, B => n25481, ZN => n18173);
   U11114 : NAND3_X1 port map( A1 => n16027, A2 => n2062, A3 => n4970, ZN => 
                           n4969);
   U11117 : OAI21_X1 port map( B1 => n24089, B2 => n6965, A => n4973, ZN => 
                           n7184);
   U11118 : NAND2_X1 port map( A1 => n19109, A2 => n25052, ZN => n4977);
   U11119 : XNOR2_X1 port map( A => n21463, B => n25040, ZN => n4978);
   U11120 : NOR2_X1 port map( A1 => n14168, A2 => n13742, ZN => n4980);
   U11122 : NAND2_X1 port map( A1 => n4982, A2 => n4981, ZN => n16950);
   U11123 : NAND2_X1 port map( A1 => n4984, A2 => n4983, ZN => n4982);
   U11124 : NAND2_X1 port map( A1 => n1382, A2 => n16417, ZN => n4983);
   U11125 : NAND2_X1 port map( A1 => n17289, A2 => n4986, ZN => n17541);
   U11126 : NAND3_X1 port map( A1 => n23079, A2 => n23064, A3 => n25024, ZN => 
                           n4989);
   U11129 : NAND2_X1 port map( A1 => n4991, A2 => n24338, ZN => n19873);
   U11130 : NAND2_X1 port map( A1 => n13171, A2 => n3688, ZN => n4992);
   U11131 : INV_X1 port map( A => n10534, ZN => n11884);
   U11132 : NAND4_X1 port map( A1 => n6808, A2 => n6807, A3 => n6809, A4 => 
                           n4994, ZN => n6810);
   U11133 : XNOR2_X1 port map( A => n12106, B => n11849, ZN => n4996);
   U11134 : NAND2_X1 port map( A1 => n1357, A2 => n10534, ZN => n10308);
   U11135 : NAND2_X1 port map( A1 => n1357, A2 => n4997, ZN => n10965);
   U11136 : AND2_X1 port map( A1 => n10534, A2 => n24479, ZN => n4997);
   U11138 : OR2_X1 port map( A1 => n6392, A2 => n6238, ZN => n5002);
   U11139 : XNOR2_X2 port map( A => n18210, B => n18211, ZN => n19526);
   U11140 : NAND2_X1 port map( A1 => n19523, A2 => n19284, ZN => n5496);
   U11141 : NAND2_X1 port map( A1 => n19526, A2 => n19522, ZN => n5003);
   U11142 : INV_X1 port map( A => n9064, ZN => n10058);
   U11143 : INV_X1 port map( A => n10052, ZN => n5004);
   U11144 : NAND2_X1 port map( A1 => n19433, A2 => n25423, ZN => n5006);
   U11145 : NAND2_X1 port map( A1 => n19438, A2 => n18834, ZN => n19433);
   U11147 : NAND2_X1 port map( A1 => n21958, A2 => n21959, ZN => n21961);
   U11149 : XNOR2_X1 port map( A => n295, B => n15244, ZN => n5009);
   U11150 : NAND2_X1 port map( A1 => n13064, A2 => n5011, ZN => n5010);
   U11151 : XNOR2_X1 port map( A => n8595, B => n8594, ZN => n9481);
   U11152 : XNOR2_X1 port map( A => n5014, B => n2241, ZN => n8777);
   U11153 : XNOR2_X1 port map( A => n8446, B => n5014, ZN => n8447);
   U11154 : XNOR2_X1 port map( A => n8172, B => n5014, ZN => n8174);
   U11158 : INV_X1 port map( A => n14188, ZN => n5020);
   U11160 : OR2_X1 port map( A1 => n12694, A2 => n13292, ZN => n5021);
   U11161 : NAND2_X1 port map( A1 => n19691, A2 => n20316, ZN => n19692);
   U11163 : NAND2_X1 port map( A1 => n12650, A2 => n12505, ZN => n5022);
   U11164 : INV_X1 port map( A => n17607, ZN => n16942);
   U11165 : NAND2_X1 port map( A1 => n5066, A2 => n5065, ZN => n5064);
   U11166 : NAND2_X1 port map( A1 => n10090, A2 => n24505, ZN => n5026);
   U11168 : MUX2_X1 port map( A => n13294, B => n13295, S => n12827, Z => 
                           n13296);
   U11172 : NAND2_X1 port map( A1 => n5033, A2 => n5030, ZN => n5029);
   U11173 : NOR2_X1 port map( A1 => n23089, A2 => n5131, ZN => n5030);
   U11174 : NAND4_X1 port map( A1 => n5035, A2 => n24941, A3 => n20975, A4 => 
                           n5037, ZN => n5031);
   U11175 : OR2_X1 port map( A1 => n23112, A2 => n24993, ZN => n5037);
   U11176 : NAND3_X1 port map( A1 => n23089, A2 => n24498, A3 => n5131, ZN => 
                           n5032);
   U11177 : NAND2_X1 port map( A1 => n5040, A2 => n5038, ZN => n16486);
   U11178 : NAND2_X1 port map( A1 => n16482, A2 => n15951, ZN => n5040);
   U11179 : AND2_X1 port map( A1 => n13231, A2 => n5041, ZN => n13232);
   U11180 : NAND2_X1 port map( A1 => n9443, A2 => n10584, ZN => n5042);
   U11181 : NAND2_X1 port map( A1 => n5042, A2 => n10317, ZN => n10319);
   U11182 : OAI22_X1 port map( A1 => n5042, A2 => n25507, B1 => n10370, B2 => 
                           n10372, ZN => n9215);
   U11183 : OAI211_X1 port map( C1 => n20426, C2 => n276, A => n24883, B => 
                           n5044, ZN => n5043);
   U11186 : OR2_X1 port map( A1 => n22592, A2 => n22317, ZN => n5046);
   U11187 : NAND2_X1 port map( A1 => n21378, A2 => n274, ZN => n5047);
   U11189 : NAND3_X1 port map( A1 => n23143, A2 => n1349, A3 => n22442, ZN => 
                           n5049);
   U11190 : NAND2_X1 port map( A1 => n7129, A2 => n7606, ZN => n5050);
   U11191 : INV_X1 port map( A => n7893, ZN => n5051);
   U11192 : NOR2_X1 port map( A1 => n16844, A2 => n5052, ZN => n17467);
   U11193 : NAND2_X1 port map( A1 => n5054, A2 => n5051, ZN => n5053);
   U11194 : NAND2_X1 port map( A1 => n7609, A2 => n7604, ZN => n7889);
   U11195 : NAND2_X1 port map( A1 => n7894, A2 => n7893, ZN => n5055);
   U11196 : NOR2_X1 port map( A1 => n5056, A2 => n17130, ZN => n17129);
   U11197 : INV_X1 port map( A => n25225, ZN => n5056);
   U11199 : NOR2_X1 port map( A1 => n10487, A2 => n10486, ZN => n5060);
   U11200 : NAND2_X1 port map( A1 => n10488, A2 => n5060, ZN => n5059);
   U11201 : NAND2_X1 port map( A1 => n5730, A2 => n10614, ZN => n5061);
   U11202 : NAND2_X1 port map( A1 => n10531, A2 => n304, ZN => n5063);
   U11203 : NAND3_X1 port map( A1 => n10465, A2 => n10855, A3 => n10858, ZN => 
                           n10466);
   U11204 : NAND2_X1 port map( A1 => n9456, A2 => n9565, ZN => n5065);
   U11206 : NOR2_X1 port map( A1 => n16832, A2 => n17152, ZN => n16834);
   U11210 : NAND2_X1 port map( A1 => n18734, A2 => n19477, ZN => n5070);
   U11211 : OAI21_X1 port map( B1 => n20173, B2 => n19803, A => n5071, ZN => 
                           n19508);
   U11212 : NAND2_X1 port map( A1 => n19507, A2 => n20173, ZN => n5071);
   U11213 : NAND2_X1 port map( A1 => n5072, A2 => n16980, ZN => n5073);
   U11214 : INV_X1 port map( A => n17450, ZN => n5072);
   U11216 : INV_X1 port map( A => n23765, ZN => n23766);
   U11217 : NAND2_X1 port map( A1 => n23779, A2 => n23757, ZN => n23765);
   U11219 : NAND2_X1 port map( A1 => n21793, A2 => n22231, ZN => n5076);
   U11220 : NAND2_X1 port map( A1 => n5077, A2 => n1481, ZN => n5078);
   U11221 : NAND2_X1 port map( A1 => n5078, A2 => n11127, ZN => n12219);
   U11222 : NAND2_X1 port map( A1 => n13953, A2 => n13954, ZN => n5079);
   U11223 : INV_X1 port map( A => n13954, ZN => n5080);
   U11224 : NAND2_X1 port map( A1 => n395, A2 => n13953, ZN => n13718);
   U11225 : NAND2_X1 port map( A1 => n14156, A2 => n395, ZN => n13719);
   U11226 : NAND2_X1 port map( A1 => n5081, A2 => n23256, ZN => n22649);
   U11227 : NAND2_X1 port map( A1 => n425, A2 => n25454, ZN => n9298);
   U11228 : OR2_X1 port map( A1 => n5082, A2 => n1348, ZN => n8574);
   U11229 : NAND2_X1 port map( A1 => n5083, A2 => n10089, ZN => n10091);
   U11230 : NAND2_X1 port map( A1 => n9779, A2 => n8571, ZN => n5083);
   U11231 : OAI21_X1 port map( B1 => n9780, B2 => n25454, A => n425, ZN => 
                           n9674);
   U11232 : INV_X1 port map( A => n5084, ZN => n21885);
   U11233 : NAND2_X1 port map( A1 => n5084, A2 => n22396, ZN => n22267);
   U11234 : NOR2_X1 port map( A1 => n22261, A2 => n5084, ZN => n22264);
   U11235 : AOI21_X1 port map( B1 => n22398, B2 => n5084, A => n22265, ZN => 
                           n21914);
   U11236 : MUX2_X1 port map( A => n22400, B => n5084, S => n25381, Z => n22136
                           );
   U11237 : AND2_X1 port map( A1 => n7023, A2 => n7025, ZN => n5088);
   U11238 : NAND2_X1 port map( A1 => n5089, A2 => n7027, ZN => n5086);
   U11241 : XNOR2_X1 port map( A => n18290, B => n24886, ZN => n17792);
   U11242 : XNOR2_X1 port map( A => n24886, B => n2319, ZN => n18460);
   U11243 : NAND2_X1 port map( A1 => n10772, A2 => n11101, ZN => n10218);
   U11244 : NAND2_X1 port map( A1 => n11031, A2 => n10772, ZN => n11034);
   U11245 : OAI22_X1 port map( A1 => n1552, A2 => n10772, B1 => n24753, B2 => 
                           n415, ZN => n11035);
   U11246 : NAND2_X1 port map( A1 => n23194, A2 => n24889, ZN => n5090);
   U11247 : INV_X1 port map( A => n11684, ZN => n12891);
   U11248 : NAND2_X1 port map( A1 => n19442, A2 => n20588, ZN => n5091);
   U11249 : NAND2_X1 port map( A1 => n5094, A2 => n5093, ZN => n5092);
   U11251 : AND3_X2 port map( A1 => n5670, A2 => n19416, A3 => n5669, ZN => 
                           n20586);
   U11252 : NAND3_X1 port map( A1 => n5218, A2 => n23974, A3 => n5095, ZN => 
                           n5217);
   U11253 : NAND2_X1 port map( A1 => n1488, A2 => n24440, ZN => n5095);
   U11254 : NAND2_X1 port map( A1 => n5098, A2 => n5096, ZN => n16234);
   U11255 : NOR2_X1 port map( A1 => n16491, A2 => n16232, ZN => n5097);
   U11256 : NAND2_X1 port map( A1 => n16233, A2 => n16232, ZN => n5098);
   U11258 : NAND2_X1 port map( A1 => n5100, A2 => n16100, ZN => n16104);
   U11261 : NAND2_X1 port map( A1 => n15576, A2 => n5104, ZN => n5103);
   U11262 : OAI211_X1 port map( C1 => n10699, C2 => n2754, A => n5109, B => 
                           n10955, ZN => n5108);
   U11263 : NAND2_X1 port map( A1 => n10699, A2 => n10548, ZN => n5109);
   U11264 : NAND2_X1 port map( A1 => n5111, A2 => n5110, ZN => n14172);
   U11265 : NAND2_X1 port map( A1 => n5113, A2 => n5112, ZN => n5110);
   U11266 : NAND2_X1 port map( A1 => n12441, A2 => n12737, ZN => n5111);
   U11268 : NAND2_X1 port map( A1 => n5115, A2 => n20060, ZN => n5114);
   U11270 : NOR2_X1 port map( A1 => n7221, A2 => n5117, ZN => n5116);
   U11271 : INV_X1 port map( A => n7222, ZN => n5117);
   U11273 : NAND2_X1 port map( A1 => n11062, A2 => n11070, ZN => n5119);
   U11274 : XNOR2_X1 port map( A => n5120, B => n2743, ZN => n18570);
   U11275 : XNOR2_X1 port map( A => n5120, B => n18295, ZN => n18087);
   U11276 : XNOR2_X1 port map( A => n5120, B => n18188, ZN => n15810);
   U11277 : NAND2_X1 port map( A1 => n13227, A2 => n13224, ZN => n13225);
   U11278 : INV_X1 port map( A => n25367, ZN => n20822);
   U11279 : NOR2_X1 port map( A1 => n20803, A2 => n21928, ZN => n5121);
   U11280 : XNOR2_X1 port map( A => n21647, B => n21106, ZN => n21184);
   U11282 : XNOR2_X1 port map( A => n21184, B => n5124, ZN => n20978);
   U11283 : XNOR2_X1 port map( A => n21332, B => n5125, ZN => n5124);
   U11284 : NAND2_X1 port map( A1 => n5127, A2 => n5129, ZN => n5125);
   U11285 : OAI21_X1 port map( B1 => n19260, B2 => n5131, A => n5126, ZN => 
                           n5128);
   U11286 : NAND3_X1 port map( A1 => n276, A2 => n24463, A3 => n20975, ZN => 
                           n5126);
   U11287 : INV_X1 port map( A => n5128, ZN => n5127);
   U11288 : NAND2_X1 port map( A1 => n5130, A2 => n19260, ZN => n5129);
   U11289 : NAND2_X1 port map( A1 => n19260, A2 => n5132, ZN => n21583);
   U11291 : OAI21_X1 port map( B1 => n19589, B2 => n5134, A => n19588, ZN => 
                           n19593);
   U11292 : NOR2_X1 port map( A1 => n24422, A2 => n13323, ZN => n13326);
   U11293 : OAI21_X1 port map( B1 => n12062, B2 => n5140, A => n5137, ZN => 
                           n5141);
   U11294 : NOR2_X1 port map( A1 => n3256, A2 => n13323, ZN => n5138);
   U11295 : INV_X1 port map( A => n24422, ZN => n5139);
   U11296 : NAND3_X1 port map( A1 => n416, A2 => n10941, A3 => n3760, ZN => 
                           n10379);
   U11297 : INV_X1 port map( A => n441, ZN => n5144);
   U11298 : XNOR2_X1 port map( A => n21455, B => n1891, ZN => n21260);
   U11300 : OAI21_X2 port map( B1 => n5148, B2 => n5146, A => n5145, ZN => 
                           n7628);
   U11301 : NAND2_X1 port map( A1 => n5147, A2 => n7007, ZN => n5146);
   U11302 : NAND2_X1 port map( A1 => n6647, A2 => n7008, ZN => n5147);
   U11303 : INV_X1 port map( A => n18428, ZN => n5149);
   U11304 : NAND2_X1 port map( A1 => n19164, A2 => n18788, ZN => n18428);
   U11305 : XNOR2_X1 port map( A => n18388, B => n17663, ZN => n18413);
   U11306 : INV_X1 port map( A => n14327, ZN => n5151);
   U11307 : NAND3_X1 port map( A1 => n5151, A2 => n13864, A3 => n14044, ZN => 
                           n5150);
   U11308 : AOI21_X1 port map( B1 => n25072, B2 => n1443, A => n5153, ZN => 
                           n5152);
   U11309 : NOR2_X1 port map( A1 => n280, A2 => n19578, ZN => n5153);
   U11310 : NAND2_X1 port map( A1 => n12931, A2 => n12897, ZN => n5156);
   U11311 : XNOR2_X1 port map( A => n8297, B => n8034, ZN => n5157);
   U11313 : OAI21_X1 port map( B1 => n19476, B2 => n18734, A => n19478, ZN => 
                           n17640);
   U11315 : XNOR2_X1 port map( A => n18372, B => n17710, ZN => n5160);
   U11316 : NAND2_X1 port map( A1 => n311, A2 => n7604, ZN => n7324);
   U11318 : NOR2_X2 port map( A1 => n15678, A2 => n5164, ZN => n17326);
   U11319 : NAND2_X1 port map( A1 => n5166, A2 => n5165, ZN => n5164);
   U11320 : NAND2_X1 port map( A1 => n15675, A2 => n16328, ZN => n5166);
   U11321 : INV_X1 port map( A => n16232, ZN => n15933);
   U11322 : OAI21_X1 port map( B1 => n5169, B2 => n15932, A => n5168, ZN => 
                           n5167);
   U11323 : AOI21_X1 port map( B1 => n5405, B2 => n20134, A => n5566, ZN => 
                           n5404);
   U11324 : NAND3_X1 port map( A1 => n12873, A2 => n12872, A3 => n13123, ZN => 
                           n5170);
   U11325 : NAND2_X1 port map( A1 => n12875, A2 => n5624, ZN => n5172);
   U11326 : OAI21_X1 port map( B1 => n13305, B2 => n12555, A => n5173, ZN => 
                           n5175);
   U11327 : NAND2_X1 port map( A1 => n12555, A2 => n12611, ZN => n5173);
   U11328 : NAND2_X1 port map( A1 => n16115, A2 => n16120, ZN => n5177);
   U11329 : XNOR2_X1 port map( A => n5179, B => n8755, ZN => n5255);
   U11330 : XNOR2_X1 port map( A => n5179, B => n9052, ZN => n9054);
   U11331 : XNOR2_X1 port map( A => n5179, B => n8754, ZN => n8559);
   U11332 : XNOR2_X1 port map( A => n5179, B => n9190, ZN => n8121);
   U11334 : MUX2_X1 port map( A => n20118, B => n25514, S => n19883, Z => 
                           n19718);
   U11335 : INV_X1 port map( A => n11433, ZN => n12376);
   U11336 : XNOR2_X1 port map( A => n5180, B => n10689, ZN => n11343);
   U11337 : XNOR2_X1 port map( A => n5181, B => n10689, ZN => n11658);
   U11338 : XNOR2_X1 port map( A => n10689, B => n5182, ZN => n12011);
   U11339 : XNOR2_X1 port map( A => n5183, B => n8734, ZN => n7310);
   U11340 : INV_X1 port map( A => n8329, ZN => n5183);
   U11341 : XNOR2_X1 port map( A => n8734, B => n5184, ZN => n8357);
   U11343 : NAND2_X1 port map( A1 => n20410, A2 => n20411, ZN => n5187);
   U11344 : NAND2_X1 port map( A1 => n20409, A2 => n20264, ZN => n5188);
   U11345 : INV_X1 port map( A => n22452, ZN => n5190);
   U11346 : NAND2_X1 port map( A1 => n5191, A2 => n12626, ZN => n12627);
   U11347 : MUX2_X1 port map( A => n16100, B => n16101, S => n15583, Z => 
                           n16103);
   U11348 : NAND2_X1 port map( A1 => n8005, A2 => n7292, ZN => n7541);
   U11349 : XNOR2_X1 port map( A => n22006, B => n2805, ZN => n21752);
   U11350 : NAND2_X1 port map( A1 => n20362, A2 => n24078, ZN => n5193);
   U11354 : INV_X1 port map( A => n24909, ZN => n5196);
   U11355 : OAI21_X1 port map( B1 => n17764, B2 => n5196, A => n17763, ZN => 
                           n17765);
   U11356 : INV_X1 port map( A => n10505, ZN => n5198);
   U11357 : NAND2_X1 port map( A1 => n9809, A2 => n9338, ZN => n5199);
   U11358 : INV_X1 port map( A => n5200, ZN => n15374);
   U11359 : XNOR2_X1 port map( A => n5200, B => n14454, ZN => n14456);
   U11360 : OAI21_X1 port map( B1 => n12816, B2 => n12815, A => n12814, ZN => 
                           n5200);
   U11361 : XNOR2_X1 port map( A => n15374, B => n3232, ZN => n14547);
   U11362 : NAND3_X1 port map( A1 => n24908, A2 => n19389, A3 => n25052, ZN => 
                           n19111);
   U11363 : OAI21_X1 port map( B1 => n5202, B2 => n432, A => n5201, ZN => n5204
                           );
   U11364 : NAND2_X1 port map( A1 => n432, A2 => n7292, ZN => n5201);
   U11365 : XNOR2_X1 port map( A => n21043, B => n641, ZN => n5339);
   U11366 : XNOR2_X1 port map( A => n5210, B => n15477, ZN => n5513);
   U11367 : XNOR2_X1 port map( A => n5210, B => n14374, ZN => n14375);
   U11368 : XNOR2_X1 port map( A => n5210, B => n13691, ZN => n13710);
   U11369 : NOR2_X1 port map( A1 => n15646, A2 => n24061, ZN => n5211);
   U11370 : OAI21_X1 port map( B1 => n19326, B2 => n24516, A => n19329, ZN => 
                           n17945);
   U11371 : OAI211_X1 port map( C1 => n19328, C2 => n18933, A => n19326, B => 
                           n24516, ZN => n17498);
   U11373 : AOI21_X1 port map( B1 => n19330, B2 => n24516, A => n5213, ZN => 
                           n19332);
   U11374 : NAND2_X1 port map( A1 => n18938, A2 => n24583, ZN => n18853);
   U11377 : INV_X1 port map( A => n13532, ZN => n5216);
   U11378 : XNOR2_X1 port map( A => n5217, B => n450, ZN => Ciphertext(186));
   U11379 : NAND2_X1 port map( A1 => n5220, A2 => n5219, ZN => n5218);
   U11380 : NAND2_X1 port map( A1 => n23984, A2 => n24014, ZN => n5219);
   U11381 : OAI21_X1 port map( B1 => n24448, B2 => n23978, A => n23993, ZN => 
                           n5220);
   U11382 : NAND2_X1 port map( A1 => n22322, A2 => n24496, ZN => n5222);
   U11383 : NAND2_X1 port map( A1 => n23228, A2 => n23227, ZN => n23221);
   U11384 : INV_X1 port map( A => n21766, ZN => n22064);
   U11386 : NAND2_X1 port map( A1 => n15958, A2 => n5229, ZN => n17434);
   U11387 : AND2_X1 port map( A1 => n16170, A2 => n16426, ZN => n5229);
   U11388 : NAND2_X1 port map( A1 => n15958, A2 => n16170, ZN => n16172);
   U11389 : NAND2_X1 port map( A1 => n21917, A2 => n1352, ZN => n5231);
   U11390 : NOR2_X1 port map( A1 => n329, A2 => n22455, ZN => n21917);
   U11391 : NAND2_X1 port map( A1 => n9468, A2 => n9963, ZN => n5232);
   U11392 : NAND2_X1 port map( A1 => n19036, A2 => n19451, ZN => n5234);
   U11393 : OAI211_X2 port map( C1 => n17561, C2 => n5238, A => n5237, B => 
                           n17560, ZN => n20316);
   U11394 : NAND3_X1 port map( A1 => n4554, A2 => n5243, A3 => n5242, ZN => 
                           n5241);
   U11395 : AOI21_X1 port map( B1 => n16100, B2 => n16101, A => n15583, ZN => 
                           n15632);
   U11396 : NAND2_X1 port map( A1 => n15780, A2 => n15583, ZN => n16681);
   U11397 : NAND2_X1 port map( A1 => n5458, A2 => n5245, ZN => n5459);
   U11398 : INV_X1 port map( A => n10623, ZN => n10669);
   U11399 : NAND2_X1 port map( A1 => n5824, A2 => n6473, ZN => n5249);
   U11401 : NAND2_X1 port map( A1 => n13392, A2 => n13975, ZN => n5252);
   U11402 : AOI21_X1 port map( B1 => n13391, B2 => n13974, A => n13390, ZN => 
                           n5253);
   U11403 : OAI21_X2 port map( B1 => n5254, B2 => n9316, A => n9317, ZN => 
                           n11128);
   U11404 : OAI21_X1 port map( B1 => n422, B2 => n9989, A => n25444, ZN => 
                           n5254);
   U11405 : XNOR2_X1 port map( A => n5255, B => n8672, ZN => n8679);
   U11406 : NAND2_X1 port map( A1 => n14320, A2 => n13868, ZN => n5256);
   U11408 : NAND2_X1 port map( A1 => n22591, A2 => n21921, ZN => n5258);
   U11409 : OAI211_X2 port map( C1 => n20311, C2 => n25101, A => n5262, B => 
                           n5261, ZN => n21324);
   U11410 : NAND3_X1 port map( A1 => n20309, A2 => n25101, A3 => n20549, ZN => 
                           n5261);
   U11412 : NAND2_X1 port map( A1 => n20309, A2 => n20549, ZN => n20544);
   U11413 : INV_X1 port map( A => n7175, ZN => n5264);
   U11414 : NAND2_X1 port map( A1 => n7418, A2 => n7789, ZN => n7175);
   U11415 : NAND2_X1 port map( A1 => n5264, A2 => n7782, ZN => n5263);
   U11416 : NAND3_X1 port map( A1 => n5267, A2 => n5266, A3 => n7783, ZN => 
                           n5265);
   U11417 : NAND2_X1 port map( A1 => n7784, A2 => n7787, ZN => n5267);
   U11418 : NAND2_X1 port map( A1 => n7420, A2 => n7419, ZN => n5268);
   U11419 : AOI21_X1 port map( B1 => n6468, B2 => n6469, A => n6467, ZN => 
                           n5270);
   U11420 : NAND3_X1 port map( A1 => n7638, A2 => n312, A3 => n7915, ZN => 
                           n7396);
   U11421 : NAND2_X1 port map( A1 => n9670, A2 => n9669, ZN => n5273);
   U11422 : NOR2_X1 port map( A1 => n9730, A2 => n9729, ZN => n5275);
   U11423 : NAND2_X1 port map( A1 => n10020, A2 => n5275, ZN => n5274);
   U11424 : NAND2_X1 port map( A1 => n9650, A2 => n9730, ZN => n5276);
   U11425 : NAND2_X1 port map( A1 => n9730, A2 => n25475, ZN => n5278);
   U11426 : NOR2_X1 port map( A1 => n5280, A2 => n20388, ZN => n20387);
   U11427 : NOR2_X1 port map( A1 => n5280, A2 => n19490, ZN => n19349);
   U11428 : NAND3_X1 port map( A1 => n25473, A2 => n19490, A3 => n5280, ZN => 
                           n19492);
   U11429 : OAI21_X1 port map( B1 => n23728, B2 => n24381, A => n5286, ZN => 
                           n5283);
   U11430 : NAND3_X1 port map( A1 => n22091, A2 => n5282, A3 => n5281, ZN => 
                           n5285);
   U11431 : NAND3_X1 port map( A1 => n5284, A2 => n24374, A3 => n23714, ZN => 
                           n5281);
   U11432 : INV_X1 port map( A => n5283, ZN => n5282);
   U11434 : OR2_X1 port map( A1 => n22091, A2 => Key(60), ZN => n5287);
   U11435 : NAND2_X1 port map( A1 => n5289, A2 => n9372, ZN => n5288);
   U11436 : NAND2_X1 port map( A1 => n19302, A2 => n19128, ZN => n5290);
   U11438 : NAND2_X1 port map( A1 => n7053, A2 => n7803, ZN => n5291);
   U11439 : OAI211_X2 port map( C1 => n7434, C2 => n7054, A => n5294, B => 
                           n5292, ZN => n8896);
   U11440 : OR2_X1 port map( A1 => n5293, A2 => n7795, ZN => n5292);
   U11441 : NAND2_X1 port map( A1 => n7798, A2 => n7166, ZN => n5293);
   U11442 : NAND2_X1 port map( A1 => n7166, A2 => n6280, ZN => n7053);
   U11443 : NAND2_X1 port map( A1 => n17173, A2 => n16434, ZN => n16432);
   U11444 : NAND2_X1 port map( A1 => n13478, A2 => n5299, ZN => n5298);
   U11445 : XNOR2_X1 port map( A => n5300, B => n16037, ZN => n5302);
   U11446 : XNOR2_X1 port map( A => n18374, B => n18513, ZN => n5304);
   U11447 : NAND2_X1 port map( A1 => n16970, A2 => n16969, ZN => n5305);
   U11448 : NOR2_X1 port map( A1 => n22506, A2 => n22528, ZN => n5306);
   U11449 : NAND2_X1 port map( A1 => n3240, A2 => n19849, ZN => n19855);
   U11450 : INV_X1 port map( A => n12683, ZN => n5311);
   U11452 : NOR2_X1 port map( A1 => n2561, A2 => n5316, ZN => n5315);
   U11453 : NAND2_X1 port map( A1 => n5318, A2 => n7761, ZN => n5689);
   U11454 : INV_X1 port map( A => n13094, ZN => n12649);
   U11455 : XNOR2_X2 port map( A => n9680, B => n9679, ZN => n13094);
   U11456 : NAND2_X1 port map( A1 => n5319, A2 => n5325, ZN => n13675);
   U11457 : NAND2_X1 port map( A1 => n5320, A2 => n5323, ZN => n5319);
   U11458 : NAND2_X1 port map( A1 => n5322, A2 => n5321, ZN => n5320);
   U11459 : NAND2_X1 port map( A1 => n12649, A2 => n12648, ZN => n5322);
   U11460 : INV_X1 port map( A => n12648, ZN => n5324);
   U11461 : NOR2_X2 port map( A1 => n13791, A2 => n5330, ZN => n15484);
   U11463 : XNOR2_X1 port map( A => n14898, B => n1411, ZN => n5331);
   U11464 : NAND2_X1 port map( A1 => n5333, A2 => n5709, ZN => n5332);
   U11465 : AND2_X1 port map( A1 => n13565, A2 => n14108, ZN => n5709);
   U11466 : NAND2_X1 port map( A1 => n19061, A2 => n24982, ZN => n5337);
   U11467 : NAND2_X1 port map( A1 => n9390, A2 => n9389, ZN => n5341);
   U11468 : NAND2_X1 port map( A1 => n25203, A2 => n11069, ZN => n5342);
   U11469 : XNOR2_X1 port map( A => n5344, B => n7161, ZN => n8430);
   U11470 : XNOR2_X1 port map( A => n5346, B => n7161, ZN => n8149);
   U11471 : INV_X1 port map( A => n22493, ZN => n5347);
   U11472 : NAND3_X1 port map( A1 => n5349, A2 => n22528, A3 => n23443, ZN => 
                           n5348);
   U11473 : NAND2_X1 port map( A1 => n22491, A2 => n22733, ZN => n5350);
   U11474 : NAND2_X1 port map( A1 => n23442, A2 => n25042, ZN => n22527);
   U11475 : INV_X1 port map( A => n10871, ZN => n5352);
   U11476 : OAI21_X1 port map( B1 => n11115, B2 => n11117, A => n5351, ZN => 
                           n10878);
   U11477 : NAND2_X1 port map( A1 => n5357, A2 => n10120, ZN => n5356);
   U11478 : NAND2_X1 port map( A1 => n24096, A2 => n5359, ZN => n11837);
   U11479 : NAND3_X1 port map( A1 => n23810, A2 => n25391, A3 => n23811, ZN => 
                           n22540);
   U11480 : NAND2_X1 port map( A1 => n10114, A2 => n9338, ZN => n5362);
   U11482 : NOR2_X1 port map( A1 => n20600, A2 => n5364, ZN => n5363);
   U11483 : NOR2_X1 port map( A1 => n276, A2 => n5365, ZN => n5364);
   U11484 : NAND2_X1 port map( A1 => n266, A2 => n17356, ZN => n5367);
   U11485 : INV_X1 port map( A => n12533, ZN => n5368);
   U11486 : XNOR2_X1 port map( A => n24337, B => n18499, ZN => n18225);
   U11487 : XNOR2_X1 port map( A => n17850, B => n18289, ZN => n5369);
   U11488 : OAI211_X1 port map( C1 => n19322, C2 => n19472, A => n19467, B => 
                           n18959, ZN => n19323);
   U11489 : NAND2_X1 port map( A1 => n18959, A2 => n17872, ZN => n18962);
   U11490 : OAI21_X1 port map( B1 => n19467, B2 => n18959, A => n19466, ZN => 
                           n19468);
   U11492 : AND2_X1 port map( A1 => n19314, A2 => n5370, ZN => n19320);
   U11493 : NAND3_X1 port map( A1 => n19309, A2 => n24912, A3 => n5371, ZN => 
                           n5370);
   U11494 : NAND2_X1 port map( A1 => n5372, A2 => n9493, ZN => n10776);
   U11496 : NAND2_X1 port map( A1 => n5372, A2 => n9732, ZN => n9733);
   U11497 : INV_X1 port map( A => n18397, ZN => n18284);
   U11498 : XNOR2_X1 port map( A => n18397, B => n5374, ZN => n5373);
   U11499 : INV_X1 port map( A => n16551, ZN => n5375);
   U11500 : AOI22_X1 port map( A1 => n16554, A2 => n16553, B1 => n16552, B2 => 
                           n5376, ZN => n17680);
   U11501 : INV_X1 port map( A => n5378, ZN => n22370);
   U11502 : NAND2_X1 port map( A1 => n5378, A2 => n22769, ZN => n21292);
   U11503 : NAND2_X1 port map( A1 => n22680, A2 => n5378, ZN => n20605);
   U11504 : AOI21_X1 port map( B1 => n5378, B2 => n22770, A => n22769, ZN => 
                           n22775);
   U11505 : AOI21_X1 port map( B1 => n22773, B2 => n22772, A => n5378, ZN => 
                           n5611);
   U11507 : NAND3_X1 port map( A1 => n1552, A2 => n415, A3 => n11101, ZN => 
                           n5379);
   U11508 : OAI21_X1 port map( B1 => n11101, B2 => n5380, A => n10912, ZN => 
                           n5381);
   U11509 : NAND2_X1 port map( A1 => n1552, A2 => n10772, ZN => n5380);
   U11511 : NAND3_X1 port map( A1 => n15773, A2 => n16024, A3 => n5383, ZN => 
                           n15776);
   U11512 : NAND2_X1 port map( A1 => n5385, A2 => n16923, ZN => n5384);
   U11513 : NOR2_X1 port map( A1 => n17320, A2 => n16927, ZN => n5385);
   U11514 : AND2_X1 port map( A1 => n16809, A2 => n17077, ZN => n5386);
   U11515 : AND2_X1 port map( A1 => n7364, A2 => n7909, ZN => n5387);
   U11517 : NAND2_X1 port map( A1 => n7365, A2 => n7908, ZN => n5389);
   U11519 : NAND2_X1 port map( A1 => n10574, A2 => n11039, ZN => n5393);
   U11520 : AOI21_X1 port map( B1 => n25071, B2 => n24893, A => n323, ZN => 
                           n5396);
   U11521 : AOI22_X1 port map( A1 => n22710, A2 => n323, B1 => n5397, B2 => 
                           n5396, ZN => n5398);
   U11522 : XNOR2_X1 port map( A => n5398, B => n3798, ZN => Ciphertext(110));
   U11523 : XNOR2_X1 port map( A => n5399, B => n21079, ZN => Ciphertext(125));
   U11524 : OAI211_X1 port map( C1 => n21078, C2 => n23650, A => n5401, B => 
                           n5400, ZN => n5399);
   U11525 : NAND3_X1 port map( A1 => n23637, A2 => n23640, A3 => n23629, ZN => 
                           n5400);
   U11526 : NAND2_X1 port map( A1 => n23651, A2 => n23649, ZN => n5401);
   U11530 : NAND2_X1 port map( A1 => n15259, A2 => n25323, ZN => n5407);
   U11531 : NAND2_X1 port map( A1 => n16191, A2 => n16197, ZN => n15901);
   U11532 : INV_X1 port map( A => n17424, ZN => n5409);
   U11533 : OAI21_X1 port map( B1 => n12861, B2 => n12636, A => n5410, ZN => 
                           n12638);
   U11534 : NAND2_X1 port map( A1 => n12636, A2 => n13345, ZN => n5410);
   U11535 : NAND2_X1 port map( A1 => n5731, A2 => n5412, ZN => n5411);
   U11536 : OR2_X1 port map( A1 => n7583, A2 => n7584, ZN => n5490);
   U11537 : NAND3_X1 port map( A1 => n7475, A2 => n7952, A3 => n5413, ZN => 
                           n7424);
   U11538 : OAI21_X1 port map( B1 => n23206, B2 => n22820, A => n5769, ZN => 
                           n5415);
   U11539 : NOR2_X1 port map( A1 => n13988, A2 => n13987, ZN => n13917);
   U11540 : NAND2_X1 port map( A1 => n13242, A2 => n5417, ZN => n5416);
   U11541 : INV_X1 port map( A => n13248, ZN => n5417);
   U11542 : INV_X1 port map( A => n13211, ZN => n5418);
   U11543 : OAI211_X1 port map( C1 => n25004, C2 => n24341, A => n5420, B => 
                           n25081, ZN => n5419);
   U11544 : NAND2_X1 port map( A1 => n5421, A2 => n24342, ZN => n5420);
   U11545 : INV_X1 port map( A => n22932, ZN => n5421);
   U11546 : NAND2_X1 port map( A1 => n22931, A2 => n22499, ZN => n5422);
   U11547 : NAND2_X1 port map( A1 => n343, A2 => n20499, ZN => n5423);
   U11548 : NAND2_X1 port map( A1 => n16572, A2 => n5429, ZN => n5428);
   U11550 : NAND2_X1 port map( A1 => n16303, A2 => n24506, ZN => n16305);
   U11552 : XNOR2_X1 port map( A => n24568, B => n5433, ZN => n16784);
   U11553 : INV_X1 port map( A => n17065, ZN => n5434);
   U11554 : NAND2_X1 port map( A1 => n5436, A2 => n13347, ZN => n12973);
   U11555 : NAND2_X1 port map( A1 => n1328, A2 => n5437, ZN => n23586);
   U11556 : NAND3_X1 port map( A1 => n1328, A2 => n23592, A3 => n22633, ZN => 
                           n21777);
   U11558 : AND2_X1 port map( A1 => n19255, A2 => n19596, ZN => n5439);
   U11559 : INV_X1 port map( A => n14317, ZN => n5440);
   U11560 : NOR2_X1 port map( A1 => n13601, A2 => n13600, ZN => n13604);
   U11561 : NAND2_X1 port map( A1 => n18724, A2 => n19367, ZN => n19222);
   U11562 : NOR2_X1 port map( A1 => n24366, A2 => n5447, ZN => n5446);
   U11563 : INV_X1 port map( A => n16268, ZN => n5447);
   U11564 : INV_X1 port map( A => n9296, ZN => n5448);
   U11566 : XNOR2_X1 port map( A => n12073, B => n12005, ZN => n10421);
   U11570 : NAND3_X1 port map( A1 => n5454, A2 => n25474, A3 => n240, ZN => 
                           n5456);
   U11572 : XNOR2_X1 port map( A => n5457, B => n21139, ZN => n21140);
   U11573 : XNOR2_X1 port map( A => n1461, B => n21664, ZN => n5457);
   U11574 : XNOR2_X1 port map( A => n24305, B => n21138, ZN => n21664);
   U11576 : NAND3_X1 port map( A1 => n5460, A2 => n7924, A3 => n7923, ZN => 
                           n7373);
   U11577 : NAND2_X1 port map( A1 => n5461, A2 => n24424, ZN => n19100);
   U11578 : AND2_X1 port map( A1 => n25382, A2 => n22901, ZN => n22482);
   U11579 : NOR2_X1 port map( A1 => n5463, A2 => n22907, ZN => n22908);
   U11580 : NAND2_X1 port map( A1 => n22921, A2 => n5465, ZN => n23008);
   U11582 : AOI21_X1 port map( B1 => n19121, B2 => n20054, A => n25089, ZN => 
                           n5467);
   U11583 : OAI22_X1 port map( A1 => n5469, A2 => n13628, B1 => n14079, B2 => 
                           n14083, ZN => n12705);
   U11584 : MUX2_X1 port map( A => n14077, B => n13852, S => n14075, Z => n5469
                           );
   U11585 : NAND2_X1 port map( A1 => n5476, A2 => n5474, ZN => n20259);
   U11586 : NAND2_X1 port map( A1 => n5477, A2 => n19531, ZN => n5476);
   U11588 : NAND2_X1 port map( A1 => n19530, A2 => n19145, ZN => n5478);
   U11590 : OR2_X1 port map( A1 => n19531, A2 => n19534, ZN => n5481);
   U11591 : NAND2_X1 port map( A1 => n5487, A2 => n5484, ZN => n5482);
   U11592 : NAND2_X1 port map( A1 => n14397, A2 => n5484, ZN => n5483);
   U11594 : NAND2_X1 port map( A1 => n5486, A2 => n2215, ZN => n5485);
   U11595 : INV_X1 port map( A => n14397, ZN => n5486);
   U11596 : OAI22_X1 port map( A1 => n10178, A2 => n9832, B1 => n10175, B2 => 
                           n10177, ZN => n9385);
   U11597 : NAND2_X1 port map( A1 => n6600, A2 => n7019, ZN => n5488);
   U11598 : XNOR2_X1 port map( A => n21208, B => n21209, ZN => n21210);
   U11602 : OAI21_X1 port map( B1 => n19521, B2 => n19523, A => n5496, ZN => 
                           n18894);
   U11603 : XNOR2_X2 port map( A => n18194, B => n18193, ZN => n19523);
   U11605 : INV_X1 port map( A => n13924, ZN => n5497);
   U11606 : NOR2_X1 port map( A1 => n14250, A2 => n13924, ZN => n5498);
   U11607 : MUX2_X1 port map( A => n14008, B => n14254, S => n13924, Z => 
                           n14012);
   U11608 : NAND3_X1 port map( A1 => n15655, A2 => n16381, A3 => n15656, ZN => 
                           n5502);
   U11609 : NOR2_X1 port map( A1 => n20054, A2 => n20055, ZN => n20471);
   U11610 : OAI21_X1 port map( B1 => n13336, B2 => n12958, A => n5505, ZN => 
                           n13342);
   U11611 : AND2_X1 port map( A1 => n23670, A2 => n5506, ZN => n23668);
   U11612 : OR3_X1 port map( A1 => n23667, A2 => n5508, A3 => n23679, ZN => 
                           n5507);
   U11613 : NOR2_X1 port map( A1 => n22157, A2 => n25018, ZN => n5508);
   U11614 : INV_X1 port map( A => n7798, ZN => n7167);
   U11615 : NAND3_X1 port map( A1 => n7432, A2 => n7167, A3 => n7166, ZN => 
                           n7168);
   U11616 : OAI211_X1 port map( C1 => n17214, C2 => n17216, A => n17212, B => 
                           n5510, ZN => n5509);
   U11618 : AOI21_X1 port map( B1 => n12694, B2 => n13289, A => n12824, ZN => 
                           n11804);
   U11619 : NAND2_X1 port map( A1 => n5533, A2 => n10060, ZN => n5519);
   U11620 : INV_X1 port map( A => n10060, ZN => n5518);
   U11621 : OAI21_X2 port map( B1 => n13727, B2 => n5520, A => n13726, ZN => 
                           n15074);
   U11622 : NAND2_X1 port map( A1 => n16766, A2 => n5522, ZN => n5521);
   U11623 : NAND3_X1 port map( A1 => n9897, A2 => n24083, A3 => n5524, ZN => 
                           n8138);
   U11624 : OR2_X1 port map( A1 => n9944, A2 => n9899, ZN => n5523);
   U11625 : NAND2_X1 port map( A1 => n9896, A2 => n5524, ZN => n9902);
   U11626 : INV_X1 port map( A => n9899, ZN => n5524);
   U11627 : NAND2_X1 port map( A1 => n24995, A2 => n13569, ZN => n5525);
   U11628 : NAND2_X1 port map( A1 => n6255, A2 => n5903, ZN => n6953);
   U11629 : NOR2_X1 port map( A1 => n25550, A2 => n23275, ZN => n5531);
   U11630 : NAND2_X1 port map( A1 => n5531, A2 => n24907, ZN => n5530);
   U11632 : NAND2_X1 port map( A1 => n309, A2 => n9218, ZN => n5533);
   U11633 : OAI21_X1 port map( B1 => n10062, B2 => n5533, A => n9220, ZN => 
                           n9128);
   U11634 : MUX2_X1 port map( A => n5533, B => n9414, S => n10060, Z => n9415);
   U11635 : NAND2_X1 port map( A1 => n9519, A2 => n5536, ZN => n5535);
   U11636 : NAND2_X1 port map( A1 => n5537, A2 => n10176, ZN => n5536);
   U11637 : NAND2_X1 port map( A1 => n10186, A2 => n10179, ZN => n5537);
   U11638 : AOI21_X1 port map( B1 => n13210, B2 => n13212, A => n13213, ZN => 
                           n5538);
   U11639 : NAND2_X1 port map( A1 => n23165, A2 => n23181, ZN => n22552);
   U11640 : NAND2_X1 port map( A1 => n22336, A2 => n24415, ZN => n5539);
   U11642 : NAND2_X1 port map( A1 => n20156, A2 => n24558, ZN => n5541);
   U11643 : OAI21_X1 port map( B1 => n12433, B2 => n13140, A => n5542, ZN => 
                           n5545);
   U11644 : NAND2_X1 port map( A1 => n11109, A2 => n12455, ZN => n5542);
   U11645 : INV_X1 port map( A => n12455, ZN => n12729);
   U11646 : INV_X1 port map( A => n11109, ZN => n13139);
   U11647 : NAND2_X1 port map( A1 => n5545, A2 => n13143, ZN => n5544);
   U11648 : NAND2_X1 port map( A1 => n15720, A2 => n5546, ZN => n15721);
   U11649 : XNOR2_X1 port map( A => n8506, B => n9011, ZN => n8250);
   U11650 : NAND2_X1 port map( A1 => n5550, A2 => n7591, ZN => n5547);
   U11651 : NOR2_X1 port map( A1 => n5549, A2 => n5972, ZN => n5548);
   U11652 : NAND2_X1 port map( A1 => n5552, A2 => n5551, ZN => n5550);
   U11653 : NAND2_X1 port map( A1 => n5971, A2 => n7592, ZN => n5551);
   U11654 : XNOR2_X1 port map( A => n5553, B => n8739, ZN => n8489);
   U11655 : XNOR2_X1 port map( A => n5554, B => n8739, ZN => n9062);
   U11656 : INV_X1 port map( A => n9146, ZN => n5554);
   U11657 : XNOR2_X1 port map( A => n18326, B => n18214, ZN => n18576);
   U11659 : NAND2_X1 port map( A1 => n16513, A2 => n16708, ZN => n5557);
   U11660 : XNOR2_X1 port map( A => n12214, B => n12324, ZN => n11088);
   U11661 : NAND2_X1 port map( A1 => n11083, A2 => n5559, ZN => n5558);
   U11662 : OAI21_X1 port map( B1 => n6949, B2 => n25437, A => n24994, ZN => 
                           n5560);
   U11663 : NAND2_X1 port map( A1 => n5561, A2 => n12535, ZN => n13757);
   U11664 : NAND2_X1 port map( A1 => n20507, A2 => n25224, ZN => n20511);
   U11666 : OAI211_X1 port map( C1 => n3554, C2 => n15557, A => n16312, B => 
                           n15556, ZN => n16641);
   U11667 : NAND2_X1 port map( A1 => n20017, A2 => n25242, ZN => n5564);
   U11668 : NAND2_X1 port map( A1 => n5570, A2 => n5568, ZN => n20256);
   U11669 : INV_X1 port map( A => n6721, ZN => n5576);
   U11670 : NAND2_X1 port map( A1 => n6727, A2 => n6723, ZN => n5575);
   U11671 : NAND2_X1 port map( A1 => n5575, A2 => n5576, ZN => n5574);
   U11673 : INV_X1 port map( A => n12233, ZN => n5577);
   U11674 : INV_X1 port map( A => n12089, ZN => n5578);
   U11675 : XNOR2_X1 port map( A => n11907, B => n5577, ZN => n12236);
   U11676 : XNOR2_X1 port map( A => n5578, B => n11907, ZN => n12091);
   U11677 : XNOR2_X1 port map( A => n11907, B => n24514, ZN => n11911);
   U11679 : OAI211_X1 port map( C1 => n15958, C2 => n707, A => n5579, B => 
                           n15825, ZN => n5581);
   U11680 : NAND2_X1 port map( A1 => n16424, A2 => n707, ZN => n5579);
   U11681 : NAND2_X1 port map( A1 => n15958, A2 => n1329, ZN => n15962);
   U11683 : NAND2_X1 port map( A1 => n5585, A2 => n22456, ZN => n5582);
   U11684 : INV_X1 port map( A => n22451, ZN => n5585);
   U11686 : NAND2_X1 port map( A1 => n18908, A2 => n19565, ZN => n5586);
   U11687 : NAND2_X1 port map( A1 => n5589, A2 => n13350, ZN => n5588);
   U11688 : NAND2_X1 port map( A1 => n12349, A2 => n13124, ZN => n5589);
   U11689 : NOR2_X1 port map( A1 => n5591, A2 => n20401, ZN => n20402);
   U11690 : NAND2_X1 port map( A1 => n20419, A2 => n5591, ZN => n19291);
   U11691 : AOI21_X1 port map( B1 => n20419, B2 => n20415, A => n25108, ZN => 
                           n19860);
   U11694 : NAND2_X1 port map( A1 => n4463, A2 => n10838, ZN => n11135);
   U11695 : XNOR2_X1 port map( A => n17817, B => n8347, ZN => n18575);
   U11696 : XNOR2_X1 port map( A => n17817, B => n5598, ZN => n18701);
   U11697 : XNOR2_X1 port map( A => n8428, B => n8690, ZN => n9124);
   U11698 : NAND3_X1 port map( A1 => n7736, A2 => n7734, A3 => n7735, ZN => 
                           n5600);
   U11699 : NAND3_X1 port map( A1 => n25151, A2 => n7736, A3 => n7731, ZN => 
                           n5601);
   U11700 : NAND2_X1 port map( A1 => n7730, A2 => n7733, ZN => n5602);
   U11701 : NAND2_X1 port map( A1 => n7165, A2 => n5603, ZN => n8428);
   U11702 : INV_X1 port map( A => n7642, ZN => n7736);
   U11703 : NOR2_X1 port map( A1 => n7924, A2 => n7923, ZN => n5605);
   U11704 : INV_X1 port map( A => n7932, ZN => n7372);
   U11705 : NAND2_X1 port map( A1 => n5613, A2 => n5612, ZN => n20374);
   U11706 : NAND2_X1 port map( A1 => n19545, A2 => n279, ZN => n5612);
   U11707 : NAND2_X1 port map( A1 => n19544, A2 => n19543, ZN => n5613);
   U11708 : XNOR2_X1 port map( A => n5614, B => n21662, ZN => n8599);
   U11709 : XNOR2_X1 port map( A => n8313, B => n5614, ZN => n7379);
   U11710 : XNOR2_X1 port map( A => n8517, B => n5614, ZN => n8519);
   U11711 : XNOR2_X1 port map( A => n8223, B => n5614, ZN => n8793);
   U11712 : XNOR2_X1 port map( A => n9008, B => n5614, ZN => n9009);
   U11713 : NAND3_X1 port map( A1 => n14315, A2 => n13460, A3 => n14311, ZN => 
                           n14312);
   U11714 : NAND2_X1 port map( A1 => n13901, A2 => n13460, ZN => n13458);
   U11715 : NAND2_X1 port map( A1 => n13904, A2 => n5615, ZN => n15103);
   U11716 : OR2_X1 port map( A1 => n13905, A2 => n13460, ZN => n5615);
   U11717 : NAND2_X1 port map( A1 => n25021, A2 => n9945, ZN => n5616);
   U11718 : INV_X1 port map( A => n9893, ZN => n9946);
   U11720 : NAND3_X1 port map( A1 => n1429, A2 => n5618, A3 => n19169, ZN => 
                           n5617);
   U11721 : INV_X1 port map( A => n19408, ZN => n19171);
   U11722 : NAND2_X1 port map( A1 => n19412, A2 => n19408, ZN => n5618);
   U11723 : XNOR2_X1 port map( A => n9092, B => n1414, ZN => n5619);
   U11724 : OR2_X1 port map( A1 => n10063, A2 => n10064, ZN => n9702);
   U11725 : MUX2_X1 port map( A => n14059, B => n14278, S => n14850, Z => n5620
                           );
   U11726 : XNOR2_X1 port map( A => n18659, B => n18334, ZN => n17092);
   U11727 : NAND2_X1 port map( A1 => n7365, A2 => n7629, ZN => n5623);
   U11728 : OAI22_X1 port map( A1 => n406, A2 => n13125, B1 => n13126, B2 => 
                           n5626, ZN => n13127);
   U11729 : OAI21_X1 port map( B1 => n10623, B2 => n10810, A => n3868, ZN => 
                           n5630);
   U11731 : INV_X1 port map( A => n19273, ZN => n5633);
   U11732 : NAND2_X1 port map( A1 => n19570, A2 => n5634, ZN => n19567);
   U11733 : OAI21_X1 port map( B1 => n1053, B2 => n19191, A => n5631, ZN => 
                           n18909);
   U11734 : NAND2_X1 port map( A1 => n5633, A2 => n19192, ZN => n5631);
   U11736 : NAND3_X1 port map( A1 => n20545, A2 => n20546, A3 => n20124, ZN => 
                           n5637);
   U11738 : XNOR2_X1 port map( A => n14858, B => n15056, ZN => n15427);
   U11739 : NAND2_X1 port map( A1 => n14140, A2 => n5641, ZN => n5640);
   U11740 : NAND3_X1 port map( A1 => n14142, A2 => n14141, A3 => n5641, ZN => 
                           n5642);
   U11741 : NAND2_X1 port map( A1 => n12933, A2 => n12934, ZN => n5643);
   U11742 : NOR2_X1 port map( A1 => n20480, A2 => n20476, ZN => n19628);
   U11743 : OAI211_X1 port map( C1 => n19413, C2 => n19173, A => n5647, B => 
                           n19170, ZN => n5646);
   U11744 : NAND2_X1 port map( A1 => n19173, A2 => n19171, ZN => n5647);
   U11745 : OAI211_X1 port map( C1 => n6909, C2 => n6918, A => n6774, B => 
                           n24037, ZN => n5649);
   U11746 : OR2_X1 port map( A1 => n6773, A2 => n6770, ZN => n5651);
   U11747 : NAND2_X1 port map( A1 => n5650, A2 => n5649, ZN => n7974);
   U11748 : NOR2_X1 port map( A1 => n24393, A2 => n19531, ZN => n5655);
   U11749 : NAND4_X2 port map( A1 => n19271, A2 => n5652, A3 => n5654, A4 => 
                           n5653, ZN => n20400);
   U11750 : NAND2_X1 port map( A1 => n5655, A2 => n19269, ZN => n5653);
   U11751 : AND2_X1 port map( A1 => n5924, A2 => n6956, ZN => n5656);
   U11752 : NAND2_X1 port map( A1 => n5658, A2 => n23326, ZN => n23328);
   U11753 : NAND2_X1 port map( A1 => n5660, A2 => n5659, ZN => n5658);
   U11755 : NAND2_X1 port map( A1 => n21956, A2 => n5663, ZN => n5662);
   U11756 : INV_X1 port map( A => n22128, ZN => n5663);
   U11758 : NAND2_X1 port map( A1 => n338, A2 => n21467, ZN => n5665);
   U11759 : NAND3_X1 port map( A1 => n407, A2 => n25015, A3 => n12680, ZN => 
                           n12608);
   U11760 : MUX2_X1 port map( A => n13266, B => n13264, S => n12680, Z => 
                           n13271);
   U11761 : NAND2_X1 port map( A1 => n19414, A2 => n19413, ZN => n5669);
   U11762 : NAND3_X1 port map( A1 => n5673, A2 => n13283, A3 => n12899, ZN => 
                           n12700);
   U11763 : NAND2_X1 port map( A1 => n25191, A2 => n12897, ZN => n5673);
   U11764 : NAND3_X2 port map( A1 => n16735, A2 => n5675, A3 => n5674, ZN => 
                           n18190);
   U11765 : NAND2_X1 port map( A1 => n5676, A2 => n16730, ZN => n5675);
   U11766 : NOR2_X1 port map( A1 => n16731, A2 => n369, ZN => n5676);
   U11767 : MUX2_X1 port map( A => n23278, B => n23281, S => n24349, Z => 
                           n22537);
   U11768 : INV_X1 port map( A => n11025, ZN => n5679);
   U11769 : XNOR2_X1 port map( A => n11310, B => n12234, ZN => n11851);
   U11770 : NAND2_X1 port map( A1 => n19225, A2 => n5680, ZN => n19226);
   U11771 : NAND2_X1 port map( A1 => n20193, A2 => n20576, ZN => n5680);
   U11772 : NAND2_X1 port map( A1 => n5682, A2 => n25243, ZN => n5681);
   U11773 : NAND2_X1 port map( A1 => n5683, A2 => n7962, ZN => n7963);
   U11774 : NAND2_X1 port map( A1 => n5684, A2 => n7961, ZN => n5683);
   U11775 : NAND2_X1 port map( A1 => n18848, A2 => n19477, ZN => n5686);
   U11776 : NAND3_X1 port map( A1 => n18848, A2 => n19482, A3 => n19477, ZN => 
                           n18973);
   U11777 : INV_X1 port map( A => n9231, ZN => n9763);
   U11778 : OAI21_X1 port map( B1 => n10070, B2 => n9231, A => n5688, ZN => 
                           n9622);
   U11780 : NAND2_X1 port map( A1 => n9622, A2 => n1330, ZN => n9413);
   U11781 : XNOR2_X1 port map( A => n8616, B => n5690, ZN => n8102);
   U11782 : NAND2_X1 port map( A1 => n15937, A2 => n387, ZN => n15934);
   U11785 : OAI21_X1 port map( B1 => n5697, B2 => n6323, A => n5696, ZN => 
                           n5695);
   U11787 : NOR2_X1 port map( A1 => n25398, A2 => n943, ZN => n5697);
   U11788 : AOI21_X1 port map( B1 => n5700, B2 => n5699, A => n23528, ZN => 
                           n23534);
   U11789 : NAND3_X1 port map( A1 => n23533, A2 => n23531, A3 => n23532, ZN => 
                           n5699);
   U11790 : NAND2_X1 port map( A1 => n5701, A2 => n5702, ZN => n5700);
   U11791 : NAND2_X1 port map( A1 => n23505, A2 => n24351, ZN => n5702);
   U11794 : INV_X1 port map( A => n11761, ZN => n11913);
   U11796 : NOR2_X1 port map( A1 => n13373, A2 => n15888, ZN => n5706);
   U11797 : NAND2_X1 port map( A1 => n17413, A2 => n17225, ZN => n5707);
   U11798 : INV_X1 port map( A => n14108, ZN => n13582);
   U11799 : INV_X1 port map( A => n20471, ZN => n5710);
   U11800 : NAND2_X1 port map( A1 => n25088, A2 => n20060, ZN => n20468);
   U11801 : INV_X1 port map( A => n22770, ZN => n5712);
   U11802 : MUX2_X1 port map( A => n22370, B => n22774, S => n21856, Z => 
                           n22371);
   U11803 : OR2_X1 port map( A1 => n7434, A2 => n7800, ZN => n5713);
   U11804 : OAI21_X1 port map( B1 => n7799, B2 => n7794, A => n5715, ZN => 
                           n5714);
   U11805 : NAND2_X1 port map( A1 => n7794, A2 => n7802, ZN => n5715);
   U11806 : INV_X1 port map( A => n16100, ZN => n16085);
   U11807 : INV_X1 port map( A => n15584, ZN => n5716);
   U11808 : NAND2_X1 port map( A1 => n5716, A2 => n16101, ZN => n15582);
   U11809 : NAND2_X1 port map( A1 => n16957, A2 => n17414, ZN => n16954);
   U11812 : NAND2_X1 port map( A1 => n6638, A2 => n6848, ZN => n5719);
   U11813 : NAND2_X1 port map( A1 => n6109, A2 => n250, ZN => n5720);
   U11816 : XNOR2_X1 port map( A => n5722, B => n18509, ZN => n18165);
   U11817 : INV_X1 port map( A => n18218, ZN => n5722);
   U11818 : AOI21_X1 port map( B1 => n18782, B2 => n18783, A => n19411, ZN => 
                           n18787);
   U11819 : NAND3_X1 port map( A1 => n12759, A2 => n13030, A3 => n13024, ZN => 
                           n5723);
   U11820 : NAND2_X1 port map( A1 => n12760, A2 => n13028, ZN => n5724);
   U11823 : NAND2_X1 port map( A1 => n10190, A2 => n25230, ZN => n10857);
   U11824 : NAND2_X1 port map( A1 => n10190, A2 => n5727, ZN => n10865);
   U11825 : AND3_X1 port map( A1 => n22587, A2 => n22804, A3 => n22586, ZN => 
                           n22588);
   U11827 : OR2_X1 port map( A1 => n19313, A2 => n19312, ZN => n18842);
   U11829 : OR2_X1 port map( A1 => n20450, A2 => n20377, ZN => n19772);
   U11830 : OR2_X1 port map( A1 => n20401, A2 => n20414, ZN => n20203);
   U11831 : AND2_X1 port map( A1 => n20414, A2 => n20401, ZN => n19857);
   U11832 : XNOR2_X1 port map( A => n16960, B => n18089, ZN => n17562);
   U11834 : XNOR2_X1 port map( A => n20639, B => n20638, ZN => n22139);
   U11835 : OAI21_X1 port map( B1 => n21413, B2 => n22932, A => n24309, ZN => 
                           n21428);
   U11836 : INV_X1 port map( A => n19560, ZN => n19141);
   U11837 : INV_X1 port map( A => n23305, ZN => n22762);
   U11839 : NOR2_X1 port map( A1 => n19238, A2 => n25086, ZN => n18546);
   U11840 : AND2_X1 port map( A1 => n22027, A2 => n24932, ZN => n22934);
   U11843 : AND2_X1 port map( A1 => n14327, A2 => n14325, ZN => n13525);
   U11844 : OR2_X1 port map( A1 => n21806, A2 => n23779, ZN => n21807);
   U11845 : OR2_X1 port map( A1 => n21467, A2 => n22968, ZN => n21486);
   U11849 : AND2_X1 port map( A1 => n23958, A2 => n22826, ZN => n22827);
   U11850 : AND2_X1 port map( A1 => n22940, A2 => n22938, ZN => n22831);
   U11852 : OAI211_X1 port map( C1 => n22675, C2 => n22674, A => n22673, B => 
                           n22672, ZN => n23958);
   U11854 : AND2_X1 port map( A1 => n25479, A2 => n25070, ZN => n22190);
   U11855 : OR2_X1 port map( A1 => n7541, A2 => n7757, ZN => n7546);
   U11856 : AND2_X1 port map( A1 => n22983, A2 => n23860, ZN => n22984);
   U11857 : MUX2_X2 port map( A => n18760, B => n18759, S => n19265, Z => 
                           n20343);
   U11858 : INV_X1 port map( A => n11955, ZN => n11400);
   U11859 : NOR2_X1 port map( A1 => n13828, A2 => n14116, ZN => n13833);
   U11860 : INV_X1 port map( A => n23612, ZN => n23648);
   U11861 : OAI21_X1 port map( B1 => n12874, B2 => n13352, A => n12330, ZN => 
                           n13354);
   U11862 : XNOR2_X1 port map( A => n18471, B => n18470, ZN => n19578);
   U11863 : INV_X1 port map( A => n23361, ZN => n23362);
   U11864 : OAI211_X1 port map( C1 => n24941, C2 => n24059, A => n23123, B => 
                           n23091, ZN => n23096);
   U11865 : INV_X1 port map( A => n17572, ZN => n17371);
   U11866 : XNOR2_X1 port map( A => n7063, B => n7062, ZN => n7183);
   U11867 : AND2_X1 port map( A1 => n18009, A2 => n19210, ZN => n19042);
   U11869 : AND2_X1 port map( A1 => n20556, A2 => n3480, ZN => n19700);
   U11870 : NOR2_X1 port map( A1 => n14318, A2 => n14317, ZN => n14323);
   U11873 : AOI21_X1 port map( B1 => n406, B2 => n13351, A => n25430, ZN => 
                           n12621);
   U11875 : XNOR2_X2 port map( A => n21991, B => n21990, ZN => n22893);
   U11876 : OR2_X1 port map( A1 => n9531, A2 => n9805, ZN => n10117);
   U11877 : OAI21_X1 port map( B1 => n19616, B2 => n18546, A => n19613, ZN => 
                           n18547);
   U11878 : XNOR2_X1 port map( A => n11786, B => n11785, ZN => n12911);
   U11879 : AOI22_X1 port map( A1 => n9360, A2 => n9950, B1 => n2876, B2 => 
                           n9270, ZN => n10192);
   U11880 : AND2_X1 port map( A1 => n19279, A2 => n19526, ZN => n19282);
   U11881 : AND2_X1 port map( A1 => n18795, A2 => n19526, ZN => n18897);
   U11882 : OR2_X1 port map( A1 => n10280, A2 => n10190, ZN => n9268);
   U11883 : OR2_X1 port map( A1 => n23157, A2 => n23129, ZN => n23133);
   U11884 : INV_X1 port map( A => n19986, ZN => n19684);
   U11885 : XNOR2_X1 port map( A => n20735, B => n21110, ZN => n22453);
   U11886 : OR2_X1 port map( A1 => n25375, A2 => n22728, ZN => n20892);
   U11887 : OR2_X1 port map( A1 => n9462, A2 => n9461, ZN => n9464);
   U11890 : OR2_X1 port map( A1 => n13358, A2 => n12976, ZN => n12584);
   U11891 : XNOR2_X2 port map( A => n18339, B => n18338, ZN => n19192);
   U11892 : NOR2_X2 port map( A1 => n14197, A2 => n14196, ZN => n15282);
   U11893 : MUX2_X2 port map( A => n10581, B => n10580, S => n10922, Z => 
                           n12129);
   U11894 : NOR2_X1 port map( A1 => n13272, A2 => n13275, ZN => n12835);
   U11895 : OAI21_X2 port map( B1 => n22716, B2 => n22715, A => n22714, ZN => 
                           n23479);
   U11896 : MUX2_X2 port map( A => n13362, B => n13361, S => n13364, Z => 
                           n13683);
   U11898 : OR2_X1 port map( A1 => n22842, A2 => n22847, ZN => n21692);
   U11899 : OR2_X1 port map( A1 => n24475, A2 => n7657, ZN => n7660);
   U11900 : OR2_X1 port map( A1 => n23720, A2 => n23714, ZN => n22147);
   U11901 : OR2_X1 port map( A1 => n20289, A2 => n20131, ZN => n5728);
   U11902 : AND2_X1 port map( A1 => n6621, A2 => n6619, ZN => n5729);
   U11903 : AND2_X1 port map( A1 => n10489, A2 => n10613, ZN => n5730);
   U11904 : AND2_X1 port map( A1 => n13347, A2 => n13348, ZN => n5731);
   U11905 : OR3_X1 port map( A1 => n23805, A2 => n21837, A3 => n24895, ZN => 
                           n5732);
   U11906 : OR2_X1 port map( A1 => n20062, A2 => n20055, ZN => n5734);
   U11907 : AND2_X1 port map( A1 => n11057, A2 => n11009, ZN => n5735);
   U11908 : AND2_X1 port map( A1 => n18933, A2 => n19327, ZN => n5736);
   U11909 : OR2_X1 port map( A1 => n7464, A2 => n7590, ZN => n5737);
   U11910 : AND2_X1 port map( A1 => n7278, A2 => n8021, ZN => n5738);
   U11911 : INV_X1 port map( A => n9991, ZN => n9657);
   U11912 : OR2_X1 port map( A1 => n10127, A2 => n10132, ZN => n5740);
   U11913 : OR3_X1 port map( A1 => n9837, A2 => n10094, A3 => n10098, ZN => 
                           n5741);
   U11914 : AND2_X1 port map( A1 => n9820, A2 => n25463, ZN => n5742);
   U11915 : XOR2_X1 port map( A => n9061, B => n9060, Z => n5743);
   U11916 : INV_X1 port map( A => n11069, ZN => n10347);
   U11917 : XOR2_X1 port map( A => n11838, B => n1835, Z => n5745);
   U11918 : AND2_X1 port map( A1 => n10364, A2 => n10682, ZN => n5746);
   U11919 : OR2_X1 port map( A1 => n13228, A2 => n12995, ZN => n5747);
   U11920 : OR2_X1 port map( A1 => n12794, A2 => n12792, ZN => n5748);
   U11921 : INV_X1 port map( A => n12800, ZN => n11580);
   U11922 : OR2_X1 port map( A1 => n14326, A2 => n5230, ZN => n5750);
   U11923 : NOR2_X1 port map( A1 => n14127, A2 => n1331, ZN => n5751);
   U11924 : AND2_X1 port map( A1 => n14439, A2 => n13974, ZN => n5752);
   U11925 : INV_X1 port map( A => n14439, ZN => n14440);
   U11926 : AND4_X1 port map( A1 => n13666, A2 => n13665, A3 => n14000, A4 => 
                           n13664, ZN => n5753);
   U11927 : AND2_X1 port map( A1 => n25033, A2 => n13132, ZN => n5754);
   U11928 : OR2_X1 port map( A1 => n13796, A2 => n13795, ZN => n5755);
   U11929 : OR2_X1 port map( A1 => n16067, A2 => n16060, ZN => n5756);
   U11930 : XOR2_X1 port map( A => n15499, B => n13405, Z => n5757);
   U11931 : AND2_X1 port map( A1 => n15977, A2 => n16394, ZN => n5758);
   U11932 : OR2_X1 port map( A1 => n17368, A2 => n17572, ZN => n5759);
   U11933 : AND2_X1 port map( A1 => n17069, A2 => n17067, ZN => n5761);
   U11934 : XNOR2_X1 port map( A => n17999, B => n17998, ZN => n19041);
   U11935 : OR2_X1 port map( A1 => n21370, A2 => n22615, ZN => n5765);
   U11936 : AND2_X1 port map( A1 => n22837, A2 => n22836, ZN => n5766);
   U11937 : AND2_X1 port map( A1 => n22333, A2 => n22137, ZN => n5767);
   U11939 : AND2_X1 port map( A1 => n21816, A2 => n22688, ZN => n5770);
   U11940 : OR3_X1 port map( A1 => n22939, A2 => n22832, A3 => n22027, ZN => 
                           n5771);
   U11941 : OR2_X1 port map( A1 => n23394, A2 => n24449, ZN => n5772);
   U11942 : AND2_X1 port map( A1 => n24954, A2 => n24011, ZN => n5773);
   U11943 : OR2_X1 port map( A1 => n24067, A2 => n4199, ZN => n6261);
   U11944 : OR2_X1 port map( A1 => n6919, A2 => n6915, ZN => n5846);
   U11945 : INV_X1 port map( A => n6812, ZN => n6371);
   U11946 : BUF_X1 port map( A => n6392, Z => n6730);
   U11947 : OR2_X1 port map( A1 => n6334, A2 => n6209, ZN => n5949);
   U11948 : OAI22_X1 port map( A1 => n6946, A2 => n6253, B1 => n5903, B2 => 
                           n5904, ZN => n6526);
   U11949 : OR2_X1 port map( A1 => n5863, A2 => n6531, ZN => n6012);
   U11950 : OR2_X1 port map( A1 => n6817, A2 => n6893, ZN => n5830);
   U11951 : NOR2_X1 port map( A1 => n6445, A2 => n6195, ZN => n6344);
   U11952 : BUF_X1 port map( A => n6184, Z => n6457);
   U11953 : OR2_X1 port map( A1 => n7031, A2 => n7035, ZN => n6227);
   U11954 : OR2_X1 port map( A1 => n8514, A2 => n17960, ZN => n8212);
   U11955 : BUF_X1 port map( A => n6497, Z => n6503);
   U11956 : BUF_X1 port map( A => n6280, Z => n7802);
   U11960 : AND2_X1 port map( A1 => n6852, A2 => n6853, ZN => n6854);
   U11961 : OR2_X1 port map( A1 => n7821, A2 => n7820, ZN => n7822);
   U11962 : INV_X1 port map( A => n8596, ZN => n8597);
   U11963 : OR2_X1 port map( A1 => n7345, A2 => n7256, ZN => n7260);
   U11964 : INV_X1 port map( A => n8786, ZN => n8552);
   U11966 : INV_X1 port map( A => n9711, ZN => n9713);
   U11967 : OR2_X1 port map( A1 => n24222, A2 => n10104, ZN => n10106);
   U11968 : OR2_X1 port map( A1 => n8534, A2 => n7667, ZN => n7668);
   U11969 : XNOR2_X1 port map( A => n7706, B => n7705, ZN => n9345);
   U11970 : XNOR2_X1 port map( A => n8300, B => n8299, ZN => n8327);
   U11971 : AND2_X1 port map( A1 => n9285, A2 => n9898, ZN => n9288);
   U11972 : XNOR2_X1 port map( A => n8992, B => n8993, ZN => n9696);
   U11974 : AND2_X1 port map( A1 => n9945, A2 => n9899, ZN => n9445);
   U11976 : OR2_X1 port map( A1 => n9934, A2 => n9599, ZN => n9205);
   U11978 : INV_X1 port map( A => n9972, ZN => n9975);
   U11980 : XNOR2_X1 port map( A => n8267, B => n8266, ZN => n8523);
   U11981 : OR2_X1 port map( A1 => n9458, A2 => n9916, ZN => n9275);
   U11982 : OR2_X1 port map( A1 => n2953, A2 => n8142, ZN => n8143);
   U11983 : OR2_X1 port map( A1 => n10176, A2 => n10177, ZN => n9830);
   U11984 : AND2_X1 port map( A1 => n11298, A2 => n11297, ZN => n11299);
   U11985 : BUF_X1 port map( A => n9462, Z => n9920);
   U11986 : INV_X1 port map( A => n10836, ZN => n9279);
   U11987 : OR2_X1 port map( A1 => n10163, A2 => n24984, ZN => n9593);
   U11988 : OR2_X1 port map( A1 => n9864, A2 => n9860, ZN => n9556);
   U11989 : INV_X1 port map( A => n9762, ZN => n10072);
   U11990 : INV_X1 port map( A => n11143, ZN => n11885);
   U11991 : INV_X1 port map( A => n9955, ZN => n9959);
   U11992 : AND2_X1 port map( A1 => n2244, A2 => n11122, ZN => n11126);
   U11993 : INV_X1 port map( A => n10444, ZN => n10749);
   U11994 : AND2_X1 port map( A1 => n10969, A2 => n10967, ZN => n9903);
   U11995 : INV_X1 port map( A => n10590, ZN => n10372);
   U11996 : INV_X1 port map( A => n10405, ZN => n10927);
   U11997 : OR2_X1 port map( A1 => n11092, A2 => n11297, ZN => n10895);
   U11998 : AND2_X1 port map( A1 => n11059, A2 => n5735, ZN => n10978);
   U11999 : NAND4_X1 port map( A1 => n10965, A2 => n10964, A3 => n10963, A4 => 
                           n10962, ZN => n12101);
   U12000 : OR2_X1 port map( A1 => n10243, A2 => n10800, ZN => n10249);
   U12002 : OAI21_X1 port map( B1 => n11306, B2 => n11305, A => n11304, ZN => 
                           n11308);
   U12003 : INV_X1 port map( A => n13207, ZN => n11360);
   U12004 : XNOR2_X1 port map( A => n11839, B => n5745, ZN => n11844);
   U12006 : XNOR2_X1 port map( A => n10640, B => n10639, ZN => n12663);
   U12008 : INV_X1 port map( A => n11965, ZN => n13272);
   U12009 : AND2_X1 port map( A1 => n12462, A2 => n13077, ZN => n12709);
   U12010 : INV_X1 port map( A => n12892, ZN => n12895);
   U12011 : OR2_X1 port map( A1 => n4587, A2 => n12991, ZN => n12998);
   U12012 : XNOR2_X1 port map( A => n11780, B => n11779, ZN => n12594);
   U12013 : INV_X1 port map( A => n14362, ZN => n13088);
   U12014 : OR2_X1 port map( A1 => n13648, A2 => n13647, ZN => n13649);
   U12015 : INV_X1 port map( A => n14000, ZN => n13487);
   U12017 : INV_X1 port map( A => n13236, ZN => n13237);
   U12018 : OR2_X1 port map( A1 => n13990, A2 => n13989, ZN => n13991);
   U12019 : INV_X1 port map( A => n14153, ZN => n13805);
   U12020 : OR2_X1 port map( A1 => n13829, A2 => n13830, ZN => n13401);
   U12022 : AND2_X1 port map( A1 => n13997, A2 => n13995, ZN => n14232);
   U12023 : INV_X1 port map( A => n2847, ZN => n14879);
   U12026 : INV_X1 port map( A => n14880, ZN => n15417);
   U12027 : OR2_X1 port map( A1 => n13573, A2 => n13089, ZN => n13091);
   U12029 : INV_X1 port map( A => n15454, ZN => n15069);
   U12030 : XNOR2_X1 port map( A => n14985, B => n14984, ZN => n15774);
   U12031 : XNOR2_X1 port map( A => n15529, B => n15530, ZN => n15707);
   U12032 : OR2_X1 port map( A1 => n16131, A2 => n15801, ZN => n15595);
   U12034 : XNOR2_X1 port map( A => n15223, B => n15002, ZN => n15331);
   U12035 : OR2_X1 port map( A1 => n16393, A2 => n16391, ZN => n15980);
   U12036 : OR2_X1 port map( A1 => n16030, A2 => n16029, ZN => n16276);
   U12037 : OR2_X1 port map( A1 => n16449, A2 => n16451, ZN => n16239);
   U12038 : OR2_X1 port map( A1 => n24366, A2 => n16266, ZN => n16005);
   U12039 : INV_X1 port map( A => n17208, ZN => n17207);
   U12040 : AND2_X1 port map( A1 => n16422, A2 => n707, ZN => n16174);
   U12041 : AOI21_X1 port map( B1 => n15541, B2 => n294, A => n15540, ZN => 
                           n15542);
   U12042 : NOR2_X1 port map( A1 => n16897, A2 => n17081, ZN => n16898);
   U12043 : OR2_X1 port map( A1 => n2636, A2 => n16241, ZN => n15711);
   U12044 : OR2_X1 port map( A1 => n17051, A2 => n17053, ZN => n17002);
   U12045 : AOI22_X1 port map( A1 => n15989, A2 => n15988, B1 => n15987, B2 => 
                           n16414, ZN => n16765);
   U12046 : NOR2_X1 port map( A1 => n16899, A2 => n16898, ZN => n16900);
   U12047 : OAI21_X1 port map( B1 => n17242, B2 => n17241, A => n15314, ZN => 
                           n16781);
   U12048 : OR2_X1 port map( A1 => n17141, A2 => n17138, ZN => n16694);
   U12049 : XNOR2_X1 port map( A => n18146, B => n17772, ZN => n17577);
   U12052 : AND2_X1 port map( A1 => n20386, A2 => n19485, ZN => n19344);
   U12053 : XNOR2_X1 port map( A => n17577, B => n17578, ZN => n17579);
   U12054 : INV_X1 port map( A => n19061, ZN => n19056);
   U12055 : XNOR2_X1 port map( A => n18362, B => n18361, ZN => n18596);
   U12056 : XNOR2_X1 port map( A => n18664, B => n18663, ZN => n18690);
   U12057 : XNOR2_X1 port map( A => n18209, B => n18208, ZN => n18210);
   U12058 : XNOR2_X1 port map( A => n18059, B => n18058, ZN => n19587);
   U12059 : XNOR2_X1 port map( A => n18504, B => n18503, ZN => n19065);
   U12062 : AND2_X1 port map( A1 => n19560, A2 => n19290, ZN => n18752);
   U12063 : XNOR2_X1 port map( A => n18464, B => n18463, ZN => n18471);
   U12064 : OR2_X1 port map( A1 => n20359, A2 => n20484, ZN => n20487);
   U12065 : NOR2_X1 port map( A1 => n24940, A2 => n20192, ZN => n19744);
   U12066 : AND2_X1 port map( A1 => n20560, A2 => n19731, ZN => n19732);
   U12067 : NOR2_X1 port map( A1 => n25012, A2 => n19065, ZN => n19612);
   U12068 : OR2_X1 port map( A1 => n19680, A2 => n19035, ZN => n19050);
   U12070 : XNOR2_X1 port map( A => n17685, B => n17684, ZN => n19353);
   U12071 : NOR2_X1 port map( A1 => n20409, A2 => n20411, ZN => n19910);
   U12072 : OR2_X1 port map( A1 => n19288, A2 => n19857, ZN => n19292);
   U12073 : OAI21_X1 port map( B1 => n19671, B2 => n24581, A => n5728, ZN => 
                           n19672);
   U12074 : OAI21_X1 port map( B1 => n20337, B2 => n19708, A => n19707, ZN => 
                           n19712);
   U12075 : OAI211_X1 port map( C1 => n18855, C2 => n18934, A => n18854, B => 
                           n18853, ZN => n19195);
   U12076 : INV_X1 port map( A => n20173, ZN => n20170);
   U12077 : INV_X1 port map( A => n20354, ZN => n20355);
   U12078 : OR2_X1 port map( A1 => n20141, A2 => n19975, ZN => n20144);
   U12079 : XNOR2_X1 port map( A => n24434, B => n21431, ZN => n21432);
   U12081 : INV_X1 port map( A => n20222, ZN => n19927);
   U12082 : INV_X1 port map( A => n22798, ZN => n22584);
   U12085 : OR2_X1 port map( A1 => n21920, A2 => n22752, ZN => n22561);
   U12086 : BUF_X1 port map( A => n21908, Z => n21910);
   U12087 : NOR2_X1 port map( A1 => n22947, A2 => n22282, ZN => n22945);
   U12089 : AND2_X1 port map( A1 => n22209, A2 => n24333, ZN => n20932);
   U12090 : AOI211_X1 port map( C1 => n22800, C2 => n24559, A => n22803, B => 
                           n22798, ZN => n22476);
   U12091 : BUF_X1 port map( A => n20776, Z => n22400);
   U12092 : AND2_X1 port map( A1 => n22952, A2 => n22954, ZN => n22857);
   U12093 : NOR2_X1 port map( A1 => n22726, A2 => n22725, ZN => n23470);
   U12094 : AND3_X1 port map( A1 => n22187, A2 => n22929, A3 => n22111, ZN => 
                           n22112);
   U12095 : OR2_X1 port map( A1 => n20940, A2 => n22066, ZN => n20941);
   U12097 : OR2_X1 port map( A1 => n22794, A2 => n24953, ZN => n22795);
   U12098 : AND2_X1 port map( A1 => n23052, A2 => n23040, ZN => n22643);
   U12102 : INV_X1 port map( A => n23499, ZN => n23484);
   U12103 : AND2_X1 port map( A1 => n23647, A2 => n20896, ZN => n20981);
   U12104 : OAI21_X1 port map( B1 => n22598, B2 => n21855, A => n21854, ZN => 
                           n23869);
   U12106 : OAI21_X1 port map( B1 => n22304, B2 => n5772, A => n22303, ZN => 
                           n22305);
   U12107 : OR2_X1 port map( A1 => n23386, A2 => n24879, ZN => n22884);
   U12109 : INV_X1 port map( A => n187, ZN => n22049);
   U12110 : XNOR2_X1 port map( A => Key(76), B => Plaintext(76), ZN => n6744);
   U12111 : XNOR2_X1 port map( A => Key(73), B => Plaintext(73), ZN => n6050);
   U12112 : XNOR2_X1 port map( A => Key(72), B => Plaintext(72), ZN => n6407);
   U12113 : NAND2_X1 port map( A1 => n6630, A2 => n6407, ZN => n5776);
   U12114 : OAI21_X1 port map( B1 => n453, B2 => n6630, A => n5776, ZN => n5777
                           );
   U12116 : INV_X1 port map( A => n6051, ZN => n6628);
   U12117 : INV_X1 port map( A => Plaintext(90), ZN => n5778);
   U12118 : XNOR2_X1 port map( A => n5778, B => Key(90), ZN => n6235);
   U12119 : INV_X1 port map( A => Plaintext(91), ZN => n5779);
   U12120 : NAND2_X1 port map( A1 => n6235, A2 => n6712, ZN => n6112);
   U12121 : INV_X1 port map( A => Plaintext(95), ZN => n5780);
   U12123 : INV_X1 port map( A => Plaintext(92), ZN => n5781);
   U12124 : XNOR2_X1 port map( A => n5781, B => Key(92), ZN => n6234);
   U12125 : INV_X1 port map( A => n6234, ZN => n6232);
   U12126 : INV_X1 port map( A => Plaintext(94), ZN => n5782);
   U12128 : INV_X1 port map( A => n6233, ZN => n6714);
   U12130 : INV_X1 port map( A => Plaintext(93), ZN => n5783);
   U12131 : NAND2_X1 port map( A1 => n24051, A2 => n6712, ZN => n5784);
   U12132 : INV_X1 port map( A => Plaintext(84), ZN => n5787);
   U12133 : XNOR2_X1 port map( A => n5787, B => Key(84), ZN => n5795);
   U12134 : INV_X1 port map( A => Plaintext(87), ZN => n5788);
   U12135 : XNOR2_X1 port map( A => n5788, B => Key(87), ZN => n5794);
   U12136 : NAND2_X1 port map( A1 => n6619, A2 => n6623, ZN => n5793);
   U12137 : INV_X1 port map( A => Plaintext(88), ZN => n5789);
   U12138 : INV_X1 port map( A => Plaintext(86), ZN => n5790);
   U12139 : NAND2_X1 port map( A1 => n6622, A2 => n6049, ZN => n5792);
   U12140 : INV_X1 port map( A => Plaintext(89), ZN => n5791);
   U12141 : INV_X1 port map( A => n6114, ZN => n6723);
   U12142 : MUX2_X1 port map( A => n5793, B => n5792, S => n6723, Z => n5799);
   U12143 : INV_X1 port map( A => n5795, ZN => n6724);
   U12144 : MUX2_X1 port map( A => n6722, B => n6243, S => n6724, Z => n5797);
   U12145 : NAND2_X1 port map( A1 => n5797, A2 => n5796, ZN => n5798);
   U12149 : OAI21_X1 port map( B1 => n443, B2 => n6963, A => n5800, ZN => n5802
                           );
   U12151 : NAND2_X1 port map( A1 => n6965, A2 => n6964, ZN => n5801);
   U12152 : XNOR2_X1 port map( A => Key(69), B => Plaintext(69), ZN => n6577);
   U12153 : INV_X1 port map( A => Plaintext(67), ZN => n5803);
   U12154 : NAND2_X1 port map( A1 => n6752, A2 => n271, ZN => n6754);
   U12155 : XNOR2_X1 port map( A => Key(70), B => Plaintext(70), ZN => n6757);
   U12156 : AND2_X1 port map( A1 => n6757, A2 => n6578, ZN => n5808);
   U12157 : XNOR2_X1 port map( A => Key(66), B => Plaintext(66), ZN => n6751);
   U12159 : NAND3_X1 port map( A1 => n6675, A2 => n5804, A3 => n6578, ZN => 
                           n5807);
   U12160 : XNOR2_X1 port map( A => Key(68), B => Plaintext(68), ZN => n6400);
   U12161 : NAND2_X1 port map( A1 => n5805, A2 => n6755, ZN => n5806);
   U12162 : NAND2_X1 port map( A1 => n7576, A2 => n7579, ZN => n5809);
   U12163 : XNOR2_X1 port map( A => Key(83), B => Plaintext(83), ZN => n6060);
   U12164 : INV_X1 port map( A => n6060, ZN => n6393);
   U12165 : INV_X1 port map( A => Plaintext(81), ZN => n5810);
   U12166 : XNOR2_X1 port map( A => n5810, B => Key(81), ZN => n6062);
   U12167 : INV_X1 port map( A => n6062, ZN => n6729);
   U12169 : NAND2_X1 port map( A1 => n6729, A2 => n6396, ZN => n6736);
   U12171 : XNOR2_X1 port map( A => Key(80), B => Plaintext(80), ZN => n6392);
   U12172 : NAND2_X1 port map( A1 => n6732, A2 => n6392, ZN => n5812);
   U12173 : NAND2_X1 port map( A1 => n5812, A2 => n6393, ZN => n5811);
   U12174 : OAI21_X1 port map( B1 => n6393, B2 => n6736, A => n5811, ZN => 
                           n5814);
   U12175 : INV_X1 port map( A => n6392, ZN => n6615);
   U12176 : XNOR2_X1 port map( A => Key(82), B => Plaintext(82), ZN => n6238);
   U12177 : NAND3_X1 port map( A1 => n6393, A2 => n6615, A3 => n6238, ZN => 
                           n6242);
   U12178 : NOR2_X1 port map( A1 => n5812, A2 => n2119, ZN => n5813);
   U12179 : OR2_X1 port map( A1 => n7577, A2 => n7576, ZN => n7483);
   U12180 : MUX2_X1 port map( A => n4136, B => n5815, S => n7483, Z => n5816);
   U12181 : XNOR2_X1 port map( A => Key(131), B => Plaintext(131), ZN => n6071)
                           ;
   U12182 : INV_X1 port map( A => n6071, ZN => n6815);
   U12183 : XNOR2_X1 port map( A => Key(130), B => Plaintext(130), ZN => n6369)
                           ;
   U12184 : INV_X1 port map( A => n6369, ZN => n6999);
   U12185 : INV_X1 port map( A => Plaintext(126), ZN => n5817);
   U12186 : XNOR2_X1 port map( A => Key(129), B => Plaintext(129), ZN => n6368)
                           ;
   U12187 : AOI21_X1 port map( B1 => n7003, B2 => n439, A => n6997, ZN => n5821
                           );
   U12189 : XNOR2_X1 port map( A => Key(127), B => Plaintext(127), ZN => n6996)
                           ;
   U12190 : AOI21_X1 port map( B1 => n5819, B2 => n5818, A => n6999, ZN => 
                           n5820);
   U12191 : INV_X1 port map( A => Plaintext(146), ZN => n5822);
   U12192 : INV_X1 port map( A => Plaintext(149), ZN => n5823);
   U12193 : XNOR2_X1 port map( A => n5823, B => Key(149), ZN => n6375);
   U12194 : NAND2_X1 port map( A1 => n6377, A2 => n6375, ZN => n6789);
   U12195 : XNOR2_X1 port map( A => Key(147), B => Plaintext(147), ZN => n6473)
                           ;
   U12196 : INV_X1 port map( A => n6377, ZN => n6374);
   U12197 : NAND3_X1 port map( A1 => n6473, A2 => n6373, A3 => n6906, ZN => 
                           n5825);
   U12198 : INV_X1 port map( A => n7887, ZN => n5861);
   U12199 : XNOR2_X1 port map( A => Key(132), B => Plaintext(132), ZN => n6890)
                           ;
   U12200 : INV_X1 port map( A => n6890, ZN => n6819);
   U12201 : XNOR2_X1 port map( A => Key(133), B => Plaintext(133), ZN => n6086)
                           ;
   U12202 : INV_X1 port map( A => n6086, ZN => n6818);
   U12203 : NAND2_X1 port map( A1 => n6819, A2 => n6818, ZN => n6817);
   U12204 : INV_X1 port map( A => Plaintext(137), ZN => n5826);
   U12205 : INV_X1 port map( A => Plaintext(136), ZN => n5827);
   U12206 : XNOR2_X1 port map( A => n5827, B => Key(136), ZN => n6651);
   U12207 : INV_X1 port map( A => Plaintext(135), ZN => n5828);
   U12208 : XNOR2_X2 port map( A => n5828, B => Key(135), ZN => n6895);
   U12209 : INV_X1 port map( A => Plaintext(134), ZN => n5829);
   U12211 : INV_X1 port map( A => n6076, ZN => n6882);
   U12212 : INV_X1 port map( A => Plaintext(142), ZN => n5831);
   U12213 : INV_X1 port map( A => n6795, ZN => n6884);
   U12214 : XNOR2_X1 port map( A => Key(143), B => Plaintext(143), ZN => n5833)
                           ;
   U12215 : BUF_X2 port map( A => n5833, Z => n6885);
   U12216 : INV_X1 port map( A => n5833, ZN => n6881);
   U12217 : INV_X1 port map( A => Plaintext(141), ZN => n5834);
   U12218 : XNOR2_X1 port map( A => n5834, B => Key(141), ZN => n5835);
   U12219 : NAND3_X1 port map( A1 => n6881, A2 => n6793, A3 => n6794, ZN => 
                           n5838);
   U12220 : INV_X1 port map( A => n5835, ZN => n6075);
   U12221 : INV_X1 port map( A => Key(140), ZN => n23151);
   U12222 : INV_X1 port map( A => Plaintext(140), ZN => n5836);
   U12223 : NAND4_X1 port map( A1 => n6075, A2 => n6885, A3 => n23151, A4 => 
                           n5836, ZN => n5837);
   U12224 : AND2_X1 port map( A1 => n5837, A2 => n5838, ZN => n5843);
   U12225 : INV_X1 port map( A => Plaintext(138), ZN => n5839);
   U12226 : NAND3_X1 port map( A1 => n5833, A2 => Key(140), A3 => 
                           Plaintext(140), ZN => n5840);
   U12227 : OAI21_X1 port map( B1 => n6078, B2 => n6885, A => n5840, ZN => 
                           n5841);
   U12228 : NAND2_X1 port map( A1 => n5841, A2 => n6075, ZN => n5842);
   U12229 : OAI21_X1 port map( B1 => n7879, B2 => n7585, A => n7313, ZN => 
                           n5860);
   U12230 : INV_X1 port map( A => Plaintext(160), ZN => n5844);
   U12231 : XNOR2_X1 port map( A => Key(156), B => Plaintext(156), ZN => n6917)
                           ;
   U12232 : INV_X1 port map( A => n6917, ZN => n6916);
   U12233 : AOI21_X1 port map( B1 => n5846, B2 => n5845, A => n6918, ZN => 
                           n5850);
   U12234 : INV_X1 port map( A => Plaintext(161), ZN => n5847);
   U12235 : NAND3_X1 port map( A1 => n6912, A2 => n6770, A3 => n6919, ZN => 
                           n5848);
   U12236 : OAI21_X1 port map( B1 => n6916, B2 => n24037, A => n5848, ZN => 
                           n5849);
   U12237 : INV_X1 port map( A => Plaintext(154), ZN => n5851);
   U12238 : XNOR2_X1 port map( A => Key(155), B => Plaintext(155), ZN => n6081)
                           ;
   U12239 : NAND2_X1 port map( A1 => n6767, A2 => n6876, ZN => n5855);
   U12240 : INV_X1 port map( A => Plaintext(150), ZN => n5852);
   U12241 : XNOR2_X1 port map( A => n5852, B => Key(150), ZN => n6083);
   U12242 : INV_X1 port map( A => n6083, ZN => n6875);
   U12243 : INV_X1 port map( A => Plaintext(151), ZN => n5853);
   U12244 : XNOR2_X1 port map( A => n5853, B => Key(151), ZN => n6310);
   U12245 : INV_X1 port map( A => n6310, ZN => n6870);
   U12246 : NAND2_X1 port map( A1 => n6875, A2 => n6870, ZN => n5854);
   U12247 : XNOR2_X1 port map( A => Key(152), B => Plaintext(152), ZN => n6871)
                           ;
   U12249 : NAND2_X1 port map( A1 => n5856, A2 => n6083, ZN => n5857);
   U12250 : AND2_X1 port map( A1 => n5858, A2 => n5857, ZN => n7584);
   U12252 : XNOR2_X1 port map( A => n8596, B => n8666, ZN => n8249);
   U12253 : INV_X1 port map( A => Plaintext(28), ZN => n5862);
   U12254 : INV_X1 port map( A => n6532, ZN => n5863);
   U12255 : INV_X1 port map( A => Plaintext(24), ZN => n5864);
   U12256 : XNOR2_X1 port map( A => n5864, B => Key(24), ZN => n6013);
   U12257 : INV_X1 port map( A => n6013, ZN => n6538);
   U12258 : AOI21_X1 port map( B1 => n6012, B2 => n6538, A => n6530, ZN => 
                           n5869);
   U12259 : INV_X1 port map( A => Plaintext(26), ZN => n5865);
   U12260 : INV_X1 port map( A => n6531, ZN => n6259);
   U12262 : NAND2_X1 port map( A1 => n4199, A2 => n6530, ZN => n5866);
   U12263 : AOI21_X1 port map( B1 => n5867, B2 => n5866, A => n6532, ZN => 
                           n5868);
   U12264 : INV_X1 port map( A => Plaintext(46), ZN => n5870);
   U12266 : XNOR2_X1 port map( A => Key(43), B => Plaintext(43), ZN => n6703);
   U12267 : XNOR2_X1 port map( A => Key(47), B => Plaintext(47), ZN => n6705);
   U12268 : INV_X1 port map( A => n6705, ZN => n6960);
   U12269 : INV_X1 port map( A => Plaintext(42), ZN => n5871);
   U12270 : INV_X1 port map( A => n5924, ZN => n6957);
   U12271 : XNOR2_X2 port map( A => Key(45), B => Plaintext(45), ZN => n6959);
   U12273 : XNOR2_X1 port map( A => Key(57), B => Plaintext(57), ZN => n6066);
   U12274 : INV_X1 port map( A => n6066, ZN => n6971);
   U12275 : INV_X1 port map( A => Plaintext(55), ZN => n5872);
   U12278 : INV_X1 port map( A => Plaintext(56), ZN => n5873);
   U12279 : INV_X1 port map( A => Plaintext(58), ZN => n5874);
   U12282 : NAND2_X1 port map( A1 => n6692, A2 => n6977, ZN => n5875);
   U12283 : INV_X1 port map( A => Plaintext(30), ZN => n5877);
   U12284 : INV_X1 port map( A => n6529, ZN => n6946);
   U12285 : INV_X1 port map( A => Plaintext(31), ZN => n5878);
   U12286 : XNOR2_X1 port map( A => n5878, B => Key(31), ZN => n5902);
   U12287 : INV_X1 port map( A => n5902, ZN => n6253);
   U12288 : INV_X1 port map( A => Plaintext(32), ZN => n5879);
   U12289 : INV_X1 port map( A => n5904, ZN => n6255);
   U12290 : XNOR2_X1 port map( A => Key(33), B => Plaintext(33), ZN => n6948);
   U12291 : NAND2_X1 port map( A1 => n6253, A2 => n6948, ZN => n6139);
   U12292 : INV_X1 port map( A => n6139, ZN => n5882);
   U12293 : INV_X1 port map( A => Plaintext(34), ZN => n5880);
   U12295 : AOI22_X1 port map( A1 => n6526, A2 => n6953, B1 => n5882, B2 => 
                           n5881, ZN => n7327);
   U12296 : XNOR2_X1 port map( A => Key(39), B => Plaintext(39), ZN => n5887);
   U12297 : INV_X1 port map( A => n5887, ZN => n6684);
   U12298 : XNOR2_X1 port map( A => Key(37), B => Plaintext(37), ZN => n5910);
   U12299 : INV_X1 port map( A => n5910, ZN => n6680);
   U12300 : XNOR2_X1 port map( A => Key(36), B => Plaintext(36), ZN => n6146);
   U12301 : NOR2_X1 port map( A1 => n6684, A2 => n6146, ZN => n5883);
   U12302 : XNOR2_X1 port map( A => Key(41), B => Plaintext(41), ZN => n5888);
   U12303 : INV_X1 port map( A => n5888, ZN => n6944);
   U12304 : OAI21_X1 port map( B1 => n5884, B2 => n5883, A => n6944, ZN => 
                           n5890);
   U12305 : INV_X1 port map( A => Plaintext(38), ZN => n5885);
   U12306 : XNOR2_X1 port map( A => n5885, B => Key(38), ZN => n5908);
   U12307 : INV_X1 port map( A => Plaintext(40), ZN => n5886);
   U12309 : INV_X1 port map( A => n5908, ZN => n6281);
   U12310 : INV_X1 port map( A => Plaintext(51), ZN => n5891);
   U12311 : XNOR2_X1 port map( A => n5891, B => Key(51), ZN => n6414);
   U12313 : XNOR2_X1 port map( A => Key(49), B => Plaintext(49), ZN => n6694);
   U12314 : INV_X1 port map( A => n6694, ZN => n5893);
   U12315 : INV_X1 port map( A => Plaintext(48), ZN => n5892);
   U12316 : INV_X1 port map( A => n6556, ZN => n6693);
   U12317 : MUX2_X1 port map( A => n6695, B => n5893, S => n6693, Z => n5900);
   U12318 : INV_X1 port map( A => Plaintext(50), ZN => n5894);
   U12319 : NAND2_X1 port map( A1 => n6695, A2 => n6556, ZN => n5898);
   U12320 : INV_X1 port map( A => Plaintext(52), ZN => n5895);
   U12321 : INV_X1 port map( A => Plaintext(53), ZN => n5896);
   U12322 : MUX2_X1 port map( A => n5898, B => n5897, S => n6934, Z => n5899);
   U12323 : XNOR2_X1 port map( A => n8412, B => n860, ZN => n5930);
   U12324 : INV_X1 port map( A => n5903, ZN => n6528);
   U12325 : INV_X1 port map( A => n6948, ZN => n6947);
   U12326 : NAND2_X1 port map( A1 => n5908, A2 => n6683, ZN => n5909);
   U12327 : MUX2_X1 port map( A => n7250, B => n8508, S => n8512, Z => n8209);
   U12328 : INV_X1 port map( A => Plaintext(18), ZN => n5913);
   U12329 : XNOR2_X1 port map( A => Key(21), B => Plaintext(21), ZN => n6267);
   U12330 : INV_X1 port map( A => Plaintext(19), ZN => n5914);
   U12331 : XNOR2_X1 port map( A => n5914, B => Key(19), ZN => n5915);
   U12332 : INV_X1 port map( A => n5915, ZN => n6539);
   U12333 : XNOR2_X1 port map( A => Key(23), B => Plaintext(23), ZN => n6133);
   U12334 : INV_X1 port map( A => n6267, ZN => n7103);
   U12335 : XNOR2_X1 port map( A => Key(22), B => Plaintext(22), ZN => n7101);
   U12336 : INV_X1 port map( A => n5916, ZN => n6266);
   U12338 : NAND2_X1 port map( A1 => n127, A2 => n6164, ZN => n5917);
   U12339 : NAND2_X1 port map( A1 => n6530, A2 => n6533, ZN => n5918);
   U12340 : AOI21_X1 port map( B1 => n5918, B2 => n24067, A => n6531, ZN => 
                           n5923);
   U12341 : NAND3_X1 port map( A1 => n4199, A2 => n25014, A3 => n6531, ZN => 
                           n5921);
   U12342 : NAND2_X1 port map( A1 => n5921, A2 => n5920, ZN => n5922);
   U12343 : AND2_X1 port map( A1 => n7350, A2 => n7346, ZN => n5929);
   U12344 : NAND2_X1 port map( A1 => n6956, A2 => n24405, ZN => n6137);
   U12345 : INV_X1 port map( A => n6959, ZN => n6553);
   U12346 : NAND2_X1 port map( A1 => n6553, A2 => n6705, ZN => n5925);
   U12347 : NAND2_X1 port map( A1 => n24405, A2 => n6959, ZN => n6954);
   U12348 : NAND3_X1 port map( A1 => n5925, A2 => n6954, A3 => n5924, ZN => 
                           n5927);
   U12349 : NAND3_X1 port map( A1 => n3926, A2 => n6703, A3 => n3922, ZN => 
                           n5926);
   U12350 : OAI211_X1 port map( C1 => n6137, C2 => n6960, A => n5927, B => 
                           n5926, ZN => n7348);
   U12351 : OAI21_X1 port map( B1 => n7250, B2 => n5929, A => n5928, ZN => 
                           n8514);
   U12352 : OAI21_X1 port map( B1 => n8209, B2 => n7350, A => n8514, ZN => 
                           n9175);
   U12353 : INV_X1 port map( A => n6445, ZN => n6019);
   U12354 : XNOR2_X1 port map( A => Key(186), B => Plaintext(186), ZN => n6444)
                           ;
   U12355 : INV_X1 port map( A => n6444, ZN => n6345);
   U12356 : INV_X1 port map( A => n6021, ZN => n5935);
   U12358 : INV_X1 port map( A => n6452, ZN => n6341);
   U12359 : OAI21_X1 port map( B1 => n6345, B2 => n6195, A => n6341, ZN => 
                           n5934);
   U12360 : XNOR2_X1 port map( A => Key(190), B => Plaintext(190), ZN => n6447)
                           ;
   U12361 : INV_X1 port map( A => n6447, ZN => n6196);
   U12362 : NAND2_X1 port map( A1 => n6196, A2 => n6452, ZN => n5932);
   U12363 : INV_X1 port map( A => Plaintext(191), ZN => n5931);
   U12365 : INV_X1 port map( A => n6187, ZN => n6449);
   U12366 : MUX2_X1 port map( A => n6021, B => n5932, S => n6449, Z => n5933);
   U12367 : INV_X1 port map( A => n7464, ZN => n7587);
   U12368 : INV_X1 port map( A => Plaintext(3), ZN => n5936);
   U12370 : INV_X1 port map( A => Plaintext(1), ZN => n5937);
   U12371 : AND2_X1 port map( A1 => n6513, A2 => n6456, ZN => n6183);
   U12372 : INV_X1 port map( A => n6183, ZN => n5939);
   U12373 : INV_X1 port map( A => n6455, ZN => n6454);
   U12374 : INV_X1 port map( A => Plaintext(2), ZN => n5938);
   U12375 : XNOR2_X1 port map( A => n5938, B => Key(2), ZN => n6184);
   U12376 : INV_X1 port map( A => n6184, ZN => n6509);
   U12377 : AOI21_X1 port map( B1 => n5939, B2 => n6454, A => n6509, ZN => 
                           n5942);
   U12378 : INV_X1 port map( A => Plaintext(5), ZN => n5940);
   U12379 : NAND2_X1 port map( A1 => n6509, A2 => n6510, ZN => n6030);
   U12380 : XNOR2_X1 port map( A => Key(4), B => Plaintext(4), ZN => n6512);
   U12381 : NOR2_X1 port map( A1 => n7587, A2 => n7590, ZN => n5970);
   U12382 : INV_X1 port map( A => Plaintext(182), ZN => n5943);
   U12383 : INV_X1 port map( A => Plaintext(181), ZN => n5944);
   U12385 : INV_X1 port map( A => n6297, ZN => n6209);
   U12386 : INV_X1 port map( A => Plaintext(184), ZN => n5945);
   U12387 : XNOR2_X1 port map( A => n5945, B => Key(184), ZN => n6332);
   U12388 : NAND2_X1 port map( A1 => n6335, A2 => n6332, ZN => n6173);
   U12389 : XNOR2_X1 port map( A => Key(180), B => Plaintext(180), ZN => n6208)
                           ;
   U12390 : INV_X1 port map( A => n6335, ZN => n6439);
   U12391 : XNOR2_X2 port map( A => Key(173), B => Plaintext(173), ZN => n6493)
                           ;
   U12392 : INV_X1 port map( A => Plaintext(170), ZN => n5950);
   U12394 : INV_X1 port map( A => Plaintext(171), ZN => n5951);
   U12395 : INV_X1 port map( A => n6427, ZN => n6301);
   U12396 : INV_X1 port map( A => Plaintext(169), ZN => n5952);
   U12397 : INV_X1 port map( A => n6488, ZN => n6304);
   U12398 : NAND2_X1 port map( A1 => n6781, A2 => n5953, ZN => n5956);
   U12399 : INV_X1 port map( A => Plaintext(172), ZN => n5954);
   U12401 : INV_X1 port map( A => n6490, ZN => n6780);
   U12402 : NAND2_X1 port map( A1 => n6493, A2 => n6780, ZN => n5955);
   U12403 : NAND2_X1 port map( A1 => n5956, A2 => n5955, ZN => n5960);
   U12404 : INV_X1 port map( A => Plaintext(168), ZN => n5957);
   U12405 : XNOR2_X1 port map( A => n5957, B => Key(168), ZN => n6784);
   U12406 : NAND2_X1 port map( A1 => n6784, A2 => n6488, ZN => n6782);
   U12407 : INV_X1 port map( A => n6782, ZN => n5958);
   U12408 : NAND2_X1 port map( A1 => n5958, A2 => n6493, ZN => n5959);
   U12409 : NAND2_X1 port map( A1 => n5960, A2 => n5959, ZN => n7335);
   U12410 : XNOR2_X1 port map( A => Key(162), B => Plaintext(162), ZN => n6777)
                           ;
   U12411 : INV_X1 port map( A => Plaintext(163), ZN => n5961);
   U12412 : INV_X1 port map( A => Plaintext(164), ZN => n5962);
   U12413 : INV_X1 port map( A => Plaintext(166), ZN => n5963);
   U12414 : XNOR2_X1 port map( A => n5963, B => Key(166), ZN => n6776);
   U12415 : INV_X1 port map( A => Plaintext(177), ZN => n5965);
   U12416 : INV_X1 port map( A => n5966, ZN => n6315);
   U12418 : INV_X1 port map( A => Plaintext(174), ZN => n5967);
   U12419 : XNOR2_X1 port map( A => n5967, B => Key(174), ZN => n6470);
   U12420 : INV_X1 port map( A => n6470, ZN => n6329);
   U12421 : INV_X1 port map( A => Plaintext(175), ZN => n5968);
   U12422 : NAND2_X1 port map( A1 => n4621, A2 => n6426, ZN => n6471);
   U12423 : INV_X1 port map( A => Plaintext(179), ZN => n5969);
   U12424 : NOR2_X1 port map( A1 => n7593, A2 => n5971, ZN => n5972);
   U12425 : XNOR2_X1 port map( A => Key(110), B => Plaintext(110), ZN => n6245)
                           ;
   U12426 : AND2_X1 port map( A1 => n6245, A2 => n6244, ZN => n5975);
   U12427 : XNOR2_X1 port map( A => Key(113), B => Plaintext(113), ZN => n6122)
                           ;
   U12428 : XNOR2_X1 port map( A => Key(108), B => Plaintext(108), ZN => n6119)
                           ;
   U12429 : NAND2_X1 port map( A1 => n6122, A2 => n6119, ZN => n5973);
   U12430 : NAND2_X1 port map( A1 => n5973, A2 => n6987, ZN => n5974);
   U12431 : INV_X1 port map( A => n6245, ZN => n6841);
   U12432 : XNOR2_X1 port map( A => Key(112), B => Plaintext(112), ZN => n6640)
                           ;
   U12433 : INV_X1 port map( A => n5975, ZN => n5976);
   U12434 : INV_X1 port map( A => n6122, ZN => n6986);
   U12435 : NAND3_X1 port map( A1 => n6639, A2 => n5976, A3 => n6986, ZN => 
                           n5977);
   U12436 : INV_X1 port map( A => Plaintext(121), ZN => n5979);
   U12437 : INV_X1 port map( A => Plaintext(120), ZN => n5980);
   U12438 : XNOR2_X1 port map( A => n5980, B => Key(120), ZN => n6647);
   U12439 : AND2_X1 port map( A1 => n6647, A2 => n7004, ZN => n6384);
   U12440 : XNOR2_X1 port map( A => Key(124), B => Plaintext(124), ZN => n6094)
                           ;
   U12441 : INV_X1 port map( A => n6094, ZN => n6650);
   U12442 : NAND2_X1 port map( A1 => n6384, A2 => n6650, ZN => n5985);
   U12443 : NAND3_X1 port map( A1 => n7006, A2 => n7004, A3 => n448, ZN => 
                           n5984);
   U12444 : INV_X1 port map( A => Plaintext(125), ZN => n5981);
   U12445 : AND2_X1 port map( A1 => n7007, A2 => n6648, ZN => n6836);
   U12446 : NAND2_X1 port map( A1 => n6836, A2 => n6650, ZN => n5983);
   U12447 : INV_X1 port map( A => n6647, ZN => n7009);
   U12449 : NAND3_X1 port map( A1 => n24051, A2 => n6233, A3 => n24500, ZN => 
                           n5988);
   U12450 : NAND3_X1 port map( A1 => n6234, A2 => n24501, A3 => n6714, ZN => 
                           n5987);
   U12451 : INV_X1 port map( A => n24050, ZN => n6611);
   U12452 : NAND3_X1 port map( A1 => n6712, A2 => n6611, A3 => n6714, ZN => 
                           n5986);
   U12453 : INV_X1 port map( A => n5992, ZN => n7019);
   U12454 : INV_X1 port map( A => Plaintext(102), ZN => n5989);
   U12455 : XNOR2_X1 port map( A => n5989, B => Key(102), ZN => n6598);
   U12456 : INV_X1 port map( A => Plaintext(105), ZN => n5990);
   U12457 : INV_X1 port map( A => n6823, ZN => n7015);
   U12458 : NAND3_X1 port map( A1 => n7019, A2 => n6598, A3 => n7015, ZN => 
                           n5996);
   U12459 : INV_X1 port map( A => Plaintext(104), ZN => n5991);
   U12460 : NAND2_X1 port map( A1 => n25044, A2 => n5992, ZN => n5995);
   U12461 : NAND2_X1 port map( A1 => n6823, A2 => n5992, ZN => n5994);
   U12462 : INV_X1 port map( A => Plaintext(103), ZN => n5993);
   U12463 : XNOR2_X1 port map( A => Key(106), B => Plaintext(106), ZN => n7013)
                           ;
   U12464 : NAND2_X1 port map( A1 => n6100, A2 => n6824, ZN => n5997);
   U12466 : INV_X1 port map( A => n7026, ZN => n6846);
   U12467 : XNOR2_X1 port map( A => Key(117), B => Plaintext(117), ZN => n6845)
                           ;
   U12468 : INV_X1 port map( A => n6845, ZN => n7022);
   U12469 : INV_X1 port map( A => Plaintext(119), ZN => n5999);
   U12470 : XNOR2_X1 port map( A => n5999, B => Key(119), ZN => n6381);
   U12471 : INV_X1 port map( A => Plaintext(116), ZN => n6000);
   U12473 : INV_X1 port map( A => n7021, ZN => n7024);
   U12474 : NAND2_X1 port map( A1 => n7024, A2 => n7026, ZN => n6001);
   U12475 : INV_X1 port map( A => Plaintext(118), ZN => n6002);
   U12476 : INV_X1 port map( A => n6849, ZN => n7023);
   U12477 : NAND3_X1 port map( A1 => n6848, A2 => n7023, A3 => n442, ZN => 
                           n6003);
   U12479 : XNOR2_X1 port map( A => Key(98), B => Plaintext(98), ZN => n6104);
   U12480 : INV_X1 port map( A => Plaintext(101), ZN => n6004);
   U12481 : OAI21_X1 port map( B1 => n7032, B2 => n6588, A => n6005, ZN => 
                           n6740);
   U12483 : NAND2_X1 port map( A1 => n6740, A2 => n7031, ZN => n6006);
   U12484 : NAND2_X1 port map( A1 => n6006, A2 => n6225, ZN => n6009);
   U12485 : INV_X1 port map( A => n6740, ZN => n6007);
   U12486 : NAND3_X1 port map( A1 => n6007, A2 => n7033, A3 => n7035, ZN => 
                           n6008);
   U12487 : NAND2_X1 port map( A1 => n24067, A2 => n6538, ZN => n6011);
   U12488 : OAI21_X1 port map( B1 => n6012, B2 => n24592, A => n6011, ZN => 
                           n6017);
   U12489 : NAND2_X1 port map( A1 => n6532, A2 => n25014, ZN => n6014);
   U12490 : AOI21_X1 port map( B1 => n6015, B2 => n6014, A => n24254, ZN => 
                           n6016);
   U12491 : OR2_X2 port map( A1 => n6017, A2 => n6016, ZN => n7600);
   U12493 : INV_X1 port map( A => n6195, ZN => n6450);
   U12494 : NAND2_X1 port map( A1 => n6450, A2 => n6445, ZN => n6018);
   U12495 : AOI21_X1 port map( B1 => n6448, B2 => n6018, A => n6196, ZN => 
                           n6022);
   U12496 : INV_X1 port map( A => Plaintext(17), ZN => n6023);
   U12498 : INV_X1 port map( A => Plaintext(16), ZN => n6024);
   U12499 : XNOR2_X1 port map( A => n6024, B => Key(16), ZN => n6324);
   U12500 : INV_X1 port map( A => Plaintext(15), ZN => n6025);
   U12501 : INV_X1 port map( A => n6519, ZN => n6156);
   U12502 : INV_X1 port map( A => Plaintext(12), ZN => n6026);
   U12503 : XNOR2_X1 port map( A => n6026, B => Key(12), ZN => n6179);
   U12504 : INV_X1 port map( A => n6179, ZN => n6323);
   U12505 : INV_X1 port map( A => n6518, ZN => n6027);
   U12506 : INV_X1 port map( A => n6275, ZN => n6274);
   U12507 : NAND2_X1 port map( A1 => n6027, A2 => n6274, ZN => n6029);
   U12508 : XNOR2_X1 port map( A => Key(13), B => Plaintext(13), ZN => n6523);
   U12509 : NAND2_X1 port map( A1 => n7595, A2 => n7602, ZN => n6802);
   U12510 : NOR2_X1 port map( A1 => n7135, A2 => n7602, ZN => n6039);
   U12511 : INV_X1 port map( A => n6510, ZN => n6459);
   U12513 : INV_X1 port map( A => n6512, ZN => n6460);
   U12514 : NOR2_X1 port map( A1 => n6513, A2 => n6456, ZN => n6506);
   U12515 : OAI21_X1 port map( B1 => n6510, B2 => n6460, A => n6506, ZN => 
                           n6031);
   U12516 : NOR2_X1 port map( A1 => n7595, A2 => n7257, ZN => n6038);
   U12517 : INV_X1 port map( A => Plaintext(10), ZN => n6033);
   U12518 : XNOR2_X1 port map( A => n6033, B => Key(10), ZN => n6496);
   U12519 : NAND2_X1 port map( A1 => n6271, A2 => n6034, ZN => n6169);
   U12520 : INV_X1 port map( A => Plaintext(7), ZN => n6035);
   U12521 : OAI21_X1 port map( B1 => n6351, B2 => n6498, A => n6168, ZN => 
                           n6037);
   U12522 : INV_X1 port map( A => Plaintext(11), ZN => n6036);
   U12523 : XNOR2_X1 port map( A => n6036, B => Key(11), ZN => n6497);
   U12524 : OAI21_X1 port map( B1 => n6039, B2 => n6038, A => n7598, ZN => 
                           n6045);
   U12525 : INV_X1 port map( A => n6133, ZN => n6136);
   U12526 : OAI211_X1 port map( C1 => n6136, C2 => n6164, A => n6265, B => 
                           n7097, ZN => n6043);
   U12527 : NAND2_X1 port map( A1 => n6266, A2 => n6539, ZN => n6040);
   U12528 : NAND3_X1 port map( A1 => n7255, A2 => n24772, A3 => n7597, ZN => 
                           n6044);
   U12529 : XNOR2_X1 port map( A => n310, B => n9181, ZN => n6046);
   U12530 : XNOR2_X1 port map( A => n9011, B => n6046, ZN => n6047);
   U12531 : XNOR2_X1 port map( A => n6048, B => n6047, ZN => n9460);
   U12532 : OAI211_X1 port map( C1 => n6750, C2 => n6409, A => n6054, B => 
                           n6053, ZN => n6056);
   U12533 : NAND3_X1 port map( A1 => n6630, A2 => n6407, A3 => n6051, ZN => 
                           n6055);
   U12534 : OAI21_X1 port map( B1 => n6964, B2 => n6963, A => n6057, ZN => 
                           n6967);
   U12536 : NAND2_X1 port map( A1 => n6570, A2 => n24089, ZN => n6576);
   U12537 : NAND2_X1 port map( A1 => n5800, A2 => n6963, ZN => n6572);
   U12538 : NAND2_X1 port map( A1 => n4754, A2 => n6575, ZN => n6059);
   U12539 : MUX2_X1 port map( A => n7747, B => n8021, S => n8022, Z => n6070);
   U12540 : NAND2_X1 port map( A1 => n6393, A2 => n6396, ZN => n6061);
   U12543 : MUX2_X1 port map( A => n6729, B => n6732, S => n6396, Z => n6063);
   U12544 : NAND2_X1 port map( A1 => n6692, A2 => n6975, ZN => n6069);
   U12545 : INV_X1 port map( A => n6976, ZN => n6568);
   U12547 : AND2_X1 port map( A1 => n6368, A2 => n6996, ZN => n6657);
   U12548 : NAND2_X1 port map( A1 => n6815, A2 => n6072, ZN => n6073);
   U12549 : NAND2_X1 port map( A1 => n6075, A2 => n6794, ZN => n6883);
   U12550 : INV_X1 port map( A => n6794, ZN => n6644);
   U12551 : NAND2_X1 port map( A1 => n6644, A2 => n6885, ZN => n6077);
   U12552 : NAND3_X1 port map( A1 => n6882, A2 => n6881, A3 => n6795, ZN => 
                           n6080);
   U12553 : INV_X1 port map( A => n6078, ZN => n6792);
   U12554 : NAND3_X1 port map( A1 => n6075, A2 => n6885, A3 => n6792, ZN => 
                           n6079);
   U12555 : NOR2_X1 port map( A1 => n7754, A2 => n7292, ZN => n7755);
   U12556 : INV_X1 port map( A => n6081, ZN => n6768);
   U12557 : NAND2_X1 port map( A1 => n6768, A2 => n6871, ZN => n6873);
   U12558 : AND2_X1 port map( A1 => n6083, A2 => n6310, ZN => n6477);
   U12559 : INV_X1 port map( A => n6477, ZN => n6082);
   U12560 : NAND2_X1 port map( A1 => n6873, A2 => n6082, ZN => n6085);
   U12561 : OAI21_X1 port map( B1 => n6874, B2 => n6870, A => n6083, ZN => 
                           n6084);
   U12562 : OAI21_X1 port map( B1 => n2522, B2 => n7542, A => n432, ZN => n6098
                           );
   U12563 : INV_X1 port map( A => n6373, ZN => n6088);
   U12564 : NAND2_X1 port map( A1 => n6087, A2 => n6377, ZN => n6093);
   U12565 : INV_X1 port map( A => n6473, ZN => n6902);
   U12567 : MUX2_X1 port map( A => n6091, B => n6090, S => n6906, Z => n6092);
   U12568 : NAND2_X1 port map( A1 => n7006, A2 => n7007, ZN => n6383);
   U12569 : INV_X1 port map( A => n6383, ZN => n6096);
   U12570 : INV_X1 port map( A => n7004, ZN => n6832);
   U12571 : OAI21_X1 port map( B1 => n6096, B2 => n6095, A => n6094, ZN => 
                           n6097);
   U12572 : XNOR2_X1 port map( A => n8674, B => n8604, ZN => n8256);
   U12573 : INV_X1 port map( A => n6602, ZN => n7012);
   U12574 : INV_X1 port map( A => n6827, ZN => n7014);
   U12575 : NAND2_X1 port map( A1 => n7012, A2 => n7014, ZN => n6101);
   U12576 : INV_X1 port map( A => n6598, ZN => n6601);
   U12577 : MUX2_X1 port map( A => n6101, B => n6099, S => n7015, Z => n6103);
   U12578 : NAND3_X1 port map( A1 => n6826, A2 => n6101, A3 => n7019, ZN => 
                           n6102);
   U12579 : NAND2_X1 port map( A1 => n6104, A2 => n7029, ZN => n6593);
   U12580 : NAND2_X1 port map( A1 => n6593, A2 => n6105, ZN => n6108);
   U12581 : NAND2_X1 port map( A1 => n7029, A2 => n7032, ZN => n6106);
   U12582 : OAI21_X1 port map( B1 => n7030, B2 => n7029, A => n6106, ZN => 
                           n6107);
   U12583 : AND2_X1 port map( A1 => n7768, A2 => n7526, ZN => n6113);
   U12584 : OAI21_X1 port map( B1 => n6845, B2 => n7021, A => n6846, ZN => 
                           n6109);
   U12585 : INV_X1 port map( A => n6715, ZN => n6610);
   U12586 : INV_X1 port map( A => n6712, ZN => n6606);
   U12587 : NAND2_X1 port map( A1 => n5796, A2 => n6114, ZN => n6728);
   U12588 : AOI21_X1 port map( B1 => n6728, B2 => n6115, A => n6622, ZN => 
                           n6118);
   U12589 : NAND2_X1 port map( A1 => n6622, A2 => n6114, ZN => n6116);
   U12590 : AOI21_X1 port map( B1 => n6116, B2 => n6724, A => n6722, ZN => 
                           n6117);
   U12591 : NOR2_X1 port map( A1 => n7768, A2 => n7527, ZN => n6126);
   U12592 : INV_X1 port map( A => n6987, ZN => n6991);
   U12593 : INV_X1 port map( A => n6119, ZN => n6988);
   U12594 : INV_X1 port map( A => n6642, ZN => n6120);
   U12595 : NAND2_X1 port map( A1 => n6120, A2 => n6990, ZN => n6125);
   U12596 : OAI21_X1 port map( B1 => n6988, B2 => n6244, A => n6841, ZN => 
                           n6121);
   U12597 : INV_X1 port map( A => n6640, ZN => n6838);
   U12598 : INV_X1 port map( A => n6989, ZN => n6123);
   U12600 : INV_X1 port map( A => n24592, ZN => n6128);
   U12602 : AOI21_X1 port map( B1 => n6264, B2 => n6130, A => n6531, ZN => 
                           n6131);
   U12603 : AOI21_X1 port map( B1 => n5916, B2 => n6543, A => n6539, ZN => 
                           n6135);
   U12604 : NAND2_X1 port map( A1 => n6136, A2 => n6165, ZN => n6540);
   U12605 : INV_X1 port map( A => n7384, ZN => n7618);
   U12606 : OAI21_X1 port map( B1 => n7385, B2 => n7618, A => n7386, ZN => 
                           n6152);
   U12607 : NAND2_X1 port map( A1 => n6950, A2 => n25437, ZN => n6138);
   U12608 : AND3_X1 port map( A1 => n6139, A2 => n6528, A3 => n6138, ZN => 
                           n6158);
   U12609 : INV_X1 port map( A => n6158, ZN => n6140);
   U12610 : AND2_X1 port map( A1 => n6540, A2 => n6140, ZN => n6143);
   U12611 : NAND3_X1 port map( A1 => n25437, A2 => n6948, A3 => n24994, ZN => 
                           n6141);
   U12612 : INV_X1 port map( A => n6157, ZN => n6142);
   U12613 : MUX2_X1 port map( A => n6145, B => n6144, S => n6281, Z => n6149);
   U12614 : INV_X1 port map( A => n6146, ZN => n6678);
   U12615 : NAND2_X1 port map( A1 => n7385, A2 => n7619, ZN => n6150);
   U12616 : NAND3_X1 port map( A1 => n6152, A2 => n6151, A3 => n6150, ZN => 
                           n6160);
   U12617 : NAND2_X1 port map( A1 => n1509, A2 => n6156, ZN => n6153);
   U12618 : NAND3_X1 port map( A1 => n7622, A2 => n1895, A3 => n7386, ZN => 
                           n6159);
   U12619 : XNOR2_X1 port map( A => n9194, B => n8824, ZN => n6161);
   U12620 : XNOR2_X1 port map( A => n8256, B => n6161, ZN => n6222);
   U12621 : OAI21_X1 port map( B1 => n6164, B2 => n6539, A => n5916, ZN => 
                           n6166);
   U12622 : INV_X1 port map( A => n6165, ZN => n6542);
   U12623 : INV_X1 port map( A => n7761, ZN => n7307);
   U12624 : OAI22_X1 port map( A1 => n6351, A2 => n6169, B1 => n6168, B2 => 
                           n6503, ZN => n6172);
   U12625 : NAND2_X1 port map( A1 => n6351, A2 => n6034, ZN => n6170);
   U12626 : INV_X1 port map( A => n6497, ZN => n6350);
   U12627 : INV_X1 port map( A => n7760, ZN => n7305);
   U12628 : AOI21_X1 port map( B1 => n6173, B2 => n6296, A => n6438, ZN => 
                           n6178);
   U12629 : NAND2_X1 port map( A1 => n6297, A2 => n6438, ZN => n6175);
   U12630 : AOI21_X1 port map( B1 => n6176, B2 => n6175, A => n6332, ZN => 
                           n6177);
   U12631 : NAND2_X1 port map( A1 => n6524, A2 => n944, ZN => n6181);
   U12632 : NOR2_X1 port map( A1 => n25427, A2 => n6455, ZN => n6182);
   U12633 : OAI21_X1 port map( B1 => n6183, B2 => n6182, A => n6510, ZN => 
                           n6186);
   U12634 : NAND2_X1 port map( A1 => n6457, A2 => n6512, ZN => n6338);
   U12635 : OAI211_X1 port map( C1 => n25427, C2 => n6457, A => n6338, B => 
                           n6459, ZN => n6185);
   U12637 : INV_X1 port map( A => n7647, ZN => n6191);
   U12638 : NAND2_X1 port map( A1 => n6187, A2 => n6452, ZN => n6188);
   U12639 : NAND2_X1 port map( A1 => n6449, A2 => n6447, ZN => n6189);
   U12640 : NAND2_X1 port map( A1 => n6191, A2 => n7651, ZN => n6190);
   U12641 : NAND3_X1 port map( A1 => n6191, A2 => n7651, A3 => n7760, ZN => 
                           n6192);
   U12642 : OAI211_X1 port map( C1 => n7307, C2 => n6194, A => n6193, B => 
                           n6192, ZN => n9196);
   U12643 : OAI21_X1 port map( B1 => n6344, B2 => n6444, A => n6341, ZN => 
                           n6197);
   U12644 : NAND2_X1 port map( A1 => n25401, A2 => n6488, ZN => n6785);
   U12645 : INV_X1 port map( A => n6493, ZN => n6429);
   U12646 : NAND2_X1 port map( A1 => n6489, A2 => n6490, ZN => n6303);
   U12647 : INV_X1 port map( A => n6777, ZN => n6925);
   U12648 : INV_X1 port map( A => n7294, ZN => n7749);
   U12649 : NAND2_X1 port map( A1 => n6915, A2 => n6918, ZN => n6774);
   U12650 : INV_X1 port map( A => n6915, ZN => n6910);
   U12651 : NAND2_X1 port map( A1 => n6910, A2 => n24509, ZN => n6201);
   U12652 : INV_X1 port map( A => n6912, ZN => n6771);
   U12653 : NAND2_X1 port map( A1 => n24037, A2 => n6771, ZN => n6200);
   U12654 : NOR2_X1 port map( A1 => n6910, A2 => n6771, ZN => n6202);
   U12655 : NAND2_X1 port map( A1 => n7749, A2 => n7537, ZN => n6206);
   U12657 : INV_X1 port map( A => n6467, ZN => n6326);
   U12658 : NAND2_X1 port map( A1 => n6326, A2 => n6315, ZN => n6204);
   U12659 : MUX2_X1 port map( A => n6204, B => n6203, S => n5451, Z => n6205);
   U12660 : MUX2_X1 port map( A => n6207, B => n6206, S => n8014, Z => n6215);
   U12661 : INV_X1 port map( A => n6208, ZN => n6294);
   U12662 : NAND2_X1 port map( A1 => n6294, A2 => n6438, ZN => n6298);
   U12663 : NAND2_X1 port map( A1 => n6298, A2 => n6335, ZN => n6443);
   U12665 : INV_X1 port map( A => n6332, ZN => n6295);
   U12666 : NAND3_X1 port map( A1 => n6212, A2 => n6334, A3 => n6211, ZN => 
                           n6213);
   U12667 : XNOR2_X1 port map( A => n8935, B => n9196, ZN => n8034);
   U12668 : INV_X1 port map( A => n7347, ZN => n6216);
   U12669 : NAND2_X1 port map( A1 => n6216, A2 => n7346, ZN => n6217);
   U12670 : OAI21_X1 port map( B1 => n8508, B2 => n7346, A => n6217, ZN => 
                           n6218);
   U12671 : XNOR2_X1 port map( A => n8341, B => n1863, ZN => n6220);
   U12672 : XNOR2_X1 port map( A => n8034, B => n6220, ZN => n6221);
   U12673 : INV_X1 port map( A => n7619, ZN => n7617);
   U12674 : MUX2_X1 port map( A => n7617, B => n7382, S => n7615, Z => n6224);
   U12676 : MUX2_X2 port map( A => n6224, B => n6223, S => n7380, Z => n8333);
   U12677 : NAND3_X1 port map( A1 => n6226, A2 => n6225, A3 => n6104, ZN => 
                           n6229);
   U12678 : NAND3_X1 port map( A1 => n7032, A2 => n7029, A3 => n7033, ZN => 
                           n6228);
   U12679 : NAND2_X1 port map( A1 => n6823, A2 => n6598, ZN => n6829);
   U12680 : INV_X1 port map( A => n7013, ZN => n6822);
   U12681 : NAND3_X1 port map( A1 => n6829, A2 => n25044, A3 => n6230, ZN => 
                           n6231);
   U12682 : NAND2_X1 port map( A1 => n6234, A2 => n6233, ZN => n6609);
   U12683 : INV_X1 port map( A => n6235, ZN => n6718);
   U12685 : INV_X1 port map( A => n6238, ZN => n6395);
   U12686 : INV_X1 port map( A => n6732, ZN => n6397);
   U12687 : NAND3_X1 port map( A1 => n6397, A2 => n6729, A3 => n6238, ZN => 
                           n6241);
   U12688 : INV_X1 port map( A => n6396, ZN => n6239);
   U12689 : NAND2_X1 port map( A1 => n6733, A2 => n6239, ZN => n6240);
   U12690 : INV_X1 port map( A => n6622, ZN => n6727);
   U12691 : MUX2_X1 port map( A => n7732, B => n7731, S => n7733, Z => n6250);
   U12692 : NAND2_X1 port map( A1 => n6986, A2 => n6245, ZN => n6246);
   U12693 : AOI21_X1 port map( B1 => n6840, B2 => n6246, A => n6640, ZN => 
                           n6249);
   U12694 : AOI21_X1 port map( B1 => n6247, B2 => n6988, A => n6245, ZN => 
                           n6248);
   U12695 : INV_X1 port map( A => n8806, ZN => n6252);
   U12696 : XNOR2_X1 port map( A => n8333, B => n6252, ZN => n8398);
   U12697 : INV_X1 port map( A => n8398, ZN => n6322);
   U12698 : NAND2_X1 port map( A1 => n6253, A2 => n24994, ZN => n6254);
   U12699 : NAND3_X1 port map( A1 => n6255, A2 => n6947, A3 => n6529, ZN => 
                           n6257);
   U12700 : NAND3_X1 port map( A1 => n6952, A2 => n25437, A3 => n6528, ZN => 
                           n6256);
   U12702 : NAND3_X1 port map( A1 => n6530, A2 => n6531, A3 => n6538, ZN => 
                           n6262);
   U12703 : OAI211_X1 port map( C1 => n6264, C2 => n24067, A => n6263, B => 
                           n6262, ZN => n6280);
   U12704 : NAND2_X1 port map( A1 => n6164, A2 => n6266, ZN => n6544);
   U12705 : NAND2_X1 port map( A1 => n7103, A2 => n6539, ZN => n6268);
   U12706 : NAND2_X1 port map( A1 => n6544, A2 => n6268, ZN => n6269);
   U12708 : MUX2_X1 port map( A => n7798, B => n7802, S => n7800, Z => n6285);
   U12709 : INV_X1 port map( A => n6280, ZN => n7432);
   U12710 : NAND2_X1 port map( A1 => n6351, A2 => n441, ZN => n6272);
   U12711 : MUX2_X1 port map( A => n6434, B => n6272, S => n6498, Z => n6273);
   U12712 : NAND2_X1 port map( A1 => n7432, A2 => n7803, ZN => n7797);
   U12713 : AND2_X1 port map( A1 => n440, A2 => n6274, ZN => n6279);
   U12714 : NAND2_X1 port map( A1 => n6275, A2 => n6521, ZN => n6276);
   U12715 : NAND2_X1 port map( A1 => n7797, A2 => n7053, ZN => n6284);
   U12717 : AOI21_X1 port map( B1 => n6945, B2 => n6943, A => n6939, ZN => 
                           n6283);
   U12718 : INV_X1 port map( A => n6770, ZN => n6911);
   U12719 : AND2_X1 port map( A1 => n6771, A2 => n6911, ZN => n6289);
   U12720 : INV_X1 port map( A => n6918, ZN => n6286);
   U12722 : NAND2_X1 port map( A1 => n6909, A2 => n24037, ZN => n6287);
   U12723 : OAI211_X2 port map( C1 => n6289, C2 => n6774, A => n6288, B => 
                           n6287, ZN => n7707);
   U12724 : INV_X1 port map( A => n7707, ZN => n7867);
   U12726 : NAND2_X1 port map( A1 => n6925, A2 => n6775, ZN => n6291);
   U12727 : NAND2_X1 port map( A1 => n6294, A2 => n6297, ZN => n6336);
   U12728 : AOI21_X1 port map( B1 => n6334, B2 => n6336, A => n6295, ZN => 
                           n6300);
   U12729 : INV_X1 port map( A => n6784, ZN => n6487);
   U12730 : MUX2_X1 port map( A => n6303, B => n6302, S => n6493, Z => n6307);
   U12731 : INV_X1 port map( A => n7863, ZN => n7860);
   U12732 : INV_X1 port map( A => n6767, ZN => n6309);
   U12733 : OAI21_X1 port map( B1 => n6876, B2 => n6309, A => n6875, ZN => 
                           n6308);
   U12734 : NAND2_X1 port map( A1 => n6308, A2 => n4922, ZN => n6313);
   U12735 : NAND3_X1 port map( A1 => n6310, A2 => n6874, A3 => n6309, ZN => 
                           n6311);
   U12736 : NAND2_X1 port map( A1 => n3570, A2 => n7861, ZN => n6319);
   U12737 : NAND3_X1 port map( A1 => n6315, A2 => n6329, A3 => n25404, ZN => 
                           n6317);
   U12738 : NAND3_X1 port map( A1 => n6326, A2 => n5451, A3 => n5966, ZN => 
                           n6316);
   U12740 : XNOR2_X1 port map( A => n9155, B => n25235, ZN => n6321);
   U12741 : XNOR2_X1 port map( A => n6322, B => n6321, ZN => n6423);
   U12742 : AOI21_X1 port map( B1 => n6519, B2 => n1509, A => n6323, ZN => 
                           n6325);
   U12743 : OAI21_X1 port map( B1 => n6328, B2 => n5451, A => n6327, ZN => 
                           n6331);
   U12744 : NAND3_X1 port map( A1 => n6440, A2 => n6209, A3 => n6438, ZN => 
                           n6333);
   U12745 : OAI211_X1 port map( C1 => n6336, C2 => n6335, A => n6334, B => 
                           n6333, ZN => n7057);
   U12746 : INV_X1 port map( A => n6456, ZN => n6339);
   U12747 : NAND3_X1 port map( A1 => n25428, A2 => n6339, A3 => n6509, ZN => 
                           n6340);
   U12748 : MUX2_X1 port map( A => n9066, B => n7057, S => n9067, Z => n6355);
   U12749 : NAND2_X1 port map( A1 => n6341, A2 => n6447, ZN => n6343);
   U12750 : NAND2_X1 port map( A1 => n6452, A2 => n6445, ZN => n6342);
   U12751 : AND2_X1 port map( A1 => n6343, A2 => n6342, ZN => n6349);
   U12752 : INV_X1 port map( A => n6344, ZN => n6346);
   U12753 : NOR2_X1 port map( A1 => n7809, A2 => n8219, ZN => n7814);
   U12754 : NAND2_X1 port map( A1 => n6496, A2 => n6350, ZN => n6353);
   U12755 : INV_X1 port map( A => n6351, ZN => n6499);
   U12757 : NOR2_X1 port map( A1 => n7813, A2 => n8219, ZN => n7196);
   U12758 : INV_X1 port map( A => n9067, ZN => n7738);
   U12759 : OAI22_X1 port map( A1 => n7814, A2 => n7196, B1 => n7738, B2 => 
                           n7809, ZN => n6354);
   U12760 : OAI21_X2 port map( B1 => n6355, B2 => n7812, A => n6354, ZN => 
                           n8278);
   U12761 : NAND2_X1 port map( A1 => n6818, A2 => n6893, ZN => n6356);
   U12762 : AOI21_X1 port map( B1 => n6357, B2 => n6356, A => n6358, ZN => 
                           n6361);
   U12763 : NAND3_X1 port map( A1 => n6651, A2 => n6358, A3 => n6893, ZN => 
                           n6360);
   U12764 : OR3_X1 port map( A1 => n6819, A2 => n6895, A3 => n6893, ZN => n6359
                           );
   U12765 : NAND2_X1 port map( A1 => n6793, A2 => n6078, ZN => n6363);
   U12766 : INV_X1 port map( A => n6363, ZN => n6366);
   U12767 : OAI21_X1 port map( B1 => n6078, B2 => n6794, A => n6882, ZN => 
                           n6365);
   U12768 : MUX2_X1 port map( A => n6363, B => n6362, S => n6885, Z => n6364);
   U12771 : OAI21_X1 port map( B1 => n6072, B2 => n6369, A => n6071, ZN => 
                           n6370);
   U12772 : OAI21_X1 port map( B1 => n6899, B2 => n6373, A => n6377, ZN => 
                           n6378);
   U12774 : OAI21_X1 port map( B1 => n6848, B2 => n7021, A => n6845, ZN => 
                           n6380);
   U12775 : NAND2_X1 port map( A1 => n7022, A2 => n7026, ZN => n6379);
   U12776 : NAND3_X1 port map( A1 => n7025, A2 => n250, A3 => n4643, ZN => 
                           n6382);
   U12777 : AND2_X1 port map( A1 => n6094, A2 => n7005, ZN => n6387);
   U12778 : NAND2_X1 port map( A1 => n6832, A2 => n7008, ZN => n6386);
   U12779 : OAI21_X1 port map( B1 => n6384, B2 => n7007, A => n6383, ZN => 
                           n6385);
   U12780 : XNOR2_X1 port map( A => n8278, B => n8615, ZN => n6421);
   U12781 : OAI21_X1 port map( B1 => n6975, B2 => n1149, A => n24395, ZN => 
                           n6391);
   U12782 : AND2_X1 port map( A1 => n1149, A2 => n6688, ZN => n6389);
   U12783 : NAND2_X1 port map( A1 => n6393, A2 => n6392, ZN => n6394);
   U12784 : AOI21_X1 port map( B1 => n6397, B2 => n6733, A => n6396, ZN => 
                           n6398);
   U12785 : NAND2_X1 port map( A1 => n271, A2 => n6400, ZN => n6403);
   U12786 : INV_X1 port map( A => n6400, ZN => n6674);
   U12787 : NAND2_X1 port map( A1 => n6674, A2 => n6757, ZN => n6401);
   U12788 : NAND2_X1 port map( A1 => n7563, A2 => n7721, ZN => n7858);
   U12789 : NAND2_X1 port map( A1 => n6965, A2 => n6963, ZN => n6405);
   U12790 : NAND2_X1 port map( A1 => n6964, A2 => n5800, ZN => n6404);
   U12791 : OAI21_X1 port map( B1 => n7184, B2 => n4752, A => n6406, ZN => 
                           n6413);
   U12792 : INV_X1 port map( A => n6630, ZN => n6565);
   U12793 : INV_X1 port map( A => n6407, ZN => n6746);
   U12794 : NAND2_X1 port map( A1 => n453, A2 => n6407, ZN => n6408);
   U12795 : INV_X1 port map( A => n7853, ZN => n7564);
   U12796 : INV_X1 port map( A => n7563, ZN => n7854);
   U12797 : INV_X1 port map( A => n6414, ZN => n6698);
   U12798 : NAND2_X1 port map( A1 => n6698, A2 => n6694, ZN => n6558);
   U12799 : INV_X1 port map( A => n6697, ZN => n6559);
   U12800 : NOR2_X1 port map( A1 => n6695, A2 => n6559, ZN => n6416);
   U12801 : NOR2_X1 port map( A1 => n7857, A2 => n7721, ZN => n7849);
   U12802 : NAND2_X1 port map( A1 => n7849, A2 => n7563, ZN => n6418);
   U12803 : OAI211_X1 port map( C1 => n24072, C2 => n7858, A => n6419, B => 
                           n6418, ZN => n8588);
   U12804 : XNOR2_X1 port map( A => n8588, B => n1739, ZN => n6420);
   U12805 : XNOR2_X1 port map( A => n6421, B => n6420, ZN => n6422);
   U12806 : XNOR2_X1 port map( A => n6423, B => n6422, ZN => n9462);
   U12809 : NAND2_X1 port map( A1 => n6470, A2 => n6426, ZN => n6469);
   U12810 : NAND2_X1 port map( A1 => n25401, A2 => n6784, ZN => n6494);
   U12811 : NAND2_X1 port map( A1 => n6429, A2 => n6490, ZN => n6428);
   U12812 : AOI21_X1 port map( B1 => n6494, B2 => n6428, A => n6301, ZN => 
                           n6433);
   U12813 : NAND2_X1 port map( A1 => n6429, A2 => n6489, ZN => n6431);
   U12814 : AOI21_X1 port map( B1 => n6431, B2 => n6430, A => n6490, ZN => 
                           n6432);
   U12816 : NAND2_X1 port map( A1 => n6497, A2 => n6034, ZN => n6501);
   U12817 : OAI21_X1 port map( B1 => n6499, B2 => n6498, A => n24466, ZN => 
                           n6436);
   U12818 : NOR2_X1 port map( A1 => n6438, A2 => n6209, ZN => n6442);
   U12819 : NAND2_X1 port map( A1 => n7085, A2 => n433, ZN => n6466);
   U12820 : NAND3_X1 port map( A1 => n6445, A2 => n6449, A3 => n6444, ZN => 
                           n6446);
   U12821 : OAI21_X1 port map( B1 => n6448, B2 => n6447, A => n6446, ZN => 
                           n7689);
   U12823 : NOR2_X1 port map( A1 => n7689, A2 => n7691, ZN => n7147);
   U12824 : INV_X1 port map( A => n7147, ZN => n8317);
   U12825 : NOR2_X1 port map( A1 => n8317, A2 => n8315, ZN => n6465);
   U12826 : INV_X1 port map( A => n25428, ZN => n6464);
   U12827 : NAND2_X1 port map( A1 => n6454, A2 => n6510, ZN => n6463);
   U12828 : NAND2_X1 port map( A1 => n6456, A2 => n6455, ZN => n6458);
   U12829 : OAI211_X1 port map( C1 => n6455, C2 => n6464, A => n6458, B => 
                           n6457, ZN => n6462);
   U12830 : NAND3_X1 port map( A1 => n6460, A2 => n6459, A3 => n6509, ZN => 
                           n6461);
   U12833 : INV_X1 port map( A => n9147, ZN => n8152);
   U12834 : AOI21_X1 port map( B1 => n6471, B2 => n6470, A => n5966, ZN => 
                           n6472);
   U12835 : NAND2_X1 port map( A1 => n6372, A2 => n6473, ZN => n6474);
   U12836 : NAND2_X1 port map( A1 => n6477, A2 => n6876, ZN => n6478);
   U12837 : AND2_X1 port map( A1 => n6874, A2 => n6870, ZN => n6879);
   U12838 : NOR2_X1 port map( A1 => n6480, A2 => n6775, ZN => n6479);
   U12839 : NAND2_X1 port map( A1 => n6915, A2 => n24509, ZN => n6769);
   U12840 : NAND2_X1 port map( A1 => n24037, A2 => n6915, ZN => n6483);
   U12841 : OAI211_X1 port map( C1 => n6912, C2 => n24037, A => n6483, B => 
                           n6911, ZN => n6484);
   U12842 : NAND2_X1 port map( A1 => n7638, A2 => n7917, ZN => n7635);
   U12843 : INV_X1 port map( A => n6489, ZN => n6783);
   U12844 : NAND3_X1 port map( A1 => n6490, A2 => n6783, A3 => n6493, ZN => 
                           n6491);
   U12845 : XNOR2_X1 port map( A => n8152, B => n8908, ZN => n8050);
   U12846 : OR2_X1 port map( A1 => n6497, A2 => n6496, ZN => n6500);
   U12848 : INV_X1 port map( A => n6506, ZN => n6508);
   U12849 : NAND2_X1 port map( A1 => n6508, A2 => n6507, ZN => n6516);
   U12850 : NAND2_X1 port map( A1 => n6509, A2 => n6512, ZN => n6511);
   U12851 : NAND2_X1 port map( A1 => n6511, A2 => n6510, ZN => n6515);
   U12852 : NOR2_X1 port map( A1 => n25427, A2 => n6512, ZN => n6514);
   U12853 : INV_X1 port map( A => n6806, ZN => n8531);
   U12854 : NAND2_X1 port map( A1 => n6519, A2 => n25398, ZN => n6520);
   U12855 : NAND2_X1 port map( A1 => n6524, A2 => n6523, ZN => n6525);
   U12856 : NAND3_X1 port map( A1 => n6947, A2 => n5903, A3 => n6950, ZN => 
                           n6527);
   U12857 : OAI21_X1 port map( B1 => n7087, B2 => n8531, A => n6548, ZN => 
                           n6860);
   U12858 : NAND2_X1 port map( A1 => n6532, A2 => n6531, ZN => n6536);
   U12859 : NAND2_X1 port map( A1 => n24254, A2 => n6538, ZN => n6535);
   U12860 : MUX2_X1 port map( A => n6536, B => n6535, S => n24067, Z => n6537);
   U12861 : MUX2_X1 port map( A => n6540, B => n7098, S => n6539, Z => n6547);
   U12862 : MUX2_X1 port map( A => n6545, B => n6544, S => n6543, Z => n6546);
   U12863 : OAI211_X1 port map( C1 => n8531, C2 => n7663, A => n6549, B => 
                           n6548, ZN => n6550);
   U12867 : NAND2_X1 port map( A1 => n6553, A2 => n5924, ZN => n6555);
   U12868 : NAND3_X1 port map( A1 => n3923, A2 => n6702, A3 => n6959, ZN => 
                           n6554);
   U12870 : INV_X1 port map( A => n6933, ZN => n6557);
   U12871 : NAND2_X1 port map( A1 => n6557, A2 => n6556, ZN => n6563);
   U12872 : INV_X1 port map( A => n6558, ZN => n6937);
   U12873 : NAND2_X1 port map( A1 => n6560, A2 => n2008, ZN => n6561);
   U12874 : NAND2_X1 port map( A1 => n7445, A2 => n7444, ZN => n7262);
   U12875 : NAND2_X1 port map( A1 => n6746, A2 => n453, ZN => n6564);
   U12876 : AOI21_X1 port map( B1 => n6748, B2 => n6564, A => n6744, ZN => 
                           n7928);
   U12877 : NAND2_X1 port map( A1 => n6565, A2 => n453, ZN => n6566);
   U12878 : OR2_X1 port map( A1 => n7262, A2 => n5607, ZN => n6586);
   U12879 : AOI21_X1 port map( B1 => n24579, B2 => n6688, A => n6687, ZN => 
                           n6974);
   U12880 : OAI211_X1 port map( C1 => n6977, C2 => n6568, A => n6567, B => 
                           n24395, ZN => n6569);
   U12881 : NAND3_X1 port map( A1 => n6572, A2 => n6969, A3 => n6571, ZN => 
                           n6574);
   U12882 : NAND3_X1 port map( A1 => n4754, A2 => n6964, A3 => n5800, ZN => 
                           n6573);
   U12883 : OAI211_X2 port map( C1 => n6576, C2 => n6575, A => n6574, B => 
                           n6573, ZN => n7932);
   U12884 : NOR2_X1 port map( A1 => n7444, A2 => n7932, ZN => n6583);
   U12885 : NAND2_X1 port map( A1 => n6583, A2 => n5607, ZN => n6585);
   U12886 : INV_X1 port map( A => n6577, ZN => n6758);
   U12887 : NAND2_X1 port map( A1 => n6675, A2 => n6758, ZN => n6580);
   U12888 : INV_X1 port map( A => n6757, ZN => n6673);
   U12889 : MUX2_X1 port map( A => n6580, B => n6579, S => n6578, Z => n6581);
   U12890 : NAND2_X1 port map( A1 => n6583, A2 => n7924, ZN => n6584);
   U12891 : XNOR2_X1 port map( A => n8484, B => n8634, ZN => n6587);
   U12892 : XNOR2_X1 port map( A => n8050, B => n6587, ZN => n6666);
   U12893 : INV_X1 port map( A => n7035, ZN => n6739);
   U12894 : NAND2_X1 port map( A1 => n6588, A2 => n7032, ZN => n6590);
   U12895 : MUX2_X1 port map( A => n6591, B => n6590, S => n25424, Z => n6595);
   U12896 : INV_X1 port map( A => n7032, ZN => n6592);
   U12898 : NAND2_X1 port map( A1 => n6597, A2 => n25045, ZN => n6605);
   U12901 : NAND2_X1 port map( A1 => n24090, A2 => n6822, ZN => n6604);
   U12902 : NAND2_X1 port map( A1 => n25044, A2 => n6601, ZN => n6603);
   U12903 : INV_X1 port map( A => n6609, ZN => n6612);
   U12904 : NAND2_X1 port map( A1 => n6393, A2 => n6615, ZN => n6616);
   U12905 : INV_X1 port map( A => n7787, ZN => n6618);
   U12906 : NAND2_X1 port map( A1 => n6619, A2 => n6722, ZN => n6620);
   U12907 : AOI21_X1 port map( B1 => n6621, B2 => n6620, A => n6723, ZN => 
                           n6627);
   U12908 : NAND2_X1 port map( A1 => n6622, A2 => n5796, ZN => n6625);
   U12909 : AOI21_X1 port map( B1 => n6625, B2 => n6624, A => n6114, ZN => 
                           n6626);
   U12910 : INV_X1 port map( A => n7789, ZN => n7783);
   U12911 : NAND2_X1 port map( A1 => n6629, A2 => n6628, ZN => n6632);
   U12912 : AND2_X1 port map( A1 => n6630, A2 => n4696, ZN => n6631);
   U12913 : AOI22_X1 port map( A1 => n7783, A2 => n7418, B1 => n7787, B2 => 
                           n7788, ZN => n7045);
   U12916 : NAND2_X1 port map( A1 => n7025, A2 => n250, ZN => n6637);
   U12917 : NAND2_X1 port map( A1 => n442, A2 => n4643, ZN => n6636);
   U12918 : INV_X1 port map( A => n7908, ZN => n7450);
   U12919 : NAND2_X1 port map( A1 => n7450, A2 => n7629, ZN => n7626);
   U12920 : OAI21_X1 port map( B1 => n6794, B2 => n6792, A => n6643, ZN => 
                           n6889);
   U12921 : NAND2_X1 port map( A1 => n6889, A2 => n6795, ZN => n6646);
   U12922 : AOI21_X1 port map( B1 => n6793, B2 => n6644, A => n6792, ZN => 
                           n6645);
   U12923 : NAND2_X1 port map( A1 => n6648, A2 => n7008, ZN => n6649);
   U12924 : MUX2_X1 port map( A => n6895, B => n6818, S => n6890, Z => n6656);
   U12925 : NAND2_X1 port map( A1 => n6819, A2 => n6895, ZN => n6654);
   U12926 : INV_X1 port map( A => n6893, ZN => n6652);
   U12927 : MUX2_X1 port map( A => n6654, B => n6653, S => n6652, Z => n6655);
   U12928 : OAI21_X1 port map( B1 => n6656, B2 => n313, A => n6655, ZN => n7909
                           );
   U12929 : NAND3_X1 port map( A1 => n6658, A2 => n6997, A3 => n439, ZN => 
                           n6659);
   U12930 : XNOR2_X1 port map( A => n8635, B => n8699, ZN => n6664);
   U12931 : INV_X1 port map( A => n7801, ZN => n7799);
   U12932 : NAND3_X1 port map( A1 => n7799, A2 => n7803, A3 => n7166, ZN => 
                           n6662);
   U12933 : INV_X1 port map( A => n7166, ZN => n7794);
   U12934 : OAI211_X1 port map( C1 => n7801, C2 => n7798, A => n7432, B => 
                           n7794, ZN => n6661);
   U12935 : NAND2_X1 port map( A1 => n7800, A2 => n7801, ZN => n6660);
   U12936 : NAND3_X1 port map( A1 => n6662, A2 => n6661, A3 => n6660, ZN => 
                           n8361);
   U12937 : XNOR2_X1 port map( A => n8361, B => n447, ZN => n6663);
   U12938 : XNOR2_X1 port map( A => n6664, B => n6663, ZN => n6665);
   U12939 : XNOR2_X1 port map( A => n6666, B => n6665, ZN => n9463);
   U12940 : NAND2_X1 port map( A1 => n24944, A2 => n9463, ZN => n9921);
   U12941 : INV_X1 port map( A => n6964, ZN => n6668);
   U12942 : OAI21_X1 port map( B1 => n6668, B2 => n6963, A => n24089, ZN => 
                           n6671);
   U12943 : NAND2_X1 port map( A1 => n443, A2 => n6969, ZN => n6669);
   U12944 : AOI22_X1 port map( A1 => n6673, A2 => n6675, B1 => n6758, B2 => 
                           n6674, ZN => n6677);
   U12945 : NAND3_X1 port map( A1 => n6680, A2 => n6679, A3 => n6939, ZN => 
                           n6681);
   U12946 : AND2_X1 port map( A1 => n7414, A2 => n7415, ZN => n6711);
   U12947 : NAND3_X1 port map( A1 => n6688, A2 => n6975, A3 => n6687, ZN => 
                           n6689);
   U12948 : INV_X1 port map( A => n7413, ZN => n7998);
   U12949 : NAND2_X1 port map( A1 => n6695, A2 => n6694, ZN => n6696);
   U12950 : AND2_X1 port map( A1 => n6696, A2 => n6935, ZN => n6701);
   U12951 : OAI21_X1 port map( B1 => n6699, B2 => n6698, A => n6936, ZN => 
                           n6700);
   U12954 : NAND2_X1 port map( A1 => n6960, A2 => n24405, ZN => n6707);
   U12955 : NAND3_X1 port map( A1 => n3923, A2 => n5924, A3 => n6705, ZN => 
                           n6706);
   U12956 : NAND3_X1 port map( A1 => n6708, A2 => n6707, A3 => n6706, ZN => 
                           n7412);
   U12957 : INV_X1 port map( A => n7412, ZN => n7990);
   U12958 : NOR2_X1 port map( A1 => n7413, A2 => n7990, ZN => n6709);
   U12959 : OAI21_X1 port map( B1 => n7498, B2 => n6709, A => n7357, ZN => 
                           n6710);
   U12960 : INV_X1 port map( A => n8846, ZN => n8576);
   U12961 : NOR2_X1 port map( A1 => n24501, A2 => n6714, ZN => n6716);
   U12962 : NAND3_X1 port map( A1 => n6724, A2 => n6723, A3 => n6722, ZN => 
                           n6725);
   U12963 : NAND2_X1 port map( A1 => n6869, A2 => n25251, ZN => n6743);
   U12964 : INV_X1 port map( A => n6868, ZN => n6738);
   U12965 : NAND2_X1 port map( A1 => n6733, A2 => n6732, ZN => n6735);
   U12966 : INV_X1 port map( A => n6867, ZN => n6737);
   U12967 : NAND4_X1 port map( A1 => n7506, A2 => n6738, A3 => n1379, A4 => 
                           n6737, ZN => n7672);
   U12968 : AOI21_X1 port map( B1 => n7030, B2 => n454, A => n7032, ZN => n6742
                           );
   U12969 : AOI21_X1 port map( B1 => n6743, B2 => n7672, A => n7676, ZN => 
                           n6761);
   U12970 : INV_X1 port map( A => n25251, ZN => n7677);
   U12971 : AND2_X1 port map( A1 => n6744, A2 => n6051, ZN => n6749);
   U12972 : NAND2_X1 port map( A1 => n7677, A2 => n7674, ZN => n6759);
   U12973 : OAI22_X1 port map( A1 => n6869, A2 => n6759, B1 => n7677, B2 => 
                           n3275, ZN => n6760);
   U12975 : NAND2_X1 port map( A1 => n7591, A2 => n7590, ZN => n7337);
   U12976 : OAI21_X1 port map( B1 => n7464, B2 => n7592, A => n7462, ZN => 
                           n6762);
   U12977 : OAI21_X1 port map( B1 => n6876, B2 => n6875, A => n6874, ZN => 
                           n6766);
   U12978 : NAND3_X1 port map( A1 => n6768, A2 => n4922, A3 => n6870, ZN => 
                           n6765);
   U12979 : INV_X1 port map( A => n6769, ZN => n6773);
   U12980 : NAND3_X1 port map( A1 => n6292, A2 => n6290, A3 => n6777, ZN => 
                           n6778);
   U12981 : AOI21_X1 port map( B1 => n6785, B2 => n6784, A => n6783, ZN => 
                           n6786);
   U12982 : INV_X1 port map( A => n7977, ZN => n7820);
   U12984 : INV_X1 port map( A => n7975, ZN => n7816);
   U12985 : NAND3_X1 port map( A1 => n7973, A2 => n7972, A3 => n7816, ZN => 
                           n6799);
   U12986 : NAND2_X1 port map( A1 => n6793, A2 => n6795, ZN => n6791);
   U12987 : NAND2_X1 port map( A1 => n6793, A2 => n6792, ZN => n6797);
   U12988 : OAI21_X1 port map( B1 => n6795, B2 => n6794, A => n6075, ZN => 
                           n6796);
   U12989 : AOI22_X1 port map( A1 => n6798, A2 => n6881, B1 => n6797, B2 => 
                           n6796, ZN => n7976);
   U12990 : INV_X1 port map( A => n7976, ZN => n7819);
   U12991 : NAND2_X1 port map( A1 => n7819, A2 => n7974, ZN => n7821);
   U12992 : XNOR2_X1 port map( A => n8913, B => n9140, ZN => n6800);
   U12993 : XNOR2_X1 port map( A => n8628, B => n6800, ZN => n6859);
   U12995 : AOI22_X1 port map( A1 => n7598, A2 => n7600, B1 => n25037, B2 => 
                           n7257, ZN => n6804);
   U12996 : NAND3_X1 port map( A1 => n7597, A2 => n7600, A3 => n7602, ZN => 
                           n6801);
   U12997 : AND2_X1 port map( A1 => n6802, A2 => n6801, ZN => n6803);
   U12998 : OAI21_X2 port map( B1 => n6804, B2 => n7597, A => n6803, ZN => 
                           n9141);
   U12999 : XNOR2_X1 port map( A => n9141, B => n2318, ZN => n6857);
   U13000 : NAND2_X1 port map( A1 => n7665, A2 => n8527, ZN => n6809);
   U13001 : NAND2_X1 port map( A1 => n6805, A2 => n7667, ZN => n6808);
   U13002 : NAND2_X1 port map( A1 => n7664, A2 => n8528, ZN => n6807);
   U13003 : NAND2_X1 port map( A1 => n6999, A2 => n6072, ZN => n6814);
   U13006 : NAND2_X1 port map( A1 => n6818, A2 => n6895, ZN => n6820);
   U13007 : AOI21_X1 port map( B1 => n6820, B2 => n6819, A => n313, ZN => n6821
                           );
   U13008 : INV_X1 port map( A => n7985, ZN => n7828);
   U13009 : NAND2_X1 port map( A1 => n6823, A2 => n6822, ZN => n6825);
   U13010 : AOI21_X1 port map( B1 => n6826, B2 => n6825, A => n6824, ZN => 
                           n6831);
   U13011 : INV_X1 port map( A => n7984, ZN => n7825);
   U13012 : MUX2_X1 port map( A => n6834, B => n6833, S => n7011, Z => n6837);
   U13013 : AND2_X1 port map( A1 => n7009, A2 => n7008, ZN => n6835);
   U13014 : OAI21_X1 port map( B1 => n6840, B2 => n6986, A => n6839, ZN => 
                           n6844);
   U13015 : NAND2_X1 port map( A1 => n6244, A2 => n6987, ZN => n6842);
   U13016 : AOI21_X1 port map( B1 => n6842, B2 => n6841, A => n6990, ZN => 
                           n6843);
   U13017 : NOR2_X1 port map( A1 => n6844, A2 => n6843, ZN => n7409);
   U13018 : INV_X1 port map( A => n7409, ZN => n7046);
   U13019 : NAND3_X1 port map( A1 => n7989, A2 => n7048, A3 => n7046, ZN => 
                           n6853);
   U13020 : NAND2_X1 port map( A1 => n6846, A2 => n6845, ZN => n6847);
   U13021 : OAI211_X1 port map( C1 => n7027, C2 => n7021, A => n6847, B => 
                           n7025, ZN => n6851);
   U13022 : OAI211_X1 port map( C1 => n250, C2 => n7027, A => n7028, B => n442,
                           ZN => n6850);
   U13023 : XNOR2_X1 port map( A => n8353, B => n8687, ZN => n6856);
   U13024 : XNOR2_X1 port map( A => n6857, B => n6856, ZN => n6858);
   U13025 : XNOR2_X1 port map( A => n6859, B => n6858, ZN => n9459);
   U13026 : NAND2_X1 port map( A1 => n9461, A2 => n9459, ZN => n9913);
   U13027 : NAND2_X1 port map( A1 => n9921, A2 => n9913, ZN => n7043);
   U13028 : NAND2_X1 port map( A1 => n6860, A2 => n7664, ZN => n6863);
   U13029 : NOR2_X1 port map( A1 => n7087, A2 => n7662, ZN => n6861);
   U13030 : AOI22_X1 port map( A1 => n6861, A2 => n8530, B1 => n269, B2 => 
                           n8531, ZN => n6862);
   U13031 : AOI21_X1 port map( B1 => n8317, B2 => n8315, A => n8314, ZN => 
                           n6866);
   U13032 : XNOR2_X1 port map( A => n8987, B => n9167, ZN => n8058);
   U13033 : NAND2_X1 port map( A1 => n6871, A2 => n6870, ZN => n6872);
   U13034 : AND2_X1 port map( A1 => n6873, A2 => n6872, ZN => n6880);
   U13035 : NAND2_X1 port map( A1 => n6875, A2 => n6874, ZN => n6877);
   U13036 : NAND2_X1 port map( A1 => n6882, A2 => n6881, ZN => n6888);
   U13037 : INV_X1 port map( A => n6883, ZN => n6887);
   U13038 : NAND2_X1 port map( A1 => n6885, A2 => n6884, ZN => n6886);
   U13039 : NAND2_X1 port map( A1 => n6895, A2 => n6890, ZN => n6891);
   U13040 : NAND2_X1 port map( A1 => n6892, A2 => n6891, ZN => n6898);
   U13041 : NOR2_X1 port map( A1 => n6895, A2 => n6894, ZN => n6896);
   U13042 : AOI21_X2 port map( B1 => n6897, B2 => n6898, A => n6896, ZN => 
                           n7657);
   U13043 : INV_X1 port map( A => n6899, ZN => n6901);
   U13044 : NAND2_X1 port map( A1 => n6901, A2 => n6900, ZN => n6908);
   U13045 : OAI21_X1 port map( B1 => n6905, B2 => n6904, A => n6903, ZN => 
                           n6907);
   U13046 : MUX2_X2 port map( A => n6908, B => n6907, S => n6906, Z => n7943);
   U13047 : NAND3_X1 port map( A1 => n6910, A2 => n6909, A3 => n6916, ZN => 
                           n6914);
   U13048 : NAND3_X1 port map( A1 => n6912, A2 => n24037, A3 => n6911, ZN => 
                           n6913);
   U13049 : NAND2_X1 port map( A1 => n6916, A2 => n6915, ZN => n6921);
   U13050 : NAND2_X1 port map( A1 => n6918, A2 => n24509, ZN => n6920);
   U13051 : NAND3_X1 port map( A1 => n7945, A2 => n7657, A3 => n7942, ZN => 
                           n6930);
   U13052 : AOI21_X1 port map( B1 => n6926, B2 => n6925, A => n6924, ZN => 
                           n6927);
   U13055 : INV_X1 port map( A => n6938, ZN => n6942);
   U13056 : NAND2_X1 port map( A1 => n6940, A2 => n6939, ZN => n6941);
   U13057 : NAND3_X1 port map( A1 => n6950, A2 => n6949, A3 => n6948, ZN => 
                           n6951);
   U13058 : OAI21_X1 port map( B1 => n6956, B2 => n24257, A => n6954, ZN => 
                           n6962);
   U13059 : OAI21_X1 port map( B1 => n3923, B2 => n6959, A => n6958, ZN => 
                           n6961);
   U13060 : INV_X1 port map( A => n6963, ZN => n6966);
   U13061 : AOI21_X1 port map( B1 => n6966, B2 => n6965, A => n6964, ZN => 
                           n6970);
   U13062 : NAND2_X1 port map( A1 => n6967, A2 => n443, ZN => n6968);
   U13064 : NOR2_X1 port map( A1 => n6971, A2 => n6977, ZN => n6973);
   U13065 : OAI21_X1 port map( B1 => n6973, B2 => n6974, A => n24579, ZN => 
                           n6981);
   U13066 : NAND2_X1 port map( A1 => n6976, A2 => n24395, ZN => n6978);
   U13067 : MUX2_X1 port map( A => n6979, B => n6978, S => n6977, Z => n6980);
   U13068 : INV_X1 port map( A => n7897, ZN => n6985);
   U13069 : NAND2_X1 port map( A1 => n6982, A2 => n7232, ZN => n6983);
   U13070 : NAND2_X1 port map( A1 => n6983, A2 => n24861, ZN => n6984);
   U13071 : XNOR2_X1 port map( A => n8499, B => n8088, ZN => n7040);
   U13072 : OAI21_X1 port map( B1 => n6838, B2 => n6986, A => n6989, ZN => 
                           n6995);
   U13073 : AOI21_X1 port map( B1 => n6988, B2 => n6987, A => n6990, ZN => 
                           n6994);
   U13074 : OAI21_X1 port map( B1 => n6244, B2 => n6990, A => n6989, ZN => 
                           n6992);
   U13075 : NAND2_X1 port map( A1 => n6992, A2 => n6991, ZN => n6993);
   U13076 : INV_X1 port map( A => n7961, ZN => n7070);
   U13077 : OAI21_X1 port map( B1 => n6368, B2 => n6996, A => n6367, ZN => 
                           n6998);
   U13078 : NAND2_X1 port map( A1 => n6998, A2 => n7002, ZN => n7001);
   U13079 : NAND2_X1 port map( A1 => n7070, A2 => n7962, ZN => n7069);
   U13080 : OAI21_X1 port map( B1 => n7009, B2 => n7008, A => n7007, ZN => 
                           n7010);
   U13081 : NAND2_X1 port map( A1 => n5992, A2 => n7013, ZN => n7016);
   U13082 : OAI21_X1 port map( B1 => n7033, B2 => n7035, A => n7032, ZN => 
                           n7034);
   U13083 : NAND2_X1 port map( A1 => n7036, A2 => n7961, ZN => n7038);
   U13084 : AND2_X1 port map( A1 => n7234, A2 => n7965, ZN => n7960);
   U13085 : NAND2_X1 port map( A1 => n7960, A2 => n7683, ZN => n7037);
   U13086 : OAI211_X2 port map( C1 => n7069, C2 => n7235, A => n7038, B => 
                           n7037, ZN => n8813);
   U13087 : XNOR2_X1 port map( A => n8813, B => n2772, ZN => n7039);
   U13088 : XNOR2_X1 port map( A => n7040, B => n7039, ZN => n7041);
   U13089 : AOI21_X1 port map( B1 => n7046, B2 => n7826, A => n7825, ZN => 
                           n7047);
   U13090 : XNOR2_X1 port map( A => n8812, B => n24056, ZN => n8459);
   U13091 : AOI21_X1 port map( B1 => n7517, B2 => n7516, A => n7972, ZN => 
                           n7051);
   U13092 : NAND2_X1 port map( A1 => n7816, A2 => n7974, ZN => n7049);
   U13093 : XNOR2_X1 port map( A => n8764, B => n8406, ZN => n7052);
   U13094 : XNOR2_X1 port map( A => n8459, B => n7052, ZN => n7063);
   U13095 : INV_X1 port map( A => n7800, ZN => n7054);
   U13096 : NAND2_X1 port map( A1 => n7801, A2 => n7798, ZN => n7434);
   U13097 : INV_X1 port map( A => n3118, ZN => n23448);
   U13098 : XNOR2_X1 port map( A => n8896, B => n23448, ZN => n7061);
   U13099 : AND2_X1 port map( A1 => n7412, A2 => n7358, ZN => n7499);
   U13100 : AOI22_X1 port map( A1 => n7499, A2 => n7991, B1 => n7992, B2 => 
                           n7415, ZN => n7056);
   U13101 : NAND3_X1 port map( A1 => n7992, A2 => n7413, A3 => n7412, ZN => 
                           n7055);
   U13102 : OAI211_X1 port map( C1 => n7414, C2 => n7992, A => n7056, B => 
                           n7055, ZN => n8285);
   U13103 : NAND2_X1 port map( A1 => n7813, A2 => n8219, ZN => n7059);
   U13104 : NAND3_X1 port map( A1 => n7813, A2 => n9068, A3 => n9066, ZN => 
                           n7058);
   U13105 : XNOR2_X1 port map( A => n8285, B => n9044, ZN => n7060);
   U13106 : XNOR2_X1 port map( A => n7061, B => n7060, ZN => n7062);
   U13107 : INV_X1 port map( A => n7183, ZN => n9951);
   U13108 : NOR2_X1 port map( A1 => n7421, A2 => n7474, ZN => n7064);
   U13109 : NAND2_X1 port map( A1 => n7423, A2 => n7477, ZN => n7067);
   U13110 : MUX2_X1 port map( A => n7067, B => n7066, S => n7476, Z => n7068);
   U13111 : OAI211_X1 port map( C1 => n7071, C2 => n7070, A => n7485, B => 
                           n7069, ZN => n7072);
   U13112 : OR2_X1 port map( A1 => n7078, A2 => n7674, ZN => n7076);
   U13113 : OAI21_X1 port map( B1 => n7076, B2 => n7224, A => n7075, ZN => 
                           n7077);
   U13114 : NAND3_X1 port map( A1 => n434, A2 => n7677, A3 => n7078, ZN => 
                           n7079);
   U13115 : INV_X1 port map( A => n8452, ZN => n8820);
   U13116 : INV_X1 port map( A => n7947, ZN => n7946);
   U13117 : NAND2_X1 port map( A1 => n7946, A2 => n7942, ZN => n7081);
   U13118 : NOR2_X1 port map( A1 => n7945, A2 => n7657, ZN => n7080);
   U13119 : XNOR2_X1 port map( A => n8820, B => n8787, ZN => n7082);
   U13120 : XNOR2_X1 port map( A => n7083, B => n7082, ZN => n7095);
   U13121 : NAND2_X1 port map( A1 => n8317, A2 => n8316, ZN => n7149);
   U13122 : NAND2_X1 port map( A1 => n8315, A2 => n8314, ZN => n7084);
   U13123 : NAND3_X1 port map( A1 => n7149, A2 => n7085, A3 => n7084, ZN => 
                           n7086);
   U13124 : OAI211_X1 port map( C1 => n7149, C2 => n7217, A => n7086, B => 
                           n8319, ZN => n9073);
   U13125 : NAND3_X1 port map( A1 => n8530, A2 => n7667, A3 => n8528, ZN => 
                           n7091);
   U13126 : NAND3_X1 port map( A1 => n7665, A2 => n7667, A3 => n269, ZN => 
                           n7090);
   U13128 : NAND3_X1 port map( A1 => n7664, A2 => n7666, A3 => n7662, ZN => 
                           n7088);
   U13129 : NAND4_X2 port map( A1 => n7088, A2 => n7091, A3 => n7090, A4 => 
                           n7089, ZN => n8651);
   U13130 : XNOR2_X1 port map( A => n9073, B => n8651, ZN => n7093);
   U13131 : INV_X1 port map( A => n21204, ZN => n22150);
   U13132 : XNOR2_X1 port map( A => n8412, B => n22150, ZN => n7092);
   U13133 : XNOR2_X1 port map( A => n7093, B => n7092, ZN => n7094);
   U13134 : XNOR2_X1 port map( A => n7095, B => n7094, ZN => n9950);
   U13135 : NAND2_X1 port map( A1 => n9951, A2 => n9950, ZN => n9387);
   U13137 : NOR2_X1 port map( A1 => n7098, A2 => n7097, ZN => n7099);
   U13138 : NAND4_X1 port map( A1 => n7105, A2 => n7347, A3 => n7349, A4 => 
                           n7104, ZN => n7106);
   U13139 : XNOR2_X1 port map( A => n8333, B => n8280, ZN => n7113);
   U13140 : NAND2_X1 port map( A1 => n7526, A2 => n7771, ZN => n7110);
   U13141 : NAND2_X1 port map( A1 => n7284, A2 => n7527, ZN => n7109);
   U13142 : INV_X1 port map( A => n7768, ZN => n7288);
   U13143 : MUX2_X1 port map( A => n7110, B => n7109, S => n7288, Z => n7112);
   U13145 : AOI22_X1 port map( A1 => n7522, A2 => n23, B1 => n7525, B2 => n7767
                           , ZN => n7111);
   U13147 : XNOR2_X1 port map( A => n8891, B => n8807, ZN => n8444);
   U13148 : XNOR2_X1 port map( A => n8444, B => n7113, ZN => n7120);
   U13149 : NAND2_X1 port map( A1 => n7754, A2 => n7292, ZN => n8006);
   U13150 : NAND2_X1 port map( A1 => n7760, A2 => n7651, ZN => n7115);
   U13151 : NOR2_X1 port map( A1 => n7761, A2 => n7646, ZN => n7116);
   U13152 : OAI21_X1 port map( B1 => n7391, B2 => n7116, A => n7305, ZN => 
                           n7117);
   U13153 : XNOR2_X1 port map( A => n8400, B => n923, ZN => n7118);
   U13154 : XNOR2_X1 port map( A => n25020, B => n7118, ZN => n7119);
   U13155 : OAI21_X1 port map( B1 => n7592, B2 => n7590, A => n268, ZN => n7122
                           );
   U13156 : NAND3_X1 port map( A1 => n7462, A2 => n2035, A3 => n5971, ZN => 
                           n7121);
   U13157 : INV_X1 port map( A => n7882, ZN => n7126);
   U13159 : INV_X1 port map( A => n7313, ZN => n7123);
   U13160 : INV_X1 port map( A => n7585, ZN => n7125);
   U13161 : NAND3_X1 port map( A1 => n7126, A2 => n7125, A3 => n7582, ZN => 
                           n7127);
   U13162 : INV_X1 port map( A => n7604, ZN => n7128);
   U13163 : NOR2_X1 port map( A1 => n7604, A2 => n7323, ZN => n7129);
   U13164 : INV_X1 port map( A => n7579, ZN => n7318);
   U13165 : NAND2_X1 port map( A1 => n7577, A2 => n7318, ZN => n7320);
   U13166 : NAND3_X1 port map( A1 => n7577, A2 => n4136, A3 => n7576, ZN => 
                           n7130);
   U13169 : NAND2_X1 port map( A1 => n7600, A2 => n7597, ZN => n7132);
   U13171 : NAND2_X1 port map( A1 => n7596, A2 => n7255, ZN => n7133);
   U13172 : NAND3_X1 port map( A1 => n25037, A2 => n24772, A3 => n7135, ZN => 
                           n7138);
   U13173 : NAND3_X1 port map( A1 => n7255, A2 => n7600, A3 => n7257, ZN => 
                           n7137);
   U13174 : XNOR2_X1 port map( A => n8647, B => n8341, ZN => n8387);
   U13175 : NAND2_X1 port map( A1 => n248, A2 => n7230, ZN => n7139);
   U13176 : NAND2_X1 port map( A1 => n7140, A2 => n24861, ZN => n7142);
   U13177 : NOR2_X1 port map( A1 => n7230, A2 => n7232, ZN => n7141);
   U13178 : INV_X1 port map( A => n8168, ZN => n8270);
   U13179 : XNOR2_X1 port map( A => n8270, B => n3089, ZN => n7144);
   U13180 : XNOR2_X1 port map( A => n8387, B => n7144, ZN => n7145);
   U13181 : XNOR2_X1 port map( A => n7146, B => n7145, ZN => n9134);
   U13182 : INV_X1 port map( A => n9134, ZN => n9389);
   U13183 : NAND3_X1 port map( A1 => n7699, A2 => n7688, A3 => n8315, ZN => 
                           n7150);
   U13186 : XNOR2_X1 port map( A => n24547, B => n8353, ZN => n8421);
   U13187 : INV_X1 port map( A => n7909, ZN => n7625);
   U13188 : NAND2_X1 port map( A1 => n7625, A2 => n7628, ZN => n7154);
   U13189 : NAND2_X1 port map( A1 => n7365, A2 => n7909, ZN => n7153);
   U13190 : NAND3_X1 port map( A1 => n7154, A2 => n7153, A3 => n7364, ZN => 
                           n7158);
   U13194 : XNOR2_X1 port map( A => n7161, B => n9082, ZN => n8689);
   U13195 : INV_X1 port map( A => n8689, ZN => n7162);
   U13196 : XNOR2_X1 port map( A => n7162, B => n8421, ZN => n7182);
   U13197 : NOR2_X1 port map( A1 => n7163, A2 => n7932, ZN => n7164);
   U13198 : INV_X1 port map( A => n7924, ZN => n7261);
   U13199 : AOI22_X1 port map( A1 => n7164, A2 => n7261, B1 => n7445, B2 => 
                           n7932, ZN => n7165);
   U13200 : NAND2_X1 port map( A1 => n7167, A2 => n7801, ZN => n7169);
   U13201 : OAI21_X1 port map( B1 => n7169, B2 => n7800, A => n7168, ZN => 
                           n7171);
   U13202 : AOI21_X1 port map( B1 => n7434, B2 => n7795, A => n7432, ZN => 
                           n7170);
   U13203 : OR2_X1 port map( A1 => n7171, A2 => n7170, ZN => n8237);
   U13204 : XNOR2_X1 port map( A => n8428, B => n8237, ZN => n7180);
   U13205 : NAND2_X1 port map( A1 => n7782, A2 => n7418, ZN => n7172);
   U13206 : NAND2_X1 port map( A1 => n7172, A2 => n2620, ZN => n7173);
   U13207 : NAND2_X1 port map( A1 => n7173, A2 => n7781, ZN => n7178);
   U13208 : NAND3_X1 port map( A1 => n7419, A2 => n7174, A3 => n7787, ZN => 
                           n7177);
   U13209 : XNOR2_X1 port map( A => n8917, B => n2120, ZN => n7179);
   U13210 : XNOR2_X1 port map( A => n7180, B => n7179, ZN => n7181);
   U13211 : XNOR2_X1 port map( A => n7182, B => n7181, ZN => n9269);
   U13212 : OR2_X1 port map( A1 => n9133, A2 => n9951, ZN => n7210);
   U13213 : NAND2_X1 port map( A1 => n7184, A2 => n4754, ZN => n7185);
   U13214 : OAI21_X1 port map( B1 => n24072, B2 => n7857, A => n7562, ZN => 
                           n7245);
   U13215 : INV_X1 port map( A => n7246, ZN => n7565);
   U13216 : NAND2_X1 port map( A1 => n7565, A2 => n7563, ZN => n7186);
   U13219 : NAND2_X1 port map( A1 => n24578, A2 => n7732, ZN => n7187);
   U13220 : XNOR2_X1 port map( A => n9107, B => n8909, ZN => n7195);
   U13221 : NAND3_X1 port map( A1 => n3570, A2 => n7867, A3 => n7865, ZN => 
                           n7190);
   U13222 : NAND3_X1 port map( A1 => n7860, A2 => n7867, A3 => n7862, ZN => 
                           n7189);
   U13223 : NAND2_X1 port map( A1 => n7271, A2 => n4536, ZN => n7188);
   U13224 : NAND2_X1 port map( A1 => n7843, A2 => n24577, ZN => n7191);
   U13225 : NAND2_X1 port map( A1 => n7719, A2 => n7191, ZN => n7192);
   U13226 : NAND2_X1 port map( A1 => n7843, A2 => n8368, ZN => n7716);
   U13227 : OAI21_X1 port map( B1 => n7193, B2 => n7843, A => n7716, ZN => 
                           n7194);
   U13228 : XNOR2_X1 port map( A => n8772, B => n9059, ZN => n8696);
   U13229 : XNOR2_X1 port map( A => n8696, B => n7195, ZN => n7207);
   U13230 : OR2_X1 port map( A1 => n9067, A2 => n7057, ZN => n7430);
   U13231 : OAI21_X1 port map( B1 => n7812, B2 => n7809, A => n7430, ZN => 
                           n7198);
   U13232 : INV_X1 port map( A => n7057, ZN => n7810);
   U13233 : NAND2_X1 port map( A1 => n7196, A2 => n7810, ZN => n7197);
   U13235 : INV_X1 port map( A => n8361, ZN => n7200);
   U13236 : XNOR2_X1 port map( A => n8633, B => n7200, ZN => n8395);
   U13237 : INV_X1 port map( A => n8395, ZN => n7205);
   U13238 : NAND2_X1 port map( A1 => n7615, A2 => n7380, ZN => n7620);
   U13239 : XNOR2_X1 port map( A => n7205, B => n7204, ZN => n7206);
   U13240 : NAND2_X1 port map( A1 => n9134, A2 => n9388, ZN => n9132);
   U13241 : OAI21_X1 port map( B1 => n9949, B2 => n9388, A => n9132, ZN => 
                           n7208);
   U13242 : NAND2_X1 port map( A1 => n7208, A2 => n9959, ZN => n7209);
   U13243 : NOR2_X1 port map( A1 => n7666, A2 => n8527, ZN => n7212);
   U13244 : INV_X1 port map( A => n8533, ZN => n7213);
   U13246 : OAI21_X1 port map( B1 => n8315, B2 => n7217, A => n8317, ZN => 
                           n7218);
   U13247 : OAI21_X1 port map( B1 => n7698, B2 => n8317, A => n7218, ZN => 
                           n7219);
   U13248 : XNOR2_X1 port map( A => n24946, B => n8172, ZN => n7448);
   U13249 : OAI21_X1 port map( B1 => n7423, B2 => n4144, A => n7220, ZN => 
                           n7223);
   U13250 : INV_X1 port map( A => n7674, ZN => n7225);
   U13251 : XNOR2_X1 port map( A => n8491, B => n9159, ZN => n8947);
   U13252 : XNOR2_X1 port map( A => n8947, B => n7448, ZN => n7241);
   U13253 : INV_X1 port map( A => n7230, ZN => n7898);
   U13254 : XNOR2_X1 port map( A => n8867, B => n8612, ZN => n7239);
   U13255 : XNOR2_X1 port map( A => n8980, B => n1767, ZN => n7238);
   U13256 : XNOR2_X1 port map( A => n7239, B => n7238, ZN => n7240);
   U13257 : AOI21_X1 port map( B1 => n7773, B2 => n7769, A => n7776, ZN => 
                           n7244);
   U13258 : NAND2_X1 port map( A1 => n7768, A2 => n7767, ZN => n7242);
   U13259 : AOI21_X1 port map( B1 => n7242, B2 => n7527, A => n7526, ZN => 
                           n7243);
   U13260 : NAND2_X1 port map( A1 => n7245, A2 => n7853, ZN => n7249);
   U13261 : INV_X1 port map( A => n7850, ZN => n7725);
   U13262 : AOI21_X1 port map( B1 => n7725, B2 => n7721, A => n7857, ZN => 
                           n7247);
   U13263 : XNOR2_X1 port map( A => n8460, B => n8501, ZN => n8703);
   U13264 : NAND2_X1 port map( A1 => n8511, A2 => n7350, ZN => n7252);
   U13265 : NAND2_X1 port map( A1 => n7255, A2 => n7600, ZN => n7344);
   U13266 : NAND2_X1 port map( A1 => n7595, A2 => n7257, ZN => n7345);
   U13267 : INV_X1 port map( A => n7597, ZN => n7256);
   U13269 : XNOR2_X1 port map( A => n8542, B => n8345, ZN => n7471);
   U13270 : NAND2_X1 port map( A1 => n7444, A2 => n7932, ZN => n7263);
   U13271 : AOI21_X1 port map( B1 => n7445, B2 => n7263, A => n7923, ZN => 
                           n7264);
   U13272 : XNOR2_X1 port map( A => n8899, B => n20995, ZN => n7276);
   U13273 : INV_X1 port map( A => n8368, ZN => n7714);
   U13274 : NAND2_X1 port map( A1 => n7714, A2 => n7843, ZN => n7267);
   U13275 : INV_X1 port map( A => n7713, ZN => n7561);
   U13276 : AOI21_X1 port map( B1 => n7267, B2 => n7266, A => n7561, ZN => 
                           n7270);
   U13277 : AOI21_X1 port map( B1 => n7268, B2 => n8370, A => n7714, ZN => 
                           n7269);
   U13278 : NAND2_X1 port map( A1 => n7553, A2 => n7865, ZN => n7275);
   U13279 : NAND2_X1 port map( A1 => n7868, A2 => n24576, ZN => n7274);
   U13280 : NAND3_X1 port map( A1 => n7863, A2 => n24576, A3 => n7707, ZN => 
                           n7273);
   U13281 : NAND2_X1 port map( A1 => n7271, A2 => n7865, ZN => n7272);
   U13282 : XNOR2_X1 port map( A => n8989, B => n8875, ZN => n8112);
   U13283 : NAND2_X1 port map( A1 => n7279, A2 => n7350, ZN => n7280);
   U13284 : NAND3_X1 port map( A1 => n7347, A2 => n5468, A3 => n7351, ZN => 
                           n7282);
   U13285 : NAND3_X1 port map( A1 => n8511, A2 => n5468, A3 => n7349, ZN => 
                           n7281);
   U13286 : XNOR2_X1 port map( A => n9139, B => n8952, ZN => n7291);
   U13287 : INV_X1 port map( A => n7776, ZN => n7283);
   U13288 : AOI21_X1 port map( B1 => n7283, B2 => n25252, A => n7527, ZN => 
                           n7289);
   U13289 : NAND3_X1 port map( A1 => n23, A2 => n7776, A3 => n7284, ZN => n7286
                           );
   U13290 : XNOR2_X1 port map( A => n8798, B => n2743, ZN => n7290);
   U13291 : XNOR2_X1 port map( A => n7291, B => n7290, ZN => n7311);
   U13292 : INV_X1 port map( A => n7293, ZN => n7297);
   U13293 : INV_X1 port map( A => n8014, ZN => n7295);
   U13294 : NAND2_X1 port map( A1 => n7295, A2 => n8015, ZN => n7296);
   U13295 : NAND2_X1 port map( A1 => n8014, A2 => n8016, ZN => n7298);
   U13296 : NAND2_X1 port map( A1 => n7299, A2 => n7298, ZN => n7300);
   U13298 : XNOR2_X1 port map( A => n8147, B => n8132, ZN => n8734);
   U13299 : OAI21_X1 port map( B1 => n7385, B2 => n7617, A => n7380, ZN => 
                           n7304);
   U13300 : NAND3_X1 port map( A1 => n1895, A2 => n7619, A3 => n7618, ZN => 
                           n7302);
   U13301 : NAND2_X1 port map( A1 => n7390, A2 => n7760, ZN => n7306);
   U13302 : NAND3_X1 port map( A1 => n7760, A2 => n7307, A3 => n7648, ZN => 
                           n7308);
   U13304 : XNOR2_X1 port map( A => n8799, B => n8916, ZN => n8329);
   U13307 : NOR2_X1 port map( A1 => n7575, A2 => n7580, ZN => n7321);
   U13308 : XNOR2_X1 port map( A => n8853, B => n8959, ZN => n8363);
   U13309 : INV_X1 port map( A => n8363, ZN => n7334);
   U13310 : INV_X1 port map( A => n7323, ZN => n7605);
   U13311 : AND2_X1 port map( A1 => n7898, A2 => n248, ZN => n7328);
   U13312 : NAND2_X1 port map( A1 => n7328, A2 => n3469, ZN => n7333);
   U13313 : NAND2_X1 port map( A1 => n7329, A2 => n24103, ZN => n7331);
   U13314 : NAND4_X2 port map( A1 => n7332, A2 => n7333, A3 => n7331, A4 => 
                           n7330, ZN => n8962);
   U13315 : XNOR2_X1 port map( A => n8771, B => n8962, ZN => n8192);
   U13316 : XNOR2_X1 port map( A => n7334, B => n8192, ZN => n7356);
   U13317 : NAND2_X1 port map( A1 => n7335, A2 => n7461, ZN => n7463);
   U13318 : NAND2_X1 port map( A1 => n7463, A2 => n2035, ZN => n7336);
   U13319 : NAND2_X1 port map( A1 => n7337, A2 => n7336, ZN => n7340);
   U13320 : NAND2_X1 port map( A1 => n5737, A2 => n7338, ZN => n7339);
   U13321 : NAND2_X1 port map( A1 => n7340, A2 => n7339, ZN => n8360);
   U13322 : OAI211_X1 port map( C1 => n7600, C2 => n7597, A => n25037, B => 
                           n7341, ZN => n7343);
   U13323 : XNOR2_X1 port map( A => n8964, B => n8360, ZN => n7518);
   U13324 : OAI211_X1 port map( C1 => n7349, C2 => n7348, A => n7347, B => 
                           n7346, ZN => n7353);
   U13325 : INV_X1 port map( A => n7350, ZN => n8509);
   U13326 : OAI211_X1 port map( C1 => n8508, C2 => n8511, A => n7353, B => 
                           n7352, ZN => n8638);
   U13327 : XNOR2_X1 port map( A => n8638, B => n187, ZN => n7354);
   U13328 : XNOR2_X1 port map( A => n7518, B => n7354, ZN => n7355);
   U13329 : AND2_X1 port map( A1 => n7358, A2 => n7413, ZN => n7359);
   U13330 : AOI21_X1 port map( B1 => n7994, B2 => n7360, A => n3549, ZN => 
                           n7361);
   U13331 : NOR2_X2 port map( A1 => n7362, A2 => n7361, ZN => n8313);
   U13332 : NAND2_X1 port map( A1 => n7363, A2 => n7364, ZN => n7369);
   U13333 : NAND3_X1 port map( A1 => n7909, A2 => n7911, A3 => n7628, ZN => 
                           n7368);
   U13334 : NAND3_X1 port map( A1 => n7913, A2 => n7910, A3 => n7908, ZN => 
                           n7367);
   U13335 : NAND3_X1 port map( A1 => n7913, A2 => n7365, A3 => n7629, ZN => 
                           n7366);
   U13336 : INV_X1 port map( A => n7923, ZN => n7370);
   U13337 : NAND2_X1 port map( A1 => n7370, A2 => n7163, ZN => n7375);
   U13338 : NAND2_X1 port map( A1 => n7372, A2 => n7923, ZN => n7371);
   U13339 : OAI211_X1 port map( C1 => n7372, C2 => n5607, A => n7371, B => 
                           n7445, ZN => n7374);
   U13341 : NAND2_X1 port map( A1 => n5595, A2 => n7640, ZN => n7378);
   U13342 : NAND2_X1 port map( A1 => n7734, A2 => n7733, ZN => n7376);
   U13343 : NAND3_X1 port map( A1 => n7641, A2 => n24578, A3 => n7642, ZN => 
                           n7377);
   U13344 : XNOR2_X1 port map( A => n9182, B => n8517, ZN => n8940);
   U13345 : XNOR2_X1 port map( A => n8940, B => n7379, ZN => n7402);
   U13348 : NAND3_X1 port map( A1 => n7622, A2 => n7385, A3 => n7384, ZN => 
                           n7388);
   U13349 : NAND3_X1 port map( A1 => n7617, A2 => n7386, A3 => n7615, ZN => 
                           n7387);
   U13350 : NAND3_X2 port map( A1 => n7389, A2 => n7388, A3 => n7387, ZN => 
                           n8786);
   U13351 : NAND2_X1 port map( A1 => n7391, A2 => n7648, ZN => n7394);
   U13352 : OAI211_X1 port map( C1 => n7647, C2 => n7760, A => n7392, B => 
                           n7646, ZN => n7393);
   U13353 : XNOR2_X1 port map( A => n8375, B => n8786, ZN => n7400);
   U13354 : NAND3_X1 port map( A1 => n7634, A2 => n3347, A3 => n7917, ZN => 
                           n7397);
   U13355 : NAND3_X1 port map( A1 => n7449, A2 => n25253, A3 => n7918, ZN => 
                           n7395);
   U13356 : XNOR2_X1 port map( A => n8860, B => n21169, ZN => n7399);
   U13357 : XNOR2_X1 port map( A => n7400, B => n7399, ZN => n7401);
   U13358 : XNOR2_X1 port map( A => n7402, B => n7401, ZN => n10129);
   U13359 : NOR2_X1 port map( A1 => n7819, A2 => n7974, ZN => n7403);
   U13360 : AOI22_X1 port map( A1 => n7404, A2 => n7816, B1 => n7403, B2 => 
                           n7820, ZN => n7408);
   U13361 : NAND2_X1 port map( A1 => n7975, A2 => n7974, ZN => n7406);
   U13362 : NAND2_X1 port map( A1 => n7829, A2 => n7983, ZN => n7987);
   U13363 : OAI21_X1 port map( B1 => n7983, B2 => n7982, A => n7987, ZN => 
                           n7410);
   U13364 : NAND2_X1 port map( A1 => n7410, A2 => n7985, ZN => n7411);
   U13365 : XNOR2_X1 port map( A => n9015, B => n8476, ZN => n8117);
   U13366 : OR2_X1 port map( A1 => n7413, A2 => n7412, ZN => n7502);
   U13367 : OAI211_X1 port map( C1 => n7990, C2 => n7993, A => n7502, B => 
                           n3549, ZN => n7417);
   U13368 : INV_X1 port map( A => n7993, ZN => n7500);
   U13369 : NAND3_X1 port map( A1 => n7500, A2 => n7415, A3 => n7998, ZN => 
                           n7416);
   U13370 : INV_X1 port map( A => n7418, ZN => n7784);
   U13371 : NOR2_X1 port map( A1 => n7788, A2 => n7418, ZN => n7420);
   U13372 : XNOR2_X1 port map( A => n8119, B => n8477, ZN => n8937);
   U13373 : INV_X1 port map( A => n8937, ZN => n8672);
   U13374 : XNOR2_X1 port map( A => n8672, B => n8117, ZN => n7436);
   U13375 : INV_X1 port map( A => n7421, ZN => n7422);
   U13376 : OAI21_X1 port map( B1 => n7422, B2 => n7476, A => n7423, ZN => 
                           n7426);
   U13377 : OAI211_X1 port map( C1 => n7954, C2 => n7426, A => n7425, B => 
                           n7424, ZN => n8296);
   U13378 : INV_X1 port map( A => n3131, ZN => n23347);
   U13379 : XNOR2_X1 port map( A => n8296, B => n23347, ZN => n7435);
   U13380 : NAND2_X1 port map( A1 => n7809, A2 => n7813, ZN => n7429);
   U13381 : MUX2_X1 port map( A => n7429, B => n7428, S => n7812, Z => n7431);
   U13382 : INV_X1 port map( A => n7809, ZN => n9071);
   U13383 : NAND3_X1 port map( A1 => n7795, A2 => n7432, A3 => n7799, ZN => 
                           n7433);
   U13384 : XNOR2_X1 port map( A => n8754, B => n8339, ZN => n7552);
   U13385 : MUX2_X1 port map( A => n7781, B => n7782, S => n7789, Z => n7442);
   U13386 : MUX2_X1 port map( A => n7443, B => n7442, S => n7784, Z => n8780);
   U13387 : MUX2_X1 port map( A => n7445, B => n7444, S => n7932, Z => n7447);
   U13388 : XNOR2_X1 port map( A => n8780, B => n8492, ZN => n8279);
   U13389 : XNOR2_X1 port map( A => n7448, B => n8279, ZN => n7454);
   U13390 : INV_X1 port map( A => n9034, ZN => n7451);
   U13391 : XNOR2_X1 port map( A => n7451, B => n8613, ZN => n8399);
   U13392 : XNOR2_X1 port map( A => n9155, B => n3125, ZN => n7452);
   U13393 : XNOR2_X1 port map( A => n8399, B => n7452, ZN => n7453);
   U13394 : AOI21_X1 port map( B1 => n7322, B2 => n7890, A => n7605, ZN => 
                           n7456);
   U13395 : INV_X1 port map( A => n7577, ZN => n7574);
   U13396 : AOI21_X1 port map( B1 => n7574, B2 => n7579, A => n7576, ZN => 
                           n7458);
   U13397 : XNOR2_X1 port map( A => n8499, B => n1789, ZN => n7459);
   U13398 : XNOR2_X1 port map( A => n8287, B => n7459, ZN => n7473);
   U13399 : OAI211_X1 port map( C1 => n7462, C2 => n7592, A => n7591, B => 
                           n7461, ZN => n7466);
   U13400 : INV_X1 port map( A => n7463, ZN => n7465);
   U13401 : AOI22_X1 port map( A1 => n7467, A2 => n7466, B1 => n7465, B2 => 
                           n7464, ZN => n8620);
   U13402 : INV_X1 port map( A => n8620, ZN => n8988);
   U13403 : INV_X1 port map( A => n7584, ZN => n7884);
   U13404 : NAND2_X1 port map( A1 => n7581, A2 => n7882, ZN => n7468);
   U13405 : NAND2_X1 port map( A1 => n7468, A2 => n7585, ZN => n7469);
   U13407 : XNOR2_X1 port map( A => n8988, B => n25228, ZN => n8405);
   U13408 : XNOR2_X1 port map( A => n8405, B => n7471, ZN => n7472);
   U13409 : NOR2_X1 port map( A1 => n7475, A2 => n7474, ZN => n7479);
   U13410 : NAND2_X1 port map( A1 => n7477, A2 => n7476, ZN => n7478);
   U13411 : INV_X1 port map( A => n9141, ZN => n7480);
   U13412 : XNOR2_X1 port map( A => n7480, B => n8238, ZN => n8467);
   U13413 : NAND3_X1 port map( A1 => n7481, A2 => n7577, A3 => n7579, ZN => 
                           n7482);
   U13414 : AND2_X1 port map( A1 => n7483, A2 => n7482, ZN => n7484);
   U13415 : XNOR2_X1 port map( A => n8795, B => n8147, ZN => n8580);
   U13416 : XNOR2_X1 port map( A => n8467, B => n8580, ZN => n7497);
   U13417 : NAND2_X1 port map( A1 => n7485, A2 => n7962, ZN => n7488);
   U13418 : INV_X1 port map( A => n7966, ZN => n7486);
   U13419 : XNOR2_X1 port map( A => n9081, B => n8799, ZN => n7495);
   U13420 : INV_X1 port map( A => n7942, ZN => n7490);
   U13421 : NAND3_X1 port map( A1 => n7943, A2 => n7490, A3 => n7947, ZN => 
                           n7492);
   U13422 : NAND2_X1 port map( A1 => n24475, A2 => n7657, ZN => n7491);
   U13423 : XNOR2_X1 port map( A => n7495, B => n7494, ZN => n7496);
   U13424 : XNOR2_X1 port map( A => n8484, B => n21623, ZN => n7511);
   U13425 : INV_X1 port map( A => n7502, ZN => n7503);
   U13426 : OAI21_X1 port map( B1 => n7991, B2 => n7993, A => n7503, ZN => 
                           n7504);
   U13427 : NAND2_X1 port map( A1 => n7505, A2 => n7504, ZN => n8093);
   U13428 : INV_X1 port map( A => n8093, ZN => n8485);
   U13429 : NOR2_X1 port map( A1 => n25251, A2 => n7674, ZN => n7508);
   U13430 : XNOR2_X1 port map( A => n8485, B => n8769, ZN => n8265);
   U13431 : XNOR2_X1 port map( A => n7511, B => n8265, ZN => n7520);
   U13432 : OAI211_X1 port map( C1 => n7985, C2 => n7829, A => n7989, B => 
                           n7982, ZN => n7512);
   U13433 : OAI211_X1 port map( C1 => n7977, C2 => n7514, A => n7975, B => 
                           n7973, ZN => n7515);
   U13434 : OAI211_X1 port map( C1 => n7517, C2 => n7977, A => n7516, B => 
                           n7515, ZN => n8639);
   U13435 : XNOR2_X1 port map( A => n9058, B => n8639, ZN => n8391);
   U13436 : XNOR2_X1 port map( A => n7518, B => n8391, ZN => n7519);
   U13437 : XNOR2_X1 port map( A => n7520, B => n7519, ZN => n8141);
   U13438 : OAI22_X1 port map( A1 => n9962, A2 => n9468, B1 => n9964, B2 => 
                           n9961, ZN => n8140);
   U13439 : INV_X1 port map( A => n7527, ZN => n7521);
   U13440 : NAND2_X1 port map( A1 => n3013, A2 => n7521, ZN => n7524);
   U13442 : XNOR2_X1 port map( A => n8790, B => n8506, ZN => n8291);
   U13443 : XNOR2_X1 port map( A => n9175, B => n8786, ZN => n7534);
   U13444 : XNOR2_X1 port map( A => n7534, B => n8291, ZN => n7550);
   U13445 : NOR2_X1 port map( A1 => n8014, A2 => n8012, ZN => n7536);
   U13446 : NAND3_X1 port map( A1 => n8014, A2 => n8016, A3 => n25451, ZN => 
                           n7539);
   U13447 : NAND3_X1 port map( A1 => n7543, A2 => n7542, A3 => n7758, ZN => 
                           n7545);
   U13449 : XNOR2_X1 port map( A => n9007, B => n9075, ZN => n8411);
   U13450 : XNOR2_X1 port map( A => n8375, B => n763, ZN => n7548);
   U13451 : XNOR2_X1 port map( A => n8411, B => n7548, ZN => n7549);
   U13452 : XNOR2_X1 port map( A => n9194, B => n16574, ZN => n7551);
   U13453 : XNOR2_X1 port map( A => n7552, B => n7551, ZN => n7571);
   U13454 : AOI22_X1 port map( A1 => n7710, A2 => n24576, B1 => n7553, B2 => 
                           n7707, ZN => n7556);
   U13455 : NAND2_X1 port map( A1 => n7867, A2 => n7864, ZN => n7554);
   U13457 : INV_X1 port map( A => n7843, ZN => n7718);
   U13458 : INV_X1 port map( A => n8370, ZN => n7715);
   U13459 : OAI211_X1 port map( C1 => n8371, C2 => n7843, A => n7558, B => 
                           n7714, ZN => n7559);
   U13460 : XNOR2_X1 port map( A => n9016, B => n8880, ZN => n8385);
   U13461 : INV_X1 port map( A => n7857, ZN => n7722);
   U13462 : NAND3_X1 port map( A1 => n7565, A2 => n7564, A3 => n7563, ZN => 
                           n7724);
   U13463 : INV_X1 port map( A => n7730, ZN => n7568);
   U13464 : XNOR2_X1 port map( A => n8478, B => n9191, ZN => n8269);
   U13465 : XNOR2_X1 port map( A => n8269, B => n8385, ZN => n7570);
   U13466 : NAND3_X1 port map( A1 => n7887, A2 => n7585, A3 => n7883, ZN => 
                           n7586);
   U13467 : XNOR2_X1 port map( A => n7594, B => n8889, ZN => n7614);
   U13469 : NOR2_X1 port map( A1 => n7600, A2 => n7597, ZN => n7599);
   U13470 : XNOR2_X1 port map( A => n8280, B => n8446, ZN => n7612);
   U13471 : NAND2_X1 port map( A1 => n7890, A2 => n7604, ZN => n7892);
   U13472 : AND2_X1 port map( A1 => n7605, A2 => n7604, ZN => n7607);
   U13474 : XNOR2_X1 port map( A => n8682, B => n1810, ZN => n7611);
   U13475 : XNOR2_X1 port map( A => n7612, B => n7611, ZN => n7613);
   U13476 : OAI22_X1 port map( A1 => n7622, A2 => n7621, B1 => n7620, B2 => 
                           n7619, ZN => n7623);
   U13477 : XNOR2_X1 port map( A => n8285, B => n8458, ZN => n8230);
   U13478 : AOI21_X1 port map( B1 => n7627, B2 => n7626, A => n7625, ZN => 
                           n7632);
   U13479 : AOI21_X1 port map( B1 => n7630, B2 => n7629, A => n7628, ZN => 
                           n7631);
   U13481 : XNOR2_X1 port map( A => n8899, B => n8706, ZN => n7633);
   U13482 : XNOR2_X1 port map( A => n8230, B => n7633, ZN => n7655);
   U13483 : AOI21_X1 port map( B1 => n7634, B2 => n3348, A => n25253, ZN => 
                           n7639);
   U13484 : NAND2_X1 port map( A1 => n7636, A2 => n7635, ZN => n7637);
   U13485 : NAND3_X1 port map( A1 => n7731, A2 => n7642, A3 => n7732, ZN => 
                           n7643);
   U13486 : XNOR2_X1 port map( A => n8760, B => n8898, ZN => n7653);
   U13487 : NAND2_X1 port map( A1 => n7760, A2 => n7647, ZN => n7650);
   U13488 : INV_X1 port map( A => n1754, ZN => n23225);
   U13489 : XNOR2_X1 port map( A => n9043, B => n23225, ZN => n7652);
   U13490 : XNOR2_X1 port map( A => n7653, B => n7652, ZN => n7654);
   U13491 : NOR2_X1 port map( A1 => n24474, A2 => n7945, ZN => n7661);
   U13492 : INV_X1 port map( A => n7943, ZN => n7656);
   U13493 : NAND2_X1 port map( A1 => n7943, A2 => n7942, ZN => n7659);
   U13494 : XNOR2_X1 port map( A => n8721, B => n8673, ZN => n7681);
   U13495 : OAI211_X1 port map( C1 => n7675, C2 => n7674, A => n7673, B => 
                           n7672, ZN => n7679);
   U13496 : NAND3_X1 port map( A1 => n7677, A2 => n7676, A3 => n3275, ZN => 
                           n7678);
   U13497 : XNOR2_X1 port map( A => n8116, B => n8296, ZN => n9020);
   U13498 : INV_X1 port map( A => n9020, ZN => n7680);
   U13499 : XNOR2_X1 port map( A => n7680, B => n7681, ZN => n7706);
   U13500 : MUX2_X1 port map( A => n7685, B => n7684, S => n7962, Z => n7686);
   U13501 : OAI21_X2 port map( B1 => n7687, B2 => n7961, A => n7686, ZN => 
                           n8675);
   U13502 : XNOR2_X1 port map( A => n8270, B => n8675, ZN => n7704);
   U13503 : NOR2_X1 port map( A1 => n7217, A2 => n7688, ZN => n7697);
   U13504 : NOR2_X1 port map( A1 => n7690, A2 => n7689, ZN => n7695);
   U13505 : INV_X1 port map( A => n7691, ZN => n7694);
   U13506 : INV_X1 port map( A => n7692, ZN => n7693);
   U13507 : NAND2_X1 port map( A1 => n8315, A2 => n7217, ZN => n7696);
   U13508 : NAND3_X1 port map( A1 => n7700, A2 => n7699, A3 => n8314, ZN => 
                           n7701);
   U13509 : XNOR2_X1 port map( A => n8203, B => n23620, ZN => n7703);
   U13510 : XNOR2_X1 port map( A => n7704, B => n7703, ZN => n7705);
   U13511 : MUX2_X1 port map( A => n25217, B => n9599, S => n9927, Z => n7839);
   U13512 : NAND2_X1 port map( A1 => n7860, A2 => n7707, ZN => n7709);
   U13513 : AOI21_X1 port map( B1 => n7709, B2 => n7708, A => n7865, ZN => 
                           n7712);
   U13514 : NAND2_X1 port map( A1 => n7714, A2 => n7713, ZN => n7844);
   U13515 : OAI211_X1 port map( C1 => n7718, C2 => n7844, A => n7717, B => 
                           n7716, ZN => n7720);
   U13516 : NAND2_X1 port map( A1 => n7722, A2 => n7721, ZN => n7723);
   U13517 : AND2_X1 port map( A1 => n7724, A2 => n7723, ZN => n7729);
   U13519 : MUX2_X1 port map( A => n7727, B => n7858, S => n7853, Z => n7728);
   U13520 : XNOR2_X1 port map( A => n8914, B => n8916, ZN => n8995);
   U13521 : XNOR2_X1 port map( A => n8797, B => n8995, ZN => n7744);
   U13522 : NAND2_X1 port map( A1 => n7733, A2 => n7732, ZN => n7737);
   U13523 : XNOR2_X1 port map( A => n8237, B => n8690, ZN => n7742);
   U13524 : INV_X1 port map( A => n7813, ZN => n7739);
   U13525 : NAND3_X1 port map( A1 => n7813, A2 => n8219, A3 => n9067, ZN => 
                           n7740);
   U13526 : INV_X1 port map( A => n2881, ZN => n23283);
   U13527 : XNOR2_X1 port map( A => n8691, B => n23283, ZN => n7741);
   U13528 : XNOR2_X1 port map( A => n7742, B => n7741, ZN => n7743);
   U13530 : INV_X1 port map( A => n9925, ZN => n9346);
   U13531 : NOR2_X1 port map( A1 => n25217, A2 => n9925, ZN => n9929);
   U13532 : XNOR2_X1 port map( A => n9002, B => n8638, ZN => n8907);
   U13533 : OR2_X1 port map( A1 => n7748, A2 => n8015, ZN => n7752);
   U13534 : OAI21_X1 port map( B1 => n25451, B2 => n8012, A => n8015, ZN => 
                           n7751);
   U13536 : NAND2_X1 port map( A1 => n5202, A2 => n7757, ZN => n7756);
   U13537 : OR2_X1 port map( A1 => n7758, A2 => n7757, ZN => n8004);
   U13538 : XNOR2_X1 port map( A => n9057, B => n8965, ZN => n8191);
   U13539 : INV_X1 port map( A => n8191, ZN => n7759);
   U13540 : XNOR2_X1 port map( A => n7759, B => n8907, ZN => n7780);
   U13541 : NOR2_X1 port map( A1 => n7760, A2 => n4880, ZN => n7764);
   U13542 : NAND2_X1 port map( A1 => n7762, A2 => n7761, ZN => n7763);
   U13543 : AOI22_X1 port map( A1 => n7766, A2 => n7765, B1 => n7764, B2 => 
                           n7763, ZN => n8244);
   U13544 : NOR2_X1 port map( A1 => n7768, A2 => n7767, ZN => n7772);
   U13545 : INV_X1 port map( A => n7772, ZN => n7775);
   U13546 : OAI21_X1 port map( B1 => n7772, B2 => n7771, A => n7770, ZN => 
                           n7774);
   U13548 : XNOR2_X1 port map( A => n9106, B => n3155, ZN => n7777);
   U13549 : XNOR2_X1 port map( A => n7778, B => n7777, ZN => n7779);
   U13550 : NAND2_X1 port map( A1 => n7781, A2 => n7788, ZN => n7786);
   U13551 : NAND2_X1 port map( A1 => n7783, A2 => n7782, ZN => n7785);
   U13552 : MUX2_X1 port map( A => n7786, B => n7785, S => n7784, Z => n7793);
   U13553 : NOR2_X1 port map( A1 => n7788, A2 => n7787, ZN => n7790);
   U13554 : OAI21_X1 port map( B1 => n7791, B2 => n7790, A => n7789, ZN => 
                           n7792);
   U13555 : XNOR2_X1 port map( A => n8313, B => n8366, ZN => n9010);
   U13556 : INV_X1 port map( A => n9010, ZN => n7808);
   U13557 : NAND2_X1 port map( A1 => n7795, A2 => n7794, ZN => n7796);
   U13558 : AOI21_X1 port map( B1 => n7797, B2 => n7796, A => n7800, ZN => 
                           n7807);
   U13559 : NAND3_X1 port map( A1 => n7800, A2 => n7799, A3 => n7798, ZN => 
                           n7805);
   U13560 : NAND3_X1 port map( A1 => n7803, A2 => n7802, A3 => n7801, ZN => 
                           n7804);
   U13561 : NAND2_X1 port map( A1 => n7805, A2 => n7804, ZN => n7806);
   U13562 : XNOR2_X1 port map( A => n7808, B => n8252, ZN => n7837);
   U13563 : OAI21_X1 port map( B1 => n7810, B2 => n9066, A => n7809, ZN => 
                           n8220);
   U13564 : NAND2_X1 port map( A1 => n7814, A2 => n7813, ZN => n9070);
   U13565 : OAI21_X1 port map( B1 => n7819, B2 => n7816, A => n7971, ZN => 
                           n7818);
   U13566 : NAND2_X1 port map( A1 => n7818, A2 => n7817, ZN => n7824);
   U13567 : NAND3_X1 port map( A1 => n7819, A2 => n7973, A3 => n7971, ZN => 
                           n7823);
   U13568 : NAND3_X2 port map( A1 => n7824, A2 => n7823, A3 => n7822, ZN => 
                           n8746);
   U13569 : XNOR2_X1 port map( A => n8746, B => n8507, ZN => n7835);
   U13570 : NAND3_X1 port map( A1 => n7989, A2 => n7983, A3 => n7984, ZN => 
                           n7833);
   U13571 : NAND3_X1 port map( A1 => n7983, A2 => n7982, A3 => n7825, ZN => 
                           n7832);
   U13573 : XNOR2_X1 port map( A => n8667, B => n1891, ZN => n7834);
   U13574 : XNOR2_X1 port map( A => n7835, B => n7834, ZN => n7836);
   U13575 : INV_X1 port map( A => n9599, ZN => n9604);
   U13576 : NOR2_X1 port map( A1 => n9603, A2 => n9604, ZN => n7838);
   U13577 : NOR2_X1 port map( A1 => n7840, A2 => n7714, ZN => n7845);
   U13578 : OAI21_X1 port map( B1 => n7844, B2 => n7843, A => n7842, ZN => 
                           n8374);
   U13579 : INV_X1 port map( A => n9176, ZN => n7846);
   U13580 : XNOR2_X1 port map( A => n7846, B => n8507, ZN => n7848);
   U13581 : XNOR2_X1 port map( A => n8786, B => n8517, ZN => n7847);
   U13582 : XNOR2_X1 port map( A => n7848, B => n7847, ZN => n7876);
   U13583 : INV_X1 port map( A => n8450, ZN => n8126);
   U13584 : INV_X1 port map( A => n7849, ZN => n7852);
   U13585 : NAND2_X1 port map( A1 => n7857, A2 => n24072, ZN => n7851);
   U13586 : AOI21_X1 port map( B1 => n7852, B2 => n7851, A => n7855, ZN => 
                           n7859);
   U13587 : NAND3_X1 port map( A1 => n7855, A2 => n7854, A3 => n7853, ZN => 
                           n7856);
   U13588 : XNOR2_X1 port map( A => n8126, B => n8789, ZN => n7874);
   U13589 : NAND3_X1 port map( A1 => n4537, A2 => n7862, A3 => n7861, ZN => 
                           n7871);
   U13590 : NAND3_X1 port map( A1 => n7865, A2 => n4536, A3 => n7864, ZN => 
                           n7870);
   U13591 : NAND3_X1 port map( A1 => n7868, A2 => n7867, A3 => n24576, ZN => 
                           n7869);
   U13592 : XNOR2_X1 port map( A => n9179, B => n20284, ZN => n7873);
   U13593 : XNOR2_X1 port map( A => n7874, B => n7873, ZN => n7875);
   U13594 : XNOR2_X1 port map( A => n8952, B => n8799, ZN => n7878);
   U13595 : XNOR2_X1 port map( A => n8691, B => n21711, ZN => n7877);
   U13596 : XNOR2_X1 port map( A => n7878, B => n7877, ZN => n7907);
   U13598 : INV_X1 port map( A => n7892, ZN => n7894);
   U13599 : XNOR2_X1 port map( A => n7895, B => n8951, ZN => n9138);
   U13602 : INV_X1 port map( A => n8468, ZN => n7904);
   U13603 : XNOR2_X1 port map( A => n8796, B => n7904, ZN => n7905);
   U13604 : XNOR2_X1 port map( A => n9138, B => n7905, ZN => n7906);
   U13605 : XNOR2_X1 port map( A => n8673, B => n9188, ZN => n7922);
   U13606 : AND2_X1 port map( A1 => n7915, A2 => n7918, ZN => n7916);
   U13607 : MUX2_X1 port map( A => n430, B => n7916, S => n7917, Z => n7921);
   U13608 : NAND2_X1 port map( A1 => n7917, A2 => n3348, ZN => n7919);
   U13609 : AOI21_X1 port map( B1 => n7920, B2 => n7919, A => n7918, ZN => 
                           n8078);
   U13610 : XNOR2_X1 port map( A => n9189, B => n2191, ZN => n8268);
   U13611 : XNOR2_X1 port map( A => n8268, B => n7922, ZN => n7940);
   U13612 : INV_X1 port map( A => n7933, ZN => n7936);
   U13613 : OAI21_X1 port map( B1 => n7924, B2 => n7923, A => n5607, ZN => 
                           n7935);
   U13614 : NOR2_X1 port map( A1 => n7927, A2 => n7926, ZN => n7931);
   U13615 : INV_X1 port map( A => n7928, ZN => n7929);
   U13616 : XNOR2_X1 port map( A => n8203, B => n24445, ZN => n7938);
   U13617 : XNOR2_X1 port map( A => n8754, B => n1777, ZN => n7937);
   U13618 : XNOR2_X1 port map( A => n7938, B => n7937, ZN => n7939);
   U13619 : XNOR2_X1 port map( A => n7940, B => n7939, ZN => n7941);
   U13620 : MUX2_X1 port map( A => n9939, B => n9449, S => n9276, Z => n8030);
   U13621 : INV_X1 port map( A => n7941, ZN => n9908);
   U13622 : OAI22_X1 port map( A1 => n7944, A2 => n24474, B1 => n7946, B2 => 
                           n7943, ZN => n7951);
   U13623 : XNOR2_X1 port map( A => n9149, B => n8959, ZN => n8263);
   U13624 : INV_X1 port map( A => n7954, ZN => n7955);
   U13625 : INV_X1 port map( A => n9057, ZN => n7958);
   U13626 : XNOR2_X1 port map( A => n8770, B => n7958, ZN => n7959);
   U13627 : XNOR2_X1 port map( A => n8263, B => n7959, ZN => n7970);
   U13629 : XNOR2_X1 port map( A => n8698, B => n8961, ZN => n7968);
   U13630 : XNOR2_X1 port map( A => n8964, B => n20825, ZN => n7967);
   U13631 : XNOR2_X1 port map( A => n7968, B => n7967, ZN => n7969);
   U13632 : XNOR2_X1 port map( A => n7969, B => n7970, ZN => n9907);
   U13633 : AND2_X1 port map( A1 => n9907, A2 => n9908, ZN => n9937);
   U13634 : MUX2_X1 port map( A => n7976, B => n7975, S => n7974, Z => n7978);
   U13635 : XNOR2_X1 port map( A => n24946, B => n8069, ZN => n7981);
   U13636 : XNOR2_X1 port map( A => n7981, B => n7980, ZN => n8002);
   U13637 : NAND2_X1 port map( A1 => n7989, A2 => n7984, ZN => n7986);
   U13638 : MUX2_X1 port map( A => n7987, B => n7986, S => n7985, Z => n7988);
   U13639 : MUX2_X1 port map( A => n7992, B => n7990, S => n7993, Z => n7997);
   U13640 : NAND2_X1 port map( A1 => n7992, A2 => n7991, ZN => n7995);
   U13642 : XNOR2_X1 port map( A => n8779, B => n9158, ZN => n8000);
   U13643 : XNOR2_X1 port map( A => n8446, B => n1757, ZN => n7999);
   U13644 : XNOR2_X1 port map( A => n8000, B => n7999, ZN => n8001);
   U13645 : MUX2_X1 port map( A => n9905, B => n9908, S => n9939, Z => n8029);
   U13646 : AOI21_X1 port map( B1 => n8004, B2 => n8003, A => n5202, ZN => 
                           n8008);
   U13647 : AOI21_X1 port map( B1 => n8006, B2 => n8005, A => n432, ZN => n8007
                           );
   U13648 : XNOR2_X1 port map( A => n8458, B => n8970, ZN => n8010);
   U13649 : XNOR2_X1 port map( A => n9043, B => n92, ZN => n8009);
   U13650 : XNOR2_X1 port map( A => n8010, B => n8009, ZN => n8028);
   U13652 : NAND3_X1 port map( A1 => n8013, A2 => n8014, A3 => n8015, ZN => 
                           n8018);
   U13653 : XNOR2_X1 port map( A => n9169, B => n8501, ZN => n8288);
   U13654 : NAND3_X1 port map( A1 => n3615, A2 => n8024, A3 => n8023, ZN => 
                           n8025);
   U13655 : XNOR2_X1 port map( A => n8542, B => n9040, ZN => n8766);
   U13656 : XNOR2_X1 port map( A => n8288, B => n8766, ZN => n8027);
   U13658 : OAI21_X1 port map( B1 => n10369, B2 => n10363, A => n8031, ZN => 
                           n8032);
   U13660 : XNOR2_X1 port map( A => n8826, B => n8675, ZN => n8297);
   U13661 : XNOR2_X1 port map( A => n8647, B => n3178, ZN => n8035);
   U13662 : XNOR2_X1 port map( A => n8036, B => n8035, ZN => n8037);
   U13663 : XNOR2_X1 port map( A => n8746, B => n2033, ZN => n8038);
   U13664 : XNOR2_X1 port map( A => n8038, B => n8313, ZN => n8040);
   U13665 : XNOR2_X1 port map( A => n9114, B => n8040, ZN => n8043);
   U13666 : XNOR2_X1 port map( A => n9181, B => n8651, ZN => n8041);
   U13667 : XNOR2_X1 port map( A => n9011, B => n8041, ZN => n8042);
   U13668 : XNOR2_X1 port map( A => n8782, B => n25235, ZN => n8044);
   U13669 : XNOR2_X1 port map( A => n8807, B => n8682, ZN => n9092);
   U13670 : XNOR2_X1 port map( A => n9092, B => n8044, ZN => n8048);
   U13671 : XNOR2_X1 port map( A => n8278, B => n8612, ZN => n8046);
   U13672 : XNOR2_X1 port map( A => n8400, B => n2042, ZN => n8045);
   U13673 : XNOR2_X1 port map( A => n8046, B => n8045, ZN => n8047);
   U13675 : XNOR2_X1 port map( A => n8965, B => n1758, ZN => n8049);
   U13676 : XNOR2_X1 port map( A => n9106, B => n8638, ZN => n8052);
   U13677 : INV_X1 port map( A => n9107, ZN => n8051);
   U13678 : XNOR2_X1 port map( A => n8052, B => n8051, ZN => n8310);
   U13679 : XNOR2_X1 port map( A => n8053, B => n8310, ZN => n9856);
   U13680 : XNOR2_X1 port map( A => n8913, B => n8730, ZN => n8953);
   U13681 : XNOR2_X1 port map( A => n8953, B => n9124, ZN => n8057);
   U13682 : XNOR2_X1 port map( A => n24547, B => n9140, ZN => n8055);
   U13683 : XNOR2_X1 port map( A => n8916, B => n20046, ZN => n8054);
   U13684 : XNOR2_X1 port map( A => n8055, B => n8054, ZN => n8056);
   U13685 : XNOR2_X1 port map( A => n8057, B => n8056, ZN => n9560);
   U13686 : MUX2_X1 port map( A => n9856, B => n9560, S => n238, Z => n8063);
   U13687 : XNOR2_X1 port map( A => n8812, B => n8706, ZN => n9095);
   U13688 : XNOR2_X1 port map( A => n8058, B => n9095, ZN => n8062);
   U13689 : XNOR2_X1 port map( A => n8899, B => n8760, ZN => n8060);
   U13690 : INV_X1 port map( A => n16, ZN => n21861);
   U13691 : XNOR2_X1 port map( A => n8896, B => n21861, ZN => n8059);
   U13692 : XNOR2_X1 port map( A => n8060, B => n8059, ZN => n8061);
   U13693 : XNOR2_X1 port map( A => n8062, B => n8061, ZN => n9554);
   U13695 : MUX2_X1 port map( A => n9905, B => n24511, S => n9276, Z => n8068);
   U13696 : NAND2_X1 port map( A1 => n9449, A2 => n9907, ZN => n8066);
   U13697 : NAND2_X1 port map( A1 => n9939, A2 => n24511, ZN => n8065);
   U13698 : MUX2_X1 port map( A => n8066, B => n8065, S => n9905, Z => n8067);
   U13699 : OAI21_X1 port map( B1 => n8068, B2 => n9449, A => n8067, ZN => 
                           n10990);
   U13700 : XNOR2_X1 port map( A => n8865, B => n8714, ZN => n8073);
   U13701 : XNOR2_X1 port map( A => n8071, B => n8070, ZN => n8072);
   U13702 : XNOR2_X1 port map( A => n8073, B => n8072, ZN => n9694);
   U13703 : XNOR2_X1 port map( A => n8478, B => n8824, ZN => n8720);
   U13704 : OAI21_X1 port map( B1 => n8076, B2 => n435, A => n8075, ZN => n8077
                           );
   U13705 : NOR2_X1 port map( A1 => n8078, A2 => n8077, ZN => n8079);
   U13706 : XNOR2_X1 port map( A => n8341, B => n8079, ZN => n8882);
   U13707 : XNOR2_X1 port map( A => n8720, B => n8882, ZN => n8083);
   U13708 : XNOR2_X1 port map( A => n8674, B => n8339, ZN => n8081);
   U13709 : XNOR2_X1 port map( A => n8203, B => n23883, ZN => n8080);
   U13710 : XNOR2_X1 port map( A => n8081, B => n8080, ZN => n8082);
   U13711 : XNOR2_X1 port map( A => n8666, B => n8507, ZN => n8085);
   U13712 : XNOR2_X1 port map( A => n8084, B => n8085, ZN => n8087);
   U13713 : XNOR2_X1 port map( A => n8375, B => n19392, ZN => n8086);
   U13714 : XNOR2_X1 port map( A => n9179, B => n8412, ZN => n8862);
   U13715 : XNOR2_X1 port map( A => n8498, B => n8813, ZN => n8726);
   U13716 : XNOR2_X1 port map( A => n8088, B => n9169, ZN => n8872);
   U13717 : XNOR2_X1 port map( A => n8726, B => n8872, ZN => n8092);
   U13718 : XNOR2_X1 port map( A => n8345, B => n8897, ZN => n8090);
   U13719 : XNOR2_X1 port map( A => n9043, B => n853, ZN => n8089);
   U13720 : XNOR2_X1 port map( A => n8090, B => n8089, ZN => n8091);
   U13721 : XNOR2_X1 port map( A => n8635, B => n8093, ZN => n8741);
   U13722 : XNOR2_X1 port map( A => n9149, B => n8361, ZN => n8855);
   U13723 : INV_X1 port map( A => n8855, ZN => n8585);
   U13724 : XNOR2_X1 port map( A => n8585, B => n8741, ZN => n8097);
   U13725 : XNOR2_X1 port map( A => n8360, B => n9057, ZN => n8095);
   U13726 : XNOR2_X1 port map( A => n8699, B => n912, ZN => n8094);
   U13727 : XNOR2_X1 port map( A => n8095, B => n8094, ZN => n8096);
   U13729 : XNOR2_X1 port map( A => n8353, B => n9121, ZN => n8844);
   U13730 : INV_X1 port map( A => n8844, ZN => n8578);
   U13731 : XNOR2_X1 port map( A => n8578, B => n8731, ZN => n8101);
   U13732 : XNOR2_X1 port map( A => n8468, B => n8687, ZN => n8099);
   U13733 : XNOR2_X1 port map( A => n8147, B => n3158, ZN => n8098);
   U13734 : XNOR2_X1 port map( A => n8099, B => n8098, ZN => n8100);
   U13735 : XNOR2_X1 port map( A => n8980, B => n9035, ZN => n8103);
   U13736 : XNOR2_X1 port map( A => n8103, B => n8102, ZN => n8104);
   U13737 : XNOR2_X1 port map( A => n8698, B => n9002, ZN => n8106);
   U13738 : INV_X1 port map( A => n2211, ZN => n23432);
   U13739 : XNOR2_X1 port map( A => n8962, B => n23432, ZN => n8105);
   U13740 : XNOR2_X1 port map( A => n8106, B => n8105, ZN => n8111);
   U13741 : XNOR2_X1 port map( A => n25407, B => n9059, ZN => n8109);
   U13742 : INV_X1 port map( A => n8853, ZN => n8107);
   U13743 : XNOR2_X1 port map( A => n8107, B => n8771, ZN => n8108);
   U13744 : XNOR2_X1 port map( A => n8108, B => n8109, ZN => n8110);
   U13745 : XNOR2_X1 port map( A => n8460, B => n8458, ZN => n8113);
   U13746 : INV_X1 port map( A => n2040, ZN => n22635);
   U13747 : XNOR2_X1 port map( A => n8896, B => n22635, ZN => n8115);
   U13748 : XNOR2_X1 port map( A => n8898, B => n9044, ZN => n8114);
   U13749 : INV_X1 port map( A => n8116, ZN => n8340);
   U13750 : XNOR2_X1 port map( A => n8340, B => n8673, ZN => n8118);
   U13751 : XNOR2_X1 port map( A => n8118, B => n8117, ZN => n8123);
   U13752 : XNOR2_X1 port map( A => n8647, B => n2746, ZN => n8120);
   U13753 : XNOR2_X1 port map( A => n8121, B => n8120, ZN => n8122);
   U13754 : INV_X1 port map( A => n9182, ZN => n8124);
   U13755 : XNOR2_X1 port map( A => n8366, B => n8124, ZN => n8216);
   U13756 : XNOR2_X1 port map( A => n8125, B => n8216, ZN => n8130);
   U13757 : XNOR2_X1 port map( A => n8126, B => n8651, ZN => n8128);
   U13758 : XNOR2_X1 port map( A => n8860, B => n3129, ZN => n8127);
   U13759 : XNOR2_X1 port map( A => n8128, B => n8127, ZN => n8129);
   U13760 : XNOR2_X1 port map( A => n8131, B => n8198, ZN => n8136);
   U13761 : XNOR2_X1 port map( A => n8132, B => n9082, ZN => n8134);
   U13762 : XNOR2_X1 port map( A => n8691, B => n2228, ZN => n8133);
   U13763 : XNOR2_X1 port map( A => n8134, B => n8133, ZN => n8135);
   U13764 : NAND3_X1 port map( A1 => n9945, A2 => n227, A3 => n24054, ZN => 
                           n8137);
   U13765 : INV_X1 port map( A => n10993, ZN => n10327);
   U13766 : NOR2_X1 port map( A1 => n10924, A2 => n10327, ZN => n8145);
   U13767 : NAND2_X1 port map( A1 => n8140, A2 => n9281, ZN => n8144);
   U13768 : INV_X1 port map( A => n8141, ZN => n9469);
   U13769 : MUX2_X1 port map( A => n8146, B => n8145, S => n10405, Z => n8181);
   U13770 : XNOR2_X1 port map( A => n8846, B => n8917, ZN => n8236);
   U13771 : XNOR2_X1 port map( A => n8147, B => n2190, ZN => n8148);
   U13772 : XNOR2_X1 port map( A => n8149, B => n8148, ZN => n8150);
   U13773 : XNOR2_X1 port map( A => n8634, B => n8909, ZN => n8852);
   U13774 : INV_X1 port map( A => n9111, ZN => n8151);
   U13775 : XNOR2_X1 port map( A => n8151, B => n8852, ZN => n8156);
   U13776 : XNOR2_X1 port map( A => n8772, B => n8152, ZN => n8154);
   U13777 : INV_X1 port map( A => n3133, ZN => n23072);
   U13778 : XNOR2_X1 port map( A => n8360, B => n23072, ZN => n8153);
   U13779 : XNOR2_X1 port map( A => n8154, B => n8153, ZN => n8155);
   U13780 : XNOR2_X1 port map( A => n8285, B => n8620, ZN => n9096);
   U13781 : INV_X1 port map( A => n9096, ZN => n8158);
   U13782 : XNOR2_X1 port map( A => n8158, B => n8301, ZN => n8162);
   U13783 : XNOR2_X1 port map( A => n9167, B => n8345, ZN => n8160);
   U13784 : XNOR2_X1 port map( A => n24056, B => n4233, ZN => n8159);
   U13785 : XNOR2_X1 port map( A => n8160, B => n8159, ZN => n8161);
   U13786 : XNOR2_X2 port map( A => n8162, B => n8161, ZN => n9886);
   U13787 : XNOR2_X1 port map( A => n8596, B => n8923, ZN => n8859);
   U13788 : XNOR2_X1 port map( A => n8859, B => n9115, ZN => n8166);
   U13789 : XNOR2_X1 port map( A => n8787, B => n8375, ZN => n8164);
   U13790 : INV_X1 port map( A => n2087, ZN => n22745);
   U13791 : XNOR2_X1 port map( A => n9181, B => n22745, ZN => n8163);
   U13792 : XNOR2_X1 port map( A => n8164, B => n8163, ZN => n8165);
   U13793 : INV_X1 port map( A => Key(44), ZN => n21942);
   U13794 : INV_X1 port map( A => n21942, ZN => n21944);
   U13795 : XNOR2_X1 port map( A => n8755, B => n21944, ZN => n8167);
   U13796 : XNOR2_X1 port map( A => n8167, B => n8339, ZN => n8169);
   U13797 : XNOR2_X1 port map( A => n9016, B => n8168, ZN => n9101);
   U13798 : XNOR2_X1 port map( A => n8169, B => n9101, ZN => n8171);
   U13799 : XNOR2_X1 port map( A => n8928, B => n9196, ZN => n8170);
   U13800 : XNOR2_X1 port map( A => n8604, B => n8170, ZN => n8884);
   U13801 : XNOR2_X1 port map( A => n8171, B => n8884, ZN => n9454);
   U13802 : NAND2_X1 port map( A1 => n9454, A2 => n25069, ZN => n8177);
   U13803 : XNOR2_X1 port map( A => n8891, B => n8588, ZN => n8868);
   U13804 : XNOR2_X1 port map( A => n8868, B => n9089, ZN => n8176);
   U13805 : XNOR2_X1 port map( A => n8278, B => n641, ZN => n8173);
   U13806 : XNOR2_X1 port map( A => n8174, B => n8173, ZN => n8175);
   U13807 : XNOR2_X2 port map( A => n8176, B => n8175, ZN => n9565);
   U13809 : AOI21_X1 port map( B1 => n8177, B2 => n9565, A => n9563, ZN => 
                           n8178);
   U13810 : INV_X1 port map( A => n10994, ZN => n10326);
   U13811 : AND2_X1 port map( A1 => n10326, A2 => n10405, ZN => n10925);
   U13813 : NOR2_X2 port map( A1 => n8181, A2 => n8180, ZN => n12378);
   U13814 : XNOR2_X1 port map( A => n11914, B => n12378, ZN => n11061);
   U13815 : XNOR2_X1 port map( A => n9155, B => n8782, ZN => n8713);
   U13818 : XNOR2_X1 port map( A => n8807, B => n2222, ZN => n8184);
   U13819 : XNOR2_X1 port map( A => n8778, B => n8184, ZN => n8185);
   U13820 : XNOR2_X1 port map( A => n8185, B => n8186, ZN => n9843);
   U13821 : INV_X1 port map( A => n8460, ZN => n8971);
   U13822 : XNOR2_X1 port map( A => n8971, B => n8499, ZN => n9165);
   U13823 : XNOR2_X1 port map( A => n8989, B => n9043, ZN => n8503);
   U13824 : XNOR2_X1 port map( A => n9165, B => n8503, ZN => n8190);
   U13825 : XNOR2_X1 port map( A => n8812, B => n8898, ZN => n8188);
   U13826 : INV_X1 port map( A => n2050, ZN => n21309);
   U13827 : XNOR2_X1 port map( A => n8760, B => n21309, ZN => n8187);
   U13828 : XNOR2_X1 port map( A => n8188, B => n8187, ZN => n8189);
   U13829 : XNOR2_X1 port map( A => n8191, B => n8192, ZN => n8196);
   U13830 : XNOR2_X1 port map( A => n8484, B => n9107, ZN => n8194);
   U13831 : XNOR2_X1 port map( A => n9002, B => n836, ZN => n8193);
   U13832 : XNOR2_X1 port map( A => n8193, B => n8194, ZN => n8195);
   U13833 : XNOR2_X1 port map( A => n8797, B => n8197, ZN => n8202);
   U13834 : INV_X1 port map( A => n8198, ZN => n8200);
   U13835 : XNOR2_X1 port map( A => n9141, B => n22702, ZN => n8199);
   U13836 : XNOR2_X1 port map( A => n8200, B => n8199, ZN => n8201);
   U13837 : XNOR2_X1 port map( A => n8721, B => n8340, ZN => n8204);
   U13838 : XNOR2_X1 port map( A => n8203, B => n9015, ZN => n8753);
   U13840 : XNOR2_X1 port map( A => n8826, B => n9190, ZN => n8206);
   U13841 : XNOR2_X1 port map( A => n9194, B => n21335, ZN => n8205);
   U13843 : INV_X1 port map( A => n8209, ZN => n8211);
   U13844 : INV_X1 port map( A => n17960, ZN => n23750);
   U13845 : AOI21_X1 port map( B1 => n8211, B2 => n8509, A => n23750, ZN => 
                           n8210);
   U13846 : NAND2_X1 port map( A1 => n8210, A2 => n8514, ZN => n8214);
   U13847 : NAND3_X1 port map( A1 => n8211, A2 => n8509, A3 => n23750, ZN => 
                           n8213);
   U13848 : NAND3_X1 port map( A1 => n8214, A2 => n8213, A3 => n8212, ZN => 
                           n8215);
   U13849 : XNOR2_X1 port map( A => n8820, B => n8215, ZN => n8218);
   U13850 : INV_X1 port map( A => n8216, ZN => n8217);
   U13851 : NAND2_X1 port map( A1 => n8221, A2 => n8219, ZN => n9069);
   U13852 : OAI211_X1 port map( C1 => n8221, C2 => n8220, A => n9070, B => 
                           n9069, ZN => n8222);
   U13853 : XNOR2_X1 port map( A => n8222, B => n8746, ZN => n8223);
   U13854 : AND2_X1 port map( A1 => n25486, A2 => n9845, ZN => n10122);
   U13855 : XNOR2_X1 port map( A => n8492, B => n25235, ZN => n8226);
   U13856 : XNOR2_X1 port map( A => n8868, B => n8226, ZN => n8229);
   U13857 : XNOR2_X1 port map( A => n8615, B => n8446, ZN => n8684);
   U13858 : XNOR2_X1 port map( A => n8280, B => n688, ZN => n8227);
   U13859 : XNOR2_X1 port map( A => n8684, B => n8227, ZN => n8228);
   U13860 : XNOR2_X1 port map( A => n8498, B => n8897, ZN => n8231);
   U13861 : XNOR2_X1 port map( A => n8231, B => n8230, ZN => n8235);
   U13862 : XNOR2_X1 port map( A => n8987, B => n8874, ZN => n8233);
   U13863 : XNOR2_X1 port map( A => n24056, B => n859, ZN => n8232);
   U13864 : XNOR2_X1 port map( A => n8233, B => n8232, ZN => n8234);
   U13865 : XNOR2_X1 port map( A => n8235, B => n8234, ZN => n9829);
   U13866 : NAND2_X1 port map( A1 => n9832, A2 => n9829, ZN => n10185);
   U13867 : INV_X1 port map( A => n8236, ZN => n8239);
   U13868 : XNOR2_X1 port map( A => n8238, B => n8237, ZN => n8274);
   U13869 : XNOR2_X1 port map( A => n8239, B => n8274, ZN => n8243);
   U13870 : XNOR2_X1 port map( A => n8913, B => n8687, ZN => n8241);
   U13871 : XNOR2_X1 port map( A => n8691, B => n20744, ZN => n8240);
   U13872 : XNOR2_X1 port map( A => n8241, B => n8240, ZN => n8242);
   U13873 : XNOR2_X1 port map( A => n8243, B => n8242, ZN => n10175);
   U13874 : XNOR2_X1 port map( A => n9001, B => n8852, ZN => n8248);
   U13875 : XNOR2_X1 port map( A => n8699, B => n2834, ZN => n8245);
   U13876 : XNOR2_X1 port map( A => n8246, B => n8245, ZN => n8247);
   U13877 : XNOR2_X1 port map( A => n8250, B => n8249, ZN => n8254);
   U13878 : XNOR2_X1 port map( A => n8923, B => n876, ZN => n8251);
   U13879 : XNOR2_X1 port map( A => n8251, B => n8252, ZN => n8253);
   U13880 : NAND2_X1 port map( A1 => n10186, A2 => n10178, ZN => n8262);
   U13881 : XNOR2_X1 port map( A => n8928, B => n8478, ZN => n8255);
   U13882 : XNOR2_X1 port map( A => n8256, B => n8255, ZN => n8260);
   U13883 : XNOR2_X1 port map( A => n8935, B => n23476, ZN => n8258);
   U13884 : XNOR2_X1 port map( A => n8673, B => n8270, ZN => n8257);
   U13885 : XNOR2_X1 port map( A => n8258, B => n8257, ZN => n8259);
   U13886 : NAND2_X1 port map( A1 => n10176, A2 => n10177, ZN => n10181);
   U13887 : INV_X1 port map( A => n10181, ZN => n8261);
   U13888 : XNOR2_X1 port map( A => n9147, B => n9058, ZN => n8851);
   U13889 : XNOR2_X1 port map( A => n8265, B => n8264, ZN => n8266);
   U13890 : INV_X1 port map( A => n8523, ZN => n9804);
   U13891 : XNOR2_X1 port map( A => n9196, B => n8880, ZN => n8827);
   U13892 : XNOR2_X1 port map( A => n8270, B => n2735, ZN => n8271);
   U13893 : XNOR2_X1 port map( A => n8271, B => n8827, ZN => n8272);
   U13894 : XNOR2_X1 port map( A => n8952, B => n681, ZN => n8273);
   U13895 : XNOR2_X1 port map( A => n9140, B => n9081, ZN => n8843);
   U13896 : XNOR2_X1 port map( A => n8843, B => n8273, ZN => n8277);
   U13897 : XNOR2_X1 port map( A => n9121, B => n8795, ZN => n8275);
   U13898 : XNOR2_X1 port map( A => n8275, B => n8274, ZN => n8276);
   U13899 : XNOR2_X1 port map( A => n8277, B => n8276, ZN => n9531);
   U13900 : INV_X1 port map( A => n9531, ZN => n9533);
   U13901 : XNOR2_X1 port map( A => n8278, B => n9034, ZN => n8866);
   U13902 : INV_X1 port map( A => n8866, ZN => n8805);
   U13903 : XNOR2_X1 port map( A => n8805, B => n8279, ZN => n8284);
   U13904 : XNOR2_X1 port map( A => n8491, B => n8069, ZN => n8282);
   U13905 : XNOR2_X1 port map( A => n8280, B => n1935, ZN => n8281);
   U13906 : XNOR2_X1 port map( A => n8282, B => n8281, ZN => n8283);
   U13908 : XNOR2_X1 port map( A => n8285, B => n2126, ZN => n8286);
   U13909 : XNOR2_X1 port map( A => n8287, B => n8286, ZN => n8290);
   U13910 : XNOR2_X1 port map( A => n25228, B => n9167, ZN => n8873);
   U13911 : XNOR2_X1 port map( A => n8873, B => n8288, ZN => n8289);
   U13912 : OAI22_X1 port map( A1 => n9531, A2 => n8523, B1 => n10113, B2 => 
                           n9806, ZN => n9809);
   U13913 : XNOR2_X1 port map( A => n8292, B => n8291, ZN => n8295);
   U13914 : XNOR2_X1 port map( A => n9181, B => n9075, ZN => n8858);
   U13915 : INV_X1 port map( A => n1875, ZN => n21500);
   U13916 : XNOR2_X1 port map( A => n9179, B => n21500, ZN => n8293);
   U13917 : XNOR2_X1 port map( A => n8858, B => n8293, ZN => n8294);
   U13918 : XNOR2_X1 port map( A => n8295, B => n8294, ZN => n9807);
   U13919 : INV_X1 port map( A => n9807, ZN => n9338);
   U13920 : XNOR2_X1 port map( A => n8604, B => n8296, ZN => n8648);
   U13921 : XNOR2_X1 port map( A => n8671, B => n8648, ZN => n8300);
   U13922 : XNOR2_X1 port map( A => n8754, B => n2137, ZN => n8298);
   U13923 : XNOR2_X1 port map( A => n8297, B => n8298, ZN => n8299);
   U13924 : INV_X1 port map( A => n8327, ZN => n9817);
   U13925 : INV_X1 port map( A => n8301, ZN => n8302);
   U13926 : XNOR2_X1 port map( A => n8302, B => n9095, ZN => n8306);
   U13927 : XNOR2_X1 port map( A => n8899, B => n9044, ZN => n8304);
   U13928 : XNOR2_X1 port map( A => n8542, B => n896, ZN => n8303);
   U13929 : XNOR2_X1 port map( A => n8304, B => n8303, ZN => n8305);
   U13930 : XNOR2_X2 port map( A => n8306, B => n8305, ZN => n10169);
   U13931 : NAND2_X1 port map( A1 => n9817, A2 => n10169, ZN => n10172);
   U13932 : XNOR2_X1 port map( A => n8964, B => n1855, ZN => n8308);
   U13933 : INV_X1 port map( A => n8634, ZN => n8307);
   U13934 : XNOR2_X1 port map( A => n8308, B => n8307, ZN => n8309);
   U13935 : XNOR2_X1 port map( A => n8309, B => n8696, ZN => n8312);
   U13936 : INV_X1 port map( A => n8310, ZN => n8311);
   U13938 : XNOR2_X1 port map( A => n8596, B => n8313, ZN => n8652);
   U13939 : XNOR2_X1 port map( A => n9114, B => n8652, ZN => n8324);
   U13940 : MUX2_X1 port map( A => n8317, B => n8315, S => n8314, Z => n8320);
   U13941 : NAND3_X1 port map( A1 => n8317, A2 => n8316, A3 => n433, ZN => 
                           n8318);
   U13942 : XNOR2_X1 port map( A => n8551, B => n20690, ZN => n8322);
   U13943 : XNOR2_X1 port map( A => n8787, B => n8786, ZN => n8321);
   U13944 : XNOR2_X1 port map( A => n8322, B => n8321, ZN => n8323);
   U13945 : XNOR2_X1 port map( A => n8324, B => n8323, ZN => n10170);
   U13946 : INV_X1 port map( A => n10170, ZN => n9814);
   U13947 : XNOR2_X1 port map( A => n8781, B => n8612, ZN => n8325);
   U13948 : XNOR2_X1 port map( A => n25020, B => n8325, ZN => n8326);
   U13949 : XNOR2_X1 port map( A => n8846, B => n20609, ZN => n8328);
   U13950 : XNOR2_X1 port map( A => n8689, B => n8328, ZN => n8331);
   U13951 : XNOR2_X1 port map( A => n8329, B => n9124, ZN => n8330);
   U13953 : XNOR2_X1 port map( A => n8333, B => n8867, ZN => n8335);
   U13954 : XNOR2_X1 port map( A => n8491, B => n1827, ZN => n8334);
   U13955 : XNOR2_X1 port map( A => n8335, B => n8334, ZN => n8338);
   U13956 : XNOR2_X1 port map( A => n8779, B => n8981, ZN => n8539);
   U13957 : XNOR2_X1 port map( A => n8336, B => n9158, ZN => n8715);
   U13958 : XNOR2_X1 port map( A => n8715, B => n8539, ZN => n8337);
   U13959 : XNOR2_X1 port map( A => n8339, B => n9188, ZN => n8719);
   U13960 : XNOR2_X1 port map( A => n8340, B => n9195, ZN => n8558);
   U13961 : XNOR2_X1 port map( A => n8558, B => n8719, ZN => n8344);
   U13962 : XNOR2_X1 port map( A => n8341, B => n23679, ZN => n8342);
   U13963 : BUF_X2 port map( A => n10100, Z => n10095);
   U13965 : XNOR2_X1 port map( A => n8501, B => n8406, ZN => n8346);
   U13966 : XNOR2_X1 port map( A => n8725, B => n8346, ZN => n8350);
   U13967 : XNOR2_X1 port map( A => n9040, B => n8898, ZN => n8544);
   U13968 : INV_X1 port map( A => n663, ZN => n8347);
   U13969 : XNOR2_X1 port map( A => n8875, B => n8347, ZN => n8348);
   U13970 : XNOR2_X1 port map( A => n8544, B => n8348, ZN => n8349);
   U13971 : XNOR2_X1 port map( A => n8350, B => n8349, ZN => n9515);
   U13972 : XNOR2_X1 port map( A => n8354, B => n8353, ZN => n8356);
   U13973 : XNOR2_X1 port map( A => n8796, B => n8914, ZN => n8561);
   U13974 : INV_X1 port map( A => n8561, ZN => n8355);
   U13975 : XNOR2_X1 port map( A => n8355, B => n8356, ZN => n8358);
   U13976 : XNOR2_X1 port map( A => n8358, B => n8357, ZN => n8359);
   U13977 : XNOR2_X1 port map( A => n8961, B => n8360, ZN => n8738);
   U13978 : XNOR2_X1 port map( A => n8361, B => n2761, ZN => n8362);
   U13979 : XNOR2_X1 port map( A => n8738, B => n8362, ZN => n8365);
   U13980 : XNOR2_X1 port map( A => n8770, B => n9002, ZN => n8567);
   U13981 : XNOR2_X1 port map( A => n8363, B => n8567, ZN => n8364);
   U13982 : XNOR2_X2 port map( A => n8365, B => n8364, ZN => n10099);
   U13984 : NAND2_X1 port map( A1 => n24878, A2 => n8370, ZN => n8369);
   U13985 : OAI211_X1 port map( C1 => n8371, C2 => n8370, A => n8369, B => 
                           n8368, ZN => n8372);
   U13986 : INV_X1 port map( A => n8372, ZN => n8373);
   U13987 : OR2_X1 port map( A1 => n8374, A2 => n8373, ZN => n8376);
   U13988 : XNOR2_X1 port map( A => n8376, B => n8375, ZN => n8745);
   U13989 : XNOR2_X1 port map( A => n8745, B => n8549, ZN => n8380);
   U13990 : XNOR2_X1 port map( A => n8517, B => n8860, ZN => n8378);
   U13991 : XNOR2_X1 port map( A => n8412, B => n1896, ZN => n8377);
   U13992 : XNOR2_X1 port map( A => n8378, B => n8377, ZN => n8379);
   U13994 : INV_X1 port map( A => n8385, ZN => n8386);
   U13995 : XNOR2_X1 port map( A => n8720, B => n8386, ZN => n8390);
   U13996 : XNOR2_X1 port map( A => n9195, B => n2236, ZN => n8388);
   U13997 : XNOR2_X1 port map( A => n8388, B => n8387, ZN => n8389);
   U13998 : XNOR2_X1 port map( A => n8770, B => n2990, ZN => n8393);
   U13999 : INV_X1 port map( A => n8391, ZN => n8392);
   U14000 : XNOR2_X1 port map( A => n8393, B => n8392, ZN => n8397);
   U14001 : INV_X1 port map( A => n8741, ZN => n8394);
   U14002 : XNOR2_X1 port map( A => n8394, B => n8395, ZN => n8396);
   U14003 : XNOR2_X1 port map( A => n8396, B => n8397, ZN => n9384);
   U14004 : INV_X1 port map( A => n9384, ZN => n9849);
   U14005 : NOR2_X1 port map( A1 => n10161, A2 => n9849, ZN => n8420);
   U14006 : XNOR2_X1 port map( A => n8398, B => n8399, ZN => n8404);
   U14007 : XNOR2_X1 port map( A => n8779, B => n8492, ZN => n8402);
   U14008 : XNOR2_X1 port map( A => n8400, B => n881, ZN => n8401);
   U14009 : XNOR2_X1 port map( A => n8402, B => n8401, ZN => n8403);
   U14010 : XNOR2_X1 port map( A => n8403, B => n8404, ZN => n10158);
   U14011 : XNOR2_X1 port map( A => n8405, B => n8726, ZN => n8410);
   U14012 : XNOR2_X1 port map( A => n9040, B => n8406, ZN => n8408);
   U14013 : XNOR2_X1 port map( A => n8896, B => n3115, ZN => n8407);
   U14014 : XNOR2_X1 port map( A => n8408, B => n8407, ZN => n8409);
   U14015 : INV_X1 port map( A => n9348, ZN => n9592);
   U14017 : XNOR2_X1 port map( A => n8789, B => n8651, ZN => n8414);
   U14018 : XNOR2_X1 port map( A => n8412, B => n1826, ZN => n8413);
   U14019 : XNOR2_X1 port map( A => n8414, B => n8413, ZN => n8415);
   U14022 : NAND2_X1 port map( A1 => n8417, A2 => n9851, ZN => n8418);
   U14023 : XNOR2_X1 port map( A => n8796, B => n9081, ZN => n8423);
   U14024 : XNOR2_X1 port map( A => n8423, B => n8422, ZN => n8424);
   U14025 : XNOR2_X1 port map( A => n8425, B => n8424, ZN => n9349);
   U14026 : NAND3_X1 port map( A1 => n2311, A2 => n24470, A3 => n10935, ZN => 
                           n8426);
   U14027 : INV_X1 port map( A => n11464, ZN => n8664);
   U14028 : XNOR2_X1 port map( A => n8427, B => n8428, ZN => n8831);
   U14029 : XNOR2_X1 port map( A => n8994, B => n8831, ZN => n8432);
   U14030 : XNOR2_X1 port map( A => n8917, B => n2031, ZN => n8429);
   U14031 : XNOR2_X1 port map( A => n8430, B => n8429, ZN => n8431);
   U14032 : XNOR2_X1 port map( A => n8432, B => n8431, ZN => n10080);
   U14033 : XNOR2_X1 port map( A => n8635, B => n9107, ZN => n8835);
   U14034 : INV_X1 port map( A => n8772, ZN => n8433);
   U14035 : XNOR2_X1 port map( A => n8433, B => n8909, ZN => n8434);
   U14036 : XNOR2_X1 port map( A => n8835, B => n8434, ZN => n8438);
   U14037 : XNOR2_X1 port map( A => n8962, B => n673, ZN => n8435);
   U14038 : XNOR2_X1 port map( A => n8436, B => n8435, ZN => n8437);
   U14039 : XNOR2_X1 port map( A => n8439, B => n8824, ZN => n8440);
   U14040 : XNOR2_X1 port map( A => n8440, B => n8441, ZN => n8443);
   U14041 : XNOR2_X1 port map( A => n8755, B => n8935, ZN => n8442);
   U14042 : XNOR2_X1 port map( A => n8442, B => n8673, ZN => n9021);
   U14043 : XNOR2_X1 port map( A => n8443, B => n9021, ZN => n9787);
   U14044 : XNOR2_X1 port map( A => n8445, B => n8444, ZN => n8448);
   U14045 : XNOR2_X1 port map( A => n8447, B => n25235, ZN => n8983);
   U14047 : NAND2_X1 port map( A1 => n24575, A2 => n4256, ZN => n8456);
   U14048 : XNOR2_X1 port map( A => n9182, B => n21553, ZN => n8449);
   U14049 : XNOR2_X1 port map( A => n8449, B => n8923, ZN => n8451);
   U14050 : XNOR2_X1 port map( A => n8452, B => n8818, ZN => n8453);
   U14051 : XNOR2_X1 port map( A => n8453, B => n9011, ZN => n8454);
   U14052 : INV_X1 port map( A => n10082, ZN => n9306);
   U14053 : NAND2_X1 port map( A1 => n8456, A2 => n8455, ZN => n8465);
   U14054 : XNOR2_X1 port map( A => n8458, B => n8457, ZN => n8985);
   U14055 : INV_X1 port map( A => n8985, ZN => n8704);
   U14056 : XNOR2_X1 port map( A => n8704, B => n8459, ZN => n8464);
   U14057 : XNOR2_X1 port map( A => n8460, B => n8987, ZN => n8462);
   U14058 : INV_X1 port map( A => n869, ZN => n22440);
   U14059 : XNOR2_X1 port map( A => n8813, B => n22440, ZN => n8461);
   U14060 : XNOR2_X1 port map( A => n8462, B => n8461, ZN => n8463);
   U14061 : MUX2_X2 port map( A => n8466, B => n8465, S => n10088, Z => n11178)
                           ;
   U14062 : INV_X1 port map( A => n8467, ZN => n8470);
   U14063 : XNOR2_X1 port map( A => n8468, B => n8845, ZN => n9080);
   U14064 : INV_X1 port map( A => n9080, ZN => n8469);
   U14065 : XNOR2_X1 port map( A => n8470, B => n8469, ZN => n8474);
   U14066 : XNOR2_X1 port map( A => n8798, B => n8952, ZN => n8472);
   U14067 : XNOR2_X1 port map( A => n8690, B => n2215, ZN => n8471);
   U14068 : XNOR2_X1 port map( A => n8472, B => n8471, ZN => n8473);
   U14069 : XNOR2_X1 port map( A => n8474, B => n8473, ZN => n8483);
   U14070 : INV_X1 port map( A => n8483, ZN => n9797);
   U14071 : XNOR2_X1 port map( A => n8475, B => n8476, ZN => n8722);
   U14072 : INV_X1 port map( A => n8722, ZN => n9051);
   U14073 : XNOR2_X1 port map( A => n9051, B => n8753, ZN => n8482);
   U14074 : XNOR2_X1 port map( A => n8477, B => n8478, ZN => n8480);
   U14075 : XNOR2_X1 port map( A => n8675, B => n2757, ZN => n8479);
   U14076 : XNOR2_X1 port map( A => n8480, B => n8479, ZN => n8481);
   U14077 : NAND2_X1 port map( A1 => n9797, A2 => n246, ZN => n8497);
   U14078 : XNOR2_X1 port map( A => n8484, B => n8853, ZN => n8739);
   U14079 : XNOR2_X1 port map( A => n8771, B => n9057, ZN => n8487);
   U14080 : XNOR2_X1 port map( A => n8485, B => n5286, ZN => n8486);
   U14081 : XNOR2_X1 port map( A => n8487, B => n8486, ZN => n8488);
   U14082 : XNOR2_X1 port map( A => n8489, B => n8488, ZN => n9998);
   U14083 : INV_X1 port map( A => n9998, ZN => n9796);
   U14084 : INV_X1 port map( A => n9796, ZN => n9669);
   U14085 : INV_X1 port map( A => n9155, ZN => n8490);
   U14086 : XNOR2_X1 port map( A => n8867, B => n8490, ZN => n9033);
   U14087 : XNOR2_X1 port map( A => n9033, B => n8778, ZN => n8496);
   U14088 : XNOR2_X1 port map( A => n8492, B => n8491, ZN => n8494);
   U14089 : XNOR2_X1 port map( A => n8682, B => n494, ZN => n8493);
   U14090 : XNOR2_X1 port map( A => n8494, B => n8493, ZN => n8495);
   U14091 : INV_X1 port map( A => n9798, ZN => n9310);
   U14092 : XNOR2_X1 port map( A => n8498, B => n8706, ZN => n8500);
   U14093 : XNOR2_X1 port map( A => n8499, B => n8875, ZN => n9042);
   U14094 : XNOR2_X1 port map( A => n9042, B => n8500, ZN => n8505);
   U14095 : INV_X1 port map( A => n891, ZN => n21359);
   U14096 : XNOR2_X1 port map( A => n8501, B => n21359, ZN => n8502);
   U14097 : XNOR2_X1 port map( A => n8503, B => n8502, ZN => n8504);
   U14098 : INV_X1 port map( A => n8521, ZN => n9671);
   U14099 : NAND2_X1 port map( A1 => n1796, A2 => n9671, ZN => n8522);
   U14100 : XNOR2_X1 port map( A => n8506, B => n8507, ZN => n8516);
   U14101 : NAND2_X1 port map( A1 => n8508, A2 => n8512, ZN => n8510);
   U14102 : OAI211_X1 port map( C1 => n8512, C2 => n8511, A => n8510, B => 
                           n8509, ZN => n8513);
   U14103 : NAND2_X1 port map( A1 => n8514, A2 => n8513, ZN => n8515);
   U14104 : XNOR2_X1 port map( A => n8515, B => n8860, ZN => n8748);
   U14105 : INV_X1 port map( A => n8748, ZN => n9065);
   U14106 : XNOR2_X1 port map( A => n8516, B => n9065, ZN => n8520);
   U14107 : XNOR2_X1 port map( A => n8667, B => n3062, ZN => n8518);
   U14108 : NOR2_X1 port map( A1 => n11178, A2 => n24591, ZN => n8611);
   U14109 : OAI21_X1 port map( B1 => n9533, B2 => n9338, A => n9805, ZN => 
                           n8526);
   U14110 : INV_X1 port map( A => n9806, ZN => n10116);
   U14111 : NOR2_X1 port map( A1 => n9805, A2 => n9530, ZN => n8524);
   U14112 : OAI21_X1 port map( B1 => n9339, B2 => n8524, A => n9807, ZN => 
                           n8525);
   U14113 : NAND2_X1 port map( A1 => n8530, A2 => n8527, ZN => n8529);
   U14114 : OAI211_X1 port map( C1 => n8531, C2 => n8530, A => n8529, B => 
                           n8528, ZN => n8532);
   U14115 : OAI211_X1 port map( C1 => n269, C2 => n8534, A => n8533, B => n8532
                           , ZN => n8535);
   U14116 : XNOR2_X1 port map( A => n9035, B => n8535, ZN => n8536);
   U14117 : XNOR2_X1 port map( A => n8537, B => n8536, ZN => n8950);
   U14118 : INV_X1 port map( A => n8950, ZN => n8541);
   U14119 : XNOR2_X1 port map( A => n8682, B => n21423, ZN => n8538);
   U14120 : INV_X1 port map( A => n9495, ZN => n9782);
   U14121 : XNOR2_X1 port map( A => n8543, B => n8760, ZN => n8977);
   U14122 : XNOR2_X1 port map( A => n8977, B => n8544, ZN => n8547);
   U14123 : XNOR2_X1 port map( A => n24056, B => n886, ZN => n8545);
   U14124 : XNOR2_X1 port map( A => n8706, B => n8545, ZN => n8546);
   U14126 : XNOR2_X1 port map( A => n8667, B => n2039, ZN => n8548);
   U14127 : XNOR2_X1 port map( A => n8548, B => n8923, ZN => n8550);
   U14128 : XNOR2_X1 port map( A => n8549, B => n8550, ZN => n8555);
   U14129 : XNOR2_X1 port map( A => n8746, B => n8551, ZN => n8553);
   U14130 : XNOR2_X1 port map( A => n8553, B => n8552, ZN => n8941);
   U14131 : INV_X1 port map( A => n8941, ZN => n8554);
   U14132 : XNOR2_X1 port map( A => n8554, B => n8555, ZN => n9297);
   U14133 : NAND2_X1 port map( A1 => n9676, A2 => n9780, ZN => n8575);
   U14134 : XNOR2_X1 port map( A => n8675, B => n2100, ZN => n8556);
   U14135 : XNOR2_X1 port map( A => n8730, B => n8690, ZN => n8560);
   U14136 : XNOR2_X1 port map( A => n8561, B => n8560, ZN => n8564);
   U14137 : XNOR2_X1 port map( A => n9082, B => n8799, ZN => n8955);
   U14138 : XNOR2_X1 port map( A => n8917, B => n1856, ZN => n8562);
   U14139 : XNOR2_X1 port map( A => n8955, B => n8562, ZN => n8563);
   U14140 : XNOR2_X1 port map( A => n8563, B => n8564, ZN => n9496);
   U14141 : INV_X1 port map( A => n9496, ZN => n9295);
   U14142 : INV_X1 port map( A => n9059, ZN => n8565);
   U14143 : XNOR2_X1 port map( A => n8565, B => n8909, ZN => n8566);
   U14144 : XNOR2_X1 port map( A => n8964, B => n9106, ZN => n8569);
   U14145 : XNOR2_X1 port map( A => n8965, B => n1833, ZN => n8568);
   U14146 : XNOR2_X1 port map( A => n8569, B => n8568, ZN => n8570);
   U14148 : NAND3_X1 port map( A1 => n9782, A2 => n25454, A3 => n1348, ZN => 
                           n8573);
   U14149 : NOR2_X1 port map( A1 => n11168, A2 => n24957, ZN => n8610);
   U14150 : XNOR2_X1 port map( A => n8576, B => n8951, ZN => n8577);
   U14152 : XNOR2_X1 port map( A => n8798, B => n14398, ZN => n8579);
   U14153 : XNOR2_X1 port map( A => n8580, B => n8579, ZN => n8581);
   U14154 : XNOR2_X1 port map( A => n8582, B => n8581, ZN => n9485);
   U14155 : XNOR2_X1 port map( A => n8771, B => n8634, ZN => n8583);
   U14156 : XNOR2_X1 port map( A => n8738, B => n8583, ZN => n8587);
   U14157 : XNOR2_X1 port map( A => n8769, B => n677, ZN => n8584);
   U14158 : XNOR2_X1 port map( A => n8585, B => n8584, ZN => n8586);
   U14159 : XNOR2_X1 port map( A => n8586, B => n8587, ZN => n9484);
   U14160 : XNOR2_X1 port map( A => n8588, B => n8780, ZN => n8614);
   U14161 : XNOR2_X1 port map( A => n8865, B => n8614, ZN => n8591);
   U14162 : XNOR2_X1 port map( A => n8980, B => n925, ZN => n8589);
   U14163 : XNOR2_X1 port map( A => n8715, B => n8589, ZN => n8590);
   U14164 : XNOR2_X1 port map( A => n1337, B => n8725, ZN => n8595);
   U14165 : XNOR2_X1 port map( A => n8874, B => n9041, ZN => n8593);
   U14166 : XNOR2_X1 port map( A => n8989, B => n2739, ZN => n8592);
   U14167 : XNOR2_X1 port map( A => n8593, B => n8592, ZN => n8594);
   U14168 : OAI22_X1 port map( A1 => n9485, A2 => n9484, B1 => n10006, B2 => 
                           n10008, ZN => n10012);
   U14169 : XNOR2_X1 port map( A => n8790, B => n8597, ZN => n8598);
   U14170 : XNOR2_X1 port map( A => n8745, B => n8598, ZN => n8601);
   U14171 : XNOR2_X1 port map( A => n8599, B => n8862, ZN => n8600);
   U14172 : XNOR2_X1 port map( A => n8601, B => n8600, ZN => n9299);
   U14173 : INV_X1 port map( A => n9299, ZN => n9724);
   U14174 : INV_X1 port map( A => n9485, ZN => n9725);
   U14175 : INV_X1 port map( A => n8719, ZN => n8602);
   U14176 : XNOR2_X1 port map( A => n8602, B => n8882, ZN => n8608);
   U14177 : INV_X1 port map( A => n9191, ZN => n8603);
   U14178 : XNOR2_X1 port map( A => n8604, B => n8603, ZN => n8606);
   U14179 : XNOR2_X1 port map( A => n9015, B => n23983, ZN => n8605);
   U14180 : XNOR2_X1 port map( A => n8606, B => n8605, ZN => n8607);
   U14181 : INV_X1 port map( A => n9484, ZN => n9301);
   U14182 : MUX2_X1 port map( A => n8611, B => n8610, S => n1338, Z => n8663);
   U14183 : XNOR2_X1 port map( A => n8613, B => n8612, ZN => n8982);
   U14184 : XNOR2_X1 port map( A => n8982, B => n8614, ZN => n8619);
   U14185 : XNOR2_X1 port map( A => n8806, B => n2826, ZN => n8617);
   U14186 : XNOR2_X1 port map( A => n8617, B => n9090, ZN => n8618);
   U14187 : XNOR2_X1 port map( A => n8619, B => n8618, ZN => n9772);
   U14188 : INV_X1 port map( A => n9772, ZN => n8644);
   U14189 : XNOR2_X1 port map( A => n8622, B => n8621, ZN => n8626);
   U14190 : XNOR2_X1 port map( A => n8899, B => n8896, ZN => n8624);
   U14191 : XNOR2_X1 port map( A => n8813, B => n2744, ZN => n8623);
   U14192 : XNOR2_X1 port map( A => n8624, B => n8623, ZN => n8625);
   U14193 : XNOR2_X1 port map( A => n24547, B => n8687, ZN => n9122);
   U14194 : XNOR2_X1 port map( A => n9122, B => n8628, ZN => n8632);
   U14195 : XNOR2_X1 port map( A => n8795, B => n8916, ZN => n8630);
   U14196 : INV_X1 port map( A => Key(119), ZN => n21533);
   U14197 : XNOR2_X1 port map( A => n8630, B => n8629, ZN => n8631);
   U14198 : XNOR2_X1 port map( A => n8633, B => n8699, ZN => n9110);
   U14199 : INV_X1 port map( A => n9110, ZN => n8637);
   U14200 : XNOR2_X1 port map( A => n8635, B => n8634, ZN => n8636);
   U14201 : XNOR2_X1 port map( A => n8637, B => n8636, ZN => n8642);
   U14202 : XNOR2_X1 port map( A => n8639, B => n8638, ZN => n9003);
   U14203 : XNOR2_X1 port map( A => n8769, B => n1745, ZN => n8640);
   U14204 : XNOR2_X1 port map( A => n9003, B => n8640, ZN => n8641);
   U14205 : OAI21_X1 port map( B1 => n8644, B2 => n4254, A => n8643, ZN => 
                           n9525);
   U14206 : NAND2_X1 port map( A1 => n8644, A2 => n10109, ZN => n8659);
   U14207 : XNOR2_X1 port map( A => n8824, B => n9016, ZN => n8646);
   U14208 : XNOR2_X1 port map( A => n9191, B => n3190, ZN => n8645);
   U14209 : XNOR2_X1 port map( A => n8646, B => n8645, ZN => n8650);
   U14210 : XNOR2_X1 port map( A => n8647, B => n8674, ZN => n9102);
   U14211 : XNOR2_X1 port map( A => n9102, B => n8648, ZN => n8649);
   U14212 : XNOR2_X1 port map( A => n8649, B => n8650, ZN => n9328);
   U14213 : INV_X1 port map( A => n9328, ZN => n9775);
   U14214 : INV_X1 port map( A => n10104, ZN => n9526);
   U14215 : NOR2_X1 port map( A1 => n9775, A2 => n9526, ZN => n8658);
   U14216 : XNOR2_X1 port map( A => n8666, B => n8651, ZN => n9117);
   U14217 : INV_X1 port map( A => n9117, ZN => n8922);
   U14218 : XNOR2_X1 port map( A => n8652, B => n8922, ZN => n8656);
   U14219 : XNOR2_X1 port map( A => n8790, B => n8818, ZN => n8654);
   U14220 : XNOR2_X1 port map( A => n9007, B => n1724, ZN => n8653);
   U14221 : XNOR2_X1 port map( A => n8654, B => n8653, ZN => n8655);
   U14222 : NAND2_X1 port map( A1 => n25393, A2 => n4254, ZN => n8657);
   U14223 : AOI22_X1 port map( A1 => n9525, A2 => n8659, B1 => n8658, B2 => 
                           n8657, ZN => n8660);
   U14224 : INV_X1 port map( A => n8660, ZN => n11170);
   U14225 : NOR2_X1 port map( A1 => n11170, A2 => n24957, ZN => n10937);
   U14226 : INV_X1 port map( A => n11172, ZN => n11175);
   U14227 : OAI21_X1 port map( B1 => n8660, B2 => n11175, A => n11178, ZN => 
                           n8661);
   U14228 : NOR2_X1 port map( A1 => n10937, A2 => n8661, ZN => n8662);
   U14230 : XNOR2_X1 port map( A => n8664, B => n11840, ZN => n11435);
   U14231 : XNOR2_X1 port map( A => n8666, B => n9073, ZN => n8669);
   U14232 : XNOR2_X1 port map( A => n8667, B => n887, ZN => n8668);
   U14233 : XNOR2_X1 port map( A => n8669, B => n8668, ZN => n8670);
   U14234 : INV_X1 port map( A => n9664, ZN => n9221);
   U14235 : XNOR2_X1 port map( A => n8675, B => n2005, ZN => n8676);
   U14236 : XNOR2_X1 port map( A => n8677, B => n8676, ZN => n8678);
   U14237 : INV_X1 port map( A => n9981, ZN => n9736);
   U14239 : XNOR2_X1 port map( A => n24598, B => n8947, ZN => n8686);
   U14240 : XNOR2_X1 port map( A => n8682, B => n1768, ZN => n8683);
   U14241 : XNOR2_X1 port map( A => n8684, B => n8683, ZN => n8685);
   U14242 : XNOR2_X1 port map( A => n8686, B => n8685, ZN => n9429);
   U14243 : MUX2_X1 port map( A => n9221, B => n9736, S => n3799, Z => n8712);
   U14244 : XNOR2_X1 port map( A => n8687, B => n8952, ZN => n8688);
   U14245 : XNOR2_X1 port map( A => n8689, B => n8688, ZN => n8695);
   U14246 : XNOR2_X1 port map( A => n9139, B => n8690, ZN => n8693);
   U14247 : XNOR2_X1 port map( A => n8691, B => n2747, ZN => n8692);
   U14248 : XNOR2_X1 port map( A => n8693, B => n8692, ZN => n8694);
   U14250 : INV_X1 port map( A => n9980, ZN => n9984);
   U14251 : XNOR2_X1 port map( A => n8698, B => n8962, ZN => n8701);
   U14252 : XNOR2_X1 port map( A => n8699, B => n1364, ZN => n8700);
   U14253 : XNOR2_X1 port map( A => n8701, B => n8700, ZN => n8702);
   U14254 : MUX2_X1 port map( A => n9984, B => n9982, S => n9981, Z => n8711);
   U14255 : INV_X1 port map( A => n8703, ZN => n8705);
   U14256 : XNOR2_X1 port map( A => n8704, B => n8705, ZN => n8710);
   U14257 : XNOR2_X1 port map( A => n8897, B => n8706, ZN => n8708);
   U14258 : XNOR2_X1 port map( A => n9044, B => n2970, ZN => n8707);
   U14259 : XOR2_X1 port map( A => n8708, B => n8707, Z => n8709);
   U14260 : XNOR2_X2 port map( A => n8710, B => n8709, ZN => n9985);
   U14262 : XNOR2_X1 port map( A => n8714, B => n8713, ZN => n8718);
   U14263 : XNOR2_X1 port map( A => n8867, B => n1815, ZN => n8716);
   U14264 : XNOR2_X1 port map( A => n8716, B => n8715, ZN => n8717);
   U14265 : XNOR2_X1 port map( A => n8720, B => n8719, ZN => n8724);
   U14266 : XNOR2_X1 port map( A => n8723, B => n8724, ZN => n10069);
   U14267 : NOR2_X1 port map( A1 => n427, A2 => n25457, ZN => n9232);
   U14268 : INV_X1 port map( A => n10069, ZN => n10075);
   U14269 : XNOR2_X1 port map( A => n8726, B => n8725, ZN => n8729);
   U14270 : XNOR2_X1 port map( A => n8760, B => n812, ZN => n8727);
   U14271 : XNOR2_X1 port map( A => n9042, B => n8727, ZN => n8728);
   U14272 : XNOR2_X1 port map( A => n8729, B => n8728, ZN => n8744);
   U14273 : INV_X1 port map( A => n8744, ZN => n9620);
   U14274 : XNOR2_X1 port map( A => n8730, B => n8951, ZN => n8732);
   U14275 : XNOR2_X1 port map( A => n8731, B => n8732, ZN => n8736);
   U14276 : XNOR2_X1 port map( A => n9141, B => n2036, ZN => n8733);
   U14277 : XNOR2_X1 port map( A => n8734, B => n8733, ZN => n8735);
   U14278 : XNOR2_X1 port map( A => n8736, B => n8735, ZN => n10068);
   U14279 : INV_X1 port map( A => n10068, ZN => n9764);
   U14280 : OAI21_X1 port map( B1 => n10075, B2 => n9620, A => n9764, ZN => 
                           n8737);
   U14281 : NOR2_X1 port map( A1 => n9232, A2 => n8737, ZN => n8752);
   U14282 : NAND2_X1 port map( A1 => n427, A2 => n10068, ZN => n9766);
   U14283 : XNOR2_X1 port map( A => n8739, B => n8738, ZN => n8743);
   U14284 : XNOR2_X1 port map( A => n8965, B => n3084, ZN => n8740);
   U14285 : XNOR2_X1 port map( A => n8741, B => n8740, ZN => n8742);
   U14286 : XNOR2_X1 port map( A => n8746, B => n1804, ZN => n8747);
   U14287 : XOR2_X1 port map( A => n8748, B => n8747, Z => n8749);
   U14288 : NAND3_X1 port map( A1 => n1330, A2 => n10070, A3 => n9762, ZN => 
                           n8751);
   U14289 : XNOR2_X1 port map( A => n9191, B => n24445, ZN => n9050);
   U14290 : XNOR2_X1 port map( A => n9050, B => n8753, ZN => n8759);
   U14291 : XNOR2_X1 port map( A => n8754, B => n3183, ZN => n8757);
   U14292 : XNOR2_X1 port map( A => n8756, B => n8757, ZN => n8758);
   U14293 : XNOR2_X1 port map( A => n8759, B => n8758, ZN => n9419);
   U14294 : INV_X1 port map( A => n9419, ZN => n9617);
   U14295 : XNOR2_X1 port map( A => n9043, B => n8760, ZN => n8763);
   U14296 : INV_X1 port map( A => n173, ZN => n8761);
   U14297 : XNOR2_X1 port map( A => n8989, B => n8761, ZN => n8762);
   U14298 : XNOR2_X1 port map( A => n8763, B => n8762, ZN => n8768);
   U14299 : XNOR2_X1 port map( A => n9041, B => n8764, ZN => n8765);
   U14300 : XNOR2_X1 port map( A => n8766, B => n8765, ZN => n8767);
   U14301 : XNOR2_X1 port map( A => n8770, B => n8769, ZN => n9146);
   U14302 : XNOR2_X1 port map( A => n8771, B => n8772, ZN => n9000);
   U14303 : XNOR2_X1 port map( A => n9146, B => n9000, ZN => n8776);
   U14304 : XNOR2_X1 port map( A => n8964, B => n9057, ZN => n8774);
   U14305 : XNOR2_X1 port map( A => n8965, B => n1924, ZN => n8773);
   U14306 : XNOR2_X1 port map( A => n8774, B => n8773, ZN => n8775);
   U14307 : XNOR2_X1 port map( A => n8776, B => n8775, ZN => n9613);
   U14308 : MUX2_X1 port map( A => n9617, B => n25005, S => n9613, Z => n8804);
   U14309 : XNOR2_X1 port map( A => n8778, B => n8777, ZN => n8785);
   U14310 : XNOR2_X1 port map( A => n8779, B => n8780, ZN => n9154);
   U14311 : XNOR2_X1 port map( A => n8782, B => n8781, ZN => n8783);
   U14312 : XNOR2_X1 port map( A => n9154, B => n8783, ZN => n8784);
   U14313 : XNOR2_X1 port map( A => n8786, B => n3164, ZN => n8788);
   U14314 : XNOR2_X1 port map( A => n8788, B => n8787, ZN => n8792);
   U14315 : XNOR2_X1 port map( A => n8790, B => n8789, ZN => n9177);
   U14316 : INV_X1 port map( A => n9177, ZN => n8791);
   U14317 : XNOR2_X1 port map( A => n8791, B => n8792, ZN => n8794);
   U14318 : XNOR2_X1 port map( A => n8794, B => n8793, ZN => n9977);
   U14319 : INV_X1 port map( A => n9977, ZN => n9757);
   U14320 : XNOR2_X1 port map( A => n9137, B => n8797, ZN => n8802);
   U14321 : INV_X1 port map( A => n2240, ZN => n20864);
   U14322 : XNOR2_X1 port map( A => n8799, B => n20864, ZN => n8800);
   U14323 : XNOR2_X1 port map( A => n8997, B => n8800, ZN => n8801);
   U14324 : XNOR2_X1 port map( A => n8802, B => n8801, ZN => n9753);
   U14325 : INV_X1 port map( A => n9753, ZN => n9974);
   U14326 : NAND3_X1 port map( A1 => n9617, A2 => n9974, A3 => n25005, ZN => 
                           n8803);
   U14327 : XNOR2_X1 port map( A => n8805, B => n9089, ZN => n8811);
   U14328 : XNOR2_X1 port map( A => n9158, B => n1874, ZN => n8809);
   U14329 : XNOR2_X1 port map( A => n8806, B => n8807, ZN => n8808);
   U14330 : XNOR2_X1 port map( A => n8809, B => n8808, ZN => n8810);
   U14332 : INV_X1 port map( A => n8970, ZN => n9168);
   U14333 : XNOR2_X1 port map( A => n9168, B => n8812, ZN => n8815);
   U14334 : XNOR2_X1 port map( A => n8813, B => Key(172), ZN => n8814);
   U14335 : XNOR2_X1 port map( A => n8815, B => n8814, ZN => n8817);
   U14336 : XNOR2_X1 port map( A => n8873, B => n9096, ZN => n8816);
   U14337 : NAND2_X1 port map( A1 => n10020, A2 => n24495, ZN => n9732);
   U14338 : INV_X1 port map( A => n9732, ZN => n8842);
   U14339 : XNOR2_X1 port map( A => n8818, B => n4034, ZN => n8819);
   U14340 : XNOR2_X1 port map( A => n8858, B => n8819, ZN => n8823);
   U14341 : XNOR2_X1 port map( A => n8820, B => n9176, ZN => n8821);
   U14342 : XNOR2_X1 port map( A => n8821, B => n9115, ZN => n8822);
   U14343 : INV_X1 port map( A => n10018, ZN => n9730);
   U14344 : XNOR2_X1 port map( A => n8824, B => n9188, ZN => n8825);
   U14345 : XNOR2_X1 port map( A => n9101, B => n8825, ZN => n8830);
   U14346 : XNOR2_X1 port map( A => n8826, B => n23699, ZN => n8828);
   U14347 : XNOR2_X1 port map( A => n8828, B => n8827, ZN => n8829);
   U14348 : XNOR2_X1 port map( A => n8830, B => n8829, ZN => n8839);
   U14349 : XNOR2_X1 port map( A => n8951, B => n21703, ZN => n8832);
   U14350 : XNOR2_X1 port map( A => n8832, B => n8831, ZN => n8834);
   U14351 : XNOR2_X1 port map( A => n8833, B => n8834, ZN => n10019);
   U14352 : INV_X1 port map( A => n10019, ZN => n9320);
   U14353 : OAI211_X1 port map( C1 => n9729, C2 => n9730, A => n8839, B => 
                           n9320, ZN => n8841);
   U14354 : INV_X1 port map( A => n9729, ZN => n9493);
   U14355 : XNOR2_X1 port map( A => n8961, B => n1952, ZN => n8836);
   U14356 : XNOR2_X1 port map( A => n9111, B => n8836, ZN => n8837);
   U14357 : INV_X1 port map( A => n8839, ZN => n9731);
   U14358 : XNOR2_X1 port map( A => n8843, B => n8844, ZN => n8850);
   U14359 : XNOR2_X1 port map( A => n8846, B => n8845, ZN => n8848);
   U14360 : XNOR2_X1 port map( A => n8917, B => n2989, ZN => n8847);
   U14361 : XNOR2_X1 port map( A => n8848, B => n8847, ZN => n8849);
   U14362 : XNOR2_X1 port map( A => n8850, B => n8849, ZN => n9634);
   U14363 : XNOR2_X1 port map( A => n8852, B => n8851, ZN => n8857);
   U14364 : XNOR2_X1 port map( A => n8853, B => n921, ZN => n8854);
   U14365 : XNOR2_X1 port map( A => n8855, B => n8854, ZN => n8856);
   U14366 : XNOR2_X1 port map( A => n8857, B => n8856, ZN => n9435);
   U14368 : XNOR2_X1 port map( A => n8858, B => n8859, ZN => n8864);
   U14369 : XNOR2_X1 port map( A => n8860, B => n2745, ZN => n8861);
   U14370 : XNOR2_X1 port map( A => n8862, B => n8861, ZN => n8863);
   U14371 : XNOR2_X1 port map( A => n8864, B => n8863, ZN => n9711);
   U14372 : OR2_X1 port map( A1 => n10038, A2 => n9711, ZN => n8888);
   U14373 : XNOR2_X1 port map( A => n8866, B => n8865, ZN => n8871);
   U14374 : XNOR2_X1 port map( A => n8867, B => n899, ZN => n8869);
   U14375 : XNOR2_X1 port map( A => n8868, B => n8869, ZN => n8870);
   U14376 : XNOR2_X1 port map( A => n8873, B => n8872, ZN => n8879);
   U14377 : XNOR2_X1 port map( A => n8874, B => n24056, ZN => n8877);
   U14378 : XNOR2_X1 port map( A => n8875, B => n4189, ZN => n8876);
   U14379 : XNOR2_X1 port map( A => n8877, B => n8876, ZN => n8878);
   U14380 : XNOR2_X1 port map( A => n8879, B => n8878, ZN => n10037);
   U14381 : NOR2_X1 port map( A1 => n9635, A2 => n10037, ZN => n9228);
   U14382 : NAND2_X1 port map( A1 => n9228, A2 => n9713, ZN => n8887);
   U14383 : INV_X1 port map( A => n9634, ZN => n9718);
   U14384 : XNOR2_X1 port map( A => n8880, B => n1854, ZN => n8881);
   U14385 : XNOR2_X1 port map( A => n8883, B => n8882, ZN => n8885);
   U14387 : INV_X1 port map( A => n9433, ZN => n9710);
   U14388 : INV_X1 port map( A => n9090, ZN => n8890);
   U14389 : XNOR2_X1 port map( A => n8890, B => n8889, ZN => n8895);
   U14390 : XNOR2_X1 port map( A => n9034, B => n25235, ZN => n8893);
   U14391 : XNOR2_X1 port map( A => n8891, B => n2805, ZN => n8892);
   U14392 : XNOR2_X1 port map( A => n8893, B => n8892, ZN => n8894);
   U14393 : XNOR2_X1 port map( A => n8897, B => n8896, ZN => n9098);
   U14394 : XNOR2_X1 port map( A => n8899, B => n8898, ZN => n8986);
   U14395 : XNOR2_X1 port map( A => n9098, B => n8986, ZN => n8905);
   U14396 : XNOR2_X1 port map( A => n25228, B => n8987, ZN => n8903);
   U14398 : XNOR2_X1 port map( A => n24056, B => n24280, ZN => n8902);
   U14399 : XNOR2_X1 port map( A => n8903, B => n8902, ZN => n8904);
   U14400 : XNOR2_X2 port map( A => n8905, B => n8904, ZN => n9990);
   U14401 : INV_X1 port map( A => n9990, ZN => n9996);
   U14402 : XNOR2_X1 port map( A => n9058, B => n1726, ZN => n8906);
   U14403 : XNOR2_X1 port map( A => n8907, B => n8906, ZN => n8912);
   U14404 : XNOR2_X1 port map( A => n8908, B => n8909, ZN => n8910);
   U14405 : XNOR2_X1 port map( A => n9110, B => n8910, ZN => n8911);
   U14406 : XNOR2_X1 port map( A => n8913, B => n8914, ZN => n8915);
   U14407 : XNOR2_X1 port map( A => n9122, B => n8915, ZN => n8921);
   U14408 : XNOR2_X1 port map( A => n9081, B => n8916, ZN => n8919);
   U14409 : XNOR2_X1 port map( A => n8917, B => n21964, ZN => n8918);
   U14410 : XNOR2_X1 port map( A => n8919, B => n8918, ZN => n8920);
   U14411 : XNOR2_X1 port map( A => n8921, B => n8920, ZN => n9658);
   U14412 : INV_X1 port map( A => n9658, ZN => n9745);
   U14413 : AOI21_X1 port map( B1 => n9745, B2 => n9989, A => n9990, ZN => 
                           n9316);
   U14414 : XNOR2_X1 port map( A => n8922, B => n9011, ZN => n8927);
   U14415 : XNOR2_X1 port map( A => n9075, B => n21742, ZN => n8924);
   U14416 : XNOR2_X1 port map( A => n8924, B => n8923, ZN => n8925);
   U14417 : XNOR2_X1 port map( A => n9010, B => n8925, ZN => n8926);
   U14418 : XNOR2_X1 port map( A => n8926, B => n8927, ZN => n9423);
   U14419 : XNOR2_X1 port map( A => n9102, B => n9020, ZN => n8932);
   U14420 : XNOR2_X1 port map( A => n8928, B => n8880, ZN => n8930);
   U14421 : XNOR2_X1 port map( A => n8935, B => n3152, ZN => n8929);
   U14422 : XNOR2_X1 port map( A => n8930, B => n8929, ZN => n8931);
   U14423 : XNOR2_X2 port map( A => n8932, B => n8931, ZN => n9991);
   U14424 : OAI211_X1 port map( C1 => n25444, C2 => n9990, A => n9657, B => 
                           n9747, ZN => n8933);
   U14425 : OAI21_X1 port map( B1 => n9425, B2 => n9316, A => n8933, ZN => 
                           n11519);
   U14426 : INV_X1 port map( A => n25060, ZN => n10384);
   U14427 : XNOR2_X1 port map( A => n8935, B => n2049, ZN => n8936);
   U14428 : XNOR2_X1 port map( A => n8940, B => n8941, ZN => n8944);
   U14429 : XNOR2_X1 port map( A => n9176, B => n1870, ZN => n8942);
   U14430 : XNOR2_X1 port map( A => n9011, B => n8942, ZN => n8943);
   U14431 : XNOR2_X1 port map( A => n9158, B => n1951, ZN => n8946);
   U14432 : XNOR2_X1 port map( A => n8946, B => n25235, ZN => n8948);
   U14433 : XNOR2_X1 port map( A => n8948, B => n8947, ZN => n8949);
   U14434 : INV_X1 port map( A => n9550, ZN => n9682);
   U14435 : MUX2_X1 port map( A => n260, B => n10046, S => n9682, Z => n8979);
   U14436 : XNOR2_X1 port map( A => n8952, B => n8951, ZN => n8954);
   U14437 : XNOR2_X1 port map( A => n8954, B => n8953, ZN => n8958);
   U14438 : XNOR2_X1 port map( A => n9139, B => n3093, ZN => n8956);
   U14439 : XNOR2_X1 port map( A => n8956, B => n8955, ZN => n8957);
   U14440 : XNOR2_X1 port map( A => n8960, B => n8959, ZN => n8963);
   U14441 : XNOR2_X1 port map( A => n8962, B => n8961, ZN => n9144);
   U14442 : XNOR2_X1 port map( A => n9144, B => n8963, ZN => n8969);
   U14443 : XNOR2_X1 port map( A => n9059, B => n8964, ZN => n8967);
   U14444 : XNOR2_X1 port map( A => n8965, B => n2717, ZN => n8966);
   U14445 : XNOR2_X1 port map( A => n8967, B => n8966, ZN => n8968);
   U14446 : XNOR2_X1 port map( A => n8969, B => n8968, ZN => n10045);
   U14447 : INV_X1 port map( A => n10045, ZN => n9627);
   U14448 : AND2_X1 port map( A1 => n261, A2 => n9627, ZN => n9684);
   U14449 : XNOR2_X1 port map( A => n8970, B => n765, ZN => n8972);
   U14450 : XNOR2_X1 port map( A => n8971, B => n8972, ZN => n8975);
   U14451 : XNOR2_X1 port map( A => n8987, B => n8973, ZN => n8974);
   U14452 : XNOR2_X1 port map( A => n8975, B => n8974, ZN => n8976);
   U14453 : MUX2_X2 port map( A => n8979, B => n8978, S => n9681, Z => n11038);
   U14454 : INV_X1 port map( A => n11038, ZN => n10570);
   U14455 : XNOR2_X1 port map( A => n8985, B => n8986, ZN => n8993);
   U14456 : XNOR2_X1 port map( A => n8987, B => n8988, ZN => n8991);
   U14457 : XNOR2_X1 port map( A => n8989, B => n24287, ZN => n8990);
   U14458 : XNOR2_X1 port map( A => n8991, B => n8990, ZN => n8992);
   U14459 : INV_X1 port map( A => n9696, ZN => n9699);
   U14460 : XNOR2_X1 port map( A => n8994, B => n8995, ZN => n8999);
   U14461 : XNOR2_X1 port map( A => n8997, B => n8996, ZN => n8998);
   U14462 : XNOR2_X1 port map( A => n8998, B => n8999, ZN => n10029);
   U14463 : INV_X1 port map( A => n10029, ZN => n9695);
   U14464 : XNOR2_X1 port map( A => n9000, B => n9001, ZN => n9006);
   U14465 : XNOR2_X1 port map( A => n9002, B => n2795, ZN => n9004);
   U14466 : XNOR2_X1 port map( A => n9003, B => n9004, ZN => n9005);
   U14467 : NOR2_X1 port map( A1 => n9639, A2 => n24332, ZN => n10028);
   U14468 : XNOR2_X1 port map( A => n9007, B => n2882, ZN => n9008);
   U14469 : XNOR2_X1 port map( A => n9010, B => n9009, ZN => n9014);
   U14470 : XNOR2_X1 port map( A => n9012, B => n9011, ZN => n9013);
   U14471 : INV_X1 port map( A => n9016, ZN => n9017);
   U14472 : XNOR2_X1 port map( A => n9018, B => n9017, ZN => n9019);
   U14473 : INV_X1 port map( A => n10026, ZN => n9022);
   U14474 : OAI211_X1 port map( C1 => n9699, C2 => n10027, A => n10031, B => 
                           n9022, ZN => n9023);
   U14475 : OAI21_X1 port map( B1 => n9565, B2 => n9563, A => n9024, ZN => 
                           n9026);
   U14476 : OAI21_X1 port map( B1 => n9454, B2 => n9885, A => n9567, ZN => 
                           n9025);
   U14477 : AOI21_X1 port map( B1 => n10570, B2 => n10944, A => n10942, ZN => 
                           n9131);
   U14478 : NAND3_X1 port map( A1 => n4993, A2 => n9872, A3 => n9875, ZN => 
                           n9031);
   U14479 : NAND2_X1 port map( A1 => n9694, A2 => n9028, ZN => n9030);
   U14480 : NAND3_X1 port map( A1 => n9875, A2 => n307, A3 => n9251, ZN => 
                           n9029);
   U14482 : XNOR2_X1 port map( A => n9033, B => n9154, ZN => n9039);
   U14483 : XNOR2_X1 port map( A => n9035, B => n1792, ZN => n9036);
   U14484 : XNOR2_X1 port map( A => n9037, B => n9036, ZN => n9038);
   U14485 : XNOR2_X1 port map( A => n9040, B => n9041, ZN => n9164);
   U14486 : XNOR2_X1 port map( A => n9164, B => n9042, ZN => n9049);
   U14487 : XNOR2_X1 port map( A => n9043, B => n62, ZN => n9047);
   U14488 : XNOR2_X1 port map( A => n25228, B => n9044, ZN => n9046);
   U14489 : XNOR2_X1 port map( A => n9047, B => n9046, ZN => n9048);
   U14490 : XNOR2_X1 port map( A => n9049, B => n9048, ZN => n9244);
   U14492 : XNOR2_X1 port map( A => n9051, B => n9050, ZN => n9056);
   U14493 : XNOR2_X1 port map( A => n8880, B => n2903, ZN => n9053);
   U14494 : XNOR2_X1 port map( A => n9054, B => n9053, ZN => n9055);
   U14495 : NAND2_X1 port map( A1 => n10058, A2 => n24092, ZN => n9063);
   U14496 : XNOR2_X1 port map( A => n9058, B => n9057, ZN => n9061);
   U14497 : XNOR2_X1 port map( A => n9059, B => n1801, ZN => n9060);
   U14498 : XNOR2_X2 port map( A => n9062, B => n5743, ZN => n10053);
   U14499 : XNOR2_X1 port map( A => n9065, B => n9177, ZN => n9079);
   U14500 : MUX2_X1 port map( A => n9068, B => n9067, S => n9066, Z => n9072);
   U14501 : OAI211_X1 port map( C1 => n9072, C2 => n9071, A => n9070, B => 
                           n9069, ZN => n9074);
   U14502 : XNOR2_X1 port map( A => n9074, B => n9073, ZN => n9077);
   U14503 : XNOR2_X1 port map( A => n9075, B => n2044, ZN => n9076);
   U14504 : XNOR2_X1 port map( A => n9077, B => n9076, ZN => n9078);
   U14505 : XNOR2_X1 port map( A => n9137, B => n9080, ZN => n9085);
   U14506 : XNOR2_X1 port map( A => n9081, B => n9141, ZN => n9084);
   U14507 : XNOR2_X1 port map( A => n9082, B => n2782, ZN => n9083);
   U14508 : MUX2_X1 port map( A => n9539, B => n9086, S => n9244, Z => n9087);
   U14509 : XNOR2_X1 port map( A => n9089, B => n9090, ZN => n9094);
   U14510 : XNOR2_X1 port map( A => n8069, B => n1835, ZN => n9091);
   U14511 : XNOR2_X1 port map( A => n9092, B => n9091, ZN => n9093);
   U14512 : XNOR2_X1 port map( A => n9096, B => n9095, ZN => n9100);
   U14513 : XNOR2_X1 port map( A => n9169, B => n1920, ZN => n9097);
   U14514 : XNOR2_X1 port map( A => n9098, B => n9097, ZN => n9099);
   U14515 : XNOR2_X1 port map( A => n9100, B => n9099, ZN => n9218);
   U14516 : NAND2_X1 port map( A1 => n10060, A2 => n10065, ZN => n9703);
   U14517 : XNOR2_X1 port map( A => n9102, B => n9101, ZN => n9105);
   U14518 : XNOR2_X1 port map( A => n9189, B => n3073, ZN => n9103);
   U14519 : XNOR2_X1 port map( A => n8297, B => n9103, ZN => n9104);
   U14520 : XNOR2_X1 port map( A => n9106, B => n9107, ZN => n9109);
   U14521 : XNOR2_X1 port map( A => n9149, B => n2208, ZN => n9108);
   U14522 : XNOR2_X1 port map( A => n9109, B => n9108, ZN => n9113);
   U14523 : XNOR2_X1 port map( A => n9110, B => n9111, ZN => n9112);
   U14524 : NAND2_X1 port map( A1 => n9127, A2 => n9704, ZN => n9120);
   U14525 : XNOR2_X1 port map( A => n9179, B => n2477, ZN => n9116);
   U14526 : XNOR2_X1 port map( A => n9117, B => n9116, ZN => n9118);
   U14527 : XNOR2_X1 port map( A => n9119, B => n9118, ZN => n10061);
   U14528 : AOI21_X1 port map( B1 => n9703, B2 => n9120, A => n309, ZN => n9129
                           );
   U14529 : XNOR2_X1 port map( A => n9121, B => n2991, ZN => n9123);
   U14530 : XNOR2_X1 port map( A => n9122, B => n9123, ZN => n9126);
   U14531 : XNOR2_X1 port map( A => n9125, B => n9126, ZN => n10063);
   U14533 : INV_X1 port map( A => n9460, ZN => n9919);
   U14534 : INV_X1 port map( A => n9459, ZN => n9271);
   U14535 : INV_X1 port map( A => n9918, ZN => n9914);
   U14536 : INV_X1 port map( A => n9463, ZN => n9916);
   U14538 : NOR2_X1 port map( A1 => n10583, A2 => n10371, ZN => n9210);
   U14539 : XNOR2_X1 port map( A => n9140, B => n9139, ZN => n9143);
   U14542 : INV_X1 port map( A => n9144, ZN => n9145);
   U14543 : XNOR2_X1 port map( A => n9145, B => n9146, ZN => n9153);
   U14544 : XNOR2_X1 port map( A => n9147, B => n8484, ZN => n9151);
   U14545 : XNOR2_X1 port map( A => n9149, B => n1865, ZN => n9150);
   U14546 : XNOR2_X1 port map( A => n9151, B => n9150, ZN => n9152);
   U14547 : INV_X1 port map( A => n24025, ZN => n10140);
   U14548 : NOR2_X1 port map( A1 => n10146, A2 => n10140, ZN => n9187);
   U14549 : INV_X1 port map( A => n9154, ZN => n9157);
   U14550 : XNOR2_X1 port map( A => n9155, B => n8069, ZN => n9156);
   U14551 : XNOR2_X1 port map( A => n9157, B => n9156, ZN => n9163);
   U14552 : XNOR2_X1 port map( A => n9159, B => n9158, ZN => n9161);
   U14553 : XNOR2_X1 port map( A => n8278, B => n2726, ZN => n9160);
   U14554 : XNOR2_X1 port map( A => n9161, B => n9160, ZN => n9162);
   U14555 : INV_X1 port map( A => n9164, ZN => n9166);
   U14556 : XNOR2_X1 port map( A => n9165, B => n9166, ZN => n9173);
   U14557 : XNOR2_X1 port map( A => n9167, B => n9168, ZN => n9171);
   U14558 : XNOR2_X1 port map( A => n9169, B => n1746, ZN => n9170);
   U14559 : XNOR2_X1 port map( A => n9171, B => n9170, ZN => n9172);
   U14562 : INV_X1 port map( A => n9174, ZN => n9397);
   U14563 : XNOR2_X1 port map( A => n9175, B => n9176, ZN => n9178);
   U14564 : XNOR2_X1 port map( A => n9177, B => n9178, ZN => n9186);
   U14565 : INV_X1 port map( A => n9179, ZN => n9180);
   U14566 : XNOR2_X1 port map( A => n9181, B => n9180, ZN => n9184);
   U14567 : INV_X1 port map( A => n22986, ZN => n20805);
   U14568 : XNOR2_X1 port map( A => n9182, B => n20805, ZN => n9183);
   U14569 : XNOR2_X1 port map( A => n9184, B => n9183, ZN => n9185);
   U14570 : XNOR2_X1 port map( A => n9186, B => n9185, ZN => n9820);
   U14571 : XNOR2_X1 port map( A => n9189, B => n9188, ZN => n9193);
   U14572 : XNOR2_X1 port map( A => n9190, B => n9191, ZN => n9192);
   U14573 : XNOR2_X1 port map( A => n9193, B => n9192, ZN => n9200);
   U14574 : XNOR2_X1 port map( A => n9194, B => n24445, ZN => n9198);
   U14575 : XNOR2_X1 port map( A => n9196, B => n5131, ZN => n9197);
   U14576 : XNOR2_X1 port map( A => n9198, B => n9197, ZN => n9199);
   U14578 : NOR2_X1 port map( A1 => n10584, A2 => n10585, ZN => n9209);
   U14579 : INV_X1 port map( A => n25216, ZN => n9928);
   U14580 : NAND2_X1 port map( A1 => n9930, A2 => n9928, ZN => n9208);
   U14581 : INV_X1 port map( A => n9345, ZN => n9600);
   U14586 : NAND2_X1 port map( A1 => n2565, A2 => n10254, ZN => n10252);
   U14587 : NAND2_X1 port map( A1 => n10250, A2 => n9372, ZN => n9213);
   U14589 : INV_X1 port map( A => n9218, ZN => n9705);
   U14590 : NAND2_X1 port map( A1 => n309, A2 => n9705, ZN => n9219);
   U14591 : NAND2_X1 port map( A1 => n9221, A2 => n9985, ZN => n9225);
   U14592 : NAND3_X1 port map( A1 => n9984, A2 => n9742, A3 => n9981, ZN => 
                           n9223);
   U14593 : OAI21_X1 port map( B1 => n9664, B2 => n9982, A => n9736, ZN => 
                           n9222);
   U14594 : NOR2_X1 port map( A1 => n9635, A2 => n9435, ZN => n9227);
   U14595 : INV_X1 port map( A => n10037, ZN => n9633);
   U14596 : NOR2_X1 port map( A1 => n9634, A2 => n9633, ZN => n9226);
   U14597 : MUX2_X1 port map( A => n9227, B => n9226, S => n9433, Z => n9230);
   U14598 : INV_X1 port map( A => n9228, ZN => n9229);
   U14599 : INV_X1 port map( A => n9435, ZN => n9709);
   U14600 : MUX2_X1 port map( A => n9231, B => n10068, S => n10075, Z => n9235)
                           ;
   U14601 : INV_X1 port map( A => n9232, ZN => n9234);
   U14602 : AOI21_X1 port map( B1 => n427, B2 => n10072, A => n9620, ZN => 
                           n9233);
   U14604 : INV_X1 port map( A => n10848, ZN => n11125);
   U14605 : INV_X1 port map( A => n10027, ZN => n9240);
   U14606 : AOI21_X1 port map( B1 => n9697, B2 => n10026, A => n10029, ZN => 
                           n9238);
   U14607 : OR2_X1 port map( A1 => n9238, A2 => n9639, ZN => n9239);
   U14608 : NAND2_X1 port map( A1 => n11121, A2 => n11123, ZN => n10847);
   U14609 : INV_X1 port map( A => n10847, ZN => n9241);
   U14610 : NAND2_X1 port map( A1 => n24446, A2 => n10050, ZN => n9867);
   U14611 : INV_X1 port map( A => n9245, ZN => n9246);
   U14612 : INV_X1 port map( A => n9564, ZN => n9456);
   U14613 : INV_X1 port map( A => n9565, ZN => n9883);
   U14614 : NAND2_X1 port map( A1 => n9883, A2 => n9885, ZN => n9249);
   U14615 : MUX2_X1 port map( A => n9249, B => n9248, S => n9887, Z => n9250);
   U14616 : INV_X1 port map( A => n9255, ZN => n9628);
   U14617 : AOI22_X1 port map( A1 => n9682, A2 => n9681, B1 => n9628, B2 => 
                           n10045, ZN => n9257);
   U14618 : NAND2_X1 port map( A1 => n261, A2 => n9681, ZN => n9256);
   U14619 : MUX2_X1 port map( A => n9257, B => n9256, S => n10046, Z => n9258);
   U14620 : INV_X1 port map( A => n10740, ZN => n10856);
   U14621 : NAND2_X1 port map( A1 => n10856, A2 => n10861, ZN => n10743);
   U14622 : INV_X1 port map( A => n9864, ZN => n9559);
   U14623 : INV_X1 port map( A => n9554, ZN => n9860);
   U14624 : INV_X1 port map( A => n9560, ZN => n9858);
   U14625 : NAND2_X1 port map( A1 => n9857, A2 => n9860, ZN => n9260);
   U14626 : INV_X1 port map( A => n9856, ZN => n9474);
   U14627 : NAND2_X1 port map( A1 => n9474, A2 => n9858, ZN => n9259);
   U14628 : MUX2_X1 port map( A => n9260, B => n9259, S => n9864, Z => n9261);
   U14629 : NAND3_X1 port map( A1 => n10740, A2 => n10737, A3 => n10858, ZN => 
                           n9267);
   U14630 : AOI21_X1 port map( B1 => n9942, B2 => n25021, A => n227, ZN => 
                           n9265);
   U14631 : NOR2_X1 port map( A1 => n9893, A2 => n9943, ZN => n9263);
   U14632 : OAI21_X1 port map( B1 => n9289, B2 => n9263, A => n9897, ZN => 
                           n9264);
   U14633 : AND2_X1 port map( A1 => n25229, A2 => n10737, ZN => n10862);
   U14634 : NAND2_X1 port map( A1 => n10862, A2 => n10190, ZN => n9266);
   U14635 : NAND4_X2 port map( A1 => n9268, A2 => n9266, A3 => n10743, A4 => 
                           n9267, ZN => n12364);
   U14636 : XNOR2_X1 port map( A => n12364, B => n12089, ZN => n11734);
   U14638 : INV_X1 port map( A => n9269, ZN => n9952);
   U14639 : INV_X1 port map( A => n9388, ZN => n9948);
   U14640 : OAI21_X1 port map( B1 => n9389, B2 => n9388, A => n9952, ZN => 
                           n9270);
   U14641 : INV_X1 port map( A => n10192, ZN => n10831);
   U14642 : INV_X1 port map( A => n9462, ZN => n9354);
   U14643 : NAND2_X1 port map( A1 => n9354, A2 => n9459, ZN => n9458);
   U14644 : NAND3_X1 port map( A1 => n9354, A2 => n9271, A3 => n9461, ZN => 
                           n9273);
   U14645 : NAND3_X1 port map( A1 => n24944, A2 => n9271, A3 => n9355, ZN => 
                           n9272);
   U14646 : NAND4_X1 port map( A1 => n9275, A2 => n9274, A3 => n9273, A4 => 
                           n9272, ZN => n10277);
   U14647 : AND2_X1 port map( A1 => n10277, A2 => n10831, ZN => n10834);
   U14648 : INV_X1 port map( A => n9449, ZN => n9906);
   U14649 : INV_X1 port map( A => n9907, ZN => n9904);
   U14650 : MUX2_X1 port map( A => n9906, B => n9904, S => n9276, Z => n9278);
   U14651 : MUX2_X1 port map( A => n9939, B => n9276, S => n9905, Z => n9277);
   U14652 : NAND2_X1 port map( A1 => n10834, A2 => n9279, ZN => n9293);
   U14653 : INV_X1 port map( A => n9857, ZN => n9555);
   U14654 : NAND2_X1 port map( A1 => n9555, A2 => n9558, ZN => n9280);
   U14655 : NAND3_X1 port map( A1 => n3292, A2 => n9468, A3 => n9964, ZN => 
                           n9284);
   U14656 : NAND2_X1 port map( A1 => n9469, A2 => n9468, ZN => n9282);
   U14657 : INV_X1 port map( A => n9944, ZN => n9285);
   U14658 : OAI22_X1 port map( A1 => n9288, A2 => n9287, B1 => n9286, B2 => 
                           n227, ZN => n9290);
   U14659 : NOR2_X2 port map( A1 => n9290, A2 => n9289, ZN => n10518);
   U14661 : INV_X1 port map( A => n10275, ZN => n10833);
   U14662 : OAI22_X1 port map( A1 => n10090, A2 => n24505, B1 => n9295, B2 => 
                           n25454, ZN => n9296);
   U14664 : AND2_X1 port map( A1 => n9781, A2 => n10093, ZN => n9498);
   U14665 : NOR2_X1 port map( A1 => n9652, A2 => n9299, ZN => n9653);
   U14666 : NOR2_X1 port map( A1 => n9725, A2 => n25043, ZN => n9300);
   U14667 : MUX2_X1 port map( A => n9653, B => n9300, S => n10008, Z => n9304);
   U14668 : INV_X1 port map( A => n10007, ZN => n9721);
   U14669 : MUX2_X1 port map( A => n9721, B => n10008, S => n9301, Z => n9302);
   U14670 : NOR2_X1 port map( A1 => n9302, A2 => n2922, ZN => n9303);
   U14673 : INV_X1 port map( A => n10080, ZN => n9326);
   U14674 : NAND3_X1 port map( A1 => n4256, A2 => n10079, A3 => n9306, ZN => 
                           n9308);
   U14675 : NAND4_X1 port map( A1 => n9309, A2 => n10087, A3 => n9308, A4 => 
                           n9307, ZN => n11130);
   U14676 : OAI21_X1 port map( B1 => n9796, B2 => n8521, A => n1796, ZN => 
                           n9313);
   U14677 : NAND2_X1 port map( A1 => n9671, A2 => n246, ZN => n9668);
   U14678 : INV_X1 port map( A => n10714, ZN => n10839);
   U14679 : OAI21_X1 port map( B1 => n9657, B2 => n9747, A => n9745, ZN => 
                           n9315);
   U14680 : NAND2_X1 port map( A1 => n9315, A2 => n24534, ZN => n9317);
   U14681 : NOR2_X1 port map( A1 => n10019, A2 => n25475, ZN => n9319);
   U14682 : NOR2_X1 port map( A1 => n9729, A2 => n24495, ZN => n9318);
   U14684 : MUX2_X1 port map( A => n9319, B => n9318, S => n25007, Z => n9323);
   U14685 : NAND2_X1 port map( A1 => n10020, A2 => n9731, ZN => n9321);
   U14687 : AOI21_X1 port map( B1 => n9321, B2 => n10015, A => n9320, ZN => 
                           n9322);
   U14688 : INV_X1 port map( A => n10470, ZN => n11129);
   U14689 : XNOR2_X1 port map( A => n24328, B => n11356, ZN => n9409);
   U14690 : OAI21_X1 port map( B1 => n4256, B2 => n9507, A => n9326, ZN => 
                           n9325);
   U14693 : NOR2_X1 port map( A1 => n9774, A2 => n4254, ZN => n9329);
   U14694 : INV_X1 port map( A => n9773, ZN => n9503);
   U14698 : INV_X1 port map( A => n10113, ZN => n9529);
   U14699 : NAND2_X1 port map( A1 => n9529, A2 => n8523, ZN => n9336);
   U14700 : INV_X1 port map( A => n9805, ZN => n10112);
   U14701 : MUX2_X1 port map( A => n9336, B => n9335, S => n10112, Z => n10873)
                           ;
   U14702 : NOR2_X1 port map( A1 => n9806, A2 => n9530, ZN => n9337);
   U14703 : INV_X1 port map( A => n9845, ZN => n10156);
   U14708 : AND2_X1 port map( A1 => n9384, A2 => n10161, ZN => n10159);
   U14709 : OAI21_X1 port map( B1 => n10159, B2 => n9349, A => n3305, ZN => 
                           n9350);
   U14712 : NOR2_X1 port map( A1 => n9950, A2 => n9951, ZN => n9363);
   U14713 : NAND2_X1 port map( A1 => n9389, A2 => n9388, ZN => n9362);
   U14714 : NAND2_X1 port map( A1 => n9955, A2 => n9951, ZN => n9359);
   U14715 : NAND2_X1 port map( A1 => n9360, A2 => n9359, ZN => n9361);
   U14716 : INV_X1 port map( A => n9365, ZN => n9368);
   U14719 : NAND2_X1 port map( A1 => n9365, A2 => n24025, ZN => n9366);
   U14720 : INV_X1 port map( A => n10137, ZN => n10134);
   U14721 : NAND3_X1 port map( A1 => n9368, A2 => n25463, A3 => n10136, ZN => 
                           n9369);
   U14722 : OR2_X1 port map( A1 => n9380, A2 => n10128, ZN => n9373);
   U14723 : INV_X1 port map( A => n10129, ZN => n10132);
   U14724 : NAND2_X1 port map( A1 => n10756, A2 => n10757, ZN => n9374);
   U14725 : INV_X1 port map( A => n12249, ZN => n9376);
   U14726 : XNOR2_X1 port map( A => n25090, B => n9376, ZN => n9407);
   U14727 : NAND2_X1 port map( A1 => n9378, A2 => n9377, ZN => n9381);
   U14728 : INV_X1 port map( A => n10729, ZN => n10731);
   U14729 : NOR2_X1 port map( A1 => n3305, A2 => n10157, ZN => n9383);
   U14730 : INV_X1 port map( A => n10175, ZN => n9585);
   U14731 : NAND2_X1 port map( A1 => n9830, A2 => n9585, ZN => n9386);
   U14732 : NAND2_X1 port map( A1 => n9387, A2 => n9947, ZN => n9391);
   U14733 : NOR2_X1 port map( A1 => n9950, A2 => n9388, ZN => n9390);
   U14734 : INV_X1 port map( A => n10734, ZN => n10271);
   U14735 : INV_X1 port map( A => n9603, ZN => n9926);
   U14736 : OAI211_X1 port map( C1 => n9926, C2 => n9604, A => n9600, B => 
                           n9934, ZN => n9396);
   U14737 : NAND2_X1 port map( A1 => n25217, A2 => n9604, ZN => n9395);
   U14738 : NAND3_X1 port map( A1 => n9925, A2 => n24084, A3 => n9599, ZN => 
                           n9394);
   U14739 : NAND3_X1 port map( A1 => n10271, A2 => n4951, A3 => n10482, ZN => 
                           n9405);
   U14740 : INV_X1 port map( A => n9398, ZN => n10142);
   U14741 : NAND3_X1 port map( A1 => n10146, A2 => n10142, A3 => n10134, ZN => 
                           n9399);
   U14742 : OAI21_X1 port map( B1 => n9174, B2 => n10140, A => n9399, ZN => 
                           n9402);
   U14743 : NOR2_X1 port map( A1 => n10142, A2 => n24026, ZN => n9400);
   U14744 : AOI21_X1 port map( B1 => n10291, B2 => n10757, A => n10753, ZN => 
                           n9410);
   U14745 : NAND2_X1 port map( A1 => n9760, A2 => n427, ZN => n9412);
   U14746 : AOI21_X1 port map( B1 => n9704, B2 => n429, A => n10063, ZN => 
                           n9414);
   U14747 : NAND2_X1 port map( A1 => n9417, A2 => n9416, ZN => n9422);
   U14748 : NAND2_X1 port map( A1 => n9418, A2 => n9754, ZN => n9421);
   U14749 : NAND2_X1 port map( A1 => n9617, A2 => n9753, ZN => n9751);
   U14750 : AND2_X1 port map( A1 => n9972, A2 => n9752, ZN => n9420);
   U14751 : NAND2_X1 port map( A1 => n11084, A2 => n10890, ZN => n9428);
   U14752 : NOR2_X1 port map( A1 => n9991, A2 => n9747, ZN => n9424);
   U14753 : OAI21_X1 port map( B1 => n9425, B2 => n9424, A => n9746, ZN => 
                           n9427);
   U14754 : AND2_X1 port map( A1 => n9423, A2 => n9990, ZN => n9993);
   U14755 : OAI21_X1 port map( B1 => n9993, B2 => n9745, A => n9991, ZN => 
                           n9426);
   U14756 : NAND2_X1 port map( A1 => n9427, A2 => n9426, ZN => n10889);
   U14757 : AOI21_X1 port map( B1 => n11082, B2 => n9428, A => n418, ZN => 
                           n9439);
   U14758 : INV_X1 port map( A => n9985, ZN => n9978);
   U14759 : NAND2_X1 port map( A1 => n10890, A2 => n418, ZN => n10441);
   U14760 : INV_X1 port map( A => n9635, ZN => n9434);
   U14761 : INV_X1 port map( A => n10439, ZN => n9437);
   U14762 : OAI22_X1 port map( A1 => n10891, A2 => n10441, B1 => n9437, B2 => 
                           n10767, ZN => n9438);
   U14763 : XNOR2_X1 port map( A => n11295, B => n12108, ZN => n9480);
   U14765 : AND2_X1 port map( A1 => n10375, A2 => n10584, ZN => n10589);
   U14766 : NAND2_X1 port map( A1 => n10589, A2 => n10585, ZN => n9442);
   U14767 : NOR2_X1 port map( A1 => n10583, A2 => n10584, ZN => n9440);
   U14768 : NAND2_X1 port map( A1 => n10590, A2 => n9440, ZN => n9441);
   U14769 : MUX2_X1 port map( A => n25021, B => n9946, S => n9945, Z => n9448);
   U14770 : NOR2_X1 port map( A1 => n9899, A2 => n9944, ZN => n9446);
   U14771 : NOR2_X1 port map( A1 => n9446, A2 => n9445, ZN => n9447);
   U14772 : MUX2_X1 port map( A => n9908, B => n24511, S => n9904, Z => n9453);
   U14773 : INV_X1 port map( A => n9905, ZN => n9935);
   U14774 : NAND3_X1 port map( A1 => n9449, A2 => n24511, A3 => n9908, ZN => 
                           n9452);
   U14775 : INV_X1 port map( A => n9450, ZN => n9938);
   U14776 : NAND3_X1 port map( A1 => n9935, A2 => n9939, A3 => n9938, ZN => 
                           n9451);
   U14777 : INV_X1 port map( A => n9454, ZN => n9882);
   U14778 : INV_X1 port map( A => n25069, ZN => n9455);
   U14779 : NAND3_X1 port map( A1 => n9564, A2 => n9882, A3 => n9886, ZN => 
                           n9457);
   U14780 : OAI21_X1 port map( B1 => n9460, B2 => n9912, A => n9458, ZN => 
                           n9467);
   U14781 : AOI21_X1 port map( B1 => n9465, B2 => n9464, A => n9463, ZN => 
                           n9466);
   U14782 : NOR2_X1 port map( A1 => n3290, A2 => n9469, ZN => n9470);
   U14783 : NAND3_X1 port map( A1 => n24168, A2 => n24345, A3 => n10302, ZN => 
                           n9479);
   U14784 : NAND2_X1 port map( A1 => n9474, A2 => n239, ZN => n9473);
   U14785 : NAND3_X1 port map( A1 => n9558, A2 => n9560, A3 => n9860, ZN => 
                           n9475);
   U14786 : XNOR2_X1 port map( A => n9480, B => n11167, ZN => n9573);
   U14787 : OAI21_X1 port map( B1 => n25043, B2 => n9652, A => n9723, ZN => 
                           n9482);
   U14788 : NAND2_X1 port map( A1 => n9482, A2 => n9725, ZN => n9490);
   U14789 : NAND2_X1 port map( A1 => n9724, A2 => n10008, ZN => n9483);
   U14790 : NAND2_X1 port map( A1 => n9483, A2 => n9652, ZN => n9488);
   U14791 : NAND2_X1 port map( A1 => n9485, A2 => n9484, ZN => n9486);
   U14792 : OAI21_X1 port map( B1 => n9731, B2 => n426, A => n10019, ZN => 
                           n9494);
   U14794 : NOR2_X1 port map( A1 => n24505, A2 => n8571, ZN => n9497);
   U14795 : OR3_X1 port map( A1 => n9798, A2 => n9998, A3 => n8521, ZN => n9499
                           );
   U14796 : INV_X1 port map( A => n10775, ZN => n9502);
   U14797 : NOR2_X1 port map( A1 => n9797, A2 => n9671, ZN => n9501);
   U14798 : NOR2_X1 port map( A1 => n9775, A2 => n10104, ZN => n9504);
   U14799 : AOI22_X1 port map( A1 => n9504, A2 => n25393, B1 => n9775, B2 => 
                           n9503, ZN => n9505);
   U14800 : OAI21_X1 port map( B1 => n10080, B2 => n9786, A => n10079, ZN => 
                           n9506);
   U14801 : NAND3_X1 port map( A1 => n4256, A2 => n9507, A3 => n10082, ZN => 
                           n9508);
   U14802 : NAND2_X1 port map( A1 => n10100, A2 => n10099, ZN => n9514);
   U14803 : OAI21_X2 port map( B1 => n9517, B2 => n9518, A => n9516, ZN => 
                           n11298);
   U14804 : INV_X1 port map( A => n10176, ZN => n9831);
   U14805 : OAI211_X1 port map( C1 => n10186, C2 => n10178, A => n9831, B => 
                           n10175, ZN => n9519);
   U14806 : MUX2_X1 port map( A => n11301, B => n11298, S => n10762, Z => n9536
                           );
   U14809 : NAND2_X1 port map( A1 => n9841, A2 => n25207, ZN => n9521);
   U14810 : NAND2_X1 port map( A1 => n9525, A2 => n9524, ZN => n9528);
   U14811 : AOI21_X1 port map( B1 => n9526, B2 => n9775, A => n9773, ZN => 
                           n9527);
   U14812 : NAND2_X1 port map( A1 => n9532, A2 => n10113, ZN => n9535);
   U14813 : NAND3_X1 port map( A1 => n9533, A2 => n9805, A3 => n10116, ZN => 
                           n9534);
   U14814 : XNOR2_X1 port map( A => n11396, B => n9537, ZN => n11420);
   U14815 : NAND2_X1 port map( A1 => n4096, A2 => n24446, ZN => n9538);
   U14816 : MUX2_X1 port map( A => n9539, B => n9538, S => n9866, Z => n9540);
   U14817 : INV_X1 port map( A => n10028, ZN => n9543);
   U14818 : NAND2_X1 port map( A1 => n10031, A2 => n10026, ZN => n9542);
   U14819 : AOI21_X1 port map( B1 => n9543, B2 => n9542, A => n10027, ZN => 
                           n9546);
   U14820 : NAND2_X1 port map( A1 => n9697, A2 => n9695, ZN => n9643);
   U14821 : NAND3_X1 port map( A1 => n9697, A2 => n9699, A3 => n10027, ZN => 
                           n9544);
   U14822 : NAND2_X1 port map( A1 => n9643, A2 => n9544, ZN => n9545);
   U14823 : NAND3_X1 port map( A1 => n1517, A2 => n307, A3 => n9692, ZN => 
                           n9548);
   U14824 : OAI211_X2 port map( C1 => n9549, C2 => n4993, A => n9548, B => 
                           n9547, ZN => n10904);
   U14825 : NAND2_X1 port map( A1 => n10445, A2 => n10904, ZN => n9553);
   U14826 : NAND2_X1 port map( A1 => n10044, A2 => n10045, ZN => n9625);
   U14827 : OAI211_X1 port map( C1 => n10046, C2 => n9681, A => n9628, B => 
                           n9627, ZN => n9552);
   U14828 : NAND2_X1 port map( A1 => n10048, A2 => n9681, ZN => n9551);
   U14829 : NAND2_X1 port map( A1 => n9558, A2 => n9560, ZN => n9557);
   U14830 : NAND3_X1 port map( A1 => n10445, A2 => n10907, A3 => n10904, ZN => 
                           n9572);
   U14831 : NAND3_X1 port map( A1 => n9882, A2 => n9886, A3 => n9567, ZN => 
                           n9569);
   U14832 : OAI211_X1 port map( C1 => n25069, C2 => n9567, A => n9566, B => 
                           n9565, ZN => n9568);
   U14833 : NAND3_X1 port map( A1 => n10902, A2 => n10747, A3 => n10901, ZN => 
                           n9571);
   U14834 : INV_X1 port map( A => n12402, ZN => n12067);
   U14835 : NOR2_X1 port map( A1 => n10885, A2 => n10886, ZN => n9574);
   U14836 : AOI22_X1 port map( A1 => n10884, A2 => n9574, B1 => n10301, B2 => 
                           n10885, ZN => n9575);
   U14837 : OAI22_X1 port map( A1 => n10902, A2 => n10747, B1 => n4341, B2 => 
                           n10904, ZN => n9579);
   U14838 : INV_X1 port map( A => n10901, ZN => n9578);
   U14839 : NAND2_X1 port map( A1 => n10444, A2 => n10905, ZN => n9577);
   U14840 : XNOR2_X1 port map( A => n11845, B => n12150, ZN => n11087);
   U14841 : INV_X1 port map( A => n11087, ZN => n9612);
   U14843 : INV_X1 port map( A => n10284, ZN => n10286);
   U14844 : INV_X1 port map( A => n11385, ZN => n9611);
   U14845 : INV_X1 port map( A => n10617, ZN => n10610);
   U14846 : INV_X1 port map( A => n9832, ZN => n10182);
   U14847 : OAI211_X1 port map( C1 => n9832, C2 => n9831, A => n9585, B => 
                           n9584, ZN => n9587);
   U14848 : NAND3_X1 port map( A1 => n9832, A2 => n10177, A3 => n10175, ZN => 
                           n9586);
   U14849 : INV_X1 port map( A => n10612, ZN => n10341);
   U14850 : NAND2_X1 port map( A1 => n9814, A2 => n10166, ZN => n9590);
   U14851 : NAND2_X1 port map( A1 => n10341, A2 => n10411, ZN => n9610);
   U14852 : INV_X1 port map( A => n10161, ZN => n9850);
   U14853 : INV_X1 port map( A => n10157, ZN => n9851);
   U14854 : NAND3_X1 port map( A1 => n3305, A2 => n10162, A3 => n9851, ZN => 
                           n9594);
   U14855 : INV_X1 port map( A => n10486, ZN => n10410);
   U14856 : NOR2_X1 port map( A1 => n10129, A2 => n10128, ZN => n9598);
   U14857 : NAND2_X1 port map( A1 => n9595, A2 => n10127, ZN => n9596);
   U14858 : NAND3_X1 port map( A1 => n10410, A2 => n10614, A3 => n10341, ZN => 
                           n9609);
   U14859 : OAI21_X1 port map( B1 => n9927, B2 => n9934, A => n9603, ZN => 
                           n9602);
   U14860 : OAI21_X1 port map( B1 => n9600, B2 => n9599, A => n9926, ZN => 
                           n9601);
   U14861 : NAND3_X1 port map( A1 => n9928, A2 => n9604, A3 => n9603, ZN => 
                           n9606);
   U14862 : NAND2_X1 port map( A1 => n9927, A2 => n9925, ZN => n9605);
   U14864 : XNOR2_X1 port map( A => n9611, B => n12143, ZN => n11446);
   U14865 : XNOR2_X1 port map( A => n11446, B => n9612, ZN => n9680);
   U14866 : AOI21_X1 port map( B1 => n9757, B2 => n9752, A => n9753, ZN => 
                           n9618);
   U14867 : INV_X1 port map( A => n9613, ZN => n9749);
   U14868 : NOR2_X1 port map( A1 => n9754, A2 => n9749, ZN => n9614);
   U14869 : OAI21_X1 port map( B1 => n9615, B2 => n9614, A => n9977, ZN => 
                           n9616);
   U14870 : NOR2_X1 port map( A1 => n9762, A2 => n9620, ZN => n9619);
   U14871 : MUX2_X1 port map( A => n10068, B => n9619, S => n9231, Z => n9623);
   U14872 : NAND2_X1 port map( A1 => n1330, A2 => n9620, ZN => n9621);
   U14873 : OAI21_X2 port map( B1 => n9623, B2 => n9622, A => n9621, ZN => 
                           n11338);
   U14874 : NAND2_X1 port map( A1 => n10062, A2 => n9705, ZN => n9624);
   U14875 : INV_X1 port map( A => n9625, ZN => n9626);
   U14877 : OAI21_X1 port map( B1 => n9628, B2 => n9627, A => n10044, ZN => 
                           n9629);
   U14878 : NAND2_X1 port map( A1 => n9629, A2 => n9682, ZN => n9631);
   U14879 : NAND3_X1 port map( A1 => n10048, A2 => n9681, A3 => n10046, ZN => 
                           n9630);
   U14880 : MUX2_X1 port map( A => n9635, B => n9634, S => n9633, Z => n9638);
   U14881 : INV_X1 port map( A => n9714, ZN => n9636);
   U14882 : AND2_X1 port map( A1 => n9711, A2 => n10037, ZN => n10043);
   U14883 : AOI22_X1 port map( A1 => n9636, A2 => n9709, B1 => n9635, B2 => 
                           n10043, ZN => n9637);
   U14884 : OAI21_X1 port map( B1 => n9638, B2 => n9710, A => n9637, ZN => 
                           n10632);
   U14885 : INV_X1 port map( A => n9639, ZN => n10034);
   U14886 : NAND2_X1 port map( A1 => n10029, A2 => n10026, ZN => n9640);
   U14887 : NAND3_X1 port map( A1 => n9643, A2 => n10034, A3 => n9640, ZN => 
                           n9642);
   U14888 : NAND3_X1 port map( A1 => n9639, A2 => n24332, A3 => n10027, ZN => 
                           n9641);
   U14890 : NAND2_X1 port map( A1 => n10233, A2 => n10633, ZN => n9644);
   U14891 : NAND2_X1 port map( A1 => n25025, A2 => n11207, ZN => n11340);
   U14892 : OAI21_X2 port map( B1 => n9644, B2 => n9645, A => n11340, ZN => 
                           n12409);
   U14893 : NAND2_X1 port map( A1 => n413, A2 => n10831, ZN => n9649);
   U14894 : AND2_X1 port map( A1 => n10515, A2 => n9646, ZN => n9648);
   U14895 : XNOR2_X1 port map( A => n24980, B => n12409, ZN => n9678);
   U14896 : NOR2_X1 port map( A1 => n10019, A2 => n8839, ZN => n9650);
   U14897 : NOR2_X1 port map( A1 => n9721, A2 => n10005, ZN => n9651);
   U14898 : NAND2_X1 port map( A1 => n9996, A2 => n9991, ZN => n9660);
   U14900 : NOR2_X1 port map( A1 => n9746, A2 => n9990, ZN => n9661);
   U14902 : NAND3_X1 port map( A1 => n9980, A2 => n9737, A3 => n9664, ZN => 
                           n9665);
   U14903 : NAND2_X1 port map( A1 => n9737, A2 => n9981, ZN => n9666);
   U14904 : AOI21_X1 port map( B1 => n9980, B2 => n9666, A => n9740, ZN => 
                           n9667);
   U14905 : NOR2_X1 port map( A1 => n25453, A2 => n9671, ZN => n9672);
   U14906 : NAND2_X1 port map( A1 => n9672, A2 => n9796, ZN => n9673);
   U14907 : NOR2_X1 port map( A1 => n9798, A2 => n8521, ZN => n9795);
   U14908 : OAI211_X1 port map( C1 => n9781, C2 => n10093, A => n9295, B => 
                           n1348, ZN => n9675);
   U14909 : NOR2_X1 port map( A1 => n11201, A2 => n11196, ZN => n10788);
   U14910 : XNOR2_X1 port map( A => n12102, B => n859, ZN => n9677);
   U14911 : XNOR2_X1 port map( A => n9678, B => n9677, ZN => n9679);
   U14912 : AOI21_X1 port map( B1 => n12648, B2 => n12871, A => n13094, ZN => 
                           n10201);
   U14913 : OAI21_X1 port map( B1 => n9682, B2 => n10045, A => n9681, ZN => 
                           n9687);
   U14914 : NAND2_X1 port map( A1 => n9684, A2 => n10048, ZN => n9685);
   U14915 : MUX2_X1 port map( A => n9689, B => n9688, S => n4096, Z => n9690);
   U14916 : NOR2_X1 port map( A1 => n10026, A2 => n24332, ZN => n9698);
   U14917 : NOR2_X1 port map( A1 => n9639, A2 => n9699, ZN => n9700);
   U14918 : NAND2_X1 port map( A1 => n10061, A2 => n9705, ZN => n9706);
   U14919 : NAND2_X1 port map( A1 => n9708, A2 => n9707, ZN => n11143);
   U14920 : NAND2_X1 port map( A1 => n10304, A2 => n11151, ZN => n9719);
   U14922 : OR2_X1 port map( A1 => n9712, A2 => n9713, ZN => n9717);
   U14923 : INV_X1 port map( A => n10039, ZN => n9716);
   U14924 : NAND2_X1 port map( A1 => n9714, A2 => n9713, ZN => n9715);
   U14925 : OR2_X1 port map( A1 => n9718, A2 => n9433, ZN => n11146);
   U14926 : MUX2_X1 port map( A => n9723, B => n9722, S => n9299, Z => n9728);
   U14927 : NOR2_X1 port map( A1 => n9724, A2 => n10008, ZN => n9726);
   U14929 : NAND2_X1 port map( A1 => n9730, A2 => n9729, ZN => n10016);
   U14930 : INV_X1 port map( A => n10016, ZN => n9735);
   U14931 : NAND2_X1 port map( A1 => n9731, A2 => n426, ZN => n9734);
   U14932 : OAI21_X1 port map( B1 => n9735, B2 => n9734, A => n9733, ZN => 
                           n11159);
   U14933 : NAND3_X1 port map( A1 => n9740, A2 => n9737, A3 => n9985, ZN => 
                           n9738);
   U14934 : AND2_X1 port map( A1 => n9739, A2 => n9738, ZN => n9744);
   U14935 : NAND2_X1 port map( A1 => n9982, A2 => n9981, ZN => n9741);
   U14936 : MUX2_X1 port map( A => n9742, B => n9741, S => n9740, Z => n9743);
   U14937 : NAND2_X2 port map( A1 => n9743, A2 => n9744, ZN => n11157);
   U14938 : MUX2_X1 port map( A => n1358, B => n4737, S => n11157, Z => n9768);
   U14940 : NAND2_X1 port map( A1 => n9751, A2 => n9750, ZN => n9756);
   U14941 : AND3_X1 port map( A1 => n9753, A2 => n9754, A3 => n9752, ZN => 
                           n9755);
   U14942 : AOI21_X1 port map( B1 => n9756, B2 => n9973, A => n9755, ZN => 
                           n10675);
   U14943 : NAND2_X1 port map( A1 => n9758, A2 => n9757, ZN => n10673);
   U14944 : NAND2_X1 port map( A1 => n10985, A2 => n11160, ZN => n9759);
   U14945 : OAI21_X1 port map( B1 => n11160, B2 => n11157, A => n9759, ZN => 
                           n9767);
   U14946 : NOR2_X1 port map( A1 => n10075, A2 => n9231, ZN => n9761);
   U14947 : NAND3_X1 port map( A1 => n9764, A2 => n9763, A3 => n9762, ZN => 
                           n9765);
   U14948 : XNOR2_X1 port map( A => n12002, B => n11967, ZN => n11642);
   U14949 : INV_X1 port map( A => n11642, ZN => n11725);
   U14950 : OAI21_X1 port map( B1 => n10681, B2 => n24622, A => n11003, ZN => 
                           n9771);
   U14951 : MUX2_X2 port map( A => n9771, B => n9770, S => n10685, Z => n11289)
                           ;
   U14952 : MUX2_X1 port map( A => n10108, B => n9774, S => n9772, Z => n9776);
   U14953 : NAND2_X1 port map( A1 => n9774, A2 => n9773, ZN => n10110);
   U14954 : NAND2_X1 port map( A1 => n9775, A2 => n10104, ZN => n10107);
   U14955 : NAND2_X1 port map( A1 => n1348, A2 => n10089, ZN => n9778);
   U14956 : NAND2_X1 port map( A1 => n8571, A2 => n9295, ZN => n9777);
   U14957 : NAND3_X1 port map( A1 => n10090, A2 => n9778, A3 => n9777, ZN => 
                           n9785);
   U14958 : NAND3_X1 port map( A1 => n9782, A2 => n24505, A3 => n9780, ZN => 
                           n9783);
   U14959 : NOR2_X1 port map( A1 => n11054, A2 => n11009, ZN => n9803);
   U14960 : NOR2_X1 port map( A1 => n10094, A2 => n10099, ZN => n9790);
   U14961 : INV_X1 port map( A => n10094, ZN => n9791);
   U14962 : NAND2_X1 port map( A1 => n9791, A2 => n10098, ZN => n9792);
   U14963 : OAI22_X1 port map( A1 => n9838, A2 => n10095, B1 => n9792, B2 => 
                           n9837, ZN => n9793);
   U14964 : NOR3_X1 port map( A1 => n9811, A2 => n11052, A3 => n9810, ZN => 
                           n9802);
   U14965 : NOR2_X1 port map( A1 => n9997, A2 => n9998, ZN => n9799);
   U14966 : OAI21_X1 port map( B1 => n9799, B2 => n9999, A => n9798, ZN => 
                           n9800);
   U14967 : INV_X1 port map( A => n11440, ZN => n9812);
   U14968 : XNOR2_X1 port map( A => n11289, B => n9812, ZN => n9813);
   U14969 : XNOR2_X1 port map( A => n11725, B => n9813, ZN => n9971);
   U14970 : INV_X1 port map( A => n9820, ZN => n9821);
   U14971 : NAND2_X1 port map( A1 => n25463, A2 => n9821, ZN => n9824);
   U14972 : NAND3_X1 port map( A1 => n10136, A2 => n9820, A3 => n25463, ZN => 
                           n9823);
   U14974 : OAI211_X1 port map( C1 => n10138, C2 => n9824, A => n9823, B => 
                           n9822, ZN => n9826);
   U14975 : INV_X1 port map( A => n9827, ZN => n9828);
   U14976 : NAND2_X1 port map( A1 => n9828, A2 => n10176, ZN => n9835);
   U14977 : OAI211_X1 port map( C1 => n9831, C2 => n10175, A => n9830, B => 
                           n9829, ZN => n9834);
   U14978 : NAND3_X1 port map( A1 => n10186, A2 => n9832, A3 => n10178, ZN => 
                           n9833);
   U14979 : INV_X1 port map( A => n10703, ZN => n10699);
   U14980 : OAI21_X1 port map( B1 => n25206, B2 => n25486, A => n9841, ZN => 
                           n9848);
   U14981 : NAND2_X1 port map( A1 => n9844, A2 => n10148, ZN => n9847);
   U14982 : NAND3_X1 port map( A1 => n1210, A2 => n24085, A3 => n9845, ZN => 
                           n9846);
   U14983 : OAI211_X1 port map( C1 => n9851, C2 => n10162, A => n9850, B => 
                           n9849, ZN => n9852);
   U14984 : OAI21_X1 port map( B1 => n9854, B2 => n9853, A => n9852, ZN => 
                           n10953);
   U14985 : INV_X1 port map( A => n11637, ZN => n9855);
   U14986 : XNOR2_X1 port map( A => n9855, B => n2761, ZN => n9969);
   U14987 : MUX2_X1 port map( A => n239, B => n9860, S => n9856, Z => n9865);
   U14988 : NAND2_X1 port map( A1 => n9857, A2 => n9864, ZN => n9862);
   U14989 : MUX2_X1 port map( A => n9862, B => n9861, S => n9860, Z => n9863);
   U14991 : INV_X1 port map( A => n10971, ZN => n9871);
   U14992 : INV_X1 port map( A => n9867, ZN => n9868);
   U14993 : NAND2_X1 port map( A1 => n9871, A2 => n10970, ZN => n10608);
   U14994 : NAND3_X1 port map( A1 => n9875, A2 => n24549, A3 => n9027, ZN => 
                           n9878);
   U14995 : INV_X1 port map( A => n9876, ZN => n9877);
   U14996 : NAND2_X1 port map( A1 => n25497, A2 => n10968, ZN => n9881);
   U14997 : NAND2_X1 port map( A1 => n10608, A2 => n9881, ZN => n9911);
   U14998 : NAND2_X1 port map( A1 => n8157, A2 => n9886, ZN => n9888);
   U14999 : NAND2_X1 port map( A1 => n9891, A2 => n9890, ZN => n9892);
   U15000 : INV_X1 port map( A => n9892, ZN => n10967);
   U15001 : NAND2_X1 port map( A1 => n227, A2 => n9943, ZN => n9894);
   U15002 : NAND2_X1 port map( A1 => n9895, A2 => n9894, ZN => n9896);
   U15003 : NAND3_X1 port map( A1 => n9899, A2 => n24054, A3 => n9897, ZN => 
                           n9901);
   U15004 : NAND3_X1 port map( A1 => n9942, A2 => n9946, A3 => n24083, ZN => 
                           n9900);
   U15005 : NOR2_X1 port map( A1 => n10818, A2 => n9903, ZN => n9910);
   U15006 : OAI21_X1 port map( B1 => n9908, B2 => n9907, A => n9906, ZN => 
                           n9909);
   U15007 : INV_X1 port map( A => n9912, ZN => n9917);
   U15008 : INV_X1 port map( A => n9913, ZN => n9915);
   U15009 : AOI22_X1 port map( A1 => n9917, A2 => n9916, B1 => n9915, B2 => 
                           n9914, ZN => n9924);
   U15010 : NAND2_X1 port map( A1 => n24844, A2 => n9918, ZN => n9922);
   U15012 : INV_X1 port map( A => n9929, ZN => n9933);
   U15013 : INV_X1 port map( A => n9930, ZN => n9932);
   U15015 : OAI21_X1 port map( B1 => n9939, B2 => n9938, A => n9937, ZN => 
                           n9940);
   U15016 : NAND2_X1 port map( A1 => n10804, A2 => n411, ZN => n9968);
   U15017 : NAND3_X1 port map( A1 => n10798, A2 => n10799, A3 => n10648, ZN => 
                           n9967);
   U15018 : MUX2_X1 port map( A => n9953, B => n9948, S => n9947, Z => n9960);
   U15019 : NAND2_X1 port map( A1 => n9950, A2 => n9949, ZN => n9956);
   U15020 : OAI21_X1 port map( B1 => n9956, B2 => n9955, A => n9954, ZN => 
                           n9957);
   U15021 : INV_X1 port map( A => n9957, ZN => n9958);
   U15022 : OAI21_X1 port map( B1 => n9960, B2 => n9959, A => n9958, ZN => 
                           n10426);
   U15023 : INV_X1 port map( A => n10426, ZN => n10649);
   U15024 : NOR2_X1 port map( A1 => n10649, A2 => n10648, ZN => n10803);
   U15025 : INV_X1 port map( A => n10651, ZN => n10801);
   U15026 : INV_X1 port map( A => n10245, ZN => n10244);
   U15027 : XNOR2_X1 port map( A => n11194, B => n9969, ZN => n9970);
   U15028 : OAI21_X1 port map( B1 => n9975, B2 => n9974, A => n9973, ZN => 
                           n9976);
   U15029 : NAND2_X1 port map( A1 => n9978, A2 => n9981, ZN => n9979);
   U15031 : MUX2_X1 port map( A => n9991, B => n9990, S => n9989, Z => n9994);
   U15032 : INV_X1 port map( A => n11045, ZN => n10642);
   U15033 : AOI21_X1 port map( B1 => n2680, B2 => n11046, A => n10642, ZN => 
                           n10014);
   U15034 : NAND2_X1 port map( A1 => n10006, A2 => n10005, ZN => n10011);
   U15035 : NOR2_X1 port map( A1 => n25043, A2 => n9301, ZN => n10010);
   U15036 : NAND2_X1 port map( A1 => n9299, A2 => n10008, ZN => n10009);
   U15037 : AOI22_X1 port map( A1 => n10012, A2 => n10011, B1 => n10010, B2 => 
                           n10009, ZN => n11051);
   U15038 : MUX2_X1 port map( A => n10020, B => n10019, S => n10018, Z => 
                           n10021);
   U15039 : NOR2_X1 port map( A1 => n10021, A2 => n8839, ZN => n10022);
   U15040 : NAND2_X1 port map( A1 => n11044, A2 => n10416, ZN => n11050);
   U15041 : NAND2_X1 port map( A1 => n10801, A2 => n10648, ZN => n10025);
   U15042 : OAI21_X1 port map( B1 => n10426, B2 => n10245, A => n10799, ZN => 
                           n10023);
   U15043 : NOR2_X1 port map( A1 => n10023, A2 => n411, ZN => n10024);
   U15044 : AOI21_X2 port map( B1 => n10427, B2 => n10025, A => n10024, ZN => 
                           n11542);
   U15045 : XNOR2_X1 port map( A => n11542, B => n12082, ZN => n10124);
   U15046 : MUX2_X1 port map( A => n10031, B => n24332, S => n10026, Z => 
                           n10035);
   U15047 : NAND2_X1 port map( A1 => n10028, A2 => n10027, ZN => n10033);
   U15048 : NAND3_X1 port map( A1 => n10031, A2 => n24332, A3 => n10029, ZN => 
                           n10032);
   U15049 : OAI211_X2 port map( C1 => n10035, C2 => n10034, A => n10033, B => 
                           n10032, ZN => n11064);
   U15050 : NAND2_X1 port map( A1 => n9433, A2 => n9709, ZN => n10042);
   U15051 : NAND2_X1 port map( A1 => n10038, A2 => n10037, ZN => n10040);
   U15052 : NAND2_X1 port map( A1 => n10040, A2 => n10039, ZN => n10041);
   U15053 : NOR2_X1 port map( A1 => n11064, A2 => n11069, ZN => n10665);
   U15054 : MUX2_X1 port map( A => n10045, B => n260, S => n10044, Z => n10049)
                           ;
   U15055 : OAI21_X1 port map( B1 => n10052, B2 => n10051, A => n10050, ZN => 
                           n10056);
   U15056 : MUX2_X1 port map( A => n10064, B => n10063, S => n9127, Z => n10066
                           );
   U15057 : OAI22_X1 port map( A1 => n1330, A2 => n10070, B1 => n25457, B2 => 
                           n9231, ZN => n10073);
   U15058 : NAND2_X1 port map( A1 => n10073, A2 => n10072, ZN => n10074);
   U15060 : INV_X1 port map( A => n11062, ZN => n11071);
   U15061 : NOR2_X1 port map( A1 => n11070, A2 => n11071, ZN => n10078);
   U15062 : INV_X1 port map( A => n10665, ZN => n10077);
   U15063 : NAND2_X1 port map( A1 => n10080, A2 => n10079, ZN => n10081);
   U15064 : NAND2_X1 port map( A1 => n10087, A2 => n10081, ZN => n10085);
   U15065 : NAND2_X1 port map( A1 => n10082, A2 => n10088, ZN => n10084);
   U15066 : MUX2_X1 port map( A => n10085, B => n10084, S => n24575, Z => 
                           n10086);
   U15067 : NAND2_X1 port map( A1 => n10091, A2 => n10090, ZN => n10092);
   U15068 : NAND3_X1 port map( A1 => n10100, A2 => n10094, A3 => n10099, ZN => 
                           n10096);
   U15069 : OAI21_X1 port map( B1 => n421, B2 => n10097, A => n10096, ZN => 
                           n10103);
   U15072 : NOR2_X1 port map( A1 => n10110, A2 => n10109, ZN => n10111);
   U15073 : OAI22_X1 port map( A1 => n10114, A2 => n1406, B1 => n10113, B2 => 
                           n10112, ZN => n10119);
   U15074 : NAND3_X1 port map( A1 => n10117, A2 => n10116, A3 => n10115, ZN => 
                           n10118);
   U15075 : XNOR2_X1 port map( A => n12053, B => n11424, ZN => n11391);
   U15076 : XNOR2_X1 port map( A => n11391, B => n10124, ZN => n10198);
   U15077 : NAND2_X1 port map( A1 => n10127, A2 => n10126, ZN => n10133);
   U15078 : NAND2_X1 port map( A1 => n10129, A2 => n10128, ZN => n10130);
   U15080 : INV_X1 port map( A => n10559, ZN => n10659);
   U15082 : NOR2_X1 port map( A1 => n9398, A2 => n24026, ZN => n10139);
   U15083 : OAI21_X1 port map( B1 => n10139, B2 => n10138, A => n25463, ZN => 
                           n10144);
   U15084 : NAND2_X1 port map( A1 => n10659, A2 => n10654, ZN => n10314);
   U15085 : NOR2_X1 port map( A1 => n25206, A2 => n10148, ZN => n10152);
   U15086 : NOR2_X1 port map( A1 => n10149, A2 => n10148, ZN => n10151);
   U15087 : NOR2_X1 port map( A1 => n10158, A2 => n10157, ZN => n10160);
   U15088 : OAI22_X1 port map( A1 => n3305, A2 => n10162, B1 => n10161, B2 => 
                           n9349, ZN => n10164);
   U15089 : OAI21_X1 port map( B1 => n10165, B2 => n25250, A => n10657, ZN => 
                           n10189);
   U15090 : NOR2_X1 port map( A1 => n10170, A2 => n10169, ZN => n10171);
   U15091 : NOR2_X1 port map( A1 => n10172, A2 => n1577, ZN => n10173);
   U15092 : NAND3_X1 port map( A1 => n10176, A2 => n10178, A3 => n10175, ZN => 
                           n10184);
   U15093 : INV_X1 port map( A => n10177, ZN => n10179);
   U15094 : NOR2_X1 port map( A1 => n10654, A2 => n10660, ZN => n10187);
   U15095 : OAI21_X1 port map( B1 => n10661, B2 => n25250, A => n10187, ZN => 
                           n10188);
   U15096 : NAND2_X1 port map( A1 => n10189, A2 => n10188, ZN => n11660);
   U15097 : INV_X1 port map( A => n25229, ZN => n10854);
   U15099 : INV_X1 port map( A => n10737, ZN => n10465);
   U15100 : OAI211_X1 port map( C1 => n10831, C2 => n10277, A => n10830, B => 
                           n10518, ZN => n10194);
   U15101 : XNOR2_X1 port map( A => n12255, B => n22702, ZN => n10195);
   U15102 : XNOR2_X1 port map( A => n10196, B => n10195, ZN => n10197);
   U15103 : INV_X1 port map( A => n14158, ZN => n10396);
   U15104 : NOR2_X1 port map( A1 => n10756, A2 => n10757, ZN => n10203);
   U15105 : NOR2_X1 port map( A1 => n11298, A2 => n11301, ZN => n10205);
   U15106 : NAND2_X1 port map( A1 => n10895, A2 => n10205, ZN => n10207);
   U15107 : NAND3_X1 port map( A1 => n11091, A2 => n11301, A3 => n10762, ZN => 
                           n10206);
   U15108 : XNOR2_X1 port map( A => n12314, B => n11263, ZN => n11829);
   U15109 : INV_X1 port map( A => n10208, ZN => n10211);
   U15110 : INV_X1 port map( A => n10209, ZN => n10210);
   U15111 : NAND3_X1 port map( A1 => n10211, A2 => n10538, A3 => n10210, ZN => 
                           n10212);
   U15112 : NAND2_X1 port map( A1 => n10585, A2 => n10371, ZN => n10317);
   U15113 : INV_X1 port map( A => n10584, ZN => n10582);
   U15114 : AND2_X1 port map( A1 => n10587, A2 => n25507, ZN => n10215);
   U15115 : OAI21_X1 port map( B1 => n10590, B2 => n10584, A => n10215, ZN => 
                           n10216);
   U15116 : NAND2_X1 port map( A1 => n10217, A2 => n10216, ZN => n11747);
   U15117 : XNOR2_X1 port map( A => n12218, B => n11747, ZN => n11481);
   U15118 : XNOR2_X1 port map( A => n11829, B => n11481, ZN => n10226);
   U15119 : INV_X1 port map( A => n10891, ZN => n11081);
   U15120 : NAND2_X1 port map( A1 => n10767, A2 => n412, ZN => n10766);
   U15122 : XNOR2_X1 port map( A => n11616, B => n12313, ZN => n10224);
   U15123 : INV_X1 port map( A => n10904, ZN => n10899);
   U15124 : XNOR2_X1 port map( A => n12159, B => n2228, ZN => n10223);
   U15125 : XNOR2_X1 port map( A => n10224, B => n10223, ZN => n10225);
   U15126 : XNOR2_X1 port map( A => n10226, B => n10225, ZN => n12724);
   U15127 : INV_X1 port map( A => n12724, ZN => n13176);
   U15129 : NAND2_X1 port map( A1 => n44, A2 => n11199, ZN => n10228);
   U15130 : NAND2_X1 port map( A1 => n11201, A2 => n11196, ZN => n10227);
   U15132 : INV_X1 port map( A => n10789, ZN => n11195);
   U15133 : OAI211_X1 port map( C1 => n10793, C2 => n11195, A => n10477, B => 
                           n10229, ZN => n10230);
   U15134 : AND2_X1 port map( A1 => n10632, A2 => n11338, ZN => n10232);
   U15135 : INV_X1 port map( A => n10411, ZN => n10489);
   U15136 : AOI22_X1 port map( A1 => n10617, A2 => n10616, B1 => n10489, B2 => 
                           n10614, ZN => n10237);
   U15137 : NOR2_X1 port map( A1 => n10614, A2 => n10486, ZN => n10234);
   U15138 : NAND2_X1 port map( A1 => n10610, A2 => n10234, ZN => n10236);
   U15139 : NOR3_X1 port map( A1 => n10486, A2 => n10411, A3 => n10613, ZN => 
                           n10235);
   U15140 : NAND3_X1 port map( A1 => n233, A2 => n11212, A3 => n11216, ZN => 
                           n10238);
   U15141 : XNOR2_X1 port map( A => n10239, B => n12046, ZN => n10270);
   U15142 : INV_X1 port map( A => n10968, ZN => n10607);
   U15143 : OAI21_X1 port map( B1 => n10497, B2 => n10607, A => n10606, ZN => 
                           n10240);
   U15144 : NOR2_X1 port map( A1 => n25497, A2 => n10968, ZN => n10496);
   U15145 : NOR2_X1 port map( A1 => n10606, A2 => n10969, ZN => n10242);
   U15146 : NOR2_X1 port map( A1 => n25497, A2 => n10970, ZN => n10241);
   U15147 : NAND3_X1 port map( A1 => n10805, A2 => n10799, A3 => n10244, ZN => 
                           n10247);
   U15148 : NAND4_X2 port map( A1 => n10246, A2 => n10248, A3 => n10249, A4 => 
                           n10247, ZN => n12201);
   U15149 : XNOR2_X1 port map( A => n12122, B => n12201, ZN => n12242);
   U15150 : INV_X1 port map( A => n10256, ZN => n10258);
   U15151 : AND2_X1 port map( A1 => n10257, A2 => n10258, ZN => n10260);
   U15152 : NAND4_X1 port map( A1 => n10261, A2 => n10480, A3 => n10260, A4 => 
                           n10259, ZN => n10265);
   U15153 : INV_X1 port map( A => n10262, ZN => n10263);
   U15154 : NAND2_X1 port map( A1 => n10263, A2 => n11190, ZN => n10264);
   U15156 : XNOR2_X1 port map( A => n12383, B => n3125, ZN => n10268);
   U15157 : XNOR2_X1 port map( A => n12242, B => n10268, ZN => n10269);
   U15158 : INV_X1 port map( A => n12459, ZN => n13177);
   U15159 : NAND2_X1 port map( A1 => n11189, A2 => n11190, ZN => n11371);
   U15160 : NOR2_X1 port map( A1 => n11190, A2 => n10728, ZN => n11185);
   U15161 : NAND2_X1 port map( A1 => n11371, A2 => n11370, ZN => n11809);
   U15163 : MUX2_X1 port map( A => n10464, B => n10272, S => n11123, Z => 
                           n10274);
   U15164 : INV_X1 port map( A => n11123, ZN => n10720);
   U15165 : AND2_X1 port map( A1 => n10850, A2 => n2244, ZN => n10851);
   U15166 : AOI22_X1 port map( A1 => n10851, A2 => n11124, B1 => n10722, B2 => 
                           n10848, ZN => n10273);
   U15167 : XNOR2_X1 port map( A => n11809, B => n11492, ZN => n12303);
   U15168 : NAND2_X1 port map( A1 => n10829, A2 => n10277, ZN => n10514);
   U15169 : NOR2_X1 port map( A1 => n9279, A2 => n10514, ZN => n10278);
   U15170 : NOR2_X2 port map( A1 => n10279, A2 => n10278, ZN => n12184);
   U15171 : OAI21_X1 port map( B1 => n10860, B2 => n10861, A => n10854, ZN => 
                           n10281);
   U15172 : XNOR2_X1 port map( A => n12184, B => n12128, ZN => n12269);
   U15174 : MUX2_X1 port map( A => n10284, B => n24574, S => n11117, Z => 
                           n10289);
   U15175 : INV_X1 port map( A => n10285, ZN => n10287);
   U15176 : NAND2_X1 port map( A1 => n10287, A2 => n10727, ZN => n10288);
   U15177 : INV_X1 port map( A => n10451, ZN => n10752);
   U15178 : XNOR2_X1 port map( A => n11966, B => n12186, ZN => n10298);
   U15179 : NAND2_X1 port map( A1 => n10713, A2 => n11128, ZN => n10296);
   U15180 : AND2_X1 port map( A1 => n11128, A2 => n11130, ZN => n10712);
   U15181 : INV_X1 port map( A => n10712, ZN => n10292);
   U15183 : XNOR2_X1 port map( A => n11698, B => n20825, ZN => n10297);
   U15184 : XNOR2_X1 port map( A => n10298, B => n10297, ZN => n10299);
   U15185 : AOI21_X1 port map( B1 => n10541, B2 => n10885, A => n10887, ZN => 
                           n10303);
   U15186 : INV_X1 port map( A => n10304, ZN => n10305);
   U15187 : NAND3_X1 port map( A1 => n714, A2 => n11143, A3 => n1357, ZN => 
                           n10307);
   U15188 : XNOR2_X1 port map( A => n11310, B => n11776, ZN => n11536);
   U15189 : INV_X1 port map( A => n11157, ZN => n10676);
   U15190 : OAI21_X1 port map( B1 => n10676, B2 => n4737, A => n11158, ZN => 
                           n10309);
   U15191 : XNOR2_X1 port map( A => n11607, B => n21204, ZN => n10310);
   U15192 : NAND2_X1 port map( A1 => n10548, A2 => n2754, ZN => n10311);
   U15193 : OAI211_X1 port map( C1 => n10548, C2 => n10950, A => n10312, B => 
                           n10311, ZN => n12297);
   U15194 : NAND2_X1 port map( A1 => n11170, A2 => n11168, ZN => n10940);
   U15196 : OAI21_X1 port map( B1 => n10587, B2 => n25507, A => n10585, ZN => 
                           n10318);
   U15197 : XNOR2_X1 port map( A => n12248, B => n25371, ZN => n11489);
   U15198 : XNOR2_X1 port map( A => n11489, B => n12028, ZN => n10320);
   U15199 : NOR2_X1 port map( A1 => n10360, A2 => n12724, ZN => n10361);
   U15200 : INV_X1 port map( A => n11005, ZN => n10365);
   U15201 : MUX2_X1 port map( A => n5746, B => n10321, S => n10685, Z => n10324
                           );
   U15202 : NAND2_X1 port map( A1 => n10684, A2 => n24622, ZN => n10322);
   U15203 : AOI21_X1 port map( B1 => n11003, B2 => n10322, A => n10369, ZN => 
                           n10323);
   U15205 : INV_X1 port map( A => n10924, ZN => n10989);
   U15207 : NAND3_X1 port map( A1 => n24118, A2 => n10405, A3 => n10990, ZN => 
                           n10325);
   U15208 : NAND2_X1 port map( A1 => n10924, A2 => n10993, ZN => n10407);
   U15209 : OAI21_X1 port map( B1 => n10407, B2 => n24118, A => n10328, ZN => 
                           n10329);
   U15210 : XNOR2_X1 port map( A => n12109, B => n12189, ZN => n12274);
   U15211 : AOI21_X1 port map( B1 => n11052, B2 => n11057, A => n11054, ZN => 
                           n11500);
   U15212 : NAND2_X1 port map( A1 => n11500, A2 => n11059, ZN => n10335);
   U15213 : NAND2_X1 port map( A1 => n11500, A2 => n11052, ZN => n10334);
   U15214 : INV_X1 port map( A => n11052, ZN => n10694);
   U15216 : OR2_X1 port map( A1 => n11059, A2 => n10331, ZN => n10333);
   U15217 : NOR2_X1 port map( A1 => n11499, A2 => n11009, ZN => n10332);
   U15218 : NAND2_X1 port map( A1 => n11054, A2 => n10332, ZN => n11501);
   U15219 : NAND4_X1 port map( A1 => n10335, A2 => n10334, A3 => n10333, A4 => 
                           n11501, ZN => n11274);
   U15220 : OAI22_X1 port map( A1 => n10337, A2 => n10398, B1 => n10658, B2 => 
                           n10559, ZN => n10340);
   U15221 : OR2_X1 port map( A1 => n10559, A2 => n10660, ZN => n10400);
   U15222 : INV_X1 port map( A => n10654, ZN => n10557);
   U15223 : NAND2_X1 port map( A1 => n10559, A2 => n10557, ZN => n10338);
   U15224 : AOI21_X1 port map( B1 => n10400, B2 => n10338, A => n10558, ZN => 
                           n10339);
   U15226 : XNOR2_X1 port map( A => n11622, B => n11274, ZN => n12063);
   U15227 : XNOR2_X1 port map( A => n12274, B => n12063, ZN => n10359);
   U15228 : AND2_X1 port map( A1 => n10486, A2 => n10613, ZN => n10342);
   U15229 : NOR2_X1 port map( A1 => n10488, A2 => n10613, ZN => n10343);
   U15230 : NOR3_X1 port map( A1 => n10343, A2 => n10342, A3 => n10610, ZN => 
                           n10344);
   U15231 : MUX2_X1 port map( A => n11068, B => n11062, S => n11064, Z => 
                           n10346);
   U15232 : NAND2_X1 port map( A1 => n10346, A2 => n25203, ZN => n10350);
   U15233 : NAND3_X1 port map( A1 => n11070, A2 => n11071, A3 => n11067, ZN => 
                           n10349);
   U15234 : INV_X1 port map( A => n25203, ZN => n10662);
   U15235 : AND3_X2 port map( A1 => n10350, A2 => n10349, A3 => n10348, ZN => 
                           n12333);
   U15236 : XNOR2_X1 port map( A => n11951, B => n12333, ZN => n10357);
   U15237 : NOR2_X1 port map( A1 => n11045, A2 => n2680, ZN => n10352);
   U15238 : NOR2_X1 port map( A1 => n10642, A2 => n11044, ZN => n10351);
   U15239 : OAI21_X1 port map( B1 => n10352, B2 => n10351, A => n11012, ZN => 
                           n10355);
   U15240 : NAND3_X1 port map( A1 => n11044, A2 => n2680, A3 => n10641, ZN => 
                           n10354);
   U15241 : NAND3_X1 port map( A1 => n10355, A2 => n10354, A3 => n10353, ZN => 
                           n11686);
   U15242 : XNOR2_X1 port map( A => n11686, B => n1863, ZN => n10356);
   U15243 : XNOR2_X1 port map( A => n10357, B => n10356, ZN => n10358);
   U15244 : XNOR2_X1 port map( A => n10359, B => n10358, ZN => n12725);
   U15245 : INV_X1 port map( A => n12460, ZN => n12651);
   U15246 : OAI22_X1 port map( A1 => n10362, A2 => n10361, B1 => n12651, B2 => 
                           n12506, ZN => n10395);
   U15247 : NAND3_X1 port map( A1 => n10365, A2 => n10681, A3 => n11004, ZN => 
                           n10366);
   U15249 : XNOR2_X1 port map( A => n11960, B => n4233, ZN => n10378);
   U15250 : INV_X1 port map( A => n10370, ZN => n10374);
   U15251 : AND2_X1 port map( A1 => n10587, A2 => n10371, ZN => n10373);
   U15252 : OAI21_X1 port map( B1 => n10374, B2 => n10373, A => n10372, ZN => 
                           n10377);
   U15253 : AOI22_X1 port map( A1 => n10589, A2 => n10590, B1 => n10375, B2 => 
                           n10585, ZN => n10376);
   U15254 : XNOR2_X1 port map( A => n10378, B => n12324, ZN => n10381);
   U15255 : INV_X1 port map( A => n10942, ZN => n10574);
   U15256 : OAI21_X1 port map( B1 => n10406, B2 => n10990, A => n10927, ZN => 
                           n10380);
   U15257 : XNOR2_X1 port map( A => n12151, B => n12207, ZN => n12288);
   U15258 : XNOR2_X1 port map( A => n12288, B => n10381, ZN => n10392);
   U15259 : NAND3_X1 port map( A1 => n11175, A2 => n11171, A3 => n24957, ZN => 
                           n10383);
   U15260 : AOI21_X1 port map( B1 => n11529, B2 => n11520, A => n10922, ZN => 
                           n10386);
   U15261 : OAI21_X1 port map( B1 => n10384, B2 => n11525, A => n11522, ZN => 
                           n10385);
   U15262 : OAI22_X1 port map( A1 => n10386, A2 => n10385, B1 => n11520, B2 => 
                           n11525, ZN => n10387);
   U15263 : XNOR2_X1 port map( A => n11959, B => n10387, ZN => n10391);
   U15264 : NOR2_X1 port map( A1 => n10935, A2 => n10931, ZN => n10389);
   U15265 : NOR2_X1 port map( A1 => n10931, A2 => n10505, ZN => n10388);
   U15266 : AOI22_X1 port map( A1 => n10936, A2 => n10389, B1 => n10388, B2 => 
                           n24470, ZN => n10390);
   U15267 : INV_X1 port map( A => n10594, ZN => n10595);
   U15268 : XNOR2_X1 port map( A => n10391, B => n12213, ZN => n11284);
   U15270 : OAI21_X1 port map( B1 => n10398, B2 => n10558, A => n10397, ZN => 
                           n10402);
   U15271 : NAND2_X1 port map( A1 => n10400, A2 => n10399, ZN => n10401);
   U15272 : MUX2_X1 port map( A => n11067, B => n11064, S => n11070, Z => 
                           n10404);
   U15273 : MUX2_X1 port map( A => n25203, B => n11069, S => n11064, Z => 
                           n10403);
   U15274 : MUX2_X1 port map( A => n10404, B => n10403, S => n11062, Z => 
                           n12130);
   U15275 : MUX2_X1 port map( A => n10994, B => n10406, S => n10405, Z => 
                           n10409);
   U15276 : OAI21_X1 port map( B1 => n10993, B2 => n10409, A => n10408, ZN => 
                           n12351);
   U15277 : XNOR2_X1 port map( A => n12130, B => n12351, ZN => n12005);
   U15278 : NAND2_X1 port map( A1 => n10410, A2 => n10489, ZN => n10414);
   U15279 : NOR2_X1 port map( A1 => n10411, A2 => n10612, ZN => n10487);
   U15280 : NAND2_X1 port map( A1 => n10617, A2 => n10487, ZN => n10413);
   U15281 : XNOR2_X1 port map( A => n11237, B => n11289, ZN => n11494);
   U15282 : NOR2_X1 port map( A1 => n11011, A2 => n10415, ZN => n10417);
   U15283 : XNOR2_X1 port map( A => n11771, B => n673, ZN => n10419);
   U15284 : XNOR2_X1 port map( A => n11494, B => n10419, ZN => n10420);
   U15285 : NOR2_X1 port map( A1 => n10594, A2 => n10505, ZN => n10422);
   U15286 : OAI21_X1 port map( B1 => n10422, B2 => n2311, A => n10936, ZN => 
                           n10424);
   U15287 : NAND3_X1 port map( A1 => n10934, A2 => n5198, A3 => n10931, ZN => 
                           n10423);
   U15288 : OAI211_X1 port map( C1 => n10936, C2 => n10425, A => n10424, B => 
                           n10423, ZN => n12233);
   U15291 : NAND2_X2 port map( A1 => n10429, A2 => n10430, ZN => n12362);
   U15292 : XNOR2_X1 port map( A => n12233, B => n12362, ZN => n10432);
   U15293 : XNOR2_X1 port map( A => n10432, B => n10431, ZN => n10450);
   U15294 : NAND2_X1 port map( A1 => n11301, A2 => n10762, ZN => n10433);
   U15295 : NAND2_X1 port map( A1 => n10434, A2 => n10433, ZN => n10437);
   U15297 : NAND2_X1 port map( A1 => n10435, A2 => n10762, ZN => n10436);
   U15298 : XNOR2_X1 port map( A => n11414, B => n11646, ZN => n12087);
   U15299 : NAND2_X1 port map( A1 => n10439, A2 => n10767, ZN => n10440);
   U15302 : NAND2_X1 port map( A1 => n10443, A2 => n10751, ZN => n10448);
   U15303 : NAND3_X1 port map( A1 => n10445, A2 => n10746, A3 => n10901, ZN => 
                           n10446);
   U15304 : XNOR2_X1 port map( A => n11908, B => n11412, ZN => n11355);
   U15305 : XNOR2_X1 port map( A => n12087, B => n11355, ZN => n10449);
   U15307 : NAND2_X1 port map( A1 => n10752, A2 => n10757, ZN => n10453);
   U15309 : XNOR2_X1 port map( A => n12209, B => n11782, ZN => n11515);
   U15310 : NAND2_X1 port map( A1 => n10729, A2 => n10457, ZN => n10456);
   U15311 : NAND2_X1 port map( A1 => n10456, A2 => n10481, ZN => n10459);
   U15312 : NOR2_X1 port map( A1 => n10457, A2 => n11190, ZN => n10458);
   U15313 : XNOR2_X1 port map( A => n11515, B => n11848, ZN => n10476);
   U15314 : OAI21_X1 port map( B1 => n10850, B2 => n11122, A => n10460, ZN => 
                           n10463);
   U15316 : NAND2_X1 port map( A1 => n10740, A2 => n10860, ZN => n10469);
   U15317 : NAND2_X1 port map( A1 => n10862, A2 => n10860, ZN => n10468);
   U15318 : NAND3_X1 port map( A1 => n10465, A2 => n10861, A3 => n25230, ZN => 
                           n10467);
   U15319 : XNOR2_X1 port map( A => n12147, B => n11741, ZN => n11992);
   U15320 : AOI21_X1 port map( B1 => n11129, B2 => n11128, A => n11130, ZN => 
                           n10473);
   U15321 : AND2_X1 port map( A1 => n11128, A2 => n10714, ZN => n10841);
   U15322 : NAND2_X1 port map( A1 => n10841, A2 => n10470, ZN => n10471);
   U15323 : XNOR2_X1 port map( A => n12286, B => n663, ZN => n10474);
   U15324 : XNOR2_X1 port map( A => n11992, B => n10474, ZN => n10475);
   U15325 : XNOR2_X1 port map( A => n10475, B => n10476, ZN => n13170);
   U15326 : INV_X1 port map( A => n13170, ZN => n10502);
   U15329 : XNOR2_X1 port map( A => n11542, B => n12257, ZN => n10485);
   U15330 : NAND2_X1 port map( A1 => n10729, A2 => n10481, ZN => n10483);
   U15331 : XNOR2_X1 port map( A => n12224, B => n4164, ZN => n10484);
   U15332 : XNOR2_X1 port map( A => n10485, B => n10484, ZN => n10501);
   U15333 : XNOR2_X1 port map( A => n10490, B => n11659, ZN => n11861);
   U15334 : OAI21_X1 port map( B1 => n11340, B2 => n11338, A => n10493, ZN => 
                           n10494);
   U15335 : NAND2_X1 port map( A1 => n11935, A2 => n10494, ZN => n10499);
   U15336 : NAND2_X1 port map( A1 => n10970, A2 => n10968, ZN => n10604);
   U15337 : NAND2_X1 port map( A1 => n10496, A2 => n10495, ZN => n10498);
   U15338 : NAND2_X1 port map( A1 => n10497, A2 => n10606, ZN => n10605);
   U15339 : OAI211_X1 port map( C1 => n10497, C2 => n10604, A => n10498, B => 
                           n10605, ZN => n11746);
   U15340 : XNOR2_X1 port map( A => n10499, B => n11746, ZN => n11429);
   U15341 : XNOR2_X1 port map( A => n11861, B => n11429, ZN => n10500);
   U15342 : XNOR2_X2 port map( A => n10501, B => n10500, ZN => n13167);
   U15343 : NAND2_X1 port map( A1 => n10951, A2 => n10952, ZN => n10504);
   U15344 : NAND3_X1 port map( A1 => n5107, A2 => n10698, A3 => n10702, ZN => 
                           n10503);
   U15345 : NAND2_X1 port map( A1 => n10934, A2 => n24470, ZN => n10507);
   U15346 : NAND2_X1 port map( A1 => n2311, A2 => n10505, ZN => n10506);
   U15347 : AOI21_X1 port map( B1 => n10507, B2 => n10506, A => n10596, ZN => 
                           n10511);
   U15349 : XNOR2_X1 port map( A => n11672, B => n11396, ZN => n12110);
   U15350 : XNOR2_X1 port map( A => n11504, B => n12110, ZN => n10530);
   U15351 : NOR2_X1 port map( A1 => n11036, A2 => n10941, ZN => n10512);
   U15352 : OAI22_X1 port map( A1 => n10515, A2 => n10829, B1 => n10836, B2 => 
                           n10514, ZN => n10522);
   U15353 : NAND3_X1 port map( A1 => n10518, A2 => n10517, A3 => n10516, ZN => 
                           n10519);
   U15354 : AOI21_X1 port map( B1 => n10520, B2 => n10519, A => n9279, ZN => 
                           n10521);
   U15355 : NOR2_X1 port map( A1 => n10522, A2 => n10521, ZN => n11756);
   U15356 : XNOR2_X1 port map( A => n12276, B => n11756, ZN => n11975);
   U15357 : MUX2_X1 port map( A => n11518, B => n11519, S => n10523, Z => 
                           n10527);
   U15358 : NOR2_X1 port map( A1 => n11520, A2 => n11524, ZN => n10524);
   U15359 : XNOR2_X1 port map( A => n12277, B => n2757, ZN => n10528);
   U15360 : XNOR2_X1 port map( A => n11975, B => n10528, ZN => n10529);
   U15361 : INV_X1 port map( A => n13165, ZN => n11597);
   U15362 : OAI21_X1 port map( B1 => n10532, B2 => n10531, A => n11597, ZN => 
                           n10569);
   U15363 : NAND2_X1 port map( A1 => n11151, A2 => n11143, ZN => n10536);
   U15364 : AND2_X1 port map( A1 => n10885, A2 => n10886, ZN => n10540);
   U15365 : NOR2_X1 port map( A1 => n10884, A2 => n24345, ZN => n10539);
   U15367 : OR2_X2 port map( A1 => n10546, A2 => n10545, ZN => n11433);
   U15368 : XNOR2_X1 port map( A => n12241, B => n11433, ZN => n11995);
   U15369 : NAND2_X1 port map( A1 => n5107, A2 => n25233, ZN => n10705);
   U15370 : NOR2_X1 port map( A1 => n10951, A2 => n25231, ZN => n10701);
   U15371 : INV_X1 port map( A => n10701, ZN => n10547);
   U15372 : NAND2_X1 port map( A1 => n10955, A2 => n2754, ZN => n10550);
   U15373 : NAND2_X1 port map( A1 => n10548, A2 => n10698, ZN => n10549);
   U15374 : XNOR2_X1 port map( A => n11840, B => n11838, ZN => n12094);
   U15375 : XNOR2_X1 port map( A => n11995, B => n12094, ZN => n10566);
   U15376 : AND2_X1 port map( A1 => n10552, A2 => n11157, ZN => n10554);
   U15377 : NOR2_X1 port map( A1 => n11157, A2 => n11158, ZN => n10555);
   U15378 : NOR2_X1 port map( A1 => n10661, A2 => n10558, ZN => n10562);
   U15379 : OAI21_X1 port map( B1 => n10556, B2 => n10654, A => n25250, ZN => 
                           n10561);
   U15380 : NAND3_X1 port map( A1 => n10558, A2 => n10557, A3 => n10660, ZN => 
                           n10560);
   U15381 : INV_X1 port map( A => n10660, ZN => n10655);
   U15382 : XNOR2_X1 port map( A => n12200, B => n21423, ZN => n10563);
   U15383 : XNOR2_X1 port map( A => n10564, B => n10563, ZN => n10565);
   U15384 : NOR3_X1 port map( A1 => n24373, A2 => n12719, A3 => n13167, ZN => 
                           n10567);
   U15385 : NOR2_X1 port map( A1 => n24373, A2 => n13170, ZN => n13168);
   U15386 : NOR2_X1 port map( A1 => n10567, A2 => n13168, ZN => n10568);
   U15387 : INV_X1 port map( A => n10572, ZN => n10573);
   U15388 : MUX2_X2 port map( A => n10576, B => n10575, S => n10574, Z => 
                           n12019);
   U15389 : XNOR2_X1 port map( A => n12019, B => n12351, ZN => n12302);
   U15390 : MUX2_X1 port map( A => n11171, B => n24957, S => n11178, Z => 
                           n10578);
   U15391 : MUX2_X1 port map( A => n11168, B => n11170, S => n24957, Z => 
                           n10577);
   U15392 : XNOR2_X1 port map( A => n11289, B => n11638, ZN => n10579);
   U15393 : XNOR2_X1 port map( A => n12302, B => n10579, ZN => n10603);
   U15394 : NAND2_X1 port map( A1 => n10585, A2 => n10584, ZN => n10586);
   U15395 : NAND2_X1 port map( A1 => n10589, A2 => n25507, ZN => n10592);
   U15396 : XNOR2_X1 port map( A => n12129, B => n12127, ZN => n10601);
   U15397 : NAND3_X1 port map( A1 => n10934, A2 => n24470, A3 => n10508, ZN => 
                           n10599);
   U15398 : XNOR2_X1 port map( A => n10602, B => n10603, ZN => n13132);
   U15399 : NAND2_X1 port map( A1 => n10605, A2 => n10604, ZN => n10609);
   U15400 : INV_X1 port map( A => n10969, ZN => n10966);
   U15401 : XNOR2_X1 port map( A => n12031, B => n12362, ZN => n12293);
   U15402 : AOI21_X1 port map( B1 => n10613, B2 => n10611, A => n10610, ZN => 
                           n10619);
   U15403 : NAND3_X1 port map( A1 => n10614, A2 => n10613, A3 => n10612, ZN => 
                           n10615);
   U15404 : OAI21_X1 port map( B1 => n10617, B2 => n10616, A => n10615, ZN => 
                           n10618);
   U15406 : NAND3_X1 port map( A1 => n24340, A2 => n3868, A3 => n11216, ZN => 
                           n10625);
   U15407 : XNOR2_X1 port map( A => n12370, B => n10627, ZN => n11986);
   U15408 : XNOR2_X1 port map( A => n11986, B => n12293, ZN => n10640);
   U15409 : NOR2_X1 port map( A1 => n10793, A2 => n11201, ZN => n11204);
   U15410 : OAI21_X1 port map( B1 => n11204, B2 => n11196, A => n11199, ZN => 
                           n10629);
   U15412 : INV_X1 port map( A => n10632, ZN => n11210);
   U15413 : NAND3_X1 port map( A1 => n11205, A2 => n11207, A3 => n11338, ZN => 
                           n10635);
   U15414 : OAI21_X1 port map( B1 => n11205, B2 => n10819, A => n10635, ZN => 
                           n10636);
   U15415 : XNOR2_X1 port map( A => n12167, B => n3164, ZN => n10637);
   U15416 : XNOR2_X1 port map( A => n10638, B => n10637, ZN => n10639);
   U15417 : XNOR2_X1 port map( A => n24980, B => n886, ZN => n10647);
   U15418 : NAND2_X1 port map( A1 => n10642, A2 => n11012, ZN => n10644);
   U15419 : AND2_X1 port map( A1 => n10643, A2 => n10644, ZN => n10645);
   U15420 : INV_X1 port map( A => n12144, ZN => n10646);
   U15421 : NAND2_X1 port map( A1 => n10655, A2 => n10654, ZN => n10656);
   U15422 : XNOR2_X1 port map( A => n12146, B => n12414, ZN => n11991);
   U15423 : INV_X1 port map( A => n11067, ZN => n10667);
   U15424 : AND2_X1 port map( A1 => n11064, A2 => n10662, ZN => n10664);
   U15425 : NOR2_X1 port map( A1 => n11068, A2 => n11067, ZN => n10663);
   U15426 : OAI22_X1 port map( A1 => n10665, A2 => n10664, B1 => n10663, B2 => 
                           n11071, ZN => n10666);
   U15427 : OAI21_X1 port map( B1 => n10667, B2 => n11064, A => n10666, ZN => 
                           n11243);
   U15428 : INV_X1 port map( A => n11243, ZN => n12039);
   U15430 : NAND2_X1 port map( A1 => n11215, A2 => n11216, ZN => n10670);
   U15431 : XNOR2_X1 port map( A => n12152, B => n12322, ZN => n10671);
   U15432 : XNOR2_X1 port map( A => n10672, B => n10671, ZN => n12498);
   U15433 : NAND2_X1 port map( A1 => n11163, A2 => n11158, ZN => n10680);
   U15434 : NAND3_X1 port map( A1 => n10674, A2 => n1453, A3 => n10673, ZN => 
                           n10678);
   U15435 : INV_X1 port map( A => n10675, ZN => n10677);
   U15436 : OAI21_X1 port map( B1 => n10678, B2 => n10677, A => n10676, ZN => 
                           n10679);
   U15437 : INV_X1 port map( A => n11007, ZN => n10688);
   U15438 : OAI211_X1 port map( C1 => n2306, C2 => n24420, A => n24622, B => 
                           n10681, ZN => n10687);
   U15439 : INV_X1 port map( A => n10682, ZN => n10684);
   U15440 : NAND2_X1 port map( A1 => n11006, A2 => n10685, ZN => n10686);
   U15441 : XNOR2_X1 port map( A => n11717, B => n10689, ZN => n12156);
   U15442 : NAND2_X1 port map( A1 => n11149, A2 => n11151, ZN => n11888);
   U15443 : NAND3_X1 port map( A1 => n714, A2 => n11884, A3 => n11143, ZN => 
                           n10692);
   U15444 : NAND3_X1 port map( A1 => n10690, A2 => n11147, A3 => n11885, ZN => 
                           n10691);
   U15445 : NAND3_X1 port map( A1 => n11888, A2 => n10692, A3 => n10691, ZN => 
                           n11247);
   U15446 : XNOR2_X1 port map( A => n11247, B => n11746, ZN => n12311);
   U15447 : XNOR2_X1 port map( A => n12156, B => n12311, ZN => n10709);
   U15448 : NAND2_X1 port map( A1 => n11054, A2 => n11499, ZN => n10696);
   U15449 : NOR2_X1 port map( A1 => n11057, A2 => n11009, ZN => n10693);
   U15450 : NAND2_X1 port map( A1 => n11059, A2 => n10693, ZN => n10695);
   U15451 : INV_X1 port map( A => n11499, ZN => n11053);
   U15452 : INV_X1 port map( A => n10698, ZN => n10954);
   U15453 : XNOR2_X1 port map( A => n10707, B => n10706, ZN => n10708);
   U15454 : NOR2_X1 port map( A1 => n12498, A2 => n13130, ZN => n10710);
   U15455 : NOR2_X1 port map( A1 => n5754, A2 => n10710, ZN => n12426);
   U15456 : INV_X1 port map( A => n12663, ZN => n10711);
   U15457 : NAND2_X1 port map( A1 => n10713, A2 => n10712, ZN => n10718);
   U15459 : NAND3_X1 port map( A1 => n10838, A2 => n420, A3 => n10714, ZN => 
                           n10715);
   U15460 : NAND4_X2 port map( A1 => n10716, A2 => n10717, A3 => n10715, A4 => 
                           n10718, ZN => n11795);
   U15461 : XNOR2_X1 port map( A => n11795, B => n2005, ZN => n10719);
   U15463 : AND2_X1 port map( A1 => n10720, A2 => n11121, ZN => n10721);
   U15465 : NAND2_X1 port map( A1 => n11110, A2 => n10875, ZN => n10726);
   U15466 : MUX2_X1 port map( A => n10729, B => n10728, S => n11190, Z => 
                           n10735);
   U15467 : NAND2_X1 port map( A1 => n11184, A2 => n10729, ZN => n10733);
   U15468 : NAND3_X1 port map( A1 => n10731, A2 => n10730, A3 => n10734, ZN => 
                           n10732);
   U15469 : XNOR2_X1 port map( A => n12404, B => n25236, ZN => n11981);
   U15470 : AND2_X1 port map( A1 => n10860, A2 => n25230, ZN => n10739);
   U15471 : NOR2_X1 port map( A1 => n10861, A2 => n25230, ZN => n10738);
   U15472 : AOI22_X1 port map( A1 => n10739, A2 => n10740, B1 => n10738, B2 => 
                           n10737, ZN => n10742);
   U15473 : NAND3_X1 port map( A1 => n10740, A2 => n10855, A3 => n10861, ZN => 
                           n10741);
   U15474 : XNOR2_X1 port map( A => n12066, B => n11756, ZN => n12338);
   U15475 : XNOR2_X1 port map( A => n11981, B => n12338, ZN => n10744);
   U15476 : INV_X1 port map( A => n13150, ZN => n13157);
   U15477 : NOR2_X1 port map( A1 => n10904, A2 => n10907, ZN => n10748);
   U15478 : AOI22_X1 port map( A1 => n10749, A2 => n10751, B1 => n10748, B2 => 
                           n10905, ZN => n10750);
   U15479 : NOR2_X1 port map( A1 => n10753, A2 => n10752, ZN => n10754);
   U15480 : INV_X1 port map( A => n10756, ZN => n10758);
   U15481 : NOR2_X2 port map( A1 => n10761, A2 => n10760, ZN => n11581);
   U15482 : INV_X1 port map( A => n11301, ZN => n11089);
   U15483 : INV_X1 port map( A => n10762, ZN => n11305);
   U15484 : MUX2_X1 port map( A => n10764, B => n10763, S => n11091, Z => 
                           n10765);
   U15485 : XNOR2_X1 port map( A => n11581, B => n12375, ZN => n11996);
   U15486 : XNOR2_X1 port map( A => n12341, B => n11996, ZN => n10786);
   U15487 : NOR2_X1 port map( A1 => n11084, A2 => n10891, ZN => n10768);
   U15488 : NOR2_X2 port map( A1 => n10770, A2 => n10769, ZN => n12121);
   U15489 : XNOR2_X1 port map( A => n10771, B => n12121, ZN => n10784);
   U15490 : OAI21_X1 port map( B1 => n11101, B2 => n10911, A => n10772, ZN => 
                           n10781);
   U15491 : INV_X1 port map( A => n10773, ZN => n10774);
   U15492 : NOR2_X1 port map( A1 => n10775, A2 => n10774, ZN => n10777);
   U15493 : NAND4_X1 port map( A1 => n10778, A2 => n415, A3 => n10777, A4 => 
                           n10776, ZN => n10780);
   U15494 : OAI211_X2 port map( C1 => n10781, C2 => n10782, A => n10780, B => 
                           n10779, ZN => n11765);
   U15495 : XNOR2_X1 port map( A => n11765, B => n2805, ZN => n10783);
   U15496 : XNOR2_X1 port map( A => n10784, B => n10783, ZN => n10785);
   U15497 : XNOR2_X1 port map( A => n10786, B => n10785, ZN => n13151);
   U15499 : OAI211_X1 port map( C1 => n13157, C2 => n13152, A => n13148, B => 
                           n13130, ZN => n10787);
   U15500 : NAND2_X1 port map( A1 => n10788, A2 => n11195, ZN => n10797);
   U15501 : INV_X1 port map( A => n10789, ZN => n10790);
   U15502 : INV_X1 port map( A => n11196, ZN => n10792);
   U15503 : NAND3_X1 port map( A1 => n11201, A2 => n11199, A3 => n10792, ZN => 
                           n10795);
   U15504 : NAND3_X1 port map( A1 => n10793, A2 => n11196, A3 => n11199, ZN => 
                           n10794);
   U15505 : XNOR2_X1 port map( A => n11951, B => n12401, ZN => n10809);
   U15506 : MUX2_X1 port map( A => n10800, B => n10799, S => n10798, Z => 
                           n10802);
   U15507 : MUX2_X1 port map( A => n10803, B => n10802, S => n10801, Z => 
                           n10807);
   U15508 : NOR2_X2 port map( A1 => n10807, A2 => n10806, ZN => n12334);
   U15509 : INV_X1 port map( A => n12334, ZN => n10808);
   U15510 : XNOR2_X1 port map( A => n10809, B => n10808, ZN => n10828);
   U15512 : XNOR2_X1 port map( A => n11619, B => n25236, ZN => n10826);
   U15513 : NOR2_X1 port map( A1 => n10967, A2 => n10969, ZN => n10815);
   U15514 : NOR2_X1 port map( A1 => n10970, A2 => n10968, ZN => n10814);
   U15515 : NAND2_X1 port map( A1 => n10816, A2 => n10970, ZN => n10817);
   U15516 : XNOR2_X1 port map( A => n12112, B => n2903, ZN => n10824);
   U15517 : MUX2_X1 port map( A => n11342, B => n10819, S => n25025, Z => 
                           n10823);
   U15518 : INV_X1 port map( A => n11205, ZN => n11339);
   U15519 : NAND2_X1 port map( A1 => n11342, A2 => n11207, ZN => n10820);
   U15520 : MUX2_X1 port map( A => n10821, B => n10820, S => n10819, Z => 
                           n10822);
   U15521 : OAI21_X2 port map( B1 => n10823, B2 => n11339, A => n10822, ZN => 
                           n12397);
   U15522 : XNOR2_X1 port map( A => n10824, B => n12397, ZN => n10825);
   U15523 : XNOR2_X1 port map( A => n10825, B => n10826, ZN => n10827);
   U15524 : XNOR2_X1 port map( A => n10827, B => n10828, ZN => n12740);
   U15525 : INV_X1 port map( A => n12740, ZN => n13101);
   U15526 : AOI22_X1 port map( A1 => n10836, A2 => n10834, B1 => n10833, B2 => 
                           n10832, ZN => n10835);
   U15527 : OAI21_X1 port map( B1 => n10837, B2 => n10836, A => n10835, ZN => 
                           n12344);
   U15528 : XNOR2_X1 port map( A => n12344, B => n11581, ZN => n11666);
   U15529 : NAND2_X1 port map( A1 => n10841, A2 => n11129, ZN => n10842);
   U15530 : XNOR2_X1 port map( A => n12381, B => n1951, ZN => n10845);
   U15531 : XNOR2_X1 port map( A => n11666, B => n10845, ZN => n10883);
   U15532 : OR2_X1 port map( A1 => n10848, A2 => n2244, ZN => n10849);
   U15533 : OAI211_X1 port map( C1 => n11125, C2 => n10850, A => n10849, B => 
                           n11124, ZN => n10852);
   U15534 : NAND3_X1 port map( A1 => n10856, A2 => n10855, A3 => n10854, ZN => 
                           n10866);
   U15536 : NAND2_X1 port map( A1 => n10862, A2 => n10861, ZN => n10863);
   U15537 : XNOR2_X1 port map( A => n11703, B => n12096, ZN => n11602);
   U15539 : NAND4_X1 port map( A1 => n10873, A2 => n10870, A3 => n10867, A4 => 
                           n9340, ZN => n11115);
   U15540 : INV_X1 port map( A => n10870, ZN => n10872);
   U15541 : NOR2_X1 port map( A1 => n10872, A2 => n10871, ZN => n10874);
   U15542 : NAND4_X1 port map( A1 => n10875, A2 => n1494, A3 => n10874, A4 => 
                           n10873, ZN => n10876);
   U15543 : OAI21_X2 port map( B1 => n10877, B2 => n10878, A => n10876, ZN => 
                           n11766);
   U15544 : INV_X1 port map( A => n12383, ZN => n10879);
   U15545 : XNOR2_X1 port map( A => n10879, B => n11766, ZN => n10880);
   U15547 : MUX2_X1 port map( A => n10887, B => n10886, S => n10885, Z => 
                           n10888);
   U15548 : XNOR2_X1 port map( A => n12306, B => n12127, ZN => n11639);
   U15549 : INV_X1 port map( A => n11966, ZN => n11457);
   U15550 : INV_X1 port map( A => n11086, ZN => n10893);
   U15551 : NOR2_X1 port map( A1 => n11085, A2 => n10891, ZN => n10892);
   U15552 : XNOR2_X1 port map( A => n11457, B => n12020, ZN => n12354);
   U15553 : NAND2_X1 port map( A1 => n11302, A2 => n11298, ZN => n10897);
   U15554 : OAI21_X1 port map( B1 => n10902, B2 => n10901, A => n10900, ZN => 
                           n10909);
   U15555 : OAI21_X1 port map( B1 => n10905, B2 => n10904, A => n10903, ZN => 
                           n10906);
   U15556 : INV_X1 port map( A => n10906, ZN => n10908);
   U15558 : XNOR2_X1 port map( A => n11627, B => n12183, ZN => n10916);
   U15559 : NAND3_X1 port map( A1 => n11099, A2 => n10911, A3 => n11101, ZN => 
                           n10912);
   U15560 : INV_X1 port map( A => n2795, ZN => n23191);
   U15561 : XNOR2_X1 port map( A => n12357, B => n23191, ZN => n10915);
   U15562 : XNOR2_X1 port map( A => n10916, B => n10915, ZN => n10917);
   U15563 : MUX2_X1 port map( A => n13101, B => n13102, S => n13185, Z => 
                           n11021);
   U15564 : NAND2_X1 port map( A1 => n10922, A2 => n11520, ZN => n10919);
   U15566 : INV_X1 port map( A => n2991, ZN => n21079);
   U15567 : XNOR2_X1 port map( A => n12388, B => n21079, ZN => n10923);
   U15568 : INV_X1 port map( A => n11747, ZN => n11942);
   U15569 : NAND2_X1 port map( A1 => n10925, A2 => n10924, ZN => n10929);
   U15570 : OAI21_X1 port map( B1 => n10927, B2 => n10990, A => n10926, ZN => 
                           n10928);
   U15571 : INV_X1 port map( A => n10931, ZN => n10932);
   U15572 : NAND2_X1 port map( A1 => n10932, A2 => n10935, ZN => n10933);
   U15573 : OAI21_X1 port map( B1 => n11171, B2 => n11175, A => n10937, ZN => 
                           n10938);
   U15574 : XNOR2_X1 port map( A => n11749, B => n12389, ZN => n10947);
   U15575 : INV_X1 port map( A => n11040, ZN => n10946);
   U15576 : NAND2_X1 port map( A1 => n416, A2 => n10942, ZN => n10943);
   U15577 : XNOR2_X1 port map( A => n10947, B => n24915, ZN => n10948);
   U15578 : XNOR2_X1 port map( A => n10949, B => n10948, ZN => n13187);
   U15579 : NAND3_X1 port map( A1 => n10955, A2 => n10954, A3 => n25232, ZN => 
                           n10956);
   U15581 : XNOR2_X1 port map( A => n24401, B => n812, ZN => n10959);
   U15582 : INV_X1 port map( A => n12146, ZN => n11555);
   U15583 : XNOR2_X1 port map( A => n10959, B => n11555, ZN => n10977);
   U15584 : NAND2_X1 port map( A1 => n714, A2 => n24480, ZN => n10964);
   U15585 : NOR2_X1 port map( A1 => n10961, A2 => n11884, ZN => n10960);
   U15587 : INV_X1 port map( A => n10961, ZN => n11148);
   U15588 : NOR2_X1 port map( A1 => n25497, A2 => n10969, ZN => n10976);
   U15589 : OAI21_X1 port map( B1 => n10967, B2 => n10966, A => n10497, ZN => 
                           n10975);
   U15590 : NAND2_X1 port map( A1 => n10969, A2 => n10968, ZN => n10973);
   U15591 : INV_X1 port map( A => n10970, ZN => n10972);
   U15592 : MUX2_X1 port map( A => n10973, B => n10972, S => n25497, Z => 
                           n10974);
   U15593 : XNOR2_X1 port map( A => n11897, B => n12325, ZN => n12210);
   U15594 : XNOR2_X1 port map( A => n10977, B => n12210, ZN => n10988);
   U15595 : NOR2_X1 port map( A1 => n11059, A2 => n11052, ZN => n11498);
   U15596 : NOR2_X1 port map( A1 => n10978, A2 => n11498, ZN => n10981);
   U15597 : AOI21_X1 port map( B1 => n11054, B2 => n11009, A => n11053, ZN => 
                           n10979);
   U15598 : OAI21_X1 port map( B1 => n11009, B2 => n410, A => n10979, ZN => 
                           n10980);
   U15599 : NAND2_X1 port map( A1 => n417, A2 => n11157, ZN => n11166);
   U15600 : NOR2_X1 port map( A1 => n4737, A2 => n11157, ZN => n10982);
   U15601 : AOI22_X1 port map( A1 => n10982, A2 => n10985, B1 => n11158, B2 => 
                           n11157, ZN => n10984);
   U15602 : NAND3_X1 port map( A1 => n417, A2 => n10985, A3 => n11160, ZN => 
                           n10983);
   U15603 : OAI211_X2 port map( C1 => n11166, C2 => n10985, A => n10984, B => 
                           n10983, ZN => n12413);
   U15604 : XNOR2_X1 port map( A => n11960, B => n12413, ZN => n10986);
   U15605 : XNOR2_X1 port map( A => n12410, B => n10986, ZN => n10987);
   U15606 : NOR2_X1 port map( A1 => n10989, A2 => n10994, ZN => n10991);
   U15607 : OAI21_X1 port map( B1 => n10992, B2 => n10991, A => n10990, ZN => 
                           n10999);
   U15608 : NOR3_X1 port map( A1 => n24118, A2 => n3606, A3 => n10993, ZN => 
                           n10997);
   U15609 : NOR2_X1 port map( A1 => n10997, A2 => n10996, ZN => n10998);
   U15610 : NAND3_X1 port map( A1 => n11068, A2 => n11069, A3 => n11064, ZN => 
                           n11000);
   U15611 : XNOR2_X1 port map( A => n11907, B => n25234, ZN => n11608);
   U15612 : XNOR2_X1 port map( A => n11563, B => n12295, ZN => n11648);
   U15613 : XNOR2_X1 port map( A => n11608, B => n11648, ZN => n11019);
   U15614 : XNOR2_X1 port map( A => n11736, B => n19392, ZN => n11017);
   U15615 : AOI21_X1 port map( B1 => n11010, B2 => n11050, A => n11046, ZN => 
                           n11015);
   U15616 : AOI21_X1 port map( B1 => n11013, B2 => n11012, A => n11044, ZN => 
                           n11014);
   U15617 : NOR2_X2 port map( A1 => n11015, A2 => n11014, ZN => n12363);
   U15618 : XNOR2_X1 port map( A => n12363, B => n25371, ZN => n11016);
   U15619 : XNOR2_X1 port map( A => n11017, B => n11016, ZN => n11018);
   U15622 : NAND3_X1 port map( A1 => n11026, A2 => n11525, A3 => n25060, ZN => 
                           n11028);
   U15623 : NAND3_X1 port map( A1 => n11529, A2 => n1332, A3 => n11524, ZN => 
                           n11027);
   U15624 : XNOR2_X1 port map( A => n12234, B => n17960, ZN => n11030);
   U15625 : XNOR2_X1 port map( A => n12249, B => n12297, ZN => n11029);
   U15626 : XNOR2_X1 port map( A => n11030, B => n11029, ZN => n11043);
   U15627 : XNOR2_X1 port map( A => n12233, B => n11561, ZN => n11692);
   U15628 : XNOR2_X1 port map( A => n11983, B => n12365, ZN => n11041);
   U15629 : XNOR2_X1 port map( A => n11692, B => n11041, ZN => n11042);
   U15630 : XNOR2_X2 port map( A => n11042, B => n11043, ZN => n13144);
   U15631 : INV_X1 port map( A => n13144, ZN => n13138);
   U15632 : OAI21_X1 port map( B1 => n11045, B2 => n4531, A => n11044, ZN => 
                           n11048);
   U15633 : NAND3_X1 port map( A1 => n11059, A2 => n11053, A3 => n11052, ZN => 
                           n11056);
   U15634 : XNOR2_X1 port map( A => n12197, B => n11706, ZN => n11060);
   U15635 : XNOR2_X1 port map( A => n11060, B => n11061, ZN => n11080);
   U15636 : NAND2_X1 port map( A1 => n10347, A2 => n11064, ZN => n11066);
   U15637 : OR3_X1 port map( A1 => n11064, A2 => n25203, A3 => n11062, ZN => 
                           n11065);
   U15639 : NAND2_X1 port map( A1 => n11068, A2 => n11067, ZN => n11073);
   U15640 : NAND2_X1 port map( A1 => n11070, A2 => n11069, ZN => n11072);
   U15641 : AOI21_X1 port map( B1 => n11073, B2 => n11072, A => n11071, ZN => 
                           n11074);
   U15642 : INV_X1 port map( A => n11076, ZN => n12343);
   U15643 : XNOR2_X1 port map( A => n12343, B => n12196, ZN => n11078);
   U15644 : XNOR2_X1 port map( A => n12200, B => n688, ZN => n11077);
   U15645 : XNOR2_X1 port map( A => n11078, B => n11077, ZN => n11079);
   U15646 : XNOR2_X1 port map( A => n11079, B => n11080, ZN => n13140);
   U15647 : INV_X1 port map( A => n13140, ZN => n12728);
   U15648 : NOR2_X1 port map( A1 => n3119, A2 => n11081, ZN => n11083);
   U15649 : XNOR2_X1 port map( A => n11087, B => n11088, ZN => n11108);
   U15650 : OAI21_X1 port map( B1 => n11089, B2 => n11092, A => n419, ZN => 
                           n11095);
   U15651 : OAI211_X1 port map( C1 => n11090, C2 => n11091, A => n11305, B => 
                           n11298, ZN => n11094);
   U15652 : NOR2_X1 port map( A1 => n11092, A2 => n11091, ZN => n11093);
   U15653 : XNOR2_X1 port map( A => n24027, B => n12209, ZN => n11900);
   U15654 : NAND2_X1 port map( A1 => n11096, A2 => n1552, ZN => n11098);
   U15655 : NAND2_X1 port map( A1 => n11099, A2 => n415, ZN => n11097);
   U15657 : NAND2_X1 port map( A1 => n11100, A2 => n11099, ZN => n11104);
   U15658 : XNOR2_X1 port map( A => n12212, B => n1754, ZN => n11106);
   U15659 : XNOR2_X1 port map( A => n11900, B => n11106, ZN => n11107);
   U15660 : XNOR2_X1 port map( A => n11108, B => n11107, ZN => n11109);
   U15661 : NAND2_X1 port map( A1 => n12728, A2 => n11109, ZN => n12437);
   U15662 : AOI21_X1 port map( B1 => n11117, B2 => n11111, A => n11110, ZN => 
                           n11120);
   U15663 : AOI21_X1 port map( B1 => n11116, B2 => n11112, A => n11113, ZN => 
                           n11119);
   U15664 : OAI211_X1 port map( C1 => n11117, C2 => n11116, A => n11115, B => 
                           n11114, ZN => n11118);
   U15665 : XNOR2_X1 port map( A => n12314, B => n11715, ZN => n11137);
   U15666 : AOI22_X1 port map( A1 => n11126, A2 => n11125, B1 => n11124, B2 => 
                           n11123, ZN => n11127);
   U15667 : NOR2_X1 port map( A1 => n11129, A2 => n11128, ZN => n11134);
   U15668 : INV_X1 port map( A => n11131, ZN => n11132);
   U15669 : OAI211_X2 port map( C1 => n11135, C2 => n11134, A => n11133, B => 
                           n11132, ZN => n12221);
   U15670 : XNOR2_X1 port map( A => n12221, B => n12219, ZN => n11136);
   U15671 : XNOR2_X1 port map( A => n11137, B => n11136, ZN => n11141);
   U15672 : XNOR2_X1 port map( A => n12391, B => n12224, ZN => n11139);
   U15673 : XNOR2_X1 port map( A => n12255, B => n1869, ZN => n11138);
   U15674 : XNOR2_X1 port map( A => n11139, B => n11138, ZN => n11140);
   U15675 : XNOR2_X1 port map( A => n11141, B => n11140, ZN => n13136);
   U15676 : INV_X1 port map( A => n13136, ZN => n13143);
   U15677 : NAND2_X1 port map( A1 => n13139, A2 => n13143, ZN => n11142);
   U15679 : NAND3_X1 port map( A1 => n11145, A2 => n11146, A3 => n11143, ZN => 
                           n11144);
   U15680 : OAI21_X1 port map( B1 => n11147, B2 => n11145, A => n11144, ZN => 
                           n11156);
   U15681 : OAI21_X1 port map( B1 => n11147, B2 => n11146, A => n4998, ZN => 
                           n11155);
   U15682 : NOR2_X1 port map( A1 => n11148, A2 => n11151, ZN => n11150);
   U15683 : NAND2_X1 port map( A1 => n11150, A2 => n11149, ZN => n11154);
   U15684 : NAND3_X1 port map( A1 => n714, A2 => n24479, A3 => n11151, ZN => 
                           n11153);
   U15685 : NOR2_X1 port map( A1 => n1358, A2 => n11157, ZN => n11162);
   U15686 : NOR2_X1 port map( A1 => n11159, A2 => n11158, ZN => n11161);
   U15687 : OAI21_X1 port map( B1 => n11162, B2 => n11161, A => n11160, ZN => 
                           n11165);
   U15688 : XNOR2_X1 port map( A => n12065, B => n11977, ZN => n12193);
   U15689 : XNOR2_X1 port map( A => n11167, B => n12193, ZN => n11183);
   U15691 : AND2_X1 port map( A1 => n11171, A2 => n1338, ZN => n11173);
   U15692 : NAND2_X1 port map( A1 => n11178, A2 => n11173, ZN => n11177);
   U15693 : OAI211_X2 port map( C1 => n11179, C2 => n11178, A => n11177, B => 
                           n11176, ZN => n11689);
   U15696 : XNOR2_X1 port map( A => n11181, B => n11180, ZN => n11182);
   U15698 : NAND2_X1 port map( A1 => n13138, A2 => n12455, ZN => n11222);
   U15699 : INV_X1 port map( A => n11370, ZN => n11191);
   U15700 : INV_X1 port map( A => n11184, ZN => n11187);
   U15701 : INV_X1 port map( A => n11185, ZN => n11186);
   U15702 : NAND2_X1 port map( A1 => n11187, A2 => n11186, ZN => n11188);
   U15703 : OAI22_X1 port map( A1 => n11191, A2 => n11190, B1 => n11189, B2 => 
                           n11188, ZN => n11192);
   U15704 : XNOR2_X1 port map( A => n11192, B => n2990, ZN => n11193);
   U15705 : XNOR2_X1 port map( A => n11194, B => n11193, ZN => n11221);
   U15706 : INV_X1 port map( A => n11201, ZN => n11197);
   U15707 : OAI21_X1 port map( B1 => n11197, B2 => n11196, A => n10790, ZN => 
                           n11203);
   U15709 : NAND2_X1 port map( A1 => n25025, A2 => n11205, ZN => n11206);
   U15710 : NAND2_X1 port map( A1 => n11210, A2 => n11207, ZN => n11208);
   U15711 : MUX2_X1 port map( A => n11214, B => n24340, S => n11212, Z => 
                           n11219);
   U15712 : XNOR2_X1 port map( A => n12181, B => n11880, ZN => n11220);
   U15713 : XNOR2_X1 port map( A => n11220, B => n11221, ZN => n12433);
   U15715 : INV_X1 port map( A => n14156, ZN => n13780);
   U15717 : XNOR2_X1 port map( A => n12189, B => n12397, ZN => n12064);
   U15718 : XNOR2_X1 port map( A => n11619, B => n11795, ZN => n11759);
   U15719 : XNOR2_X1 port map( A => n12064, B => n11759, ZN => n11227);
   U15720 : XNOR2_X1 port map( A => n12066, B => n12401, ZN => n11816);
   U15721 : INV_X1 port map( A => n23476, ZN => n20840);
   U15722 : XNOR2_X1 port map( A => n11816, B => n11225, ZN => n11226);
   U15723 : XNOR2_X1 port map( A => n11227, B => n11226, ZN => n12541);
   U15724 : XNOR2_X1 port map( A => n12031, B => n12363, ZN => n11833);
   U15725 : INV_X1 port map( A => n11833, ZN => n11228);
   U15726 : XNOR2_X1 port map( A => n12248, B => n25234, ZN => n12030);
   U15727 : XNOR2_X1 port map( A => n11228, B => n12030, ZN => n11231);
   U15728 : XNOR2_X1 port map( A => n12233, B => n11736, ZN => n11535);
   U15729 : XNOR2_X1 port map( A => n11735, B => n20690, ZN => n11229);
   U15730 : XNOR2_X1 port map( A => n11535, B => n11229, ZN => n11230);
   U15731 : INV_X1 port map( A => n11703, ZN => n12377);
   U15732 : XNOR2_X1 port map( A => n12377, B => n11766, ZN => n11232);
   U15733 : XNOR2_X1 port map( A => n11232, B => n11812, ZN => n11236);
   U15734 : XNOR2_X1 port map( A => n11765, B => n12201, ZN => n11234);
   U15735 : XNOR2_X1 port map( A => n12200, B => n881, ZN => n11233);
   U15736 : XNOR2_X1 port map( A => n11234, B => n11233, ZN => n11235);
   U15737 : XNOR2_X1 port map( A => n11627, B => n11638, ZN => n11724);
   U15738 : XNOR2_X1 port map( A => n12019, B => n12357, ZN => n11456);
   U15739 : XNOR2_X1 port map( A => n11456, B => n11724, ZN => n11241);
   U15740 : XNOR2_X1 port map( A => n12184, B => n12020, ZN => n11239);
   U15741 : INV_X1 port map( A => n11237, ZN => n12180);
   U15742 : XNOR2_X1 port map( A => n12180, B => n1865, ZN => n11238);
   U15743 : XNOR2_X1 port map( A => n11239, B => n11238, ZN => n11240);
   U15744 : XNOR2_X1 port map( A => n11240, B => n11241, ZN => n12540);
   U15745 : XNOR2_X1 port map( A => n24401, B => n11242, ZN => n11745);
   U15746 : XNOR2_X1 port map( A => n12410, B => n11243, ZN => n11822);
   U15747 : XNOR2_X1 port map( A => n11822, B => n11745, ZN => n11246);
   U15748 : XNOR2_X1 port map( A => n12209, B => n3118, ZN => n11244);
   U15749 : XNOR2_X1 port map( A => n12413, B => n12207, ZN => n12038);
   U15750 : XNOR2_X1 port map( A => n12038, B => n11244, ZN => n11245);
   U15751 : XNOR2_X1 port map( A => n12218, B => n12388, ZN => n11718);
   U15752 : XNOR2_X1 port map( A => n11718, B => n11827, ZN => n11250);
   U15753 : XNOR2_X1 port map( A => n11749, B => n12224, ZN => n11545);
   U15754 : XNOR2_X1 port map( A => n11248, B => n11545, ZN => n11249);
   U15755 : MUX2_X1 port map( A => n13217, B => n13216, S => n12767, Z => 
                           n11251);
   U15756 : NOR2_X1 port map( A1 => n11251, A2 => n24512, ZN => n11252);
   U15757 : XNOR2_X1 port map( A => n11253, B => n11914, ZN => n11842);
   U15758 : XNOR2_X1 port map( A => n12096, B => n11582, ZN => n12198);
   U15759 : XNOR2_X1 port map( A => n11842, B => n12198, ZN => n11257);
   U15760 : XNOR2_X1 port map( A => n11838, B => n1831, ZN => n11255);
   U15761 : XNOR2_X1 port map( A => n11704, B => n12381, ZN => n11254);
   U15762 : XNOR2_X1 port map( A => n11255, B => n11254, ZN => n11256);
   U15763 : XNOR2_X1 port map( A => n12249, B => n11776, ZN => n11905);
   U15764 : XNOR2_X1 port map( A => n11607, B => n11907, ZN => n11693);
   U15765 : XNOR2_X1 port map( A => n11693, B => n11905, ZN => n11261);
   U15766 : XNOR2_X1 port map( A => n12363, B => n3062, ZN => n11259);
   U15767 : XNOR2_X1 port map( A => n11646, B => n11564, ZN => n11258);
   U15768 : XNOR2_X1 port map( A => n11259, B => n11258, ZN => n11260);
   U15769 : XNOR2_X1 port map( A => n11261, B => n11260, ZN => n11287);
   U15770 : INV_X1 port map( A => n11616, ZN => n11262);
   U15771 : XNOR2_X1 port map( A => n12226, B => n11262, ZN => n11716);
   U15772 : XNOR2_X1 port map( A => n12313, B => n12255, ZN => n11893);
   U15773 : XNOR2_X1 port map( A => n11716, B => n11893, ZN => n11267);
   U15774 : XNOR2_X1 port map( A => n11659, B => n12389, ZN => n11265);
   U15775 : XNOR2_X1 port map( A => n12225, B => n681, ZN => n11264);
   U15776 : XNOR2_X1 port map( A => n11265, B => n11264, ZN => n11266);
   U15777 : XNOR2_X1 port map( A => n11267, B => n11266, ZN => n13011);
   U15778 : XNOR2_X1 port map( A => n12186, B => n11640, ZN => n11269);
   U15779 : XNOR2_X1 port map( A => n11268, B => n11492, ZN => n11878);
   U15780 : INV_X1 port map( A => n11878, ZN => n11858);
   U15781 : XNOR2_X1 port map( A => n11858, B => n11269, ZN => n11273);
   U15782 : XNOR2_X1 port map( A => n12183, B => n12357, ZN => n11271);
   U15783 : XNOR2_X1 port map( A => n11698, B => n1745, ZN => n11270);
   U15784 : XNOR2_X1 port map( A => n11271, B => n11270, ZN => n11272);
   U15785 : INV_X1 port map( A => n13013, ZN => n13017);
   U15787 : XNOR2_X1 port map( A => n12333, B => n12275, ZN => n11924);
   U15788 : INV_X1 port map( A => n11924, ZN => n11275);
   U15789 : XNOR2_X1 port map( A => n25027, B => n11274, ZN => n12190);
   U15790 : XNOR2_X1 port map( A => n11275, B => n12190, ZN => n11279);
   U15791 : INV_X1 port map( A => n11686, ZN => n11618);
   U15792 : XNOR2_X1 port map( A => n11672, B => n11618, ZN => n11277);
   U15793 : XNOR2_X1 port map( A => n12401, B => n2100, ZN => n11276);
   U15794 : XNOR2_X1 port map( A => n11277, B => n11276, ZN => n11278);
   U15795 : XNOR2_X2 port map( A => n11279, B => n11278, ZN => n13245);
   U15796 : XNOR2_X1 port map( A => n12101, B => n2050, ZN => n11280);
   U15797 : XNOR2_X1 port map( A => n11280, B => n12410, ZN => n11283);
   U15798 : INV_X1 port map( A => n11653, ZN => n11281);
   U15799 : XNOR2_X1 port map( A => n12283, B => n11281, ZN => n11282);
   U15800 : XNOR2_X1 port map( A => n11282, B => n11283, ZN => n11286);
   U15801 : INV_X1 port map( A => n11284, ZN => n11285);
   U15802 : XNOR2_X1 port map( A => n11285, B => n11286, ZN => n12560);
   U15803 : INV_X1 port map( A => n12560, ZN => n12808);
   U15804 : NOR2_X1 port map( A1 => n25199, A2 => n13246, ZN => n11288);
   U15805 : XNOR2_X1 port map( A => n12003, B => n11289, ZN => n12074);
   U15807 : XNOR2_X1 port map( A => n11637, B => n11568, ZN => n11439);
   U15808 : XNOR2_X1 port map( A => n24990, B => n11439, ZN => n11293);
   U15809 : XNOR2_X1 port map( A => n12023, B => n12128, ZN => n11856);
   U15810 : XNOR2_X1 port map( A => n11698, B => n1364, ZN => n11291);
   U15811 : XNOR2_X1 port map( A => n11856, B => n11291, ZN => n11292);
   U15812 : XNOR2_X1 port map( A => n11292, B => n11293, ZN => n13228);
   U15814 : XNOR2_X1 port map( A => n11689, B => n729, ZN => n11294);
   U15815 : XNOR2_X1 port map( A => n11294, B => n11618, ZN => n11296);
   U15816 : XNOR2_X1 port map( A => n11296, B => n12114, ZN => n11309);
   U15817 : NOR2_X1 port map( A1 => n11302, A2 => n11301, ZN => n11303);
   U15818 : NAND2_X1 port map( A1 => n11303, A2 => n11305, ZN => n11304);
   U15819 : XNOR2_X1 port map( A => n12065, B => n12134, ZN => n11868);
   U15820 : XNOR2_X1 port map( A => n25090, B => n11561, ZN => n11413);
   U15821 : XNOR2_X1 port map( A => n12088, B => n11413, ZN => n11313);
   U15822 : XNOR2_X1 port map( A => n11607, B => n2745, ZN => n11311);
   U15823 : XNOR2_X1 port map( A => n11851, B => n11311, ZN => n11312);
   U15824 : INV_X1 port map( A => n12197, ZN => n11314);
   U15825 : XNOR2_X1 port map( A => n11314, B => n12122, ZN => n11510);
   U15826 : INV_X1 port map( A => n11510, ZN => n11839);
   U15827 : XNOR2_X1 port map( A => n11839, B => n12095, ZN => n11318);
   U15828 : XNOR2_X1 port map( A => n11704, B => n11706, ZN => n11316);
   U15829 : XNOR2_X1 port map( A => n11316, B => n11315, ZN => n11317);
   U15830 : NOR2_X1 port map( A1 => n12993, A2 => n24750, ZN => n11319);
   U15832 : XNOR2_X1 port map( A => n25087, B => n11959, ZN => n11320);
   U15833 : XNOR2_X1 port map( A => n12151, B => n12212, ZN => n11516);
   U15834 : INV_X1 port map( A => n11516, ZN => n11849);
   U15835 : INV_X1 port map( A => n11782, ZN => n11322);
   U15836 : XNOR2_X1 port map( A => n12214, B => n11322, ZN => n12106);
   U15837 : INV_X1 port map( A => n12159, ZN => n12260);
   U15838 : XNOR2_X1 port map( A => n12221, B => n12260, ZN => n11863);
   U15840 : XNOR2_X1 port map( A => n11616, B => n21964, ZN => n11324);
   U15841 : XNOR2_X1 port map( A => n25048, B => n11324, ZN => n11327);
   U15842 : XNOR2_X1 port map( A => n11715, B => n11660, ZN => n11426);
   U15843 : XNOR2_X1 port map( A => n11787, B => n11426, ZN => n11326);
   U15844 : NOR2_X1 port map( A1 => n4587, A2 => n12791, ZN => n11329);
   U15845 : NAND2_X1 port map( A1 => n11329, A2 => n25080, ZN => n11330);
   U15846 : INV_X1 port map( A => n11771, ZN => n11879);
   U15847 : XNOR2_X1 port map( A => n11879, B => n12130, ZN => n12267);
   U15848 : XNOR2_X1 port map( A => n11628, B => n11440, ZN => n11332);
   U15849 : XNOR2_X1 port map( A => n12267, B => n11332, ZN => n11335);
   U15850 : XNOR2_X1 port map( A => n12355, B => n12127, ZN => n11570);
   U15851 : XNOR2_X1 port map( A => n12023, B => n1801, ZN => n11333);
   U15852 : XNOR2_X1 port map( A => n11570, B => n11333, ZN => n11334);
   U15853 : XNOR2_X2 port map( A => n11335, B => n11334, ZN => n13211);
   U15854 : XNOR2_X1 port map( A => n11892, B => n12391, ZN => n11789);
   U15855 : XNOR2_X1 port map( A => n11336, B => n11424, ZN => n11337);
   U15856 : XNOR2_X1 port map( A => n11337, B => n11789, ZN => n11345);
   U15857 : MUX2_X1 port map( A => n11340, B => n11339, S => n11338, Z => 
                           n11939);
   U15858 : INV_X1 port map( A => n11935, ZN => n11341);
   U15859 : AOI21_X1 port map( B1 => n11939, B2 => n11342, A => n11341, ZN => 
                           n12263);
   U15860 : INV_X1 port map( A => n12263, ZN => n12161);
   U15861 : XNOR2_X1 port map( A => n11343, B => n12161, ZN => n11344);
   U15862 : XNOR2_X1 port map( A => n11345, B => n11344, ZN => n11350);
   U15863 : XNOR2_X1 port map( A => n12065, B => n11396, ZN => n11347);
   U15864 : XNOR2_X1 port map( A => n12277, B => n21944, ZN => n11346);
   U15865 : XNOR2_X1 port map( A => n12276, B => n12396, ZN => n12136);
   U15866 : INV_X1 port map( A => n12136, ZN => n11348);
   U15867 : XNOR2_X1 port map( A => n11349, B => n25047, ZN => n11684);
   U15868 : AOI21_X1 port map( B1 => n13211, B2 => n13206, A => n11684, ZN => 
                           n11367);
   U15869 : INV_X1 port map( A => n11350, ZN => n13004);
   U15870 : XNOR2_X1 port map( A => n12282, B => n11385, ZN => n11351);
   U15871 : XNOR2_X1 port map( A => n11351, B => n11991, ZN => n11354);
   U15872 : XNOR2_X1 port map( A => n12212, B => n1920, ZN => n11352);
   U15873 : INV_X1 port map( A => n12150, ZN => n12408);
   U15874 : XNOR2_X1 port map( A => n12408, B => n12286, ZN => n11781);
   U15875 : XNOR2_X1 port map( A => n11352, B => n11781, ZN => n11353);
   U15876 : XNOR2_X1 port map( A => n11353, B => n11354, ZN => n13000);
   U15877 : NAND2_X1 port map( A1 => n13004, A2 => n13000, ZN => n11361);
   U15878 : INV_X1 port map( A => n11355, ZN => n12247);
   U15879 : XNOR2_X1 port map( A => n12247, B => n11356, ZN => n11359);
   U15880 : XNOR2_X1 port map( A => n12234, B => n2033, ZN => n11357);
   U15881 : XNOR2_X1 port map( A => n11986, B => n11357, ZN => n11358);
   U15882 : NAND2_X1 port map( A1 => n11361, A2 => n11360, ZN => n12892);
   U15883 : XNOR2_X1 port map( A => n11581, B => n12241, ZN => n12124);
   U15884 : XNOR2_X1 port map( A => n12197, B => n888, ZN => n11362);
   U15885 : XNOR2_X1 port map( A => n12124, B => n11362, ZN => n11365);
   U15886 : XNOR2_X1 port map( A => n11761, B => n12378, ZN => n11800);
   U15887 : XNOR2_X1 port map( A => n12375, B => n25016, ZN => n11363);
   U15888 : XNOR2_X1 port map( A => n11800, B => n11363, ZN => n11364);
   U15889 : OAI21_X1 port map( B1 => n13213, B2 => n13206, A => n13000, ZN => 
                           n11366);
   U15890 : INV_X1 port map( A => n11411, ZN => n14290);
   U15891 : AOI21_X1 port map( B1 => n13951, B2 => n14294, A => n14290, ZN => 
                           n11368);
   U15892 : NAND2_X1 port map( A1 => n11369, A2 => n11368, ZN => n14686);
   U15893 : XNOR2_X1 port map( A => n11628, B => n12129, ZN => n11375);
   U15894 : AND3_X1 port map( A1 => n24913, A2 => n11371, A3 => n2211, ZN => 
                           n11373);
   U15895 : AOI21_X1 port map( B1 => n11371, B2 => n24913, A => n2211, ZN => 
                           n11372);
   U15896 : NOR2_X1 port map( A1 => n11373, A2 => n11372, ZN => n11374);
   U15897 : XNOR2_X1 port map( A => n11375, B => n11374, ZN => n11379);
   U15898 : XNOR2_X1 port map( A => n11638, B => n12306, ZN => n11377);
   U15899 : XNOR2_X1 port map( A => n11440, B => n11967, ZN => n11376);
   U15900 : XNOR2_X1 port map( A => n11376, B => n11377, ZN => n11378);
   U15901 : XNOR2_X1 port map( A => n11414, B => n12364, ZN => n11380);
   U15902 : XNOR2_X1 port map( A => n11946, B => n11380, ZN => n11383);
   U15903 : XNOR2_X1 port map( A => n11735, B => n860, ZN => n11381);
   U15904 : XNOR2_X1 port map( A => n12370, B => n12297, ZN => n11610);
   U15905 : XNOR2_X1 port map( A => n11610, B => n11381, ZN => n11382);
   U15906 : INV_X1 port map( A => n13027, ZN => n13030);
   U15907 : XNOR2_X1 port map( A => n12414, B => n853, ZN => n11384);
   U15908 : XNOR2_X1 port map( A => n11384, B => n12152, ZN => n11387);
   U15909 : XNOR2_X1 port map( A => n11385, B => n12324, ZN => n11386);
   U15910 : XNOR2_X1 port map( A => n11387, B => n11386, ZN => n11389);
   U15911 : XNOR2_X1 port map( A => n11388, B => n12409, ZN => n11956);
   U15913 : XNOR2_X1 port map( A => n11717, B => n12315, ZN => n11941);
   U15914 : XNOR2_X1 port map( A => n11941, B => n11614, ZN => n11393);
   U15915 : XNOR2_X1 port map( A => n11661, B => n20046, ZN => n11390);
   U15916 : XNOR2_X1 port map( A => n11391, B => n11390, ZN => n11392);
   U15917 : XNOR2_X1 port map( A => n11393, B => n11392, ZN => n13023);
   U15918 : INV_X1 port map( A => n12494, ZN => n11410);
   U15919 : XNOR2_X1 port map( A => n12334, B => n12067, ZN => n11394);
   U15920 : XNOR2_X1 port map( A => n11394, B => n24970, ZN => n11955);
   U15921 : XNOR2_X1 port map( A => n11795, B => n16574, ZN => n11395);
   U15922 : XNOR2_X1 port map( A => n12404, B => n11395, ZN => n11398);
   U15923 : XNOR2_X1 port map( A => n11396, B => n11622, ZN => n11397);
   U15924 : XNOR2_X1 port map( A => n11398, B => n11397, ZN => n11399);
   U15925 : XNOR2_X1 port map( A => n12343, B => n12375, ZN => n11604);
   U15926 : INV_X1 port map( A => n11401, ZN => n12382);
   U15927 : XNOR2_X1 port map( A => n12382, B => n25016, ZN => n11402);
   U15928 : XNOR2_X1 port map( A => n11402, B => n11604, ZN => n11405);
   U15929 : XNOR2_X1 port map( A => n12344, B => n12121, ZN => n11931);
   U15930 : XNOR2_X1 port map( A => n11765, B => n1757, ZN => n11403);
   U15931 : XNOR2_X1 port map( A => n11931, B => n11403, ZN => n11404);
   U15932 : INV_X1 port map( A => n13028, ZN => n13024);
   U15933 : INV_X1 port map( A => n13023, ZN => n12758);
   U15934 : OAI21_X1 port map( B1 => n13029, B2 => n13027, A => n11406, ZN => 
                           n11409);
   U15935 : NOR2_X1 port map( A1 => n12784, A2 => n13030, ZN => n11408);
   U15936 : INV_X1 port map( A => n11406, ZN => n11407);
   U15938 : NOR2_X1 port map( A1 => n13907, A2 => n11411, ZN => n11453);
   U15939 : XNOR2_X1 port map( A => n12168, B => n12089, ZN => n11985);
   U15940 : XNOR2_X1 port map( A => n11985, B => n11413, ZN => n11418);
   U15941 : XNOR2_X1 port map( A => n11414, B => n12362, ZN => n11416);
   U15942 : XNOR2_X1 port map( A => n25371, B => n2044, ZN => n11415);
   U15943 : XNOR2_X1 port map( A => n11416, B => n11415, ZN => n11417);
   U15945 : XNOR2_X1 port map( A => n11951, B => n12108, ZN => n11419);
   U15946 : XNOR2_X1 port map( A => n11419, B => n11420, ZN => n11423);
   U15947 : XNOR2_X1 port map( A => n11689, B => n2049, ZN => n11421);
   U15948 : XNOR2_X1 port map( A => n11975, B => n11421, ZN => n11422);
   U15949 : XNOR2_X1 port map( A => n11423, B => n11422, ZN => n13056);
   U15951 : XNOR2_X1 port map( A => n11425, B => n11942, ZN => n11427);
   U15952 : XNOR2_X1 port map( A => n11427, B => n11426, ZN => n11430);
   U15953 : INV_X1 port map( A => n12082, ZN => n11428);
   U15954 : XNOR2_X1 port map( A => n11429, B => n11428, ZN => n12013);
   U15955 : INV_X1 port map( A => n13057, ZN => n13054);
   U15956 : XNOR2_X1 port map( A => n12383, B => n21046, ZN => n11431);
   U15957 : XNOR2_X1 port map( A => n11432, B => n11431, ZN => n11437);
   U15958 : XNOR2_X1 port map( A => n11433, B => n11706, ZN => n11434);
   U15959 : XNOR2_X1 port map( A => n11435, B => n11434, ZN => n11436);
   U15960 : XNOR2_X1 port map( A => n12005, B => n11439, ZN => n11444);
   U15961 : XNOR2_X1 port map( A => n11457, B => n11440, ZN => n11442);
   U15962 : INV_X1 port map( A => n12002, ZN => n12075);
   U15963 : XNOR2_X1 port map( A => n12075, B => n2208, ZN => n11441);
   U15964 : XNOR2_X1 port map( A => n11442, B => n11441, ZN => n11443);
   U15965 : NOR2_X1 port map( A1 => n303, A2 => n13056, ZN => n12751);
   U15966 : XNOR2_X1 port map( A => n12147, B => n11960, ZN => n11445);
   U15967 : XNOR2_X1 port map( A => n11446, B => n11445, ZN => n11450);
   U15968 : XNOR2_X1 port map( A => n11741, B => n12102, ZN => n11448);
   U15969 : XNOR2_X1 port map( A => n11448, B => n11447, ZN => n11449);
   U15970 : XNOR2_X1 port map( A => n11450, B => n11449, ZN => n13052);
   U15971 : INV_X1 port map( A => n13052, ZN => n13055);
   U15972 : AND2_X1 port map( A1 => n13053, A2 => n13055, ZN => n12485);
   U15973 : AOI21_X1 port map( B1 => n12751, B2 => n25085, A => n12485, ZN => 
                           n11451);
   U15974 : NAND2_X1 port map( A1 => n11452, A2 => n11451, ZN => n14289);
   U15975 : INV_X1 port map( A => n12184, ZN => n11455);
   U15976 : XNOR2_X1 port map( A => n11455, B => n12129, ZN => n11701);
   U15977 : XNOR2_X1 port map( A => n11701, B => n11456, ZN => n11461);
   U15978 : XNOR2_X1 port map( A => n11457, B => n11637, ZN => n11459);
   U15979 : XNOR2_X1 port map( A => n12356, B => n912, ZN => n11458);
   U15980 : XNOR2_X1 port map( A => n11459, B => n11458, ZN => n11460);
   U15981 : XNOR2_X1 port map( A => n11461, B => n11460, ZN => n12462);
   U15982 : INV_X1 port map( A => n12462, ZN => n12713);
   U15985 : XNOR2_X1 port map( A => n11812, B => n11463, ZN => n11468);
   U15986 : XNOR2_X1 port map( A => n11464, B => n12201, ZN => n11466);
   U15987 : XNOR2_X1 port map( A => n24964, B => n641, ZN => n11465);
   U15988 : XNOR2_X1 port map( A => n11466, B => n11465, ZN => n11467);
   U15989 : XNOR2_X2 port map( A => n11468, B => n11467, ZN => n12483);
   U15990 : NOR2_X1 port map( A1 => n12713, A2 => n12483, ZN => n12464);
   U15991 : XNOR2_X1 port map( A => n11469, B => n11816, ZN => n11473);
   U15992 : XNOR2_X1 port map( A => n12404, B => n12189, ZN => n11471);
   U15993 : XNOR2_X1 port map( A => n11951, B => n3178, ZN => n11470);
   U15994 : XNOR2_X1 port map( A => n11471, B => n11470, ZN => n11472);
   U15995 : XNOR2_X1 port map( A => n11473, B => n11472, ZN => n12715);
   U15996 : INV_X1 port map( A => n12715, ZN => n13078);
   U15997 : NOR2_X1 port map( A1 => n12462, A2 => n13078, ZN => n11474);
   U15998 : NOR2_X1 port map( A1 => n12464, A2 => n11474, ZN => n11589);
   U15999 : INV_X1 port map( A => n11960, ZN => n11475);
   U16000 : XNOR2_X1 port map( A => n12144, B => n11475, ZN => n11476);
   U16001 : XNOR2_X1 port map( A => n11822, B => n11476, ZN => n11480);
   U16002 : XNOR2_X1 port map( A => n12414, B => n12207, ZN => n11478);
   U16003 : XNOR2_X1 port map( A => n25087, B => n24287, ZN => n11477);
   U16004 : XNOR2_X1 port map( A => n11478, B => n11477, ZN => n11479);
   U16006 : XNOR2_X1 port map( A => n11717, B => n11660, ZN => n11482);
   U16007 : XNOR2_X1 port map( A => n11482, B => n11481, ZN => n11485);
   U16008 : XNOR2_X1 port map( A => n11827, B => n11483, ZN => n11484);
   U16009 : XNOR2_X1 port map( A => n11485, B => n11484, ZN => n12707);
   U16010 : MUX2_X1 port map( A => n12710, B => n12707, S => n12483, Z => 
                           n11592);
   U16011 : XNOR2_X1 port map( A => n25090, B => n11486, ZN => n11488);
   U16012 : XNOR2_X1 port map( A => n12370, B => n3129, ZN => n11487);
   U16013 : XNOR2_X1 port map( A => n11488, B => n11487, ZN => n11491);
   U16014 : XNOR2_X1 port map( A => n11489, B => n11833, ZN => n11490);
   U16016 : MUX2_X2 port map( A => n11589, B => n11592, S => n24573, Z => 
                           n14362);
   U16017 : INV_X1 port map( A => n11492, ZN => n11770);
   U16018 : XNOR2_X1 port map( A => n11770, B => n12186, ZN => n11493);
   U16019 : XNOR2_X1 port map( A => n11494, B => n11493, ZN => n11497);
   U16020 : XNOR2_X1 port map( A => n11627, B => n836, ZN => n11495);
   U16021 : XNOR2_X1 port map( A => n11856, B => n11495, ZN => n11496);
   U16022 : MUX2_X1 port map( A => n11500, B => n11499, S => n11498, Z => 
                           n11503);
   U16023 : INV_X1 port map( A => n11501, ZN => n11502);
   U16024 : NOR2_X1 port map( A1 => n11503, A2 => n11502, ZN => n11577);
   U16025 : XNOR2_X1 port map( A => n11619, B => n11577, ZN => n11505);
   U16026 : XNOR2_X1 port map( A => n12333, B => n2735, ZN => n11506);
   U16027 : XNOR2_X1 port map( A => n11868, B => n11506, ZN => n11507);
   U16028 : XNOR2_X1 port map( A => n11508, B => n11507, ZN => n12469);
   U16029 : NOR2_X1 port map( A1 => n13067, A2 => n12469, ZN => n11541);
   U16030 : XNOR2_X1 port map( A => n11915, B => n11766, ZN => n11509);
   U16031 : XNOR2_X1 port map( A => n11510, B => n11509, ZN => n11514);
   U16032 : XNOR2_X1 port map( A => n12200, B => n1827, ZN => n11511);
   U16033 : XNOR2_X1 port map( A => n11511, B => n11512, ZN => n11513);
   U16034 : INV_X1 port map( A => n11515, ZN => n11517);
   U16035 : XNOR2_X1 port map( A => n24401, B => n12040, ZN => n11531);
   U16036 : NAND2_X1 port map( A1 => n11520, A2 => n11524, ZN => n11528);
   U16037 : INV_X1 port map( A => n11518, ZN => n11521);
   U16038 : NAND3_X1 port map( A1 => n11521, A2 => n11520, A3 => n11519, ZN => 
                           n11523);
   U16039 : AND2_X1 port map( A1 => n11522, A2 => n11523, ZN => n11527);
   U16040 : NAND3_X1 port map( A1 => n11525, A2 => n1332, A3 => n11524, ZN => 
                           n11526);
   U16042 : XNOR2_X1 port map( A => n12323, B => n3115, ZN => n11530);
   U16043 : XNOR2_X1 port map( A => n11531, B => n11530, ZN => n11532);
   U16044 : INV_X1 port map( A => n12471, ZN => n13072);
   U16045 : XNOR2_X1 port map( A => n12234, B => n1724, ZN => n11534);
   U16046 : XNOR2_X1 port map( A => n11535, B => n11534, ZN => n11540);
   U16047 : INV_X1 port map( A => n11536, ZN => n11538);
   U16048 : XNOR2_X1 port map( A => n11538, B => n11537, ZN => n11539);
   U16049 : XNOR2_X1 port map( A => n11542, B => n12313, ZN => n11544);
   U16050 : XNOR2_X1 port map( A => n11544, B => n11543, ZN => n11547);
   U16051 : XNOR2_X1 port map( A => n11863, B => n11545, ZN => n11546);
   U16052 : INV_X1 port map( A => n12773, ZN => n13071);
   U16053 : NOR2_X1 port map( A1 => n13071, A2 => n12471, ZN => n11548);
   U16054 : NOR3_X1 port map( A1 => n11549, A2 => n13070, A3 => n11548, ZN => 
                           n11550);
   U16055 : NOR2_X2 port map( A1 => n11551, A2 => n11550, ZN => n14361);
   U16056 : NAND2_X1 port map( A1 => n14362, A2 => n14361, ZN => n13711);
   U16057 : XNOR2_X1 port map( A => n11715, B => n11659, ZN => n12259);
   U16058 : XNOR2_X1 port map( A => n11789, B => n12259, ZN => n11554);
   U16059 : XNOR2_X1 port map( A => n12225, B => n2215, ZN => n11552);
   U16060 : XNOR2_X1 port map( A => n12011, B => n11552, ZN => n11553);
   U16061 : XNOR2_X1 port map( A => n11554, B => n11553, ZN => n13038);
   U16062 : INV_X1 port map( A => n13038, ZN => n12476);
   U16063 : XNOR2_X1 port map( A => n11555, B => n12214, ZN => n11557);
   U16064 : XNOR2_X1 port map( A => n24027, B => n11653, ZN => n12284);
   U16065 : XNOR2_X1 port map( A => n11557, B => n12284, ZN => n11560);
   U16066 : XNOR2_X1 port map( A => n12040, B => n869, ZN => n11558);
   U16067 : XNOR2_X1 port map( A => n11781, B => n11558, ZN => n11559);
   U16068 : XNOR2_X1 port map( A => n11560, B => n11559, ZN => n13037);
   U16069 : INV_X1 port map( A => n13037, ZN => n12798);
   U16072 : XNOR2_X1 port map( A => n11563, B => n12365, ZN => n12166);
   U16073 : XNOR2_X1 port map( A => n12246, B => n12166, ZN => n11567);
   U16074 : XNOR2_X1 port map( A => n11564, B => n11983, ZN => n12230);
   U16075 : XNOR2_X1 port map( A => n11908, B => n887, ZN => n11565);
   U16076 : XNOR2_X1 port map( A => n12230, B => n11565, ZN => n11566);
   U16077 : XNOR2_X1 port map( A => n11879, B => n12186, ZN => n11569);
   U16078 : XNOR2_X1 port map( A => n11568, B => n11640, ZN => n12268);
   U16079 : XNOR2_X1 port map( A => n11569, B => n12268, ZN => n11573);
   U16080 : XNOR2_X1 port map( A => n11570, B => n11571, ZN => n11572);
   U16081 : XNOR2_X1 port map( A => n12277, B => n12396, ZN => n11792);
   U16082 : XNOR2_X1 port map( A => n11792, B => n25236, ZN => n11575);
   U16083 : XNOR2_X1 port map( A => n11672, B => n11689, ZN => n12273);
   U16084 : XNOR2_X1 port map( A => n11575, B => n12273, ZN => n11579);
   U16085 : XNOR2_X1 port map( A => n11977, B => n3152, ZN => n11576);
   U16086 : XNOR2_X1 port map( A => n11577, B => n11576, ZN => n11578);
   U16087 : XNOR2_X1 port map( A => n11579, B => n11578, ZN => n12800);
   U16088 : XNOR2_X1 port map( A => n12239, B => n11800, ZN => n11586);
   U16089 : XNOR2_X1 port map( A => n11581, B => n11582, ZN => n11584);
   U16090 : XNOR2_X1 port map( A => n12196, B => n1874, ZN => n11583);
   U16091 : XNOR2_X1 port map( A => n11584, B => n11583, ZN => n11585);
   U16092 : XNOR2_X1 port map( A => n11586, B => n11585, ZN => n12519);
   U16093 : INV_X1 port map( A => n12519, ZN => n13039);
   U16094 : NOR2_X1 port map( A1 => n13039, A2 => n13038, ZN => n11588);
   U16095 : INV_X1 port map( A => n13041, ZN => n11587);
   U16096 : OAI21_X1 port map( B1 => n11588, B2 => n13044, A => n11587, ZN => 
                           n11590);
   U16097 : INV_X1 port map( A => n11590, ZN => n11591);
   U16098 : AOI21_X1 port map( B1 => n11592, B2 => n24573, A => n11591, ZN => 
                           n11593);
   U16099 : NAND2_X1 port map( A1 => n11594, A2 => n11593, ZN => n11601);
   U16100 : INV_X1 port map( A => n11595, ZN => n11600);
   U16101 : INV_X1 port map( A => n13169, ZN => n12718);
   U16102 : OAI22_X1 port map( A1 => n12716, A2 => n11597, B1 => n12719, B2 => 
                           n10502, ZN => n11598);
   U16103 : XNOR2_X1 port map( A => n11914, B => n1810, ZN => n11603);
   U16104 : XNOR2_X1 port map( A => n11602, B => n11603, ZN => n11606);
   U16105 : XNOR2_X1 port map( A => n11704, B => n11766, ZN => n12342);
   U16106 : XNOR2_X1 port map( A => n12342, B => n11604, ZN => n11605);
   U16107 : XNOR2_X1 port map( A => n11736, B => n11607, ZN => n12292);
   U16108 : XNOR2_X1 port map( A => n11608, B => n12292, ZN => n11612);
   U16109 : XNOR2_X1 port map( A => n12249, B => n22986, ZN => n11609);
   U16110 : XNOR2_X1 port map( A => n11610, B => n11609, ZN => n11611);
   U16112 : XNOR2_X1 port map( A => n12388, B => n2318, ZN => n11613);
   U16113 : XNOR2_X1 port map( A => n11613, B => n12255, ZN => n11615);
   U16114 : XNOR2_X1 port map( A => n11749, B => n11616, ZN => n12312);
   U16115 : XNOR2_X1 port map( A => n12312, B => n24915, ZN => n11617);
   U16116 : XNOR2_X1 port map( A => n11618, B => n11619, ZN => n12339);
   U16117 : XNOR2_X1 port map( A => n12112, B => n3131, ZN => n11620);
   U16118 : XNOR2_X1 port map( A => n11620, B => n12397, ZN => n11621);
   U16119 : XNOR2_X1 port map( A => n11621, B => n12339, ZN => n11625);
   U16120 : XNOR2_X1 port map( A => n11622, B => n12275, ZN => n11623);
   U16121 : XNOR2_X1 port map( A => n12404, B => n11623, ZN => n11624);
   U16122 : XNOR2_X1 port map( A => n11699, B => n11626, ZN => n11631);
   U16123 : XNOR2_X1 port map( A => n11698, B => n11627, ZN => n12307);
   U16124 : XNOR2_X1 port map( A => n11628, B => n11809, ZN => n11629);
   U16125 : XNOR2_X1 port map( A => n12307, B => n11629, ZN => n11630);
   U16127 : XNOR2_X1 port map( A => n12283, B => n12324, ZN => n11632);
   U16128 : XNOR2_X1 port map( A => n11632, B => n12320, ZN => n11636);
   U16129 : XNOR2_X1 port map( A => n11897, B => n12413, ZN => n11634);
   U16130 : XNOR2_X1 port map( A => n12414, B => n92, ZN => n11633);
   U16131 : XNOR2_X1 port map( A => n11634, B => n11633, ZN => n11635);
   U16132 : XNOR2_X1 port map( A => n12132, B => n11639, ZN => n11644);
   U16133 : XNOR2_X1 port map( A => n11640, B => n1924, ZN => n11641);
   U16134 : XNOR2_X1 port map( A => n11642, B => n11641, ZN => n11643);
   U16135 : XNOR2_X1 port map( A => n25090, B => n11735, ZN => n12165);
   U16136 : XNOR2_X1 port map( A => n11734, B => n12165, ZN => n11650);
   U16137 : XNOR2_X1 port map( A => n11646, B => n2477, ZN => n11647);
   U16138 : XNOR2_X1 port map( A => n11648, B => n11647, ZN => n11649);
   U16139 : INV_X1 port map( A => Key(172), ZN => n23271);
   U16140 : XNOR2_X1 port map( A => n12325, B => n23271, ZN => n11651);
   U16141 : XNOR2_X1 port map( A => n11651, B => n12146, ZN => n11652);
   U16142 : XNOR2_X1 port map( A => n12409, B => n12102, ZN => n11743);
   U16143 : XNOR2_X1 port map( A => n11652, B => n11743, ZN => n11656);
   U16144 : XNOR2_X1 port map( A => n25087, B => n11653, ZN => n11654);
   U16145 : XNOR2_X1 port map( A => n12152, B => n11654, ZN => n11655);
   U16148 : XNOR2_X1 port map( A => n12053, B => n2747, ZN => n11657);
   U16149 : XNOR2_X1 port map( A => n11658, B => n11657, ZN => n11664);
   U16150 : XNOR2_X1 port map( A => n11659, B => n12082, ZN => n11662);
   U16151 : XNOR2_X1 port map( A => n11661, B => n11660, ZN => n12157);
   U16152 : XNOR2_X1 port map( A => n12157, B => n11662, ZN => n11663);
   U16153 : XNOR2_X1 port map( A => n11666, B => n11665, ZN => n11669);
   U16154 : XNOR2_X1 port map( A => n11765, B => n11464, ZN => n11798);
   U16155 : XNOR2_X1 port map( A => n11838, B => n1815, ZN => n11667);
   U16156 : XNOR2_X1 port map( A => n11798, B => n11667, ZN => n11668);
   U16157 : XNOR2_X1 port map( A => n11668, B => n11669, ZN => n12454);
   U16158 : NOR2_X1 port map( A1 => n13063, A2 => n13061, ZN => n11678);
   U16159 : XNOR2_X1 port map( A => n11795, B => n1854, ZN => n11670);
   U16160 : XNOR2_X1 port map( A => n11670, B => n12334, ZN => n11671);
   U16161 : XNOR2_X1 port map( A => n12108, B => n12402, ZN => n11758);
   U16162 : XNOR2_X1 port map( A => n11671, B => n11758, ZN => n11676);
   U16163 : INV_X1 port map( A => n11672, ZN => n11673);
   U16164 : XNOR2_X1 port map( A => n11673, B => n25236, ZN => n11674);
   U16165 : XNOR2_X1 port map( A => n11796, B => n11674, ZN => n11675);
   U16166 : XNOR2_X1 port map( A => n11676, B => n11675, ZN => n12439);
   U16167 : INV_X1 port map( A => n12439, ZN => n13163);
   U16168 : NAND2_X1 port map( A1 => n13163, A2 => n1353, ZN => n11677);
   U16169 : NAND2_X1 port map( A1 => n13394, A2 => n13568, ZN => n11679);
   U16170 : OR2_X1 port map( A1 => n13712, A2 => n11679, ZN => n11680);
   U16171 : XNOR2_X1 port map( A => n11682, B => n15401, ZN => n14884);
   U16172 : NAND2_X1 port map( A1 => n13211, A2 => n11684, ZN => n12551);
   U16173 : NAND3_X1 port map( A1 => n13213, A2 => n11684, A3 => n13004, ZN => 
                           n11683);
   U16174 : OAI21_X1 port map( B1 => n12551, B2 => n11360, A => n11683, ZN => 
                           n11685);
   U16175 : INV_X1 port map( A => n13000, ZN => n13212);
   U16176 : XNOR2_X1 port map( A => n11686, B => n23699, ZN => n11687);
   U16177 : XNOR2_X1 port map( A => n11687, B => n24969, ZN => n11688);
   U16178 : XNOR2_X1 port map( A => n12064, B => n11688, ZN => n11691);
   U16179 : XNOR2_X1 port map( A => n11689, B => n11690, ZN => n11926);
   U16180 : XNOR2_X1 port map( A => n11691, B => n11926, ZN => n12613);
   U16181 : INV_X1 port map( A => n11692, ZN => n11906);
   U16182 : XNOR2_X1 port map( A => n11906, B => n12030, ZN => n11697);
   U16183 : INV_X1 port map( A => n11693, ZN => n11695);
   U16184 : XNOR2_X1 port map( A => n12167, B => n21742, ZN => n11694);
   U16185 : XNOR2_X1 port map( A => n11695, B => n11694, ZN => n11696);
   U16187 : NAND2_X1 port map( A1 => n12613, A2 => n13305, ZN => n12558);
   U16188 : XNOR2_X1 port map( A => n11698, B => n5286, ZN => n11700);
   U16189 : INV_X1 port map( A => n11701, ZN => n11702);
   U16190 : XNOR2_X1 port map( A => n11703, B => n12201, ZN => n12045);
   U16191 : XNOR2_X1 port map( A => n11704, B => n925, ZN => n11705);
   U16192 : XNOR2_X1 port map( A => n12096, B => n12200, ZN => n11707);
   U16193 : XNOR2_X1 port map( A => n11706, B => n11707, ZN => n11918);
   U16194 : XNOR2_X1 port map( A => n11708, B => n11918, ZN => n12611);
   U16196 : XNOR2_X1 port map( A => n11959, B => n2744, ZN => n11709);
   U16197 : XNOR2_X1 port map( A => n25418, B => n11709, ZN => n11713);
   U16198 : XNOR2_X1 port map( A => n11897, B => n12144, ZN => n11711);
   U16199 : XNOR2_X1 port map( A => n11711, B => n11900, ZN => n11712);
   U16200 : OAI21_X1 port map( B1 => n12558, B2 => n12915, A => n11714, ZN => 
                           n11723);
   U16201 : XNOR2_X1 port map( A => n11715, B => n12224, ZN => n11890);
   U16202 : XNOR2_X1 port map( A => n11716, B => n11890, ZN => n11721);
   U16203 : XNOR2_X1 port map( A => n11717, B => n1856, ZN => n11719);
   U16204 : INV_X1 port map( A => n11718, ZN => n12058);
   U16205 : XNOR2_X1 port map( A => n11719, B => n12058, ZN => n11720);
   U16206 : INV_X1 port map( A => n11724, ZN => n11726);
   U16207 : XNOR2_X1 port map( A => n11725, B => n11726, ZN => n11731);
   U16208 : XNOR2_X1 port map( A => n11771, B => n11966, ZN => n11729);
   U16209 : INV_X1 port map( A => n12351, ZN => n11727);
   U16210 : XNOR2_X1 port map( A => n11727, B => n768, ZN => n11728);
   U16211 : XNOR2_X1 port map( A => n11729, B => n11728, ZN => n11730);
   U16213 : XNOR2_X1 port map( A => n12362, B => n24514, ZN => n11733);
   U16214 : XNOR2_X1 port map( A => n11734, B => n11733, ZN => n11740);
   U16215 : INV_X1 port map( A => n21169, ZN => n22556);
   U16216 : XNOR2_X1 port map( A => n11735, B => n22556, ZN => n11738);
   U16217 : XNOR2_X1 port map( A => n11736, B => n25371, ZN => n11737);
   U16218 : XNOR2_X1 port map( A => n11738, B => n11737, ZN => n11739);
   U16219 : XNOR2_X1 port map( A => n11741, B => n11960, ZN => n12416);
   U16220 : XNOR2_X1 port map( A => n12286, B => n2040, ZN => n11742);
   U16221 : XNOR2_X1 port map( A => n12416, B => n11742, ZN => n11744);
   U16222 : INV_X1 port map( A => n13227, ZN => n11754);
   U16223 : XNOR2_X1 port map( A => n12053, B => n11746, ZN => n11748);
   U16224 : XNOR2_X1 port map( A => n11747, B => n11748, ZN => n12395);
   U16225 : XNOR2_X1 port map( A => n11749, B => n2847, ZN => n11750);
   U16226 : XNOR2_X1 port map( A => n12257, B => n12082, ZN => n11751);
   U16227 : XNOR2_X1 port map( A => n11752, B => n11751, ZN => n11753);
   U16228 : NOR2_X1 port map( A1 => n13221, A2 => n11755, ZN => n12920);
   U16229 : XNOR2_X1 port map( A => n11756, B => n11951, ZN => n12400);
   U16230 : XNOR2_X1 port map( A => n12277, B => n23620, ZN => n11757);
   U16231 : XNOR2_X1 port map( A => n11759, B => n11758, ZN => n11760);
   U16232 : XNOR2_X1 port map( A => n11761, B => n923, ZN => n11762);
   U16233 : XNOR2_X1 port map( A => n12376, B => n11762, ZN => n11763);
   U16234 : XNOR2_X1 port map( A => n11765, B => n24964, ZN => n11767);
   U16235 : XNOR2_X1 port map( A => n11767, B => n11766, ZN => n11768);
   U16236 : INV_X1 port map( A => n12569, ZN => n12924);
   U16237 : OAI211_X1 port map( C1 => n13223, C2 => n12885, A => n12924, B => 
                           n13224, ZN => n11769);
   U16238 : OAI21_X1 port map( B1 => n13010, B2 => n12920, A => n11769, ZN => 
                           n13965);
   U16239 : XNOR2_X1 port map( A => n12132, B => n12074, ZN => n11775);
   U16240 : XNOR2_X1 port map( A => n11771, B => n11770, ZN => n11773);
   U16241 : XNOR2_X1 port map( A => n12355, B => n1758, ZN => n11772);
   U16242 : XNOR2_X1 port map( A => n11773, B => n11772, ZN => n11774);
   U16243 : XNOR2_X1 port map( A => n12165, B => n12088, ZN => n11780);
   U16244 : XNOR2_X1 port map( A => n12296, B => n12365, ZN => n11778);
   U16245 : XNOR2_X1 port map( A => n11908, B => n763, ZN => n11777);
   U16246 : XNOR2_X1 port map( A => n11778, B => n11777, ZN => n11779);
   U16247 : INV_X1 port map( A => n12594, ZN => n12597);
   U16248 : XNOR2_X1 port map( A => n24980, B => n12323, ZN => n11784);
   U16249 : XNOR2_X1 port map( A => n25087, B => n62, ZN => n11783);
   U16250 : XNOR2_X1 port map( A => n11784, B => n11783, ZN => n11785);
   U16252 : XNOR2_X1 port map( A => n12157, B => n11787, ZN => n11791);
   U16253 : XNOR2_X1 port map( A => n12313, B => n2190, ZN => n11788);
   U16254 : XNOR2_X1 port map( A => n11789, B => n11788, ZN => n11790);
   U16255 : XNOR2_X1 port map( A => n11790, B => n11791, ZN => n13288);
   U16257 : XNOR2_X1 port map( A => n12333, B => n1777, ZN => n11793);
   U16258 : XNOR2_X1 port map( A => n11792, B => n11793, ZN => n11794);
   U16260 : XNOR2_X1 port map( A => n11796, B => n11795, ZN => n12141);
   U16261 : XNOR2_X1 port map( A => n12095, B => n11800, ZN => n11801);
   U16262 : XNOR2_X1 port map( A => n11802, B => n11801, ZN => n12593);
   U16263 : BUF_X2 port map( A => n12593, Z => n12827);
   U16264 : NOR2_X1 port map( A1 => n11804, A2 => n11803, ZN => n11805);
   U16265 : INV_X1 port map( A => n11805, ZN => n13884);
   U16267 : XNOR2_X1 port map( A => n12019, B => n12002, ZN => n11808);
   U16268 : XNOR2_X1 port map( A => n12357, B => n1855, ZN => n11807);
   U16269 : XNOR2_X1 port map( A => n11808, B => n11807, ZN => n11811);
   U16270 : XNOR2_X1 port map( A => n12186, B => n11809, ZN => n12025);
   U16271 : XNOR2_X1 port map( A => n12306, B => n12129, ZN => n11970);
   U16272 : XNOR2_X1 port map( A => n12025, B => n11970, ZN => n11810);
   U16273 : XNOR2_X1 port map( A => n11812, B => n12046, ZN => n11815);
   U16274 : XNOR2_X1 port map( A => n11931, B => n11813, ZN => n11814);
   U16276 : XNOR2_X1 port map( A => n12334, B => n12138, ZN => n11817);
   U16277 : XNOR2_X1 port map( A => n11816, B => n11817, ZN => n11820);
   U16278 : XNOR2_X1 port map( A => n12108, B => n23679, ZN => n11818);
   U16279 : XNOR2_X1 port map( A => n12063, B => n11818, ZN => n11819);
   U16280 : XNOR2_X1 port map( A => n12144, B => n12324, ZN => n11821);
   U16281 : XNOR2_X1 port map( A => n11822, B => n11821, ZN => n11826);
   U16282 : XNOR2_X1 port map( A => n12040, B => n12102, ZN => n11824);
   U16283 : XNOR2_X1 port map( A => n12325, B => n1746, ZN => n11823);
   U16284 : XNOR2_X1 port map( A => n11824, B => n11823, ZN => n11825);
   U16285 : XNOR2_X1 port map( A => n11826, B => n11825, ZN => n12935);
   U16287 : XNOR2_X1 port map( A => n12082, B => n20744, ZN => n11828);
   U16288 : XNOR2_X1 port map( A => n11827, B => n11828, ZN => n11831);
   U16289 : INV_X1 port map( A => n11829, ZN => n12057);
   U16290 : XNOR2_X1 port map( A => n11941, B => n12057, ZN => n11830);
   U16291 : INV_X1 port map( A => n13298, ZN => n12936);
   U16292 : XNOR2_X1 port map( A => n12089, B => n1875, ZN => n11832);
   U16293 : XNOR2_X1 port map( A => n11832, B => n11946, ZN => n11835);
   U16294 : XNOR2_X1 port map( A => n11833, B => n12028, ZN => n11834);
   U16295 : XNOR2_X1 port map( A => n12377, B => n25016, ZN => n11841);
   U16296 : XNOR2_X1 port map( A => n11842, B => n11841, ZN => n11843);
   U16298 : XNOR2_X1 port map( A => n12413, B => n11845, ZN => n11847);
   U16299 : XNOR2_X1 port map( A => n12323, B => n2970, ZN => n11846);
   U16300 : INV_X1 port map( A => n11848, ZN => n12105);
   U16301 : XNOR2_X1 port map( A => n11849, B => n12105, ZN => n11850);
   U16302 : XNOR2_X1 port map( A => n25234, B => n1870, ZN => n11853);
   U16303 : INV_X1 port map( A => n11851, ZN => n11852);
   U16304 : XNOR2_X1 port map( A => n11852, B => n11853, ZN => n11855);
   U16305 : XNOR2_X1 port map( A => n12087, B => n11905, ZN => n11854);
   U16308 : XNOR2_X1 port map( A => n12073, B => n11856, ZN => n11860);
   U16309 : XNOR2_X1 port map( A => n12020, B => n921, ZN => n11857);
   U16310 : XNOR2_X1 port map( A => n11858, B => n11857, ZN => n11859);
   U16311 : INV_X1 port map( A => n11861, ZN => n12080);
   U16312 : XNOR2_X1 port map( A => n12388, B => n2036, ZN => n11862);
   U16313 : XNOR2_X1 port map( A => n12080, B => n11862, ZN => n11865);
   U16314 : XNOR2_X1 port map( A => n11863, B => n11893, ZN => n11864);
   U16315 : XNOR2_X1 port map( A => n11865, B => n11864, ZN => n12900);
   U16316 : NAND2_X1 port map( A1 => n12899, A2 => n12900, ZN => n11866);
   U16317 : NAND3_X1 port map( A1 => n11867, A2 => n5672, A3 => n11866, ZN => 
                           n11875);
   U16318 : XNOR2_X1 port map( A => n11924, B => n12110, ZN => n11872);
   U16319 : XNOR2_X1 port map( A => n12397, B => n1864, ZN => n11870);
   U16320 : INV_X1 port map( A => n11868, ZN => n11869);
   U16321 : XNOR2_X1 port map( A => n11870, B => n11869, ZN => n11871);
   U16322 : NAND3_X1 port map( A1 => n12928, A2 => n12897, A3 => n11873, ZN => 
                           n11874);
   U16323 : XNOR2_X1 port map( A => n12183, B => n2717, ZN => n11877);
   U16324 : XNOR2_X1 port map( A => n11878, B => n11877, ZN => n11883);
   U16325 : XNOR2_X1 port map( A => n11879, B => n12019, ZN => n11881);
   U16326 : XNOR2_X1 port map( A => n11881, B => n11880, ZN => n11882);
   U16327 : NAND2_X1 port map( A1 => n714, A2 => n11884, ZN => n11887);
   U16328 : NAND2_X1 port map( A1 => n10690, A2 => n11147, ZN => n11886);
   U16329 : MUX2_X1 port map( A => n11887, B => n11886, S => n11885, Z => 
                           n11889);
   U16330 : NAND2_X1 port map( A1 => n11889, A2 => n11888, ZN => n12055);
   U16331 : XNOR2_X1 port map( A => n12055, B => n12226, ZN => n11891);
   U16332 : XNOR2_X1 port map( A => n11891, B => n11890, ZN => n11896);
   U16333 : XNOR2_X1 port map( A => n11892, B => n889, ZN => n11894);
   U16334 : XNOR2_X1 port map( A => n11894, B => n11893, ZN => n11895);
   U16335 : XNOR2_X1 port map( A => n11895, B => n11896, ZN => n12942);
   U16336 : INV_X1 port map( A => n12101, ZN => n11898);
   U16337 : XNOR2_X1 port map( A => n12283, B => n11898, ZN => n11899);
   U16338 : XNOR2_X1 port map( A => n11899, B => n11900, ZN => n11904);
   U16339 : XNOR2_X1 port map( A => n12039, B => n12286, ZN => n11902);
   U16340 : XNOR2_X1 port map( A => n12323, B => n4189, ZN => n11901);
   U16341 : XNOR2_X1 port map( A => n11902, B => n11901, ZN => n11903);
   U16342 : INV_X1 port map( A => n12031, ZN => n11909);
   U16343 : XNOR2_X1 port map( A => n11909, B => n22745, ZN => n11910);
   U16344 : XNOR2_X1 port map( A => n11911, B => n11910, ZN => n11912);
   U16345 : XNOR2_X2 port map( A => n5749, B => n11912, ZN => n13317);
   U16346 : NOR2_X1 port map( A1 => n12945, A2 => n13317, ZN => n11920);
   U16347 : XNOR2_X1 port map( A => n11916, B => n11915, ZN => n11917);
   U16348 : MUX2_X1 port map( A => n11921, B => n11920, S => n25499, Z => 
                           n11928);
   U16349 : XNOR2_X1 port map( A => n12277, B => n23883, ZN => n11923);
   U16350 : INV_X1 port map( A => n12066, ZN => n11922);
   U16352 : INV_X1 port map( A => n13318, ZN => n12580);
   U16353 : INV_X1 port map( A => n12942, ZN => n13316);
   U16354 : OAI22_X1 port map( A1 => n13321, A2 => n12580, B1 => n12687, B2 => 
                           n13316, ZN => n11927);
   U16355 : XNOR2_X1 port map( A => n12382, B => n12241, ZN => n11930);
   U16356 : XNOR2_X1 port map( A => n24964, B => n2826, ZN => n11929);
   U16357 : XNOR2_X1 port map( A => n11930, B => n11929, ZN => n11933);
   U16358 : XNOR2_X1 port map( A => n12342, B => n11931, ZN => n11932);
   U16359 : XNOR2_X1 port map( A => n11932, B => n11933, ZN => n12600);
   U16360 : NAND2_X1 port map( A1 => n11935, A2 => n4711, ZN => n11938);
   U16361 : NAND2_X1 port map( A1 => n11939, A2 => n11934, ZN => n11937);
   U16362 : MUX2_X1 port map( A => n4711, B => n1495, S => n11935, Z => n11936)
                           ;
   U16363 : OAI211_X1 port map( C1 => n11939, C2 => n11938, A => n11937, B => 
                           n11936, ZN => n11940);
   U16364 : XNOR2_X1 port map( A => n11941, B => n11940, ZN => n11945);
   U16365 : XNOR2_X1 port map( A => n12053, B => n11942, ZN => n11944);
   U16366 : INV_X1 port map( A => n12312, ZN => n11943);
   U16367 : NOR2_X1 port map( A1 => n12966, A2 => n12963, ZN => n11974);
   U16368 : XNOR2_X1 port map( A => n12292, B => n11946, ZN => n11950);
   U16369 : XNOR2_X1 port map( A => n12364, B => n25371, ZN => n11948);
   U16370 : XNOR2_X1 port map( A => n12168, B => n2039, ZN => n11947);
   U16371 : XNOR2_X1 port map( A => n11948, B => n11947, ZN => n11949);
   U16372 : XNOR2_X1 port map( A => n11950, B => n11949, ZN => n11965);
   U16373 : XNOR2_X1 port map( A => n12276, B => n2058, ZN => n11952);
   U16374 : XNOR2_X1 port map( A => n11952, B => n11951, ZN => n11953);
   U16375 : XNOR2_X1 port map( A => n11953, B => n12339, ZN => n11954);
   U16376 : XNOR2_X1 port map( A => n11954, B => n11955, ZN => n13275);
   U16377 : INV_X1 port map( A => n11956, ZN => n11964);
   U16378 : XNOR2_X1 port map( A => n11957, B => n896, ZN => n11958);
   U16379 : XNOR2_X1 port map( A => n12282, B => n11958, ZN => n11962);
   U16380 : XNOR2_X1 port map( A => n11960, B => n11959, ZN => n11961);
   U16381 : XNOR2_X1 port map( A => n11962, B => n11961, ZN => n11963);
   U16382 : XNOR2_X1 port map( A => n11966, B => n12130, ZN => n11969);
   U16383 : INV_X1 port map( A => n11967, ZN => n12352);
   U16384 : XNOR2_X1 port map( A => n12352, B => n2193, ZN => n11968);
   U16385 : XNOR2_X1 port map( A => n11969, B => n11968, ZN => n11973);
   U16386 : INV_X1 port map( A => n11970, ZN => n11971);
   U16387 : XNOR2_X1 port map( A => n12307, B => n11971, ZN => n11972);
   U16388 : NOR2_X1 port map( A1 => n24588, A2 => n13945, ZN => n13890);
   U16389 : XNOR2_X1 port map( A => n12401, B => n2236, ZN => n11976);
   U16390 : XNOR2_X1 port map( A => n11975, B => n11976, ZN => n11980);
   U16391 : INV_X1 port map( A => n12108, ZN => n11978);
   U16392 : XNOR2_X1 port map( A => n11977, B => n11978, ZN => n11979);
   U16393 : XNOR2_X1 port map( A => n12363, B => n11983, ZN => n11984);
   U16394 : XNOR2_X1 port map( A => n11985, B => n11984, ZN => n11989);
   U16395 : XNOR2_X1 port map( A => n12362, B => n876, ZN => n11987);
   U16396 : XNOR2_X1 port map( A => n11986, B => n11987, ZN => n11988);
   U16398 : XNOR2_X1 port map( A => n12102, B => n2772, ZN => n11990);
   U16399 : XNOR2_X1 port map( A => n11992, B => n12410, ZN => n11993);
   U16400 : XNOR2_X1 port map( A => n11994, B => n11993, ZN => n12680);
   U16401 : INV_X1 port map( A => n11995, ZN => n11997);
   U16402 : XNOR2_X1 port map( A => n11997, B => n11996, ZN => n12001);
   U16403 : XNOR2_X1 port map( A => n12196, B => n2726, ZN => n11998);
   U16404 : XNOR2_X1 port map( A => n11999, B => n11998, ZN => n12000);
   U16405 : XNOR2_X1 port map( A => n12002, B => n25396, ZN => n12004);
   U16406 : XNOR2_X1 port map( A => n12005, B => n12004, ZN => n12009);
   U16407 : XNOR2_X1 port map( A => n12357, B => n187, ZN => n12007);
   U16408 : XNOR2_X1 port map( A => n12356, B => n12127, ZN => n12006);
   U16409 : XNOR2_X1 port map( A => n12006, B => n12007, ZN => n12008);
   U16410 : XNOR2_X1 port map( A => n12008, B => n12009, ZN => n12934);
   U16411 : XNOR2_X1 port map( A => n12010, B => n12389, ZN => n12012);
   U16412 : XNOR2_X1 port map( A => n12012, B => n12011, ZN => n12015);
   U16413 : INV_X1 port map( A => n12013, ZN => n12014);
   U16414 : NAND2_X1 port map( A1 => n25015, A2 => n13264, ZN => n12016);
   U16415 : AOI21_X1 port map( B1 => n12829, B2 => n12016, A => n13265, ZN => 
                           n12017);
   U16416 : NOR2_X1 port map( A1 => n13890, A2 => n12018, ZN => n12177);
   U16417 : INV_X1 port map( A => n12019, ZN => n12022);
   U16418 : XNOR2_X1 port map( A => n12020, B => n12352, ZN => n12021);
   U16419 : XNOR2_X1 port map( A => n12022, B => n12021, ZN => n12027);
   U16420 : XNOR2_X1 port map( A => n12023, B => n1726, ZN => n12024);
   U16421 : XNOR2_X1 port map( A => n12029, B => n12030, ZN => n12035);
   U16422 : XNOR2_X1 port map( A => n12031, B => n12364, ZN => n12033);
   U16423 : XNOR2_X1 port map( A => n12234, B => n1804, ZN => n12032);
   U16424 : XNOR2_X1 port map( A => n12033, B => n12032, ZN => n12034);
   U16425 : INV_X1 port map( A => n12324, ZN => n12036);
   U16426 : XNOR2_X1 port map( A => n12036, B => n12409, ZN => n12037);
   U16427 : XNOR2_X1 port map( A => n12038, B => n12037, ZN => n12044);
   U16428 : XNOR2_X1 port map( A => n12039, B => n12212, ZN => n12042);
   U16429 : XNOR2_X1 port map( A => n12040, B => n891, ZN => n12041);
   U16430 : XNOR2_X1 port map( A => n12042, B => n12041, ZN => n12043);
   U16431 : INV_X1 port map( A => n12045, ZN => n12047);
   U16432 : XNOR2_X1 port map( A => n12047, B => n12046, ZN => n12052);
   U16433 : XNOR2_X1 port map( A => n12382, B => n12197, ZN => n12050);
   U16434 : XNOR2_X1 port map( A => n12048, B => n1768, ZN => n12049);
   U16435 : XNOR2_X1 port map( A => n12050, B => n12049, ZN => n12051);
   U16436 : XNOR2_X1 port map( A => n12052, B => n12051, ZN => n13328);
   U16437 : NAND2_X1 port map( A1 => n12684, A2 => n24422, ZN => n12062);
   U16438 : INV_X1 port map( A => n12053, ZN => n12054);
   U16439 : XNOR2_X1 port map( A => n12055, B => n12054, ZN => n12056);
   U16440 : XNOR2_X1 port map( A => n12056, B => n12057, ZN => n12061);
   U16441 : XNOR2_X1 port map( A => n12221, B => n21703, ZN => n12059);
   U16442 : XNOR2_X1 port map( A => n12058, B => n12059, ZN => n12060);
   U16443 : XNOR2_X1 port map( A => n12060, B => n12061, ZN => n12951);
   U16444 : INV_X1 port map( A => n12951, ZN => n13330);
   U16445 : XNOR2_X1 port map( A => n12064, B => n12063, ZN => n12071);
   U16446 : XNOR2_X1 port map( A => n12065, B => n12066, ZN => n12069);
   U16447 : XNOR2_X1 port map( A => n12067, B => n3183, ZN => n12068);
   U16448 : XNOR2_X1 port map( A => n12069, B => n12068, ZN => n12070);
   U16449 : NAND2_X1 port map( A1 => n24588, A2 => n14306, ZN => n12120);
   U16450 : XNOR2_X1 port map( A => n12074, B => n12073, ZN => n12079);
   U16451 : XNOR2_X1 port map( A => n12075, B => n12183, ZN => n12077);
   U16452 : XNOR2_X1 port map( A => n12128, B => n21623, ZN => n12076);
   U16453 : XNOR2_X1 port map( A => n12077, B => n12076, ZN => n12078);
   U16454 : XNOR2_X1 port map( A => n12080, B => n12081, ZN => n12086);
   U16455 : XNOR2_X1 port map( A => n12082, B => n12226, ZN => n12084);
   U16456 : XNOR2_X1 port map( A => n12159, B => n21711, ZN => n12083);
   U16457 : XNOR2_X1 port map( A => n12084, B => n12083, ZN => n12085);
   U16458 : XNOR2_X1 port map( A => n12086, B => n12085, ZN => n12840);
   U16459 : INV_X1 port map( A => n12840, ZN => n13338);
   U16460 : NOR2_X1 port map( A1 => n231, A2 => n13338, ZN => n12107);
   U16461 : XNOR2_X1 port map( A => n12087, B => n12088, ZN => n12093);
   U16462 : XNOR2_X1 port map( A => n24323, B => n1891, ZN => n12090);
   U16463 : XNOR2_X1 port map( A => n12091, B => n12090, ZN => n12092);
   U16464 : XNOR2_X1 port map( A => n12092, B => n12093, ZN => n12576);
   U16465 : XNOR2_X1 port map( A => n12095, B => n12094, ZN => n12100);
   U16466 : XNOR2_X1 port map( A => n12122, B => n1739, ZN => n12097);
   U16467 : XNOR2_X1 port map( A => n12098, B => n12097, ZN => n12099);
   U16468 : XNOR2_X1 port map( A => n12151, B => n11897, ZN => n12104);
   U16470 : AOI21_X1 port map( B1 => n13335, B2 => n13341, A => n231, ZN => 
                           n12119);
   U16471 : INV_X1 port map( A => n12839, ZN => n12118);
   U16472 : XNOR2_X1 port map( A => n12109, B => n12108, ZN => n12111);
   U16473 : XNOR2_X1 port map( A => n12110, B => n12111, ZN => n12116);
   U16474 : XNOR2_X1 port map( A => n25027, B => n3089, ZN => n12113);
   U16475 : NAND2_X1 port map( A1 => n231, A2 => n12956, ZN => n12642);
   U16476 : INV_X1 port map( A => n12642, ZN => n12117);
   U16477 : XNOR2_X1 port map( A => n12122, B => n1776, ZN => n12123);
   U16478 : XNOR2_X1 port map( A => n12124, B => n12123, ZN => n12125);
   U16479 : XNOR2_X1 port map( A => n12130, B => n12129, ZN => n12131);
   U16480 : INV_X1 port map( A => n12132, ZN => n12133);
   U16481 : INV_X1 port map( A => n13358, ZN => n13366);
   U16482 : XNOR2_X1 port map( A => n12134, B => n21335, ZN => n12135);
   U16483 : XNOR2_X1 port map( A => n12136, B => n12135, ZN => n12140);
   U16484 : XNOR2_X1 port map( A => n24970, B => n25236, ZN => n12139);
   U16485 : XNOR2_X1 port map( A => n12140, B => n12139, ZN => n12142);
   U16486 : XNOR2_X1 port map( A => n12142, B => n12141, ZN => n12625);
   U16487 : XNOR2_X1 port map( A => n12143, B => n20995, ZN => n12145);
   U16488 : XNOR2_X1 port map( A => n12145, B => n12144, ZN => n12149);
   U16489 : XNOR2_X1 port map( A => n12147, B => n12146, ZN => n12148);
   U16490 : XNOR2_X1 port map( A => n12149, B => n12148, ZN => n12155);
   U16491 : XNOR2_X1 port map( A => n12151, B => n25032, ZN => n12153);
   U16492 : XNOR2_X1 port map( A => n12152, B => n12153, ZN => n12154);
   U16493 : XNOR2_X2 port map( A => n12155, B => n12154, ZN => n12980);
   U16494 : INV_X1 port map( A => n12980, ZN => n13359);
   U16495 : AOI22_X1 port map( A1 => n24552, A2 => n13366, B1 => n12625, B2 => 
                           n13359, ZN => n12175);
   U16496 : INV_X1 port map( A => n12156, ZN => n12158);
   U16497 : XNOR2_X1 port map( A => n12157, B => n12158, ZN => n12164);
   U16498 : XNOR2_X1 port map( A => n12159, B => n22886, ZN => n12160);
   U16499 : XNOR2_X1 port map( A => n12160, B => n12391, ZN => n12162);
   U16500 : XNOR2_X1 port map( A => n12161, B => n12162, ZN => n12163);
   U16501 : XNOR2_X1 port map( A => n12164, B => n12163, ZN => n12583);
   U16503 : XNOR2_X1 port map( A => n12165, B => n12166, ZN => n12172);
   U16504 : XNOR2_X1 port map( A => n12167, B => n24323, ZN => n12170);
   U16505 : XNOR2_X1 port map( A => n12168, B => n1896, ZN => n12169);
   U16506 : XNOR2_X1 port map( A => n12170, B => n12169, ZN => n12171);
   U16507 : NAND2_X1 port map( A1 => n13358, A2 => n12976, ZN => n12626);
   U16508 : INV_X1 port map( A => n12626, ZN => n12173);
   U16509 : AOI22_X1 port map( A1 => n12173, A2 => n12878, B1 => n13366, B2 => 
                           n12980, ZN => n12174);
   U16510 : OAI21_X1 port map( B1 => n12175, B2 => n12977, A => n12174, ZN => 
                           n13453);
   U16511 : INV_X1 port map( A => n13453, ZN => n13947);
   U16512 : MUX2_X2 port map( A => n12177, B => n12176, S => n13947, Z => 
                           n15416);
   U16513 : XNOR2_X1 port map( A => n15416, B => n14732, ZN => n14691);
   U16514 : INV_X1 port map( A => n14691, ZN => n15176);
   U16515 : INV_X1 port map( A => n12178, ZN => n13093);
   U16516 : INV_X1 port map( A => n14311, ZN => n13733);
   U16517 : XNOR2_X1 port map( A => n12182, B => n12181, ZN => n12188);
   U16518 : XNOR2_X1 port map( A => n12184, B => n12183, ZN => n12185);
   U16519 : XNOR2_X1 port map( A => n12186, B => n12185, ZN => n12187);
   U16520 : INV_X1 port map( A => n12854, ZN => n13107);
   U16521 : XNOR2_X1 port map( A => n12334, B => n12189, ZN => n12191);
   U16522 : XNOR2_X1 port map( A => n12191, B => n12190, ZN => n12195);
   U16523 : XNOR2_X1 port map( A => n12193, B => n12192, ZN => n12194);
   U16524 : XNOR2_X1 port map( A => n12195, B => n12194, ZN => n13112);
   U16525 : INV_X1 port map( A => n13112, ZN => n12673);
   U16526 : XNOR2_X1 port map( A => n12197, B => n12196, ZN => n12199);
   U16527 : XNOR2_X1 port map( A => n12198, B => n12199, ZN => n12205);
   U16528 : XNOR2_X1 port map( A => n12344, B => n2042, ZN => n12203);
   U16529 : XNOR2_X1 port map( A => n12203, B => n12202, ZN => n12204);
   U16530 : NAND2_X1 port map( A1 => n3827, A2 => n12856, ZN => n12633);
   U16531 : XNOR2_X1 port map( A => n12209, B => n12208, ZN => n12211);
   U16532 : XNOR2_X1 port map( A => n12210, B => n12211, ZN => n12217);
   U16533 : XNOR2_X1 port map( A => n12214, B => n12215, ZN => n12216);
   U16534 : XNOR2_X1 port map( A => n12217, B => n12216, ZN => n12672);
   U16535 : INV_X1 port map( A => n12672, ZN => n13109);
   U16536 : XNOR2_X1 port map( A => n12219, B => n12220, ZN => n12223);
   U16537 : XNOR2_X1 port map( A => n12221, B => n12315, ZN => n12222);
   U16538 : XNOR2_X1 port map( A => n12223, B => n12222, ZN => n12229);
   U16539 : XNOR2_X1 port map( A => n12225, B => n12224, ZN => n12227);
   U16540 : XNOR2_X1 port map( A => n24915, B => n12227, ZN => n12228);
   U16541 : INV_X1 port map( A => n12230, ZN => n12232);
   U16542 : XNOR2_X1 port map( A => n12248, B => n12295, ZN => n12231);
   U16543 : XNOR2_X1 port map( A => n12232, B => n12231, ZN => n12238);
   U16544 : XNOR2_X1 port map( A => n12234, B => n20284, ZN => n12235);
   U16545 : XNOR2_X1 port map( A => n12236, B => n12235, ZN => n12237);
   U16546 : INV_X1 port map( A => n13110, ZN => n12674);
   U16547 : INV_X1 port map( A => n12239, ZN => n12240);
   U16548 : XNOR2_X1 port map( A => n12241, B => n1767, ZN => n12243);
   U16549 : XNOR2_X1 port map( A => n12243, B => n12242, ZN => n12244);
   U16550 : XNOR2_X1 port map( A => n12245, B => n12244, ZN => n12868);
   U16551 : XNOR2_X1 port map( A => n12247, B => n12246, ZN => n12254);
   U16552 : XNOR2_X1 port map( A => n12249, B => n12248, ZN => n12252);
   U16553 : XNOR2_X1 port map( A => n24323, B => n1826, ZN => n12251);
   U16554 : XNOR2_X1 port map( A => n12251, B => n12252, ZN => n12253);
   U16555 : XNOR2_X1 port map( A => n12255, B => n2120, ZN => n12256);
   U16556 : XNOR2_X1 port map( A => n12256, B => n12257, ZN => n12258);
   U16557 : XNOR2_X1 port map( A => n12258, B => n12259, ZN => n12265);
   U16558 : XNOR2_X1 port map( A => n12260, B => n24987, ZN => n12262);
   U16559 : XNOR2_X1 port map( A => n12263, B => n12262, ZN => n12264);
   U16561 : XNOR2_X1 port map( A => n12267, B => n12266, ZN => n12271);
   U16562 : INV_X1 port map( A => n12268, ZN => n12270);
   U16563 : NOR2_X1 port map( A1 => n12865, A2 => n12272, ZN => n12659);
   U16564 : XNOR2_X1 port map( A => n12274, B => n12273, ZN => n12281);
   U16565 : XNOR2_X1 port map( A => n12276, B => n12275, ZN => n12279);
   U16566 : XNOR2_X1 port map( A => n12277, B => n5131, ZN => n12278);
   U16567 : XNOR2_X1 port map( A => n12279, B => n12278, ZN => n12280);
   U16568 : XNOR2_X1 port map( A => n12281, B => n12280, ZN => n12864);
   U16569 : INV_X1 port map( A => n12864, ZN => n12503);
   U16570 : XNOR2_X1 port map( A => n12282, B => n12283, ZN => n12285);
   U16571 : XNOR2_X1 port map( A => n12285, B => n12284, ZN => n12290);
   U16572 : XNOR2_X1 port map( A => n12286, B => n1789, ZN => n12287);
   U16573 : XNOR2_X1 port map( A => n12288, B => n12287, ZN => n12289);
   U16574 : NOR2_X1 port map( A1 => n13114, A2 => n3327, ZN => n12291);
   U16575 : INV_X1 port map( A => n12292, ZN => n12294);
   U16576 : XNOR2_X1 port map( A => n12294, B => n12293, ZN => n12301);
   U16577 : XNOR2_X1 port map( A => n12295, B => n12296, ZN => n12299);
   U16578 : XNOR2_X1 port map( A => n12297, B => n2882, ZN => n12298);
   U16579 : XNOR2_X1 port map( A => n12299, B => n12298, ZN => n12300);
   U16580 : INV_X1 port map( A => n13123, ZN => n12874);
   U16581 : INV_X1 port map( A => n12302, ZN => n12305);
   U16582 : INV_X1 port map( A => n12303, ZN => n12304);
   U16583 : XNOR2_X1 port map( A => n12304, B => n12305, ZN => n12310);
   U16584 : XNOR2_X1 port map( A => n12306, B => n3084, ZN => n12308);
   U16585 : XNOR2_X1 port map( A => n12308, B => n12307, ZN => n12309);
   U16587 : XNOR2_X1 port map( A => n12312, B => n12311, ZN => n12319);
   U16588 : XNOR2_X1 port map( A => n12314, B => n12313, ZN => n12317);
   U16589 : XNOR2_X1 port map( A => n12315, B => n2240, ZN => n12316);
   U16590 : XNOR2_X1 port map( A => n12317, B => n12316, ZN => n12318);
   U16591 : XNOR2_X1 port map( A => n12319, B => n12318, ZN => n12349);
   U16592 : INV_X1 port map( A => n12320, ZN => n12321);
   U16593 : XNOR2_X1 port map( A => n12321, B => n12322, ZN => n12329);
   U16594 : XNOR2_X1 port map( A => n12324, B => n12323, ZN => n12327);
   U16595 : XNOR2_X1 port map( A => n12325, B => n1797, ZN => n12326);
   U16596 : XNOR2_X1 port map( A => n12327, B => n12326, ZN => n12328);
   U16597 : INV_X1 port map( A => n13354, ZN => n12332);
   U16598 : NAND2_X1 port map( A1 => n13352, A2 => n13123, ZN => n13122);
   U16599 : INV_X1 port map( A => n13122, ZN => n12331);
   U16600 : XNOR2_X1 port map( A => n12334, B => n12333, ZN => n12337);
   U16601 : XNOR2_X1 port map( A => n12335, B => n3073, ZN => n12336);
   U16602 : XNOR2_X1 port map( A => n12339, B => n12338, ZN => n12340);
   U16603 : XNOR2_X1 port map( A => n12343, B => n11915, ZN => n12346);
   U16604 : XNOR2_X1 port map( A => n12344, B => n899, ZN => n12345);
   U16605 : XNOR2_X1 port map( A => n12346, B => n12345, ZN => n12347);
   U16606 : INV_X1 port map( A => n12349, ZN => n13351);
   U16607 : NAND2_X1 port map( A1 => n406, A2 => n13351, ZN => n12350);
   U16608 : XNOR2_X1 port map( A => n12351, B => n12352, ZN => n12353);
   U16609 : XNOR2_X1 port map( A => n12354, B => n12353, ZN => n12361);
   U16610 : XNOR2_X1 port map( A => n12356, B => n12355, ZN => n12359);
   U16611 : XNOR2_X1 port map( A => n12357, B => n1833, ZN => n12358);
   U16612 : XNOR2_X1 port map( A => n12359, B => n12358, ZN => n12360);
   U16613 : XNOR2_X1 port map( A => n12362, B => n12363, ZN => n12367);
   U16614 : XNOR2_X1 port map( A => n12364, B => n12365, ZN => n12366);
   U16615 : XNOR2_X1 port map( A => n12366, B => n12367, ZN => n12374);
   U16616 : XNOR2_X1 port map( A => n12370, B => n4034, ZN => n12371);
   U16617 : XNOR2_X1 port map( A => n12372, B => n12371, ZN => n12373);
   U16618 : XNOR2_X1 port map( A => n12375, B => n12376, ZN => n12380);
   U16619 : XNOR2_X1 port map( A => n12378, B => n12377, ZN => n12379);
   U16620 : XNOR2_X1 port map( A => n12379, B => n12380, ZN => n12387);
   U16622 : XNOR2_X1 port map( A => n24964, B => n494, ZN => n12384);
   U16623 : XNOR2_X1 port map( A => n12385, B => n12384, ZN => n12386);
   U16624 : XNOR2_X1 port map( A => n12387, B => n12386, ZN => n12859);
   U16625 : XNOR2_X1 port map( A => n12388, B => n2031, ZN => n12390);
   U16626 : XNOR2_X1 port map( A => n12390, B => n12389, ZN => n12393);
   U16627 : XNOR2_X1 port map( A => n12393, B => n12392, ZN => n12394);
   U16629 : NAND2_X1 port map( A1 => n12859, A2 => n13344, ZN => n12407);
   U16630 : XNOR2_X1 port map( A => n12396, B => n23983, ZN => n12398);
   U16631 : XNOR2_X1 port map( A => n12398, B => n12397, ZN => n12399);
   U16632 : XNOR2_X1 port map( A => n12400, B => n12399, ZN => n12406);
   U16633 : XNOR2_X1 port map( A => n12402, B => n12401, ZN => n12403);
   U16634 : XNOR2_X1 port map( A => n12404, B => n12403, ZN => n12405);
   U16635 : XNOR2_X1 port map( A => n12406, B => n12405, ZN => n13347);
   U16636 : NAND2_X1 port map( A1 => n13347, A2 => n12636, ZN => n12419);
   U16637 : XNOR2_X1 port map( A => n12408, B => n2126, ZN => n12412);
   U16638 : XNOR2_X1 port map( A => n12412, B => n12411, ZN => n12418);
   U16639 : XNOR2_X1 port map( A => n12414, B => n12413, ZN => n12415);
   U16640 : XNOR2_X1 port map( A => n12416, B => n12415, ZN => n12417);
   U16642 : AOI21_X1 port map( B1 => n12419, B2 => n13345, A => n12859, ZN => 
                           n12420);
   U16643 : NOR2_X1 port map( A1 => n12421, A2 => n12420, ZN => n13903);
   U16644 : INV_X1 port map( A => n12422, ZN => n12424);
   U16645 : NOR3_X1 port map( A1 => n13903, A2 => n12424, A3 => n12423, ZN => 
                           n14310);
   U16646 : INV_X1 port map( A => n14310, ZN => n12425);
   U16647 : OAI21_X1 port map( B1 => n13959, B2 => n13958, A => n12425, ZN => 
                           n12427);
   U16648 : INV_X1 port map( A => n13132, ZN => n13129);
   U16649 : INV_X1 port map( A => n12498, ZN => n13131);
   U16650 : INV_X1 port map( A => n12483, ZN => n12712);
   U16651 : INV_X1 port map( A => n12707, ZN => n12711);
   U16652 : INV_X1 port map( A => n12710, ZN => n12431);
   U16653 : INV_X1 port map( A => n12433, ZN => n13145);
   U16654 : NAND3_X1 port map( A1 => n13145, A2 => n12729, A3 => n13144, ZN => 
                           n12438);
   U16655 : NAND2_X1 port map( A1 => n13144, A2 => n12455, ZN => n13146);
   U16656 : INV_X1 port map( A => n13146, ZN => n12434);
   U16657 : NAND2_X1 port map( A1 => n12434, A2 => n12728, ZN => n12436);
   U16658 : NAND3_X1 port map( A1 => n13140, A2 => n12729, A3 => n13143, ZN => 
                           n12435);
   U16659 : MUX2_X1 port map( A => n24601, B => n13061, S => n13063, Z => 
                           n12441);
   U16660 : NAND3_X1 port map( A1 => n13049, A2 => n12490, A3 => n12535, ZN => 
                           n12442);
   U16661 : NOR2_X1 port map( A1 => n14166, A2 => n14168, ZN => n12445);
   U16662 : INV_X1 port map( A => n12774, ZN => n13068);
   U16663 : NAND2_X1 port map( A1 => n13068, A2 => n12773, ZN => n12472);
   U16664 : NOR2_X1 port map( A1 => n13067, A2 => n12470, ZN => n12530);
   U16665 : INV_X1 port map( A => n12469, ZN => n12778);
   U16666 : OAI21_X1 port map( B1 => n12530, B2 => n1439, A => n12778, ZN => 
                           n12446);
   U16667 : AND2_X1 port map( A1 => n14165, A2 => n13744, ZN => n13745);
   U16668 : AOI21_X1 port map( B1 => n12718, B2 => n12447, A => n304, ZN => 
                           n12448);
   U16669 : NAND2_X1 port map( A1 => n13745, A2 => n13742, ZN => n13529);
   U16671 : MUX2_X1 port map( A => n13165, B => n24930, S => n24373, Z => 
                           n12453);
   U16672 : NAND2_X1 port map( A1 => n13170, A2 => n24930, ZN => n12452);
   U16673 : NAND2_X1 port map( A1 => n13137, A2 => n13144, ZN => n12458);
   U16674 : OAI211_X1 port map( C1 => n13144, C2 => n12455, A => n13140, B => 
                           n13136, ZN => n12457);
   U16675 : NAND3_X1 port map( A1 => n11109, A2 => n13138, A3 => n13143, ZN => 
                           n12456);
   U16676 : AOI21_X1 port map( B1 => n1355, B2 => n14049, A => n14050, ZN => 
                           n12468);
   U16677 : NAND2_X1 port map( A1 => n12462, A2 => n12715, ZN => n12482);
   U16678 : OAI21_X1 port map( B1 => n12710, B2 => n12707, A => n12713, ZN => 
                           n12461);
   U16679 : OAI21_X1 port map( B1 => n12712, B2 => n24573, A => n12710, ZN => 
                           n12463);
   U16680 : AOI22_X1 port map( A1 => n12490, A2 => n12534, B1 => n25408, B2 => 
                           n13049, ZN => n12466);
   U16681 : OAI21_X2 port map( B1 => n12466, B2 => n13048, A => n12465, ZN => 
                           n14054);
   U16682 : AND2_X1 port map( A1 => n14054, A2 => n13521, ZN => n13611);
   U16683 : NAND2_X1 port map( A1 => n14049, A2 => n14048, ZN => n12820);
   U16684 : INV_X1 port map( A => n12820, ZN => n12467);
   U16685 : XNOR2_X1 port map( A => n15054, B => n2005, ZN => n12518);
   U16686 : AND2_X1 port map( A1 => n12774, A2 => n12470, ZN => n13073);
   U16687 : AND2_X1 port map( A1 => n12469, A2 => n12470, ZN => n12532);
   U16688 : AOI21_X1 port map( B1 => n12774, B2 => n12471, A => n12470, ZN => 
                           n12473);
   U16689 : AND2_X1 port map( A1 => n12472, A2 => n12473, ZN => n12474);
   U16690 : INV_X1 port map( A => n12520, ZN => n12478);
   U16691 : NAND2_X1 port map( A1 => n12478, A2 => n12476, ZN => n12477);
   U16693 : NAND3_X1 port map( A1 => n12799, A2 => n12478, A3 => n13044, ZN => 
                           n12479);
   U16694 : NAND2_X1 port map( A1 => n12796, A2 => n12484, ZN => n12488);
   U16695 : NOR2_X1 port map( A1 => n25085, A2 => n409, ZN => n12486);
   U16696 : AOI22_X1 port map( A1 => n3065, A2 => n12486, B1 => n12485, B2 => 
                           n25085, ZN => n12487);
   U16697 : AOI22_X1 port map( A1 => n14241, A2 => n25209, B1 => n13931, B2 => 
                           n13200, ZN => n12497);
   U16698 : OAI211_X1 port map( C1 => n12534, C2 => n12535, A => n25494, B => 
                           n13048, ZN => n12492);
   U16699 : NAND3_X1 port map( A1 => n12490, A2 => n12489, A3 => n13051, ZN => 
                           n12491);
   U16700 : INV_X1 port map( A => n14244, ZN => n12496);
   U16702 : NAND2_X1 port map( A1 => n25369, A2 => n12786, ZN => n12493);
   U16703 : AOI22_X1 port map( A1 => n12494, A2 => n13029, B1 => n12493, B2 => 
                           n302, ZN => n13635);
   U16704 : INV_X1 port map( A => n13635, ZN => n14240);
   U16706 : NOR2_X1 port map( A1 => n13132, A2 => n13150, ZN => n12500);
   U16707 : NOR2_X1 port map( A1 => n13151, A2 => n12498, ZN => n12499);
   U16708 : NAND2_X1 port map( A1 => n13145, A2 => n13139, ZN => n12502);
   U16709 : NAND2_X1 port map( A1 => n14090, A2 => n13533, ZN => n12509);
   U16710 : AOI22_X1 port map( A1 => n12659, A2 => n12864, B1 => n13119, B2 => 
                           n13114, ZN => n13536);
   U16711 : NAND3_X1 port map( A1 => n3328, A2 => n12864, A3 => n12660, ZN => 
                           n12504);
   U16712 : NAND2_X1 port map( A1 => n5324, A2 => n13092, ZN => n12650);
   U16713 : MUX2_X1 port map( A => n12506, B => n10360, S => n12459, Z => 
                           n12508);
   U16714 : NAND2_X1 port map( A1 => n12652, A2 => n12724, ZN => n12507);
   U16715 : AOI21_X1 port map( B1 => n12509, B2 => n12817, A => n14018, ZN => 
                           n12515);
   U16717 : NAND2_X1 port map( A1 => n13102, A2 => n13187, ZN => n13183);
   U16718 : INV_X1 port map( A => n13187, ZN => n13103);
   U16719 : NAND2_X1 port map( A1 => n13103, A2 => n12656, ZN => n13191);
   U16720 : NAND3_X1 port map( A1 => n13183, A2 => n13185, A3 => n13191, ZN => 
                           n13535);
   U16721 : AOI21_X1 port map( B1 => n14085, B2 => n12513, A => n14090, ZN => 
                           n12514);
   U16722 : NOR2_X2 port map( A1 => n12515, A2 => n12514, ZN => n15056);
   U16723 : INV_X1 port map( A => n15056, ZN => n12516);
   U16724 : XNOR2_X1 port map( A => n14377, B => n12516, ZN => n12517);
   U16725 : XNOR2_X1 port map( A => n12518, B => n12517, ZN => n12620);
   U16726 : MUX2_X1 port map( A => n12800, B => n12523, S => n13041, Z => 
                           n12522);
   U16727 : NOR2_X1 port map( A1 => n13044, A2 => n12523, ZN => n12521);
   U16728 : NAND2_X1 port map( A1 => n12523, A2 => n13040, ZN => n13045);
   U16731 : NOR2_X1 port map( A1 => n12753, A2 => n25085, ZN => n12528);
   U16732 : NOR2_X2 port map( A1 => n12529, A2 => n12528, ZN => n13840);
   U16733 : NAND2_X1 port map( A1 => n12774, A2 => n13071, ZN => n12531);
   U16734 : NOR2_X1 port map( A1 => n13840, A2 => n397, ZN => n12537);
   U16735 : MUX2_X1 port map( A => n13023, B => n13028, S => n12786, Z => 
                           n12538);
   U16736 : NAND2_X1 port map( A1 => n12786, A2 => n13028, ZN => n13025);
   U16737 : INV_X1 port map( A => n13623, ZN => n12543);
   U16738 : AOI22_X1 port map( A1 => n12543, A2 => n13839, B1 => n12542, B2 => 
                           n13837, ZN => n12544);
   U16739 : NOR2_X1 port map( A1 => n12546, A2 => n13298, ZN => n12549);
   U16740 : NAND2_X1 port map( A1 => n13301, A2 => n12902, ZN => n12903);
   U16741 : NAND2_X1 port map( A1 => n12546, A2 => n12903, ZN => n13239);
   U16742 : NOR2_X1 port map( A1 => n13239, A2 => n405, ZN => n13853);
   U16743 : INV_X1 port map( A => n13211, ZN => n13205);
   U16744 : OAI21_X1 port map( B1 => n13205, B2 => n13207, A => n13213, ZN => 
                           n12550);
   U16745 : AND2_X1 port map( A1 => n13000, A2 => n13207, ZN => n13001);
   U16746 : NOR2_X1 port map( A1 => n12551, A2 => n13207, ZN => n12552);
   U16747 : NOR2_X2 port map( A1 => n12553, A2 => n12552, ZN => n12704);
   U16748 : INV_X1 port map( A => n12704, ZN => n14074);
   U16749 : OAI21_X1 port map( B1 => n12611, B2 => n12555, A => n12914, ZN => 
                           n12554);
   U16750 : NAND2_X1 port map( A1 => n24487, A2 => n12554, ZN => n12557);
   U16751 : INV_X1 port map( A => n13245, ZN => n12559);
   U16752 : NAND3_X1 port map( A1 => n13244, A2 => n13011, A3 => n12559, ZN => 
                           n12562);
   U16753 : NAND2_X1 port map( A1 => n12563, A2 => n13246, ZN => n12564);
   U16756 : NAND2_X1 port map( A1 => n13009, A2 => n13222, ZN => n12568);
   U16757 : OAI211_X1 port map( C1 => n24965, C2 => n13009, A => n24490, B => 
                           n12568, ZN => n12572);
   U16758 : OAI21_X1 port map( B1 => n14075, B2 => n14076, A => n14077, ZN => 
                           n12573);
   U16759 : NAND2_X1 port map( A1 => n12573, A2 => n12704, ZN => n12574);
   U16760 : XNOR2_X1 port map( A => n14857, B => n15169, ZN => n15408);
   U16761 : NOR2_X1 port map( A1 => n12838, A2 => n13336, ZN => n12579);
   U16764 : NAND2_X1 port map( A1 => n12577, A2 => n12839, ZN => n12578);
   U16765 : INV_X1 port map( A => n12688, ZN => n12947);
   U16766 : MUX2_X1 port map( A => n25053, B => n12980, S => n12976, Z => 
                           n12586);
   U16767 : INV_X1 port map( A => n24554, ZN => n13365);
   U16768 : AOI21_X1 port map( B1 => n12586, B2 => n13365, A => n12585, ZN => 
                           n13847);
   U16770 : OAI21_X1 port map( B1 => n13108, B2 => n12856, A => n12672, ZN => 
                           n12587);
   U16771 : NOR3_X1 port map( A1 => n13109, A2 => n13112, A3 => n13108, ZN => 
                           n12588);
   U16772 : MUX2_X1 port map( A => n25430, B => n13123, S => n13124, Z => 
                           n12590);
   U16773 : INV_X1 port map( A => n14064, ZN => n13426);
   U16775 : NOR2_X1 port map( A1 => n13291, A2 => n12593, ZN => n12596);
   U16778 : AND2_X1 port map( A1 => n12600, A2 => n13272, ZN => n12965);
   U16779 : NAND2_X1 port map( A1 => n13275, A2 => n12695, ZN => n12602);
   U16780 : NAND2_X1 port map( A1 => n12834, A2 => n13274, ZN => n12601);
   U16781 : MUX2_X1 port map( A => n12602, B => n12601, S => n24346, Z => 
                           n12603);
   U16782 : INV_X1 port map( A => n13325, ZN => n12683);
   U16783 : OAI21_X1 port map( B1 => n12955, B2 => n12604, A => n13329, ZN => 
                           n12605);
   U16784 : NAND2_X1 port map( A1 => n14849, A2 => n14852, ZN => n12617);
   U16785 : INV_X1 port map( A => n12900, ZN => n13282);
   U16787 : AND2_X1 port map( A1 => n12900, A2 => n11873, ZN => n12925);
   U16788 : NAND2_X1 port map( A1 => n12614, A2 => n24572, ZN => n12616);
   U16789 : AND2_X1 port map( A1 => n14059, A2 => n14278, ZN => n14280);
   U16790 : NAND2_X1 port map( A1 => n14280, A2 => n14849, ZN => n12615);
   U16791 : OAI211_X1 port map( C1 => n24572, C2 => n12617, A => n12616, B => 
                           n12615, ZN => n14721);
   U16793 : XNOR2_X1 port map( A => n14699, B => n15408, ZN => n12619);
   U16794 : INV_X1 port map( A => n13350, ZN => n13125);
   U16795 : NAND2_X1 port map( A1 => n5624, A2 => n12349, ZN => n12622);
   U16797 : INV_X1 port map( A => n12976, ZN => n13364);
   U16799 : INV_X1 port map( A => n12625, ZN => n13357);
   U16800 : INV_X1 port map( A => n12865, ZN => n13117);
   U16801 : INV_X1 port map( A => n12660, ZN => n13116);
   U16802 : OAI21_X1 port map( B1 => n3328, B2 => n13116, A => n13114, ZN => 
                           n12630);
   U16803 : NAND2_X1 port map( A1 => n12854, A2 => n13108, ZN => n12634);
   U16804 : NAND3_X1 port map( A1 => n12673, A2 => n4923, A3 => n13107, ZN => 
                           n12635);
   U16805 : NAND2_X1 port map( A1 => n3889, A2 => n3888, ZN => n12646);
   U16806 : NOR2_X1 port map( A1 => n25415, A2 => n25366, ZN => n12637);
   U16807 : INV_X1 port map( A => n14198, ZN => n14946);
   U16808 : MUX2_X1 port map( A => n13335, B => n12956, S => n13341, Z => 
                           n12644);
   U16809 : INV_X1 port map( A => n12960, ZN => n12643);
   U16810 : NAND2_X1 port map( A1 => n13336, A2 => n12956, ZN => n12640);
   U16811 : NAND2_X1 port map( A1 => n13337, A2 => n12640, ZN => n12641);
   U16813 : NAND2_X1 port map( A1 => n2570, A2 => n2684, ZN => n12645);
   U16814 : OAI21_X1 port map( B1 => n12646, B2 => n14946, A => n12645, ZN => 
                           n12647);
   U16815 : INV_X1 port map( A => n14988, ZN => n12679);
   U16817 : INV_X1 port map( A => n14003, ZN => n13484);
   U16818 : INV_X1 port map( A => n13102, ZN => n12744);
   U16819 : NAND2_X1 port map( A1 => n12744, A2 => n12656, ZN => n12655);
   U16820 : OAI211_X1 port map( C1 => n12744, C2 => n12742, A => n12655, B => 
                           n12654, ZN => n12658);
   U16821 : NAND3_X1 port map( A1 => n13185, A2 => n12656, A3 => n12740, ZN => 
                           n12657);
   U16822 : INV_X1 port map( A => n12668, ZN => n13486);
   U16823 : INV_X1 port map( A => n12659, ZN => n12662);
   U16824 : NOR2_X1 port map( A1 => n12868, A2 => n12660, ZN => n12661);
   U16825 : INV_X1 port map( A => n13130, ZN => n13149);
   U16826 : NOR2_X1 port map( A1 => n13129, A2 => n13149, ZN => n12665);
   U16827 : NOR2_X1 port map( A1 => n13131, A2 => n13152, ZN => n12664);
   U16828 : INV_X1 port map( A => n5754, ZN => n12667);
   U16829 : OAI22_X1 port map( A1 => n13158, A2 => n13150, B1 => n12667, B2 => 
                           n13130, ZN => n13660);
   U16830 : NAND2_X1 port map( A1 => n14002, A2 => n12669, ZN => n12670);
   U16832 : INV_X1 port map( A => n13262, ZN => n12676);
   U16833 : MUX2_X1 port map( A => n13265, B => n13266, S => n5361, Z => n12682
                           );
   U16835 : NAND2_X1 port map( A1 => n13329, A2 => n13323, ZN => n12685);
   U16836 : NAND2_X1 port map( A1 => n13788, A2 => n14143, ZN => n12703);
   U16839 : OAI21_X1 port map( B1 => n13316, B2 => n25499, A => n12945, ZN => 
                           n12689);
   U16840 : NOR2_X1 port map( A1 => n12827, A2 => n24476, ZN => n12691);
   U16841 : OAI21_X1 port map( B1 => n12692, B2 => n12691, A => n12690, ZN => 
                           n12693);
   U16842 : INV_X1 port map( A => n13275, ZN => n12964);
   U16843 : NOR2_X1 port map( A1 => n13785, A2 => n14143, ZN => n13789);
   U16844 : OAI21_X1 port map( B1 => n12897, B2 => n13282, A => n24988, ZN => 
                           n12699);
   U16845 : OAI21_X1 port map( B1 => n13789, B2 => n14142, A => n24347, ZN => 
                           n12701);
   U16848 : XNOR2_X1 port map( A => n15070, B => n15185, ZN => n12783);
   U16849 : MUX2_X1 port map( A => n12721, B => n12720, S => n24930, Z => 
                           n12722);
   U16851 : NOR2_X1 port map( A1 => n14440, A2 => n24556, ZN => n13257);
   U16853 : OAI211_X1 port map( C1 => n3974, C2 => n13178, A => n13177, B => 
                           n12724, ZN => n12727);
   U16855 : NAND2_X1 port map( A1 => n12728, A2 => n13136, ZN => n12731);
   U16857 : MUX2_X1 port map( A => n12731, B => n12730, S => n13138, Z => 
                           n12732);
   U16858 : OAI22_X1 port map( A1 => n24571, A2 => n24713, B1 => n14440, B2 => 
                           n14510, ZN => n12739);
   U16859 : NAND2_X1 port map( A1 => n12439, A2 => n1353, ZN => n12738);
   U16860 : NAND2_X1 port map( A1 => n25061, A2 => n13061, ZN => n12736);
   U16861 : NAND2_X1 port map( A1 => n12742, A2 => n24640, ZN => n12743);
   U16863 : INV_X1 port map( A => n13188, ZN => n12745);
   U16864 : AND2_X2 port map( A1 => n12746, A2 => n12745, ZN => n13693);
   U16865 : INV_X1 port map( A => n13693, ZN => n14507);
   U16866 : NOR2_X1 port map( A1 => n24556, A2 => n14507, ZN => n13260);
   U16867 : XNOR2_X1 port map( A => n14911, B => n1896, ZN => n12781);
   U16868 : NAND2_X1 port map( A1 => n14052, A2 => n14054, ZN => n12749);
   U16869 : NAND3_X1 port map( A1 => n13521, A2 => n14054, A3 => n1355, ZN => 
                           n12747);
   U16870 : INV_X1 port map( A => n15184, ZN => n12780);
   U16871 : NOR2_X1 port map( A1 => n12796, A2 => n13053, ZN => n12750);
   U16872 : NOR2_X1 port map( A1 => n12751, A2 => n12750, ZN => n12755);
   U16873 : NAND2_X1 port map( A1 => n13053, A2 => n13057, ZN => n12752);
   U16874 : AND2_X1 port map( A1 => n12753, A2 => n12752, ZN => n12754);
   U16875 : MUX2_X2 port map( A => n12755, B => n12754, S => n25085, Z => 
                           n14178);
   U16876 : NAND2_X1 port map( A1 => n12560, A2 => n13011, ZN => n12756);
   U16877 : INV_X1 port map( A => n13011, ZN => n13243);
   U16878 : OAI21_X1 port map( B1 => n13244, B2 => n13243, A => n13015, ZN => 
                           n12757);
   U16879 : AOI22_X1 port map( A1 => n13242, A2 => n13245, B1 => n13017, B2 => 
                           n12757, ZN => n13578);
   U16880 : INV_X1 port map( A => n12761, ZN => n12760);
   U16881 : INV_X1 port map( A => n12786, ZN => n12759);
   U16883 : NAND3_X1 port map( A1 => n2793, A2 => n12761, A3 => n13027, ZN => 
                           n12762);
   U16884 : NAND2_X1 port map( A1 => n24949, A2 => n13792, ZN => n12771);
   U16885 : NOR2_X1 port map( A1 => n4651, A2 => n13215, ZN => n12764);
   U16886 : NAND2_X1 port map( A1 => n12764, A2 => n13220, ZN => n12766);
   U16887 : NAND2_X1 port map( A1 => n12766, A2 => n12765, ZN => n12770);
   U16888 : INV_X1 port map( A => n13217, ZN => n12768);
   U16889 : INV_X1 port map( A => n12772, ZN => n13769);
   U16890 : AOI21_X1 port map( B1 => n13797, B2 => n12771, A => n13769, ZN => 
                           n12779);
   U16891 : AOI22_X1 port map( A1 => n13067, A2 => n13066, B1 => n12774, B2 => 
                           n12773, ZN => n12777);
   U16892 : NAND2_X1 port map( A1 => n12775, A2 => n13068, ZN => n12776);
   U16893 : XNOR2_X1 port map( A => n14669, B => n12780, ZN => n15367);
   U16894 : XNOR2_X1 port map( A => n15367, B => n12781, ZN => n12782);
   U16895 : XNOR2_X1 port map( A => n12783, B => n12782, ZN => n15822);
   U16897 : AND2_X1 port map( A1 => n12787, A2 => n25369, ZN => n12789);
   U16898 : NOR2_X1 port map( A1 => n14327, A2 => n14041, ZN => n12804);
   U16899 : NAND2_X1 port map( A1 => n12800, A2 => n12799, ZN => n12802);
   U16900 : NOR2_X1 port map( A1 => n13045, A2 => n11580, ZN => n12801);
   U16901 : AOI22_X1 port map( A1 => n5230, A2 => n12804, B1 => n14327, B2 => 
                           n12803, ZN => n12816);
   U16902 : MUX2_X1 port map( A => n25198, B => n13011, S => n12808, Z => 
                           n12805);
   U16904 : MUX2_X1 port map( A => n12810, B => n12809, S => n24512, Z => 
                           n12813);
   U16905 : NOR3_X1 port map( A1 => n298, A2 => n14330, A3 => n14324, ZN => 
                           n12815);
   U16906 : NAND2_X1 port map( A1 => n13741, A2 => n13742, ZN => n12818);
   U16907 : INV_X1 port map( A => n13742, ZN => n14169);
   U16908 : NAND3_X1 port map( A1 => n13526, A2 => n14169, A3 => n14167, ZN => 
                           n12819);
   U16909 : XNOR2_X1 port map( A => n14900, B => n1797, ZN => n12852);
   U16910 : NAND2_X1 port map( A1 => n12825, A2 => n13292, ZN => n13507);
   U16911 : NOR2_X1 port map( A1 => n12827, A2 => n13288, ZN => n12826);
   U16912 : NAND2_X1 port map( A1 => n13507, A2 => n13502, ZN => n13877);
   U16913 : INV_X1 port map( A => n12830, ZN => n12831);
   U16914 : OAI21_X1 port map( B1 => n12832, B2 => n2632, A => n12831, ZN => 
                           n12833);
   U16915 : MUX2_X1 port map( A => n13278, B => n13273, S => n1200, Z => n12837
                           );
   U16916 : AOI22_X1 port map( A1 => n12835, A2 => n13278, B1 => n13274, B2 => 
                           n12965, ZN => n12836);
   U16917 : INV_X1 port map( A => n12956, ZN => n12842);
   U16919 : OAI21_X1 port map( B1 => n12840, B2 => n13341, A => n13335, ZN => 
                           n12841);
   U16920 : INV_X1 port map( A => n14339, ZN => n14334);
   U16921 : NOR2_X1 port map( A1 => n14333, A2 => n14339, ZN => n14337);
   U16922 : NAND2_X1 port map( A1 => n13318, A2 => n12844, ZN => n12843);
   U16923 : INV_X1 port map( A => n13323, ZN => n12952);
   U16925 : NOR2_X1 port map( A1 => n13325, A2 => n3256, ZN => n12849);
   U16929 : XNOR2_X1 port map( A => n12852, B => n15347, ZN => n12908);
   U16931 : NAND3_X1 port map( A1 => n13109, A2 => n4923, A3 => n12856, ZN => 
                           n12857);
   U16932 : INV_X1 port map( A => n13344, ZN => n12860);
   U16933 : NOR2_X1 port map( A1 => n14321, A2 => n13871, ZN => n14457);
   U16934 : INV_X1 port map( A => n13114, ZN => n12869);
   U16935 : MUX2_X1 port map( A => n3328, B => n13116, S => n12869, Z => n12867
                           );
   U16936 : NOR2_X1 port map( A1 => n12864, A2 => n13113, ZN => n12866);
   U16937 : INV_X1 port map( A => n14460, ZN => n12883);
   U16938 : NAND2_X1 port map( A1 => n13124, A2 => n13351, ZN => n12872);
   U16939 : NOR2_X1 port map( A1 => n24552, A2 => n12977, ZN => n12876);
   U16940 : INV_X1 port map( A => n12981, ZN => n12877);
   U16941 : NAND2_X1 port map( A1 => n12877, A2 => n12878, ZN => n12880);
   U16942 : NAND2_X1 port map( A1 => n13366, A2 => n12976, ZN => n12879);
   U16943 : NAND2_X1 port map( A1 => n3401, A2 => n13868, ZN => n12881);
   U16944 : OAI22_X1 port map( A1 => n14459, A2 => n13868, B1 => n12881, B2 => 
                           n14321, ZN => n12882);
   U16945 : NOR2_X1 port map( A1 => n12884, A2 => n12924, ZN => n12888);
   U16946 : INV_X1 port map( A => n13223, ZN => n12919);
   U16948 : NAND2_X1 port map( A1 => n13208, A2 => n12891, ZN => n12896);
   U16949 : NOR2_X1 port map( A1 => n5418, A2 => n11360, ZN => n12894);
   U16950 : INV_X1 port map( A => n13208, ZN => n12893);
   U16951 : NOR2_X1 port map( A1 => n12899, A2 => n13282, ZN => n12898);
   U16952 : AOI21_X1 port map( B1 => n13283, B2 => n12900, A => n12899, ZN => 
                           n12901);
   U16953 : INV_X1 port map( A => n13806, ZN => n12905);
   U16954 : NOR2_X1 port map( A1 => n3859, A2 => n13305, ZN => n12904);
   U16955 : NOR2_X1 port map( A1 => n12905, A2 => n13513, ZN => n12906);
   U16956 : NOR2_X2 port map( A1 => n12907, A2 => n12906, ZN => n14936);
   U16957 : XNOR2_X1 port map( A => n14936, B => n14992, ZN => n14714);
   U16958 : XNOR2_X1 port map( A => n12908, B => n14714, ZN => n12909);
   U16959 : AOI21_X1 port map( B1 => n12911, B2 => n24476, A => n12910, ZN => 
                           n12912);
   U16960 : NOR3_X1 port map( A1 => n12824, A2 => n13292, A3 => n13291, ZN => 
                           n12913);
   U16961 : OAI21_X1 port map( B1 => n13307, B2 => n13304, A => n12915, ZN => 
                           n12916);
   U16962 : AND2_X1 port map( A1 => n12918, A2 => n13227, ZN => n12923);
   U16963 : NOR2_X1 port map( A1 => n12569, A2 => n13224, ZN => n12921);
   U16964 : OAI21_X1 port map( B1 => n12921, B2 => n12920, A => n12919, ZN => 
                           n12922);
   U16965 : INV_X1 port map( A => n12925, ZN => n12926);
   U16966 : NAND2_X1 port map( A1 => n12926, A2 => n12928, ZN => n12930);
   U16970 : NAND2_X1 port map( A1 => n12935, A2 => n13298, ZN => n13236);
   U16972 : NAND2_X1 port map( A1 => n25193, A2 => n14130, ZN => n12939);
   U16973 : INV_X1 port map( A => n13826, ZN => n12938);
   U16974 : AOI21_X1 port map( B1 => n13896, B2 => n12939, A => n12938, ZN => 
                           n12940);
   U16975 : NOR2_X2 port map( A1 => n12941, A2 => n12940, ZN => n14928);
   U16976 : NOR2_X1 port map( A1 => n12942, A2 => n12688, ZN => n12943);
   U16977 : MUX2_X1 port map( A => n12944, B => n12943, S => n13317, Z => 
                           n12950);
   U16979 : NOR2_X1 port map( A1 => n12948, A2 => n12947, ZN => n12949);
   U16980 : OAI211_X1 port map( C1 => n13329, C2 => n12952, A => n12951, B => 
                           n24422, ZN => n12954);
   U16981 : NAND3_X1 port map( A1 => n13330, A2 => n13327, A3 => n13323, ZN => 
                           n12953);
   U16982 : OR2_X1 port map( A1 => n14208, A2 => n14205, ZN => n12975);
   U16983 : NOR2_X1 port map( A1 => n231, A2 => n12956, ZN => n12957);
   U16984 : NOR3_X1 port map( A1 => n12960, A2 => n12959, A3 => n12958, ZN => 
                           n12961);
   U16985 : NAND3_X1 port map( A1 => n13278, A2 => n13272, A3 => n12964, ZN => 
                           n12970);
   U16986 : NAND2_X1 port map( A1 => n13273, A2 => n12966, ZN => n12967);
   U16987 : AND4_X2 port map( A1 => n12970, A2 => n12969, A3 => n12968, A4 => 
                           n12967, ZN => n13549);
   U16988 : NAND2_X1 port map( A1 => n14206, A2 => n13549, ZN => n12974);
   U16989 : AOI21_X1 port map( B1 => n398, B2 => n25415, A => n13345, ZN => 
                           n12971);
   U16990 : MUX2_X1 port map( A => n12975, B => n12974, S => n14123, Z => 
                           n12983);
   U16991 : NOR2_X1 port map( A1 => n13357, A2 => n25584, ZN => n12979);
   U16993 : NOR2_X1 port map( A1 => n12981, A2 => n12980, ZN => n13419);
   U16994 : INV_X1 port map( A => n14208, ZN => n13422);
   U16995 : NAND2_X1 port map( A1 => n12983, A2 => n12982, ZN => n14466);
   U16996 : INV_X1 port map( A => n14466, ZN => n15341);
   U16997 : XNOR2_X1 port map( A => n15341, B => n14928, ZN => n14677);
   U16998 : INV_X1 port map( A => n14222, ZN => n14218);
   U16999 : NAND2_X1 port map( A1 => n25080, A2 => n12993, ZN => n13231);
   U17000 : INV_X1 port map( A => n13231, ZN => n12996);
   U17001 : NAND2_X1 port map( A1 => n12996, A2 => n12995, ZN => n12997);
   U17002 : INV_X1 port map( A => n14219, ZN => n13032);
   U17003 : NAND2_X1 port map( A1 => n13211, A2 => n13000, ZN => n13003);
   U17004 : NAND2_X1 port map( A1 => n13001, A2 => n1335, ZN => n13002);
   U17005 : OAI21_X1 port map( B1 => n13003, B2 => n1335, A => n13002, ZN => 
                           n13008);
   U17006 : OAI22_X1 port map( A1 => n13006, A2 => n11684, B1 => n13005, B2 => 
                           n13004, ZN => n13007);
   U17007 : INV_X1 port map( A => n13830, ZN => n14223);
   U17008 : NAND2_X1 port map( A1 => n14223, A2 => n13829, ZN => n14226);
   U17009 : NOR2_X1 port map( A1 => n13011, A2 => n13014, ZN => n13021);
   U17010 : OAI21_X1 port map( B1 => n13013, B2 => n13246, A => n25199, ZN => 
                           n13020);
   U17011 : AOI22_X1 port map( A1 => n13018, A2 => n13017, B1 => n13016, B2 => 
                           n13015, ZN => n13019);
   U17012 : MUX2_X1 port map( A => n13022, B => n14226, S => n14225, Z => 
                           n13036);
   U17013 : INV_X1 port map( A => n14225, ZN => n13399);
   U17014 : NAND2_X1 port map( A1 => n13399, A2 => n13829, ZN => n13555);
   U17015 : INV_X1 port map( A => n13555, ZN => n13034);
   U17016 : NAND2_X1 port map( A1 => n13024, A2 => n13023, ZN => n13026);
   U17017 : NOR2_X1 port map( A1 => n13032, A2 => n14221, ZN => n13033);
   U17018 : AOI22_X1 port map( A1 => n13034, A2 => n14222, B1 => n14119, B2 => 
                           n13033, ZN => n13035);
   U17019 : MUX2_X1 port map( A => n13039, B => n13038, S => n13037, Z => 
                           n13043);
   U17020 : NOR2_X1 port map( A1 => n11580, A2 => n13040, ZN => n13042);
   U17022 : NOR2_X1 port map( A1 => n13045, A2 => n13044, ZN => n13046);
   U17024 : AOI21_X1 port map( B1 => n13054, B2 => n13053, A => n13052, ZN => 
                           n13060);
   U17025 : NAND2_X1 port map( A1 => n12526, A2 => n303, ZN => n13058);
   U17026 : NOR2_X1 port map( A1 => n13386, A2 => n24589, ZN => n13820);
   U17027 : NAND2_X1 port map( A1 => n24876, A2 => n13820, ZN => n13085);
   U17028 : INV_X1 port map( A => n13061, ZN => n13161);
   U17029 : INV_X1 port map( A => n13385, ZN => n13644);
   U17030 : INV_X1 port map( A => n13067, ZN => n13070);
   U17031 : NAND2_X1 port map( A1 => n13073, A2 => n13072, ZN => n13079);
   U17032 : NAND3_X1 port map( A1 => n13644, A2 => n24589, A3 => n392, ZN => 
                           n13084);
   U17033 : NOR2_X1 port map( A1 => n13074, A2 => n24573, ZN => n13075);
   U17034 : NOR2_X1 port map( A1 => n12709, A2 => n13075, ZN => n13081);
   U17035 : NAND2_X1 port map( A1 => n24589, A2 => n13647, ZN => n13082);
   U17036 : NAND3_X1 port map( A1 => n13559, A2 => n13082, A3 => n24507, ZN => 
                           n13083);
   U17037 : XNOR2_X1 port map( A => n14675, B => n15210, ZN => n15383);
   U17038 : XNOR2_X1 port map( A => n14677, B => n15383, ZN => n13199);
   U17039 : NAND2_X1 port map( A1 => n5526, A2 => n13394, ZN => n13571);
   U17040 : NOR3_X1 port map( A1 => n13087, A2 => n14360, A3 => n13086, ZN => 
                           n13573);
   U17041 : NOR2_X1 port map( A1 => n13394, A2 => n13589, ZN => n13090);
   U17042 : NAND2_X1 port map( A1 => n13712, A2 => n13090, ZN => n14366);
   U17043 : OAI211_X1 port map( C1 => n14361, C2 => n13571, A => n13091, B => 
                           n14366, ZN => n14345);
   U17044 : XNOR2_X1 port map( A => n14345, B => n3155, ZN => n13197);
   U17045 : NOR2_X1 port map( A1 => n13098, A2 => n13097, ZN => n13099);
   U17048 : NOR2_X1 port map( A1 => n13109, A2 => n13108, ZN => n13111);
   U17049 : INV_X1 port map( A => n13417, ZN => n14099);
   U17050 : MUX2_X1 port map( A => n13117, B => n13114, S => n13113, Z => 
                           n13120);
   U17051 : INV_X1 port map( A => n13115, ZN => n13118);
   U17052 : INV_X1 port map( A => n14101, ZN => n14213);
   U17053 : NAND2_X1 port map( A1 => n406, A2 => n12349, ZN => n13121);
   U17054 : AOI21_X1 port map( B1 => n13122, B2 => n13121, A => n13353, ZN => 
                           n13128);
   U17055 : NAND2_X1 port map( A1 => n13124, A2 => n13123, ZN => n13126);
   U17056 : OAI21_X1 port map( B1 => n13131, B2 => n13130, A => n13129, ZN => 
                           n13134);
   U17057 : NOR2_X1 port map( A1 => n13150, A2 => n13152, ZN => n13133);
   U17058 : NAND2_X1 port map( A1 => n12433, A2 => n13136, ZN => n13142);
   U17060 : MUX2_X1 port map( A => n13142, B => n13141, S => n13140, Z => 
                           n13193);
   U17061 : NAND2_X1 port map( A1 => n13144, A2 => n13143, ZN => n13147);
   U17062 : MUX2_X1 port map( A => n13147, B => n13146, S => n13145, Z => 
                           n13192);
   U17063 : NAND3_X1 port map( A1 => n13150, A2 => n13149, A3 => n13148, ZN => 
                           n13155);
   U17064 : AND3_X1 port map( A1 => n13155, A2 => n13154, A3 => n13153, ZN => 
                           n13156);
   U17065 : OAI21_X1 port map( B1 => n13158, B2 => n13157, A => n13156, ZN => 
                           n13565);
   U17066 : NOR2_X1 port map( A1 => n14106, A2 => n13565, ZN => n14111);
   U17067 : AOI22_X1 port map( A1 => n13168, A2 => n13167, B1 => n13166, B2 => 
                           n24373, ZN => n13173);
   U17068 : NAND2_X1 port map( A1 => n13175, A2 => n13174, ZN => n13181);
   U17069 : NAND3_X1 port map( A1 => n12459, A2 => n13176, A3 => n13178, ZN => 
                           n13180);
   U17070 : NAND3_X1 port map( A1 => n13181, A2 => n13180, A3 => n13179, ZN => 
                           n13583);
   U17071 : OAI21_X1 port map( B1 => n13566, B2 => n14105, A => n14112, ZN => 
                           n13182);
   U17072 : OAI21_X1 port map( B1 => n14111, B2 => n14112, A => n13182, ZN => 
                           n13196);
   U17073 : INV_X1 port map( A => n13183, ZN => n13186);
   U17074 : OAI21_X1 port map( B1 => n13186, B2 => n13185, A => n24640, ZN => 
                           n13190);
   U17076 : NAND3_X1 port map( A1 => n13193, A2 => n13192, A3 => n13582, ZN => 
                           n13194);
   U17077 : OAI211_X1 port map( C1 => n14112, C2 => n13582, A => n13194, B => 
                           n14105, ZN => n13195);
   U17078 : NAND2_X1 port map( A1 => n13196, A2 => n13195, ZN => n14865);
   U17079 : XNOR2_X1 port map( A => n14976, B => n14865, ZN => n15028);
   U17080 : XNOR2_X1 port map( A => n13197, B => n15028, ZN => n13198);
   U17081 : INV_X1 port map( A => n16597, ZN => n15890);
   U17082 : MUX2_X1 port map( A => n25209, B => n14244, S => n13636, Z => 
                           n13204);
   U17085 : OAI21_X1 port map( B1 => n13207, B2 => n13206, A => n5418, ZN => 
                           n13209);
   U17086 : NAND3_X1 port map( A1 => n13213, A2 => n13212, A3 => n11360, ZN => 
                           n13214);
   U17087 : NAND2_X1 port map( A1 => n4651, A2 => n13215, ZN => n13219);
   U17088 : NAND2_X1 port map( A1 => n13217, A2 => n12767, ZN => n13218);
   U17089 : AND2_X1 port map( A1 => n13988, A2 => n13981, ZN => n13241);
   U17090 : NAND2_X1 port map( A1 => n13223, A2 => n13222, ZN => n13226);
   U17091 : INV_X1 port map( A => n13918, ZN => n13653);
   U17092 : NOR2_X1 port map( A1 => n13230, A2 => n13229, ZN => n13233);
   U17093 : MUX2_X2 port map( A => n13233, B => n13232, S => n24750, Z => 
                           n13989);
   U17094 : NOR2_X1 port map( A1 => n13653, A2 => n13989, ZN => n13240);
   U17095 : MUX2_X1 port map( A => n13241, B => n13240, S => n13982, Z => 
                           n13251);
   U17096 : OAI211_X1 port map( C1 => n13246, C2 => n13245, A => n13244, B => 
                           n13243, ZN => n13247);
   U17097 : MUX2_X1 port map( A => n13987, B => n13988, S => n13981, Z => 
                           n13249);
   U17098 : INV_X1 port map( A => n13989, ZN => n13652);
   U17099 : NOR2_X1 port map( A1 => n13249, A2 => n13652, ZN => n13250);
   U17100 : NOR2_X2 port map( A1 => n13251, A2 => n13250, ZN => n14703);
   U17102 : NAND2_X1 port map( A1 => n13385, A2 => n13818, ZN => n13822);
   U17103 : INV_X1 port map( A => n13822, ZN => n13255);
   U17104 : INV_X1 port map( A => n13648, ZN => n13252);
   U17105 : NAND2_X1 port map( A1 => n13252, A2 => n13385, ZN => n13254);
   U17107 : OAI21_X1 port map( B1 => n13693, B2 => n24713, A => n24715, ZN => 
                           n13259);
   U17108 : NAND2_X1 port map( A1 => n13257, A2 => n13693, ZN => n14513);
   U17109 : NOR2_X1 port map( A1 => n14436, A2 => n14439, ZN => n14511);
   U17110 : NAND2_X1 port map( A1 => n14511, A2 => n14510, ZN => n13258);
   U17111 : OAI211_X1 port map( C1 => n13260, C2 => n13259, A => n14513, B => 
                           n13258, ZN => n13261);
   U17112 : XNOR2_X1 port map( A => n14952, B => n13261, ZN => n14287);
   U17113 : XNOR2_X1 port map( A => n15392, B => n14287, ZN => n13372);
   U17114 : XNOR2_X1 port map( A => n15062, B => n1935, ZN => n13370);
   U17115 : NAND2_X1 port map( A1 => n5361, A2 => n13265, ZN => n13269);
   U17116 : MUX2_X1 port map( A => n13269, B => n13268, S => n13267, Z => 
                           n13270);
   U17117 : OAI21_X1 port map( B1 => n5361, B2 => n13271, A => n13270, ZN => 
                           n14252);
   U17118 : NAND2_X1 port map( A1 => n13275, A2 => n13272, ZN => n13277);
   U17119 : INV_X1 port map( A => n14251, ZN => n14008);
   U17120 : NAND2_X1 port map( A1 => n24988, A2 => n12928, ZN => n13280);
   U17121 : NAND2_X1 port map( A1 => n13281, A2 => n13280, ZN => n13287);
   U17123 : INV_X1 port map( A => n13923, ZN => n14011);
   U17124 : NOR2_X1 port map( A1 => n13291, A2 => n24476, ZN => n13295);
   U17125 : NOR2_X1 port map( A1 => n25466, A2 => n12594, ZN => n13294);
   U17126 : NOR2_X2 port map( A1 => n13297, A2 => n13296, ZN => n14254);
   U17127 : NAND2_X1 port map( A1 => n545, A2 => n13298, ZN => n13300);
   U17128 : OAI22_X1 port map( A1 => n4493, A2 => n13300, B1 => n24220, B2 => 
                           n545, ZN => n13302);
   U17129 : NAND2_X1 port map( A1 => n14009, A2 => n14251, ZN => n13703);
   U17130 : OAI22_X1 port map( A1 => n13701, A2 => n14011, B1 => n14254, B2 => 
                           n13703, ZN => n13315);
   U17131 : NAND2_X1 port map( A1 => n14254, A2 => n14009, ZN => n13313);
   U17132 : INV_X1 port map( A => n14009, ZN => n14253);
   U17133 : NOR2_X1 port map( A1 => n13304, A2 => n13303, ZN => n13312);
   U17134 : OAI211_X1 port map( C1 => n13318, C2 => n13317, A => n25499, B => 
                           n13316, ZN => n13319);
   U17135 : INV_X1 port map( A => n13319, ZN => n13320);
   U17136 : NOR2_X1 port map( A1 => n13329, A2 => n13323, ZN => n13324);
   U17137 : NAND2_X1 port map( A1 => n5311, A2 => n13324, ZN => n13334);
   U17138 : NAND2_X1 port map( A1 => n13326, A2 => n13329, ZN => n13333);
   U17139 : NAND2_X1 port map( A1 => n5139, A2 => n13327, ZN => n13332);
   U17140 : NAND3_X1 port map( A1 => n13330, A2 => n4634, A3 => n24422, ZN => 
                           n13331);
   U17141 : AND2_X1 port map( A1 => n14230, A2 => n13682, ZN => n13356);
   U17142 : NAND2_X1 port map( A1 => n13345, A2 => n25415, ZN => n13346);
   U17144 : NOR2_X1 port map( A1 => n25053, A2 => n13357, ZN => n13362);
   U17145 : NOR2_X1 port map( A1 => n24552, A2 => n13359, ZN => n13361);
   U17146 : NAND3_X1 port map( A1 => n14231, A2 => n25434, A3 => n14233, ZN => 
                           n13368);
   U17147 : INV_X1 port map( A => n14231, ZN => n14234);
   U17148 : NAND3_X1 port map( A1 => n14234, A2 => n13995, A3 => n14233, ZN => 
                           n13367);
   U17149 : XNOR2_X1 port map( A => n15273, B => n15203, ZN => n14704);
   U17150 : XNOR2_X1 port map( A => n14704, B => n13370, ZN => n13371);
   U17151 : XNOR2_X1 port map( A => n13371, B => n13372, ZN => n15821);
   U17152 : NOR2_X1 port map( A1 => n24890, A2 => n24080, ZN => n13373);
   U17153 : NAND2_X1 port map( A1 => n13374, A2 => n15888, ZN => n13375);
   U17154 : INV_X1 port map( A => n14230, ZN => n13680);
   U17155 : NAND3_X1 port map( A1 => n14234, A2 => n25435, A3 => n13680, ZN => 
                           n13377);
   U17156 : OAI22_X1 port map( A1 => n25434, A2 => n24402, B1 => n14230, B2 => 
                           n13682, ZN => n13929);
   U17157 : NAND2_X1 port map( A1 => n13929, A2 => n13997, ZN => n13376);
   U17158 : NOR2_X1 port map( A1 => n13667, A2 => n14005, ZN => n13378);
   U17159 : NAND2_X1 port map( A1 => n13987, A2 => n13981, ZN => n13921);
   U17160 : AND2_X1 port map( A1 => n13988, A2 => n13987, ZN => n13655);
   U17161 : INV_X1 port map( A => n13981, ZN => n13379);
   U17163 : XNOR2_X1 port map( A => n14377, B => n14620, ZN => n13384);
   U17164 : INV_X1 port map( A => n14252, ZN => n14256);
   U17165 : NOR2_X1 port map( A1 => n14254, A2 => n13924, ZN => n13702);
   U17166 : OAI21_X1 port map( B1 => n13702, B2 => n14253, A => n14011, ZN => 
                           n13382);
   U17167 : INV_X1 port map( A => n3089, ZN => n22382);
   U17168 : XNOR2_X1 port map( A => n14694, B => n22382, ZN => n13383);
   U17169 : XNOR2_X1 port map( A => n13383, B => n13384, ZN => n13393);
   U17170 : NAND2_X1 port map( A1 => n13385, A2 => n13647, ZN => n13561);
   U17171 : NAND2_X1 port map( A1 => n25011, A2 => n13386, ZN => n13560);
   U17172 : AND2_X1 port map( A1 => n13818, A2 => n13647, ZN => n13387);
   U17173 : OAI21_X1 port map( B1 => n13387, B2 => n13644, A => n13646, ZN => 
                           n13388);
   U17174 : OAI211_X1 port map( C1 => n13561, C2 => n13824, A => n13389, B => 
                           n13388, ZN => n15229);
   U17175 : NOR2_X1 port map( A1 => n14510, A2 => n13693, ZN => n13390);
   U17176 : OAI22_X1 port map( A1 => n14436, A2 => n14507, B1 => n24556, B2 => 
                           n14510, ZN => n13392);
   U17177 : NOR2_X1 port map( A1 => n13712, A2 => n13569, ZN => n13713);
   U17179 : NOR2_X1 port map( A1 => n14361, A2 => n13394, ZN => n13395);
   U17180 : INV_X1 port map( A => n13396, ZN => n13397);
   U17182 : NOR2_X1 port map( A1 => n13829, A2 => n14219, ZN => n13404);
   U17183 : XNOR2_X1 port map( A => n14952, B => n24418, ZN => n13405);
   U17184 : NAND3_X1 port map( A1 => n14127, A2 => n1331, A3 => n4844, ZN => 
                           n13409);
   U17185 : INV_X1 port map( A => n14130, ZN => n13894);
   U17186 : NAND3_X1 port map( A1 => n13894, A2 => n13893, A3 => n14127, ZN => 
                           n13408);
   U17187 : NAND4_X2 port map( A1 => n13408, A2 => n13410, A3 => n13409, A4 => 
                           n13407, ZN => n15396);
   U17188 : XNOR2_X1 port map( A => n15396, B => n1792, ZN => n13416);
   U17189 : NAND2_X1 port map( A1 => n14106, A2 => n13565, ZN => n13413);
   U17190 : NAND2_X1 port map( A1 => n14107, A2 => n4868, ZN => n13411);
   U17191 : MUX2_X1 port map( A => n13413, B => n13411, S => n5333, Z => n13415
                           );
   U17192 : INV_X1 port map( A => n13565, ZN => n13584);
   U17193 : AOI21_X1 port map( B1 => n13584, B2 => n14108, A => n14105, ZN => 
                           n13412);
   U17194 : NAND2_X1 port map( A1 => n13413, A2 => n13412, ZN => n13414);
   U17195 : NAND2_X1 port map( A1 => n13415, A2 => n13414, ZN => n13873);
   U17196 : INV_X1 port map( A => n13873, ZN => n15199);
   U17197 : XNOR2_X1 port map( A => n13416, B => n15199, ZN => n13423);
   U17198 : OAI21_X1 port map( B1 => n13417, B2 => n14211, A => n14213, ZN => 
                           n13418);
   U17199 : NOR2_X1 port map( A1 => n14124, A2 => n13419, ZN => n13420);
   U17200 : NAND2_X1 port map( A1 => n13421, A2 => n13420, ZN => n13548);
   U17201 : XNOR2_X1 port map( A => n14834, B => n15463, ZN => n15270);
   U17202 : XNOR2_X1 port map( A => n13423, B => n15270, ZN => n13424);
   U17203 : INV_X1 port map( A => n15915, ZN => n16336);
   U17204 : INV_X1 port map( A => n13845, ZN => n13844);
   U17205 : NOR2_X1 port map( A1 => n14063, A2 => n13844, ZN => n13425);
   U17206 : NAND2_X1 port map( A1 => n13426, A2 => n13425, ZN => n13431);
   U17207 : NAND2_X1 port map( A1 => n13427, A2 => n13845, ZN => n14069);
   U17208 : NOR2_X1 port map( A1 => n13843, A2 => n13845, ZN => n13428);
   U17209 : NAND2_X1 port map( A1 => n14064, A2 => n13428, ZN => n13429);
   U17210 : NAND2_X1 port map( A1 => n13566, A2 => n14108, ZN => n13436);
   U17211 : OAI21_X1 port map( B1 => n5333, B2 => n13566, A => n13584, ZN => 
                           n13432);
   U17213 : NOR2_X1 port map( A1 => n5333, A2 => n14105, ZN => n13433);
   U17214 : NAND2_X1 port map( A1 => n13433, A2 => n13566, ZN => n13434);
   U17216 : INV_X1 port map( A => n13552, ZN => n14216);
   U17217 : NAND2_X1 port map( A1 => n14216, A2 => n24376, ZN => n13440);
   U17218 : OAI21_X1 port map( B1 => n13417, B2 => n13552, A => n25445, ZN => 
                           n13438);
   U17219 : XNOR2_X1 port map( A => n15183, B => n1870, ZN => n13441);
   U17220 : INV_X1 port map( A => n13982, ZN => n13922);
   U17221 : OAI21_X1 port map( B1 => n13918, B2 => n13989, A => n13922, ZN => 
                           n13443);
   U17222 : INV_X1 port map( A => n13988, ZN => n13656);
   U17223 : INV_X1 port map( A => n13917, ZN => n13986);
   U17224 : OAI21_X1 port map( B1 => n13656, B2 => n13981, A => n13986, ZN => 
                           n13442);
   U17228 : NAND3_X1 port map( A1 => n24572, A2 => n24958, A3 => n14852, ZN => 
                           n13446);
   U17229 : NAND3_X1 port map( A1 => n14849, A2 => n14850, A3 => n14852, ZN => 
                           n13445);
   U17231 : NOR2_X1 port map( A1 => n14271, A2 => n13840, ZN => n13761);
   U17233 : NOR3_X1 port map( A1 => n24368, A2 => n397, A3 => n14268, ZN => 
                           n13449);
   U17234 : AOI21_X1 port map( B1 => n3947, B2 => n16336, A => n290, ZN => 
                           n13547);
   U17241 : MUX2_X1 port map( A => n13459, B => n13458, S => n14307, Z => 
                           n13462);
   U17242 : XNOR2_X1 port map( A => n14477, B => n14676, ZN => n15290);
   U17243 : INV_X1 port map( A => n14289, ZN => n14293);
   U17244 : NAND3_X1 port map( A1 => n14293, A2 => n13909, A3 => n394, ZN => 
                           n13465);
   U17245 : AOI21_X1 port map( B1 => n13909, B2 => n24974, A => n14294, ZN => 
                           n13463);
   U17246 : XNOR2_X1 port map( A => n14345, B => n14468, ZN => n14933);
   U17247 : XNOR2_X1 port map( A => n15290, B => n14933, ZN => n13476);
   U17248 : NAND2_X1 port map( A1 => n14172, A2 => n14168, ZN => n13527);
   U17249 : NOR2_X1 port map( A1 => n13775, A2 => n13954, ZN => n13716);
   U17250 : AOI22_X1 port map( A1 => n13716, A2 => n14156, B1 => n13467, B2 => 
                           n13954, ZN => n13468);
   U17251 : OAI21_X2 port map( B1 => n14160, B2 => n13469, A => n13468, ZN => 
                           n15386);
   U17252 : XNOR2_X1 port map( A => n14979, B => n15386, ZN => n13474);
   U17253 : AOI22_X1 port map( A1 => n13969, A2 => n13596, B1 => n13470, B2 => 
                           n13968, ZN => n13471);
   U17254 : INV_X1 port map( A => n1726, ZN => n13472);
   U17255 : XNOR2_X1 port map( A => n15488, B => n13472, ZN => n13473);
   U17256 : XNOR2_X1 port map( A => n13474, B => n13473, ZN => n13475);
   U17258 : AND2_X1 port map( A1 => n13785, A2 => n14142, ZN => n13477);
   U17259 : AND2_X1 port map( A1 => n14144, A2 => n14199, ZN => n13481);
   U17261 : INV_X1 port map( A => n13804, ZN => n13480);
   U17262 : NOR2_X1 port map( A1 => n14200, A2 => n3888, ZN => n13479);
   U17264 : NOR2_X1 port map( A1 => n13792, A2 => n13795, ZN => n13482);
   U17265 : INV_X1 port map( A => n14178, ZN => n13580);
   U17266 : OAI21_X1 port map( B1 => n13482, B2 => n13580, A => n14182, ZN => 
                           n13483);
   U17267 : XNOR2_X1 port map( A => n14900, B => n15190, ZN => n14940);
   U17268 : INV_X1 port map( A => n14078, ZN => n14073);
   U17269 : OAI21_X1 port map( B1 => n13491, B2 => n13628, A => n13629, ZN => 
                           n13492);
   U17270 : XNOR2_X1 port map( A => n15191, B => n15514, ZN => n13497);
   U17271 : OAI211_X1 port map( C1 => n14439, C2 => n13974, A => n24556, B => 
                           n24713, ZN => n13495);
   U17272 : NAND3_X1 port map( A1 => n14440, A2 => n13693, A3 => n13975, ZN => 
                           n13494);
   U17273 : AND3_X1 port map( A1 => n13978, A2 => n13495, A3 => n13494, ZN => 
                           n14996);
   U17274 : INV_X1 port map( A => n14996, ZN => n14549);
   U17275 : XNOR2_X1 port map( A => n14549, B => n2772, ZN => n13496);
   U17276 : XNOR2_X1 port map( A => n13497, B => n13496, ZN => n13498);
   U17277 : NOR2_X1 port map( A1 => n16332, A2 => n25092, ZN => n13545);
   U17278 : INV_X1 port map( A => n14333, ZN => n13593);
   U17279 : INV_X1 port map( A => n25196, ZN => n13501);
   U17280 : INV_X1 port map( A => n13504, ZN => n13505);
   U17281 : OAI211_X1 port map( C1 => n25197, C2 => n14025, A => n14334, B => 
                           n13508, ZN => n13510);
   U17282 : NAND3_X1 port map( A1 => n14336, A2 => n13593, A3 => n14339, ZN => 
                           n13509);
   U17283 : XNOR2_X1 port map( A => n14880, B => n14815, ZN => n15281);
   U17284 : NOR2_X1 port map( A1 => n13807, A2 => n14149, ZN => n13512);
   U17285 : OAI21_X1 port map( B1 => n13515, B2 => n14153, A => n13514, ZN => 
                           n13516);
   U17286 : NOR2_X1 port map( A1 => n13614, A2 => n1355, ZN => n13520);
   U17287 : NAND2_X1 port map( A1 => n13612, A2 => n13610, ZN => n13519);
   U17289 : NOR2_X1 port map( A1 => n14325, A2 => n14041, ZN => n13590);
   U17290 : OAI21_X1 port map( B1 => n14172, B2 => n13741, A => n13526, ZN => 
                           n13531);
   U17291 : INV_X1 port map( A => n13527, ZN => n13530);
   U17292 : NAND3_X1 port map( A1 => n13741, A2 => n14164, A3 => n13744, ZN => 
                           n13528);
   U17293 : OAI211_X1 port map( C1 => n13531, C2 => n13530, A => n13529, B => 
                           n13528, ZN => n13532);
   U17294 : NAND4_X1 port map( A1 => n13538, A2 => n13537, A3 => n13536, A4 => 
                           n13535, ZN => n13539);
   U17295 : AOI21_X1 port map( B1 => n13540, B2 => n13539, A => n14088, ZN => 
                           n13541);
   U17296 : XNOR2_X1 port map( A => n15178, B => n4711, ZN => n13543);
   U17297 : XNOR2_X1 port map( A => n14964, B => n13543, ZN => n13544);
   U17298 : NOR2_X1 port map( A1 => n16331, A2 => n15667, ZN => n16337);
   U17299 : OAI21_X1 port map( B1 => n13545, B2 => n16337, A => n15915, ZN => 
                           n13546);
   U17300 : INV_X1 port map( A => n13813, ZN => n13550);
   U17302 : NOR2_X1 port map( A1 => n14101, A2 => n4894, ZN => n13554);
   U17303 : OAI21_X1 port map( B1 => n14217, B2 => n13554, A => n13553, ZN => 
                           n15194);
   U17304 : XNOR2_X1 port map( A => n14993, B => n15194, ZN => n15513);
   U17305 : OAI211_X1 port map( C1 => n14223, C2 => n13829, A => n14218, B => 
                           n14219, ZN => n13557);
   U17307 : XNOR2_X1 port map( A => n15444, B => n173, ZN => n13558);
   U17308 : XNOR2_X1 port map( A => n15513, B => n13558, ZN => n13577);
   U17309 : INV_X1 port map( A => n13561, ZN => n13564);
   U17310 : NAND2_X1 port map( A1 => n13824, A2 => n24589, ZN => n13563);
   U17311 : OAI211_X1 port map( C1 => n13561, C2 => n25011, A => n13560, B => 
                           n13559, ZN => n13562);
   U17313 : INV_X1 port map( A => n14106, ZN => n14109);
   U17314 : INV_X1 port map( A => n13581, ZN => n13567);
   U17315 : XNOR2_X1 port map( A => n14667, B => n15244, ZN => n14770);
   U17316 : AND2_X1 port map( A1 => n14132, A2 => n13895, ZN => n13575);
   U17317 : NAND3_X1 port map( A1 => n14127, A2 => n14126, A3 => n14132, ZN => 
                           n13574);
   U17318 : XNOR2_X1 port map( A => n14488, B => n15034, ZN => n14825);
   U17319 : XNOR2_X1 port map( A => n14825, B => n14770, ZN => n13576);
   U17320 : INV_X1 port map( A => n16200, ZN => n16403);
   U17321 : NOR2_X1 port map( A1 => n14178, A2 => n13578, ZN => n13793);
   U17322 : XNOR2_X1 port map( A => n15165, B => n729, ZN => n13585);
   U17323 : INV_X1 port map( A => n14361, ZN => n13586);
   U17324 : INV_X1 port map( A => n13712, ZN => n14364);
   U17325 : NAND3_X1 port map( A1 => n24995, A2 => n14364, A3 => n3701, ZN => 
                           n13588);
   U17326 : NOR2_X1 port map( A1 => n13590, A2 => n14328, ZN => n13591);
   U17327 : INV_X1 port map( A => n25413, ZN => n13592);
   U17328 : XNOR2_X1 port map( A => n15230, B => n13592, ZN => n14763);
   U17329 : INV_X1 port map( A => n14336, ZN => n14026);
   U17330 : INV_X1 port map( A => n13877, ZN => n14340);
   U17331 : OAI21_X2 port map( B1 => n13595, B2 => n14026, A => n13594, ZN => 
                           n15051);
   U17333 : XNOR2_X1 port map( A => n15051, B => n15430, ZN => n13605);
   U17335 : XNOR2_X1 port map( A => n13605, B => n25431, ZN => n14633);
   U17337 : NAND2_X1 port map( A1 => n14017, A2 => n14089, ZN => n13608);
   U17338 : NAND2_X1 port map( A1 => n14054, A2 => n14049, ZN => n13613);
   U17339 : OAI22_X1 port map( A1 => n13614, A2 => n13613, B1 => n14054, B2 => 
                           n13612, ZN => n13615);
   U17340 : XNOR2_X1 port map( A => n14755, B => n15487, ZN => n15241);
   U17341 : NOR2_X1 port map( A1 => n14059, A2 => n14852, ZN => n13617);
   U17342 : NAND2_X1 port map( A1 => n14267, A2 => n14269, ZN => n13621);
   U17343 : OR2_X1 port map( A1 => n13840, A2 => n14269, ZN => n13620);
   U17345 : AOI21_X1 port map( B1 => n13621, B2 => n13620, A => n123, ZN => 
                           n13625);
   U17346 : OAI21_X1 port map( B1 => n13839, B2 => n13623, A => n13622, ZN => 
                           n13624);
   U17348 : INV_X1 port map( A => n14678, ZN => n14756);
   U17349 : XNOR2_X1 port map( A => n14756, B => n14789, ZN => n13626);
   U17350 : XNOR2_X1 port map( A => n13626, B => n15241, ZN => n13642);
   U17351 : OAI211_X1 port map( C1 => n14076, C2 => n14078, A => n13629, B => 
                           n14074, ZN => n13630);
   U17352 : XNOR2_X1 port map( A => n15486, B => n15436, ZN => n14649);
   U17353 : NAND2_X1 port map( A1 => n14240, A2 => n14244, ZN => n13634);
   U17354 : OAI211_X1 port map( C1 => n13633, C2 => n14244, A => n4116, B => 
                           n13634, ZN => n13638);
   U17358 : XNOR2_X1 port map( A => n14792, B => n1865, ZN => n13640);
   U17359 : XNOR2_X1 port map( A => n14649, B => n13640, ZN => n13641);
   U17360 : NOR2_X1 port map( A1 => n13989, A2 => n13656, ZN => n13654);
   U17361 : INV_X1 port map( A => n13655, ZN => n13658);
   U17362 : NAND2_X1 port map( A1 => n13656, A2 => n13981, ZN => n13657);
   U17363 : XNOR2_X1 port map( A => n14644, B => n14816, ZN => n13691);
   U17364 : INV_X1 port map( A => n13659, ZN => n13666);
   U17365 : AOI21_X1 port map( B1 => n13661, B2 => n13662, A => n13660, ZN => 
                           n13665);
   U17366 : NAND2_X1 port map( A1 => n13663, A2 => n13662, ZN => n13664);
   U17367 : INV_X1 port map( A => n13668, ZN => n13673);
   U17368 : INV_X1 port map( A => n13669, ZN => n13672);
   U17369 : INV_X1 port map( A => n13670, ZN => n13671);
   U17370 : NAND3_X1 port map( A1 => n13673, A2 => n13672, A3 => n13671, ZN => 
                           n13674);
   U17371 : NAND2_X1 port map( A1 => n14003, A2 => n13676, ZN => n13677);
   U17372 : OAI21_X2 port map( B1 => n13679, B2 => n13678, A => n13677, ZN => 
                           n15175);
   U17373 : NAND2_X1 port map( A1 => n13680, A2 => n13683, ZN => n13688);
   U17374 : NAND2_X1 port map( A1 => n13680, A2 => n13681, ZN => n13687);
   U17375 : NOR2_X1 port map( A1 => n13682, A2 => n13681, ZN => n13685);
   U17376 : INV_X1 port map( A => n13683, ZN => n13684);
   U17377 : AOI21_X1 port map( B1 => n13685, B2 => n13684, A => n24402, ZN => 
                           n13686);
   U17378 : NAND3_X1 port map( A1 => n13688, A2 => n13687, A3 => n13686, ZN => 
                           n13690);
   U17379 : NOR2_X1 port map( A1 => n24556, A2 => n14439, ZN => n13692);
   U17380 : MUX2_X1 port map( A => n14511, B => n13692, S => n14510, Z => 
                           n13696);
   U17383 : OAI21_X1 port map( B1 => n14440, B2 => n14509, A => n14434, ZN => 
                           n13695);
   U17384 : NOR2_X1 port map( A1 => n13696, A2 => n13695, ZN => n13700);
   U17387 : XNOR2_X1 port map( A => n14690, B => n13700, ZN => n14781);
   U17388 : INV_X1 port map( A => n14254, ZN => n14250);
   U17389 : NAND3_X1 port map( A1 => n14250, A2 => n14008, A3 => n13923, ZN => 
                           n13706);
   U17390 : NAND2_X1 port map( A1 => n13702, A2 => n14251, ZN => n13705);
   U17392 : XNOR2_X1 port map( A => n24938, B => n20046, ZN => n13708);
   U17393 : XNOR2_X1 port map( A => n14781, B => n13708, ZN => n13709);
   U17394 : AND3_X1 port map( A1 => n14361, A2 => n13712, A3 => n14360, ZN => 
                           n13714);
   U17395 : NOR2_X1 port map( A1 => n13714, A2 => n13713, ZN => n13715);
   U17396 : INV_X1 port map( A => n13716, ZN => n13955);
   U17397 : NAND2_X1 port map( A1 => n14156, A2 => n5080, ZN => n13717);
   U17398 : NAND2_X1 port map( A1 => n13955, A2 => n13717, ZN => n13721);
   U17399 : NAND2_X1 port map( A1 => n13718, A2 => n13776, ZN => n13720);
   U17400 : XNOR2_X1 port map( A => n14671, B => n15253, ZN => n14749);
   U17401 : INV_X1 port map( A => n24973, ZN => n14292);
   U17402 : NAND2_X1 port map( A1 => n14289, A2 => n13907, ZN => n13723);
   U17403 : XNOR2_X1 port map( A => n15452, B => n15074, ZN => n14653);
   U17404 : XNOR2_X1 port map( A => n14653, B => n14749, ZN => n13738);
   U17405 : AOI21_X1 port map( B1 => n13892, B2 => n14306, A => n13947, ZN => 
                           n13729);
   U17406 : INV_X1 port map( A => n13892, ZN => n13728);
   U17407 : OAI21_X1 port map( B1 => n13959, B2 => n13900, A => n13956, ZN => 
                           n13732);
   U17408 : NAND2_X1 port map( A1 => n14311, A2 => n14307, ZN => n13730);
   U17409 : NAND2_X1 port map( A1 => n13900, A2 => n4525, ZN => n14314);
   U17410 : OAI21_X1 port map( B1 => n13730, B2 => n13958, A => n14314, ZN => 
                           n13731);
   U17411 : INV_X1 port map( A => n14168, ZN => n13743);
   U17412 : XNOR2_X1 port map( A => n14800, B => n1724, ZN => n13736);
   U17413 : XNOR2_X1 port map( A => n14389, B => n13736, ZN => n13737);
   U17414 : INV_X1 port map( A => n13785, ZN => n14191);
   U17415 : MUX2_X1 port map( A => n14189, B => n14141, S => n14190, Z => 
                           n13739);
   U17416 : NOR2_X1 port map( A1 => n25560, A2 => n13739, ZN => n13740);
   U17417 : OAI21_X1 port map( B1 => n14164, B2 => n13741, A => n14172, ZN => 
                           n13749);
   U17418 : NOR2_X1 port map( A1 => n14167, A2 => n13742, ZN => n13748);
   U17419 : NOR2_X1 port map( A1 => n13744, A2 => n13743, ZN => n13746);
   U17420 : AOI22_X1 port map( A1 => n14166, A2 => n13746, B1 => n13745, B2 => 
                           n14167, ZN => n13747);
   U17421 : XNOR2_X1 port map( A => n15318, B => n15219, ZN => n13756);
   U17422 : OR2_X1 port map( A1 => n14035, A2 => n14149, ZN => n14033);
   U17423 : OAI211_X1 port map( C1 => n297, C2 => n14034, A => n14033, B => 
                           n14153, ZN => n13751);
   U17424 : NOR2_X1 port map( A1 => n3889, A2 => n3888, ZN => n14947);
   U17425 : NAND2_X1 port map( A1 => n14947, A2 => n14946, ZN => n13755);
   U17426 : NOR2_X1 port map( A1 => n2570, A2 => n25458, ZN => n13753);
   U17427 : NOR2_X1 port map( A1 => n2684, A2 => n12629, ZN => n13752);
   U17428 : OAI21_X1 port map( B1 => n13753, B2 => n13752, A => n14198, ZN => 
                           n13754);
   U17429 : NAND3_X1 port map( A1 => n13755, A2 => n13754, A3 => n14949, ZN => 
                           n14383);
   U17430 : XNOR2_X1 port map( A => n15464, B => n14383, ZN => n14638);
   U17431 : XNOR2_X1 port map( A => n13756, B => n14638, ZN => n13784);
   U17432 : INV_X1 port map( A => n13757, ZN => n13758);
   U17433 : NOR3_X1 port map( A1 => n397, A2 => n13759, A3 => n13758, ZN => 
                           n13760);
   U17434 : NOR2_X1 port map( A1 => n13839, A2 => n13760, ZN => n13763);
   U17435 : INV_X1 port map( A => n13761, ZN => n13762);
   U17436 : NAND2_X1 port map( A1 => n13763, A2 => n13762, ZN => n13767);
   U17437 : NOR2_X1 port map( A1 => n14271, A2 => n14274, ZN => n13765);
   U17438 : AOI22_X1 port map( A1 => n13765, A2 => n24368, B1 => n13839, B2 => 
                           n13764, ZN => n13766);
   U17439 : NAND2_X1 port map( A1 => n13767, A2 => n13766, ZN => n14516);
   U17440 : NOR2_X1 port map( A1 => n14178, A2 => n14182, ZN => n13770);
   U17441 : NOR2_X1 port map( A1 => n13796, A2 => n13792, ZN => n13768);
   U17442 : AOI22_X1 port map( A1 => n13770, A2 => n13769, B1 => n13768, B2 => 
                           n14178, ZN => n13772);
   U17443 : XNOR2_X1 port map( A => n14775, B => n14516, ZN => n13782);
   U17444 : NAND2_X1 port map( A1 => n13775, A2 => n13954, ZN => n13779);
   U17445 : INV_X1 port map( A => n13776, ZN => n13777);
   U17446 : NAND2_X1 port map( A1 => n13777, A2 => n5080, ZN => n13778);
   U17447 : XNOR2_X1 port map( A => n25436, B => n1831, ZN => n13781);
   U17448 : XNOR2_X1 port map( A => n13782, B => n13781, ZN => n13783);
   U17449 : XNOR2_X1 port map( A => n13784, B => n13783, ZN => n16202);
   U17450 : INV_X1 port map( A => n16202, ZN => n16406);
   U17451 : NOR2_X1 port map( A1 => n13788, A2 => n14141, ZN => n13787);
   U17453 : NAND2_X1 port map( A1 => n13789, A2 => n13788, ZN => n13790);
   U17454 : NOR2_X1 port map( A1 => n14178, A2 => n24949, ZN => n13794);
   U17455 : MUX2_X1 port map( A => n13794, B => n13793, S => n13792, Z => 
                           n13799);
   U17456 : OAI22_X1 port map( A1 => n13797, A2 => n14179, B1 => n14182, B2 => 
                           n5755, ZN => n13798);
   U17457 : XNOR2_X1 port map( A => n15484, B => n1359, ZN => n13800);
   U17458 : XNOR2_X1 port map( A => n14979, B => n14678, ZN => n14534);
   U17459 : XNOR2_X1 port map( A => n13800, B => n14534, ZN => n13810);
   U17460 : XNOR2_X1 port map( A => n15386, B => n921, ZN => n13808);
   U17461 : NAND3_X1 port map( A1 => n14945, A2 => n14199, A3 => n25458, ZN => 
                           n13803);
   U17462 : XNOR2_X1 port map( A => n14977, B => n25013, ZN => n14608);
   U17463 : XNOR2_X1 port map( A => n13808, B => n14608, ZN => n13809);
   U17464 : XNOR2_X1 port map( A => n13810, B => n13809, ZN => n15638);
   U17465 : INV_X1 port map( A => n15638, ZN => n15973);
   U17466 : NOR2_X1 port map( A1 => n3341, A2 => n14205, ZN => n13812);
   U17467 : OAI21_X1 port map( B1 => n13813, B2 => n13812, A => n13811, ZN => 
                           n13817);
   U17468 : AOI21_X1 port map( B1 => n13815, B2 => n14209, A => n13814, ZN => 
                           n13816);
   U17469 : XNOR2_X1 port map( A => n14671, B => n15094, ZN => n13825);
   U17470 : NOR2_X1 port map( A1 => n13819, A2 => n13818, ZN => n13821);
   U17471 : OAI21_X1 port map( B1 => n13821, B2 => n13820, A => n13824, ZN => 
                           n13823);
   U17472 : OAI211_X1 port map( C1 => n13824, C2 => n13648, A => n13823, B => 
                           n13822, ZN => n14737);
   U17473 : XNOR2_X1 port map( A => n14737, B => n14654, ZN => n14986);
   U17474 : XNOR2_X1 port map( A => n14986, B => n13825, ZN => n13836);
   U17475 : NOR2_X1 port map( A1 => n13895, A2 => n1331, ZN => n13827);
   U17476 : XNOR2_X1 port map( A => n15507, B => n15183, ZN => n15368);
   U17477 : NOR2_X1 port map( A1 => n13830, A2 => n14219, ZN => n13828);
   U17478 : AND2_X1 port map( A1 => n13830, A2 => n14225, ZN => n14116);
   U17479 : NAND3_X1 port map( A1 => n14222, A2 => n13830, A3 => n14219, ZN => 
                           n13832);
   U17480 : OAI211_X2 port map( C1 => n13833, C2 => n14119, A => n13832, B => 
                           n13831, ZN => n15359);
   U17481 : XNOR2_X1 port map( A => n15359, B => n2033, ZN => n13834);
   U17482 : XNOR2_X1 port map( A => n15368, B => n13834, ZN => n13835);
   U17483 : INV_X1 port map( A => n16186, ZN => n16398);
   U17484 : NOR2_X1 port map( A1 => n15973, A2 => n16398, ZN => n13916);
   U17485 : NOR2_X1 port map( A1 => n13839, A2 => n14268, ZN => n13838);
   U17486 : AOI21_X1 port map( B1 => n13840, B2 => n13839, A => n13838, ZN => 
                           n13841);
   U17487 : MUX2_X1 port map( A => n13842, B => n13841, S => n14274, Z => 
                           n15002);
   U17488 : XNOR2_X1 port map( A => n1351, B => n15002, ZN => n13850);
   U17489 : NOR2_X1 port map( A1 => n13627, A2 => n14063, ZN => n13846);
   U17490 : NAND2_X1 port map( A1 => n14069, A2 => n13846, ZN => n13848);
   U17491 : AND2_X1 port map( A1 => n13847, A2 => n14063, ZN => n14065);
   U17493 : XNOR2_X1 port map( A => n14611, B => n15178, ZN => n14965);
   U17494 : XNOR2_X1 port map( A => n14965, B => n13850, ZN => n13862);
   U17495 : OAI21_X1 port map( B1 => n14075, B2 => n13852, A => n13851, ZN => 
                           n13857);
   U17496 : OAI21_X1 port map( B1 => n13854, B2 => n13853, A => n12704, ZN => 
                           n13856);
   U17497 : AOI21_X1 port map( B1 => n14074, B2 => n14079, A => n14078, ZN => 
                           n13855);
   U17498 : AOI21_X1 port map( B1 => n24572, B2 => n14849, A => n14852, ZN => 
                           n13858);
   U17499 : OAI21_X1 port map( B1 => n24572, B2 => n14416, A => n13858, ZN => 
                           n13859);
   U17500 : XNOR2_X1 port map( A => n24956, B => n14558, ZN => n14614);
   U17501 : XNOR2_X1 port map( A => n14690, B => n1856, ZN => n13860);
   U17502 : XNOR2_X1 port map( A => n14614, B => n13860, ZN => n13861);
   U17503 : XNOR2_X1 port map( A => n13862, B => n13861, ZN => n13940);
   U17504 : INV_X1 port map( A => n13940, ZN => n16188);
   U17505 : NOR2_X1 port map( A1 => n14325, A2 => n14328, ZN => n14043);
   U17506 : OAI21_X1 port map( B1 => n14043, B2 => n13864, A => n13863, ZN => 
                           n13866);
   U17507 : OAI21_X1 port map( B1 => n13864, B2 => n14324, A => n14328, ZN => 
                           n13865);
   U17508 : XNOR2_X1 port map( A => n13867, B => n14775, ZN => n13874);
   U17509 : OR2_X1 port map( A1 => n14319, A2 => n13868, ZN => n13870);
   U17510 : NAND3_X1 port map( A1 => n14321, A2 => n13868, A3 => n14320, ZN => 
                           n13869);
   U17511 : OAI21_X1 port map( B1 => n14317, B2 => n13870, A => n13869, ZN => 
                           n13872);
   U17512 : XNOR2_X1 port map( A => n15120, B => n13873, ZN => n14955);
   U17513 : XNOR2_X1 port map( A => n13874, B => n14955, ZN => n13887);
   U17514 : NAND2_X1 port map( A1 => n14340, A2 => n14335, ZN => n13876);
   U17515 : NAND2_X1 port map( A1 => n13877, A2 => n25197, ZN => n13875);
   U17516 : AOI21_X1 port map( B1 => n13876, B2 => n13875, A => n14333, ZN => 
                           n13882);
   U17517 : NOR2_X1 port map( A1 => n25196, A2 => n14339, ZN => n14028);
   U17518 : NAND2_X1 port map( A1 => n13878, A2 => n14336, ZN => n13879);
   U17519 : NAND2_X1 port map( A1 => n13880, A2 => n13879, ZN => n13881);
   U17520 : XNOR2_X1 port map( A => n25443, B => n15393, ZN => n14593);
   U17521 : XNOR2_X1 port map( A => n15019, B => n14593, ZN => n13886);
   U17522 : XNOR2_X1 port map( A => n13887, B => n13886, ZN => n15637);
   U17523 : INV_X1 port map( A => n15637, ZN => n16399);
   U17524 : NOR2_X1 port map( A1 => n16188, A2 => n16399, ZN => n13915);
   U17525 : OAI21_X1 port map( B1 => n13890, B2 => n3966, A => n1527, ZN => 
                           n13891);
   U17526 : NAND2_X1 port map( A1 => n13894, A2 => n4133, ZN => n13898);
   U17528 : XNOR2_X1 port map( A => n15326, B => n24423, ZN => n14619);
   U17529 : AOI21_X1 port map( B1 => n13901, B2 => n13900, A => n13903, ZN => 
                           n13905);
   U17531 : XNOR2_X1 port map( A => n14973, B => n14619, ZN => n13914);
   U17532 : XNOR2_X1 port map( A => n25413, B => n15229, ZN => n14543);
   U17533 : AOI21_X1 port map( B1 => n24974, B2 => n13907, A => n14293, ZN => 
                           n13911);
   U17534 : INV_X1 port map( A => n14294, ZN => n14291);
   U17535 : NOR2_X1 port map( A1 => n14294, A2 => n13909, ZN => n13948);
   U17536 : OAI21_X1 port map( B1 => n13911, B2 => n14291, A => n13910, ZN => 
                           n14719);
   U17537 : XNOR2_X1 port map( A => n14719, B => n2236, ZN => n13912);
   U17538 : XNOR2_X1 port map( A => n14543, B => n13912, ZN => n13913);
   U17539 : MUX2_X1 port map( A => n13916, B => n13915, S => n3630, Z => n13943
                           );
   U17540 : NAND2_X1 port map( A1 => n1846, A2 => n16186, ZN => n15639);
   U17541 : INV_X1 port map( A => n13985, ZN => n13920);
   U17542 : OAI21_X1 port map( B1 => n13918, B2 => n13922, A => n13917, ZN => 
                           n13919);
   U17543 : NOR2_X1 port map( A1 => n14008, A2 => n13923, ZN => n14255);
   U17544 : NOR2_X1 port map( A1 => n14252, A2 => n14251, ZN => n13926);
   U17545 : NAND2_X1 port map( A1 => n14254, A2 => n13924, ZN => n13925);
   U17546 : OAI22_X1 port map( A1 => n13927, A2 => n14255, B1 => n13926, B2 => 
                           n13925, ZN => n15515);
   U17547 : XNOR2_X1 port map( A => n15515, B => n15350, ZN => n14600);
   U17548 : XNOR2_X1 port map( A => n14600, B => n13928, ZN => n13939);
   U17549 : NOR2_X1 port map( A1 => n13995, A2 => n13997, ZN => n13930);
   U17550 : XNOR2_X1 port map( A => n15112, B => n14996, ZN => n13937);
   U17551 : NAND3_X1 port map( A1 => n13931, A2 => n13935, A3 => n14244, ZN => 
                           n13934);
   U17552 : NOR2_X1 port map( A1 => n25208, A2 => n14244, ZN => n13933);
   U17553 : XNOR2_X1 port map( A => n14997, B => n1746, ZN => n13936);
   U17554 : XNOR2_X1 port map( A => n13937, B => n13936, ZN => n13938);
   U17556 : AOI21_X1 port map( B1 => n15639, B2 => n13941, A => n15971, ZN => 
                           n13942);
   U17557 : AOI21_X1 port map( B1 => n24588, B2 => n24710, A => n14306, ZN => 
                           n13946);
   U17558 : INV_X1 port map( A => n13948, ZN => n13950);
   U17559 : NAND2_X1 port map( A1 => n13953, A2 => n14158, ZN => n13952);
   U17560 : XNOR2_X1 port map( A => n15111, B => n14579, ZN => n14429);
   U17561 : XNOR2_X1 port map( A => n14429, B => n14715, ZN => n13973);
   U17562 : NAND2_X1 port map( A1 => n13957, A2 => n13956, ZN => n13961);
   U17563 : OAI211_X1 port map( C1 => n14311, C2 => n14307, A => n13959, B => 
                           n13958, ZN => n13960);
   U17565 : XNOR2_X1 port map( A => n15109, B => n25008, ZN => n13971);
   U17566 : NAND3_X1 port map( A1 => n13968, A2 => n13966, A3 => n13965, ZN => 
                           n13967);
   U17567 : XNOR2_X1 port map( A => n15153, B => n1754, ZN => n13970);
   U17568 : XNOR2_X1 port map( A => n13971, B => n13970, ZN => n13972);
   U17573 : XNOR2_X1 port map( A => n15088, B => n15210, ZN => n14423);
   U17574 : INV_X1 port map( A => n14423, ZN => n13999);
   U17575 : NOR2_X1 port map( A1 => n13988, A2 => n13981, ZN => n13983);
   U17576 : NAND2_X1 port map( A1 => n13986, A2 => n13985, ZN => n13992);
   U17577 : XNOR2_X1 port map( A => n14788, B => n15483, ZN => n14532);
   U17578 : XNOR2_X1 port map( A => n13999, B => n14532, ZN => n14016);
   U17579 : AOI21_X1 port map( B1 => n299, B2 => n14000, A => n14003, ZN => 
                           n14001);
   U17580 : NOR2_X1 port map( A1 => n14009, A2 => n14251, ZN => n14010);
   U17581 : XNOR2_X1 port map( A => n14980, B => n24502, ZN => n14014);
   U17582 : XNOR2_X1 port map( A => n14792, B => n1924, ZN => n14013);
   U17583 : XNOR2_X1 port map( A => n14014, B => n14013, ZN => n14015);
   U17584 : XNOR2_X1 port map( A => n14015, B => n14016, ZN => n15640);
   U17585 : NAND2_X1 port map( A1 => n14022, A2 => n14085, ZN => n14092);
   U17586 : NOR2_X1 port map( A1 => n14018, A2 => n14022, ZN => n14019);
   U17587 : AOI21_X1 port map( B1 => n14020, B2 => n14092, A => n14019, ZN => 
                           n14024);
   U17588 : NOR3_X1 port map( A1 => n14022, A2 => n14089, A3 => n14021, ZN => 
                           n14023);
   U17589 : XNOR2_X1 port map( A => n15184, B => n15097, ZN => n14414);
   U17590 : AND2_X1 port map( A1 => n14025, A2 => n25197, ZN => n14027);
   U17591 : OAI21_X1 port map( B1 => n14337, B2 => n14027, A => n14026, ZN => 
                           n14030);
   U17592 : NAND2_X1 port map( A1 => n14028, A2 => n14336, ZN => n14029);
   U17593 : NAND2_X1 port map( A1 => n14033, A2 => n14032, ZN => n14037);
   U17594 : NOR2_X1 port map( A1 => n14150, A2 => n14034, ZN => n14036);
   U17595 : XNOR2_X1 port map( A => n15506, B => n14846, ZN => n15150);
   U17596 : NOR2_X1 port map( A1 => n14321, A2 => n3401, ZN => n14038);
   U17597 : NOR2_X1 port map( A1 => n14319, A2 => n14458, ZN => n14039);
   U17598 : OAI21_X1 port map( B1 => n14039, B2 => n14320, A => n14321, ZN => 
                           n14040);
   U17599 : NOR2_X1 port map( A1 => n14330, A2 => n14041, ZN => n14042);
   U17600 : XNOR2_X1 port map( A => n15095, B => n15298, ZN => n14046);
   U17601 : XNOR2_X1 port map( A => n14800, B => n19392, ZN => n14045);
   U17602 : XNOR2_X1 port map( A => n14046, B => n14045, ZN => n14047);
   U17603 : NAND2_X1 port map( A1 => n14050, A2 => n14049, ZN => n14051);
   U17604 : NAND2_X1 port map( A1 => n14053, A2 => n14051, ZN => n14057);
   U17605 : NOR2_X1 port map( A1 => n14052, A2 => n14054, ZN => n14056);
   U17606 : XNOR2_X1 port map( A => n15119, B => n641, ZN => n14061);
   U17607 : XNOR2_X1 port map( A => n14061, B => n15133, ZN => n14084);
   U17608 : INV_X1 port map( A => n14069, ZN => n14062);
   U17609 : NOR2_X1 port map( A1 => n14062, A2 => n14063, ZN => n14072);
   U17610 : NAND2_X1 port map( A1 => n14064, A2 => n14063, ZN => n14264);
   U17611 : INV_X1 port map( A => n14065, ZN => n14066);
   U17613 : AOI21_X1 port map( B1 => n13627, B2 => n14067, A => n300, ZN => 
                           n14068);
   U17614 : NAND2_X1 port map( A1 => n14069, A2 => n14068, ZN => n14070);
   U17616 : NAND2_X1 port map( A1 => n14074, A2 => n14073, ZN => n14082);
   U17618 : XNOR2_X1 port map( A => n15497, B => n15274, ZN => n14725);
   U17619 : XNOR2_X1 port map( A => n14084, B => n14725, ZN => n14095);
   U17620 : XNOR2_X1 port map( A => n14553, B => n14516, ZN => n14093);
   U17621 : INV_X1 port map( A => n14085, ZN => n14086);
   U17622 : NAND2_X1 port map( A1 => n14092, A2 => n14087, ZN => n14091);
   U17623 : XNOR2_X1 port map( A => n14093, B => n15321, ZN => n14094);
   U17624 : NAND2_X1 port map( A1 => n4892, A2 => n25445, ZN => n14097);
   U17625 : NOR2_X1 port map( A1 => n14101, A2 => n24376, ZN => n14102);
   U17626 : MUX2_X1 port map( A => n14107, B => n14106, S => n14105, Z => 
                           n14114);
   U17627 : NOR2_X1 port map( A1 => n14109, A2 => n14108, ZN => n14110);
   U17628 : NOR2_X1 port map( A1 => n14111, A2 => n14110, ZN => n14113);
   U17629 : XNOR2_X1 port map( A => n15082, B => n15401, ZN => n14403);
   U17630 : XNOR2_X1 port map( A => n14403, B => n14115, ZN => n14137);
   U17631 : INV_X1 port map( A => n14116, ZN => n14117);
   U17632 : NAND2_X1 port map( A1 => n14118, A2 => n14117, ZN => n14120);
   U17633 : XNOR2_X1 port map( A => n15284, B => n15480, ZN => n14731);
   U17636 : AND2_X1 port map( A1 => n14130, A2 => n1331, ZN => n14131);
   U17637 : XNOR2_X1 port map( A => n15415, B => n4164, ZN => n14135);
   U17638 : XNOR2_X1 port map( A => n14731, B => n14135, ZN => n14136);
   U17639 : XNOR2_X1 port map( A => n14137, B => n14136, ZN => n15905);
   U17640 : NOR2_X1 port map( A1 => n16368, A2 => n15905, ZN => n15641);
   U17641 : INV_X1 port map( A => n15641, ZN => n14139);
   U17642 : NAND2_X1 port map( A1 => n14139, A2 => n14138, ZN => n14176);
   U17643 : XNOR2_X1 port map( A => n14858, B => n3131, ZN => n14155);
   U17644 : NAND2_X1 port map( A1 => n14200, A2 => n3888, ZN => n14148);
   U17645 : OAI21_X1 port map( B1 => n14945, B2 => n14944, A => n2684, ZN => 
                           n14146);
   U17646 : XNOR2_X1 port map( A => n15526, B => n15055, ZN => n14541);
   U17647 : XNOR2_X1 port map( A => n14155, B => n14541, ZN => n14175);
   U17648 : NAND2_X1 port map( A1 => n14159, A2 => n14158, ZN => n14161);
   U17649 : NAND2_X1 port map( A1 => n14161, A2 => n14160, ZN => n14162);
   U17650 : NAND2_X1 port map( A1 => n14163, A2 => n14162, ZN => n14897);
   U17651 : NAND3_X1 port map( A1 => n14169, A2 => n14168, A3 => n14167, ZN => 
                           n14170);
   U17652 : XNOR2_X1 port map( A => n14809, B => n14897, ZN => n15102);
   U17653 : XNOR2_X1 port map( A => n14806, B => n15169, ZN => n14173);
   U17654 : XNOR2_X1 port map( A => n14173, B => n15102, ZN => n14174);
   U17655 : XNOR2_X1 port map( A => n14892, B => n15002, ZN => n14373);
   U17656 : MUX2_X1 port map( A => n24949, B => n14179, S => n14178, Z => 
                           n14184);
   U17657 : XNOR2_X1 port map( A => n14185, B => n14642, ZN => n14186);
   U17658 : NAND2_X1 port map( A1 => n25560, A2 => n25360, ZN => n14192);
   U17660 : NOR2_X1 port map( A1 => n25560, A2 => n14194, ZN => n14196);
   U17661 : NAND2_X1 port map( A1 => n14201, A2 => n14200, ZN => n14203);
   U17662 : OAI21_X1 port map( B1 => n14206, B2 => n14205, A => n14204, ZN => 
                           n14207);
   U17663 : AOI22_X2 port map( A1 => n14210, A2 => n14209, B1 => n14207, B2 => 
                           n2378, ZN => n15409);
   U17664 : XNOR2_X1 port map( A => n15409, B => n14377, ZN => n14972);
   U17665 : OAI21_X1 port map( B1 => n24503, B2 => n13417, A => n14211, ZN => 
                           n14214);
   U17666 : NAND2_X1 port map( A1 => n14214, A2 => n14213, ZN => n14215);
   U17667 : OAI21_X1 port map( B1 => n14217, B2 => n14216, A => n14215, ZN => 
                           n15164);
   U17668 : XNOR2_X1 port map( A => n15164, B => n15054, ZN => n14860);
   U17669 : XNOR2_X1 port map( A => n14860, B => n14972, ZN => n14229);
   U17670 : XNOR2_X1 port map( A => n14719, B => n3073, ZN => n14227);
   U17671 : OAI21_X1 port map( B1 => n14219, B2 => n14218, A => n14221, ZN => 
                           n14220);
   U17672 : NAND3_X1 port map( A1 => n14223, A2 => n14222, A3 => n14221, ZN => 
                           n14224);
   U17673 : XNOR2_X1 port map( A => n14694, B => n25384, ZN => n14896);
   U17674 : XNOR2_X1 port map( A => n14896, B => n14227, ZN => n14228);
   U17675 : XNOR2_X1 port map( A => n14845, B => n15369, ZN => n14239);
   U17676 : XNOR2_X1 port map( A => n14911, B => n14239, ZN => n14263);
   U17677 : NAND3_X1 port map( A1 => n14241, A2 => n14245, A3 => n14240, ZN => 
                           n14248);
   U17678 : NAND3_X1 port map( A1 => n14245, A2 => n13633, A3 => n14244, ZN => 
                           n14246);
   U17679 : XNOR2_X1 port map( A => n14907, B => n2039, ZN => n14249);
   U17680 : XNOR2_X1 port map( A => n14737, B => n14249, ZN => n14261);
   U17682 : OR2_X1 port map( A1 => n14254, A2 => n14253, ZN => n14258);
   U17683 : NAND2_X1 port map( A1 => n14256, A2 => n14255, ZN => n14257);
   U17684 : XNOR2_X1 port map( A => n14958, B => n15505, ZN => n15366);
   U17685 : XNOR2_X1 port map( A => n14261, B => n15366, ZN => n14262);
   U17686 : XNOR2_X1 port map( A => n295, B => n14900, ZN => n14354);
   U17687 : XNOR2_X1 port map( A => n15033, B => n15375, ZN => n14266);
   U17688 : XNOR2_X1 port map( A => n14354, B => n14266, ZN => n14286);
   U17689 : OAI21_X1 port map( B1 => n14268, B2 => n14267, A => n397, ZN => 
                           n14273);
   U17690 : NAND2_X1 port map( A1 => n14274, A2 => n14269, ZN => n14270);
   U17692 : NOR2_X2 port map( A1 => n14277, A2 => n14276, ZN => n14902);
   U17693 : XNOR2_X1 port map( A => n14902, B => n15514, ZN => n14284);
   U17694 : NOR2_X1 port map( A1 => n14850, A2 => n14278, ZN => n14279);
   U17695 : OAI21_X1 port map( B1 => n14849, B2 => n14852, A => n14279, ZN => 
                           n14282);
   U17696 : NAND2_X1 port map( A1 => n14280, A2 => n14415, ZN => n14281);
   U17697 : OAI211_X1 port map( C1 => n24572, C2 => n14415, A => n14281, B => 
                           n14282, ZN => n15378);
   U17698 : XNOR2_X1 port map( A => n15378, B => n4189, ZN => n14283);
   U17699 : XNOR2_X1 port map( A => n14284, B => n14283, ZN => n14285);
   U17700 : XNOR2_X1 port map( A => n14285, B => n14286, ZN => n14350);
   U17701 : INV_X1 port map( A => n14350, ZN => n16382);
   U17702 : OAI21_X1 port map( B1 => n15656, B2 => n25210, A => n15990, ZN => 
                           n14352);
   U17703 : XNOR2_X1 port map( A => n14724, B => n494, ZN => n14288);
   U17704 : XNOR2_X1 port map( A => n14288, B => n14287, ZN => n14316);
   U17705 : OAI21_X1 port map( B1 => n394, B2 => n14290, A => n14289, ZN => 
                           n14297);
   U17707 : NAND3_X1 port map( A1 => n14294, A2 => n14293, A3 => n14292, ZN => 
                           n14295);
   U17708 : XNOR2_X1 port map( A => n14634, B => n15396, ZN => n15495);
   U17709 : NOR2_X1 port map( A1 => n14302, A2 => n1527, ZN => n14300);
   U17710 : NOR2_X1 port map( A1 => n14301, A2 => n13888, ZN => n14299);
   U17711 : AOI22_X1 port map( A1 => n14300, A2 => n13728, B1 => n14299, B2 => 
                           n1527, ZN => n14305);
   U17712 : NAND2_X1 port map( A1 => n14302, A2 => n14301, ZN => n14303);
   U17713 : INV_X1 port map( A => n14307, ZN => n14315);
   U17714 : OAI21_X1 port map( B1 => n14310, B2 => n14309, A => n14308, ZN => 
                           n14313);
   U17715 : OAI211_X1 port map( C1 => n14315, C2 => n14314, A => n14313, B => 
                           n14312, ZN => n15204);
   U17716 : XNOR2_X1 port map( A => n15204, B => n15275, ZN => n15398);
   U17717 : NOR2_X1 port map( A1 => n14321, A2 => n14320, ZN => n14322);
   U17718 : XNOR2_X1 port map( A => n15238, B => n14982, ZN => n14332);
   U17719 : MUX2_X1 port map( A => n14325, B => n14327, S => n14324, Z => 
                           n14326);
   U17721 : XNOR2_X1 port map( A => n14332, B => n14331, ZN => n14349);
   U17722 : OAI21_X1 port map( B1 => n14335, B2 => n14334, A => n14333, ZN => 
                           n14343);
   U17723 : NAND2_X1 port map( A1 => n14337, A2 => n14336, ZN => n14342);
   U17724 : NAND3_X1 port map( A1 => n14340, A2 => n14339, A3 => n25197, ZN => 
                           n14341);
   U17725 : OAI211_X2 port map( C1 => n14344, C2 => n14343, A => n14342, B => 
                           n14341, ZN => n15387);
   U17726 : XNOR2_X1 port map( A => n14345, B => n15387, ZN => n14347);
   U17727 : XNOR2_X1 port map( A => n15488, B => n449, ZN => n14346);
   U17728 : XNOR2_X1 port map( A => n14347, B => n14346, ZN => n14348);
   U17729 : XNOR2_X1 port map( A => n14348, B => n14349, ZN => n15657);
   U17731 : OAI21_X1 port map( B1 => n16383, B2 => n16177, A => n15837, ZN => 
                           n14351);
   U17732 : INV_X1 port map( A => n14354, ZN => n14356);
   U17733 : XNOR2_X1 port map( A => n24975, B => n62, ZN => n14355);
   U17734 : XOR2_X1 port map( A => n14356, B => n14355, Z => n14358);
   U17735 : XNOR2_X1 port map( A => n15515, B => n15444, ZN => n15113);
   U17736 : XNOR2_X1 port map( A => n15113, B => n15513, ZN => n14357);
   U17737 : NAND2_X1 port map( A1 => n14359, A2 => n3701, ZN => n14367);
   U17738 : NOR2_X1 port map( A1 => n24995, A2 => n3701, ZN => n14365);
   U17739 : XNOR2_X1 port map( A => n14368, B => n15487, ZN => n14920);
   U17740 : XNOR2_X1 port map( A => n15486, B => n2193, ZN => n14369);
   U17741 : XNOR2_X1 port map( A => n14920, B => n14369, ZN => n14372);
   U17742 : XNOR2_X1 port map( A => n15436, B => n15484, ZN => n15087);
   U17743 : XNOR2_X1 port map( A => n15087, B => n14370, ZN => n14371);
   U17744 : XNOR2_X1 port map( A => n24956, B => n14644, ZN => n14780);
   U17745 : XNOR2_X1 port map( A => n14780, B => n14373, ZN => n14376);
   U17746 : XNOR2_X1 port map( A => n15284, B => n2881, ZN => n14374);
   U17747 : XNOR2_X1 port map( A => n14375, B => n14376, ZN => n16156);
   U17748 : INV_X1 port map( A => n16156, ZN => n16154);
   U17749 : XNOR2_X1 port map( A => n25431, B => n14719, ZN => n15012);
   U17750 : XNOR2_X1 port map( A => n15012, B => n15106, ZN => n14380);
   U17751 : XNOR2_X1 port map( A => n15055, B => n23883, ZN => n14378);
   U17752 : XNOR2_X1 port map( A => n14898, B => n14378, ZN => n14379);
   U17753 : NAND2_X1 port map( A1 => n16122, A2 => n15842, ZN => n14381);
   U17755 : NAND2_X1 port map( A1 => n16156, A2 => n25449, ZN => n15619);
   U17756 : INV_X1 port map( A => n15619, ZN => n14388);
   U17757 : XNOR2_X1 port map( A => n14724, B => n14383, ZN => n15016);
   U17758 : XNOR2_X1 port map( A => n15393, B => n15464, ZN => n15123);
   U17759 : XNOR2_X1 port map( A => n15274, B => n1768, ZN => n14385);
   U17760 : XNOR2_X1 port map( A => n15123, B => n14385, ZN => n14386);
   U17761 : XNOR2_X1 port map( A => n14387, B => n14386, ZN => n16123);
   U17762 : INV_X1 port map( A => n16123, ZN => n16155);
   U17763 : NAND2_X1 port map( A1 => n14388, A2 => n16155, ZN => n14395);
   U17764 : XNOR2_X1 port map( A => n15298, B => n21742, ZN => n14390);
   U17765 : XNOR2_X1 port map( A => n15504, B => n14390, ZN => n14393);
   U17766 : INV_X1 port map( A => n15507, ZN => n14391);
   U17767 : XNOR2_X1 port map( A => n14392, B => n14393, ZN => n16125);
   U17768 : NAND3_X1 port map( A1 => n24459, A2 => n381, A3 => n16122, ZN => 
                           n14394);
   U17769 : INV_X1 port map( A => n14398, ZN => n23602);
   U17770 : OAI21_X1 port map( B1 => n5487, B2 => n14397, A => n23602, ZN => 
                           n14400);
   U17771 : NAND3_X1 port map( A1 => n5486, A2 => n14398, A3 => n2556, ZN => 
                           n14399);
   U17772 : NAND2_X1 port map( A1 => n14400, A2 => n14399, ZN => n14401);
   U17773 : XNOR2_X1 port map( A => n14402, B => n14401, ZN => n14404);
   U17774 : XNOR2_X1 port map( A => n14880, B => n14642, ZN => n14891);
   U17775 : INV_X1 port map( A => n16170, ZN => n16424);
   U17776 : XNOR2_X1 port map( A => n14634, B => n15200, ZN => n14406);
   U17777 : XNOR2_X1 port map( A => n15119, B => n3125, ZN => n14405);
   U17778 : XNOR2_X1 port map( A => n14406, B => n14405, ZN => n14408);
   U17779 : XNOR2_X1 port map( A => n15273, B => n14591, ZN => n15201);
   U17780 : XNOR2_X1 port map( A => n15201, B => n15270, ZN => n14407);
   U17781 : XNOR2_X1 port map( A => n14408, B => n14407, ZN => n16426);
   U17782 : INV_X1 port map( A => n16426, ZN => n16169);
   U17783 : XNOR2_X1 port map( A => n15170, B => n15268, ZN => n14412);
   U17784 : INV_X1 port map( A => n15522, ZN => n14409);
   U17785 : XNOR2_X1 port map( A => n14409, B => n15169, ZN => n14562);
   U17786 : XNOR2_X1 port map( A => n14809, B => n2137, ZN => n14410);
   U17787 : XNOR2_X1 port map( A => n14562, B => n14410, ZN => n14411);
   U17788 : NAND2_X1 port map( A1 => n16169, A2 => n15958, ZN => n14433);
   U17789 : INV_X1 port map( A => n20284, ZN => n23523);
   U17790 : AOI21_X1 port map( B1 => n14849, B2 => n14416, A => n14415, ZN => 
                           n14417);
   U17791 : OAI21_X1 port map( B1 => n24572, B2 => n14849, A => n14417, ZN => 
                           n14418);
   U17792 : NAND2_X1 port map( A1 => n14419, A2 => n14418, ZN => n14420);
   U17793 : XNOR2_X1 port map( A => n14799, B => n14420, ZN => n15299);
   U17794 : XNOR2_X1 port map( A => n15188, B => n15299, ZN => n14421);
   U17795 : OAI21_X1 port map( B1 => n16169, B2 => n244, A => n16427, ZN => 
                           n14427);
   U17796 : XNOR2_X1 port map( A => n14928, B => n14468, ZN => n15208);
   U17797 : XNOR2_X1 port map( A => n15290, B => n15208, ZN => n14426);
   U17798 : XNOR2_X1 port map( A => n14919, B => n2795, ZN => n14424);
   U17799 : XNOR2_X1 port map( A => n14423, B => n14424, ZN => n14425);
   U17800 : NAND2_X1 port map( A1 => n14427, A2 => n1329, ZN => n14432);
   U17801 : XNOR2_X1 port map( A => n15190, B => n859, ZN => n14428);
   U17802 : INV_X1 port map( A => n16422, ZN => n15961);
   U17803 : NAND3_X1 port map( A1 => n15961, A2 => n707, A3 => n16169, ZN => 
                           n14431);
   U17804 : NOR2_X1 port map( A1 => n17283, A2 => n17229, ZN => n16952);
   U17805 : INV_X1 port map( A => n14434, ZN => n14438);
   U17806 : NOR2_X1 port map( A1 => n14438, A2 => n14437, ZN => n14441);
   U17808 : XNOR2_X1 port map( A => n15223, B => n14816, ZN => n14443);
   U17809 : XNOR2_X1 port map( A => n14442, B => n15415, ZN => n14729);
   U17810 : XNOR2_X1 port map( A => n15177, B => n15416, ZN => n14444);
   U17811 : XNOR2_X1 port map( A => n15230, B => n14806, ZN => n14446);
   U17812 : XNOR2_X1 port map( A => n15168, B => n15056, ZN => n14445);
   U17813 : XNOR2_X1 port map( A => n14446, B => n14445, ZN => n14450);
   U17814 : XNOR2_X1 port map( A => n14620, B => n14858, ZN => n14448);
   U17815 : XNOR2_X1 port map( A => n14857, B => n2049, ZN => n14447);
   U17816 : XNOR2_X1 port map( A => n14448, B => n14447, ZN => n14449);
   U17817 : XNOR2_X1 port map( A => n14450, B => n14449, ZN => n16408);
   U17818 : XNOR2_X1 port map( A => n14800, B => n21662, ZN => n14451);
   U17819 : XNOR2_X1 port map( A => n15253, B => n14669, ZN => n14452);
   U17820 : XNOR2_X1 port map( A => n14988, B => n14846, ZN => n14739);
   U17821 : XNOR2_X1 port map( A => n14739, B => n15358, ZN => n15456);
   U17822 : XNOR2_X1 port map( A => n15456, B => n14453, ZN => n16414);
   U17823 : INV_X1 port map( A => n16414, ZN => n16140);
   U17824 : XNOR2_X1 port map( A => n15244, B => n24287, ZN => n14454);
   U17825 : XNOR2_X1 port map( A => n25008, B => n15190, ZN => n14455);
   U17826 : XNOR2_X1 port map( A => n14456, B => n14455, ZN => n14465);
   U17827 : INV_X1 port map( A => n14457, ZN => n14462);
   U17828 : AND2_X1 port map( A1 => n14458, A2 => n14459, ZN => n14461);
   U17829 : XNOR2_X1 port map( A => n15153, B => n14463, ZN => n14464);
   U17830 : XNOR2_X1 port map( A => n15347, B => n14464, ZN => n15449);
   U17831 : XNOR2_X2 port map( A => n14465, B => n15449, ZN => n16412);
   U17832 : NAND2_X1 port map( A1 => n16140, A2 => n16412, ZN => n15653);
   U17833 : INV_X1 port map( A => n16408, ZN => n16416);
   U17834 : XNOR2_X1 port map( A => n15138, B => n14976, ZN => n14467);
   U17835 : XNOR2_X1 port map( A => n14467, B => n14466, ZN => n15441);
   U17836 : XNOR2_X1 port map( A => n14755, B => n14792, ZN => n14470);
   U17837 : XNOR2_X1 port map( A => n14468, B => n836, ZN => n14469);
   U17838 : XNOR2_X1 port map( A => n15441, B => n14471, ZN => n15986);
   U17839 : INV_X1 port map( A => n15986, ZN => n16409);
   U17840 : INV_X1 port map( A => n16412, ZN => n14472);
   U17841 : XNOR2_X1 port map( A => n15203, B => n14516, ZN => n14831);
   U17842 : XNOR2_X1 port map( A => n15462, B => n14831, ZN => n14476);
   U17843 : XNOR2_X1 port map( A => n14703, B => n15219, ZN => n14474);
   U17844 : XNOR2_X1 port map( A => n24418, B => n1874, ZN => n14473);
   U17845 : XNOR2_X1 port map( A => n14474, B => n14473, ZN => n14475);
   U17846 : XNOR2_X1 port map( A => n14476, B => n14475, ZN => n16417);
   U17847 : INV_X1 port map( A => n16417, ZN => n15868);
   U17848 : XNOR2_X1 port map( A => n15238, B => n15488, ZN => n15385);
   U17849 : XNOR2_X1 port map( A => n14865, B => n14792, ZN => n15293);
   U17850 : XNOR2_X1 port map( A => n15385, B => n15293, ZN => n14481);
   U17851 : XNOR2_X1 port map( A => n14977, B => n14477, ZN => n14479);
   U17852 : XNOR2_X1 port map( A => n14468, B => n673, ZN => n14478);
   U17853 : XNOR2_X1 port map( A => n14479, B => n14478, ZN => n14480);
   U17854 : XNOR2_X1 port map( A => n15359, B => n3164, ZN => n14482);
   U17855 : XNOR2_X1 port map( A => n14482, B => n15369, ZN => n14483);
   U17856 : XNOR2_X1 port map( A => n14483, B => n14909, ZN => n14486);
   U17857 : INV_X1 port map( A => n14800, ZN => n14484);
   U17858 : XNOR2_X1 port map( A => n14484, B => n14845, ZN => n15297);
   U17859 : XNOR2_X1 port map( A => n15297, B => n15188, ZN => n14485);
   U17860 : XNOR2_X1 port map( A => n15514, B => n4233, ZN => n14487);
   U17861 : XNOR2_X1 port map( A => n14487, B => n15375, ZN => n14492);
   U17862 : INV_X1 port map( A => n15033, ZN => n14489);
   U17863 : XNOR2_X1 port map( A => n14488, B => n14489, ZN => n15303);
   U17864 : XNOR2_X1 port map( A => n15280, B => n14494, ZN => n14498);
   U17865 : XNOR2_X1 port map( A => n15476, B => n15417, ZN => n14496);
   U17866 : INV_X1 port map( A => n14558, ZN => n15333);
   U17867 : XNOR2_X1 port map( A => n15333, B => n1869, ZN => n14495);
   U17868 : XNOR2_X1 port map( A => n14495, B => n14496, ZN => n14497);
   U17869 : XNOR2_X1 port map( A => n14498, B => n14497, ZN => n14499);
   U17870 : OAI21_X1 port map( B1 => n15856, B2 => n15611, A => n16118, ZN => 
                           n14522);
   U17871 : INV_X1 port map( A => n14499, ZN => n16113);
   U17873 : XNOR2_X1 port map( A => n14694, B => n2765, ZN => n15407);
   U17874 : XNOR2_X1 port map( A => n15407, B => n15267, ZN => n14504);
   U17875 : XNOR2_X1 port map( A => n15431, B => n14620, ZN => n14502);
   U17876 : XNOR2_X1 port map( A => n15326, B => n3178, ZN => n14501);
   U17877 : XNOR2_X1 port map( A => n14502, B => n14501, ZN => n14503);
   U17878 : NAND2_X1 port map( A1 => n16113, A2 => n15857, ZN => n16680);
   U17879 : OAI21_X1 port map( B1 => n16117, B2 => n15856, A => n16680, ZN => 
                           n14521);
   U17880 : INV_X1 port map( A => n15204, ZN => n14505);
   U17881 : XNOR2_X1 port map( A => n15463, B => n14505, ZN => n14873);
   U17882 : MUX2_X1 port map( A => n14512, B => n14511, S => n14510, Z => 
                           n14515);
   U17883 : INV_X1 port map( A => n14513, ZN => n14514);
   U17884 : XNOR2_X1 port map( A => n15063, B => n14516, ZN => n15271);
   U17885 : XNOR2_X1 port map( A => n15271, B => n14873, ZN => n14520);
   U17886 : XNOR2_X1 port map( A => n25443, B => n14591, ZN => n14518);
   U17887 : XNOR2_X1 port map( A => n15396, B => n1815, ZN => n14517);
   U17888 : XNOR2_X1 port map( A => n14518, B => n14517, ZN => n14519);
   U17891 : OR2_X1 port map( A1 => n16952, A2 => n16753, ZN => n14590);
   U17892 : XNOR2_X1 port map( A => n15318, B => n15274, ZN => n14833);
   U17893 : XNOR2_X1 port map( A => n14775, B => n923, ZN => n14523);
   U17894 : XNOR2_X1 port map( A => n14523, B => n15321, ZN => n14524);
   U17895 : XNOR2_X1 port map( A => n14524, B => n14833, ZN => n14527);
   U17896 : XNOR2_X1 port map( A => n14703, B => n15497, ZN => n14525);
   U17897 : XNOR2_X1 port map( A => n14525, B => n15499, ZN => n14526);
   U17898 : INV_X1 port map( A => n16389, ZN => n15848);
   U17899 : XNOR2_X1 port map( A => n14731, B => n15332, ZN => n14531);
   U17900 : XNOR2_X1 port map( A => n14690, B => n1351, ZN => n14529);
   U17901 : XNOR2_X1 port map( A => n14529, B => n14528, ZN => n14530);
   U17902 : XNOR2_X1 port map( A => n15338, B => n14532, ZN => n14536);
   U17903 : XNOR2_X1 port map( A => n14675, B => n1801, ZN => n14533);
   U17904 : XNOR2_X1 port map( A => n14533, B => n14534, ZN => n14535);
   U17905 : XNOR2_X1 port map( A => n15506, B => n15298, ZN => n14738);
   U17906 : XNOR2_X1 port map( A => n15074, B => n15095, ZN => n15355);
   U17907 : XNOR2_X1 port map( A => n14738, B => n15355, ZN => n14540);
   U17908 : XNOR2_X1 port map( A => n14671, B => n14669, ZN => n14538);
   U17909 : XNOR2_X1 port map( A => n14654, B => n860, ZN => n14537);
   U17910 : XNOR2_X1 port map( A => n14538, B => n14537, ZN => n14539);
   U17912 : INV_X1 port map( A => n15980, ZN => n14546);
   U17913 : INV_X1 port map( A => n14897, ZN => n14629);
   U17914 : XNOR2_X1 port map( A => n14629, B => n15051, ZN => n15324);
   U17915 : XNOR2_X1 port map( A => n15324, B => n14541, ZN => n14545);
   U17916 : XNOR2_X1 port map( A => n14857, B => n23679, ZN => n14542);
   U17917 : XNOR2_X1 port map( A => n14543, B => n14542, ZN => n14544);
   U17918 : XNOR2_X1 port map( A => n14545, B => n14544, ZN => n16388);
   U17919 : INV_X1 port map( A => n14715, ZN => n14548);
   U17920 : XNOR2_X1 port map( A => n14548, B => n14547, ZN => n14552);
   U17921 : XNOR2_X1 port map( A => n15034, B => n15109, ZN => n15348);
   U17922 : XNOR2_X1 port map( A => n14549, B => n2050, ZN => n14550);
   U17923 : XNOR2_X1 port map( A => n15348, B => n14550, ZN => n14551);
   U17924 : INV_X1 port map( A => n16393, ZN => n16163);
   U17925 : XNOR2_X1 port map( A => n15464, B => n1767, ZN => n14554);
   U17926 : XNOR2_X1 port map( A => n14553, B => n14554, ZN => n14555);
   U17927 : XNOR2_X1 port map( A => n14556, B => n25426, ZN => n15218);
   U17928 : INV_X1 port map( A => n16151, ZN => n14747);
   U17929 : INV_X1 port map( A => n14644, ZN => n15421);
   U17930 : XNOR2_X1 port map( A => n14642, B => n15421, ZN => n14557);
   U17931 : XNOR2_X1 port map( A => n14557, B => n14965, ZN => n14561);
   U17932 : XNOR2_X1 port map( A => n15282, B => n14558, ZN => n15225);
   U17933 : XNOR2_X1 port map( A => n15401, B => n2240, ZN => n14559);
   U17934 : XNOR2_X1 port map( A => n15225, B => n14559, ZN => n14560);
   U17935 : INV_X1 port map( A => n14562, ZN => n14564);
   U17936 : XNOR2_X1 port map( A => n15430, B => n3190, ZN => n14563);
   U17937 : XNOR2_X1 port map( A => n14564, B => n14563, ZN => n14567);
   U17938 : INV_X1 port map( A => n15409, ZN => n14565);
   U17939 : XNOR2_X1 port map( A => n14565, B => n15326, ZN => n15010);
   U17940 : XNOR2_X1 port map( A => n14973, B => n15010, ZN => n14566);
   U17941 : NAND2_X1 port map( A1 => n293, A2 => n1762, ZN => n14586);
   U17942 : INV_X1 port map( A => n14919, ZN => n14568);
   U17943 : XNOR2_X1 port map( A => n14977, B => n14568, ZN => n14569);
   U17944 : INV_X1 port map( A => n14922, ZN => n14868);
   U17945 : XNOR2_X1 port map( A => n14868, B => n15386, ZN => n14929);
   U17946 : XNOR2_X1 port map( A => n14929, B => n14569, ZN => n14573);
   U17947 : XNOR2_X1 port map( A => n15387, B => n15210, ZN => n14571);
   U17948 : XNOR2_X1 port map( A => n15436, B => n3133, ZN => n14570);
   U17949 : XNOR2_X1 port map( A => n14571, B => n14570, ZN => n14572);
   U17950 : XNOR2_X1 port map( A => n15094, B => n15183, ZN => n14961);
   U17951 : XNOR2_X1 port map( A => n15184, B => n15452, ZN => n14574);
   U17952 : XNOR2_X1 port map( A => n14961, B => n14574, ZN => n14577);
   U17953 : XNOR2_X1 port map( A => n14958, B => n15359, ZN => n15252);
   U17954 : XNOR2_X1 port map( A => n14907, B => n1891, ZN => n14575);
   U17955 : XNOR2_X1 port map( A => n15252, B => n14575, ZN => n14576);
   U17958 : XNOR2_X1 port map( A => n15378, B => n15350, ZN => n15246);
   U17959 : XNOR2_X1 port map( A => n14902, B => n15444, ZN => n14581);
   U17960 : XNOR2_X1 port map( A => n14579, B => n2126, ZN => n14580);
   U17961 : XNOR2_X1 port map( A => n14581, B => n14580, ZN => n14582);
   U17962 : NOR2_X1 port map( A1 => n16096, A2 => n16147, ZN => n14584);
   U17964 : INV_X1 port map( A => n17283, ZN => n17289);
   U17965 : NAND3_X1 port map( A1 => n17289, A2 => n17284, A3 => n17229, ZN => 
                           n14587);
   U17966 : NAND4_X1 port map( A1 => n14590, A2 => n14589, A3 => n14588, A4 => 
                           n14587, ZN => n17653);
   U17967 : XNOR2_X1 port map( A => n17653, B => n18146, ZN => n18323);
   U17968 : XNOR2_X1 port map( A => n15318, B => n24418, ZN => n14592);
   U17969 : INV_X1 port map( A => n14594, ZN => n15187);
   U17970 : XNOR2_X1 port map( A => n15094, B => n15187, ZN => n14912);
   U17971 : INV_X1 port map( A => n14912, ZN => n14598);
   U17972 : XNOR2_X1 port map( A => n15507, B => n15074, ZN => n14596);
   U17973 : XNOR2_X1 port map( A => n15359, B => n2882, ZN => n14595);
   U17974 : XNOR2_X1 port map( A => n14596, B => n14595, ZN => n14597);
   U17975 : XNOR2_X1 port map( A => n14600, B => n14940, ZN => n14604);
   U17976 : XNOR2_X1 port map( A => n15112, B => n15194, ZN => n14602);
   U17977 : XNOR2_X1 port map( A => n15034, B => n1789, ZN => n14601);
   U17978 : XNOR2_X1 port map( A => n14602, B => n14601, ZN => n14603);
   U17979 : XNOR2_X1 port map( A => n14604, B => n14603, ZN => n15262);
   U17980 : INV_X1 port map( A => n15262, ZN => n15790);
   U17981 : INV_X1 port map( A => n14789, ZN => n14605);
   U17982 : XNOR2_X1 port map( A => n14605, B => n15484, ZN => n14606);
   U17983 : XNOR2_X1 port map( A => n14606, B => n14920, ZN => n14610);
   U17984 : XNOR2_X1 port map( A => n14468, B => n1952, ZN => n14607);
   U17985 : XNOR2_X1 port map( A => n14608, B => n14607, ZN => n14609);
   U17986 : NOR2_X1 port map( A1 => n16043, A2 => n15262, ZN => n16041);
   U17987 : INV_X1 port map( A => n14611, ZN => n14889);
   U17988 : XNOR2_X1 port map( A => n14889, B => n15175, ZN => n14613);
   U17989 : XNOR2_X1 port map( A => n24937, B => n22702, ZN => n14612);
   U17990 : XNOR2_X1 port map( A => n14613, B => n14612, ZN => n14617);
   U17991 : INV_X1 port map( A => n14614, ZN => n14615);
   U17992 : XNOR2_X1 port map( A => n14615, B => n14964, ZN => n14616);
   U17993 : XNOR2_X1 port map( A => n14616, B => n14617, ZN => n14625);
   U17994 : OAI21_X1 port map( B1 => n16041, B2 => n291, A => n16038, ZN => 
                           n14627);
   U17995 : INV_X1 port map( A => n14898, ZN => n14618);
   U17996 : XNOR2_X1 port map( A => n14619, B => n14618, ZN => n14624);
   U17997 : XNOR2_X1 port map( A => n14620, B => n15051, ZN => n14622);
   U17998 : XNOR2_X1 port map( A => n15103, B => n1863, ZN => n14621);
   U17999 : XNOR2_X1 port map( A => n14622, B => n14621, ZN => n14623);
   U18000 : NAND3_X1 port map( A1 => n2251, A2 => n24430, A3 => n15789, ZN => 
                           n14626);
   U18001 : XNOR2_X1 port map( A => n15522, B => n23983, ZN => n14628);
   U18002 : XNOR2_X1 port map( A => n14858, B => n14628, ZN => n14631);
   U18003 : XNOR2_X1 port map( A => n14629, B => n24508, ZN => n15011);
   U18004 : INV_X1 port map( A => n15011, ZN => n14630);
   U18005 : XNOR2_X1 port map( A => n14631, B => n14630, ZN => n14632);
   U18006 : XNOR2_X1 port map( A => n14634, B => n1776, ZN => n14635);
   U18007 : XNOR2_X1 port map( A => n14635, B => n15321, ZN => n14637);
   U18008 : XNOR2_X1 port map( A => n15133, B => n15318, ZN => n14636);
   U18009 : XNOR2_X1 port map( A => n14637, B => n14636, ZN => n14641);
   U18010 : INV_X1 port map( A => n14638, ZN => n14639);
   U18011 : XNOR2_X1 port map( A => n14639, B => n15499, ZN => n14640);
   U18012 : XNOR2_X1 port map( A => n14642, B => n15005, ZN => n15482);
   U18013 : INV_X1 port map( A => n15332, ZN => n14643);
   U18014 : XNOR2_X1 port map( A => n14643, B => n15482, ZN => n14648);
   U18015 : XNOR2_X1 port map( A => n14644, B => n15415, ZN => n14646);
   U18016 : XNOR2_X1 port map( A => n15003, B => n889, ZN => n14645);
   U18017 : XNOR2_X1 port map( A => n14646, B => n14645, ZN => n14647);
   U18018 : XNOR2_X1 port map( A => n15138, B => n21623, ZN => n14650);
   U18019 : XNOR2_X1 port map( A => n14649, B => n14650, ZN => n14651);
   U18020 : XNOR2_X1 port map( A => n14651, B => n14652, ZN => n14664);
   U18021 : INV_X1 port map( A => n14664, ZN => n15799);
   U18022 : XNOR2_X1 port map( A => n15071, B => n15095, ZN => n14987);
   U18023 : XNOR2_X1 port map( A => n14987, B => n14653, ZN => n14657);
   U18024 : XNOR2_X1 port map( A => n14846, B => n876, ZN => n14655);
   U18025 : XNOR2_X1 port map( A => n14654, B => n14907, ZN => n15503);
   U18026 : XNOR2_X1 port map( A => n14655, B => n15503, ZN => n14656);
   U18027 : NAND2_X1 port map( A1 => n15799, A2 => n16129, ZN => n16131);
   U18028 : INV_X1 port map( A => n16129, ZN => n15800);
   U18029 : XNOR2_X1 port map( A => n14902, B => n14996, ZN => n15247);
   U18030 : INV_X1 port map( A => n15247, ZN => n15512);
   U18031 : XNOR2_X1 port map( A => n15512, B => n15348, ZN => n14661);
   U18032 : XNOR2_X1 port map( A => n14993, B => n15444, ZN => n14659);
   U18033 : XNOR2_X1 port map( A => n15153, B => n891, ZN => n14658);
   U18034 : XNOR2_X1 port map( A => n14659, B => n14658, ZN => n14660);
   U18035 : INV_X1 port map( A => n16076, ZN => n16130);
   U18036 : NAND2_X1 port map( A1 => n16131, A2 => n14662, ZN => n14663);
   U18037 : NAND2_X1 port map( A1 => n16077, A2 => n16129, ZN => n15312);
   U18038 : INV_X1 port map( A => n15312, ZN => n14665);
   U18039 : NAND2_X1 port map( A1 => n14665, A2 => n1365, ZN => n14666);
   U18040 : XNOR2_X1 port map( A => n15374, B => n14827, ZN => n15156);
   U18041 : XNOR2_X1 port map( A => n14667, B => n14826, ZN => n15447);
   U18042 : XNOR2_X1 port map( A => n15347, B => n14936, ZN => n15195);
   U18043 : XNOR2_X1 port map( A => n15514, B => n869, ZN => n14668);
   U18044 : INV_X1 port map( A => n14669, ZN => n14670);
   U18045 : XNOR2_X1 port map( A => n14670, B => n14799, ZN => n15147);
   U18046 : XNOR2_X1 port map( A => n14671, B => n15097, ZN => n15454);
   U18047 : XNOR2_X1 port map( A => n15454, B => n15147, ZN => n14674);
   U18048 : XNOR2_X1 port map( A => n15505, B => n22986, ZN => n14672);
   U18049 : XNOR2_X1 port map( A => n15185, B => n14672, ZN => n14673);
   U18050 : INV_X1 port map( A => n14676, ZN => n14791);
   U18051 : XNOR2_X1 port map( A => n1362, B => n14791, ZN => n15139);
   U18052 : XNOR2_X1 port map( A => n14677, B => n15139, ZN => n14681);
   U18053 : XNOR2_X1 port map( A => n14678, B => n15088, ZN => n15438);
   U18054 : XNOR2_X1 port map( A => n15488, B => n2211, ZN => n14679);
   U18055 : XNOR2_X1 port map( A => n15438, B => n14679, ZN => n14680);
   U18056 : INV_X1 port map( A => n14686, ZN => n14684);
   U18057 : INV_X1 port map( A => n14685, ZN => n14683);
   U18058 : INV_X1 port map( A => n2989, ZN => n14682);
   U18059 : OAI21_X1 port map( B1 => n14684, B2 => n14683, A => n14682, ZN => 
                           n14688);
   U18060 : NAND3_X1 port map( A1 => n14686, A2 => n2989, A3 => n14685, ZN => 
                           n14687);
   U18061 : NAND2_X1 port map( A1 => n14688, A2 => n14687, ZN => n14689);
   U18062 : XNOR2_X1 port map( A => n15082, B => n14690, ZN => n15420);
   U18063 : XNOR2_X1 port map( A => n15420, B => n14691, ZN => n14692);
   U18064 : NAND2_X1 port map( A1 => n24532, A2 => n16109, ZN => n14702);
   U18065 : XNOR2_X1 port map( A => n14694, B => n14805, ZN => n14696);
   U18066 : XNOR2_X1 port map( A => n14857, B => n2100, ZN => n14695);
   U18067 : XNOR2_X1 port map( A => n14696, B => n14695, ZN => n14701);
   U18068 : XNOR2_X1 port map( A => n14697, B => n14698, ZN => n15429);
   U18069 : XNOR2_X1 port map( A => n14699, B => n15429, ZN => n14700);
   U18070 : XNOR2_X1 port map( A => n14834, B => n14703, ZN => n15131);
   U18071 : XNOR2_X1 port map( A => n15131, B => n14704, ZN => n14707);
   U18072 : XNOR2_X1 port map( A => n15396, B => n881, ZN => n14705);
   U18073 : XNOR2_X1 port map( A => n15461, B => n14705, ZN => n14706);
   U18074 : NOR2_X1 port map( A1 => n16107, A2 => n15782, ZN => n14708);
   U18076 : INV_X1 port map( A => n15804, ZN => n16114);
   U18078 : XNOR2_X1 port map( A => n14755, B => n14982, ZN => n15339);
   U18079 : XNOR2_X1 port map( A => n14928, B => n14788, ZN => n15291);
   U18080 : XNOR2_X1 port map( A => n15291, B => n15339, ZN => n14713);
   U18081 : XNOR2_X1 port map( A => n15483, B => n24502, ZN => n14711);
   U18082 : XNOR2_X1 port map( A => n14976, B => n5286, ZN => n14710);
   U18083 : XNOR2_X1 port map( A => n14711, B => n14710, ZN => n14712);
   U18084 : XNOR2_X1 port map( A => n14715, B => n14714, ZN => n14718);
   U18085 : XNOR2_X1 port map( A => n15153, B => n2040, ZN => n14716);
   U18086 : XNOR2_X1 port map( A => n15351, B => n14716, ZN => n14717);
   U18087 : XNOR2_X1 port map( A => n15230, B => n14719, ZN => n15325);
   U18088 : XNOR2_X1 port map( A => n15526, B => n1777, ZN => n14720);
   U18089 : XNOR2_X1 port map( A => n15325, B => n14720, ZN => n14723);
   U18090 : XNOR2_X1 port map( A => n15427, B => n15269, ZN => n14722);
   U18091 : XNOR2_X1 port map( A => n15462, B => n15126, ZN => n14728);
   U18092 : XNOR2_X1 port map( A => n15273, B => n1835, ZN => n14726);
   U18093 : XNOR2_X1 port map( A => n14726, B => n14725, ZN => n14727);
   U18094 : XNOR2_X1 port map( A => n14728, B => n14727, ZN => n16080);
   U18095 : NAND2_X1 port map( A1 => n16080, A2 => n15584, ZN => n16082);
   U18096 : INV_X1 port map( A => n14729, ZN => n14730);
   U18097 : XNOR2_X1 port map( A => n14730, B => n15331, ZN => n14736);
   U18098 : INV_X1 port map( A => n14731, ZN => n14734);
   U18099 : XNOR2_X1 port map( A => n15285, B => n20744, ZN => n14733);
   U18100 : XNOR2_X1 port map( A => n14734, B => n14733, ZN => n14735);
   U18101 : NOR2_X1 port map( A1 => n16100, A2 => n15584, ZN => n15780);
   U18102 : XNOR2_X1 port map( A => n14737, B => n15253, ZN => n15356);
   U18103 : XNOR2_X1 port map( A => n15356, B => n14738, ZN => n14742);
   U18104 : INV_X1 port map( A => n14739, ZN => n14741);
   U18105 : XNOR2_X1 port map( A => n14960, B => n2745, ZN => n14740);
   U18106 : INV_X1 port map( A => n17273, ZN => n17254);
   U18107 : INV_X1 port map( A => n17272, ZN => n17279);
   U18108 : OAI21_X1 port map( B1 => n16151, B2 => n213, A => n16095, ZN => 
                           n14744);
   U18112 : INV_X1 port map( A => n14749, ZN => n14750);
   U18113 : XNOR2_X1 port map( A => n15093, B => n14750, ZN => n14754);
   U18114 : XNOR2_X1 port map( A => n14988, B => n15506, ZN => n14752);
   U18115 : XNOR2_X1 port map( A => n14799, B => n924, ZN => n14751);
   U18116 : XNOR2_X1 port map( A => n14752, B => n14751, ZN => n14753);
   U18117 : XNOR2_X1 port map( A => n14754, B => n14753, ZN => n15938);
   U18118 : XNOR2_X1 port map( A => n14755, B => n15484, ZN => n14758);
   U18119 : XNOR2_X1 port map( A => n14756, B => n14791, ZN => n14757);
   U18120 : XNOR2_X1 port map( A => n14757, B => n14758, ZN => n14762);
   U18121 : XNOR2_X1 port map( A => n15436, B => n15483, ZN => n14760);
   U18122 : XNOR2_X1 port map( A => n14976, B => n2761, ZN => n14759);
   U18123 : XNOR2_X1 port map( A => n14760, B => n14759, ZN => n14761);
   U18124 : XNOR2_X2 port map( A => n14762, B => n14761, ZN => n16247);
   U18125 : INV_X1 port map( A => n15526, ZN => n14764);
   U18126 : XNOR2_X1 port map( A => n14764, B => n14805, ZN => n15159);
   U18127 : XNOR2_X1 port map( A => n15056, B => n2903, ZN => n14765);
   U18128 : XNOR2_X1 port map( A => n15159, B => n14765, ZN => n14766);
   U18129 : XNOR2_X1 port map( A => n14766, B => n14767, ZN => n15764);
   U18130 : INV_X1 port map( A => n15764, ZN => n16018);
   U18131 : NAND2_X1 port map( A1 => n16247, A2 => n16018, ZN => n14787);
   U18132 : XNOR2_X1 port map( A => n14827, B => n765, ZN => n14768);
   U18133 : XNOR2_X1 port map( A => n14769, B => n14768, ZN => n14772);
   U18134 : XNOR2_X1 port map( A => n15113, B => n14770, ZN => n14771);
   U18137 : XNOR2_X1 port map( A => n14834, B => n15464, ZN => n14774);
   U18138 : XNOR2_X1 port map( A => n15062, B => n15219, ZN => n14773);
   U18139 : XNOR2_X1 port map( A => n14773, B => n14774, ZN => n14779);
   U18140 : XNOR2_X1 port map( A => n15393, B => n2805, ZN => n14777);
   U18141 : XNOR2_X1 port map( A => n15497, B => n14775, ZN => n14776);
   U18142 : XNOR2_X1 port map( A => n14776, B => n14777, ZN => n14778);
   U18143 : XNOR2_X1 port map( A => n14779, B => n14778, ZN => n15762);
   U18145 : XNOR2_X1 port map( A => n15480, B => n14815, ZN => n15141);
   U18146 : INV_X1 port map( A => n14780, ZN => n15081);
   U18147 : XNOR2_X1 port map( A => n15081, B => n15141, ZN => n14784);
   U18148 : XNOR2_X1 port map( A => n15422, B => n2120, ZN => n14782);
   U18149 : XNOR2_X1 port map( A => n14782, B => n14781, ZN => n14783);
   U18150 : XNOR2_X1 port map( A => n14789, B => n14788, ZN => n15029);
   U18151 : INV_X1 port map( A => n15029, ZN => n14790);
   U18152 : XNOR2_X1 port map( A => n15238, B => n15341, ZN => n15209);
   U18153 : XNOR2_X1 port map( A => n14790, B => n15209, ZN => n14796);
   U18154 : XNOR2_X1 port map( A => n15088, B => n14791, ZN => n14794);
   U18155 : XNOR2_X1 port map( A => n14792, B => n2717, ZN => n14793);
   U18156 : XNOR2_X1 port map( A => n14794, B => n14793, ZN => n14795);
   U18157 : XNOR2_X1 port map( A => n15097, B => n15298, ZN => n14798);
   U18158 : XNOR2_X1 port map( A => n15358, B => n15369, ZN => n14797);
   U18159 : XNOR2_X1 port map( A => n14797, B => n14798, ZN => n14804);
   U18160 : XNOR2_X1 port map( A => n14799, B => n15074, ZN => n14802);
   U18161 : XNOR2_X1 port map( A => n14800, B => n763, ZN => n14801);
   U18162 : XNOR2_X1 port map( A => n14802, B => n14801, ZN => n14803);
   U18164 : XNOR2_X1 port map( A => n15168, B => n14805, ZN => n14808);
   U18165 : XNOR2_X1 port map( A => n14806, B => n15051, ZN => n14807);
   U18166 : XNOR2_X1 port map( A => n14808, B => n14807, ZN => n14813);
   U18167 : XNOR2_X1 port map( A => n2765, B => n15055, ZN => n14811);
   U18168 : XNOR2_X1 port map( A => n14809, B => n21335, ZN => n14810);
   U18169 : XNOR2_X1 port map( A => n14811, B => n14810, ZN => n14812);
   U18170 : NAND2_X1 port map( A1 => n16491, A2 => n16232, ZN => n14823);
   U18171 : INV_X1 port map( A => n15416, ZN => n14814);
   U18172 : XNOR2_X1 port map( A => n14814, B => n14815, ZN => n14818);
   U18173 : XNOR2_X1 port map( A => n15082, B => n14816, ZN => n14817);
   U18174 : XNOR2_X1 port map( A => n14818, B => n14817, ZN => n14822);
   U18175 : XNOR2_X1 port map( A => n15174, B => n15284, ZN => n14820);
   U18176 : XNOR2_X1 port map( A => n24937, B => n21703, ZN => n14819);
   U18177 : XNOR2_X1 port map( A => n14820, B => n14819, ZN => n14821);
   U18178 : OAI22_X1 port map( A1 => n16229, A2 => n14823, B1 => n16230, B2 => 
                           n16232, ZN => n14839);
   U18179 : XNOR2_X1 port map( A => n15347, B => n15375, ZN => n14824);
   U18180 : XNOR2_X1 port map( A => n14825, B => n14824, ZN => n14830);
   U18181 : XNOR2_X1 port map( A => n24976, B => n14826, ZN => n14829);
   U18182 : INV_X1 port map( A => n896, ZN => n23798);
   U18183 : XNOR2_X1 port map( A => n14827, B => n23798, ZN => n14828);
   U18184 : INV_X1 port map( A => n14831, ZN => n14832);
   U18185 : XNOR2_X1 port map( A => n14832, B => n14833, ZN => n14838);
   U18186 : XNOR2_X1 port map( A => n15119, B => n1739, ZN => n14836);
   U18187 : XNOR2_X1 port map( A => n14834, B => n15204, ZN => n14835);
   U18188 : XNOR2_X1 port map( A => n14836, B => n14835, ZN => n14837);
   U18189 : XNOR2_X1 port map( A => n14838, B => n14837, ZN => n16231);
   U18190 : INV_X1 port map( A => n14840, ZN => n14844);
   U18191 : XNOR2_X1 port map( A => n14841, B => n15446, ZN => n14843);
   U18192 : XNOR2_X1 port map( A => n15112, B => n15375, ZN => n14842);
   U18193 : XNOR2_X1 port map( A => n14845, B => n15094, ZN => n14848);
   U18194 : XNOR2_X1 port map( A => n14846, B => n3062, ZN => n14847);
   U18195 : XNOR2_X1 port map( A => n14848, B => n14847, ZN => n14856);
   U18196 : MUX2_X1 port map( A => n24572, B => n14850, S => n14849, Z => 
                           n14853);
   U18197 : XNOR2_X1 port map( A => n15451, B => n15369, ZN => n14854);
   U18198 : XNOR2_X1 port map( A => n14854, B => n15367, ZN => n14855);
   U18199 : XNOR2_X1 port map( A => n15169, B => n1864, ZN => n14859);
   U18200 : XNOR2_X1 port map( A => n15160, B => n14859, ZN => n14863);
   U18201 : INV_X1 port map( A => n14860, ZN => n14861);
   U18202 : XNOR2_X1 port map( A => n15431, B => n15103, ZN => n14895);
   U18203 : XNOR2_X1 port map( A => n14861, B => n14895, ZN => n14862);
   U18204 : NAND2_X1 port map( A1 => n14864, A2 => n16458, ZN => n14888);
   U18206 : XNOR2_X1 port map( A => n14477, B => n14865, ZN => n14866);
   U18207 : XNOR2_X1 port map( A => n14867, B => n14866, ZN => n14872);
   U18208 : XNOR2_X1 port map( A => n14868, B => n24502, ZN => n14870);
   U18209 : XNOR2_X1 port map( A => n15210, B => n1855, ZN => n14869);
   U18210 : XNOR2_X1 port map( A => n14870, B => n14869, ZN => n14871);
   U18211 : INV_X1 port map( A => n14873, ZN => n14874);
   U18212 : XNOR2_X1 port map( A => n14874, B => n15392, ZN => n14878);
   U18213 : XNOR2_X1 port map( A => n15063, B => n15133, ZN => n14876);
   U18214 : XNOR2_X1 port map( A => n15120, B => n925, ZN => n14875);
   U18215 : XNOR2_X1 port map( A => n14876, B => n14875, ZN => n14877);
   U18216 : XNOR2_X1 port map( A => n14881, B => n15415, ZN => n14883);
   U18217 : XNOR2_X1 port map( A => n14889, B => n15174, ZN => n14882);
   U18218 : XNOR2_X1 port map( A => n14883, B => n14882, ZN => n14886);
   U18219 : INV_X1 port map( A => n14884, ZN => n14885);
   U18220 : INV_X1 port map( A => n17608, ZN => n16940);
   U18221 : INV_X1 port map( A => n15084, ZN => n14890);
   U18222 : XNOR2_X1 port map( A => n14892, B => n15175, ZN => n14894);
   U18223 : XNOR2_X1 port map( A => n15476, B => n2743, ZN => n14893);
   U18224 : XNOR2_X1 port map( A => n14895, B => n14896, ZN => n14899);
   U18225 : XNOR2_X1 port map( A => n14900, B => n853, ZN => n14901);
   U18226 : XNOR2_X1 port map( A => n14902, B => n15194, ZN => n14903);
   U18227 : INV_X1 port map( A => n15514, ZN => n14904);
   U18228 : XNOR2_X1 port map( A => n14906, B => n14905, ZN => n14926);
   U18229 : INV_X1 port map( A => n14926, ZN => n15572);
   U18230 : XNOR2_X1 port map( A => n14907, B => n887, ZN => n14908);
   U18231 : XNOR2_X1 port map( A => n14908, B => n15095, ZN => n14910);
   U18232 : XNOR2_X1 port map( A => n14909, B => n14910, ZN => n14914);
   U18233 : XNOR2_X1 port map( A => n14912, B => n14911, ZN => n14913);
   U18234 : XNOR2_X1 port map( A => n14914, B => n14913, ZN => n16028);
   U18235 : AOI22_X1 port map( A1 => n16274, A2 => n16029, B1 => n15572, B2 => 
                           n16028, ZN => n16280);
   U18236 : XNOR2_X1 port map( A => n15463, B => n15321, ZN => n14916);
   U18237 : XNOR2_X1 port map( A => n15120, B => n2241, ZN => n14917);
   U18238 : XNOR2_X1 port map( A => n14917, B => n15495, ZN => n14918);
   U18239 : XNOR2_X1 port map( A => n14477, B => n14919, ZN => n14921);
   U18240 : XNOR2_X1 port map( A => n14920, B => n14921, ZN => n14925);
   U18241 : XNOR2_X1 port map( A => n14980, B => n25013, ZN => n15090);
   U18242 : XNOR2_X1 port map( A => n15488, B => n1745, ZN => n14923);
   U18243 : XNOR2_X1 port map( A => n15090, B => n14923, ZN => n14924);
   U18244 : XNOR2_X1 port map( A => n14925, B => n14924, ZN => n15573);
   U18246 : OAI21_X1 port map( B1 => n24403, B2 => n16277, A => n16028, ZN => 
                           n14927);
   U18247 : MUX2_X1 port map( A => n17607, B => n16940, S => n17615, Z => 
                           n15026);
   U18248 : XNOR2_X1 port map( A => n14928, B => n15387, ZN => n14931);
   U18249 : INV_X1 port map( A => n14929, ZN => n14930);
   U18250 : XNOR2_X1 port map( A => n14930, B => n14931, ZN => n14935);
   U18251 : XNOR2_X1 port map( A => n15486, B => n2208, ZN => n14932);
   U18252 : XNOR2_X1 port map( A => n14933, B => n14932, ZN => n14934);
   U18253 : XNOR2_X1 port map( A => n14935, B => n14934, ZN => n14970);
   U18254 : XNOR2_X1 port map( A => n15378, B => n14936, ZN => n15306);
   U18255 : XNOR2_X1 port map( A => n14937, B => n15306, ZN => n14942);
   U18256 : INV_X1 port map( A => n14993, ZN => n14938);
   U18257 : XNOR2_X1 port map( A => n14938, B => n3115, ZN => n14939);
   U18258 : XNOR2_X1 port map( A => n14939, B => n14940, ZN => n14941);
   U18260 : NOR2_X1 port map( A1 => n16448, A2 => n16447, ZN => n14963);
   U18262 : MUX2_X1 port map( A => n14948, B => n14947, S => n14946, Z => 
                           n14951);
   U18263 : XNOR2_X1 port map( A => n14952, B => n15494, ZN => n14953);
   U18264 : XNOR2_X1 port map( A => n15201, B => n14953, ZN => n14957);
   U18265 : XNOR2_X1 port map( A => n15275, B => n1757, ZN => n14954);
   U18266 : XNOR2_X1 port map( A => n14954, B => n14955, ZN => n14956);
   U18267 : XNOR2_X1 port map( A => n14956, B => n14957, ZN => n16452);
   U18268 : INV_X1 port map( A => n14958, ZN => n14959);
   U18269 : XNOR2_X1 port map( A => n14959, B => n14960, ZN => n15296);
   U18270 : XNOR2_X1 port map( A => n15071, B => n3129, ZN => n14962);
   U18271 : AOI22_X1 port map( A1 => n14963, A2 => n16452, B1 => n223, B2 => 
                           n16448, ZN => n14975);
   U18272 : XNOR2_X1 port map( A => n14965, B => n14964, ZN => n14969);
   U18273 : XNOR2_X1 port map( A => n15282, B => n15003, ZN => n14967);
   U18274 : XNOR2_X1 port map( A => n14967, B => n14966, ZN => n14968);
   U18275 : XNOR2_X1 port map( A => n15521, B => n23476, ZN => n14971);
   U18276 : INV_X1 port map( A => n17409, ZN => n17255);
   U18279 : XNOR2_X1 port map( A => n15486, B => n15387, ZN => n14983);
   U18280 : XNOR2_X1 port map( A => n14983, B => n1359, ZN => n14984);
   U18281 : INV_X1 port map( A => n15774, ZN => n16303);
   U18282 : XNOR2_X1 port map( A => n14986, B => n14987, ZN => n14991);
   U18283 : XNOR2_X1 port map( A => n14988, B => n21204, ZN => n14989);
   U18284 : XNOR2_X1 port map( A => n15252, B => n14989, ZN => n14990);
   U18285 : INV_X1 port map( A => n16022, ZN => n16224);
   U18286 : XNOR2_X1 port map( A => n14993, B => n25416, ZN => n15032);
   U18287 : INV_X1 port map( A => n15032, ZN => n14995);
   U18288 : INV_X1 port map( A => n15246, ZN => n14994);
   U18290 : XNOR2_X1 port map( A => n15109, B => n14996, ZN => n14999);
   U18291 : XNOR2_X1 port map( A => n14997, B => n663, ZN => n14998);
   U18292 : XNOR2_X1 port map( A => n14999, B => n14998, ZN => n15000);
   U18293 : XNOR2_X1 port map( A => n15422, B => n15003, ZN => n15039);
   U18294 : XNOR2_X1 port map( A => n15039, B => n15004, ZN => n15008);
   U18295 : XNOR2_X1 port map( A => n1351, B => n2747, ZN => n15006);
   U18296 : XNOR2_X1 port map( A => n15225, B => n15006, ZN => n15007);
   U18297 : OAI21_X1 port map( B1 => n16224, B2 => n16225, A => n16226, ZN => 
                           n15024);
   U18298 : XNOR2_X1 port map( A => n15056, B => n2735, ZN => n15009);
   U18299 : XNOR2_X1 port map( A => n15010, B => n15009, ZN => n15014);
   U18300 : XNOR2_X1 port map( A => n15012, B => n15011, ZN => n15013);
   U18301 : INV_X1 port map( A => n16226, ZN => n15773);
   U18302 : XNOR2_X1 port map( A => n25443, B => n1810, ZN => n15015);
   U18303 : XNOR2_X1 port map( A => n15015, B => n15321, ZN => n15017);
   U18304 : XNOR2_X1 port map( A => n15017, B => n15016, ZN => n15021);
   U18305 : XNOR2_X1 port map( A => n15062, B => n25426, ZN => n15018);
   U18306 : XNOR2_X1 port map( A => n15019, B => n15018, ZN => n15020);
   U18307 : XNOR2_X1 port map( A => n18251, B => n18326, ZN => n17897);
   U18308 : XNOR2_X1 port map( A => n17897, B => n18323, ZN => n15555);
   U18309 : XNOR2_X1 port map( A => n15486, B => n20825, ZN => n15027);
   U18310 : XNOR2_X1 port map( A => n15028, B => n15027, ZN => n15031);
   U18311 : XNOR2_X1 port map( A => n15029, B => n15438, ZN => n15030);
   U18312 : XNOR2_X1 port map( A => n15032, B => n15447, ZN => n15038);
   U18313 : XNOR2_X1 port map( A => n24976, B => n15033, ZN => n15036);
   U18314 : XNOR2_X1 port map( A => n15034, B => n886, ZN => n15035);
   U18315 : XNOR2_X1 port map( A => n15036, B => n15035, ZN => n15037);
   U18316 : XNOR2_X1 port map( A => n15038, B => n15037, ZN => n16341);
   U18317 : INV_X1 port map( A => n16341, ZN => n16285);
   U18318 : XNOR2_X1 port map( A => n15420, B => n15039, ZN => n15050);
   U18319 : XNOR2_X1 port map( A => n24938, B => n15284, ZN => n15048);
   U18320 : INV_X1 port map( A => n15044, ZN => n15042);
   U18321 : INV_X1 port map( A => n15043, ZN => n15041);
   U18322 : OAI21_X1 port map( B1 => n15042, B2 => n15041, A => n21079, ZN => 
                           n15046);
   U18323 : NAND3_X1 port map( A1 => n15044, A2 => n2991, A3 => n15043, ZN => 
                           n15045);
   U18324 : NAND2_X1 port map( A1 => n15046, A2 => n15045, ZN => n15047);
   U18325 : XNOR2_X1 port map( A => n15048, B => n15047, ZN => n15049);
   U18327 : XNOR2_X1 port map( A => n15521, B => n15051, ZN => n15053);
   U18328 : INV_X1 port map( A => n15429, ZN => n15052);
   U18329 : XNOR2_X1 port map( A => n15052, B => n15053, ZN => n15060);
   U18330 : XNOR2_X1 port map( A => n15054, B => n2757, ZN => n15058);
   U18331 : XNOR2_X1 port map( A => n15055, B => n15056, ZN => n15057);
   U18332 : XNOR2_X1 port map( A => n15058, B => n15057, ZN => n15059);
   U18335 : NAND2_X1 port map( A1 => n1654, A2 => n16341, ZN => n15061);
   U18336 : XNOR2_X1 port map( A => n15494, B => n15318, ZN => n15065);
   U18337 : XNOR2_X1 port map( A => n15063, B => n15062, ZN => n15064);
   U18338 : XNOR2_X1 port map( A => n15065, B => n15064, ZN => n15068);
   U18339 : XNOR2_X1 port map( A => n15274, B => n688, ZN => n15066);
   U18340 : XNOR2_X1 port map( A => n15461, B => n15066, ZN => n15067);
   U18341 : XNOR2_X1 port map( A => n15067, B => n15068, ZN => n16345);
   U18342 : NAND3_X1 port map( A1 => n16345, A2 => n25441, A3 => n24539, ZN => 
                           n15080);
   U18343 : XNOR2_X1 port map( A => n15069, B => n15070, ZN => n15078);
   U18344 : INV_X1 port map( A => n15071, ZN => n15073);
   U18345 : INV_X1 port map( A => n15298, ZN => n15072);
   U18346 : XNOR2_X1 port map( A => n15074, B => n1826, ZN => n15075);
   U18348 : NAND3_X1 port map( A1 => n16342, A2 => n1122, A3 => n1654, ZN => 
                           n15079);
   U18349 : XNOR2_X1 port map( A => n15081, B => n15331, ZN => n15086);
   U18350 : XNOR2_X1 port map( A => n15082, B => n20609, ZN => n15083);
   U18351 : XNOR2_X1 port map( A => n15084, B => n15083, ZN => n15085);
   U18352 : XNOR2_X1 port map( A => n15087, B => n15339, ZN => n15092);
   U18353 : XNOR2_X1 port map( A => n15088, B => n677, ZN => n15089);
   U18354 : XNOR2_X1 port map( A => n15090, B => n15089, ZN => n15091);
   U18355 : XNOR2_X1 port map( A => n15092, B => n15091, ZN => n16355);
   U18356 : XNOR2_X1 port map( A => n15093, B => n15356, ZN => n15101);
   U18357 : XNOR2_X1 port map( A => n15094, B => n2477, ZN => n15096);
   U18358 : INV_X1 port map( A => n15097, ZN => n15098);
   U18359 : INV_X1 port map( A => n16359, ZN => n16293);
   U18360 : INV_X1 port map( A => n15102, ZN => n15105);
   U18361 : XNOR2_X1 port map( A => n15103, B => n16574, ZN => n15104);
   U18362 : XNOR2_X1 port map( A => n15105, B => n15104, ZN => n15108);
   U18363 : XNOR2_X1 port map( A => n15325, B => n15106, ZN => n15107);
   U18366 : NOR2_X1 port map( A1 => n16293, A2 => n3451, ZN => n15118);
   U18368 : XNOR2_X1 port map( A => n15109, B => n92, ZN => n15110);
   U18369 : XNOR2_X1 port map( A => n15110, B => n15351, ZN => n15116);
   U18370 : XNOR2_X1 port map( A => n15113, B => n15114, ZN => n15115);
   U18371 : NOR2_X1 port map( A1 => n16359, A2 => n16360, ZN => n15117);
   U18372 : XNOR2_X1 port map( A => n15119, B => n21046, ZN => n15122);
   U18373 : INV_X1 port map( A => n15120, ZN => n15121);
   U18374 : XNOR2_X1 port map( A => n15122, B => n15121, ZN => n15125);
   U18375 : INV_X1 port map( A => n15123, ZN => n15124);
   U18376 : XNOR2_X1 port map( A => n15125, B => n15124, ZN => n15128);
   U18377 : XNOR2_X1 port map( A => n15319, B => n15321, ZN => n15127);
   U18378 : XNOR2_X1 port map( A => n15128, B => n15127, ZN => n16357);
   U18379 : INV_X1 port map( A => n16357, ZN => n15894);
   U18380 : NOR2_X1 port map( A1 => n15894, A2 => n24456, ZN => n15129);
   U18381 : NAND2_X1 port map( A1 => n15129, A2 => n16290, ZN => n15130);
   U18382 : INV_X1 port map( A => n15131, ZN => n15132);
   U18383 : XNOR2_X1 port map( A => n15132, B => n15271, ZN => n15137);
   U18384 : XNOR2_X1 port map( A => n15133, B => n13873, ZN => n15135);
   U18385 : XNOR2_X1 port map( A => n15497, B => n899, ZN => n15134);
   U18386 : XNOR2_X1 port map( A => n15135, B => n15134, ZN => n15136);
   U18387 : INV_X1 port map( A => n15139, ZN => n15140);
   U18388 : XNOR2_X1 port map( A => n15280, B => n15141, ZN => n15145);
   U18389 : XNOR2_X1 port map( A => n15415, B => n22886, ZN => n15143);
   U18390 : XNOR2_X1 port map( A => n15178, B => n24966, ZN => n15404);
   U18391 : XNOR2_X1 port map( A => n15404, B => n15143, ZN => n15144);
   U18392 : INV_X1 port map( A => n16266, ZN => n15146);
   U18393 : MUX2_X1 port map( A => n16001, B => n24366, S => n15146, Z => 
                           n15163);
   U18394 : INV_X1 port map( A => n15147, ZN => n15148);
   U18395 : XNOR2_X1 port map( A => n15148, B => n15297, ZN => n15152);
   U18396 : XNOR2_X1 port map( A => n15183, B => n1804, ZN => n15149);
   U18397 : XNOR2_X1 port map( A => n15150, B => n15149, ZN => n15151);
   U18398 : XNOR2_X1 port map( A => n15152, B => n15151, ZN => n16002);
   U18399 : INV_X1 port map( A => n16002, ZN => n16269);
   U18400 : XNOR2_X1 port map( A => n15153, B => n16, ZN => n15154);
   U18401 : XNOR2_X1 port map( A => n15155, B => n15154, ZN => n15158);
   U18402 : XNOR2_X1 port map( A => n15156, B => n4556, ZN => n15157);
   U18403 : XNOR2_X1 port map( A => n15410, B => n2746, ZN => n15161);
   U18404 : MUX2_X1 port map( A => n17424, B => n17381, S => n17379, Z => 
                           n15261);
   U18405 : NAND2_X1 port map( A1 => n15573, A2 => n16028, ZN => n15771);
   U18407 : XNOR2_X1 port map( A => n15165, B => n2058, ZN => n15166);
   U18408 : XNOR2_X1 port map( A => n15167, B => n15166, ZN => n15173);
   U18409 : XNOR2_X1 port map( A => n15168, B => n15169, ZN => n15171);
   U18410 : XNOR2_X1 port map( A => n15170, B => n15171, ZN => n15172);
   U18411 : XNOR2_X1 port map( A => n15172, B => n15173, ZN => n16008);
   U18412 : XNOR2_X1 port map( A => n15175, B => n15174, ZN => n15226);
   U18413 : XNOR2_X1 port map( A => n15176, B => n15226, ZN => n15182);
   U18414 : XNOR2_X1 port map( A => n15177, B => n15401, ZN => n15180);
   U18415 : XNOR2_X1 port map( A => n15178, B => n2036, ZN => n15179);
   U18416 : XNOR2_X1 port map( A => n15180, B => n15179, ZN => n15181);
   U18417 : NAND2_X1 port map( A1 => n3554, A2 => n16311, ZN => n16638);
   U18418 : INV_X1 port map( A => n16638, ZN => n15216);
   U18419 : XNOR2_X1 port map( A => n15185, B => n15186, ZN => n15189);
   U18420 : XNOR2_X1 port map( A => n15369, B => n15187, ZN => n15251);
   U18421 : XNOR2_X1 port map( A => n15191, B => n15190, ZN => n15193);
   U18422 : XNOR2_X1 port map( A => n14579, B => n2744, ZN => n15192);
   U18423 : XNOR2_X1 port map( A => n15193, B => n15192, ZN => n15197);
   U18424 : XNOR2_X1 port map( A => n15375, B => n15194, ZN => n15248);
   U18425 : XNOR2_X1 port map( A => n15248, B => n15195, ZN => n15196);
   U18426 : XNOR2_X1 port map( A => n15196, B => n15197, ZN => n15556);
   U18427 : AND2_X1 port map( A1 => n15767, A2 => n24297, ZN => n15215);
   U18428 : XNOR2_X1 port map( A => n15200, B => n15199, ZN => n15202);
   U18429 : XNOR2_X1 port map( A => n15201, B => n15202, ZN => n15207);
   U18430 : INV_X1 port map( A => n15203, ZN => n15465);
   U18431 : XNOR2_X1 port map( A => n15465, B => n2726, ZN => n15205);
   U18432 : XNOR2_X1 port map( A => n25436, B => n15204, ZN => n15217);
   U18433 : XNOR2_X1 port map( A => n15205, B => n15217, ZN => n15206);
   U18435 : XNOR2_X1 port map( A => n15209, B => n15208, ZN => n15214);
   U18436 : XNOR2_X1 port map( A => n15487, B => n1758, ZN => n15212);
   U18437 : XNOR2_X1 port map( A => n15386, B => n15210, ZN => n15211);
   U18438 : XNOR2_X1 port map( A => n15212, B => n15211, ZN => n15213);
   U18439 : NAND2_X1 port map( A1 => n16945, A2 => n17424, ZN => n17378);
   U18440 : NAND2_X1 port map( A1 => n16644, A2 => n17378, ZN => n15260);
   U18441 : XNOR2_X1 port map( A => n15218, B => n15217, ZN => n15222);
   U18442 : XNOR2_X1 port map( A => n15219, B => n2222, ZN => n15220);
   U18443 : XNOR2_X1 port map( A => n15499, B => n15220, ZN => n15221);
   U18444 : XNOR2_X1 port map( A => n15223, B => n3093, ZN => n15224);
   U18445 : XNOR2_X1 port map( A => n15482, B => n15224, ZN => n15228);
   U18446 : XNOR2_X1 port map( A => n15225, B => n15226, ZN => n15227);
   U18447 : INV_X1 port map( A => n15229, ZN => n15520);
   U18448 : XNOR2_X1 port map( A => n15230, B => n15520, ZN => n15233);
   U18449 : XNOR2_X1 port map( A => n2765, B => n15409, ZN => n15232);
   U18450 : XNOR2_X1 port map( A => n15233, B => n15232, ZN => n15237);
   U18451 : XNOR2_X1 port map( A => n25384, B => n15326, ZN => n15235);
   U18452 : XNOR2_X1 port map( A => n15165, B => n23699, ZN => n15234);
   U18453 : XNOR2_X1 port map( A => n15235, B => n15234, ZN => n15236);
   U18454 : INV_X1 port map( A => n15674, ZN => n16197);
   U18455 : XNOR2_X1 port map( A => n15387, B => n768, ZN => n15240);
   U18456 : XNOR2_X1 port map( A => n15241, B => n15240, ZN => n15242);
   U18457 : INV_X1 port map( A => n16324, ZN => n15742);
   U18458 : XNOR2_X1 port map( A => n15244, B => n2739, ZN => n15245);
   U18459 : XNOR2_X1 port map( A => n15246, B => n15245, ZN => n15250);
   U18460 : XNOR2_X1 port map( A => n15248, B => n15247, ZN => n15249);
   U18461 : XNOR2_X1 port map( A => n15249, B => n15250, ZN => n16323);
   U18462 : INV_X1 port map( A => n16323, ZN => n16193);
   U18463 : XNOR2_X1 port map( A => n15251, B => n15503, ZN => n15257);
   U18468 : AND2_X1 port map( A1 => n15262, A2 => n16043, ZN => n15263);
   U18469 : OAI21_X1 port map( B1 => n15263, B2 => n15789, A => n24430, ZN => 
                           n15265);
   U18470 : INV_X1 port map( A => n15270, ZN => n15272);
   U18471 : XNOR2_X1 port map( A => n15272, B => n15271, ZN => n15279);
   U18472 : XNOR2_X1 port map( A => n15273, B => n888, ZN => n15277);
   U18473 : XNOR2_X1 port map( A => n25426, B => n15274, ZN => n15276);
   U18474 : XNOR2_X1 port map( A => n15277, B => n15276, ZN => n15278);
   U18475 : XNOR2_X1 port map( A => n15280, B => n15281, ZN => n15289);
   U18476 : INV_X1 port map( A => n15282, ZN => n15283);
   U18477 : XNOR2_X1 port map( A => n15284, B => n15283, ZN => n15287);
   U18478 : XNOR2_X1 port map( A => n15285, B => n681, ZN => n15286);
   U18479 : XNOR2_X1 port map( A => n15287, B => n15286, ZN => n15288);
   U18480 : XNOR2_X1 port map( A => n15290, B => n15291, ZN => n15295);
   U18481 : XNOR2_X1 port map( A => n15387, B => n1364, ZN => n15292);
   U18482 : XNOR2_X1 port map( A => n15293, B => n15292, ZN => n15294);
   U18483 : XNOR2_X1 port map( A => n15295, B => n15294, ZN => n15706);
   U18484 : XNOR2_X1 port map( A => n15296, B => n15297, ZN => n15302);
   U18485 : XNOR2_X1 port map( A => n15298, B => n2044, ZN => n15300);
   U18486 : XNOR2_X1 port map( A => n15300, B => n15299, ZN => n15301);
   U18487 : XNOR2_X1 port map( A => n15302, B => n15301, ZN => n15605);
   U18488 : NAND3_X1 port map( A1 => n294, A2 => n4541, A3 => n15605, ZN => 
                           n15310);
   U18489 : XNOR2_X1 port map( A => n24975, B => n3118, ZN => n15305);
   U18490 : XNOR2_X1 port map( A => n15306, B => n15305, ZN => n15307);
   U18491 : NOR2_X1 port map( A1 => n17342, A2 => n17241, ZN => n17202);
   U18493 : NAND3_X1 port map( A1 => n15802, A2 => n15799, A3 => n16076, ZN => 
                           n15311);
   U18494 : XNOR2_X1 port map( A => n15316, B => n2042, ZN => n15317);
   U18496 : XNOR2_X1 port map( A => n15465, B => n15497, ZN => n15322);
   U18497 : XNOR2_X1 port map( A => n15322, B => n15321, ZN => n15323);
   U18498 : XNOR2_X1 port map( A => n15324, B => n15325, ZN => n15330);
   U18499 : XNOR2_X1 port map( A => n15168, B => n15326, ZN => n15328);
   U18500 : XNOR2_X1 port map( A => n15526, B => n5131, ZN => n15327);
   U18501 : XNOR2_X1 port map( A => n15328, B => n15327, ZN => n15329);
   U18502 : XNOR2_X1 port map( A => n15330, B => n15329, ZN => n15696);
   U18503 : XNOR2_X1 port map( A => n15332, B => n15331, ZN => n15337);
   U18504 : XNOR2_X1 port map( A => n15416, B => n25019, ZN => n15335);
   U18505 : XNOR2_X1 port map( A => n15333, B => n2031, ZN => n15334);
   U18506 : XNOR2_X1 port map( A => n15334, B => n15335, ZN => n15336);
   U18507 : OAI21_X1 port map( B1 => n15695, B2 => n15696, A => n25238, ZN => 
                           n15952);
   U18508 : INV_X1 port map( A => n25237, ZN => n16484);
   U18509 : INV_X1 port map( A => n15338, ZN => n15340);
   U18510 : XNOR2_X1 port map( A => n15340, B => n15339, ZN => n15346);
   U18511 : XNOR2_X1 port map( A => n15342, B => n15341, ZN => n15344);
   U18512 : XNOR2_X1 port map( A => n15483, B => n3084, ZN => n15343);
   U18513 : XNOR2_X1 port map( A => n15344, B => n15343, ZN => n15345);
   U18514 : XNOR2_X1 port map( A => n15349, B => n15348, ZN => n15354);
   U18515 : XNOR2_X1 port map( A => n15350, B => n20995, ZN => n15352);
   U18516 : XNOR2_X1 port map( A => n15354, B => n15353, ZN => n16480);
   U18517 : XNOR2_X1 port map( A => n15356, B => n15355, ZN => n15363);
   U18518 : XNOR2_X1 port map( A => n15359, B => n2087, ZN => n15360);
   U18519 : XNOR2_X1 port map( A => n15361, B => n15360, ZN => n15362);
   U18520 : XNOR2_X1 port map( A => n15363, B => n15362, ZN => n16481);
   U18521 : INV_X1 port map( A => n15695, ZN => n15364);
   U18522 : NAND3_X1 port map( A1 => n15364, A2 => n16480, A3 => n16481, ZN => 
                           n15365);
   U18523 : XNOR2_X1 port map( A => n15366, B => n15367, ZN => n15373);
   U18524 : INV_X1 port map( A => n15368, ZN => n15371);
   U18525 : XNOR2_X1 port map( A => n15369, B => n17960, ZN => n15370);
   U18526 : XNOR2_X1 port map( A => n15371, B => n15370, ZN => n15372);
   U18527 : XNOR2_X1 port map( A => n15375, B => n15514, ZN => n15376);
   U18528 : XNOR2_X1 port map( A => n15376, B => n15377, ZN => n15382);
   U18529 : XNOR2_X1 port map( A => n25501, B => n14579, ZN => n15380);
   U18530 : XNOR2_X1 port map( A => n15378, B => n23271, ZN => n15379);
   U18531 : XNOR2_X1 port map( A => n15380, B => n15379, ZN => n15381);
   U18532 : INV_X1 port map( A => n15383, ZN => n15384);
   U18533 : XNOR2_X1 port map( A => n15385, B => n15384, ZN => n15391);
   U18534 : XNOR2_X1 port map( A => n15484, B => n15386, ZN => n15389);
   U18535 : XNOR2_X1 port map( A => n15387, B => n2034, ZN => n15388);
   U18536 : XNOR2_X1 port map( A => n15389, B => n15388, ZN => n15390);
   U18537 : XNOR2_X2 port map( A => n15391, B => n15390, ZN => n16064);
   U18538 : INV_X1 port map( A => n16064, ZN => n15550);
   U18539 : INV_X1 port map( A => n15392, ZN => n15395);
   U18540 : INV_X1 port map( A => n15393, ZN => n15498);
   U18541 : XNOR2_X1 port map( A => n15498, B => n13873, ZN => n15394);
   U18542 : XNOR2_X1 port map( A => n15395, B => n15394, ZN => n15400);
   U18543 : XNOR2_X1 port map( A => n15396, B => n1827, ZN => n15397);
   U18544 : XNOR2_X1 port map( A => n15398, B => n15397, ZN => n15399);
   U18545 : XNOR2_X1 port map( A => n15478, B => n2782, ZN => n15402);
   U18546 : XNOR2_X1 port map( A => n15405, B => n15406, ZN => n15549);
   U18547 : XNOR2_X1 port map( A => n15407, B => n15408, ZN => n15414);
   U18548 : XNOR2_X1 port map( A => n15409, B => n24423, ZN => n15412);
   U18549 : XNOR2_X1 port map( A => n15412, B => n15411, ZN => n15413);
   U18550 : XNOR2_X1 port map( A => n15414, B => n15413, ZN => n15548);
   U18551 : NOR2_X1 port map( A1 => n17341, A2 => n17346, ZN => n17235);
   U18552 : XNOR2_X1 port map( A => n15416, B => n15415, ZN => n15419);
   U18553 : XNOR2_X1 port map( A => n15417, B => n2190, ZN => n15418);
   U18554 : XNOR2_X1 port map( A => n15419, B => n15418, ZN => n15426);
   U18555 : INV_X1 port map( A => n15420, ZN => n15424);
   U18556 : XNOR2_X1 port map( A => n15422, B => n15421, ZN => n15423);
   U18557 : XNOR2_X1 port map( A => n15424, B => n15423, ZN => n15425);
   U18558 : XNOR2_X1 port map( A => n15425, B => n15426, ZN => n15715);
   U18559 : INV_X1 port map( A => n15427, ZN => n15428);
   U18560 : XNOR2_X1 port map( A => n15428, B => n15429, ZN => n15435);
   U18561 : XNOR2_X1 port map( A => n15430, B => n3183, ZN => n15433);
   U18562 : XNOR2_X1 port map( A => n15168, B => n15431, ZN => n15432);
   U18563 : XNOR2_X1 port map( A => n15433, B => n15432, ZN => n15434);
   U18564 : XNOR2_X1 port map( A => n15436, B => n187, ZN => n15437);
   U18565 : XNOR2_X1 port map( A => n14477, B => n15437, ZN => n15440);
   U18566 : INV_X1 port map( A => n15438, ZN => n15439);
   U18567 : XNOR2_X1 port map( A => n15440, B => n15439, ZN => n15443);
   U18568 : INV_X1 port map( A => n15441, ZN => n15442);
   U18569 : XNOR2_X1 port map( A => n15444, B => n2970, ZN => n15445);
   U18570 : XNOR2_X1 port map( A => n15445, B => n15446, ZN => n15448);
   U18571 : XNOR2_X1 port map( A => n15448, B => n15447, ZN => n15450);
   U18572 : NAND2_X1 port map( A1 => n16474, A2 => n24550, ZN => n15459);
   U18573 : XNOR2_X1 port map( A => n15451, B => n1875, ZN => n15453);
   U18574 : XNOR2_X1 port map( A => n15453, B => n15452, ZN => n15455);
   U18575 : XNOR2_X1 port map( A => n15454, B => n15455, ZN => n15458);
   U18576 : INV_X1 port map( A => n15456, ZN => n15457);
   U18577 : XNOR2_X1 port map( A => n15458, B => n15457, ZN => n15714);
   U18578 : MUX2_X1 port map( A => n15460, B => n15459, S => n16471, Z => 
                           n17237);
   U18579 : XNOR2_X1 port map( A => n15461, B => n15462, ZN => n15469);
   U18580 : XNOR2_X1 port map( A => n15464, B => n15463, ZN => n15467);
   U18581 : XNOR2_X1 port map( A => n15465, B => n2826, ZN => n15466);
   U18582 : XNOR2_X1 port map( A => n15467, B => n15466, ZN => n15468);
   U18583 : INV_X1 port map( A => n16473, ZN => n16476);
   U18584 : NOR2_X1 port map( A1 => n16476, A2 => n16472, ZN => n15471);
   U18585 : NAND2_X1 port map( A1 => n17237, A2 => n3872, ZN => n16780);
   U18586 : NOR2_X1 port map( A1 => n17241, A2 => n17346, ZN => n15472);
   U18587 : XNOR2_X1 port map( A => n18074, B => n18523, ZN => n17987);
   U18588 : MUX2_X1 port map( A => n16484, B => n24981, S => n15953, Z => 
                           n15475);
   U18589 : NOR2_X1 port map( A1 => n25238, A2 => n16480, ZN => n15474);
   U18590 : INV_X1 port map( A => n16481, ZN => n15950);
   U18591 : INV_X1 port map( A => n15872, ZN => n15534);
   U18592 : XNOR2_X1 port map( A => n15476, B => n2228, ZN => n15477);
   U18593 : INV_X1 port map( A => n24956, ZN => n15479);
   U18594 : XNOR2_X1 port map( A => n15479, B => n25019, ZN => n15481);
   U18595 : XNOR2_X1 port map( A => n15484, B => n15483, ZN => n15485);
   U18596 : XNOR2_X1 port map( A => n15486, B => n15487, ZN => n15490);
   U18597 : INV_X1 port map( A => n2990, ZN => n23239);
   U18598 : XNOR2_X1 port map( A => n15488, B => n23239, ZN => n15489);
   U18599 : XNOR2_X1 port map( A => n15490, B => n15489, ZN => n15491);
   U18600 : XNOR2_X1 port map( A => n15492, B => n15491, ZN => n15710);
   U18601 : INV_X1 port map( A => n15710, ZN => n16443);
   U18602 : XNOR2_X1 port map( A => n14384, B => n21423, ZN => n15493);
   U18603 : XNOR2_X1 port map( A => n15493, B => n15494, ZN => n15496);
   U18604 : XNOR2_X1 port map( A => n15496, B => n15495, ZN => n15502);
   U18605 : XNOR2_X1 port map( A => n15498, B => n15497, ZN => n15500);
   U18606 : XNOR2_X1 port map( A => n15500, B => n15499, ZN => n15501);
   U18607 : XNOR2_X1 port map( A => n15502, B => n15501, ZN => n16243);
   U18608 : INV_X1 port map( A => n16243, ZN => n15943);
   U18609 : XNOR2_X1 port map( A => n15505, B => n15506, ZN => n15509);
   U18610 : XNOR2_X1 port map( A => n15507, B => n21553, ZN => n15508);
   U18611 : XNOR2_X1 port map( A => n15509, B => n15508, ZN => n15510);
   U18612 : INV_X1 port map( A => n16437, ZN => n15945);
   U18613 : XNOR2_X1 port map( A => n15512, B => n15513, ZN => n15519);
   U18614 : XNOR2_X1 port map( A => n25501, B => n812, ZN => n15516);
   U18615 : XNOR2_X1 port map( A => n15517, B => n15516, ZN => n15518);
   U18616 : XNOR2_X1 port map( A => n25431, B => n15520, ZN => n15525);
   U18617 : XNOR2_X1 port map( A => n25384, B => n15523, ZN => n15524);
   U18618 : XNOR2_X1 port map( A => n15525, B => n15524, ZN => n15530);
   U18619 : XNOR2_X1 port map( A => n15526, B => n14694, ZN => n15528);
   U18620 : XNOR2_X1 port map( A => n15165, B => n1854, ZN => n15527);
   U18621 : XNOR2_X1 port map( A => n15528, B => n15527, ZN => n15529);
   U18622 : INV_X1 port map( A => n15707, ZN => n15946);
   U18624 : NOR2_X1 port map( A1 => n15952, A2 => n15695, ZN => n15871);
   U18625 : NOR2_X1 port map( A1 => n16578, A2 => n15871, ZN => n15533);
   U18626 : NAND2_X1 port map( A1 => n16043, A2 => n15790, ZN => n15537);
   U18627 : INV_X1 port map( A => n16043, ZN => n15535);
   U18628 : AND2_X1 port map( A1 => n15535, A2 => n16042, ZN => n15788);
   U18630 : NAND2_X1 port map( A1 => n16742, A2 => n15538, ZN => n16653);
   U18631 : INV_X1 port map( A => n16051, ZN => n16509);
   U18632 : NAND2_X1 port map( A1 => n15691, A2 => n16509, ZN => n15544);
   U18633 : NAND2_X1 port map( A1 => n15539, A2 => n16508, ZN => n15543);
   U18637 : MUX2_X1 port map( A => n17087, B => n17086, S => n16578, Z => 
                           n16647);
   U18638 : INV_X1 port map( A => n15548, ZN => n16062);
   U18640 : INV_X1 port map( A => n15694, ZN => n15794);
   U18641 : OAI211_X1 port map( C1 => n16062, C2 => n15794, A => n15550, B => 
                           n16067, ZN => n15551);
   U18642 : XNOR2_X1 port map( A => n18351, B => n869, ZN => n15553);
   U18643 : XNOR2_X1 port map( A => n17987, B => n15553, ZN => n15554);
   U18646 : INV_X1 port map( A => n17335, ZN => n15563);
   U18647 : MUX2_X1 port map( A => n16225, B => n16022, S => n15774, Z => 
                           n15562);
   U18649 : INV_X1 port map( A => n16917, ZN => n16727);
   U18650 : OAI21_X1 port map( B1 => n16974, B2 => n15563, A => n16727, ZN => 
                           n15578);
   U18651 : OAI21_X1 port map( B1 => n15933, B2 => n16230, A => n15565, ZN => 
                           n15566);
   U18652 : INV_X1 port map( A => n16491, ZN => n15937);
   U18653 : INV_X1 port map( A => n16016, ZN => n16251);
   U18654 : AOI21_X1 port map( B1 => n16251, B2 => n16247, A => n2605, ZN => 
                           n15571);
   U18655 : NAND2_X1 port map( A1 => n16247, A2 => n25484, ZN => n15569);
   U18656 : MUX2_X1 port map( A => n15569, B => n15568, S => n16016, Z => 
                           n15570);
   U18657 : OAI21_X1 port map( B1 => n15571, B2 => n16018, A => n15570, ZN => 
                           n17334);
   U18658 : OAI21_X1 port map( B1 => n16971, B2 => n25412, A => n16917, ZN => 
                           n15577);
   U18659 : NOR2_X1 port map( A1 => n15573, A2 => n16028, ZN => n15574);
   U18660 : AOI21_X1 port map( B1 => n17335, B2 => n376, A => n17332, ZN => 
                           n15575);
   U18661 : INV_X1 port map( A => n15579, ZN => n15581);
   U18662 : INV_X1 port map( A => n25409, ZN => n16084);
   U18663 : NAND2_X1 port map( A1 => n16084, A2 => n16105, ZN => n15580);
   U18664 : NAND2_X1 port map( A1 => n15581, A2 => n15580, ZN => n15586);
   U18665 : INV_X1 port map( A => n15582, ZN => n15585);
   U18666 : NAND2_X1 port map( A1 => n16038, A2 => n24429, ZN => n15588);
   U18667 : NAND3_X1 port map( A1 => n15789, A2 => n15790, A3 => n24430, ZN => 
                           n15587);
   U18668 : OAI21_X1 port map( B1 => n24928, B2 => n16107, A => n25030, ZN => 
                           n15591);
   U18669 : INV_X1 port map( A => n16107, ZN => n15783);
   U18671 : NAND3_X1 port map( A1 => n24826, A2 => n16077, A3 => n15801, ZN => 
                           n15597);
   U18672 : NAND3_X1 port map( A1 => n1365, A2 => n16077, A3 => n16076, ZN => 
                           n15596);
   U18674 : NAND2_X1 port map( A1 => n16067, A2 => n16060, ZN => n15599);
   U18679 : INV_X1 port map( A => n17068, ZN => n16730);
   U18680 : XNOR2_X1 port map( A => n18262, B => n18240, ZN => n17906);
   U18681 : NOR2_X1 port map( A1 => n15611, A2 => n14499, ZN => n15614);
   U18682 : NOR2_X1 port map( A1 => n15612, A2 => n15857, ZN => n15613);
   U18683 : NAND3_X1 port map( A1 => n15804, A2 => n16118, A3 => n15857, ZN => 
                           n15615);
   U18684 : OAI21_X1 port map( B1 => n16680, B2 => n16117, A => n15615, ZN => 
                           n15616);
   U18685 : INV_X1 port map( A => n24585, ZN => n15883);
   U18686 : NAND2_X1 port map( A1 => n16125, A2 => n15842, ZN => n15965);
   U18687 : NAND2_X1 port map( A1 => n15965, A2 => n16122, ZN => n15618);
   U18688 : AOI22_X1 port map( A1 => n15620, A2 => n15846, B1 => n15619, B2 => 
                           n15618, ZN => n17061);
   U18689 : INV_X1 port map( A => n17061, ZN => n16929);
   U18691 : INV_X1 port map( A => n16388, ZN => n16162);
   U18692 : NOR2_X1 port map( A1 => n16394, A2 => n16162, ZN => n15847);
   U18693 : NOR2_X1 port map( A1 => n16393, A2 => n15849, ZN => n15622);
   U18694 : OAI21_X1 port map( B1 => n15847, B2 => n15622, A => n15848, ZN => 
                           n15623);
   U18696 : AOI21_X1 port map( B1 => n293, B2 => n15625, A => n16095, ZN => 
                           n15626);
   U18697 : NAND2_X1 port map( A1 => n17059, A2 => n15631, ZN => n16935);
   U18698 : INV_X1 port map( A => n16935, ZN => n15634);
   U18699 : MUX2_X1 port map( A => n16082, B => n15632, S => n16102, Z => 
                           n15633);
   U18700 : NAND2_X1 port map( A1 => n15634, A2 => n17054, ZN => n15636);
   U18701 : NOR2_X1 port map( A1 => n16932, A2 => n24585, ZN => n15880);
   U18702 : NAND2_X1 port map( A1 => n15638, A2 => n15970, ZN => n16187);
   U18703 : NAND2_X1 port map( A1 => n17183, A2 => n15641, ZN => n15644);
   U18704 : NAND2_X1 port map( A1 => n15907, A2 => n16367, ZN => n15642);
   U18705 : NAND3_X1 port map( A1 => n17312, A2 => n17596, A3 => n17597, ZN => 
                           n15664);
   U18707 : NAND2_X1 port map( A1 => n16422, A2 => n16427, ZN => n15648);
   U18708 : MUX2_X1 port map( A => n15649, B => n15648, S => n16170, Z => 
                           n15650);
   U18709 : AOI21_X1 port map( B1 => n25492, B2 => n16412, A => n16414, ZN => 
                           n15651);
   U18710 : NAND2_X1 port map( A1 => n16417, A2 => n16408, ZN => n15984);
   U18711 : MUX2_X1 port map( A => n15651, B => n15984, S => n16413, Z => 
                           n15652);
   U18712 : NOR2_X1 port map( A1 => n17305, A2 => n17316, ZN => n17600);
   U18713 : NAND2_X1 port map( A1 => n2968, A2 => n17600, ZN => n15663);
   U18715 : NAND2_X1 port map( A1 => n16382, A2 => n25210, ZN => n15654);
   U18717 : NOR2_X1 port map( A1 => n4046, A2 => n15837, ZN => n16385);
   U18718 : NAND2_X1 port map( A1 => n16385, A2 => n25210, ZN => n15658);
   U18719 : NAND2_X1 port map( A1 => n17598, A2 => n16921, ZN => n17315);
   U18720 : INV_X1 port map( A => n17315, ZN => n15661);
   U18721 : NAND2_X1 port map( A1 => n17312, A2 => n15661, ZN => n15662);
   U18722 : NAND3_X1 port map( A1 => n17316, A2 => n24542, A3 => n16921, ZN => 
                           n17601);
   U18723 : NAND4_X1 port map( A1 => n15664, A2 => n15663, A3 => n15662, A4 => 
                           n17601, ZN => n15665);
   U18724 : XNOR2_X1 port map( A => n15665, B => n17875, ZN => n18317);
   U18725 : INV_X1 port map( A => n18317, ZN => n15666);
   U18726 : XNOR2_X1 port map( A => n15666, B => n17906, ZN => n15736);
   U18727 : INV_X1 port map( A => n16331, ZN => n15755);
   U18728 : NAND2_X1 port map( A1 => n15755, A2 => n16332, ZN => n15668);
   U18729 : INV_X1 port map( A => n16595, ZN => n15887);
   U18730 : INV_X1 port map( A => n16349, ZN => n15885);
   U18731 : AOI21_X1 port map( B1 => n16597, B2 => n15885, A => n25432, ZN => 
                           n15672);
   U18732 : NAND3_X1 port map( A1 => n17326, A2 => n15673, A3 => n4426, ZN => 
                           n15685);
   U18733 : OAI22_X1 port map( A1 => n1122, A2 => n16285, B1 => n24539, B2 => 
                           n1654, ZN => n16015);
   U18734 : NAND2_X1 port map( A1 => n24540, A2 => n25441, ZN => n16344);
   U18735 : NAND2_X1 port map( A1 => n16015, A2 => n16344, ZN => n15683);
   U18736 : NOR2_X1 port map( A1 => n16345, A2 => n25441, ZN => n15747);
   U18737 : INV_X1 port map( A => n15747, ZN => n15681);
   U18738 : INV_X1 port map( A => n15679, ZN => n15680);
   U18739 : NAND2_X1 port map( A1 => n15681, A2 => n15680, ZN => n15682);
   U18740 : NAND3_X1 port map( A1 => n15673, A2 => n17319, A3 => n16607, ZN => 
                           n15684);
   U18741 : INV_X1 port map( A => n16242, ZN => n15944);
   U18742 : NOR2_X1 port map( A1 => n16243, A2 => n15946, ZN => n16441);
   U18743 : NAND2_X1 port map( A1 => n16443, A2 => n15946, ZN => n15686);
   U18744 : OAI21_X1 port map( B1 => n16450, B2 => n16447, A => n223, ZN => 
                           n15687);
   U18745 : MUX2_X1 port map( A => n24550, B => n16471, S => n16469, Z => 
                           n15690);
   U18746 : AOI21_X1 port map( B1 => n15715, B2 => n16475, A => n16472, ZN => 
                           n15689);
   U18748 : MUX2_X1 port map( A => n15953, B => n16483, S => n16480, Z => 
                           n16485);
   U18749 : INV_X1 port map( A => n15698, ZN => n16547);
   U18750 : AOI21_X1 port map( B1 => n16547, B2 => n16795, A => n16550, ZN => 
                           n15701);
   U18751 : INV_X1 port map( A => n16549, ZN => n15699);
   U18752 : NAND2_X1 port map( A1 => n15699, A2 => n16795, ZN => n15700);
   U18753 : XNOR2_X1 port map( A => n18080, B => n18539, ZN => n15734);
   U18754 : INV_X1 port map( A => n16465, ZN => n16460);
   U18755 : AOI21_X1 port map( B1 => n5269, B2 => n16221, A => n16460, ZN => 
                           n15705);
   U18756 : INV_X1 port map( A => n15921, ZN => n16459);
   U18757 : NOR2_X1 port map( A1 => n15707, A2 => n16242, ZN => n15708);
   U18759 : NAND3_X1 port map( A1 => n16438, A2 => n16437, A3 => n16442, ZN => 
                           n15712);
   U18760 : NAND2_X1 port map( A1 => n16616, A2 => n17299, ZN => n17302);
   U18761 : NOR2_X1 port map( A1 => n16705, A2 => n17299, ZN => n15724);
   U18762 : INV_X1 port map( A => n15714, ZN => n16057);
   U18764 : NOR2_X1 port map( A1 => n16616, A2 => n17297, ZN => n15723);
   U18765 : INV_X1 port map( A => n16480, ZN => n15951);
   U18766 : NOR2_X1 port map( A1 => n15718, A2 => n15717, ZN => n15722);
   U18767 : NOR2_X1 port map( A1 => n15953, A2 => n15950, ZN => n15719);
   U18768 : NAND2_X1 port map( A1 => n15719, A2 => n24981, ZN => n15720);
   U18769 : OAI21_X1 port map( B1 => n15724, B2 => n15723, A => n16708, ZN => 
                           n15732);
   U18770 : INV_X1 port map( A => n16451, ZN => n15725);
   U18772 : XNOR2_X1 port map( A => n18382, B => n21623, ZN => n15733);
   U18773 : XNOR2_X1 port map( A => n15734, B => n15733, ZN => n15735);
   U18774 : NOR2_X1 port map( A1 => n19302, A2 => n19307, ZN => n19130);
   U18775 : NOR2_X1 port map( A1 => n15737, A2 => n16551, ZN => n15741);
   U18777 : NOR2_X2 port map( A1 => n15741, A2 => n15740, ZN => n18188);
   U18778 : INV_X1 port map( A => n16194, ZN => n15744);
   U18779 : NAND2_X1 port map( A1 => n16356, A2 => n16290, ZN => n16363);
   U18780 : OAI22_X1 port map( A1 => n16363, A2 => n25546, B1 => n15748, B2 => 
                           n16290, ZN => n15749);
   U18781 : OAI22_X1 port map( A1 => n16309, A2 => n15751, B1 => n16012, B2 => 
                           n15750, ZN => n15754);
   U18782 : NAND2_X1 port map( A1 => n15557, A2 => n3554, ZN => n15752);
   U18783 : INV_X1 port map( A => n15757, ZN => n15759);
   U18784 : INV_X1 port map( A => n16267, ZN => n15758);
   U18785 : NAND2_X1 port map( A1 => n16230, A2 => n16232, ZN => n16490);
   U18786 : NAND2_X1 port map( A1 => n16491, A2 => n15564, ZN => n16489);
   U18787 : NOR2_X1 port map( A1 => n16489, A2 => n16232, ZN => n15760);
   U18791 : NOR2_X1 port map( A1 => n16312, A2 => n15556, ZN => n16315);
   U18792 : INV_X1 port map( A => n16809, ZN => n17481);
   U18793 : NAND2_X1 port map( A1 => n16030, A2 => n16273, ZN => n15769);
   U18794 : MUX2_X1 port map( A => n15770, B => n15769, S => n16274, Z => 
                           n16810);
   U18795 : INV_X1 port map( A => n15771, ZN => n15772);
   U18796 : NAND2_X1 port map( A1 => n15772, A2 => n16029, ZN => n16808);
   U18797 : INV_X1 port map( A => n17076, ZN => n16588);
   U18798 : NAND3_X1 port map( A1 => n16302, A2 => n16022, A3 => n16023, ZN => 
                           n15775);
   U18799 : NAND3_X1 port map( A1 => n16220, A2 => n15921, A3 => n16221, ZN => 
                           n15778);
   U18800 : NAND2_X1 port map( A1 => n5269, A2 => n16465, ZN => n15777);
   U18801 : INV_X1 port map( A => n15780, ZN => n15781);
   U18802 : NOR2_X1 port map( A1 => n15781, A2 => n16102, ZN => n15787);
   U18803 : MUX2_X1 port map( A => n4678, B => n15854, S => n24586, Z => n15785
                           );
   U18804 : NOR2_X1 port map( A1 => n17134, A2 => n3458, ZN => n15809);
   U18805 : NOR2_X1 port map( A1 => n16038, A2 => n24429, ZN => n15786);
   U18806 : AOI22_X1 port map( A1 => n15788, A2 => n24430, B1 => n15786, B2 => 
                           n2251, ZN => n16576);
   U18807 : INV_X1 port map( A => n15787, ZN => n15793);
   U18808 : INV_X1 port map( A => n15788, ZN => n15792);
   U18809 : AOI21_X1 port map( B1 => n291, B2 => n15790, A => n15789, ZN => 
                           n15791);
   U18810 : NAND3_X1 port map( A1 => n16576, A2 => n15793, A3 => n16575, ZN => 
                           n15797);
   U18811 : OAI21_X1 port map( B1 => n15798, B2 => n15797, A => n17131, ZN => 
                           n15808);
   U18812 : NAND2_X1 port map( A1 => n25245, A2 => n17130, ZN => n15803);
   U18813 : XNOR2_X1 port map( A => n18289, B => n18301, ZN => n17911);
   U18814 : XNOR2_X1 port map( A => n15810, B => n17911, ZN => n15879);
   U18816 : NAND2_X1 port map( A1 => n15814, A2 => n16204, ZN => n15815);
   U18817 : NAND2_X1 port map( A1 => n15905, A2 => n17183, ZN => n16366);
   U18821 : NOR2_X1 port map( A1 => n16170, A2 => n244, ZN => n15819);
   U18823 : NOR2_X1 port map( A1 => n15890, A2 => n24587, ZN => n15823);
   U18824 : OAI21_X1 port map( B1 => n15824, B2 => n15823, A => n24080, ZN => 
                           n15827);
   U18825 : INV_X1 port map( A => n16427, ZN => n15825);
   U18826 : OAI21_X1 port map( B1 => n16422, B2 => n707, A => n15825, ZN => 
                           n15826);
   U18827 : NAND2_X1 port map( A1 => n15826, A2 => n16170, ZN => n15836);
   U18828 : AND4_X1 port map( A1 => n15835, A2 => n16598, A3 => n15827, A4 => 
                           n15836, ZN => n15834);
   U18829 : NOR2_X1 port map( A1 => n16188, A2 => n15970, ZN => n15829);
   U18830 : NAND2_X1 port map( A1 => n16400, A2 => n15970, ZN => n15831);
   U18831 : NAND3_X1 port map( A1 => n16188, A2 => n15972, A3 => n16397, ZN => 
                           n15830);
   U18832 : NAND2_X1 port map( A1 => n15831, A2 => n15830, ZN => n15832);
   U18833 : INV_X1 port map( A => n17729, ZN => n17735);
   U18834 : NOR2_X1 port map( A1 => n15837, A2 => n16177, ZN => n15838);
   U18835 : NOR3_X1 port map( A1 => n15839, A2 => n4045, A3 => n15838, ZN => 
                           n15840);
   U18837 : MUX2_X1 port map( A => n15844, B => n24654, S => n16122, Z => 
                           n15845);
   U18838 : INV_X1 port map( A => n15847, ZN => n15853);
   U18839 : NOR2_X1 port map( A1 => n16391, A2 => n15849, ZN => n16390);
   U18840 : NAND2_X1 port map( A1 => n15848, A2 => n16162, ZN => n15851);
   U18841 : INV_X1 port map( A => n15849, ZN => n16392);
   U18842 : AOI22_X2 port map( A1 => n15852, A2 => n15853, B1 => n15851, B2 => 
                           n15850, ZN => n17118);
   U18843 : INV_X1 port map( A => n17118, ZN => n17100);
   U18844 : INV_X1 port map( A => n17120, ZN => n17115);
   U18845 : OAI21_X1 port map( B1 => n890, B2 => n17100, A => n17115, ZN => 
                           n15870);
   U18846 : NOR2_X1 port map( A1 => n16114, A2 => n16118, ZN => n15859);
   U18850 : INV_X1 port map( A => n15625, ZN => n16148);
   U18851 : NAND2_X1 port map( A1 => n16409, A2 => n16412, ZN => n15865);
   U18852 : NAND2_X1 port map( A1 => n15984, A2 => n16414, ZN => n15867);
   U18853 : NOR3_X1 port map( A1 => n17088, A2 => n17086, A3 => n16578, ZN => 
                           n15874);
   U18854 : AOI21_X1 port map( B1 => n15875, B2 => n17087, A => n15874, ZN => 
                           n15876);
   U18855 : XNOR2_X1 port map( A => n18294, B => n20744, ZN => n15877);
   U18856 : XNOR2_X1 port map( A => n18305, B => n15877, ZN => n15878);
   U18857 : NAND2_X1 port map( A1 => n25031, A2 => n16929, ZN => n15884);
   U18858 : AOI21_X1 port map( B1 => n17060, B2 => n17059, A => n17054, ZN => 
                           n15881);
   U18859 : OAI22_X1 port map( A1 => n15881, A2 => n15880, B1 => n15883, B2 => 
                           n17060, ZN => n15882);
   U18860 : NAND2_X1 port map( A1 => n15885, A2 => n24467, ZN => n15886);
   U18861 : NAND3_X1 port map( A1 => n15888, A2 => n15886, A3 => n15887, ZN => 
                           n15892);
   U18862 : NAND3_X1 port map( A1 => n15890, A2 => n25432, A3 => n24467, ZN => 
                           n15891);
   U18863 : NAND2_X1 port map( A1 => n15894, A2 => n16360, ZN => n15898);
   U18864 : NAND3_X1 port map( A1 => n24841, A2 => n24456, A3 => n15894, ZN => 
                           n15896);
   U18865 : OAI211_X1 port map( C1 => n24919, C2 => n15898, A => n15897, B => 
                           n15896, ZN => n16770);
   U18866 : AOI21_X1 port map( B1 => n16196, B2 => n16328, A => n15899, ZN => 
                           n15903);
   U18867 : NAND2_X1 port map( A1 => n15901, A2 => n15900, ZN => n15902);
   U18869 : NAND3_X1 port map( A1 => n16368, A2 => n15904, A3 => n16204, ZN => 
                           n15911);
   U18870 : NOR2_X1 port map( A1 => n16367, A2 => n16206, ZN => n15906);
   U18871 : NAND2_X1 port map( A1 => n15906, A2 => n17180, ZN => n15909);
   U18872 : NAND3_X1 port map( A1 => n15907, A2 => n17183, A3 => n16367, ZN => 
                           n15908);
   U18873 : NAND4_X1 port map( A1 => n15911, A2 => n15910, A3 => n15909, A4 => 
                           n15908, ZN => n16989);
   U18874 : NAND2_X1 port map( A1 => n16406, A2 => n24061, ZN => n16402);
   U18875 : NAND2_X1 port map( A1 => n15646, A2 => n25500, ZN => n15912);
   U18876 : NAND3_X1 port map( A1 => n16406, A2 => n15646, A3 => n16403, ZN => 
                           n15913);
   U18877 : MUX2_X1 port map( A => n25455, B => n16334, S => n1123, Z => n15914
                           );
   U18878 : NAND2_X1 port map( A1 => n15914, A2 => n267, ZN => n15919);
   U18880 : NAND2_X1 port map( A1 => n17364, A2 => n25214, ZN => n15920);
   U18881 : INV_X1 port map( A => n16989, ZN => n17362);
   U18882 : NOR2_X1 port map( A1 => n16220, A2 => n16221, ZN => n15924);
   U18883 : NOR2_X1 port map( A1 => n15921, A2 => n16219, ZN => n15923);
   U18884 : INV_X1 port map( A => n15922, ZN => n16462);
   U18885 : MUX2_X1 port map( A => n15924, B => n15923, S => n16462, Z => 
                           n15927);
   U18886 : OAI22_X1 port map( A1 => n15925, A2 => n16461, B1 => n16216, B2 => 
                           n16465, ZN => n15926);
   U18887 : NOR2_X2 port map( A1 => n15927, A2 => n15926, ZN => n17048);
   U18888 : MUX2_X1 port map( A => n16447, B => n257, S => n16449, Z => n15931)
                           ;
   U18889 : NAND2_X1 port map( A1 => n16235, A2 => n16451, ZN => n15928);
   U18890 : MUX2_X1 port map( A => n15929, B => n15928, S => n16449, Z => 
                           n15930);
   U18891 : INV_X1 port map( A => n16231, ZN => n16494);
   U18892 : INV_X1 port map( A => n16230, ZN => n16492);
   U18893 : MUX2_X1 port map( A => n15935, B => n15934, S => n16492, Z => 
                           n15936);
   U18894 : INV_X1 port map( A => n15938, ZN => n16252);
   U18895 : NOR2_X1 port map( A1 => n16252, A2 => n15762, ZN => n15939);
   U18896 : AOI22_X1 port map( A1 => n15939, A2 => n16016, B1 => n16246, B2 => 
                           n16252, ZN => n15942);
   U18897 : INV_X1 port map( A => n17048, ZN => n16628);
   U18898 : OAI211_X1 port map( C1 => n15943, C2 => n15946, A => n16438, B => 
                           n16242, ZN => n15949);
   U18899 : NAND3_X1 port map( A1 => n16442, A2 => n15945, A3 => n15944, ZN => 
                           n15948);
   U18900 : MUX2_X1 port map( A => n15951, B => n15950, S => n15953, Z => 
                           n15955);
   U18901 : NAND2_X1 port map( A1 => n15952, A2 => n24981, ZN => n15954);
   U18902 : AOI22_X1 port map( A1 => n15956, A2 => n372, B1 => n17049, B2 => 
                           n16628, ZN => n15957);
   U18903 : NOR2_X1 port map( A1 => n1329, A2 => n16427, ZN => n15959);
   U18904 : MUX2_X1 port map( A => n15960, B => n15959, S => n15958, Z => 
                           n15964);
   U18905 : NOR2_X1 port map( A1 => n15962, A2 => n16422, ZN => n15963);
   U18906 : OAI21_X1 port map( B1 => n16156, B2 => n16122, A => n15965, ZN => 
                           n15966);
   U18907 : NAND2_X1 port map( A1 => n15966, A2 => n16155, ZN => n15969);
   U18908 : OAI21_X1 port map( B1 => n24459, B2 => n2996, A => n16125, ZN => 
                           n15967);
   U18909 : NAND2_X1 port map( A1 => n15967, A2 => n16156, ZN => n15968);
   U18911 : AOI21_X1 port map( B1 => n15971, B2 => n16399, A => n3630, ZN => 
                           n15975);
   U18912 : NAND2_X1 port map( A1 => n15973, A2 => n15972, ZN => n15974);
   U18913 : INV_X1 port map( A => n16391, ZN => n15978);
   U18914 : NAND2_X1 port map( A1 => n15978, A2 => n15977, ZN => n15983);
   U18915 : NAND2_X1 port map( A1 => n16391, A2 => n15849, ZN => n15979);
   U18916 : NAND2_X1 port map( A1 => n15980, A2 => n15979, ZN => n15981);
   U18917 : NAND3_X1 port map( A1 => n16394, A2 => n16162, A3 => n16389, ZN => 
                           n15982);
   U18918 : INV_X1 port map( A => n17042, ZN => n16998);
   U18919 : NAND2_X1 port map( A1 => n16418, A2 => n15984, ZN => n15989);
   U18920 : NAND2_X1 port map( A1 => n16408, A2 => n16412, ZN => n15985);
   U18921 : OAI211_X1 port map( C1 => n16412, C2 => n16409, A => n16413, B => 
                           n15985, ZN => n15988);
   U18922 : NOR2_X1 port map( A1 => n16141, A2 => n16408, ZN => n15987);
   U18924 : INV_X1 port map( A => n15992, ZN => n15993);
   U18925 : AND2_X1 port map( A1 => n15990, A2 => n25210, ZN => n15991);
   U18926 : NAND2_X1 port map( A1 => n15994, A2 => n16997, ZN => n15997);
   U18927 : OAI21_X1 port map( B1 => n16998, B2 => n374, A => n15995, ZN => 
                           n15996);
   U18928 : XNOR2_X1 port map( A => n18557, B => n18312, ZN => n15999);
   U18929 : XNOR2_X1 port map( A => n15999, B => n16000, ZN => n16093);
   U18930 : NAND2_X1 port map( A1 => n16001, A2 => n16268, ZN => n16007);
   U18931 : NOR2_X1 port map( A1 => n16002, A2 => n25009, ZN => n16003);
   U18932 : NAND2_X1 port map( A1 => n16266, A2 => n16003, ZN => n16006);
   U18933 : MUX2_X1 port map( A => n3554, B => n16309, S => n15556, Z => n16013
                           );
   U18934 : OAI22_X1 port map( A1 => n16638, A2 => n16010, B1 => n16309, B2 => 
                           n16009, ZN => n16011);
   U18935 : INV_X1 port map( A => n25406, ZN => n16844);
   U18936 : OAI21_X1 port map( B1 => n16342, B2 => n16285, A => n16286, ZN => 
                           n16014);
   U18937 : NAND2_X1 port map( A1 => n16247, A2 => n16016, ZN => n16017);
   U18938 : OAI21_X1 port map( B1 => n16253, B2 => n25284, A => n16017, ZN => 
                           n16019);
   U18939 : NAND2_X1 port map( A1 => n16019, A2 => n15762, ZN => n16020);
   U18940 : OAI22_X1 port map( A1 => n16226, A2 => n16023, B1 => n16225, B2 => 
                           n16022, ZN => n16228);
   U18941 : INV_X1 port map( A => n16024, ZN => n16026);
   U18942 : NAND2_X1 port map( A1 => n16277, A2 => n16029, ZN => n16031);
   U18943 : INV_X1 port map( A => n16032, ZN => n16033);
   U18944 : NOR2_X1 port map( A1 => n17067, A2 => n369, ZN => n16035);
   U18945 : OAI21_X1 port map( B1 => n16546, B2 => n17069, A => n17067, ZN => 
                           n16036);
   U18946 : INV_X1 port map( A => n16546, ZN => n16612);
   U18947 : INV_X1 port map( A => n16041, ZN => n16046);
   U18948 : NAND2_X1 port map( A1 => n16043, A2 => n16042, ZN => n16045);
   U18949 : INV_X1 port map( A => n16260, ZN => n16533);
   U18950 : MUX2_X1 port map( A => n16048, B => n294, S => n24352, Z => n16049)
                           ;
   U18951 : NAND2_X1 port map( A1 => n16049, A2 => n16509, ZN => n16055);
   U18952 : NOR2_X1 port map( A1 => n16050, A2 => n16508, ZN => n16052);
   U18954 : OAI21_X1 port map( B1 => n24551, B2 => n16469, A => n16057, ZN => 
                           n16058);
   U18956 : INV_X1 port map( A => n16060, ZN => n16061);
   U18957 : NOR2_X1 port map( A1 => n16062, A2 => n16061, ZN => n16066);
   U18958 : MUX2_X1 port map( A => n16066, B => n16065, S => n16064, Z => 
                           n16071);
   U18960 : NAND2_X1 port map( A1 => n16129, A2 => n16076, ZN => n16072);
   U18963 : NOR2_X1 port map( A1 => n16077, A2 => n16076, ZN => n16078);
   U18964 : OAI21_X1 port map( B1 => n1365, B2 => n16075, A => n16078, ZN => 
                           n17157);
   U18965 : INV_X1 port map( A => n17164, ZN => n16262);
   U18967 : INV_X1 port map( A => n16082, ZN => n16083);
   U18968 : NAND2_X1 port map( A1 => n16083, A2 => n16100, ZN => n16087);
   U18969 : NAND3_X1 port map( A1 => n16085, A2 => n16101, A3 => n16084, ZN => 
                           n16086);
   U18970 : OAI21_X1 port map( B1 => n16375, B2 => n25219, A => n17166, ZN => 
                           n16089);
   U18971 : XNOR2_X1 port map( A => n18375, B => n23883, ZN => n16090);
   U18972 : XNOR2_X1 port map( A => n16091, B => n16090, ZN => n16092);
   U18973 : NOR2_X1 port map( A1 => n15625, A2 => n16096, ZN => n16094);
   U18974 : OAI21_X1 port map( B1 => n16151, B2 => n16095, A => n16094, ZN => 
                           n16098);
   U18975 : NOR2_X1 port map( A1 => n16114, A2 => n16113, ZN => n16115);
   U18976 : NAND2_X1 port map( A1 => n16123, A2 => n25449, ZN => n16128);
   U18977 : INV_X1 port map( A => n24459, ZN => n16124);
   U18978 : NOR2_X1 port map( A1 => n16155, A2 => n2996, ZN => n16126);
   U18979 : AOI21_X1 port map( B1 => n16130, B2 => n16129, A => n24826, ZN => 
                           n16132);
   U18980 : MUX2_X1 port map( A => n16134, B => n16432, S => n17174, Z => 
                           n16135);
   U18981 : INV_X1 port map( A => n16780, ZN => n17348);
   U18982 : INV_X1 port map( A => n17342, ZN => n17242);
   U18984 : OAI21_X1 port map( B1 => n16778, B2 => n17346, A => n16136, ZN => 
                           n16137);
   U18985 : NOR2_X1 port map( A1 => n16777, A2 => n16137, ZN => n16138);
   U18987 : XNOR2_X1 port map( A => n25077, B => n18277, ZN => n16215);
   U18989 : NOR2_X1 port map( A1 => n16418, A2 => n16141, ZN => n16411);
   U18990 : NOR2_X1 port map( A1 => n16413, A2 => n16417, ZN => n16142);
   U18991 : NOR2_X1 port map( A1 => n16411, A2 => n16142, ZN => n16143);
   U18992 : OAI21_X1 port map( B1 => n16148, B2 => n4418, A => n16147, ZN => 
                           n16150);
   U18993 : AOI22_X1 port map( A1 => n16152, A2 => n16151, B1 => n16150, B2 => 
                           n213, ZN => n16660);
   U18994 : NOR2_X1 port map( A1 => n17399, A2 => n17031, ZN => n17397);
   U18995 : INV_X1 port map( A => n17397, ZN => n16182);
   U18998 : NAND2_X1 port map( A1 => n381, A2 => n2996, ZN => n16157);
   U18999 : MUX2_X1 port map( A => n16158, B => n16157, S => n16156, Z => 
                           n16159);
   U19001 : INV_X1 port map( A => n17395, ZN => n17196);
   U19002 : MUX2_X1 port map( A => n16163, B => n16162, S => n16392, Z => 
                           n16168);
   U19003 : INV_X1 port map( A => n16161, ZN => n16165);
   U19004 : AND3_X1 port map( A1 => n16163, A2 => n16391, A3 => n16162, ZN => 
                           n16164);
   U19005 : AOI21_X1 port map( B1 => n16165, B2 => n16167, A => n16164, ZN => 
                           n16166);
   U19006 : NAND2_X1 port map( A1 => n16169, A2 => n244, ZN => n16173);
   U19007 : NAND2_X1 port map( A1 => n16383, A2 => n16381, ZN => n16179);
   U19008 : NOR3_X1 port map( A1 => n4046, A2 => n16177, A3 => n16381, ZN => 
                           n16178);
   U19009 : NOR2_X1 port map( A1 => n17400, A2 => n17192, ZN => n17396);
   U19010 : NAND2_X1 port map( A1 => n17396, A2 => n17031, ZN => n16181);
   U19011 : NAND2_X1 port map( A1 => n16339, A2 => n16183, ZN => n16184);
   U19012 : NAND2_X1 port map( A1 => n16187, A2 => n16186, ZN => n16189);
   U19013 : NAND2_X1 port map( A1 => n16189, A2 => n16188, ZN => n16190);
   U19014 : INV_X1 port map( A => n17185, ZN => n16203);
   U19015 : NOR2_X1 port map( A1 => n16192, A2 => n16191, ZN => n16327);
   U19016 : NOR2_X1 port map( A1 => n16324, A2 => n16193, ZN => n16195);
   U19017 : NAND2_X1 port map( A1 => n16203, A2 => n17391, ZN => n16214);
   U19018 : NAND3_X1 port map( A1 => n3544, A2 => n16401, A3 => n25500, ZN => 
                           n16201);
   U19019 : MUX2_X1 port map( A => n16205, B => n17182, S => n16204, Z => 
                           n16210);
   U19020 : INV_X1 port map( A => n16366, ZN => n16209);
   U19021 : NOR2_X1 port map( A1 => n17180, A2 => n16206, ZN => n16208);
   U19022 : INV_X1 port map( A => n17387, ZN => n17186);
   U19024 : NAND2_X1 port map( A1 => n16349, A2 => n16597, ZN => n16211);
   U19025 : NAND2_X1 port map( A1 => n17389, A2 => n17185, ZN => n16212);
   U19026 : XNOR2_X1 port map( A => n17863, B => n18549, ZN => n18342);
   U19027 : XNOR2_X1 port map( A => n18342, B => n16215, ZN => n16322);
   U19028 : INV_X1 port map( A => n16216, ZN => n16218);
   U19029 : MUX2_X1 port map( A => n16218, B => n16217, S => n16462, Z => 
                           n16223);
   U19030 : NOR2_X2 port map( A1 => n16223, A2 => n16222, ZN => n17212);
   U19031 : OAI21_X1 port map( B1 => n16302, B2 => n16225, A => n16224, ZN => 
                           n16227);
   U19032 : NOR2_X1 port map( A1 => n16231, A2 => n16230, ZN => n16233);
   U19033 : OAI211_X1 port map( C1 => n16235, C2 => n385, A => n16450, B => 
                           n16447, ZN => n16238);
   U19034 : INV_X1 port map( A => n16447, ZN => n16236);
   U19035 : INV_X1 port map( A => n17017, ZN => n16240);
   U19036 : OAI22_X1 port map( A1 => n2636, A2 => n16442, B1 => n16443, B2 => 
                           n16242, ZN => n16244);
   U19037 : NAND2_X1 port map( A1 => n16244, A2 => n16243, ZN => n16245);
   U19038 : NOR2_X1 port map( A1 => n16246, A2 => n15762, ZN => n16250);
   U19043 : XNOR2_X1 port map( A => n24384, B => n3164, ZN => n16320);
   U19044 : NAND2_X1 port map( A1 => n16375, A2 => n25219, ZN => n16532);
   U19046 : INV_X1 port map( A => n25219, ZN => n17160);
   U19047 : INV_X1 port map( A => n17824, ZN => n18006);
   U19048 : AOI21_X1 port map( B1 => n25009, B2 => n16268, A => n16266, ZN => 
                           n16271);
   U19050 : NAND3_X1 port map( A1 => n16277, A2 => n16276, A3 => n24403, ZN => 
                           n16278);
   U19051 : INV_X1 port map( A => n16345, ZN => n16281);
   U19052 : NOR2_X1 port map( A1 => n16281, A2 => n24540, ZN => n16283);
   U19053 : OAI21_X1 port map( B1 => n16286, B2 => n16285, A => n24540, ZN => 
                           n16287);
   U19054 : NOR2_X1 port map( A1 => n16347, A2 => n16287, ZN => n16288);
   U19057 : INV_X1 port map( A => n16363, ZN => n16295);
   U19058 : NOR2_X1 port map( A1 => n16293, A2 => n25546, ZN => n16294);
   U19059 : OAI21_X1 port map( B1 => n16295, B2 => n16294, A => n16357, ZN => 
                           n16296);
   U19061 : INV_X1 port map( A => n16298, ZN => n16300);
   U19062 : NAND2_X1 port map( A1 => n16302, A2 => n16301, ZN => n16306);
   U19063 : MUX2_X1 port map( A => n16306, B => n16305, S => n16304, Z => 
                           n16307);
   U19064 : AOI21_X1 port map( B1 => n16311, B2 => n15557, A => n3554, ZN => 
                           n16310);
   U19065 : XNOR2_X1 port map( A => n18646, B => n18006, ZN => n16319);
   U19066 : XNOR2_X1 port map( A => n16320, B => n16319, ZN => n16321);
   U19067 : XNOR2_X1 port map( A => n16321, B => n16322, ZN => n19132);
   U19068 : NOR2_X1 port map( A1 => n25323, A2 => n16324, ZN => n16326);
   U19069 : NOR2_X1 port map( A1 => n16327, A2 => n16326, ZN => n16329);
   U19070 : OAI21_X1 port map( B1 => n3947, B2 => n16332, A => n25455, ZN => 
                           n16340);
   U19075 : NOR2_X2 port map( A1 => n16348, A2 => n16347, ZN => n17455);
   U19076 : INV_X1 port map( A => n17455, ZN => n16354);
   U19077 : NAND2_X1 port map( A1 => n24890, A2 => n24467, ZN => n16353);
   U19078 : OAI21_X1 port map( B1 => n15822, B2 => n16349, A => n16595, ZN => 
                           n16351);
   U19079 : OAI21_X1 port map( B1 => n16357, B2 => n24456, A => n16355, ZN => 
                           n16362);
   U19081 : MUX2_X1 port map( A => n16362, B => n16361, S => n16360, Z => 
                           n16364);
   U19086 : AND2_X1 port map( A1 => n17297, A2 => n17296, ZN => n16371);
   U19087 : NAND2_X1 port map( A1 => n17299, A2 => n17297, ZN => n16372);
   U19090 : XNOR2_X1 port map( A => n18532, B => n18610, ZN => n16380);
   U19091 : INV_X1 port map( A => n16375, ZN => n16838);
   U19092 : NAND3_X1 port map( A1 => n17163, A2 => n17160, A3 => n16838, ZN => 
                           n16377);
   U19093 : NAND2_X1 port map( A1 => n16533, A2 => n17166, ZN => n16376);
   U19094 : OAI211_X2 port map( C1 => n16378, C2 => n17164, A => n16377, B => 
                           n16376, ZN => n18270);
   U19095 : XNOR2_X1 port map( A => n18270, B => n1951, ZN => n16379);
   U19096 : XNOR2_X1 port map( A => n16380, B => n16379, ZN => n16503);
   U19097 : NOR2_X1 port map( A1 => n16383, A2 => n16382, ZN => n16384);
   U19098 : NOR2_X1 port map( A1 => n16385, A2 => n16384, ZN => n16386);
   U19099 : OAI21_X1 port map( B1 => n16390, B2 => n5758, A => n16389, ZN => 
                           n16396);
   U19100 : AOI21_X1 port map( B1 => n16393, B2 => n16392, A => n16391, ZN => 
                           n16395);
   U19101 : INV_X1 port map( A => n16400, ZN => n17433);
   U19102 : INV_X1 port map( A => n17439, ZN => n16828);
   U19103 : AOI21_X1 port map( B1 => n16402, B2 => n16401, A => n16404, ZN => 
                           n16407);
   U19104 : NOR2_X1 port map( A1 => n16409, A2 => n16408, ZN => n16410);
   U19105 : NOR2_X1 port map( A1 => n16413, A2 => n16412, ZN => n16415);
   U19106 : NAND2_X1 port map( A1 => n16417, A2 => n16416, ZN => n16419);
   U19107 : NOR2_X1 port map( A1 => n16419, A2 => n16418, ZN => n16420);
   U19110 : INV_X1 port map( A => n17442, ZN => n16964);
   U19111 : INV_X1 port map( A => n16432, ZN => n16433);
   U19112 : AOI21_X1 port map( B1 => n17171, B2 => n17522, A => n16433, ZN => 
                           n16436);
   U19113 : XNOR2_X1 port map( A => n24565, B => n18335, ZN => n18101);
   U19114 : AOI21_X1 port map( B1 => n16438, B2 => n16437, A => n16442, ZN => 
                           n16439);
   U19115 : NAND2_X1 port map( A1 => n16441, A2 => n16440, ZN => n16445);
   U19116 : MUX2_X1 port map( A => n385, B => n16448, S => n16447, Z => n16457)
                           ;
   U19117 : NAND2_X1 port map( A1 => n16450, A2 => n16449, ZN => n16455);
   U19118 : NAND2_X1 port map( A1 => n385, A2 => n257, ZN => n16453);
   U19119 : OAI22_X1 port map( A1 => n16455, A2 => n223, B1 => n16453, B2 => 
                           n16452, ZN => n16456);
   U19120 : INV_X1 port map( A => n16849, ZN => n17139);
   U19121 : AND2_X1 port map( A1 => n17144, A2 => n17139, ZN => n16488);
   U19123 : NOR2_X1 port map( A1 => n5269, A2 => n16464, ZN => n16467);
   U19124 : OAI21_X1 port map( B1 => n16467, B2 => n16466, A => n16465, ZN => 
                           n16468);
   U19125 : INV_X1 port map( A => n16984, ZN => n17140);
   U19126 : MUX2_X1 port map( A => n16471, B => n24550, S => n16469, Z => 
                           n16479);
   U19127 : OAI21_X1 port map( B1 => n16474, B2 => n16473, A => n16472, ZN => 
                           n16478);
   U19128 : NOR2_X1 port map( A1 => n16476, A2 => n16475, ZN => n16477);
   U19129 : INV_X1 port map( A => n16851, ZN => n17137);
   U19130 : NOR2_X1 port map( A1 => n17140, A2 => n17137, ZN => n16487);
   U19131 : NAND2_X1 port map( A1 => n16485, A2 => n16484, ZN => n16515);
   U19132 : NAND2_X1 port map( A1 => n16486, A2 => n16515, ZN => n17141);
   U19134 : NAND2_X1 port map( A1 => n16490, A2 => n16489, ZN => n16495);
   U19135 : NAND2_X1 port map( A1 => n17138, A2 => n16984, ZN => n16691);
   U19136 : NAND3_X1 port map( A1 => n16991, A2 => n287, A3 => n16499, ZN => 
                           n16501);
   U19137 : OAI21_X1 port map( B1 => n16021, B2 => n17461, A => n16991, ZN => 
                           n16500);
   U19138 : XNOR2_X1 port map( A => n17581, B => n18331, ZN => n17722);
   U19139 : XNOR2_X1 port map( A => n18101, B => n17722, ZN => n16502);
   U19140 : MUX2_X2 port map( A => n16505, B => n16504, S => n24324, Z => 
                           n20670);
   U19141 : OAI21_X1 port map( B1 => n17467, B2 => n25572, A => n16506, ZN => 
                           n16507);
   U19142 : INV_X1 port map( A => n17041, ZN => n18700);
   U19143 : NAND2_X1 port map( A1 => n16511, A2 => n16510, ZN => n16512);
   U19144 : MUX2_X1 port map( A => n16512, B => n17297, S => n17299, Z => 
                           n16514);
   U19145 : XNOR2_X1 port map( A => n18700, B => n18214, ZN => n16521);
   U19146 : NAND2_X1 port map( A1 => n16515, A2 => n17138, ZN => n16517);
   U19147 : OAI21_X1 port map( B1 => n16518, B2 => n16517, A => n16848, ZN => 
                           n16519);
   U19148 : XNOR2_X1 port map( A => n18605, B => n1797, ZN => n16520);
   U19149 : XNOR2_X1 port map( A => n16521, B => n16520, ZN => n16538);
   U19150 : AOI22_X1 port map( A1 => n16523, A2 => n17522, B1 => n16522, B2 => 
                           n17175, ZN => n16525);
   U19151 : NOR2_X1 port map( A1 => n17522, A2 => n17171, ZN => n16524);
   U19152 : MUX2_X1 port map( A => n16525, B => n16863, S => n16524, Z => 
                           n17900);
   U19153 : NOR2_X1 port map( A1 => n16526, A2 => n16980, ZN => n16530);
   U19154 : INV_X1 port map( A => n16527, ZN => n17451);
   U19155 : NOR2_X1 port map( A1 => n17455, A2 => n17450, ZN => n16528);
   U19156 : INV_X1 port map( A => n16532, ZN => n16534);
   U19157 : MUX2_X1 port map( A => n17166, B => n17163, S => n25218, Z => 
                           n16535);
   U19158 : XNOR2_X1 port map( A => n18420, B => n18451, ZN => n17974);
   U19159 : XNOR2_X1 port map( A => n17974, B => n18348, ZN => n16537);
   U19160 : XNOR2_X1 port map( A => n16537, B => n16538, ZN => n18749);
   U19161 : AOI21_X1 port map( B1 => n17474, B2 => n17473, A => n17472, ZN => 
                           n16542);
   U19162 : OAI22_X1 port map( A1 => n16540, A2 => n17633, B1 => n16901, B2 => 
                           n16902, ZN => n16541);
   U19163 : NAND2_X1 port map( A1 => n17288, A2 => n17229, ZN => n17539);
   U19164 : NAND2_X1 port map( A1 => n17540, A2 => n17539, ZN => n16755);
   U19165 : NAND2_X1 port map( A1 => n17288, A2 => n17283, ZN => n16543);
   U19166 : AOI21_X1 port map( B1 => n16543, B2 => n17229, A => n17293, ZN => 
                           n16544);
   U19167 : XNOR2_X1 port map( A => n18659, B => n17993, ZN => n18359);
   U19168 : INV_X1 port map( A => n18359, ZN => n18529);
   U19169 : INV_X1 port map( A => n17919, ZN => n16555);
   U19170 : AOI21_X1 port map( B1 => n16796, B2 => n16794, A => n5375, ZN => 
                           n16554);
   U19171 : NOR2_X1 port map( A1 => n16550, A2 => n16547, ZN => n16548);
   U19172 : NAND2_X1 port map( A1 => n16549, A2 => n16548, ZN => n16553);
   U19173 : XNOR2_X1 port map( A => n17680, B => n16555, ZN => n16937);
   U19174 : XNOR2_X1 port map( A => n18529, B => n16937, ZN => n16571);
   U19176 : OAI21_X1 port map( B1 => n17216, B2 => n17207, A => n17015, ZN => 
                           n16558);
   U19177 : NAND2_X1 port map( A1 => n16558, A2 => n17212, ZN => n16559);
   U19178 : INV_X1 port map( A => n18102, ZN => n17649);
   U19179 : XNOR2_X1 port map( A => n17649, B => n2145, ZN => n16569);
   U19180 : NAND2_X1 port map( A1 => n16942, A2 => n16940, ZN => n16564);
   U19181 : INV_X1 port map( A => n16743, ZN => n16560);
   U19182 : AOI21_X1 port map( B1 => n17224, B2 => n17413, A => n16956, ZN => 
                           n16568);
   U19183 : INV_X1 port map( A => n17419, ZN => n16565);
   U19185 : NAND3_X1 port map( A1 => n16565, A2 => n17227, A3 => n25246, ZN => 
                           n16566);
   U19187 : XNOR2_X1 port map( A => n18269, B => n18530, ZN => n18405);
   U19188 : XNOR2_X1 port map( A => n18405, B => n16569, ZN => n16570);
   U19190 : NAND2_X1 port map( A1 => n18749, A2 => n24421, ZN => n19562);
   U19192 : NOR2_X1 port map( A1 => n16572, A2 => n17120, ZN => n16573);
   U19193 : MUX2_X1 port map( A => n17134, B => n25245, S => n17132, Z => 
                           n16577);
   U19194 : OAI21_X1 port map( B1 => n16649, B2 => n17086, A => n16740, ZN => 
                           n16581);
   U19195 : NAND2_X1 port map( A1 => n17086, A2 => n16578, ZN => n16579);
   U19196 : INV_X1 port map( A => n17086, ZN => n16648);
   U19197 : OAI22_X1 port map( A1 => n17084, A2 => n16579, B1 => n16648, B2 => 
                           n371, ZN => n16580);
   U19198 : XNOR2_X1 port map( A => n17970, B => n17881, ZN => n18246);
   U19199 : XNOR2_X1 port map( A => n18246, B => n16582, ZN => n16601);
   U19200 : AOI21_X1 port map( B1 => n16901, B2 => n17472, A => n17629, ZN => 
                           n16587);
   U19201 : NAND2_X1 port map( A1 => n17633, A2 => n16539, ZN => n16583);
   U19202 : OAI21_X1 port map( B1 => n2561, B2 => n17633, A => n16583, ZN => 
                           n16586);
   U19203 : INV_X1 port map( A => n17472, ZN => n16584);
   U19204 : NAND2_X1 port map( A1 => n16584, A2 => n17633, ZN => n16585);
   U19206 : INV_X1 port map( A => n17478, ZN => n17079);
   U19207 : NAND2_X1 port map( A1 => n17479, A2 => n17079, ZN => n16589);
   U19208 : AOI21_X1 port map( B1 => n16590, B2 => n16589, A => n16588, ZN => 
                           n16593);
   U19209 : NAND2_X1 port map( A1 => n17481, A2 => n17078, ZN => n16591);
   U19211 : XNOR2_X1 port map( A => n18685, B => n18042, ZN => n16599);
   U19212 : INV_X1 port map( A => n16888, ZN => n17730);
   U19213 : INV_X1 port map( A => n17734, ZN => n17731);
   U19214 : XNOR2_X1 port map( A => n16599, B => n18370, ZN => n18520);
   U19215 : INV_X1 port map( A => n17334, ZN => n16973);
   U19216 : INV_X1 port map( A => n16726, ZN => n16606);
   U19217 : INV_X1 port map( A => n17333, ZN => n16604);
   U19218 : NOR2_X1 port map( A1 => n17335, A2 => n16602, ZN => n16603);
   U19220 : AOI22_X1 port map( A1 => n17599, A2 => n17316, B1 => n17304, B2 => 
                           n16921, ZN => n16920);
   U19221 : INV_X1 port map( A => n17316, ZN => n16715);
   U19222 : NOR2_X1 port map( A1 => n17304, A2 => n24542, ZN => n16714);
   U19223 : OAI21_X1 port map( B1 => n3783, B2 => n17316, A => n16714, ZN => 
                           n16608);
   U19224 : OAI21_X1 port map( B1 => n16920, B2 => n16716, A => n16608, ZN => 
                           n17757);
   U19225 : XNOR2_X1 port map( A => n18220, B => n18431, ZN => n16625);
   U19226 : INV_X1 port map( A => n16619, ZN => n16621);
   U19227 : NAND2_X1 port map( A1 => n16622, A2 => n16795, ZN => n16798);
   U19228 : NAND2_X1 port map( A1 => n5762, A2 => n16798, ZN => n16623);
   U19229 : XNOR2_X1 port map( A => n17476, B => n1870, ZN => n16624);
   U19230 : XNOR2_X1 port map( A => n16625, B => n16624, ZN => n16626);
   U19231 : NAND2_X1 port map( A1 => n19560, A2 => n19559, ZN => n16666);
   U19232 : NOR2_X1 port map( A1 => n17216, A2 => n25201, ZN => n16878);
   U19233 : NOR2_X1 port map( A1 => n17185, A2 => n17179, ZN => n16627);
   U19234 : XNOR2_X1 port map( A => n17515, B => n18541, ZN => n18439);
   U19235 : MUX2_X1 port map( A => n17050, B => n16628, S => n17049, Z => 
                           n16634);
   U19236 : NAND3_X1 port map( A1 => n16775, A2 => n24570, A3 => n17053, ZN => 
                           n16632);
   U19237 : INV_X1 port map( A => n17049, ZN => n16629);
   U19238 : XNOR2_X1 port map( A => n18439, B => n16635, ZN => n16665);
   U19239 : INV_X1 port map( A => n17381, ZN => n17422);
   U19240 : NOR2_X1 port map( A1 => n17379, A2 => n17422, ZN => n16637);
   U19241 : INV_X1 port map( A => n17425, ZN => n17382);
   U19242 : NOR2_X1 port map( A1 => n17382, A2 => n5409, ZN => n16636);
   U19243 : MUX2_X1 port map( A => n16637, B => n16636, S => n24330, Z => 
                           n16646);
   U19244 : NAND2_X1 port map( A1 => n16639, A2 => n16638, ZN => n16640);
   U19245 : NAND2_X1 port map( A1 => n16641, A2 => n16640, ZN => n17423);
   U19246 : INV_X1 port map( A => n17423, ZN => n16642);
   U19247 : NAND2_X1 port map( A1 => n17382, A2 => n16642, ZN => n16643);
   U19248 : AOI21_X1 port map( B1 => n16644, B2 => n16643, A => n5406, ZN => 
                           n16645);
   U19249 : NOR2_X2 port map( A1 => n16646, A2 => n16645, ZN => n18666);
   U19250 : INV_X1 port map( A => n16647, ZN => n16652);
   U19251 : NAND2_X1 port map( A1 => n16650, A2 => n16739, ZN => n16651);
   U19252 : NAND2_X1 port map( A1 => n17132, A2 => n16655, ZN => n16658);
   U19253 : NOR2_X1 port map( A1 => n25227, A2 => n3458, ZN => n16654);
   U19254 : NAND2_X1 port map( A1 => n17134, A2 => n16654, ZN => n16657);
   U19255 : OAI211_X1 port map( C1 => n17134, C2 => n16658, A => n16657, B => 
                           n16656, ZN => n16910);
   U19256 : INV_X1 port map( A => n16910, ZN => n16663);
   U19257 : NAND2_X1 port map( A1 => n17399, A2 => n17395, ZN => n16659);
   U19258 : NAND2_X1 port map( A1 => n16659, A2 => n17031, ZN => n17030);
   U19260 : NAND2_X1 port map( A1 => n17400, A2 => n17028, ZN => n16661);
   U19261 : XNOR2_X1 port map( A => n16663, B => n17840, ZN => n18381);
   U19262 : AOI21_X1 port map( B1 => n19562, B2 => n16666, A => n19555, ZN => 
                           n16701);
   U19263 : NAND2_X1 port map( A1 => n17347, A2 => n17346, ZN => n16668);
   U19264 : NAND3_X1 port map( A1 => n17241, A2 => n17343, A3 => n17236, ZN => 
                           n16667);
   U19265 : OAI21_X1 port map( B1 => n16668, B2 => n17348, A => n16667, ZN => 
                           n17206);
   U19266 : NOR2_X2 port map( A1 => n16669, A2 => n17206, ZN => n18227);
   U19267 : OAI21_X1 port map( B1 => n17051, B2 => n17050, A => n17053, ZN => 
                           n16670);
   U19268 : MUX2_X1 port map( A => n25214, B => n25058, S => n17039, Z => 
                           n16988);
   U19269 : NOR3_X1 port map( A1 => n16770, A2 => n25058, A3 => n25214, ZN => 
                           n16671);
   U19270 : NAND2_X1 port map( A1 => n266, A2 => n17351, ZN => n16672);
   U19271 : NAND2_X1 port map( A1 => n16672, A2 => n17356, ZN => n16675);
   U19272 : NOR2_X1 port map( A1 => n17014, A2 => n17351, ZN => n16876);
   U19273 : OR2_X1 port map( A1 => n16672, A2 => n4004, ZN => n16674);
   U19274 : XNOR2_X1 port map( A => n18674, B => n17663, ZN => n18501);
   U19275 : XNOR2_X1 port map( A => n17679, B => n18501, ZN => n16698);
   U19276 : NAND2_X1 port map( A1 => n374, A2 => n17368, ZN => n16676);
   U19278 : AND2_X1 port map( A1 => n17573, A2 => n17574, ZN => n16677);
   U19279 : NAND3_X1 port map( A1 => n16682, A2 => n16681, A3 => n16680, ZN => 
                           n16685);
   U19280 : INV_X1 port map( A => n16683, ZN => n16684);
   U19281 : OAI22_X1 port map( A1 => n16685, A2 => n16684, B1 => n17277, B2 => 
                           n17273, ZN => n16690);
   U19282 : NAND4_X1 port map( A1 => n16687, A2 => n17273, A3 => n16686, A4 => 
                           n17276, ZN => n16689);
   U19283 : NAND3_X1 port map( A1 => n17279, A2 => n17254, A3 => n17249, ZN => 
                           n16688);
   U19285 : AND3_X1 port map( A1 => n17145, A2 => n16985, A3 => n17137, ZN => 
                           n16693);
   U19286 : INV_X1 port map( A => n17664, ZN => n18116);
   U19287 : XNOR2_X1 port map( A => n18116, B => n21533, ZN => n16696);
   U19288 : XNOR2_X1 port map( A => n18390, B => n16696, ZN => n16697);
   U19289 : NAND2_X1 port map( A1 => n19290, A2 => n19559, ZN => n16699);
   U19290 : AOI21_X1 port map( B1 => n16699, B2 => n19560, A => n19138, ZN => 
                           n16700);
   U19291 : INV_X1 port map( A => n18678, ZN => n16713);
   U19292 : OAI21_X1 port map( B1 => n17319, B2 => n17320, A => n17321, ZN => 
                           n16712);
   U19293 : XNOR2_X1 port map( A => n16713, B => n18633, ZN => n18303);
   U19294 : INV_X1 port map( A => n18303, ZN => n17912);
   U19295 : XNOR2_X1 port map( A => n17912, B => n18226, ZN => n16738);
   U19296 : XNOR2_X1 port map( A => n18188, B => n2228, ZN => n16736);
   U19297 : NAND3_X1 port map( A1 => n17332, A2 => n17336, A3 => n17335, ZN => 
                           n16729);
   U19298 : NAND2_X1 port map( A1 => n25412, A2 => n17335, ZN => n16725);
   U19299 : XNOR2_X1 port map( A => n17788, B => n16736, ZN => n16737);
   U19301 : XNOR2_X1 port map( A => n18195, B => n1875, ZN => n16745);
   U19302 : NOR2_X1 port map( A1 => n17086, A2 => n17085, ZN => n16741);
   U19303 : NOR2_X1 port map( A1 => n17615, A2 => n17408, ZN => n16744);
   U19304 : XNOR2_X1 port map( A => n18432, B => n18693, ZN => n17785);
   U19305 : XNOR2_X1 port map( A => n17785, B => n16745, ZN => n16761);
   U19308 : INV_X1 port map( A => n17421, ZN => n16752);
   U19309 : NOR2_X1 port map( A1 => n17423, A2 => n17424, ZN => n16749);
   U19310 : OAI21_X1 port map( B1 => n17381, B2 => n17421, A => n16749, ZN => 
                           n16751);
   U19311 : NAND3_X1 port map( A1 => n17425, A2 => n16752, A3 => n17423, ZN => 
                           n16750);
   U19312 : OAI211_X1 port map( C1 => n17379, C2 => n16752, A => n16751, B => 
                           n16750, ZN => n18476);
   U19314 : NAND2_X1 port map( A1 => n17289, A2 => n17284, ZN => n17538);
   U19315 : NAND2_X1 port map( A1 => n17541, A2 => n17538, ZN => n16754);
   U19317 : OAI21_X1 port map( B1 => n16755, B2 => n16754, A => n17544, ZN => 
                           n16759);
   U19318 : NAND2_X1 port map( A1 => n17419, A2 => n25433, ZN => n16756);
   U19319 : NAND2_X1 port map( A1 => n17227, A2 => n25246, ZN => n16757);
   U19320 : XNOR2_X1 port map( A => n16759, B => n17931, ZN => n18218);
   U19321 : XNOR2_X1 port map( A => n16761, B => n16760, ZN => n19261);
   U19322 : NAND2_X1 port map( A1 => n24386, A2 => n19261, ZN => n19146);
   U19323 : INV_X1 port map( A => n17368, ZN => n17571);
   U19324 : INV_X1 port map( A => n18233, ZN => n16768);
   U19325 : XNOR2_X1 port map( A => n16768, B => n17681, ZN => n18142);
   U19326 : INV_X1 port map( A => n16770, ZN => n17040);
   U19328 : AOI22_X1 port map( A1 => n17364, A2 => n25058, B1 => n16989, B2 => 
                           n16770, ZN => n16771);
   U19331 : NAND3_X1 port map( A1 => n16775, A2 => n17049, A3 => n17050, ZN => 
                           n16776);
   U19332 : XNOR2_X1 port map( A => n18660, B => n18611, ZN => n18333);
   U19333 : XNOR2_X1 port map( A => n18142, B => n18333, ZN => n16786);
   U19334 : INV_X1 port map( A => n16778, ZN => n16779);
   U19335 : INV_X1 port map( A => n17581, ZN => n16783);
   U19336 : XNOR2_X1 port map( A => n18103, B => n16783, ZN => n18178);
   U19337 : XNOR2_X1 port map( A => n16784, B => n18178, ZN => n16785);
   U19339 : NAND2_X1 port map( A1 => n17134, A2 => n17132, ZN => n16787);
   U19340 : OAI21_X1 port map( B1 => n17134, B2 => n4684, A => n16787, ZN => 
                           n16790);
   U19343 : INV_X1 port map( A => n18208, ZN => n16800);
   U19345 : XNOR2_X1 port map( A => n18602, B => n16799, ZN => n18324);
   U19346 : INV_X1 port map( A => n18324, ZN => n17898);
   U19347 : XNOR2_X1 port map( A => n17898, B => n16800, ZN => n16821);
   U19348 : MUX2_X1 port map( A => n17100, B => n25357, S => n17114, Z => 
                           n16804);
   U19349 : NOR2_X1 port map( A1 => n16802, A2 => n16801, ZN => n16803);
   U19350 : MUX2_X2 port map( A => n16804, B => n16803, S => n2581, Z => n18446
                           );
   U19351 : XNOR2_X1 port map( A => n18446, B => n20995, ZN => n16819);
   U19352 : NAND2_X1 port map( A1 => n17081, A2 => n16809, ZN => n16896);
   U19353 : AOI21_X1 port map( B1 => n17481, B2 => n17077, A => n17078, ZN => 
                           n16807);
   U19354 : NAND2_X1 port map( A1 => n24660, A2 => n17478, ZN => n16806);
   U19356 : NAND3_X1 port map( A1 => n16810, A2 => n16809, A3 => n16808, ZN => 
                           n17477);
   U19357 : NOR2_X1 port map( A1 => n25429, A2 => n17477, ZN => n16811);
   U19359 : NAND2_X1 port map( A1 => n17729, A2 => n25472, ZN => n16817);
   U19360 : NAND2_X1 port map( A1 => n25472, A2 => n17734, ZN => n16814);
   U19361 : NOR2_X1 port map( A1 => n17728, A2 => n17485, ZN => n17094);
   U19362 : INV_X1 port map( A => n17094, ZN => n16813);
   U19364 : XNOR2_X1 port map( A => n18418, B => n18149, ZN => n18607);
   U19365 : INV_X1 port map( A => n18607, ZN => n16818);
   U19366 : XNOR2_X1 port map( A => n16819, B => n16818, ZN => n16820);
   U19367 : XNOR2_X1 port map( A => n16821, B => n16820, ZN => n17556);
   U19368 : NAND3_X1 port map( A1 => n19146, A2 => n16822, A3 => n18919, ZN => 
                           n16887);
   U19369 : INV_X1 port map( A => n17171, ZN => n17523);
   U19370 : MUX2_X1 port map( A => n16862, B => n16823, S => n17174, Z => 
                           n16825);
   U19371 : OAI21_X1 port map( B1 => n17170, B2 => n17173, A => n17523, ZN => 
                           n16824);
   U19372 : INV_X1 port map( A => n17445, ZN => n17125);
   U19374 : INV_X1 port map( A => n16826, ZN => n16827);
   U19375 : AOI22_X1 port map( A1 => n17125, A2 => n2549, B1 => n16827, B2 => 
                           n16964, ZN => n16831);
   U19376 : OAI22_X1 port map( A1 => n16831, A2 => n16830, B1 => n1612, B2 => 
                           n16829, ZN => n17905);
   U19377 : XNOR2_X1 port map( A => n17839, B => n17905, ZN => n18237);
   U19378 : INV_X1 port map( A => n16979, ZN => n17457);
   U19379 : AOI21_X1 port map( B1 => n17455, B2 => n523, A => n17457, ZN => 
                           n16833);
   U19380 : OAI21_X1 port map( B1 => n17163, B2 => n17165, A => n16836, ZN => 
                           n16837);
   U19381 : INV_X1 port map( A => n16837, ZN => n16842);
   U19382 : NAND2_X1 port map( A1 => n17164, A2 => n17166, ZN => n16840);
   U19384 : MUX2_X1 port map( A => n16840, B => n16839, S => n17163, Z => 
                           n16841);
   U19385 : XNOR2_X1 port map( A => n18124, B => n18121, ZN => n16843);
   U19386 : XNOR2_X1 port map( A => n18237, B => n16843, ZN => n16858);
   U19387 : INV_X1 port map( A => n16847, ZN => n16854);
   U19388 : AND2_X1 port map( A1 => n17144, A2 => n16985, ZN => n16850);
   U19389 : NAND3_X1 port map( A1 => n17138, A2 => n16851, A3 => n17139, ZN => 
                           n16852);
   U19391 : XNOR2_X1 port map( A => n18435, B => n18669, ZN => n16856);
   U19392 : XNOR2_X1 port map( A => n18382, B => n2208, ZN => n16855);
   U19393 : XNOR2_X1 port map( A => n16855, B => n16856, ZN => n16857);
   U19394 : XNOR2_X1 port map( A => n16858, B => n16857, ZN => n19266);
   U19395 : NAND2_X1 port map( A1 => n19263, A2 => n19266, ZN => n16886);
   U19396 : INV_X1 port map( A => n17241, ZN => n17240);
   U19397 : XNOR2_X1 port map( A => n18308, B => n3152, ZN => n16868);
   U19398 : NOR3_X1 port map( A1 => n17524, A2 => n17170, A3 => n17175, ZN => 
                           n16861);
   U19399 : NOR2_X1 port map( A1 => n16862, A2 => n16861, ZN => n17525);
   U19400 : NOR2_X1 port map( A1 => n17524, A2 => n17171, ZN => n17177);
   U19401 : NOR2_X1 port map( A1 => n16863, A2 => n16112, ZN => n16864);
   U19402 : OAI21_X1 port map( B1 => n17177, B2 => n16864, A => n17522, ZN => 
                           n16865);
   U19403 : NAND2_X1 port map( A1 => n17525, A2 => n16865, ZN => n16866);
   U19404 : XNOR2_X1 port map( A => n16867, B => n16868, ZN => n16884);
   U19405 : NOR2_X1 port map( A1 => n25003, A2 => n17192, ZN => n16870);
   U19407 : OAI22_X1 port map( A1 => n16873, A2 => n17389, B1 => n16872, B2 => 
                           n17387, ZN => n16874);
   U19408 : NAND3_X1 port map( A1 => n367, A2 => n4004, A3 => n25491, ZN => 
                           n16877);
   U19409 : NAND2_X1 port map( A1 => n16878, A2 => n24391, ZN => n16882);
   U19410 : INV_X1 port map( A => n17216, ZN => n17021);
   U19411 : NAND2_X1 port map( A1 => n17021, A2 => n17015, ZN => n16881);
   U19412 : NAND3_X1 port map( A1 => n17216, A2 => n17016, A3 => n17208, ZN => 
                           n16879);
   U19413 : XNOR2_X1 port map( A => n18129, B => n25194, ZN => n18629);
   U19414 : XNOR2_X1 port map( A => n18248, B => n18629, ZN => n16883);
   U19415 : XNOR2_X1 port map( A => n16883, B => n16884, ZN => n18914);
   U19416 : NAND3_X2 port map( A1 => n16887, A2 => n16886, A3 => n16885, ZN => 
                           n20669);
   U19419 : MUX2_X1 port map( A => n17485, B => n17728, S => n17734, Z => 
                           n16889);
   U19420 : NOR2_X1 port map( A1 => n17486, A2 => n24410, ZN => n17737);
   U19421 : MUX2_X1 port map( A => n16889, B => n17737, S => n17729, Z => 
                           n16891);
   U19422 : NOR3_X1 port map( A1 => n17728, A2 => n17730, A3 => n17731, ZN => 
                           n16890);
   U19423 : NOR2_X1 port map( A1 => n16891, A2 => n16890, ZN => n18122);
   U19424 : XNOR2_X1 port map( A => n18122, B => n18239, ZN => n16906);
   U19425 : NOR2_X1 port map( A1 => n17077, A2 => n17078, ZN => n16894);
   U19426 : NOR2_X1 port map( A1 => n16896, A2 => n17076, ZN => n16899);
   U19427 : NAND2_X1 port map( A1 => n1033, A2 => n17629, ZN => n16905);
   U19428 : OAI211_X1 port map( C1 => n17472, C2 => n16905, A => n16904, B => 
                           n16903, ZN => n18038);
   U19429 : XNOR2_X1 port map( A => n18038, B => n17595, ZN => n18667);
   U19430 : XNOR2_X1 port map( A => n16906, B => n18667, ZN => n16914);
   U19431 : MUX2_X1 port map( A => n17114, B => n17118, S => n17119, Z => 
                           n16907);
   U19432 : NAND2_X1 port map( A1 => n16907, A2 => n2580, ZN => n16909);
   U19433 : NOR2_X1 port map( A1 => n17120, A2 => n17119, ZN => n16908);
   U19434 : XNOR2_X1 port map( A => n18582, B => n836, ZN => n16912);
   U19435 : XNOR2_X1 port map( A => n17907, B => n18539, ZN => n16911);
   U19436 : XNOR2_X1 port map( A => n16912, B => n16911, ZN => n16913);
   U19437 : XNOR2_X1 port map( A => n16913, B => n16914, ZN => n19309);
   U19438 : INV_X1 port map( A => n16974, ZN => n16918);
   U19439 : OAI21_X1 port map( B1 => n17336, B2 => n16973, A => n16971, ZN => 
                           n16916);
   U19441 : INV_X1 port map( A => n16920, ZN => n16922);
   U19442 : NAND2_X1 port map( A1 => n17304, A2 => n24543, ZN => n17314);
   U19443 : XNOR2_X1 port map( A => n17720, B => n17582, ZN => n18657);
   U19444 : INV_X1 port map( A => n18657, ZN => n18176);
   U19446 : OAI21_X1 port map( B1 => n17326, B2 => n17319, A => n4426, ZN => 
                           n16925);
   U19447 : AOI22_X2 port map( A1 => n16926, A2 => n16927, B1 => n16925, B2 => 
                           n15673, ZN => n18658);
   U19448 : XNOR2_X1 port map( A => n18658, B => n18532, ZN => n18267);
   U19449 : INV_X1 port map( A => n18267, ZN => n16928);
   U19450 : XNOR2_X1 port map( A => n16928, B => n18176, ZN => n16939);
   U19451 : OAI22_X1 port map( A1 => n16932, A2 => n25031, B1 => n24585, B2 => 
                           n17059, ZN => n16930);
   U19452 : NAND2_X1 port map( A1 => n16930, A2 => n16929, ZN => n16934);
   U19453 : INV_X1 port map( A => n17059, ZN => n16931);
   U19454 : NAND2_X1 port map( A1 => n16932, A2 => n16931, ZN => n16933);
   U19455 : XNOR2_X1 port map( A => n18067, B => n923, ZN => n16936);
   U19456 : XOR2_X1 port map( A => n16937, B => n16936, Z => n16938);
   U19457 : MUX2_X1 port map( A => n4487, B => n17407, S => n16940, Z => n16943
                           );
   U19458 : NOR3_X1 port map( A1 => n17410, A2 => n17615, A3 => n17255, ZN => 
                           n17611);
   U19460 : XNOR2_X1 port map( A => n16946, B => n18677, ZN => n16949);
   U19461 : XNOR2_X1 port map( A => n18227, B => n16947, ZN => n16948);
   U19462 : XNOR2_X1 port map( A => n16949, B => n16948, ZN => n16960);
   U19463 : NAND2_X1 port map( A1 => n16952, A2 => n17230, ZN => n16953);
   U19464 : INV_X1 port map( A => n17791, ZN => n16959);
   U19465 : NOR2_X1 port map( A1 => n17227, A2 => n25433, ZN => n17416);
   U19466 : NAND3_X1 port map( A1 => n16957, A2 => n16956, A3 => n1230, ZN => 
                           n16958);
   U19467 : XNOR2_X1 port map( A => n16959, B => n18675, ZN => n18189);
   U19468 : INV_X1 port map( A => n18189, ZN => n18089);
   U19469 : BUF_X2 port map( A => n17562, Z => n18923);
   U19470 : NAND2_X1 port map( A1 => n16964, A2 => n16962, ZN => n16968);
   U19471 : INV_X1 port map( A => n17662, ZN => n16967);
   U19472 : NAND2_X1 port map( A1 => n16963, A2 => n24444, ZN => n17446);
   U19473 : INV_X1 port map( A => n17446, ZN => n17127);
   U19474 : NOR2_X1 port map( A1 => n17439, A2 => n16964, ZN => n16965);
   U19475 : INV_X1 port map( A => n17661, ZN => n16966);
   U19476 : OAI21_X1 port map( B1 => n16967, B2 => n16966, A => n23347, ZN => 
                           n16970);
   U19477 : NOR2_X1 port map( A1 => n16974, A2 => n17335, ZN => n16972);
   U19478 : NOR2_X1 port map( A1 => n16972, A2 => n16971, ZN => n16978);
   U19479 : NOR2_X1 port map( A1 => n16973, A2 => n376, ZN => n16975);
   U19480 : OAI21_X1 port map( B1 => n16976, B2 => n16975, A => n16974, ZN => 
                           n16977);
   U19481 : NOR2_X1 port map( A1 => n16979, A2 => n16980, ZN => n16983);
   U19482 : OAI21_X1 port map( B1 => n24942, B2 => n17453, A => n5072, ZN => 
                           n16982);
   U19483 : NAND3_X1 port map( A1 => n24942, A2 => n523, A3 => n17451, ZN => 
                           n16981);
   U19484 : XNOR2_X1 port map( A => n18562, B => n18172, ZN => n18687);
   U19485 : MUX2_X1 port map( A => n17141, B => n17137, S => n17139, Z => 
                           n16987);
   U19486 : OAI21_X1 port map( B1 => n16984, B2 => n17144, A => n17138, ZN => 
                           n16986);
   U19487 : INV_X1 port map( A => n19313, ZN => n19317);
   U19488 : NAND2_X1 port map( A1 => n19317, A2 => n5371, ZN => n17010);
   U19489 : NOR2_X1 port map( A1 => n25214, A2 => n16989, ZN => n16990);
   U19490 : NAND3_X1 port map( A1 => n16991, A2 => n288, A3 => n287, ZN => 
                           n16992);
   U19493 : XNOR2_X1 port map( A => n24536, B => n18220, ZN => n16996);
   U19494 : XNOR2_X1 port map( A => n18692, B => n16996, ZN => n17008);
   U19495 : NAND2_X1 port map( A1 => n17572, A2 => n16998, ZN => n16999);
   U19496 : NAND3_X1 port map( A1 => n17049, A2 => n17053, A3 => n17050, ZN => 
                           n17001);
   U19497 : XNOR2_X1 port map( A => n18200, B => n18695, ZN => n17006);
   U19498 : XNOR2_X1 port map( A => n18006, B => n2033, ZN => n17005);
   U19499 : XNOR2_X1 port map( A => n17006, B => n17005, ZN => n17007);
   U19500 : INV_X1 port map( A => n19312, ZN => n17009);
   U19501 : MUX2_X1 port map( A => n17011, B => n17010, S => n17009, Z => 
                           n17036);
   U19502 : MUX2_X1 port map( A => n17015, B => n17212, S => n25200, Z => 
                           n17022);
   U19503 : NAND2_X1 port map( A1 => n17016, A2 => n25201, ZN => n17018);
   U19504 : OAI22_X1 port map( A1 => n17018, A2 => n5512, B1 => n17216, B2 => 
                           n17017, ZN => n17019);
   U19505 : INV_X1 port map( A => n17019, ZN => n17020);
   U19506 : OAI21_X1 port map( B1 => n17186, B2 => n3602, A => n17185, ZN => 
                           n17024);
   U19507 : XNOR2_X1 port map( A => n18325, B => n18096, ZN => n18704);
   U19508 : OAI211_X1 port map( C1 => n17400, C2 => n25003, A => n17398, B => 
                           n17198, ZN => n17029);
   U19509 : INV_X1 port map( A => n17399, ZN => n17193);
   U19510 : XNOR2_X1 port map( A => n18451, B => n4189, ZN => n17033);
   U19511 : NAND2_X1 port map( A1 => n19311, A2 => n19310, ZN => n18925);
   U19512 : NOR2_X1 port map( A1 => n24567, A2 => n20336, ZN => n20672);
   U19513 : NAND2_X1 port map( A1 => n17364, A2 => n17362, ZN => n17037);
   U19514 : XNOR2_X1 port map( A => n18023, B => n17041, ZN => n18349);
   U19515 : AOI21_X1 port map( B1 => n17370, B2 => n17044, A => n17572, ZN => 
                           n17046);
   U19516 : NOR3_X1 port map( A1 => n5522, A2 => n17574, A3 => n3371, ZN => 
                           n17045);
   U19517 : OR3_X2 port map( A1 => n17576, A2 => n17046, A3 => n17045, ZN => 
                           n17748);
   U19518 : INV_X1 port map( A => n17748, ZN => n18252);
   U19519 : XNOR2_X1 port map( A => n18252, B => n18451, ZN => n17047);
   U19520 : XNOR2_X1 port map( A => n18349, B => n17047, ZN => n17074);
   U19521 : NAND2_X1 port map( A1 => n17054, A2 => n17059, ZN => n17055);
   U19522 : NAND2_X1 port map( A1 => n17056, A2 => n17055, ZN => n17058);
   U19523 : NOR2_X1 port map( A1 => n17060, A2 => n17059, ZN => n17064);
   U19524 : NOR2_X1 port map( A1 => n24585, A2 => n24398, ZN => n17063);
   U19525 : XNOR2_X1 port map( A => n17819, B => n18350, ZN => n17072);
   U19526 : NAND2_X1 port map( A1 => n17068, A2 => n369, ZN => n17066);
   U19527 : XNOR2_X1 port map( A => n18599, B => n92, ZN => n17071);
   U19528 : XNOR2_X1 port map( A => n17071, B => n17072, ZN => n17073);
   U19529 : AOI21_X1 port map( B1 => n17480, B2 => n17482, A => n17076, ZN => 
                           n17083);
   U19530 : AOI21_X1 port map( B1 => n17079, B2 => n17078, A => n17077, ZN => 
                           n17080);
   U19531 : NOR2_X1 port map( A1 => n25429, A2 => n17080, ZN => n17082);
   U19533 : XNOR2_X1 port map( A => n17680, B => n18483, ZN => n17953);
   U19534 : INV_X1 port map( A => n17084, ZN => n17091);
   U19535 : XNOR2_X1 port map( A => n17953, B => n17092, ZN => n17113);
   U19536 : AOI22_X1 port map( A1 => n17093, A2 => n17484, B1 => n17735, B2 => 
                           n17731, ZN => n17097);
   U19537 : NAND2_X1 port map( A1 => n17735, A2 => n17094, ZN => n17096);
   U19538 : OR2_X1 port map( A1 => n17690, A2 => n17486, ZN => n17095);
   U19539 : NAND2_X1 port map( A1 => n17120, A2 => n17118, ZN => n17098);
   U19540 : AND3_X1 port map( A1 => n17099, A2 => n17116, A3 => n17098, ZN => 
                           n17106);
   U19543 : NAND3_X1 port map( A1 => n17114, A2 => n16572, A3 => n25357, ZN => 
                           n17104);
   U19544 : OAI211_X2 port map( C1 => n17106, C2 => n2580, A => n17105, B => 
                           n17104, ZN => n18032);
   U19545 : XNOR2_X1 port map( A => n18356, B => n18032, ZN => n18268);
   U19547 : NAND2_X1 port map( A1 => n17132, A2 => n17131, ZN => n17109);
   U19548 : XNOR2_X1 port map( A => n17832, B => n1935, ZN => n17110);
   U19550 : NOR2_X1 port map( A1 => n18934, A2 => n17496, ZN => n17495);
   U19551 : OAI211_X1 port map( C1 => n17116, C2 => n17115, A => n17114, B => 
                           n17118, ZN => n17117);
   U19552 : INV_X1 port map( A => n17117, ZN => n17124);
   U19553 : NOR2_X1 port map( A1 => n17119, A2 => n17118, ZN => n17121);
   U19555 : OAI211_X1 port map( C1 => n17125, C2 => n24444, A => n17439, B => 
                           n17442, ZN => n17126);
   U19556 : OAI21_X1 port map( B1 => n17128, B2 => n17127, A => n17126, ZN => 
                           n18276);
   U19557 : XNOR2_X1 port map( A => n18276, B => n17958, ZN => n17136);
   U19558 : OAI211_X1 port map( C1 => n17132, C2 => n17131, A => n4684, B => 
                           n17130, ZN => n17133);
   U19559 : XNOR2_X1 port map( A => n18341, B => n1826, ZN => n17135);
   U19560 : XNOR2_X1 port map( A => n17136, B => n17135, ZN => n17154);
   U19561 : NOR2_X1 port map( A1 => n17138, A2 => n17137, ZN => n17143);
   U19562 : AOI21_X1 port map( B1 => n17145, B2 => n17140, A => n17139, ZN => 
                           n17142);
   U19563 : NOR2_X1 port map( A1 => n17145, A2 => n17144, ZN => n17146);
   U19565 : NAND2_X1 port map( A1 => n17460, A2 => n17451, ZN => n17151);
   U19566 : NAND2_X1 port map( A1 => n523, A2 => n17450, ZN => n17148);
   U19569 : XNOR2_X1 port map( A => n18694, B => n18060, ZN => n18367);
   U19570 : INV_X1 port map( A => n18367, ZN => n17693);
   U19571 : XNOR2_X1 port map( A => n17693, B => n18475, ZN => n17153);
   U19572 : XNOR2_X2 port map( A => n17153, B => n17154, ZN => n19326);
   U19573 : NAND3_X1 port map( A1 => n17158, A2 => n17157, A3 => n17156, ZN => 
                           n17162);
   U19574 : INV_X1 port map( A => n17159, ZN => n17161);
   U19576 : NAND3_X1 port map( A1 => n17165, A2 => n17164, A3 => n17163, ZN => 
                           n17168);
   U19577 : XNOR2_X1 port map( A => n25380, B => n3093, ZN => n17178);
   U19579 : XNOR2_X1 port map( A => n17178, B => n17806, ZN => n17191);
   U19580 : AND2_X1 port map( A1 => n3602, A2 => n17184, ZN => n17188);
   U19581 : NOR2_X1 port map( A1 => n17185, A2 => n17391, ZN => n17187);
   U19582 : AOI22_X1 port map( A1 => n17188, A2 => n17389, B1 => n17187, B2 => 
                           n3604, ZN => n17189);
   U19583 : OAI21_X2 port map( B1 => n17190, B2 => n16203, A => n17189, ZN => 
                           n18295);
   U19584 : XNOR2_X1 port map( A => n17191, B => n18387, ZN => n17222);
   U19585 : MUX2_X1 port map( A => n17198, B => n17195, S => n17192, Z => 
                           n17194);
   U19586 : AND2_X1 port map( A1 => n17194, A2 => n17193, ZN => n17201);
   U19587 : NAND2_X1 port map( A1 => n4039, A2 => n17400, ZN => n17199);
   U19588 : OAI22_X1 port map( A1 => n17199, A2 => n17198, B1 => n17197, B2 => 
                           n17196, ZN => n17200);
   U19589 : INV_X1 port map( A => n17202, ZN => n17204);
   U19590 : NAND2_X1 port map( A1 => n17342, A2 => n17346, ZN => n17203);
   U19591 : AOI21_X1 port map( B1 => n17204, B2 => n17203, A => n17347, ZN => 
                           n17205);
   U19592 : NOR2_X1 port map( A1 => n17206, A2 => n17205, ZN => n17220);
   U19594 : NAND2_X1 port map( A1 => n25201, A2 => n17208, ZN => n17209);
   U19595 : NAND3_X1 port map( A1 => n17210, A2 => n5512, A3 => n17209, ZN => 
                           n17219);
   U19596 : NAND3_X1 port map( A1 => n24391, A2 => n17212, A3 => n17211, ZN => 
                           n17218);
   U19597 : NAND3_X1 port map( A1 => n17216, A2 => n25201, A3 => n17214, ZN => 
                           n17217);
   U19598 : XNOR2_X1 port map( A => n17220, B => n18187, ZN => n18459);
   U19599 : XNOR2_X1 port map( A => n18290, B => n18459, ZN => n17221);
   U19600 : XNOR2_X1 port map( A => n17222, B => n17221, ZN => n17497);
   U19602 : NOR2_X1 port map( A1 => n24583, A2 => n19326, ZN => n17223);
   U19603 : NOR2_X1 port map( A1 => n17495, A2 => n17223, ZN => n17310);
   U19604 : XNOR2_X1 port map( A => n18261, B => n18666, ZN => n18380);
   U19605 : MUX2_X1 port map( A => n17288, B => n17283, S => n17229, Z => 
                           n17233);
   U19606 : NAND2_X1 port map( A1 => n17283, A2 => n17229, ZN => n17286);
   U19607 : MUX2_X1 port map( A => n17286, B => n17231, S => n17230, Z => 
                           n17232);
   U19608 : XNOR2_X1 port map( A => n18239, B => n18665, ZN => n17234);
   U19609 : XNOR2_X1 port map( A => n18380, B => n17234, ZN => n17263);
   U19610 : INV_X1 port map( A => n17235, ZN => n17239);
   U19611 : NAND2_X1 port map( A1 => n17239, A2 => n17238, ZN => n17246);
   U19612 : AND2_X1 port map( A1 => n17346, A2 => n17344, ZN => n17245);
   U19613 : MUX2_X1 port map( A => n17242, B => n17241, S => n15314, Z => 
                           n17243);
   U19614 : NAND2_X1 port map( A1 => n17347, A2 => n17243, ZN => n17244);
   U19616 : NAND3_X1 port map( A1 => n17275, A2 => n17277, A3 => n17249, ZN => 
                           n17250);
   U19617 : NAND3_X1 port map( A1 => n17407, A2 => n17607, A3 => n17408, ZN => 
                           n17256);
   U19618 : NOR2_X1 port map( A1 => n4487, A2 => n17257, ZN => n17258);
   U19619 : NOR2_X2 port map( A1 => n17259, A2 => n17258, ZN => n18489);
   U19620 : XNOR2_X1 port map( A => n18489, B => n1726, ZN => n17260);
   U19621 : XNOR2_X1 port map( A => n17261, B => n17260, ZN => n17262);
   U19622 : XNOR2_X1 port map( A => n17263, B => n17262, ZN => n17264);
   U19623 : INV_X1 port map( A => n17264, ZN => n18933);
   U19624 : NOR2_X1 port map( A1 => n17264, A2 => n17496, ZN => n19331);
   U19625 : INV_X1 port map( A => n17319, ZN => n17265);
   U19626 : NOR2_X1 port map( A1 => n17267, A2 => n17266, ZN => n17270);
   U19627 : INV_X1 port map( A => n17326, ZN => n17323);
   U19628 : NOR2_X1 port map( A1 => n17322, A2 => n17323, ZN => n17268);
   U19630 : AND2_X1 port map( A1 => n17273, A2 => n17276, ZN => n17271);
   U19631 : NAND2_X1 port map( A1 => n17272, A2 => n17271, ZN => n17281);
   U19632 : NOR2_X1 port map( A1 => n17277, A2 => n17276, ZN => n17278);
   U19633 : NAND2_X1 port map( A1 => n3855, A2 => n17278, ZN => n17280);
   U19634 : AND2_X1 port map( A1 => n17285, A2 => n17286, ZN => n17291);
   U19636 : XNOR2_X1 port map( A => n18512, B => n2058, ZN => n17294);
   U19637 : XNOR2_X1 port map( A => n17294, B => n17520, ZN => n17295);
   U19638 : XNOR2_X1 port map( A => n17295, B => n18372, ZN => n17308);
   U19639 : INV_X1 port map( A => n17296, ZN => n17298);
   U19640 : NAND2_X1 port map( A1 => n17298, A2 => n17297, ZN => n17301);
   U19642 : XNOR2_X1 port map( A => n18465, B => n25411, ZN => n17306);
   U19643 : XNOR2_X1 port map( A => n17306, B => n5300, ZN => n17307);
   U19644 : OAI21_X1 port map( B1 => n19331, B2 => n3034, A => n24583, ZN => 
                           n17309);
   U19645 : INV_X1 port map( A => n20668, ZN => n20671);
   U19646 : MUX2_X1 port map( A => n17311, B => n20672, S => n20671, Z => 
                           n17494);
   U19647 : NOR2_X1 port map( A1 => n20670, A2 => n20335, ZN => n19709);
   U19648 : NAND2_X1 port map( A1 => n17315, A2 => n17314, ZN => n17317);
   U19649 : XNOR2_X1 port map( A => n18448, B => n17819, ZN => n18422);
   U19650 : INV_X1 port map( A => n18447, ZN => n17327);
   U19651 : XNOR2_X1 port map( A => n17328, B => n17327, ZN => n17329);
   U19652 : XNOR2_X1 port map( A => n17329, B => n18422, ZN => n17340);
   U19653 : NAND2_X1 port map( A1 => n3817, A2 => n17335, ZN => n17338);
   U19654 : XNOR2_X1 port map( A => n18423, B => n18599, ZN => n17506);
   U19655 : XNOR2_X1 port map( A => n17506, B => n18214, ZN => n17657);
   U19656 : XNOR2_X1 port map( A => n17340, B => n17657, ZN => n18761);
   U19657 : AOI21_X1 port map( B1 => n17343, B2 => n17342, A => n17341, ZN => 
                           n17345);
   U19658 : NOR3_X1 port map( A1 => n17348, A2 => n17347, A3 => n17346, ZN => 
                           n17349);
   U19659 : NOR2_X1 port map( A1 => n17350, A2 => n17349, ZN => n17359);
   U19660 : NAND2_X1 port map( A1 => n17357, A2 => n17351, ZN => n17355);
   U19661 : NAND2_X1 port map( A1 => n17353, A2 => n25491, ZN => n17354);
   U19662 : OAI211_X1 port map( C1 => n17357, C2 => n17356, A => n17355, B => 
                           n17354, ZN => n17358);
   U19663 : XNOR2_X1 port map( A => n17359, B => n18123, ZN => n17642);
   U19664 : XNOR2_X1 port map( A => n17642, B => n17360, ZN => n17377);
   U19665 : NOR2_X1 port map( A1 => n17362, A2 => n25215, ZN => n17365);
   U19666 : NOR2_X1 port map( A1 => n17366, A2 => n370, ZN => n17367);
   U19667 : XNOR2_X1 port map( A => n18491, B => n18669, ZN => n17375);
   U19668 : NAND2_X1 port map( A1 => n24471, A2 => n17368, ZN => n17369);
   U19669 : NOR2_X1 port map( A1 => n24471, A2 => n17574, ZN => n17372);
   U19670 : NAND2_X1 port map( A1 => n17378, A2 => n17425, ZN => n17380);
   U19671 : MUX2_X1 port map( A => n17426, B => n17380, S => n17379, Z => 
                           n17385);
   U19672 : NAND2_X1 port map( A1 => n17423, A2 => n17381, ZN => n17383);
   U19673 : NOR2_X1 port map( A1 => n17383, A2 => n17382, ZN => n17384);
   U19674 : NOR2_X2 port map( A1 => n17385, A2 => n17384, ZN => n18407);
   U19675 : INV_X1 port map( A => n17389, ZN => n17388);
   U19676 : MUX2_X1 port map( A => n17391, B => n17390, S => n17389, Z => 
                           n17392);
   U19678 : XNOR2_X1 port map( A => n18531, B => n18102, ZN => n18232);
   U19679 : INV_X1 port map( A => n18232, ZN => n17394);
   U19680 : XNOR2_X1 port map( A => n17394, B => n17648, ZN => n17405);
   U19681 : OAI21_X1 port map( B1 => n17397, B2 => n17396, A => n17395, ZN => 
                           n17402);
   U19683 : XNOR2_X1 port map( A => n17832, B => n18484, ZN => n18404);
   U19684 : XNOR2_X1 port map( A => n18660, B => n688, ZN => n17403);
   U19685 : XNOR2_X1 port map( A => n18404, B => n17403, ZN => n17404);
   U19686 : XNOR2_X2 port map( A => n17405, B => n17404, ZN => n19531);
   U19687 : INV_X1 port map( A => n17881, ZN => n17406);
   U19688 : XNOR2_X1 port map( A => n18311, B => n17406, ZN => n17660);
   U19689 : OAI22_X1 port map( A1 => n17410, A2 => n17608, B1 => n17407, B2 => 
                           n17607, ZN => n17411);
   U19690 : INV_X1 port map( A => n17408, ZN => n17612);
   U19691 : XNOR2_X1 port map( A => n18128, B => n18308, ZN => n17412);
   U19692 : XNOR2_X1 port map( A => n17660, B => n17412, ZN => n17432);
   U19693 : NOR2_X1 port map( A1 => n17414, A2 => n17413, ZN => n17415);
   U19694 : INV_X1 port map( A => n18512, ZN => n17420);
   U19695 : XNOR2_X1 port map( A => n18466, B => n17420, ZN => n17967);
   U19697 : NAND3_X1 port map( A1 => n17423, A2 => n17422, A3 => n5409, ZN => 
                           n17428);
   U19698 : OAI21_X1 port map( B1 => n17426, B2 => n17425, A => n17424, ZN => 
                           n17427);
   U19700 : INV_X1 port map( A => n18515, ZN => n18467);
   U19701 : XNOR2_X1 port map( A => n17967, B => n17430, ZN => n17431);
   U19702 : XNOR2_X1 port map( A => n17432, B => n17431, ZN => n19145);
   U19703 : INV_X1 port map( A => n19145, ZN => n19269);
   U19704 : NOR2_X1 port map( A1 => n17439, A2 => n24444, ZN => n17443);
   U19705 : NOR2_X1 port map( A1 => n17446, A2 => n17445, ZN => n17447);
   U19706 : XNOR2_X1 port map( A => n18456, B => n17806, ZN => n18415);
   U19708 : XNOR2_X1 port map( A => n18225, B => n18415, ZN => n17471);
   U19709 : XNOR2_X1 port map( A => n24488, B => n18388, ZN => n17469);
   U19710 : XNOR2_X1 port map( A => n25379, B => n2036, ZN => n17468);
   U19711 : XNOR2_X1 port map( A => n17469, B => n17468, ZN => n17470);
   U19712 : XNOR2_X1 port map( A => n17471, B => n17470, ZN => n18762);
   U19713 : AND2_X1 port map( A1 => n19269, A2 => n19534, ZN => n19533);
   U19715 : XNOR2_X1 port map( A => n18473, B => n17476, ZN => n18219);
   U19716 : INV_X1 port map( A => n18219, ZN => n17489);
   U19717 : INV_X1 port map( A => n17477, ZN => n17483);
   U19718 : AND2_X1 port map( A1 => n25472, A2 => n17485, ZN => n17688);
   U19719 : NAND2_X1 port map( A1 => n17688, A2 => n17687, ZN => n17487);
   U19720 : NAND3_X1 port map( A1 => n17690, A2 => n17686, A3 => n17487, ZN => 
                           n17488);
   U19721 : XNOR2_X1 port map( A => n18365, B => n17488, ZN => n18478);
   U19722 : XNOR2_X1 port map( A => n17489, B => n18478, ZN => n17493);
   U19723 : XNOR2_X1 port map( A => n17958, B => n18693, ZN => n17491);
   U19724 : XNOR2_X1 port map( A => n18341, B => n21204, ZN => n17490);
   U19725 : XNOR2_X1 port map( A => n17491, B => n17490, ZN => n17492);
   U19727 : INV_X1 port map( A => n20338, ZN => n20341);
   U19731 : NAND2_X1 port map( A1 => n25566, A2 => n19329, ZN => n17944);
   U19732 : AOI21_X1 port map( B1 => n19327, B2 => n17944, A => n17495, ZN => 
                           n17500);
   U19733 : INV_X1 port map( A => n17496, ZN => n19328);
   U19734 : INV_X1 port map( A => n17498, ZN => n17499);
   U19735 : AOI21_X1 port map( B1 => n19132, B2 => n18767, A => n18766, ZN => 
                           n17503);
   U19736 : INV_X1 port map( A => n19132, ZN => n19303);
   U19737 : AND2_X1 port map( A1 => n19303, A2 => n19133, ZN => n18768);
   U19738 : INV_X1 port map( A => n18768, ZN => n17502);
   U19739 : NAND2_X1 port map( A1 => n19307, A2 => n24324, ZN => n17501);
   U19740 : XNOR2_X1 port map( A => n17504, B => n18446, ZN => n17505);
   U19741 : INV_X1 port map( A => n18420, ZN => n18022);
   U19742 : XNOR2_X1 port map( A => n18022, B => n17816, ZN => n18521);
   U19743 : XNOR2_X1 port map( A => n18521, B => n17505, ZN => n17508);
   U19744 : XNOR2_X1 port map( A => n18098, B => n17506, ZN => n17507);
   U19745 : XNOR2_X1 port map( A => n17681, B => n17993, ZN => n17833);
   U19746 : INV_X1 port map( A => n17833, ZN => n17509);
   U19747 : XNOR2_X1 port map( A => n17509, B => n17648, ZN => n17512);
   U19748 : XNOR2_X1 port map( A => n18103, B => n2241, ZN => n17510);
   U19749 : XNOR2_X1 port map( A => n18405, B => n17510, ZN => n17511);
   U19750 : XNOR2_X1 port map( A => n17726, B => n18621, ZN => n17514);
   U19751 : XNOR2_X1 port map( A => n17839, B => n18121, ZN => n17513);
   U19752 : XNOR2_X1 port map( A => n17514, B => n17513, ZN => n17519);
   U19753 : XNOR2_X1 port map( A => n17515, B => n912, ZN => n17517);
   U19754 : XNOR2_X1 port map( A => n18123, B => n18541, ZN => n17516);
   U19755 : XNOR2_X1 port map( A => n17517, B => n17516, ZN => n17518);
   U19756 : XNOR2_X1 port map( A => n17519, B => n17518, ZN => n18929);
   U19757 : NAND2_X1 port map( A1 => n3653, A2 => n18929, ZN => n17553);
   U19758 : XNOR2_X1 port map( A => n17811, B => n1854, ZN => n17521);
   U19759 : XNOR2_X1 port map( A => n18627, B => n17521, ZN => n17531);
   U19760 : OAI21_X1 port map( B1 => n17524, B2 => n17523, A => n17522, ZN => 
                           n17526);
   U19761 : OAI21_X1 port map( B1 => n17527, B2 => n17526, A => n17525, ZN => 
                           n17880);
   U19762 : XNOR2_X1 port map( A => n18370, B => n17880, ZN => n17529);
   U19763 : XNOR2_X1 port map( A => n18042, B => n18128, ZN => n18399);
   U19764 : INV_X1 port map( A => n18399, ZN => n17528);
   U19765 : XNOR2_X1 port map( A => n17529, B => n17528, ZN => n17530);
   U19766 : XNOR2_X1 port map( A => n17530, B => n17531, ZN => n19295);
   U19767 : XNOR2_X1 port map( A => n25379, B => n17532, ZN => n18635);
   U19768 : INV_X1 port map( A => n18635, ZN => n18160);
   U19769 : XNOR2_X1 port map( A => n18160, B => n17533, ZN => n17537);
   U19770 : XNOR2_X1 port map( A => n17807, B => n18388, ZN => n17535);
   U19771 : XNOR2_X1 port map( A => n18190, B => n2120, ZN => n17534);
   U19772 : XNOR2_X1 port map( A => n17535, B => n17534, ZN => n17536);
   U19773 : XNOR2_X2 port map( A => n17537, B => n17536, ZN => n19296);
   U19774 : OAI211_X1 port map( C1 => n19297, C2 => n18929, A => n24457, B => 
                           n19296, ZN => n17551);
   U19775 : INV_X1 port map( A => n18929, ZN => n18967);
   U19776 : NAND3_X1 port map( A1 => n17540, A2 => n17539, A3 => n17538, ZN => 
                           n17543);
   U19777 : INV_X1 port map( A => n17541, ZN => n17542);
   U19779 : XNOR2_X1 port map( A => n18472, B => n17757, ZN => n17827);
   U19780 : XNOR2_X1 port map( A => n18341, B => n18431, ZN => n18648);
   U19781 : INV_X1 port map( A => n18648, ZN => n17545);
   U19782 : XNOR2_X1 port map( A => n17545, B => n17827, ZN => n17549);
   U19783 : XNOR2_X1 port map( A => n18365, B => n3062, ZN => n17547);
   U19784 : XNOR2_X1 port map( A => n18198, B => n18429, ZN => n17546);
   U19785 : XNOR2_X1 port map( A => n17547, B => n17546, ZN => n17548);
   U19786 : XNOR2_X1 port map( A => n17549, B => n17548, ZN => n18927);
   U19789 : INV_X1 port map( A => n19531, ZN => n19272);
   U19790 : NOR2_X1 port map( A1 => n17559, A2 => n1299, ZN => n17555);
   U19791 : NOR2_X1 port map( A1 => n18919, A2 => n17555, ZN => n17561);
   U19792 : INV_X1 port map( A => n17556, ZN => n18756);
   U19794 : NAND2_X1 port map( A1 => n17558, A2 => n18756, ZN => n17560);
   U19795 : AND2_X1 port map( A1 => n20322, A2 => n20316, ZN => n17566);
   U19796 : INV_X1 port map( A => n17562, ZN => n19315);
   U19797 : NAND2_X1 port map( A1 => n18923, A2 => n19313, ZN => n17563);
   U19798 : INV_X1 port map( A => n19309, ZN => n18841);
   U19799 : NAND2_X1 port map( A1 => n18923, A2 => n24912, ZN => n19318);
   U19800 : XNOR2_X1 port map( A => n25202, B => n21273, ZN => n17952);
   U19801 : INV_X1 port map( A => n18074, ZN => n18600);
   U19802 : XNOR2_X1 port map( A => n18351, B => n18600, ZN => n17569);
   U19803 : XNOR2_X1 port map( A => n18325, B => n17819, ZN => n18524);
   U19804 : XNOR2_X1 port map( A => n18524, B => n17569, ZN => n17580);
   U19805 : INV_X1 port map( A => n17900, ZN => n17570);
   U19806 : XNOR2_X1 port map( A => n17570, B => n23225, ZN => n17578);
   U19807 : NOR2_X1 port map( A1 => n24471, A2 => n17572, ZN => n17575);
   U19808 : XNOR2_X1 port map( A => n17580, B => n17579, ZN => n18735);
   U19809 : INV_X1 port map( A => n18735, ZN => n19482);
   U19810 : XNOR2_X1 port map( A => n17581, B => n17919, ZN => n18360);
   U19811 : XNOR2_X1 port map( A => n17832, B => n17582, ZN => n18528);
   U19812 : XNOR2_X1 port map( A => n18360, B => n18528, ZN => n17586);
   U19813 : XNOR2_X1 port map( A => n24565, B => n18610, ZN => n17584);
   U19814 : XNOR2_X1 port map( A => n18032, B => n494, ZN => n17583);
   U19815 : XNOR2_X1 port map( A => n17584, B => n17583, ZN => n17585);
   U19816 : XNOR2_X1 port map( A => n17587, B => n18549, ZN => n17588);
   U19817 : XNOR2_X1 port map( A => n18646, B => n18695, ZN => n18196);
   U19818 : XNOR2_X1 port map( A => n18512, B => n23699, ZN => n17589);
   U19819 : XNOR2_X1 port map( A => n17589, B => n18513, ZN => n17591);
   U19820 : OAI21_X1 port map( B1 => n19482, B2 => n19477, A => n17594, ZN => 
                           n17896);
   U19821 : INV_X1 port map( A => n17601, ZN => n17602);
   U19822 : XNOR2_X1 port map( A => n16910, B => n18382, ZN => n17604);
   U19823 : INV_X1 port map( A => n18665, ZN => n17603);
   U19824 : XNOR2_X1 port map( A => n17604, B => n17603, ZN => n18040);
   U19825 : INV_X1 port map( A => n18040, ZN => n17605);
   U19826 : XNOR2_X1 port map( A => n17606, B => n17605, ZN => n18730);
   U19827 : INV_X1 port map( A => n18730, ZN => n18848);
   U19828 : NAND2_X1 port map( A1 => n17608, A2 => n17607, ZN => n17616);
   U19829 : NOR2_X1 port map( A1 => n17611, A2 => n17610, ZN => n17618);
   U19830 : NAND2_X1 port map( A1 => n17613, A2 => n17612, ZN => n17614);
   U19831 : NAND3_X1 port map( A1 => n17616, A2 => n17615, A3 => n17614, ZN => 
                           n17617);
   U19833 : XNOR2_X1 port map( A => n17619, B => n18018, ZN => n17636);
   U19834 : INV_X1 port map( A => n17620, ZN => n17621);
   U19835 : NOR2_X1 port map( A1 => n17622, A2 => n17621, ZN => n17627);
   U19836 : INV_X1 port map( A => n17623, ZN => n17625);
   U19837 : NOR2_X1 port map( A1 => n17625, A2 => n17624, ZN => n17626);
   U19838 : AOI21_X1 port map( B1 => n17627, B2 => n17626, A => n17629, ZN => 
                           n17628);
   U19839 : NAND2_X1 port map( A1 => n17628, A2 => n17632, ZN => n17631);
   U19840 : NAND3_X1 port map( A1 => n17633, A2 => n2561, A3 => n17629, ZN => 
                           n17630);
   U19841 : OAI211_X1 port map( C1 => n17633, C2 => n17632, A => n17631, B => 
                           n17630, ZN => n18017);
   U19842 : INV_X1 port map( A => n18017, ZN => n17634);
   U19843 : XOR2_X1 port map( A => n18157, B => n17634, Z => n17635);
   U19844 : XNOR2_X1 port map( A => n17636, B => n17635, ZN => n17639);
   U19845 : XNOR2_X1 port map( A => n18188, B => n24433, ZN => n17638);
   U19846 : NAND2_X1 port map( A1 => n19482, A2 => n17640, ZN => n17641);
   U19847 : XNOR2_X1 port map( A => n17905, B => n18541, ZN => n17981);
   U19848 : XNOR2_X1 port map( A => n17642, B => n17981, ZN => n17647);
   U19849 : XNOR2_X1 port map( A => n25000, B => n17643, ZN => n17645);
   U19850 : XNOR2_X1 port map( A => n17645, B => n17644, ZN => n17646);
   U19851 : XNOR2_X1 port map( A => n18233, B => n18067, ZN => n17918);
   U19852 : XNOR2_X1 port map( A => n18335, B => n1827, ZN => n17651);
   U19853 : XNOR2_X1 port map( A => n17649, B => n18530, ZN => n17650);
   U19854 : XNOR2_X1 port map( A => n17651, B => n17650, ZN => n17652);
   U19855 : XNOR2_X1 port map( A => n18149, B => n2040, ZN => n17654);
   U19857 : XNOR2_X1 port map( A => n17654, B => n18601, ZN => n17656);
   U19858 : XNOR2_X1 port map( A => n18022, B => n17899, ZN => n17655);
   U19859 : XNOR2_X1 port map( A => n17656, B => n17655, ZN => n17659);
   U19860 : INV_X1 port map( A => n17657, ZN => n17658);
   U19861 : INV_X1 port map( A => n18312, ZN => n17709);
   U19862 : XNOR2_X1 port map( A => n17709, B => n17969, ZN => n18626);
   U19863 : XNOR2_X1 port map( A => n18637, B => n17791, ZN => n17915);
   U19864 : XNOR2_X1 port map( A => n18413, B => n17915, ZN => n17668);
   U19865 : XNOR2_X1 port map( A => n25493, B => n24337, ZN => n17666);
   U19866 : XNOR2_X1 port map( A => n25380, B => n889, ZN => n17665);
   U19867 : XNOR2_X1 port map( A => n17666, B => n17665, ZN => n17667);
   U19869 : XNOR2_X1 port map( A => n18341, B => n18365, ZN => n17670);
   U19870 : XNOR2_X1 port map( A => n17476, B => n22986, ZN => n17669);
   U19871 : XNOR2_X1 port map( A => n17670, B => n17669, ZN => n17673);
   U19872 : INV_X1 port map( A => n17863, ZN => n17671);
   U19873 : XNOR2_X1 port map( A => n17671, B => n18200, ZN => n17672);
   U19874 : XNOR2_X1 port map( A => n18429, B => n17931, ZN => n17963);
   U19875 : NAND2_X1 port map( A1 => n25440, A2 => n19346, ZN => n17674);
   U19877 : XNOR2_X1 port map( A => n18456, B => n18636, ZN => n17851);
   U19878 : XNOR2_X1 port map( A => n17851, B => n17676, ZN => n17678);
   U19879 : INV_X1 port map( A => n18387, ZN => n17677);
   U19881 : XNOR2_X1 port map( A => n17681, B => n17680, ZN => n18481);
   U19884 : XNOR2_X1 port map( A => n18481, B => n17994, ZN => n17685);
   U19885 : XNOR2_X1 port map( A => n18269, B => n18335, ZN => n18616);
   U19886 : XNOR2_X1 port map( A => n18659, B => n1739, ZN => n17683);
   U19887 : XNOR2_X1 port map( A => n18616, B => n17683, ZN => n17684);
   U19889 : OAI22_X1 port map( A1 => n17689, A2 => n17688, B1 => n17687, B2 => 
                           n17733, ZN => n17691);
   U19890 : XNOR2_X1 port map( A => n18004, B => n18472, ZN => n17692);
   U19891 : XNOR2_X1 port map( A => n17693, B => n17692, ZN => n17697);
   U19892 : XNOR2_X1 port map( A => n17863, B => n18220, ZN => n17695);
   U19893 : XNOR2_X1 port map( A => n18431, B => n2087, ZN => n17694);
   U19894 : XNOR2_X1 port map( A => n17695, B => n17694, ZN => n17696);
   U19896 : INV_X1 port map( A => n18349, ZN => n17699);
   U19897 : XNOR2_X1 port map( A => n18601, B => n18446, ZN => n17698);
   U19898 : XNOR2_X1 port map( A => n17699, B => n17698, ZN => n17703);
   U19899 : XNOR2_X1 port map( A => n18605, B => n812, ZN => n17700);
   U19900 : XNOR2_X1 port map( A => n17701, B => n17700, ZN => n17702);
   U19903 : NAND2_X1 port map( A1 => n19037, A2 => n19451, ZN => n17712);
   U19904 : XNOR2_X1 port map( A => n18261, B => n1855, ZN => n17705);
   U19905 : XNOR2_X1 port map( A => n17705, B => n18666, ZN => n17706);
   U19906 : XNOR2_X1 port map( A => n17706, B => n18619, ZN => n17708);
   U19908 : XNOR2_X1 port map( A => n18397, B => n23620, ZN => n17710);
   U19910 : XNOR2_X1 port map( A => n18290, B => n18188, ZN => n17715);
   U19911 : XNOR2_X1 port map( A => n17911, B => n17715, ZN => n17719);
   U19912 : XNOR2_X1 port map( A => n17807, B => n18633, ZN => n17717);
   U19913 : XNOR2_X1 port map( A => n17716, B => n17717, ZN => n17718);
   U19914 : XNOR2_X1 port map( A => n18270, B => n18032, ZN => n18656);
   U19915 : INV_X1 port map( A => n17720, ZN => n18104);
   U19916 : XNOR2_X1 port map( A => n18104, B => n641, ZN => n17721);
   U19917 : XNOR2_X1 port map( A => n18656, B => n17721, ZN => n17725);
   U19918 : XNOR2_X1 port map( A => n17993, B => n18611, ZN => n17723);
   U19919 : XNOR2_X1 port map( A => n17723, B => n17722, ZN => n17724);
   U19920 : NOR2_X1 port map( A1 => n19389, A2 => n24451, ZN => n19109);
   U19921 : INV_X1 port map( A => n19109, ZN => n19387);
   U19922 : XNOR2_X1 port map( A => n17726, B => n18665, ZN => n17727);
   U19923 : XNOR2_X1 port map( A => n18124, B => n18240, ZN => n18318);
   U19924 : XNOR2_X1 port map( A => n18318, B => n17727, ZN => n17743);
   U19925 : MUX2_X1 port map( A => n17730, B => n17729, S => n25472, Z => 
                           n17732);
   U19926 : NOR2_X1 port map( A1 => n17732, A2 => n17731, ZN => n17739);
   U19927 : NOR2_X1 port map( A1 => n17734, A2 => n17733, ZN => n17736);
   U19928 : MUX2_X1 port map( A => n17737, B => n17736, S => n17735, Z => 
                           n17738);
   U19929 : NOR2_X1 port map( A1 => n17739, A2 => n17738, ZN => n17740);
   U19930 : XNOR2_X1 port map( A => n18262, B => n17740, ZN => n18671);
   U19931 : XNOR2_X1 port map( A => n18382, B => n3155, ZN => n17741);
   U19932 : XNOR2_X1 port map( A => n18671, B => n17741, ZN => n17742);
   U19933 : XNOR2_X1 port map( A => n17743, B => n17742, ZN => n19021);
   U19934 : XNOR2_X1 port map( A => n18172, B => n18370, ZN => n17745);
   U19935 : XNOR2_X1 port map( A => n18375, B => n2746, ZN => n17744);
   U19936 : XNOR2_X1 port map( A => n17744, B => n17745, ZN => n17747);
   U19937 : XNOR2_X1 port map( A => n18557, B => n18129, ZN => n18309);
   U19938 : XNOR2_X1 port map( A => n18309, B => n18683, ZN => n17746);
   U19939 : INV_X1 port map( A => n19217, ZN => n19388);
   U19940 : OAI22_X1 port map( A1 => n19387, A2 => n17762, B1 => n19389, B2 => 
                           n19388, ZN => n17766);
   U19941 : NAND2_X1 port map( A1 => n19390, A2 => n17762, ZN => n17764);
   U19942 : XNOR2_X1 port map( A => n17748, B => n18351, ZN => n18024);
   U19943 : INV_X1 port map( A => n18024, ZN => n17749);
   U19944 : XNOR2_X1 port map( A => n17897, B => n17749, ZN => n17754);
   U19945 : INV_X1 port map( A => n17816, ZN => n17750);
   U19946 : XNOR2_X1 port map( A => n18602, B => n17750, ZN => n17752);
   U19947 : XNOR2_X1 port map( A => n18096, B => n2739, ZN => n17751);
   U19948 : XNOR2_X1 port map( A => n17752, B => n17751, ZN => n17753);
   U19949 : INV_X1 port map( A => n18277, ZN => n17859);
   U19951 : XNOR2_X1 port map( A => n17755, B => n17859, ZN => n17932);
   U19952 : INV_X1 port map( A => n17757, ZN => n18506);
   U19953 : XNOR2_X1 port map( A => n18197, B => n18506, ZN => n17759);
   U19954 : XNOR2_X1 port map( A => n18476, B => n2477, ZN => n17758);
   U19955 : XNOR2_X1 port map( A => n17759, B => n17758, ZN => n17760);
   U19958 : INV_X1 port map( A => n18146, ZN => n17768);
   U19960 : XNOR2_X1 port map( A => n18418, B => n859, ZN => n17769);
   U19961 : XNOR2_X1 port map( A => n17769, B => n18447, ZN => n17770);
   U19962 : XNOR2_X1 port map( A => n17770, B => n18573, ZN => n17774);
   U19963 : XNOR2_X1 port map( A => n17772, B => n17771, ZN => n17773);
   U19964 : XNOR2_X2 port map( A => n17774, B => n17773, ZN => n19376);
   U19965 : INV_X1 port map( A => n18032, ZN => n17775);
   U19966 : XNOR2_X1 port map( A => n18103, B => n17775, ZN => n17776);
   U19967 : XNOR2_X1 port map( A => n24565, B => n18531, ZN => n18143);
   U19968 : XNOR2_X1 port map( A => n17776, B => n18143, ZN => n17778);
   U19969 : XNOR2_X1 port map( A => n18067, B => n1768, ZN => n17777);
   U19970 : XNOR2_X1 port map( A => n18435, B => n18491, ZN => n18238);
   U19971 : XNOR2_X1 port map( A => n18579, B => n18121, ZN => n17779);
   U19972 : XNOR2_X1 port map( A => n18238, B => n17779, ZN => n17782);
   U19973 : XNOR2_X1 port map( A => n18669, B => n18582, ZN => n18081);
   U19974 : XNOR2_X1 port map( A => n18665, B => n1801, ZN => n17780);
   U19975 : XNOR2_X1 port map( A => n18081, B => n17780, ZN => n17781);
   U19977 : INV_X1 port map( A => n19097, ZN => n18724);
   U19978 : XNOR2_X1 port map( A => n18276, B => n18549, ZN => n17783);
   U19979 : XNOR2_X1 port map( A => n18200, B => n18198, ZN => n18550);
   U19980 : XNOR2_X1 port map( A => n17783, B => n18550, ZN => n17787);
   U19981 : XNOR2_X1 port map( A => n18473, B => n2039, ZN => n17784);
   U19982 : XNOR2_X1 port map( A => n17785, B => n17784, ZN => n17786);
   U19983 : INV_X1 port map( A => n19370, ZN => n19364);
   U19987 : XNOR2_X1 port map( A => n17791, B => n18157, ZN => n18569);
   U19988 : XNOR2_X1 port map( A => n17792, B => n18569, ZN => n17793);
   U19989 : NAND3_X1 port map( A1 => n19222, A2 => n19364, A3 => n19371, ZN => 
                           n17802);
   U19990 : XNOR2_X1 port map( A => n18559, B => n18308, ZN => n17796);
   U19991 : XNOR2_X1 port map( A => n18310, B => n17880, ZN => n17795);
   U19992 : XNOR2_X1 port map( A => n17796, B => n17795, ZN => n17800);
   U19993 : XNOR2_X1 port map( A => n25411, B => n25194, ZN => n17798);
   U19994 : XNOR2_X1 port map( A => n17798, B => n17797, ZN => n17799);
   U19996 : XNOR2_X1 port map( A => n18675, B => n451, ZN => n17805);
   U19998 : XNOR2_X1 port map( A => n17807, B => n17806, ZN => n17808);
   U19999 : XNOR2_X1 port map( A => n17808, B => n18294, ZN => n18503);
   U20001 : XNOR2_X1 port map( A => n18512, B => n2903, ZN => n17810);
   U20002 : XNOR2_X1 port map( A => n17810, B => n18370, ZN => n17813);
   U20003 : XNOR2_X1 port map( A => n17811, B => n18172, ZN => n17812);
   U20004 : NAND2_X1 port map( A1 => n19460, A2 => n19457, ZN => n17887);
   U20005 : XNOR2_X1 port map( A => n17816, B => n18446, ZN => n17818);
   U20006 : XNOR2_X1 port map( A => n18350, B => n17817, ZN => n18253);
   U20007 : XNOR2_X1 port map( A => n18253, B => n17818, ZN => n17823);
   U20008 : XNOR2_X1 port map( A => n18523, B => n18096, ZN => n17821);
   U20009 : XNOR2_X1 port map( A => n17821, B => n17820, ZN => n17822);
   U20010 : XNOR2_X1 port map( A => n17823, B => n17822, ZN => n19456);
   U20011 : INV_X1 port map( A => n18430, ZN => n17826);
   U20012 : XNOR2_X1 port map( A => n18275, B => n887, ZN => n17825);
   U20013 : XNOR2_X1 port map( A => n17826, B => n17825, ZN => n17830);
   U20014 : INV_X1 port map( A => n18692, ZN => n17828);
   U20015 : XNOR2_X1 port map( A => n17828, B => n17827, ZN => n17829);
   U20016 : INV_X1 port map( A => n19457, ZN => n19028);
   U20017 : NAND2_X1 port map( A1 => n18976, A2 => n19028, ZN => n17831);
   U20018 : NAND3_X1 port map( A1 => n17887, A2 => n19456, A3 => n17831, ZN => 
                           n17848);
   U20019 : XNOR2_X1 port map( A => n17832, B => n18658, ZN => n17834);
   U20020 : XNOR2_X1 port map( A => n17833, B => n17834, ZN => n17838);
   U20021 : XNOR2_X1 port map( A => n18104, B => n18483, ZN => n17836);
   U20023 : XNOR2_X1 port map( A => n17836, B => n17835, ZN => n17837);
   U20024 : XNOR2_X1 port map( A => n17837, B => n17838, ZN => n17845);
   U20025 : INV_X1 port map( A => n17845, ZN => n18979);
   U20026 : XNOR2_X1 port map( A => n17839, B => n18122, ZN => n17841);
   U20027 : XNOR2_X1 port map( A => n17841, B => n18537, ZN => n17844);
   U20028 : XNOR2_X1 port map( A => n18038, B => n18489, ZN => n18259);
   U20029 : XNOR2_X1 port map( A => n18539, B => n20825, ZN => n17842);
   U20030 : XNOR2_X1 port map( A => n18259, B => n17842, ZN => n17843);
   U20031 : XNOR2_X1 port map( A => n17843, B => n17844, ZN => n18977);
   U20032 : INV_X1 port map( A => n18977, ZN => n19032);
   U20033 : NAND3_X1 port map( A1 => n24172, A2 => n18979, A3 => n19032, ZN => 
                           n17847);
   U20034 : NAND3_X1 port map( A1 => n19460, A2 => n19457, A3 => n19464, ZN => 
                           n17846);
   U20035 : NOR2_X1 port map( A1 => n19887, A2 => n25388, ZN => n17849);
   U20036 : XNOR2_X1 port map( A => n18190, B => n681, ZN => n17850);
   U20037 : INV_X1 port map( A => n18484, ZN => n17853);
   U20038 : XNOR2_X1 port map( A => n18103, B => n17853, ZN => n17854);
   U20039 : XNOR2_X1 port map( A => n17854, B => n18232, ZN => n17858);
   U20040 : XNOR2_X1 port map( A => n24568, B => n18335, ZN => n17856);
   U20041 : XNOR2_X1 port map( A => n18270, B => n2042, ZN => n17855);
   U20042 : XNOR2_X1 port map( A => n17856, B => n17855, ZN => n17857);
   U20043 : XNOR2_X1 port map( A => n18004, B => n17859, ZN => n17861);
   U20044 : XNOR2_X1 port map( A => n18198, B => n2882, ZN => n17860);
   U20045 : XNOR2_X1 port map( A => n17861, B => n17860, ZN => n17865);
   U20046 : XNOR2_X1 port map( A => n17862, B => n17863, ZN => n18645);
   U20047 : XNOR2_X1 port map( A => n18645, B => n18219, ZN => n17864);
   U20048 : XNOR2_X1 port map( A => n17864, B => n17865, ZN => n19321);
   U20049 : MUX2_X1 port map( A => n18959, B => n19470, S => n19321, Z => 
                           n17886);
   U20050 : XNOR2_X1 port map( A => n18251, B => n18448, ZN => n17868);
   U20051 : XNOR2_X1 port map( A => n18418, B => Key(172), ZN => n17866);
   U20054 : XNOR2_X1 port map( A => n18447, B => n18214, ZN => n17869);
   U20055 : XNOR2_X1 port map( A => n18098, B => n17869, ZN => n17870);
   U20056 : XNOR2_X1 port map( A => n17873, B => n18121, ZN => n18580);
   U20057 : XNOR2_X1 port map( A => n18580, B => n18238, ZN => n17879);
   U20058 : XNOR2_X1 port map( A => n25000, B => n4942, ZN => n17877);
   U20059 : XNOR2_X1 port map( A => n18262, B => n187, ZN => n17876);
   U20060 : XNOR2_X1 port map( A => n17877, B => n17876, ZN => n17878);
   U20061 : XNOR2_X1 port map( A => n17881, B => n17880, ZN => n18560);
   U20062 : XNOR2_X1 port map( A => n18130, B => n17882, ZN => n17885);
   U20063 : XNOR2_X1 port map( A => n18515, B => n25194, ZN => n18247);
   U20064 : XNOR2_X1 port map( A => n17883, B => n18247, ZN => n17884);
   U20065 : INV_X1 port map( A => n19466, ZN => n18960);
   U20066 : INV_X1 port map( A => n19460, ZN => n18739);
   U20067 : AND2_X1 port map( A1 => n17888, A2 => n17887, ZN => n17893);
   U20068 : NAND2_X1 port map( A1 => n19456, A2 => n18977, ZN => n19465);
   U20071 : NAND2_X1 port map( A1 => n17890, A2 => n19464, ZN => n17891);
   U20072 : OAI21_X2 port map( B1 => n17893, B2 => n17892, A => n17891, ZN => 
                           n19896);
   U20073 : NAND2_X1 port map( A1 => n19697, A2 => n19896, ZN => n17947);
   U20074 : INV_X1 port map( A => n17947, ZN => n17950);
   U20075 : NOR2_X1 port map( A1 => n18735, A2 => n19477, ZN => n19480);
   U20076 : XNOR2_X1 port map( A => n17897, B => n17898, ZN => n17904);
   U20077 : XNOR2_X1 port map( A => n17900, B => n17899, ZN => n17902);
   U20078 : XNOR2_X1 port map( A => n18149, B => n62, ZN => n17901);
   U20079 : XNOR2_X1 port map( A => n17902, B => n17901, ZN => n17903);
   U20080 : XNOR2_X1 port map( A => n18124, B => n17905, ZN => n18623);
   U20081 : XNOR2_X1 port map( A => n18623, B => n17906, ZN => n17910);
   U20082 : XNOR2_X1 port map( A => n17907, B => n673, ZN => n17908);
   U20083 : XNOR2_X1 port map( A => n17908, B => n18081, ZN => n17909);
   U20084 : XNOR2_X1 port map( A => n17909, B => n17910, ZN => n19502);
   U20085 : XNOR2_X1 port map( A => n17912, B => n17911, ZN => n17917);
   U20086 : XNOR2_X1 port map( A => n24433, B => n2240, ZN => n17914);
   U20087 : XNOR2_X1 port map( A => n17915, B => n17914, ZN => n17916);
   U20088 : INV_X1 port map( A => n18719, ZN => n19335);
   U20089 : XNOR2_X1 port map( A => n25006, B => n17918, ZN => n17923);
   U20090 : XNOR2_X1 port map( A => n24431, B => n18331, ZN => n17921);
   U20091 : XNOR2_X1 port map( A => n18270, B => n881, ZN => n17920);
   U20092 : XNOR2_X1 port map( A => n17921, B => n17920, ZN => n17922);
   U20093 : NOR2_X1 port map( A1 => n18986, A2 => n17924, ZN => n17940);
   U20094 : INV_X1 port map( A => n18559, ZN => n17925);
   U20095 : XNOR2_X1 port map( A => n17926, B => n17925, ZN => n18058);
   U20096 : INV_X1 port map( A => n18058, ZN => n17930);
   U20098 : XNOR2_X1 port map( A => n17927, B => n18374, ZN => n17928);
   U20099 : XNOR2_X1 port map( A => n17928, B => n18309, ZN => n17929);
   U20101 : NAND2_X1 port map( A1 => n19335, A2 => n19499, ZN => n18987);
   U20102 : XNOR2_X1 port map( A => n18476, B => n17931, ZN => n18644);
   U20103 : XNOR2_X1 port map( A => n17932, B => n18644, ZN => n17937);
   U20104 : XNOR2_X1 port map( A => n24536, B => n18693, ZN => n17935);
   U20105 : XNOR2_X1 port map( A => n18200, B => n860, ZN => n17934);
   U20106 : XNOR2_X1 port map( A => n17935, B => n17934, ZN => n17936);
   U20107 : XNOR2_X1 port map( A => n17937, B => n17936, ZN => n19498);
   U20108 : NAND2_X1 port map( A1 => n19497, A2 => n25459, ZN => n17938);
   U20109 : OAI21_X1 port map( B1 => n24370, B2 => n19896, A => n21033, ZN => 
                           n17949);
   U20110 : NAND3_X1 port map( A1 => n18970, A2 => n19297, A3 => n18967, ZN => 
                           n17941);
   U20111 : MUX2_X1 port map( A => n17947, B => n17946, S => n21038, Z => 
                           n17948);
   U20112 : XNOR2_X1 port map( A => n17951, B => n17952, ZN => n18712);
   U20113 : XNOR2_X1 port map( A => n17953, B => n18404, ZN => n17957);
   U20114 : XNOR2_X1 port map( A => n18233, B => n18658, ZN => n17955);
   U20115 : XNOR2_X1 port map( A => n18530, B => n21423, ZN => n17954);
   U20116 : XNOR2_X1 port map( A => n17955, B => n17954, ZN => n17956);
   U20117 : XNOR2_X1 port map( A => n18004, B => n17958, ZN => n17962);
   U20118 : INV_X1 port map( A => n17959, ZN => n18548);
   U20119 : XNOR2_X1 port map( A => n18548, B => n17960, ZN => n17961);
   U20120 : XNOR2_X1 port map( A => n17962, B => n17961, ZN => n17965);
   U20121 : XNOR2_X1 port map( A => n18475, B => n17963, ZN => n17964);
   U20122 : XNOR2_X1 port map( A => n17964, B => n17965, ZN => n18876);
   U20123 : XNOR2_X1 port map( A => n18465, B => n23983, ZN => n17966);
   U20124 : XNOR2_X1 port map( A => n17966, B => n18562, ZN => n17968);
   U20125 : XNOR2_X1 port map( A => n17968, B => n17967, ZN => n17973);
   U20126 : XNOR2_X1 port map( A => n18042, B => n17969, ZN => n17971);
   U20127 : XNOR2_X1 port map( A => n17970, B => n17971, ZN => n17972);
   U20128 : XNOR2_X1 port map( A => n17974, B => n18422, ZN => n17975);
   U20129 : INV_X1 port map( A => n19092, ZN => n18819);
   U20130 : AOI21_X1 port map( B1 => n18876, B2 => n19094, A => n18819, ZN => 
                           n17980);
   U20131 : XNOR2_X1 port map( A => n18227, B => n17663, ZN => n17976);
   U20132 : XNOR2_X1 port map( A => n17976, B => n24371, ZN => n17979);
   U20133 : XNOR2_X1 port map( A => n18637, B => n2190, ZN => n17977);
   U20134 : XNOR2_X1 port map( A => n17977, B => n18415, ZN => n17978);
   U20135 : XNOR2_X1 port map( A => n17979, B => n17978, ZN => n19382);
   U20136 : XNOR2_X1 port map( A => n17981, B => n17982, ZN => n17985);
   U20137 : XNOR2_X1 port map( A => n4942, B => n3084, ZN => n17983);
   U20138 : XNOR2_X1 port map( A => n18259, B => n17983, ZN => n17984);
   U20139 : NOR3_X1 port map( A1 => n24335, A2 => n19380, A3 => n19377, ZN => 
                           n17986);
   U20140 : INV_X1 port map( A => n17987, ZN => n17988);
   U20141 : XNOR2_X1 port map( A => n17988, B => n18348, ZN => n17992);
   U20142 : XNOR2_X1 port map( A => n18325, B => n765, ZN => n17989);
   U20143 : XNOR2_X1 port map( A => n17989, B => n17990, ZN => n17991);
   U20144 : XNOR2_X1 port map( A => n17993, B => n18610, ZN => n17995);
   U20145 : XNOR2_X1 port map( A => n17995, B => n17994, ZN => n17999);
   U20146 : XNOR2_X1 port map( A => n24431, B => n17582, ZN => n17997);
   U20147 : XNOR2_X1 port map( A => n18532, B => n2726, ZN => n17996);
   U20148 : XNOR2_X1 port map( A => n17997, B => n17996, ZN => n17998);
   U20150 : XNOR2_X1 port map( A => n18466, B => n23476, ZN => n18000);
   U20151 : XNOR2_X1 port map( A => n18000, B => n18370, ZN => n18001);
   U20152 : XNOR2_X1 port map( A => n18285, B => n18628, ZN => n18057);
   U20153 : XNOR2_X1 port map( A => n18057, B => n18001, ZN => n18003);
   U20154 : XNOR2_X1 port map( A => n18003, B => n18002, ZN => n18817);
   U20155 : XNOR2_X1 port map( A => n18196, B => n18005, ZN => n18008);
   U20156 : XNOR2_X1 port map( A => n18060, B => n18006, ZN => n18281);
   U20157 : XNOR2_X1 port map( A => n18363, B => n18281, ZN => n18007);
   U20158 : INV_X1 port map( A => n19360, ZN => n18009);
   U20159 : INV_X1 port map( A => n1745, ZN => n23508);
   U20160 : XNOR2_X1 port map( A => n18261, B => n23508, ZN => n18011);
   U20161 : XNOR2_X1 port map( A => n4942, B => n18539, ZN => n18010);
   U20162 : XNOR2_X1 port map( A => n18011, B => n18010, ZN => n18012);
   U20163 : INV_X1 port map( A => n18295, ZN => n18014);
   U20164 : XNOR2_X1 port map( A => n18014, B => n18294, ZN => n18016);
   U20165 : XNOR2_X1 port map( A => n18456, B => n2747, ZN => n18015);
   U20166 : XNOR2_X1 port map( A => n18016, B => n18015, ZN => n18020);
   U20167 : XNOR2_X1 port map( A => n18018, B => n18017, ZN => n18192);
   U20168 : XNOR2_X1 port map( A => n18192, B => n18390, ZN => n18019);
   U20170 : INV_X1 port map( A => n19878, ZN => n20329);
   U20171 : NOR2_X1 port map( A1 => n20554, A2 => n20329, ZN => n18136);
   U20172 : XNOR2_X1 port map( A => n18022, B => n18023, ZN => n18025);
   U20173 : XNOR2_X1 port map( A => n18024, B => n18025, ZN => n18030);
   U20174 : INV_X1 port map( A => n18326, ZN => n18026);
   U20175 : XNOR2_X1 port map( A => n18026, B => n3115, ZN => n18027);
   U20176 : XNOR2_X1 port map( A => n18028, B => n18027, ZN => n18029);
   U20177 : INV_X1 port map( A => n19595, ZN => n18037);
   U20178 : INV_X1 port map( A => n18360, ZN => n18031);
   U20179 : XNOR2_X1 port map( A => n18331, B => n18658, ZN => n18587);
   U20180 : XNOR2_X1 port map( A => n18031, B => n18587, ZN => n18036);
   U20181 : XNOR2_X1 port map( A => n18032, B => n18530, ZN => n18034);
   U20182 : XNOR2_X1 port map( A => n18356, B => n2805, ZN => n18033);
   U20183 : XNOR2_X1 port map( A => n18034, B => n18033, ZN => n18035);
   U20184 : AND2_X1 port map( A1 => n18037, A2 => n19598, ZN => n19257);
   U20185 : XNOR2_X1 port map( A => n18038, B => n18240, ZN => n18584);
   U20186 : XNOR2_X1 port map( A => n18039, B => n18584, ZN => n18041);
   U20187 : XNOR2_X1 port map( A => n18042, B => n3183, ZN => n18043);
   U20189 : XNOR2_X1 port map( A => n18045, B => n18429, ZN => n18047);
   U20190 : XNOR2_X1 port map( A => n18548, B => n18060, ZN => n18046);
   U20191 : XNOR2_X1 port map( A => n18047, B => n18046, ZN => n18048);
   U20192 : XNOR2_X1 port map( A => n18295, B => n2847, ZN => n18050);
   U20193 : XNOR2_X1 port map( A => n18052, B => n18051, ZN => n18830);
   U20195 : NAND2_X1 port map( A1 => n19597, A2 => n24079, ZN => n18053);
   U20196 : OAI21_X2 port map( B1 => n18054, B2 => n18055, A => n18053, ZN => 
                           n20330);
   U20197 : INV_X1 port map( A => n20330, ZN => n20556);
   U20198 : XNOR2_X1 port map( A => n18172, B => n2735, ZN => n18056);
   U20199 : XNOR2_X1 port map( A => n18197, B => n18277, ZN => n18062);
   U20200 : XNOR2_X1 port map( A => n18060, B => n18693, ZN => n18061);
   U20201 : XNOR2_X1 port map( A => n18062, B => n18061, ZN => n18066);
   U20202 : XNOR2_X1 port map( A => n18552, B => n18200, ZN => n18064);
   U20203 : XNOR2_X1 port map( A => n18432, B => n21169, ZN => n18063);
   U20204 : XNOR2_X1 port map( A => n18064, B => n18063, ZN => n18065);
   U20205 : XNOR2_X1 port map( A => n18067, B => n18610, ZN => n18588);
   U20206 : XNOR2_X1 port map( A => n18104, B => n18660, ZN => n18068);
   U20207 : XNOR2_X1 port map( A => n2052, B => n18068, ZN => n18072);
   U20208 : XNOR2_X1 port map( A => n24568, B => n18356, ZN => n18070);
   U20209 : XNOR2_X1 port map( A => n18270, B => n2222, ZN => n18069);
   U20210 : XNOR2_X1 port map( A => n18070, B => n18069, ZN => n18071);
   U20211 : AND2_X1 port map( A1 => n24483, A2 => n19080, ZN => n18093);
   U20212 : XNOR2_X1 port map( A => n18073, B => n18074, ZN => n18574);
   U20213 : INV_X1 port map( A => n18574, ZN => n18207);
   U20214 : XNOR2_X1 port map( A => n18251, B => n18254, ZN => n18075);
   U20215 : XNOR2_X1 port map( A => n18207, B => n18075, ZN => n18079);
   U20216 : XNOR2_X1 port map( A => n18418, B => n16, ZN => n18077);
   U20217 : XNOR2_X1 port map( A => n18077, B => n18076, ZN => n18078);
   U20218 : XNOR2_X1 port map( A => n18079, B => n18078, ZN => n19078);
   U20219 : INV_X1 port map( A => n19078, ZN => n19592);
   U20220 : INV_X1 port map( A => n19589, ZN => n18092);
   U20221 : INV_X1 port map( A => n18620, ZN => n18082);
   U20222 : XNOR2_X1 port map( A => n18082, B => n18081, ZN => n18084);
   U20223 : XNOR2_X1 port map( A => n18261, B => n677, ZN => n18083);
   U20224 : XNOR2_X1 port map( A => n24488, B => n2991, ZN => n18085);
   U20226 : AND2_X1 port map( A1 => n19591, A2 => n19077, ZN => n18806);
   U20227 : XNOR2_X1 port map( A => n18423, B => n173, ZN => n18094);
   U20228 : XNOR2_X1 port map( A => n18094, B => n18602, ZN => n18095);
   U20229 : XNOR2_X1 port map( A => n18095, B => n18323, ZN => n18100);
   U20230 : XNOR2_X1 port map( A => n18096, B => n18214, ZN => n18097);
   U20231 : XOR2_X1 port map( A => n18098, B => n18097, Z => n18099);
   U20232 : XNOR2_X1 port map( A => n18611, B => n18407, ZN => n18482);
   U20233 : XNOR2_X1 port map( A => n18101, B => n18482, ZN => n18108);
   U20234 : XNOR2_X1 port map( A => n18103, B => n18102, ZN => n18591);
   U20235 : INV_X1 port map( A => n18591, ZN => n18106);
   U20236 : XNOR2_X1 port map( A => n18104, B => n3125, ZN => n18105);
   U20237 : XNOR2_X1 port map( A => n18105, B => n18106, ZN => n18107);
   U20238 : XNOR2_X1 port map( A => n18197, B => n18365, ZN => n18110);
   U20239 : XNOR2_X1 port map( A => n18110, B => n18109, ZN => n18113);
   U20240 : INV_X1 port map( A => n19392, ZN => n23693);
   U20241 : XNOR2_X1 port map( A => n17476, B => n23693, ZN => n18111);
   U20242 : XNOR2_X1 port map( A => n18342, B => n18111, ZN => n18112);
   U20243 : XNOR2_X1 port map( A => n18112, B => n18113, ZN => n19607);
   U20247 : XNOR2_X1 port map( A => n18116, B => n18190, ZN => n18568);
   U20250 : XNOR2_X2 port map( A => n18118, B => n18119, ZN => n19233);
   U20251 : AOI21_X1 port map( B1 => n19607, B2 => n19112, A => n19233, ZN => 
                           n18120);
   U20252 : XNOR2_X1 port map( A => n18122, B => n18121, ZN => n18184);
   U20253 : XNOR2_X1 port map( A => n18317, B => n18125, ZN => n18126);
   U20254 : XNOR2_X1 port map( A => n18127, B => n18126, ZN => n19237);
   U20255 : XNOR2_X1 port map( A => n18310, B => n3089, ZN => n18132);
   U20256 : XNOR2_X1 port map( A => n18172, B => n18312, ZN => n18131);
   U20257 : XNOR2_X1 port map( A => n18132, B => n18131, ZN => n18133);
   U20258 : AOI21_X1 port map( B1 => n19610, B2 => n24310, A => n1404, ZN => 
                           n18134);
   U20259 : INV_X1 port map( A => n20328, ZN => n20089);
   U20260 : XNOR2_X1 port map( A => n18258, B => n18579, ZN => n18137);
   U20261 : XNOR2_X1 port map( A => n18538, B => n18137, ZN => n18141);
   U20262 : INV_X1 port map( A => n18237, ZN => n18139);
   U20263 : XNOR2_X1 port map( A => n18621, B => n2211, ZN => n18138);
   U20264 : XNOR2_X1 port map( A => n18139, B => n18138, ZN => n18140);
   U20265 : INV_X1 port map( A => n18142, ZN => n18144);
   U20266 : XNOR2_X1 port map( A => n18144, B => n18143, ZN => n18145);
   U20267 : XNOR2_X1 port map( A => n18447, B => n18700, ZN => n18522);
   U20268 : INV_X1 port map( A => n18522, ZN => n18148);
   U20269 : XNOR2_X1 port map( A => n18146, B => n18446, ZN => n18147);
   U20270 : XNOR2_X1 port map( A => n18149, B => n18599, ZN => n18151);
   U20271 : XNOR2_X1 port map( A => n18605, B => n2126, ZN => n18150);
   U20272 : XNOR2_X1 port map( A => n18151, B => n18150, ZN => n18152);
   U20273 : XNOR2_X1 port map( A => n18248, B => n18627, ZN => n18156);
   U20274 : XNOR2_X1 port map( A => n364, B => n18685, ZN => n18154);
   U20275 : XNOR2_X1 port map( A => n18154, B => n18153, ZN => n18155);
   U20276 : XNOR2_X1 port map( A => n18155, B => n18156, ZN => n19579);
   U20277 : INV_X1 port map( A => n19579, ZN => n19198);
   U20278 : XNOR2_X1 port map( A => n18674, B => n1869, ZN => n18158);
   U20279 : XNOR2_X1 port map( A => n18159, B => n18158, ZN => n18162);
   U20280 : XNOR2_X1 port map( A => n18160, B => n18226, ZN => n18161);
   U20281 : XNOR2_X1 port map( A => n18161, B => n18162, ZN => n19199);
   U20282 : NAND3_X1 port map( A1 => n3412, A2 => n24481, A3 => n19198, ZN => 
                           n18168);
   U20283 : XNOR2_X1 port map( A => n18473, B => n18694, ZN => n18509);
   U20284 : XNOR2_X1 port map( A => n18549, B => n21742, ZN => n18163);
   U20285 : XNOR2_X1 port map( A => n18163, B => n18648, ZN => n18164);
   U20286 : XNOR2_X1 port map( A => n18164, B => n18165, ZN => n18809);
   U20287 : INV_X1 port map( A => n18809, ZN => n19580);
   U20289 : XNOR2_X1 port map( A => n18465, B => n2100, ZN => n18169);
   U20290 : XNOR2_X1 port map( A => n18169, B => n18559, ZN => n18170);
   U20291 : XNOR2_X1 port map( A => n18170, B => n18171, ZN => n18175);
   U20292 : XNOR2_X1 port map( A => n18173, B => n18513, ZN => n18174);
   U20294 : XNOR2_X1 port map( A => n18483, B => n2826, ZN => n18177);
   U20295 : XNOR2_X1 port map( A => n18178, B => n18177, ZN => n18179);
   U20296 : XNOR2_X1 port map( A => n18582, B => n18382, ZN => n18182);
   U20297 : XNOR2_X1 port map( A => n18489, B => n1364, ZN => n18181);
   U20298 : XNOR2_X1 port map( A => n18182, B => n18181, ZN => n18186);
   U20299 : XNOR2_X1 port map( A => n18183, B => n18184, ZN => n18185);
   U20300 : XNOR2_X1 port map( A => n18185, B => n18186, ZN => n19518);
   U20301 : XNOR2_X1 port map( A => n18187, B => n18188, ZN => n18386);
   U20302 : XNOR2_X1 port map( A => n18386, B => n18189, ZN => n18194);
   U20303 : XNOR2_X1 port map( A => n18190, B => n2782, ZN => n18191);
   U20304 : XNOR2_X1 port map( A => n18192, B => n18191, ZN => n18193);
   U20305 : OAI21_X1 port map( B1 => n19518, B2 => n19522, A => n19279, ZN => 
                           n18205);
   U20306 : XNOR2_X1 port map( A => n25077, B => n18275, ZN => n18364);
   U20307 : XNOR2_X1 port map( A => n18364, B => n18196, ZN => n18204);
   U20308 : INV_X1 port map( A => n18197, ZN => n18199);
   U20309 : XNOR2_X1 port map( A => n18199, B => n18198, ZN => n18202);
   U20310 : XNOR2_X1 port map( A => n18200, B => n876, ZN => n18201);
   U20311 : XNOR2_X1 port map( A => n18202, B => n18201, ZN => n18203);
   U20312 : XNOR2_X1 port map( A => n18203, B => n18204, ZN => n19284);
   U20313 : MUX2_X1 port map( A => n18206, B => n18205, S => n19284, Z => 
                           n19723);
   U20314 : XNOR2_X1 port map( A => n18207, B => n18704, ZN => n18211);
   U20315 : XNOR2_X1 port map( A => n18350, B => n1789, ZN => n18209);
   U20316 : INV_X1 port map( A => n19720, ZN => n18212);
   U20318 : XNOR2_X1 port map( A => n18447, B => n18446, ZN => n18213);
   U20319 : XNOR2_X1 port map( A => n18213, B => n18607, ZN => n18217);
   U20320 : XNOR2_X1 port map( A => n18451, B => n886, ZN => n18215);
   U20321 : XNOR2_X1 port map( A => n18576, B => n18215, ZN => n18216);
   U20322 : INV_X1 port map( A => n19184, ZN => n19552);
   U20323 : XNOR2_X1 port map( A => n18219, B => n18218, ZN => n18224);
   U20324 : XNOR2_X1 port map( A => n18432, B => n18220, ZN => n18222);
   U20325 : XNOR2_X1 port map( A => n24383, B => n1804, ZN => n18221);
   U20326 : XNOR2_X1 port map( A => n18222, B => n18221, ZN => n18223);
   U20327 : XNOR2_X1 port map( A => n18226, B => n18225, ZN => n18231);
   U20328 : XNOR2_X1 port map( A => n18227, B => n24416, ZN => n18229);
   U20329 : XNOR2_X1 port map( A => n18229, B => n18228, ZN => n18230);
   U20330 : XNOR2_X1 port map( A => n18481, B => n18232, ZN => n18236);
   U20331 : XNOR2_X1 port map( A => n18331, B => n1792, ZN => n18234);
   U20332 : XNOR2_X1 port map( A => n18612, B => n18234, ZN => n18235);
   U20333 : XNOR2_X1 port map( A => n18237, B => n18238, ZN => n18244);
   U20334 : XNOR2_X1 port map( A => n18240, B => n18239, ZN => n18242);
   U20335 : XNOR2_X1 port map( A => n18242, B => n18241, ZN => n18243);
   U20336 : XNOR2_X1 port map( A => n18244, B => n18243, ZN => n19402);
   U20337 : NAND2_X1 port map( A1 => n19184, A2 => n19402, ZN => n19719);
   U20338 : XNOR2_X1 port map( A => n18557, B => n21944, ZN => n18245);
   U20339 : XNOR2_X1 port map( A => n18246, B => n18245, ZN => n18250);
   U20340 : XNOR2_X1 port map( A => n18247, B => n18248, ZN => n18249);
   U20341 : INV_X1 port map( A => n20560, ZN => n20023);
   U20342 : XNOR2_X1 port map( A => n18252, B => n18251, ZN => n18703);
   U20343 : XNOR2_X1 port map( A => n18703, B => n18253, ZN => n18257);
   U20344 : XNOR2_X1 port map( A => n18254, B => n2050, ZN => n18255);
   U20345 : XNOR2_X1 port map( A => n18523, B => n18605, ZN => n18425);
   U20346 : XNOR2_X1 port map( A => n18425, B => n18255, ZN => n18256);
   U20347 : XNOR2_X1 port map( A => n18258, B => n18665, ZN => n18260);
   U20348 : XNOR2_X1 port map( A => n18259, B => n18260, ZN => n18266);
   U20349 : XNOR2_X1 port map( A => n18261, B => n18539, ZN => n18264);
   U20350 : XNOR2_X1 port map( A => n18262, B => n3133, ZN => n18263);
   U20351 : XNOR2_X1 port map( A => n18264, B => n18263, ZN => n18265);
   U20352 : XNOR2_X1 port map( A => n18266, B => n18265, ZN => n19277);
   U20353 : XNOR2_X1 port map( A => n18268, B => n18267, ZN => n18274);
   U20354 : XNOR2_X1 port map( A => n18269, B => n18483, ZN => n18272);
   U20355 : XNOR2_X1 port map( A => n18270, B => n1815, ZN => n18271);
   U20356 : XNOR2_X1 port map( A => n18272, B => n18271, ZN => n18273);
   U20357 : OAI21_X1 port map( B1 => n5573, B2 => n1334, A => n19126, ZN => 
                           n18299);
   U20358 : XNOR2_X1 port map( A => n18548, B => n18275, ZN => n18279);
   U20359 : XNOR2_X1 port map( A => n18276, B => n18277, ZN => n18691);
   U20360 : INV_X1 port map( A => n18691, ZN => n18278);
   U20361 : XNOR2_X1 port map( A => n18279, B => n18278, ZN => n18282);
   U20362 : XNOR2_X1 port map( A => n18431, B => n21662, ZN => n18280);
   U20363 : XNOR2_X1 port map( A => n18287, B => n18288, ZN => n18772);
   U20364 : XNOR2_X1 port map( A => n18290, B => n18289, ZN => n18680);
   U20365 : INV_X1 port map( A => n18680, ZN => n18292);
   U20366 : XNOR2_X1 port map( A => n18292, B => n24371, ZN => n18298);
   U20367 : XNOR2_X1 port map( A => n18293, B => n18294, ZN => n18412);
   U20368 : XNOR2_X1 port map( A => n18295, B => n2881, ZN => n18296);
   U20369 : XNOR2_X1 port map( A => n18412, B => n18296, ZN => n18297);
   U20370 : XNOR2_X1 port map( A => n18298, B => n18297, ZN => n18902);
   U20371 : XNOR2_X1 port map( A => n25380, B => n21703, ZN => n18302);
   U20372 : XNOR2_X1 port map( A => n24416, B => n18302, ZN => n18304);
   U20373 : XNOR2_X1 port map( A => n18303, B => n18304, ZN => n18307);
   U20374 : XNOR2_X1 port map( A => n18305, B => n18677, ZN => n18306);
   U20375 : XNOR2_X1 port map( A => n18308, B => n18513, ZN => n18684);
   U20376 : XNOR2_X1 port map( A => n18309, B => n18684, ZN => n18316);
   U20377 : XNOR2_X1 port map( A => n18310, B => n5131, ZN => n18314);
   U20378 : XNOR2_X1 port map( A => n18312, B => n18311, ZN => n18313);
   U20379 : XNOR2_X1 port map( A => n18313, B => n18314, ZN => n18315);
   U20380 : NOR2_X1 port map( A1 => n19191, A2 => n19565, ZN => n18340);
   U20381 : XNOR2_X1 port map( A => n18318, B => n18317, ZN => n18322);
   U20382 : XNOR2_X1 port map( A => n18540, B => n18621, ZN => n18320);
   U20383 : XNOR2_X1 port map( A => n18669, B => n2761, ZN => n18319);
   U20384 : XNOR2_X1 port map( A => n18320, B => n18319, ZN => n18321);
   U20385 : XNOR2_X1 port map( A => n18324, B => n18323, ZN => n18330);
   U20386 : XNOR2_X1 port map( A => n18325, B => n18326, ZN => n18328);
   U20387 : XNOR2_X1 port map( A => n18599, B => n1920, ZN => n18327);
   U20388 : XNOR2_X1 port map( A => n18327, B => n18328, ZN => n18329);
   U20389 : XNOR2_X1 port map( A => n24565, B => n18331, ZN => n18332);
   U20390 : XNOR2_X1 port map( A => n25006, B => n18332, ZN => n18339);
   U20391 : XNOR2_X1 port map( A => n18334, B => n17582, ZN => n18337);
   U20392 : XNOR2_X1 port map( A => n18335, B => n1810, ZN => n18336);
   U20393 : XNOR2_X1 port map( A => n18337, B => n18336, ZN => n18338);
   U20394 : XNOR2_X1 port map( A => n18693, B => n18341, ZN => n18343);
   U20395 : XNOR2_X1 port map( A => n18342, B => n18343, ZN => n18347);
   U20396 : INV_X1 port map( A => n3129, ZN => n23825);
   U20397 : XNOR2_X1 port map( A => n18476, B => n23825, ZN => n18345);
   U20398 : XNOR2_X1 port map( A => n24384, B => n18695, ZN => n18344);
   U20399 : XNOR2_X1 port map( A => n18345, B => n18344, ZN => n18346);
   U20400 : XNOR2_X1 port map( A => n18347, B => n18346, ZN => n19273);
   U20401 : NOR2_X1 port map( A1 => n19566, A2 => n19273, ZN => n18395);
   U20403 : XNOR2_X1 port map( A => n18349, B => n18348, ZN => n18354);
   U20404 : XNOR2_X1 port map( A => n18423, B => n18350, ZN => n18453);
   U20405 : XNOR2_X1 port map( A => n18351, B => n4233, ZN => n18352);
   U20406 : XNOR2_X1 port map( A => n18453, B => n18352, ZN => n18353);
   U20407 : INV_X1 port map( A => n18407, ZN => n18355);
   U20408 : XNOR2_X1 port map( A => n18355, B => n18483, ZN => n18358);
   U20409 : XNOR2_X1 port map( A => n18356, B => n1776, ZN => n18357);
   U20410 : XNOR2_X1 port map( A => n18358, B => n18357, ZN => n18362);
   U20411 : XNOR2_X1 port map( A => n18359, B => n18360, ZN => n18361);
   U20412 : XNOR2_X1 port map( A => n18364, B => n18363, ZN => n18369);
   U20413 : XNOR2_X1 port map( A => n18365, B => n1891, ZN => n18366);
   U20414 : XNOR2_X1 port map( A => n18367, B => n18366, ZN => n18368);
   U20415 : XNOR2_X1 port map( A => n18369, B => n18368, ZN => n19176);
   U20416 : INV_X1 port map( A => n19176, ZN => n18777);
   U20417 : XNOR2_X1 port map( A => n18371, B => n18370, ZN => n18373);
   U20418 : XNOR2_X1 port map( A => n18372, B => n18373, ZN => n18379);
   U20419 : XNOR2_X1 port map( A => n18374, B => n23679, ZN => n18377);
   U20420 : XNOR2_X1 port map( A => n18465, B => n18375, ZN => n18376);
   U20421 : XNOR2_X1 port map( A => n18376, B => n18377, ZN => n18378);
   U20422 : XNOR2_X1 port map( A => n18380, B => n18381, ZN => n18384);
   U20423 : XNOR2_X1 port map( A => n18437, B => n18382, ZN => n18383);
   U20424 : XNOR2_X1 port map( A => n18387, B => n18386, ZN => n18392);
   U20425 : XNOR2_X1 port map( A => n18388, B => n2989, ZN => n18389);
   U20426 : XNOR2_X1 port map( A => n18390, B => n18389, ZN => n18391);
   U20427 : OAI21_X1 port map( B1 => n25195, B2 => n19176, A => n19428, ZN => 
                           n18393);
   U20428 : NAND2_X1 port map( A1 => n19183, A2 => n18393, ZN => n18394);
   U20429 : NOR2_X1 port map( A1 => n19730, A2 => n19729, ZN => n18445);
   U20430 : XNOR2_X1 port map( A => n18397, B => n25194, ZN => n18398);
   U20431 : XNOR2_X1 port map( A => n18399, B => n18398, ZN => n18403);
   U20432 : XNOR2_X1 port map( A => n18512, B => n2005, ZN => n18400);
   U20433 : XNOR2_X1 port map( A => n18401, B => n18400, ZN => n18402);
   U20434 : XNOR2_X1 port map( A => n18405, B => n18404, ZN => n18411);
   U20435 : XNOR2_X1 port map( A => n24568, B => n18407, ZN => n18409);
   U20436 : XNOR2_X1 port map( A => n18532, B => n1874, ZN => n18408);
   U20437 : XNOR2_X1 port map( A => n18409, B => n18408, ZN => n18410);
   U20438 : XNOR2_X1 port map( A => n18412, B => n18413, ZN => n18417);
   U20439 : XNOR2_X1 port map( A => n18415, B => n18414, ZN => n18416);
   U20440 : XNOR2_X1 port map( A => n18417, B => n18416, ZN => n19015);
   U20441 : INV_X1 port map( A => n19015, ZN => n19164);
   U20443 : XNOR2_X1 port map( A => n18422, B => n18421, ZN => n18427);
   U20444 : XNOR2_X1 port map( A => n18423, B => n1746, ZN => n18424);
   U20445 : XNOR2_X1 port map( A => n18424, B => n18425, ZN => n18426);
   U20447 : XNOR2_X1 port map( A => n18431, B => n1724, ZN => n18433);
   U20448 : XNOR2_X1 port map( A => n18432, B => n18433, ZN => n18434);
   U20449 : NOR2_X1 port map( A1 => n18788, A2 => n24326, ZN => n18442);
   U20450 : XNOR2_X1 port map( A => n18435, B => n18539, ZN => n18436);
   U20451 : XNOR2_X1 port map( A => n18439, B => n18438, ZN => n18440);
   U20452 : NOR2_X1 port map( A1 => n20094, A2 => n20567, ZN => n18444);
   U20453 : XNOR2_X1 port map( A => n21559, B => n21699, ZN => n18710);
   U20454 : XNOR2_X1 port map( A => n18602, B => n18446, ZN => n18450);
   U20455 : XNOR2_X1 port map( A => n18448, B => n18447, ZN => n18449);
   U20456 : XNOR2_X1 port map( A => n18450, B => n18449, ZN => n18455);
   U20457 : XNOR2_X1 port map( A => n18451, B => n24287, ZN => n18452);
   U20458 : XNOR2_X1 port map( A => n18453, B => n18452, ZN => n18454);
   U20459 : XNOR2_X1 port map( A => n18454, B => n18455, ZN => n19061);
   U20460 : INV_X1 port map( A => n19061, ZN => n19007);
   U20461 : XNOR2_X1 port map( A => n18458, B => n18457, ZN => n18462);
   U20462 : XNOR2_X1 port map( A => n18460, B => n18459, ZN => n18461);
   U20463 : XNOR2_X1 port map( A => n18465, B => n18466, ZN => n18469);
   U20464 : XNOR2_X1 port map( A => n18467, B => n2236, ZN => n18468);
   U20465 : XNOR2_X1 port map( A => n18469, B => n18468, ZN => n18470);
   U20466 : NAND3_X1 port map( A1 => n19007, A2 => n280, A3 => n1002, ZN => 
                           n18498);
   U20467 : XNOR2_X1 port map( A => n18473, B => n18472, ZN => n18474);
   U20468 : XNOR2_X1 port map( A => n18475, B => n18474, ZN => n18480);
   U20469 : XNOR2_X1 port map( A => n18476, B => n20284, ZN => n18477);
   U20470 : XNOR2_X1 port map( A => n18478, B => n18477, ZN => n18479);
   U20471 : OR3_X1 port map( A1 => n19061, A2 => n19575, A3 => n1002, ZN => 
                           n18497);
   U20472 : XNOR2_X1 port map( A => n18481, B => n18482, ZN => n18488);
   U20473 : XNOR2_X1 port map( A => n18483, B => n18531, ZN => n18486);
   U20474 : XNOR2_X1 port map( A => n18484, B => n1767, ZN => n18485);
   U20475 : XNOR2_X1 port map( A => n18486, B => n18485, ZN => n18487);
   U20476 : XNOR2_X1 port map( A => n18489, B => n2193, ZN => n18490);
   U20477 : XNOR2_X1 port map( A => n18493, B => n18494, ZN => n19059);
   U20478 : OR3_X1 port map( A1 => n19007, A2 => n24982, A3 => n19059, ZN => 
                           n18496);
   U20479 : NAND2_X1 port map( A1 => n1443, A2 => n1002, ZN => n18495);
   U20481 : XNOR2_X1 port map( A => n18499, B => n22702, ZN => n18500);
   U20482 : XNOR2_X1 port map( A => n18500, B => n18677, ZN => n18502);
   U20483 : XNOR2_X1 port map( A => n18502, B => n18501, ZN => n18504);
   U20484 : INV_X1 port map( A => n18505, ZN => n18511);
   U20485 : XNOR2_X1 port map( A => n18695, B => n2745, ZN => n18507);
   U20486 : XNOR2_X1 port map( A => n18507, B => n18506, ZN => n18508);
   U20487 : XNOR2_X1 port map( A => n18508, B => n18509, ZN => n18510);
   U20488 : INV_X1 port map( A => n3178, ZN => n22385);
   U20489 : XNOR2_X1 port map( A => n18512, B => n22385, ZN => n18514);
   U20490 : XNOR2_X1 port map( A => n18514, B => n18513, ZN => n18518);
   U20491 : XNOR2_X1 port map( A => n18516, B => n18515, ZN => n18517);
   U20492 : XNOR2_X1 port map( A => n18518, B => n18517, ZN => n18519);
   U20493 : XNOR2_X1 port map( A => n18522, B => n18521, ZN => n18527);
   U20494 : XNOR2_X1 port map( A => n18523, B => n891, ZN => n18525);
   U20495 : XNOR2_X1 port map( A => n18524, B => n18525, ZN => n18526);
   U20497 : XNOR2_X1 port map( A => n18529, B => n18528, ZN => n18536);
   U20498 : XNOR2_X1 port map( A => n18531, B => n18530, ZN => n18534);
   U20499 : XNOR2_X1 port map( A => n18532, B => n888, ZN => n18533);
   U20500 : XNOR2_X1 port map( A => n18534, B => n18533, ZN => n18535);
   U20501 : XNOR2_X1 port map( A => n18536, B => n18535, ZN => n19066);
   U20502 : XNOR2_X1 port map( A => n18538, B => n18537, ZN => n18545);
   U20503 : XNOR2_X1 port map( A => n18540, B => n18539, ZN => n18543);
   U20504 : XNOR2_X1 port map( A => n18541, B => n2034, ZN => n18542);
   U20505 : XNOR2_X1 port map( A => n18543, B => n18542, ZN => n18544);
   U20507 : XNOR2_X1 port map( A => n18548, B => n18549, ZN => n18551);
   U20508 : XNOR2_X1 port map( A => n18550, B => n18551, ZN => n18556);
   U20509 : XNOR2_X1 port map( A => n18552, B => n17476, ZN => n18555);
   U20511 : INV_X1 port map( A => n18557, ZN => n18558);
   U20512 : XNOR2_X1 port map( A => n18559, B => n18558, ZN => n18561);
   U20513 : XNOR2_X1 port map( A => n18560, B => n18561, ZN => n18566);
   U20514 : XNOR2_X1 port map( A => n364, B => n18562, ZN => n18564);
   U20515 : XNOR2_X1 port map( A => n25482, B => n1864, ZN => n18563);
   U20516 : XNOR2_X1 port map( A => n18564, B => n18563, ZN => n18565);
   U20517 : XNOR2_X1 port map( A => n18568, B => n18567, ZN => n18572);
   U20518 : XNOR2_X1 port map( A => n18570, B => n18569, ZN => n18571);
   U20519 : MUX2_X1 port map( A => n19084, B => n19417, S => n24584, Z => 
                           n18595);
   U20520 : XNOR2_X1 port map( A => n18574, B => n18573, ZN => n18578);
   U20521 : XNOR2_X1 port map( A => n18576, B => n18575, ZN => n18577);
   U20522 : XNOR2_X1 port map( A => n18582, B => n1758, ZN => n18583);
   U20523 : XNOR2_X1 port map( A => n18584, B => n18583, ZN => n18585);
   U20524 : INV_X1 port map( A => n19420, ZN => n19083);
   U20525 : AND2_X1 port map( A1 => n19088, A2 => n18586, ZN => n18594);
   U20526 : XNOR2_X1 port map( A => n18588, B => n18587, ZN => n18593);
   U20527 : INV_X1 port map( A => n899, ZN => n22739);
   U20528 : XNOR2_X1 port map( A => n24565, B => n22739, ZN => n18590);
   U20529 : XNOR2_X1 port map( A => n18591, B => n18590, ZN => n18592);
   U20530 : NAND3_X1 port map( A1 => n18597, A2 => n25195, A3 => n18777, ZN => 
                           n18598);
   U20531 : XNOR2_X1 port map( A => n18600, B => n18599, ZN => n18604);
   U20532 : XNOR2_X1 port map( A => n18602, B => n18601, ZN => n18603);
   U20533 : XNOR2_X1 port map( A => n18603, B => n18604, ZN => n18609);
   U20534 : XNOR2_X1 port map( A => n18605, B => n2772, ZN => n18606);
   U20535 : XNOR2_X1 port map( A => n18607, B => n18606, ZN => n18608);
   U20536 : XNOR2_X1 port map( A => n18609, B => n18608, ZN => n19436);
   U20537 : XNOR2_X1 port map( A => n18611, B => n18610, ZN => n18614);
   U20538 : XNOR2_X1 port map( A => n18613, B => n18614, ZN => n18618);
   U20539 : XNOR2_X1 port map( A => n18616, B => n18615, ZN => n18617);
   U20540 : XNOR2_X1 port map( A => n18620, B => n18619, ZN => n18625);
   U20541 : XNOR2_X1 port map( A => n18621, B => n1924, ZN => n18622);
   U20542 : XNOR2_X1 port map( A => n18623, B => n18622, ZN => n18624);
   U20543 : XNOR2_X1 port map( A => n18627, B => n18626, ZN => n18632);
   U20544 : XNOR2_X1 port map( A => n25482, B => n2757, ZN => n18630);
   U20545 : XNOR2_X1 port map( A => n18630, B => n18629, ZN => n18631);
   U20546 : INV_X1 port map( A => n19438, ZN => n18642);
   U20547 : XNOR2_X1 port map( A => n18635, B => n18634, ZN => n18641);
   U20548 : XNOR2_X1 port map( A => n18637, B => n25493, ZN => n18639);
   U20549 : XNOR2_X1 port map( A => n18639, B => n18638, ZN => n18640);
   U20550 : XNOR2_X1 port map( A => n18641, B => n18640, ZN => n18832);
   U20551 : OAI21_X1 port map( B1 => n5007, B2 => n19245, A => n18643, ZN => 
                           n18655);
   U20552 : XNOR2_X1 port map( A => n18645, B => n18644, ZN => n18650);
   U20553 : XNOR2_X1 port map( A => n18646, B => n20690, ZN => n18647);
   U20554 : XNOR2_X1 port map( A => n18648, B => n18647, ZN => n18649);
   U20555 : XNOR2_X1 port map( A => n18650, B => n18649, ZN => n18834);
   U20556 : INV_X1 port map( A => n18834, ZN => n19081);
   U20557 : OAI21_X1 port map( B1 => n19081, B2 => n25260, A => n18651, ZN => 
                           n18653);
   U20558 : NOR2_X1 port map( A1 => n18653, A2 => n19435, ZN => n18654);
   U20559 : NOR2_X1 port map( A1 => n24835, A2 => n20569, ZN => n18706);
   U20560 : XNOR2_X1 port map( A => n18656, B => n18657, ZN => n18664);
   U20561 : XNOR2_X1 port map( A => n18659, B => n18658, ZN => n18662);
   U20562 : XNOR2_X1 port map( A => n18660, B => n1757, ZN => n18661);
   U20563 : XNOR2_X1 port map( A => n18662, B => n18661, ZN => n18663);
   U20564 : INV_X1 port map( A => n18690, ZN => n19170);
   U20565 : XNOR2_X1 port map( A => n18666, B => n18665, ZN => n18668);
   U20567 : XNOR2_X1 port map( A => n18669, B => n2990, ZN => n18670);
   U20568 : XNOR2_X1 port map( A => n18671, B => n18670, ZN => n18672);
   U20569 : XNOR2_X1 port map( A => n18674, B => n18675, ZN => n18676);
   U20570 : XNOR2_X1 port map( A => n18677, B => n18676, ZN => n18682);
   U20571 : XNOR2_X1 port map( A => n18678, B => n2031, ZN => n18679);
   U20572 : XNOR2_X1 port map( A => n18684, B => n18683, ZN => n18689);
   U20573 : XNOR2_X1 port map( A => n18685, B => n1863, ZN => n18686);
   U20574 : XNOR2_X1 port map( A => n18687, B => n18686, ZN => n18688);
   U20575 : XNOR2_X1 port map( A => n18688, B => n18689, ZN => n19406);
   U20576 : INV_X1 port map( A => n19406, ZN => n19169);
   U20577 : XNOR2_X1 port map( A => n18692, B => n18691, ZN => n18699);
   U20578 : XNOR2_X1 port map( A => n18694, B => n18693, ZN => n18697);
   U20579 : XNOR2_X1 port map( A => n18695, B => n2044, ZN => n18696);
   U20580 : XNOR2_X1 port map( A => n18697, B => n18696, ZN => n18698);
   U20582 : NOR2_X1 port map( A1 => n20617, A2 => n20615, ZN => n18705);
   U20583 : AOI22_X1 port map( A1 => n18706, A2 => n20614, B1 => n24338, B2 => 
                           n18705, ZN => n18708);
   U20584 : NAND2_X1 port map( A1 => n24338, A2 => n20623, ZN => n18707);
   U20585 : OAI211_X1 port map( C1 => n20619, C2 => n24338, A => n18708, B => 
                           n18707, ZN => n20742);
   U20586 : XNOR2_X1 port map( A => n20742, B => n2190, ZN => n18709);
   U20587 : XNOR2_X1 port map( A => n18710, B => n18709, ZN => n18711);
   U20589 : NAND2_X1 port map( A1 => n19357, A2 => n19444, ZN => n18717);
   U20590 : OR3_X1 port map( A1 => n19357, A2 => n19451, A3 => n19452, ZN => 
                           n18716);
   U20591 : NAND2_X1 port map( A1 => n25002, A2 => n19446, ZN => n18714);
   U20592 : NAND2_X1 port map( A1 => n18990, A2 => n19445, ZN => n19351);
   U20593 : INV_X1 port map( A => n19498, ZN => n18718);
   U20595 : NAND3_X1 port map( A1 => n18724, A2 => n19371, A3 => n24361, ZN => 
                           n18725);
   U20596 : NAND2_X1 port map( A1 => n19345, A2 => n19346, ZN => n18728);
   U20597 : OAI21_X1 port map( B1 => n19487, B2 => n240, A => n18727, ZN => 
                           n19208);
   U20598 : NAND2_X1 port map( A1 => n19230, A2 => n18729, ZN => n18743);
   U20599 : NAND2_X1 port map( A1 => n18730, A2 => n19477, ZN => n18733);
   U20600 : INV_X1 port map( A => n19478, ZN => n18731);
   U20601 : NAND2_X1 port map( A1 => n19476, A2 => n18731, ZN => n18732);
   U20602 : MUX2_X1 port map( A => n18733, B => n18732, S => n19482, Z => 
                           n18738);
   U20603 : INV_X1 port map( A => n18734, ZN => n18974);
   U20604 : NOR2_X1 port map( A1 => n18735, A2 => n18974, ZN => n18736);
   U20605 : OAI21_X1 port map( B1 => n18971, B2 => n18736, A => n19478, ZN => 
                           n18737);
   U20606 : NAND3_X1 port map( A1 => n18739, A2 => n18979, A3 => n19028, ZN => 
                           n18740);
   U20608 : OAI21_X1 port map( B1 => n20191, B2 => n20185, A => n25478, ZN => 
                           n18742);
   U20610 : XNOR2_X1 port map( A => n21135, B => n1745, ZN => n18746);
   U20611 : NAND2_X1 port map( A1 => n20336, A2 => n20669, ZN => n18744);
   U20612 : NAND2_X1 port map( A1 => n18744, A2 => n20668, ZN => n18745);
   U20613 : NAND2_X1 port map( A1 => n19309, A2 => n19311, ZN => n18921);
   U20614 : NAND2_X1 port map( A1 => n18921, A2 => n19313, ZN => n18748);
   U20615 : NOR2_X1 port map( A1 => n19309, A2 => n19312, ZN => n18747);
   U20616 : NOR2_X1 port map( A1 => n3284, A2 => n19555, ZN => n18750);
   U20617 : INV_X1 port map( A => n19556, ZN => n19558);
   U20618 : MUX2_X1 port map( A => n18752, B => n18750, S => n19558, Z => 
                           n18754);
   U20619 : OAI21_X1 port map( B1 => n19560, B2 => n4262, A => n3284, ZN => 
                           n18751);
   U20620 : NOR2_X1 port map( A1 => n18752, A2 => n18751, ZN => n18753);
   U20621 : INV_X1 port map( A => n19266, ZN => n18917);
   U20622 : NOR2_X1 port map( A1 => n18919, A2 => n18917, ZN => n18758);
   U20623 : NOR2_X1 port map( A1 => n18756, A2 => n24386, ZN => n18757);
   U20624 : NOR2_X1 port map( A1 => n18758, A2 => n18757, ZN => n18760);
   U20625 : MUX2_X1 port map( A => n19531, B => n19534, S => n24393, Z => 
                           n18763);
   U20626 : INV_X1 port map( A => n18762, ZN => n19530);
   U20627 : NAND2_X1 port map( A1 => n19535, A2 => n19532, ZN => n18764);
   U20629 : NOR2_X1 port map( A1 => n24441, A2 => n18767, ZN => n18770);
   U20631 : INV_X1 port map( A => n18772, ZN => n19540);
   U20632 : AOI22_X1 port map( A1 => n5573, A2 => n19539, B1 => n19540, B2 => 
                           n1334, ZN => n18773);
   U20633 : MUX2_X1 port map( A => n19546, B => n19185, S => n19548, Z => 
                           n18775);
   U20635 : NAND3_X1 port map( A1 => n24758, A2 => n19177, A3 => n19179, ZN => 
                           n18781);
   U20636 : AOI21_X1 port map( B1 => n19427, B2 => n19177, A => n1361, ZN => 
                           n18776);
   U20637 : OAI21_X1 port map( B1 => n19183, B2 => n19427, A => n18776, ZN => 
                           n18780);
   U20638 : NOR2_X1 port map( A1 => n18777, A2 => n19428, ZN => n18778);
   U20639 : NAND2_X1 port map( A1 => n19183, A2 => n18778, ZN => n18779);
   U20640 : INV_X1 port map( A => n19173, ZN => n19411);
   U20641 : AND2_X1 port map( A1 => n19413, A2 => n19406, ZN => n19172);
   U20642 : INV_X1 port map( A => n19172, ZN => n18784);
   U20644 : NOR2_X1 port map( A1 => n20060, A2 => n25088, ZN => n19641);
   U20645 : NAND2_X1 port map( A1 => n20470, A2 => n19641, ZN => n18803);
   U20646 : INV_X1 port map( A => n24326, ZN => n18899);
   U20647 : INV_X1 port map( A => n18788, ZN => n19396);
   U20648 : OAI21_X1 port map( B1 => n18790, B2 => n18899, A => n18789, ZN => 
                           n18792);
   U20649 : NOR2_X1 port map( A1 => n19191, A2 => n1053, ZN => n18794);
   U20650 : NAND2_X1 port map( A1 => n19192, A2 => n19568, ZN => n18793);
   U20651 : INV_X1 port map( A => n19518, ZN => n18795);
   U20652 : AOI22_X1 port map( A1 => n18897, A2 => n19522, B1 => n19523, B2 => 
                           n19521, ZN => n18799);
   U20653 : INV_X1 port map( A => n19284, ZN => n19519);
   U20654 : NAND2_X1 port map( A1 => n19279, A2 => n19519, ZN => n18797);
   U20655 : MUX2_X1 port map( A => n18797, B => n18796, S => n19518, Z => 
                           n18798);
   U20656 : OAI21_X1 port map( B1 => n25490, B2 => n19928, A => n20062, ZN => 
                           n18800);
   U20658 : NAND2_X1 port map( A1 => n18800, A2 => n5115, ZN => n18802);
   U20659 : INV_X1 port map( A => n20060, ZN => n19121);
   U20660 : NAND3_X1 port map( A1 => n20062, A2 => n20055, A3 => n19121, ZN => 
                           n18801);
   U20661 : XNOR2_X1 port map( A => n21084, B => n21212, ZN => n21696);
   U20662 : NAND2_X1 port map( A1 => n19233, A2 => n19607, ZN => n19113);
   U20663 : NOR2_X1 port map( A1 => n19237, A2 => n19112, ZN => n18804);
   U20664 : NOR2_X1 port map( A1 => n19113, A2 => n18804, ZN => n18805);
   U20665 : INV_X1 port map( A => n20359, ZN => n20911);
   U20666 : INV_X1 port map( A => n19591, ZN => n19250);
   U20667 : INV_X1 port map( A => n18806, ZN => n18807);
   U20668 : INV_X1 port map( A => n19199, ZN => n19581);
   U20669 : MUX2_X1 port map( A => n19198, B => n18809, S => n19581, Z => 
                           n18811);
   U20670 : INV_X1 port map( A => n19105, ZN => n19582);
   U20671 : INV_X1 port map( A => n19107, ZN => n19586);
   U20672 : OAI21_X1 port map( B1 => n19582, B2 => n19581, A => n19202, ZN => 
                           n18810);
   U20673 : NOR2_X1 port map( A1 => n24909, A2 => n19021, ZN => n19108);
   U20674 : INV_X1 port map( A => n19108, ZN => n18815);
   U20676 : OAI21_X1 port map( B1 => n24931, B2 => n19389, A => n25052, ZN => 
                           n18813);
   U20677 : AND2_X1 port map( A1 => n19386, A2 => n19217, ZN => n19631);
   U20678 : INV_X1 port map( A => n19021, ZN => n19630);
   U20679 : NAND2_X1 port map( A1 => n19631, A2 => n19630, ZN => n18814);
   U20680 : AOI22_X1 port map( A1 => n20911, A2 => n20909, B1 => n20913, B2 => 
                           n20491, ZN => n20363);
   U20681 : INV_X1 port map( A => n19041, ZN => n18816);
   U20682 : NAND2_X1 port map( A1 => n18817, A2 => n25392, ZN => n18818);
   U20685 : OAI21_X1 port map( B1 => n19380, B2 => n24452, A => n18819, ZN => 
                           n18821);
   U20686 : NOR2_X1 port map( A1 => n19382, A2 => n18876, ZN => n19205);
   U20688 : NAND3_X1 port map( A1 => n25067, A2 => n24318, A3 => n19094, ZN => 
                           n18820);
   U20689 : OAI21_X1 port map( B1 => n18821, B2 => n19205, A => n18820, ZN => 
                           n18823);
   U20690 : NOR2_X1 port map( A1 => n19379, A2 => n19377, ZN => n18822);
   U20692 : NAND2_X1 port map( A1 => n20487, A2 => n20909, ZN => n18824);
   U20693 : NAND2_X1 port map( A1 => n18824, A2 => n347, ZN => n18825);
   U20695 : MUX2_X1 port map( A => n18826, B => n19406, S => n19408, Z => 
                           n18827);
   U20696 : INV_X1 port map( A => n19417, ZN => n19087);
   U20697 : NAND2_X1 port map( A1 => n19419, A2 => n19084, ZN => n18829);
   U20698 : NOR2_X1 port map( A1 => n19166, A2 => n19084, ZN => n18828);
   U20699 : NAND2_X1 port map( A1 => n25423, A2 => n361, ZN => n18833);
   U20700 : INV_X1 port map( A => n19065, ZN => n19241);
   U20701 : INV_X1 port map( A => n19066, ZN => n19615);
   U20702 : MUX2_X1 port map( A => n18837, B => n18836, S => n19615, Z => 
                           n18838);
   U20703 : INV_X1 port map( A => n20478, ZN => n18839);
   U20705 : XNOR2_X1 port map( A => n21572, B => n25073, ZN => n20954);
   U20706 : INV_X1 port map( A => n18959, ZN => n18944);
   U20708 : INV_X1 port map( A => n19470, ZN => n19322);
   U20709 : INV_X1 port map( A => n19321, ZN => n19467);
   U20710 : AOI21_X1 port map( B1 => n18842, B2 => n18925, A => n18841, ZN => 
                           n18845);
   U20711 : OAI22_X1 port map( A1 => n18923, A2 => n18843, B1 => n19317, B2 => 
                           n24912, ZN => n18844);
   U20712 : NOR2_X1 port map( A1 => n357, A2 => n19501, ZN => n18847);
   U20713 : INV_X1 port map( A => n19480, ZN => n18851);
   U20714 : NOR2_X1 port map( A1 => n18974, A2 => n19476, ZN => n18849);
   U20715 : NAND2_X1 port map( A1 => n18971, A2 => n19479, ZN => n18850);
   U20716 : AND2_X1 port map( A1 => n19658, A2 => n20068, ZN => n19194);
   U20717 : AOI21_X1 port map( B1 => n20071, B2 => n19660, A => n19194, ZN => 
                           n18859);
   U20718 : INV_X1 port map( A => n19329, ZN => n18935);
   U20719 : MUX2_X1 port map( A => n24583, B => n25566, S => n18935, Z => 
                           n18855);
   U20720 : NAND2_X1 port map( A1 => n5736, A2 => n18934, ZN => n18854);
   U20721 : AND2_X1 port map( A1 => n19329, A2 => n19328, ZN => n18938);
   U20722 : INV_X1 port map( A => n19195, ZN => n19850);
   U20723 : NAND2_X1 port map( A1 => n19297, A2 => n24427, ZN => n18856);
   U20724 : NAND3_X1 port map( A1 => n24457, A2 => n19297, A3 => n356, ZN => 
                           n18857);
   U20725 : INV_X1 port map( A => n20068, ZN => n20073);
   U20726 : AOI21_X1 port map( B1 => n19849, B2 => n19658, A => n20073, ZN => 
                           n18858);
   U20728 : XNOR2_X1 port map( A => n20954, B => n25222, ZN => n18860);
   U20730 : NAND2_X1 port map( A1 => n18865, A2 => n18864, ZN => n18866);
   U20732 : INV_X1 port map( A => n19596, ZN => n18871);
   U20733 : OAI21_X1 port map( B1 => n18037, B2 => n19601, A => n19254, ZN => 
                           n18874);
   U20734 : NAND3_X1 port map( A1 => n19071, A2 => n18871, A3 => n19601, ZN => 
                           n18872);
   U20735 : NOR2_X1 port map( A1 => n20289, A2 => n19668, ZN => n18887);
   U20736 : OAI22_X1 port map( A1 => n24335, A2 => n24318, B1 => n24452, B2 => 
                           n19094, ZN => n19206);
   U20737 : NAND2_X1 port map( A1 => n19382, A2 => n18876, ZN => n19093);
   U20740 : MUX2_X1 port map( A => n19581, B => n19580, S => n19198, Z => 
                           n18882);
   U20741 : NAND2_X1 port map( A1 => n19105, A2 => n19107, ZN => n18881);
   U20742 : INV_X1 port map( A => n21009, ZN => n20530);
   U20743 : INV_X1 port map( A => n21008, ZN => n20528);
   U20744 : INV_X1 port map( A => n19066, ZN => n18883);
   U20745 : INV_X1 port map( A => n19067, ZN => n19614);
   U20746 : NAND2_X1 port map( A1 => n18884, A2 => n19239, ZN => n18885);
   U20748 : INV_X1 port map( A => n19546, ZN => n18889);
   U20751 : INV_X1 port map( A => n19402, ZN => n19549);
   U20752 : NAND3_X1 port map( A1 => n19552, A2 => n19549, A3 => n19186, ZN => 
                           n18892);
   U20753 : NAND3_X1 port map( A1 => n24929, A2 => n18889, A3 => n1711, ZN => 
                           n18891);
   U20754 : NAND3_X1 port map( A1 => n24929, A2 => n19185, A3 => n19546, ZN => 
                           n18890);
   U20755 : NAND2_X1 port map( A1 => n18894, A2 => n19522, ZN => n18898);
   U20756 : NOR2_X1 port map( A1 => n19526, A2 => n19523, ZN => n18896);
   U20757 : NAND2_X1 port map( A1 => n20126, A2 => n20309, ZN => n20548);
   U20758 : NAND2_X1 port map( A1 => n19540, A2 => n19543, ZN => n18904);
   U20759 : OAI21_X1 port map( B1 => n1334, B2 => n19126, A => n19275, ZN => 
                           n18903);
   U20760 : INV_X1 port map( A => n19276, ZN => n18905);
   U20762 : NOR2_X1 port map( A1 => n19191, A2 => n363, ZN => n18908);
   U20763 : NAND2_X1 port map( A1 => n19555, A2 => n24421, ZN => n18912);
   U20764 : INV_X1 port map( A => n19290, ZN => n19554);
   U20765 : NAND3_X1 port map( A1 => n19554, A2 => n19559, A3 => n19555, ZN => 
                           n18911);
   U20766 : INV_X1 port map( A => n20127, ZN => n20543);
   U20767 : NAND3_X1 port map( A1 => n20130, A2 => n20545, A3 => n20543, ZN => 
                           n18913);
   U20768 : XNOR2_X1 port map( A => n21678, B => n21597, ZN => n21116);
   U20769 : INV_X1 port map( A => n19263, ZN => n19150);
   U20770 : INV_X1 port map( A => n18921, ZN => n18922);
   U20771 : NAND3_X1 port map( A1 => n18923, A2 => n5371, A3 => n19313, ZN => 
                           n18924);
   U20772 : OAI21_X1 port map( B1 => n18925, B2 => n19312, A => n18924, ZN => 
                           n18926);
   U20773 : INV_X1 port map( A => n18928, ZN => n18931);
   U20774 : AND2_X1 port map( A1 => n19297, A2 => n18929, ZN => n19301);
   U20775 : INV_X1 port map( A => n19301, ZN => n18930);
   U20776 : AOI22_X2 port map( A1 => n18968, A2 => n18932, B1 => n18930, B2 => 
                           n18931, ZN => n19785);
   U20777 : MUX2_X1 port map( A => n19684, B => n19984, S => n19785, Z => 
                           n18942);
   U20778 : NOR2_X1 port map( A1 => n18934, A2 => n18933, ZN => n18937);
   U20779 : NOR2_X2 port map( A1 => n18941, A2 => n18940, ZN => n19987);
   U20780 : NOR2_X1 port map( A1 => n18942, A2 => n24979, ZN => n18955);
   U20781 : NOR2_X1 port map( A1 => n19472, A2 => n19467, ZN => n18943);
   U20782 : MUX2_X1 port map( A => n19466, B => n18943, S => n18959, Z => 
                           n18946);
   U20783 : INV_X1 port map( A => n19472, ZN => n18956);
   U20784 : NAND2_X1 port map( A1 => n19984, A2 => n24464, ZN => n18953);
   U20786 : NAND2_X1 port map( A1 => n19303, A2 => n18947, ZN => n18948);
   U20787 : AND2_X1 port map( A1 => n19306, A2 => n18948, ZN => n18952);
   U20789 : NOR2_X1 port map( A1 => n25364, A2 => n19128, ZN => n18950);
   U20790 : AOI22_X1 port map( A1 => n24441, A2 => n18950, B1 => n18949, B2 => 
                           n24324, ZN => n18951);
   U20791 : OAI22_X1 port map( A1 => n19986, A2 => n18953, B1 => n24315, B2 => 
                           n19786, ZN => n18954);
   U20792 : NOR2_X1 port map( A1 => n18955, A2 => n18954, ZN => n20767);
   U20794 : NOR2_X1 port map( A1 => n19466, A2 => n19321, ZN => n18957);
   U20796 : AOI21_X1 port map( B1 => n18962, B2 => n18961, A => n18960, ZN => 
                           n18963);
   U20798 : NAND2_X1 port map( A1 => n19296, A2 => n24427, ZN => n18966);
   U20799 : AND2_X1 port map( A1 => n4075, A2 => n18966, ZN => n18969);
   U20801 : NAND2_X1 port map( A1 => n18971, A2 => n19476, ZN => n18972);
   U20802 : INV_X1 port map( A => n19459, ZN => n18976);
   U20803 : NAND2_X1 port map( A1 => n18976, A2 => n19457, ZN => n19030);
   U20804 : NAND3_X1 port map( A1 => n19030, A2 => n18979, A3 => n18977, ZN => 
                           n18981);
   U20805 : OAI21_X1 port map( B1 => n19030, B2 => n19464, A => n18978, ZN => 
                           n18980);
   U20806 : AOI21_X2 port map( B1 => n18980, B2 => n18981, A => n19029, ZN => 
                           n20019);
   U20807 : OAI211_X1 port map( C1 => n25459, C2 => n19501, A => n358, B => 
                           n19334, ZN => n18988);
   U20808 : NAND2_X1 port map( A1 => n19500, A2 => n18983, ZN => n18984);
   U20809 : OAI211_X1 port map( C1 => n18987, C2 => n19501, A => n18988, B => 
                           n18984, ZN => n18985);
   U20810 : NOR2_X1 port map( A1 => n20136, A2 => n20014, ZN => n18991);
   U20812 : NAND2_X1 port map( A1 => n18991, A2 => n19755, ZN => n20925);
   U20813 : XNOR2_X1 port map( A => n20767, B => n21523, ZN => n20439);
   U20814 : XNOR2_X1 port map( A => n21116, B => n20439, ZN => n19054);
   U20815 : NAND2_X1 port map( A1 => n20317, A2 => n18994, ZN => n18993);
   U20816 : INV_X1 port map( A => n19889, ZN => n20320);
   U20818 : MUX2_X1 port map( A => n18993, B => n18992, S => n20319, Z => 
                           n18997);
   U20819 : AND2_X1 port map( A1 => n19714, A2 => n20316, ZN => n18995);
   U20820 : AOI22_X1 port map( A1 => n19888, A2 => n24917, B1 => n18995, B2 => 
                           n341, ZN => n18996);
   U20822 : NOR2_X1 port map( A1 => n19417, A2 => n19418, ZN => n18999);
   U20823 : AOI22_X1 port map( A1 => n19000, A2 => n18998, B1 => n24584, B2 => 
                           n18999, ZN => n19001);
   U20824 : NOR2_X1 port map( A1 => n18385, A2 => n19177, ZN => n19180);
   U20825 : AND2_X1 port map( A1 => n19003, A2 => n19177, ZN => n19005);
   U20826 : OAI211_X1 port map( C1 => n19179, C2 => n19760, A => n19176, B => 
                           n25195, ZN => n19004);
   U20827 : NOR2_X1 port map( A1 => n20536, A2 => n20537, ZN => n19689);
   U20828 : OAI21_X1 port map( B1 => n280, B2 => n354, A => n1002, ZN => n19006
                           );
   U20830 : INV_X1 port map( A => n20537, ZN => n19011);
   U20831 : MUX2_X1 port map( A => n19413, B => n19407, S => n19170, Z => 
                           n19010);
   U20832 : NAND2_X1 port map( A1 => n19173, A2 => n19413, ZN => n19009);
   U20833 : OAI21_X1 port map( B1 => n20149, B2 => n19011, A => n20447, ZN => 
                           n19012);
   U20835 : MUX2_X1 port map( A => n18834, B => n361, S => n19438, Z => n19013)
                           ;
   U20836 : NAND2_X1 port map( A1 => n20533, A2 => n20149, ZN => n19019);
   U20837 : NAND2_X1 port map( A1 => n19397, A2 => n19164, ZN => n19014);
   U20838 : NAND2_X1 port map( A1 => n19016, A2 => n19396, ZN => n19017);
   U20839 : INV_X1 port map( A => n20445, ZN => n19018);
   U20840 : XNOR2_X1 port map( A => n21679, B => n21639, ZN => n21096);
   U20841 : NAND2_X1 port map( A1 => n24451, A2 => n19021, ZN => n19391);
   U20842 : NAND2_X1 port map( A1 => n19384, A2 => n25052, ZN => n19022);
   U20843 : OAI21_X1 port map( B1 => n19024, B2 => n19490, A => n19023, ZN => 
                           n19027);
   U20844 : MUX2_X1 port map( A => n19345, B => n240, S => n19488, Z => n19025)
                           ;
   U20845 : NOR2_X1 port map( A1 => n19025, A2 => n25473, ZN => n19026);
   U20848 : NAND2_X1 port map( A1 => n19452, A2 => n19444, ZN => n19039);
   U20849 : NOR2_X1 port map( A1 => n18816, A2 => n19210, ZN => n19043);
   U20850 : MUX2_X1 port map( A => n19043, B => n19042, S => n24312, Z => 
                           n19046);
   U20851 : NAND2_X1 port map( A1 => n19361, A2 => n19210, ZN => n19044);
   U20852 : OAI22_X1 port map( A1 => n19211, A2 => n19044, B1 => n19103, B2 => 
                           n24312, ZN => n19045);
   U20853 : NAND2_X1 port map( A1 => n19047, A2 => n20297, ZN => n19048);
   U20854 : INV_X1 port map( A => n2126, ZN => n19051);
   U20855 : XNOR2_X1 port map( A => n20870, B => n19051, ZN => n19052);
   U20856 : XNOR2_X1 port map( A => n21096, B => n19052, ZN => n19053);
   U20859 : OAI21_X1 port map( B1 => n19615, B2 => n24606, A => n355, ZN => 
                           n19070);
   U20860 : NOR2_X1 port map( A1 => n19065, A2 => n19064, ZN => n19243);
   U20861 : NAND2_X1 port map( A1 => n19243, A2 => n25086, ZN => n19069);
   U20862 : NAND2_X1 port map( A1 => n19067, A2 => n19613, ZN => n19068);
   U20863 : NOR2_X1 port map( A1 => n18037, A2 => n19602, ZN => n19076);
   U20864 : NOR3_X1 port map( A1 => n19071, A2 => n18037, A3 => n19598, ZN => 
                           n19072);
   U20865 : NOR2_X1 port map( A1 => n19073, A2 => n19072, ZN => n19074);
   U20866 : NOR2_X1 port map( A1 => n19591, A2 => n19077, ZN => n19079);
   U20867 : INV_X1 port map( A => n20497, ZN => n19904);
   U20868 : NAND3_X1 port map( A1 => n24887, A2 => n20224, A3 => n20501, ZN => 
                           n19090);
   U20869 : NAND3_X1 port map( A1 => n24584, A2 => n19084, A3 => n19083, ZN => 
                           n19086);
   U20870 : NAND3_X1 port map( A1 => n19166, A2 => n19420, A3 => n19418, ZN => 
                           n19085);
   U20871 : MUX2_X1 port map( A => n19382, B => n19381, S => n19092, Z => 
                           n19096);
   U20872 : OAI21_X1 port map( B1 => n19382, B2 => n19094, A => n19093, ZN => 
                           n19095);
   U20874 : AOI22_X1 port map( A1 => n19363, A2 => n19376, B1 => n19098, B2 => 
                           n19097, ZN => n19102);
   U20875 : NAND2_X1 port map( A1 => n19100, A2 => n25243, ZN => n19101);
   U20876 : NAND3_X1 port map( A1 => n19103, A2 => n18816, A3 => n19359, ZN => 
                           n19104);
   U20877 : NOR2_X1 port map( A1 => n19386, A2 => n25052, ZN => n19110);
   U20878 : AOI22_X1 port map( A1 => n20276, A2 => n19924, B1 => n20517, B2 => 
                           n20272, ZN => n19117);
   U20879 : OAI21_X1 port map( B1 => n19235, B2 => n19237, A => n19112, ZN => 
                           n19116);
   U20880 : OAI21_X1 port map( B1 => n19233, B2 => n19608, A => n19113, ZN => 
                           n19115);
   U20881 : INV_X1 port map( A => n19233, ZN => n19606);
   U20882 : NOR2_X1 port map( A1 => n18863, A2 => n19606, ZN => n19114);
   U20883 : NAND2_X1 port map( A1 => n20276, A2 => n20272, ZN => n19118);
   U20884 : XNOR2_X1 port map( A => n21587, B => n20826, ZN => n21448);
   U20885 : OAI21_X1 port map( B1 => n25388, B2 => n339, A => n19917, ZN => 
                           n19119);
   U20886 : AOI21_X2 port map( B1 => n19120, B2 => n19119, A => n19916, ZN => 
                           n21686);
   U20887 : XNOR2_X1 port map( A => n21686, B => n1528, ZN => n19124);
   U20888 : INV_X1 port map( A => n20062, ZN => n20472);
   U20889 : NAND2_X1 port map( A1 => n20060, A2 => n20055, ZN => n19122);
   U20890 : MUX2_X1 port map( A => n20472, B => n19122, S => n20054, Z => 
                           n19123);
   U20891 : AOI21_X1 port map( B1 => n19523, B2 => n19519, A => n19520, ZN => 
                           n19127);
   U20892 : NOR2_X1 port map( A1 => n19133, A2 => n25364, ZN => n19129);
   U20893 : OAI21_X1 port map( B1 => n19130, B2 => n19129, A => n24324, ZN => 
                           n19137);
   U20894 : NAND3_X1 port map( A1 => n19133, A2 => n19132, A3 => n25364, ZN => 
                           n19134);
   U20895 : AND2_X1 port map( A1 => n19135, A2 => n19134, ZN => n19136);
   U20896 : AOI21_X1 port map( B1 => n19743, B2 => n25421, A => n20410, ZN => 
                           n19154);
   U20897 : NAND2_X1 port map( A1 => n19290, A2 => n19138, ZN => n19139);
   U20898 : MUX2_X1 port map( A => n19562, B => n19139, S => n4262, Z => n19144
                           );
   U20899 : NOR2_X1 port map( A1 => n19290, A2 => n24421, ZN => n19142);
   U20900 : AOI22_X1 port map( A1 => n19142, A2 => n19141, B1 => n19140, B2 => 
                           n3284, ZN => n19143);
   U20901 : NOR3_X1 port map( A1 => n4172, A2 => n19537, A3 => n19531, ZN => 
                           n20257);
   U20902 : NAND2_X1 port map( A1 => n20255, A2 => n25421, ZN => n19911);
   U20903 : INV_X1 port map( A => n19911, ZN => n19152);
   U20905 : AOI21_X2 port map( B1 => n19150, B2 => n19149, A => n19148, ZN => 
                           n20262);
   U20906 : NOR2_X1 port map( A1 => n20262, A2 => n20411, ZN => n19151);
   U20907 : OAI21_X1 port map( B1 => n19152, B2 => n19151, A => n2024, ZN => 
                           n19153);
   U20908 : OAI21_X1 port map( B1 => n19154, B2 => n20263, A => n19153, ZN => 
                           n21228);
   U20910 : INV_X1 port map( A => n19697, ZN => n20103);
   U20911 : INV_X1 port map( A => n19896, ZN => n20104);
   U20912 : XNOR2_X1 port map( A => n21228, B => n21266, ZN => n19159);
   U20913 : NAND2_X1 port map( A1 => n19849, A2 => n19851, ZN => n20072);
   U20914 : NAND2_X1 port map( A1 => n19658, A2 => n19852, ZN => n19157);
   U20915 : MUX2_X1 port map( A => n20072, B => n19157, S => n19850, Z => 
                           n19158);
   U20916 : XNOR2_X1 port map( A => n19159, B => n21689, ZN => n19160);
   U20917 : NOR2_X1 port map( A1 => n18998, A2 => n19417, ZN => n19423);
   U20918 : NAND2_X1 port map( A1 => n19172, A2 => n19407, ZN => n19175);
   U20920 : NOR2_X1 port map( A1 => n19428, A2 => n19760, ZN => n19178);
   U20921 : AOI22_X1 port map( A1 => n19180, A2 => n19179, B1 => n19178, B2 => 
                           n25195, ZN => n19181);
   U20923 : INV_X1 port map( A => n19185, ZN => n19547);
   U20924 : NOR2_X1 port map( A1 => n25057, A2 => n19547, ZN => n19188);
   U20925 : NAND2_X1 port map( A1 => n19402, A2 => n19186, ZN => n19187);
   U20926 : OAI211_X1 port map( C1 => n25223, C2 => n20216, A => n25347, B => 
                           n20510, ZN => n19190);
   U20927 : NOR3_X1 port map( A1 => n25224, A2 => n20510, A3 => n20199, ZN => 
                           n19193);
   U20928 : NOR2_X1 port map( A1 => n19194, A2 => n19660, ZN => n19197);
   U20930 : OAI21_X1 port map( B1 => n19195, B2 => n19660, A => n19659, ZN => 
                           n19196);
   U20931 : XNOR2_X1 port map( A => n20780, B => n21514, ZN => n21645);
   U20932 : NAND2_X1 port map( A1 => n19584, A2 => n19198, ZN => n19200);
   U20933 : MUX2_X1 port map( A => n19200, B => n19586, S => n24481, Z => 
                           n19201);
   U20934 : OAI21_X1 port map( B1 => n19345, B2 => n19346, A => n2333, ZN => 
                           n19207);
   U20935 : NAND2_X1 port map( A1 => n19208, A2 => n5454, ZN => n19209);
   U20936 : AOI21_X1 port map( B1 => n19211, B2 => n19359, A => n19361, ZN => 
                           n19214);
   U20937 : NAND2_X1 port map( A1 => n24940, A2 => n19841, ZN => n19227);
   U20938 : NOR2_X1 port map( A1 => n19219, A2 => n19367, ZN => n19220);
   U20939 : AND2_X1 port map( A1 => n19221, A2 => n19220, ZN => n19223);
   U20940 : OAI211_X2 port map( C1 => n20583, C2 => n20433, A => n19227, B => 
                           n19226, ZN => n21728);
   U20941 : NOR2_X1 port map( A1 => n20183, A2 => n25212, ZN => n19231);
   U20943 : INV_X1 port map( A => n20182, ZN => n20041);
   U20944 : NAND2_X1 port map( A1 => n19228, A2 => n20041, ZN => n19229);
   U20945 : OAI211_X1 port map( C1 => n19231, C2 => n19662, A => n19230, B => 
                           n19229, ZN => n21515);
   U20946 : XNOR2_X1 port map( A => n21728, B => n21515, ZN => n20842);
   U20947 : INV_X1 port map( A => n20842, ZN => n19232);
   U20948 : XNOR2_X1 port map( A => n19232, B => n21645, ZN => n19342);
   U20949 : OAI21_X1 port map( B1 => n19233, B2 => n19607, A => n19608, ZN => 
                           n19234);
   U20950 : NOR2_X1 port map( A1 => n19241, A2 => n25012, ZN => n19242);
   U20951 : NOR2_X1 port map( A1 => n19243, A2 => n19242, ZN => n19244);
   U20952 : NAND3_X1 port map( A1 => n3986, A2 => n25260, A3 => n361, ZN => 
                           n19247);
   U20953 : INV_X1 port map( A => n19576, ZN => n19249);
   U20954 : MUX2_X1 port map( A => n19592, B => n2346, S => n19250, Z => n19253
                           );
   U20955 : NAND2_X1 port map( A1 => n25476, A2 => n20428, ZN => n19259);
   U20956 : NOR2_X1 port map( A1 => n19255, A2 => n19598, ZN => n19256);
   U20957 : AOI22_X1 port map( A1 => n19257, A2 => n24079, B1 => n19597, B2 => 
                           n19256, ZN => n19258);
   U20959 : NOR2_X1 port map( A1 => n19264, A2 => n19261, ZN => n19262);
   U20960 : NOR2_X1 port map( A1 => n19263, A2 => n19262, ZN => n19268);
   U20961 : NAND2_X1 port map( A1 => n19265, A2 => n19264, ZN => n19267);
   U20962 : NAND3_X1 port map( A1 => n19531, A2 => n19530, A3 => n19270, ZN => 
                           n19271);
   U20963 : INV_X1 port map( A => n19565, ZN => n19569);
   U20964 : NAND2_X1 port map( A1 => n20400, A2 => n20414, ZN => n19293);
   U20965 : NOR2_X1 port map( A1 => n19278, A2 => n19277, ZN => n19541);
   U20966 : NAND2_X1 port map( A1 => n20417, A2 => n20415, ZN => n19288);
   U20967 : INV_X1 port map( A => n19523, ZN => n19279);
   U20968 : OAI21_X1 port map( B1 => n19282, B2 => n19281, A => n19521, ZN => 
                           n19287);
   U20969 : NAND3_X1 port map( A1 => n19283, A2 => n19518, A3 => n18895, ZN => 
                           n19286);
   U20970 : NAND3_X1 port map( A1 => n19526, A2 => n19284, A3 => n19520, ZN => 
                           n19285);
   U20971 : MUX2_X1 port map( A => n3284, B => n19560, S => n19556, Z => n19289
                           );
   U20973 : MUX2_X1 port map( A => n24457, B => n18927, S => n19296, Z => 
                           n19299);
   U20974 : NOR2_X1 port map( A1 => n19300, A2 => n19296, ZN => n19298);
   U20975 : AOI21_X1 port map( B1 => n19304, B2 => n19303, A => n24441, ZN => 
                           n19305);
   U20976 : NAND3_X1 port map( A1 => n19313, A2 => n264, A3 => n19312, ZN => 
                           n19314);
   U20977 : NAND2_X1 port map( A1 => n19315, A2 => n5371, ZN => n19316);
   U20978 : NAND3_X1 port map( A1 => n19318, A2 => n19317, A3 => n19316, ZN => 
                           n19319);
   U20979 : NAND2_X1 port map( A1 => n19320, A2 => n19319, ZN => n20241);
   U20981 : INV_X1 port map( A => n19936, ZN => n20244);
   U20982 : NOR2_X1 port map( A1 => n19329, A2 => n19328, ZN => n19330);
   U20983 : INV_X1 port map( A => n19937, ZN => n20243);
   U20984 : INV_X1 port map( A => n19499, ZN => n19496);
   U20985 : OAI21_X1 port map( B1 => n19500, B2 => n357, A => n19501, ZN => 
                           n19337);
   U20986 : NOR2_X1 port map( A1 => n19502, A2 => n19497, ZN => n19336);
   U20988 : NAND3_X1 port map( A1 => n19936, A2 => n20242, A3 => n19939, ZN => 
                           n19339);
   U20989 : XNOR2_X1 port map( A => n21106, B => n2735, ZN => n19340);
   U20990 : XNOR2_X1 port map( A => n21121, B => n19340, ZN => n19341);
   U20991 : NAND2_X1 port map( A1 => n25474, A2 => n19346, ZN => n20389);
   U20992 : NAND2_X1 port map( A1 => n20389, A2 => n20388, ZN => n19347);
   U20993 : OAI21_X1 port map( B1 => n19348, B2 => n20388, A => n19347, ZN => 
                           n19350);
   U20994 : NAND2_X1 port map( A1 => n19349, A2 => n352, ZN => n20390);
   U20997 : NAND2_X1 port map( A1 => n19357, A2 => n19353, ZN => n19448);
   U20998 : INV_X1 port map( A => n19448, ZN => n19354);
   U20999 : NAND2_X1 port map( A1 => n19354, A2 => n19452, ZN => n19355);
   U21002 : NOR2_X1 port map( A1 => n19364, A2 => n2216, ZN => n19369);
   U21003 : NOR2_X1 port map( A1 => n19366, A2 => n24968, ZN => n19368);
   U21004 : AOI22_X1 port map( A1 => n19376, A2 => n19369, B1 => n19368, B2 => 
                           n19367, ZN => n19374);
   U21005 : NOR2_X1 port map( A1 => n19371, A2 => n24361, ZN => n19372);
   U21006 : AND3_X1 port map( A1 => n19382, A2 => n19381, A3 => n19380, ZN => 
                           n19383);
   U21007 : NAND2_X1 port map( A1 => n19384, A2 => n19389, ZN => n19385);
   U21008 : XNOR2_X1 port map( A => n1326, B => n19392, ZN => n19443);
   U21009 : NOR2_X1 port map( A1 => n19396, A2 => n24407, ZN => n19398);
   U21010 : OAI21_X1 port map( B1 => n19402, B2 => n1711, A => n19719, ZN => 
                           n19405);
   U21011 : NAND2_X1 port map( A1 => n19406, A2 => n19412, ZN => n19410);
   U21012 : MUX2_X1 port map( A => n19410, B => n19409, S => n19408, Z => 
                           n19416);
   U21013 : NOR2_X1 port map( A1 => n19412, A2 => n19411, ZN => n19414);
   U21014 : OAI21_X1 port map( B1 => n24584, B2 => n19418, A => n19417, ZN => 
                           n19422);
   U21015 : INV_X1 port map( A => n19761, ZN => n19431);
   U21016 : AOI21_X1 port map( B1 => n19428, B2 => n19760, A => n19427, ZN => 
                           n19429);
   U21017 : OAI21_X1 port map( B1 => n24758, B2 => n19760, A => n19429, ZN => 
                           n19430);
   U21018 : NAND2_X1 port map( A1 => n19431, A2 => n19430, ZN => n19432);
   U21019 : MUX2_X1 port map( A => n20174, B => n20586, S => n19432, Z => 
                           n19442);
   U21020 : OAI21_X1 port map( B1 => n19435, B2 => n25423, A => n19433, ZN => 
                           n19440);
   U21021 : XNOR2_X1 port map( A => n19443, B => n21505, ZN => n19514);
   U21029 : NAND2_X1 port map( A1 => n19459, A2 => n19464, ZN => n19461);
   U21030 : MUX2_X1 port map( A => n19462, B => n19461, S => n19460, Z => 
                           n19463);
   U21032 : NAND2_X1 port map( A1 => n19468, A2 => n19471, ZN => n19475);
   U21033 : OAI21_X1 port map( B1 => n17872, B2 => n19470, A => n19469, ZN => 
                           n19473);
   U21034 : NAND2_X1 port map( A1 => n19473, A2 => n19472, ZN => n19474);
   U21035 : AND2_X2 port map( A1 => n19475, A2 => n19474, ZN => n20173);
   U21036 : MUX2_X1 port map( A => n20169, B => n20235, S => n20173, Z => 
                           n19484);
   U21039 : NOR2_X1 port map( A1 => n19484, A2 => n20168, ZN => n19509);
   U21040 : OAI21_X1 port map( B1 => n19490, B2 => n240, A => n20388, ZN => 
                           n19486);
   U21042 : NAND3_X1 port map( A1 => n19490, A2 => n19345, A3 => n19488, ZN => 
                           n19491);
   U21043 : OAI211_X1 port map( C1 => n19500, C2 => n19497, A => n19496, B => 
                           n19495, ZN => n19506);
   U21044 : NAND3_X1 port map( A1 => n19500, A2 => n19499, A3 => n25459, ZN => 
                           n19505);
   U21045 : NOR2_X1 port map( A1 => n19502, A2 => n19501, ZN => n19503);
   U21046 : NOR2_X1 port map( A1 => n19494, A2 => n19777, ZN => n19507);
   U21049 : INV_X1 port map( A => n19939, ZN => n19788);
   U21050 : INV_X1 port map( A => n20242, ZN => n19513);
   U21051 : OAI21_X1 port map( B1 => n19939, B2 => n19936, A => n19937, ZN => 
                           n19511);
   U21052 : OAI21_X1 port map( B1 => n19819, B2 => n19513, A => n19512, ZN => 
                           n21616);
   U21053 : XNOR2_X1 port map( A => n21659, B => n21616, ZN => n20285);
   U21054 : XNOR2_X1 port map( A => n20285, B => n19514, ZN => n19624);
   U21055 : OR2_X1 port map( A1 => n21068, A2 => n19986, ZN => n19988);
   U21056 : MUX2_X1 port map( A => n19987, B => n19785, S => n19986, Z => 
                           n19516);
   U21057 : INV_X1 port map( A => n19983, ZN => n19751);
   U21058 : NAND2_X1 port map( A1 => n19986, A2 => n19751, ZN => n19515);
   U21059 : INV_X1 port map( A => n19520, ZN => n19521);
   U21062 : AOI22_X1 port map( A1 => n19532, A2 => n19531, B1 => n19530, B2 => 
                           n19529, ZN => n19538);
   U21063 : AOI21_X1 port map( B1 => n19535, B2 => n5480, A => n19533, ZN => 
                           n19536);
   U21064 : INV_X1 port map( A => n24454, ZN => n19962);
   U21065 : MUX2_X1 port map( A => n19540, B => n3773, S => n19539, Z => n19545
                           );
   U21067 : AOI21_X1 port map( B1 => n25057, B2 => n19547, A => n19546, ZN => 
                           n19553);
   U21069 : OAI21_X1 port map( B1 => n19553, B2 => n19552, A => n19551, ZN => 
                           n20373);
   U21070 : MUX2_X1 port map( A => n19962, B => n20368, S => n20369, Z => 
                           n19574);
   U21071 : NAND2_X1 port map( A1 => n19554, A2 => n4262, ZN => n19564);
   U21072 : INV_X1 port map( A => n19555, ZN => n19557);
   U21073 : NOR2_X1 port map( A1 => n19557, A2 => n24421, ZN => n19563);
   U21074 : NAND3_X1 port map( A1 => n19560, A2 => n19559, A3 => n19558, ZN => 
                           n19561);
   U21075 : NOR2_X1 port map( A1 => n20370, A2 => n24558, ZN => n19573);
   U21076 : NOR2_X1 port map( A1 => n19569, A2 => n1053, ZN => n19571);
   U21077 : NOR2_X1 port map( A1 => n20368, A2 => n3428, ZN => n19572);
   U21078 : INV_X1 port map( A => n20961, ZN => n20450);
   U21079 : AOI21_X1 port map( B1 => n19581, B2 => n19580, A => n19198, ZN => 
                           n19583);
   U21080 : MUX2_X1 port map( A => n19584, B => n19583, S => n19582, Z => 
                           n19585);
   U21081 : INV_X1 port map( A => n20451, ZN => n19942);
   U21082 : NAND3_X1 port map( A1 => n19587, A2 => n24483, A3 => n19591, ZN => 
                           n19588);
   U21083 : NOR2_X1 port map( A1 => n25001, A2 => n24079, ZN => n19600);
   U21084 : NOR2_X1 port map( A1 => n19597, A2 => n19596, ZN => n19599);
   U21085 : NAND2_X1 port map( A1 => n20960, A2 => n19942, ZN => n19605);
   U21086 : OAI211_X1 port map( C1 => n20450, C2 => n19942, A => n20377, B => 
                           n19605, ZN => n19621);
   U21087 : NOR2_X1 port map( A1 => n19608, A2 => n2644, ZN => n19609);
   U21088 : INV_X1 port map( A => n19612, ZN => n19619);
   U21089 : NOR2_X1 port map( A1 => n19613, A2 => n19615, ZN => n19618);
   U21090 : OAI21_X1 port map( B1 => n19616, B2 => n19615, A => n19614, ZN => 
                           n19617);
   U21091 : NOR2_X1 port map( A1 => n20377, A2 => n20448, ZN => n19620);
   U21092 : AOI22_X1 port map( A1 => n20158, A2 => n20960, B1 => n19620, B2 => 
                           n20451, ZN => n20962);
   U21093 : NAND2_X1 port map( A1 => n19621, A2 => n20962, ZN => n19622);
   U21094 : XNOR2_X1 port map( A => n24305, B => n19622, ZN => n20723);
   U21095 : XNOR2_X1 port map( A => n24898, B => n20723, ZN => n19623);
   U21098 : INV_X1 port map( A => n19629, ZN => n19632);
   U21099 : OAI21_X1 port map( B1 => n19632, B2 => n19631, A => n19630, ZN => 
                           n19633);
   U21100 : INV_X1 port map( A => n19636, ZN => n19634);
   U21101 : MUX2_X1 port map( A => n19634, B => n20484, S => n20359, Z => 
                           n19639);
   U21104 : NAND2_X1 port map( A1 => n20482, A2 => n19636, ZN => n19637);
   U21106 : NOR2_X1 port map( A1 => n25088, A2 => n19928, ZN => n19640);
   U21111 : INV_X1 port map( A => n20343, ZN => n19645);
   U21113 : NOR2_X1 port map( A1 => n20281, A2 => n1733, ZN => n19646);
   U21114 : NAND3_X1 port map( A1 => n20345, A2 => n20281, A3 => n20279, ZN => 
                           n19647);
   U21115 : NAND4_X2 port map( A1 => n19650, A2 => n19649, A3 => n19648, A4 => 
                           n19647, ZN => n21193);
   U21116 : XNOR2_X1 port map( A => n21193, B => n25265, ZN => n21715);
   U21117 : XNOR2_X1 port map( A => n21715, B => n20831, ZN => n19667);
   U21118 : NOR2_X1 port map( A1 => n24567, A2 => n20338, ZN => n19653);
   U21119 : NOR2_X1 port map( A1 => n20669, A2 => n20668, ZN => n19652);
   U21120 : MUX2_X1 port map( A => n19653, B => n19652, S => n20666, Z => 
                           n19656);
   U21121 : NOR2_X1 port map( A1 => n20669, A2 => n20336, ZN => n20349);
   U21122 : AND2_X1 port map( A1 => n20666, A2 => n20336, ZN => n19654);
   U21125 : XNOR2_X1 port map( A => n21306, B => n24916, ZN => n19665);
   U21126 : INV_X1 port map( A => n20183, ZN => n20186);
   U21127 : INV_X1 port map( A => n20181, ZN => n20038);
   U21128 : NAND3_X1 port map( A1 => n20191, A2 => n20041, A3 => n20038, ZN => 
                           n19663);
   U21129 : XNOR2_X1 port map( A => n21311, B => n869, ZN => n19664);
   U21130 : XNOR2_X1 port map( A => n19665, B => n19664, ZN => n19666);
   U21131 : XNOR2_X1 port map( A => n19667, B => n19666, ZN => n22688);
   U21135 : INV_X1 port map( A => n19675, ZN => n19677);
   U21136 : OAI211_X1 port map( C1 => n19675, C2 => n20124, A => n20130, B => 
                           n19674, ZN => n19676);
   U21137 : XNOR2_X1 port map( A => n21649, B => n21436, ZN => n21253);
   U21138 : INV_X1 port map( A => n19991, ZN => n20135);
   U21139 : OAI211_X1 port map( C1 => n20135, C2 => n20014, A => n1954, B => 
                           n20019, ZN => n19678);
   U21140 : XNOR2_X1 port map( A => n21336, B => n2058, ZN => n19679);
   U21141 : XNOR2_X1 port map( A => n21253, B => n19679, ZN => n19696);
   U21142 : INV_X1 port map( A => n20301, ZN => n20008);
   U21143 : NAND2_X1 port map( A1 => n20008, A2 => n19976, ZN => n19682);
   U21144 : INV_X1 port map( A => n19680, ZN => n19681);
   U21145 : INV_X1 port map( A => n19785, ZN => n19980);
   U21146 : OAI211_X1 port map( C1 => n19784, C2 => n19986, A => n19984, B => 
                           n19785, ZN => n19683);
   U21147 : OAI21_X1 port map( B1 => n19986, B2 => n19750, A => n19683, ZN => 
                           n19685);
   U21148 : NOR2_X1 port map( A1 => n19684, A2 => n19987, ZN => n21066);
   U21150 : XNOR2_X1 port map( A => n21332, B => n21997, ZN => n19694);
   U21151 : NAND2_X1 port map( A1 => n20539, A2 => n20147, ZN => n19690);
   U21153 : INV_X1 port map( A => n20145, ZN => n19686);
   U21154 : NAND2_X1 port map( A1 => n20145, A2 => n20149, ZN => n20534);
   U21155 : NAND2_X1 port map( A1 => n19691, A2 => n19714, ZN => n19693);
   U21156 : XNOR2_X1 port map( A => n21729, B => n21582, ZN => n21200);
   U21157 : XNOR2_X1 port map( A => n19694, B => n21200, ZN => n19695);
   U21158 : XNOR2_X1 port map( A => n19696, B => n19695, ZN => n22685);
   U21159 : OR2_X1 port map( A1 => n22688, A2 => n22685, ZN => n22352);
   U21160 : MUX2_X1 port map( A => n19896, B => n21033, S => n19155, Z => 
                           n19699);
   U21162 : NOR2_X1 port map( A1 => n19700, A2 => n19880, ZN => n19702);
   U21163 : MUX2_X1 port map( A => n3480, B => n20554, S => n20328, Z => n19701
                           );
   U21164 : MUX2_X2 port map( A => n19702, B => n19701, S => n20555, Z => 
                           n21258);
   U21165 : XNOR2_X1 port map( A => n21300, B => n21258, ZN => n19713);
   U21166 : MUX2_X1 port map( A => n20616, B => n20571, S => n20618, Z => 
                           n19706);
   U21167 : NAND3_X1 port map( A1 => n19704, A2 => n20614, A3 => n19703, ZN => 
                           n19705);
   U21168 : INV_X1 port map( A => n20669, ZN => n20337);
   U21169 : NAND2_X1 port map( A1 => n20337, A2 => n20668, ZN => n19707);
   U21170 : OAI22_X1 port map( A1 => n19710, A2 => n19709, B1 => n20337, B2 => 
                           n20670, ZN => n19711);
   U21171 : XNOR2_X1 port map( A => n21745, B => n21975, ZN => n21208);
   U21172 : XNOR2_X1 port map( A => n21208, B => n19713, ZN => n19738);
   U21173 : INV_X1 port map( A => n21506, ZN => n21979);
   U21174 : INV_X1 port map( A => n20111, ZN => n20118);
   U21177 : XNOR2_X1 port map( A => n21297, B => n21979, ZN => n19736);
   U21178 : INV_X1 port map( A => n19719, ZN => n19722);
   U21179 : INV_X1 port map( A => n19725, ZN => n19721);
   U21180 : AOI21_X1 port map( B1 => n19722, B2 => n19721, A => n19720, ZN => 
                           n19724);
   U21181 : OAI211_X1 port map( C1 => n19726, C2 => n19725, A => n19724, B => 
                           n19723, ZN => n19728);
   U21182 : INV_X1 port map( A => n19729, ZN => n19733);
   U21183 : INV_X1 port map( A => n19730, ZN => n19731);
   U21184 : NAND2_X1 port map( A1 => n19733, A2 => n19732, ZN => n19734);
   U21185 : XNOR2_X1 port map( A => n24491, B => n2033, ZN => n19735);
   U21186 : XNOR2_X1 port map( A => n19736, B => n19735, ZN => n19737);
   U21187 : INV_X1 port map( A => n21848, ZN => n21289);
   U21188 : NAND2_X1 port map( A1 => n22352, A2 => n21289, ZN => n19836);
   U21189 : INV_X1 port map( A => n20419, ZN => n20204);
   U21190 : NAND3_X1 port map( A1 => n20422, A2 => n20400, A3 => n5590, ZN => 
                           n19739);
   U21192 : INV_X1 port map( A => n20426, ZN => n20598);
   U21193 : NAND2_X1 port map( A1 => n20427, A2 => n20598, ZN => n19846);
   U21194 : INV_X1 port map( A => n25442, ZN => n19749);
   U21195 : OAI21_X1 port map( B1 => n20263, B2 => n20262, A => n20410, ZN => 
                           n19742);
   U21196 : NOR2_X1 port map( A1 => n20193, A2 => n20192, ZN => n19745);
   U21197 : NAND2_X1 port map( A1 => n20437, A2 => n19745, ZN => n19747);
   U21198 : NOR2_X1 port map( A1 => n20193, A2 => n20576, ZN => n20195);
   U21199 : NAND2_X1 port map( A1 => n20195, A2 => n24940, ZN => n19746);
   U21200 : XNOR2_X1 port map( A => n19749, B => n19748, ZN => n19769);
   U21201 : INV_X1 port map( A => n19750, ZN => n21065);
   U21202 : NAND2_X1 port map( A1 => n21065, A2 => n25579, ZN => n19754);
   U21203 : OAI21_X1 port map( B1 => n19984, B2 => n19785, A => n19751, ZN => 
                           n19752);
   U21205 : NAND3_X1 port map( A1 => n19754, A2 => n19753, A3 => n21067, ZN => 
                           n21132);
   U21206 : NOR2_X1 port map( A1 => n25242, A2 => n20134, ZN => n19759);
   U21207 : XNOR2_X1 port map( A => n21132, B => n21245, ZN => n21328);
   U21210 : INV_X1 port map( A => n20593, ZN => n20176);
   U21211 : OAI21_X1 port map( B1 => n20590, B2 => n20586, A => n20176, ZN => 
                           n19764);
   U21212 : NAND3_X1 port map( A1 => n20589, A2 => n20176, A3 => n3734, ZN => 
                           n19765);
   U21213 : OAI211_X2 port map( C1 => n19952, C2 => n20591, A => n19766, B => 
                           n19765, ZN => n21720);
   U21214 : XNOR2_X1 port map( A => n21720, B => n450, ZN => n19767);
   U21215 : XNOR2_X1 port map( A => n21328, B => n19767, ZN => n19768);
   U21217 : AND2_X1 port map( A1 => n22685, A2 => n21816, ZN => n22349);
   U21218 : INV_X1 port map( A => n22688, ZN => n22686);
   U21219 : NAND3_X1 port map( A1 => n2688, A2 => n20448, A3 => n20377, ZN => 
                           n19773);
   U21221 : XNOR2_X1 port map( A => n21750, B => n21608, ZN => n20708);
   U21222 : AND2_X1 port map( A1 => n24461, A2 => n20384, ZN => n20385);
   U21224 : NAND2_X1 port map( A1 => n20459, A2 => n20384, ZN => n19776);
   U21225 : NAND3_X1 port map( A1 => n20234, A2 => n20231, A3 => n25205, ZN => 
                           n19780);
   U21226 : OAI21_X1 port map( B1 => n20169, B2 => n20236, A => n20168, ZN => 
                           n19779);
   U21227 : NOR2_X1 port map( A1 => n20173, A2 => n20236, ZN => n19778);
   U21228 : AOI22_X1 port map( A1 => n19780, A2 => n19779, B1 => n20235, B2 => 
                           n19778, ZN => n21042);
   U21229 : XNOR2_X1 port map( A => n21267, B => n21042, ZN => n21345);
   U21230 : XNOR2_X1 port map( A => n20708, B => n21345, ZN => n19796);
   U21231 : OAI21_X1 port map( B1 => n20589, B2 => n20590, A => n20586, ZN => 
                           n19782);
   U21232 : NOR2_X1 port map( A1 => n20587, A2 => n20588, ZN => n19781);
   U21233 : AOI22_X2 port map( A1 => n19783, A2 => n19782, B1 => n20174, B2 => 
                           n19781, ZN => n21227);
   U21234 : INV_X1 port map( A => n21227, ZN => n21588);
   U21235 : OAI21_X1 port map( B1 => n19785, B2 => n19784, A => n19984, ZN => 
                           n19787);
   U21236 : XNOR2_X1 port map( A => n21588, B => n21231, ZN => n19794);
   U21238 : NAND2_X1 port map( A1 => n19788, A2 => n1344, ZN => n19791);
   U21240 : OAI211_X1 port map( C1 => n20243, C2 => n20248, A => n19789, B => 
                           n19821, ZN => n19790);
   U21241 : XNOR2_X1 port map( A => n21141, B => n2042, ZN => n19793);
   U21242 : XNOR2_X1 port map( A => n19794, B => n19793, ZN => n19795);
   U21243 : INV_X1 port map( A => n22689, ZN => n21817);
   U21244 : NAND3_X1 port map( A1 => n22686, A2 => n21816, A3 => n21817, ZN => 
                           n19835);
   U21245 : AND2_X1 port map( A1 => n3519, A2 => n19924, ZN => n19798);
   U21247 : NAND2_X1 port map( A1 => n20169, A2 => n20231, ZN => n19802);
   U21248 : AOI21_X1 port map( B1 => n19803, B2 => n19802, A => n20239, ZN => 
                           n19808);
   U21249 : NAND2_X1 port map( A1 => n20173, A2 => n20236, ZN => n19806);
   U21250 : INV_X1 port map( A => n20231, ZN => n19804);
   U21254 : NAND2_X1 port map( A1 => n19809, A2 => n20281, ZN => n19812);
   U21255 : MUX2_X1 port map( A => n20281, B => n20343, S => n20345, Z => 
                           n19810);
   U21256 : MUX2_X1 port map( A => n19810, B => n1484, S => n20279, Z => n19811
                           );
   U21257 : OAI21_X1 port map( B1 => n19645, B2 => n19812, A => n19811, ZN => 
                           n21971);
   U21258 : INV_X1 port map( A => n21971, ZN => n19813);
   U21259 : XNOR2_X1 port map( A => n21430, B => n19813, ZN => n19833);
   U21260 : NOR2_X1 port map( A1 => n20507, A2 => n20214, ZN => n20218);
   U21262 : NOR2_X1 port map( A1 => n25224, A2 => n100, ZN => n19814);
   U21264 : OAI21_X2 port map( B1 => n19816, B2 => n20199, A => n19815, ZN => 
                           n21735);
   U21265 : INV_X1 port map( A => n19817, ZN => n19820);
   U21266 : OAI211_X1 port map( C1 => n20244, C2 => n20242, A => n24077, B => 
                           n19821, ZN => n19822);
   U21267 : XNOR2_X1 port map( A => n21319, B => n2228, ZN => n19823);
   U21268 : XNOR2_X1 port map( A => n19823, B => n21735, ZN => n19831);
   U21269 : INV_X1 port map( A => n20268, ZN => n20496);
   U21270 : NAND2_X1 port map( A1 => n20501, A2 => n20496, ZN => n19827);
   U21272 : NAND3_X1 port map( A1 => n20411, A2 => n25420, A3 => n20410, ZN => 
                           n19829);
   U21273 : XNOR2_X1 port map( A => n21561, B => n21738, ZN => n21224);
   U21274 : INV_X1 port map( A => n21224, ZN => n19830);
   U21275 : XNOR2_X1 port map( A => n19830, B => n19831, ZN => n19832);
   U21276 : NOR2_X1 port map( A1 => n21847, A2 => n21816, ZN => n22690);
   U21277 : NAND2_X1 port map( A1 => n22690, A2 => n21848, ZN => n19834);
   U21278 : OAI211_X2 port map( C1 => n19836, C2 => n22349, A => n19835, B => 
                           n19834, ZN => n23865);
   U21281 : NOR2_X1 port map( A1 => n5208, A2 => n20576, ZN => n19838);
   U21282 : NAND3_X1 port map( A1 => n19843, A2 => n19842, A3 => n19841, ZN => 
                           n19844);
   U21283 : XNOR2_X1 port map( A => n20804, B => n21974, ZN => n20722);
   U21284 : NOR2_X1 port map( A1 => n20597, A2 => n20427, ZN => n20602);
   U21285 : INV_X1 port map( A => n20427, ZN => n20595);
   U21286 : NAND2_X1 port map( A1 => n20595, A2 => n20599, ZN => n19845);
   U21287 : NAND2_X1 port map( A1 => n19846, A2 => n19845, ZN => n19847);
   U21288 : XNOR2_X1 port map( A => n21660, B => n21616, ZN => n21003);
   U21289 : XNOR2_X1 port map( A => n21003, B => n20722, ZN => n19870);
   U21290 : INV_X1 port map( A => n20071, ZN => n20074);
   U21292 : NOR2_X1 port map( A1 => n20415, A2 => n20400, ZN => n20416);
   U21293 : NOR2_X1 port map( A1 => n20416, A2 => n20414, ZN => n19861);
   U21294 : INV_X1 port map( A => n20415, ZN => n20399);
   U21295 : NOR2_X1 port map( A1 => n20399, A2 => n20414, ZN => n19856);
   U21296 : NAND2_X1 port map( A1 => n19856, A2 => n1662, ZN => n19859);
   U21297 : NAND2_X1 port map( A1 => n19857, A2 => n4509, ZN => n19858);
   U21299 : XNOR2_X1 port map( A => n21301, B => n21136, ZN => n19868);
   U21300 : NAND2_X1 port map( A1 => n25212, A2 => n20039, ZN => n19863);
   U21301 : NAND2_X1 port map( A1 => n25212, A2 => n25478, ZN => n20043);
   U21302 : MUX2_X1 port map( A => n19863, B => n20043, S => n20191, Z => 
                           n19864);
   U21304 : XNOR2_X1 port map( A => n20964, B => n2044, ZN => n19867);
   U21305 : XNOR2_X1 port map( A => n19868, B => n19867, ZN => n19869);
   U21307 : OAI21_X1 port map( B1 => n20572, B2 => n3795, A => n20571, ZN => 
                           n19874);
   U21308 : NAND2_X2 port map( A1 => n19874, A2 => n19873, ZN => n21399);
   U21309 : AOI21_X1 port map( B1 => n20023, B2 => n20562, A => n20094, ZN => 
                           n19877);
   U21311 : XNOR2_X1 port map( A => n25040, B => n21399, ZN => n20816);
   U21312 : NAND2_X1 port map( A1 => n20556, A2 => n20557, ZN => n19879);
   U21313 : AND2_X1 port map( A1 => n20091, A2 => n19879, ZN => n19882);
   U21314 : OAI21_X1 port map( B1 => n19880, B2 => n20330, A => n20328, ZN => 
                           n19881);
   U21315 : NAND2_X1 port map( A1 => n19917, A2 => n25262, ZN => n20114);
   U21316 : OAI22_X1 port map( A1 => n25262, A2 => n19883, B1 => n20109, B2 => 
                           n19887, ZN => n19884);
   U21317 : NAND2_X1 port map( A1 => n19884, A2 => n20118, ZN => n19886);
   U21318 : XNOR2_X1 port map( A => n21496, B => n20816, ZN => n19903);
   U21322 : INV_X1 port map( A => n20102, ZN => n19895);
   U21323 : NAND2_X1 port map( A1 => n19895, A2 => n19896, ZN => n19913);
   U21324 : NAND2_X1 port map( A1 => n20101, A2 => n20100, ZN => n19894);
   U21325 : AOI21_X1 port map( B1 => n19913, B2 => n19894, A => n19893, ZN => 
                           n19899);
   U21326 : NAND2_X1 port map( A1 => n19895, A2 => n24378, ZN => n19897);
   U21327 : AOI21_X1 port map( B1 => n19897, B2 => n19896, A => n20100, ZN => 
                           n19898);
   U21328 : XNOR2_X1 port map( A => n20697, B => n21621, ZN => n19901);
   U21329 : XNOR2_X1 port map( A => n21247, B => n2193, ZN => n19900);
   U21330 : XNOR2_X1 port map( A => n19901, B => n19900, ZN => n19902);
   U21331 : XNOR2_X1 port map( A => n19903, B => n19902, ZN => n22227);
   U21332 : INV_X1 port map( A => n22227, ZN => n21791);
   U21333 : INV_X1 port map( A => n20501, ZN => n20226);
   U21334 : NOR2_X1 port map( A1 => n20502, A2 => n20225, ZN => n19907);
   U21335 : NOR2_X1 port map( A1 => n343, A2 => n20497, ZN => n19906);
   U21336 : OAI211_X1 port map( C1 => n19904, C2 => n20269, A => n20226, B => 
                           n24887, ZN => n19905);
   U21337 : OAI21_X1 port map( B1 => n19907, B2 => n19906, A => n19905, ZN => 
                           n21510);
   U21338 : NAND2_X1 port map( A1 => n2024, A2 => n345, ZN => n19909);
   U21339 : NAND2_X1 port map( A1 => n19909, A2 => n19910, ZN => n19912);
   U21340 : XNOR2_X1 port map( A => n21510, B => n20778, ZN => n21108);
   U21341 : MUX2_X1 port map( A => n21033, B => n19913, S => n21038, Z => 
                           n19914);
   U21342 : OAI21_X1 port map( B1 => n19915, B2 => n20099, A => n19914, ZN => 
                           n21331);
   U21343 : OAI21_X1 port map( B1 => n25034, B2 => n20118, A => n25388, ZN => 
                           n19918);
   U21345 : NAND3_X1 port map( A1 => n20117, A2 => n20118, A3 => n25514, ZN => 
                           n19920);
   U21346 : XNOR2_X1 port map( A => n21331, B => n21647, ZN => n20568);
   U21347 : XNOR2_X1 port map( A => n21108, B => n20568, ZN => n19935);
   U21348 : NAND2_X1 port map( A1 => n351, A2 => n20517, ZN => n19923);
   U21349 : NAND2_X1 port map( A1 => n20516, A2 => n19924, ZN => n19922);
   U21350 : NAND2_X1 port map( A1 => n19923, A2 => n19922, ZN => n20222);
   U21351 : INV_X1 port map( A => n19924, ZN => n20514);
   U21352 : NAND2_X1 port map( A1 => n20276, A2 => n20514, ZN => n20519);
   U21353 : OAI21_X1 port map( B1 => n20272, B2 => n20517, A => n19925, ZN => 
                           n19926);
   U21355 : XNOR2_X1 port map( A => n20780, B => n24986, ZN => n19933);
   U21356 : NAND3_X1 port map( A1 => n20468, A2 => n19928, A3 => n25490, ZN => 
                           n19931);
   U21358 : NAND2_X1 port map( A1 => n20470, A2 => n20473, ZN => n19930);
   U21359 : NAND3_X1 port map( A1 => n20062, A2 => n25088, A3 => n20055, ZN => 
                           n19929);
   U21361 : XNOR2_X1 port map( A => n20999, B => n23679, ZN => n19932);
   U21362 : XNOR2_X1 port map( A => n19933, B => n19932, ZN => n19934);
   U21363 : INV_X1 port map( A => n22226, ZN => n21836);
   U21364 : MUX2_X1 port map( A => n20243, B => n19939, S => n19936, Z => 
                           n19941);
   U21365 : NOR2_X1 port map( A1 => n19937, A2 => n20242, ZN => n19938);
   U21366 : XNOR2_X1 port map( A => n25062, B => n663, ZN => n19946);
   U21367 : INV_X1 port map( A => n20448, ZN => n20159);
   U21368 : AOI21_X1 port map( B1 => n19948, B2 => n20383, A => n20460, ZN => 
                           n19947);
   U21369 : NAND2_X1 port map( A1 => n20461, A2 => n1327, ZN => n20163);
   U21370 : NAND2_X1 port map( A1 => n19947, A2 => n20163, ZN => n19950);
   U21371 : NAND3_X1 port map( A1 => n20588, A2 => n20593, A3 => n20586, ZN => 
                           n19954);
   U21373 : NAND2_X1 port map( A1 => n25205, A2 => n20169, ZN => n19956);
   U21374 : MUX2_X1 port map( A => n19956, B => n20234, S => n20235, Z => 
                           n19961);
   U21375 : INV_X1 port map( A => n20169, ZN => n20232);
   U21377 : NAND2_X1 port map( A1 => n20173, A2 => n20231, ZN => n19957);
   U21378 : OAI22_X1 port map( A1 => n20235, A2 => n19958, B1 => n25205, B2 => 
                           n19957, ZN => n19959);
   U21379 : INV_X1 port map( A => n19959, ZN => n19960);
   U21380 : XNOR2_X1 port map( A => n20767, B => n20948, ZN => n19965);
   U21381 : NOR2_X1 port map( A1 => n20374, A2 => n20370, ZN => n19964);
   U21382 : XNOR2_X1 port map( A => n19965, B => n21115, ZN => n21642);
   U21383 : XNOR2_X1 port map( A => n19966, B => n21642, ZN => n20036);
   U21384 : NOR2_X1 port map( A1 => n20312, A2 => n20546, ZN => n19968);
   U21386 : NOR3_X1 port map( A1 => n20126, A2 => n20124, A3 => n20309, ZN => 
                           n19969);
   U21387 : NOR2_X2 port map( A1 => n19970, A2 => n19969, ZN => n21126);
   U21389 : OAI22_X1 port map( A1 => n20289, A2 => n19971, B1 => n20131, B2 => 
                           n21010, ZN => n19974);
   U21390 : XNOR2_X1 port map( A => n21534, B => n21126, ZN => n20812);
   U21391 : NAND2_X1 port map( A1 => n20301, A2 => n19976, ZN => n19977);
   U21392 : OAI21_X1 port map( B1 => n19979, B2 => n20141, A => n19978, ZN => 
                           n21967);
   U21393 : XNOR2_X1 port map( A => n20812, B => n21967, ZN => n21083);
   U21396 : NOR2_X1 port map( A1 => n19988, A2 => n24979, ZN => n19989);
   U21397 : NOR2_X2 port map( A1 => n19990, A2 => n19989, ZN => n21318);
   U21398 : INV_X1 port map( A => n20016, ZN => n19996);
   U21399 : OAI21_X1 port map( B1 => n20134, B2 => n20019, A => n25242, ZN => 
                           n19995);
   U21400 : NOR2_X1 port map( A1 => n19991, A2 => n20014, ZN => n19992);
   U21401 : INV_X1 port map( A => n3158, ZN => n23500);
   U21402 : XNOR2_X1 port map( A => n20914, B => n23500, ZN => n19997);
   U21403 : XNOR2_X1 port map( A => n19997, B => n21318, ZN => n20001);
   U21404 : NAND2_X1 port map( A1 => n20447, A2 => n20147, ZN => n20000);
   U21405 : NOR2_X1 port map( A1 => n20536, A2 => n20445, ZN => n20150);
   U21406 : NOR2_X1 port map( A1 => n20537, A2 => n19018, ZN => n19998);
   U21407 : AND2_X1 port map( A1 => n20536, A2 => n20149, ZN => n20148);
   U21408 : NAND2_X1 port map( A1 => n20148, A2 => n19018, ZN => n19999);
   U21409 : XNOR2_X1 port map( A => n20001, B => n20984, ZN => n20002);
   U21410 : AND2_X1 port map( A1 => n20036, A2 => n24905, ZN => n22232);
   U21411 : INV_X1 port map( A => n22232, ZN => n21835);
   U21412 : AOI21_X1 port map( B1 => n20478, B2 => n20003, A => n2168, ZN => 
                           n20004);
   U21414 : NOR2_X1 port map( A1 => n20486, A2 => n24275, ZN => n20005);
   U21415 : INV_X1 port map( A => n20484, ZN => n20910);
   U21416 : AND2_X1 port map( A1 => n20910, A2 => n20909, ZN => n20080);
   U21417 : AOI21_X1 port map( B1 => n20005, B2 => n20360, A => n20080, ZN => 
                           n20007);
   U21418 : NAND3_X1 port map( A1 => n24078, A2 => n20486, A3 => n20911, ZN => 
                           n20006);
   U21419 : NOR2_X1 port map( A1 => n20298, A2 => n20142, ZN => n20010);
   U21420 : OAI21_X1 port map( B1 => n20010, B2 => n20009, A => n20008, ZN => 
                           n20013);
   U21421 : INV_X1 port map( A => n20141, ZN => n20011);
   U21423 : NAND2_X1 port map( A1 => n25242, A2 => n20014, ZN => n20015);
   U21425 : NAND2_X1 port map( A1 => n20135, A2 => n1954, ZN => n20020);
   U21426 : INV_X1 port map( A => n1792, ZN => n20021);
   U21427 : NAND2_X1 port map( A1 => n275, A2 => n20022, ZN => n20026);
   U21428 : NAND3_X1 port map( A1 => n275, A2 => n20562, A3 => n20560, ZN => 
                           n20024);
   U21429 : OAI211_X1 port map( C1 => n25221, C2 => n20026, A => n20025, B => 
                           n20024, ZN => n20798);
   U21430 : NOR2_X1 port map( A1 => n20027, A2 => n3671, ZN => n20031);
   U21431 : NOR2_X1 port map( A1 => n20281, A2 => n19809, ZN => n20029);
   U21432 : NOR2_X1 port map( A1 => n19809, A2 => n1733, ZN => n20028);
   U21433 : AOI22_X1 port map( A1 => n19645, A2 => n20029, B1 => n20028, B2 => 
                           n20345, ZN => n20030);
   U21434 : OAI21_X1 port map( B1 => n20031, B2 => n20345, A => n20030, ZN => 
                           n21142);
   U21435 : XNOR2_X1 port map( A => n20798, B => n21142, ZN => n20032);
   U21436 : XNOR2_X1 port map( A => n20033, B => n20032, ZN => n20034);
   U21437 : XNOR2_X1 port map( A => n20035, B => n20034, ZN => n22225);
   U21438 : INV_X1 port map( A => n22225, ZN => n22235);
   U21439 : OAI22_X1 port map( A1 => n21835, A2 => n22228, B1 => n22235, B2 => 
                           n22233, ZN => n20037);
   U21440 : NOR2_X1 port map( A1 => n20040, A2 => n20042, ZN => n20045);
   U21441 : INV_X1 port map( A => n20046, ZN => n22697);
   U21442 : NOR2_X1 port map( A1 => n20478, A2 => n20477, ZN => n20048);
   U21443 : INV_X1 port map( A => n20476, ZN => n20049);
   U21444 : NAND2_X1 port map( A1 => n20353, A2 => n20049, ZN => n20050);
   U21445 : AND3_X1 port map( A1 => n20051, A2 => n20050, A3 => n20477, ZN => 
                           n20052);
   U21446 : INV_X1 port map( A => n25490, ZN => n20056);
   U21447 : OAI21_X1 port map( B1 => n20056, B2 => n20472, A => n5734, ZN => 
                           n20058);
   U21448 : NAND2_X1 port map( A1 => n20058, A2 => n5115, ZN => n20065);
   U21449 : NOR2_X1 port map( A1 => n20054, A2 => n25089, ZN => n20063);
   U21450 : NOR2_X1 port map( A1 => n20060, A2 => n20473, ZN => n20061);
   U21451 : AOI22_X1 port map( A1 => n20063, A2 => n20062, B1 => n20061, B2 => 
                           n20470, ZN => n20064);
   U21452 : NAND2_X1 port map( A1 => n20065, A2 => n20064, ZN => n21222);
   U21453 : XNOR2_X1 port map( A => n21704, B => n21222, ZN => n20628);
   U21454 : OAI21_X1 port map( B1 => n20909, B2 => n20359, A => n347, ZN => 
                           n20079);
   U21455 : NOR2_X1 port map( A1 => n20076, A2 => n347, ZN => n20078);
   U21456 : NOR2_X1 port map( A1 => n20483, A2 => n20486, ZN => n20077);
   U21458 : OAI21_X1 port map( B1 => n20080, B2 => n20079, A => n20912, ZN => 
                           n20626);
   U21459 : XNOR2_X1 port map( A => n25483, B => n20626, ZN => n20081);
   U21460 : XNOR2_X1 port map( A => n21971, B => n20081, ZN => n20082);
   U21461 : NOR3_X1 port map( A1 => n20616, A2 => n20615, A3 => n20614, ZN => 
                           n20086);
   U21462 : AOI21_X1 port map( B1 => n20572, B2 => n20617, A => n20086, ZN => 
                           n20087);
   U21463 : XNOR2_X1 port map( A => n21521, B => n21676, ZN => n21114);
   U21464 : INV_X1 port map( A => n20557, ZN => n20092);
   U21466 : INV_X1 port map( A => n25221, ZN => n20566);
   U21468 : XNOR2_X1 port map( A => n21192, B => n21114, ZN => n20123);
   U21471 : NAND2_X1 port map( A1 => n20104, A2 => n20103, ZN => n21034);
   U21472 : MUX2_X1 port map( A => n20105, B => n21034, S => n21038, Z => 
                           n20106);
   U21473 : XNOR2_X1 port map( A => n21469, B => n21679, ZN => n20121);
   U21474 : NAND2_X1 port map( A1 => n20111, A2 => n25262, ZN => n20112);
   U21475 : MUX2_X1 port map( A => n20113, B => n20112, S => n25034, Z => 
                           n20119);
   U21476 : NAND2_X1 port map( A1 => n339, A2 => n25388, ZN => n20116);
   U21477 : XNOR2_X1 port map( A => n21601, B => n2744, ZN => n20120);
   U21478 : XNOR2_X1 port map( A => n20121, B => n20120, ZN => n20122);
   U21479 : AND2_X1 port map( A1 => n20546, A2 => n20125, ZN => n20308);
   U21480 : INV_X1 port map( A => n20308, ZN => n20129);
   U21481 : NAND2_X1 port map( A1 => n20545, A2 => n20127, ZN => n20128);
   U21483 : XNOR2_X1 port map( A => n21665, B => n22745, ZN => n20133);
   U21484 : XNOR2_X1 port map( A => n21209, B => n20133, ZN => n20155);
   U21485 : MUX2_X1 port map( A => n20136, B => n20135, S => n25242, Z => 
                           n20138);
   U21486 : MUX2_X2 port map( A => n20139, B => n20138, S => n20137, Z => 
                           n21980);
   U21487 : INV_X1 port map( A => n20140, ZN => n20299);
   U21488 : XNOR2_X1 port map( A => n21554, B => n21980, ZN => n21030);
   U21489 : OAI211_X1 port map( C1 => n20533, C2 => n20447, A => n20147, B => 
                           n20146, ZN => n20153);
   U21490 : NAND2_X1 port map( A1 => n20148, A2 => n20537, ZN => n20152);
   U21491 : NAND2_X1 port map( A1 => n20150, A2 => n20149, ZN => n20151);
   U21493 : XNOR2_X1 port map( A => n21506, B => n21138, ZN => n20898);
   U21494 : XNOR2_X1 port map( A => n21030, B => n20898, ZN => n20154);
   U21495 : XNOR2_X2 port map( A => n20155, B => n20154, ZN => n22356);
   U21496 : MUX2_X1 port map( A => n22355, B => n22361, S => n22356, Z => 
                           n20254);
   U21497 : AND2_X1 port map( A1 => n24454, A2 => n20369, ZN => n20156);
   U21498 : NOR2_X1 port map( A1 => n20451, A2 => n20159, ZN => n20157);
   U21499 : INV_X1 port map( A => n20960, ZN => n20455);
   U21500 : AOI22_X1 port map( A1 => n20157, A2 => n20961, B1 => n20455, B2 => 
                           n20451, ZN => n20162);
   U21501 : INV_X1 port map( A => n20158, ZN => n20160);
   U21502 : NAND3_X1 port map( A1 => n20160, A2 => n20159, A3 => n20377, ZN => 
                           n20161);
   U21503 : XNOR2_X1 port map( A => n21577, B => n1381, ZN => n21199);
   U21504 : INV_X1 port map( A => n20163, ZN => n20164);
   U21505 : OAI21_X1 port map( B1 => n20395, B2 => n24460, A => n20164, ZN => 
                           n20167);
   U21506 : OAI21_X1 port map( B1 => n20458, B2 => n24461, A => n20165, ZN => 
                           n20166);
   U21507 : AND2_X1 port map( A1 => n20167, A2 => n20166, ZN => n21578);
   U21508 : NOR2_X1 port map( A1 => n20169, A2 => n20231, ZN => n20237);
   U21509 : NAND2_X1 port map( A1 => n20237, A2 => n20173, ZN => n20172);
   U21510 : OAI211_X1 port map( C1 => n20170, C2 => n20236, A => n20169, B => 
                           n20168, ZN => n20171);
   U21511 : XNOR2_X1 port map( A => n21998, B => n21578, ZN => n21061);
   U21512 : XNOR2_X1 port map( A => n21061, B => n21199, ZN => n20180);
   U21513 : XNOR2_X1 port map( A => n21997, B => n23151, ZN => n20178);
   U21514 : NAND2_X1 port map( A1 => n20174, A2 => n20588, ZN => n20175);
   U21515 : NAND3_X1 port map( A1 => n20175, A2 => n20590, A3 => n20586, ZN => 
                           n20177);
   U21516 : XNOR2_X1 port map( A => n25386, B => n21106, ZN => n21671);
   U21517 : XNOR2_X1 port map( A => n21671, B => n20178, ZN => n20179);
   U21518 : XNOR2_X1 port map( A => n20179, B => n20180, ZN => n21838);
   U21519 : AOI21_X1 port map( B1 => n20183, B2 => n25211, A => n25478, ZN => 
                           n20190);
   U21520 : OAI21_X1 port map( B1 => n20188, B2 => n20187, A => n20186, ZN => 
                           n20189);
   U21521 : XNOR2_X1 port map( A => n22007, B => n21689, ZN => n21093);
   U21522 : NAND2_X1 port map( A1 => n20195, A2 => n20194, ZN => n20196);
   U21523 : XNOR2_X1 port map( A => n20197, B => n21093, ZN => n20213);
   U21526 : MUX2_X1 port map( A => n20200, B => n20199, S => n20215, Z => 
                           n20201);
   U21527 : INV_X1 port map( A => n20203, ZN => n20205);
   U21528 : AOI22_X1 port map( A1 => n20205, A2 => n20399, B1 => n5733, B2 => 
                           n20204, ZN => n20207);
   U21529 : NAND3_X1 port map( A1 => n20415, A2 => n20401, A3 => n20400, ZN => 
                           n20206);
   U21530 : NOR2_X1 port map( A1 => n20595, A2 => n20599, ZN => n20208);
   U21531 : OAI21_X1 port map( B1 => n1667, B2 => n20426, A => n20595, ZN => 
                           n20211);
   U21532 : NOR2_X1 port map( A1 => n1667, A2 => n25397, ZN => n20210);
   U21533 : XNOR2_X1 port map( A => n20212, B => n21445, ZN => n20642);
   U21535 : MUX2_X1 port map( A => n21782, B => n21839, S => n22361, Z => 
                           n20253);
   U21536 : AOI22_X1 port map( A1 => n24327, A2 => n20215, B1 => n20216, B2 => 
                           n20214, ZN => n20220);
   U21538 : OAI21_X1 port map( B1 => n20276, B2 => n20514, A => n20516, ZN => 
                           n20221);
   U21539 : XNOR2_X1 port map( A => n21495, B => n21568, ZN => n21215);
   U21540 : OAI21_X1 port map( B1 => n3016, B2 => n20226, A => n20268, ZN => 
                           n20227);
   U21542 : NAND2_X1 port map( A1 => n20237, A2 => n20236, ZN => n20238);
   U21543 : XNOR2_X1 port map( A => n21070, B => n21694, ZN => n20251);
   U21544 : NAND3_X1 port map( A1 => n19936, A2 => n20242, A3 => n20241, ZN => 
                           n20247);
   U21548 : XNOR2_X1 port map( A => n21087, B => n673, ZN => n20250);
   U21549 : XNOR2_X1 port map( A => n20251, B => n20250, ZN => n20252);
   U21550 : OR3_X1 port map( A1 => n20255, A2 => n25420, A3 => n20411, ZN => 
                           n20267);
   U21551 : NOR2_X1 port map( A1 => n20256, A2 => n25420, ZN => n20261);
   U21552 : NOR3_X1 port map( A1 => n20259, A2 => n20258, A3 => n20257, ZN => 
                           n20260);
   U21553 : NAND2_X1 port map( A1 => n20261, A2 => n20260, ZN => n20266);
   U21554 : NAND3_X1 port map( A1 => n20411, A2 => n20262, A3 => n25421, ZN => 
                           n20265);
   U21555 : XNOR2_X1 port map( A => n21172, B => n20804, ZN => n21409);
   U21556 : MUX2_X2 port map( A => n20271, B => n20270, S => n20497, Z => 
                           n21501);
   U21557 : NAND2_X1 port map( A1 => n20515, A2 => n20272, ZN => n20273);
   U21558 : XNOR2_X1 port map( A => n21501, B => n21658, ZN => n21302);
   U21559 : XNOR2_X1 port map( A => n21409, B => n21302, ZN => n20288);
   U21560 : NOR2_X1 port map( A1 => n20280, A2 => n20343, ZN => n20282);
   U21562 : XNOR2_X1 port map( A => n20475, B => n20284, ZN => n20286);
   U21563 : XNOR2_X1 port map( A => n20285, B => n20286, ZN => n20287);
   U21564 : NAND2_X1 port map( A1 => n20289, A2 => n21008, ZN => n20293);
   U21565 : NAND2_X1 port map( A1 => n20290, A2 => n20522, ZN => n20292);
   U21566 : AOI21_X1 port map( B1 => n20293, B2 => n20292, A => n20291, ZN => 
                           n20294);
   U21568 : OAI21_X1 port map( B1 => n20298, B2 => n20297, A => n20296, ZN => 
                           n20300);
   U21569 : XNOR2_X1 port map( A => n25470, B => n21985, ZN => n20307);
   U21570 : NAND3_X1 port map( A1 => n3428, A2 => n24558, A3 => n24454, ZN => 
                           n20304);
   U21572 : XNOR2_X1 port map( A => n21569, B => n5514, ZN => n20306);
   U21573 : XNOR2_X1 port map( A => n20307, B => n20306, ZN => n20315);
   U21574 : XNOR2_X1 port map( A => n21399, B => n25222, ZN => n20313);
   U21575 : NOR2_X1 port map( A1 => n20308, A2 => n20543, ZN => n20311);
   U21576 : XNOR2_X1 port map( A => n21324, B => n21247, ZN => n20990);
   U21577 : XNOR2_X1 port map( A => n20313, B => n20990, ZN => n20314);
   U21579 : XNOR2_X1 port map( A => n21686, B => n1757, ZN => n20324);
   U21583 : INV_X1 port map( A => n20554, ZN => n20333);
   U21584 : OAI21_X1 port map( B1 => n20554, B2 => n20555, A => n20330, ZN => 
                           n20331);
   U21585 : NAND2_X1 port map( A1 => n20670, A2 => n20335, ZN => n20350);
   U21586 : NAND3_X1 port map( A1 => n20338, A2 => n20337, A3 => n20336, ZN => 
                           n20339);
   U21587 : OAI211_X1 port map( C1 => n20350, C2 => n20341, A => n20340, B => 
                           n20339, ZN => n21157);
   U21588 : XNOR2_X1 port map( A => n20798, B => n21157, ZN => n21420);
   U21589 : XNOR2_X1 port map( A => n21420, B => n21343, ZN => n20342);
   U21590 : NOR2_X1 port map( A1 => n24414, A2 => n1733, ZN => n20344);
   U21592 : OAI211_X1 port map( C1 => n24414, C2 => n19809, A => n20345, B => 
                           n1733, ZN => n20347);
   U21594 : XNOR2_X1 port map( A => n20780, B => n21334, ZN => n20358);
   U21595 : OAI21_X1 port map( B1 => n20353, B2 => n20480, A => n20352, ZN => 
                           n20357);
   U21598 : XNOR2_X1 port map( A => n21058, B => n21511, ZN => n20889);
   U21599 : XNOR2_X1 port map( A => n20358, B => n20889, ZN => n20366);
   U21600 : OAI211_X1 port map( C1 => n20360, C2 => n20491, A => n20486, B => 
                           n20359, ZN => n20361);
   U21602 : XNOR2_X1 port map( A => n21996, B => n21515, ZN => n21668);
   U21603 : XNOR2_X1 port map( A => n20999, B => n2757, ZN => n20364);
   U21604 : XNOR2_X1 port map( A => n21668, B => n20364, ZN => n20365);
   U21605 : XNOR2_X1 port map( A => n20366, B => n20365, ZN => n22655);
   U21606 : NOR2_X1 port map( A1 => n20368, A2 => n24558, ZN => n20372);
   U21607 : NOR2_X2 port map( A1 => n20376, A2 => n20375, ZN => n21429);
   U21609 : OAI21_X1 port map( B1 => n20377, B2 => n20451, A => n20961, ZN => 
                           n20381);
   U21610 : OAI21_X1 port map( B1 => n2688, B2 => n20451, A => n24357, ZN => 
                           n20379);
   U21611 : OAI21_X1 port map( B1 => n20961, B2 => n20448, A => n20960, ZN => 
                           n20378);
   U21612 : NAND2_X1 port map( A1 => n20379, A2 => n20378, ZN => n20380);
   U21613 : XNOR2_X1 port map( A => n21429, B => n21633, ZN => n21317);
   U21614 : NAND2_X1 port map( A1 => n20385, A2 => n20459, ZN => n20397);
   U21616 : AND2_X1 port map( A1 => n20388, A2 => n20389, ZN => n20391);
   U21617 : OAI21_X1 port map( B1 => n20392, B2 => n20391, A => n20390, ZN => 
                           n20393);
   U21619 : XNOR2_X1 port map( A => n21965, B => n21532, ZN => n21701);
   U21620 : XNOR2_X1 port map( A => n25495, B => n21701, ZN => n20408);
   U21621 : MUX2_X1 port map( A => n20400, B => n20399, S => n20422, Z => 
                           n20405);
   U21622 : NOR2_X1 port map( A1 => n20415, A2 => n20414, ZN => n20403);
   U21623 : AOI22_X1 port map( A1 => n20403, A2 => n20422, B1 => n20402, B2 => 
                           n20419, ZN => n20404);
   U21625 : XNOR2_X1 port map( A => n24353, B => n2847, ZN => n20406);
   U21626 : XNOR2_X1 port map( A => n20406, B => n20984, ZN => n20407);
   U21627 : XNOR2_X1 port map( A => n21600, B => n891, ZN => n20424);
   U21628 : NAND2_X1 port map( A1 => n20415, A2 => n20414, ZN => n20423);
   U21629 : NAND2_X1 port map( A1 => n20416, A2 => n20419, ZN => n20421);
   U21631 : XNOR2_X1 port map( A => n21310, B => n24936, ZN => n21415);
   U21632 : XNOR2_X1 port map( A => n21415, B => n20424, ZN => n20441);
   U21633 : NOR2_X1 port map( A1 => n20427, A2 => n20599, ZN => n20429);
   U21634 : AOI22_X1 port map( A1 => n20597, A2 => n20430, B1 => n20429, B2 => 
                           n25397, ZN => n20431);
   U21635 : NAND2_X1 port map( A1 => n20432, A2 => n20577, ZN => n20436);
   U21636 : OAI211_X1 port map( C1 => n20438, C2 => n20437, A => n20436, B => 
                           n20435, ZN => n22014);
   U21637 : XNOR2_X1 port map( A => n21308, B => n20439, ZN => n20440);
   U21638 : NAND2_X1 port map( A1 => n25075, A2 => n22655, ZN => n20442);
   U21639 : NAND2_X1 port map( A1 => n20443, A2 => n22656, ZN => n20444);
   U21640 : AOI21_X1 port map( B1 => n20537, B2 => n20536, A => n20445, ZN => 
                           n20446);
   U21641 : XNOR2_X1 port map( A => n21721, B => n25385, ZN => n20457);
   U21642 : AOI21_X1 port map( B1 => n24354, B2 => n20448, A => n20450, ZN => 
                           n20456);
   U21645 : XNOR2_X1 port map( A => n21246, B => n20457, ZN => n20467);
   U21646 : OAI211_X1 port map( C1 => n20461, C2 => n1327, A => n20460, B => 
                           n20459, ZN => n20463);
   U21647 : XNOR2_X1 port map( A => n21621, B => n21693, ZN => n21167);
   U21648 : INV_X1 port map( A => Key(60), ZN => n22089);
   U21649 : XNOR2_X1 port map( A => n21167, B => n20465, ZN => n20466);
   U21650 : XNOR2_X1 port map( A => n20466, B => n20467, ZN => n22770);
   U21651 : INV_X1 port map( A => n22770, ZN => n22680);
   U21652 : NAND2_X1 port map( A1 => n25490, A2 => n20472, ZN => n20474);
   U21653 : XNOR2_X1 port map( A => n21173, B => n20475, ZN => n21551);
   U21654 : MUX2_X1 port map( A => n20477, B => n20476, S => n20479, Z => 
                           n20481);
   U21655 : XNOR2_X1 port map( A => n21301, B => n21040, ZN => n21406);
   U21656 : XNOR2_X1 port map( A => n21551, B => n21406, ZN => n20495);
   U21657 : XNOR2_X1 port map( A => n21745, B => n3129, ZN => n20493);
   U21659 : NOR2_X1 port map( A1 => n20484, A2 => n20491, ZN => n20485);
   U21661 : INV_X1 port map( A => n20487, ZN => n20488);
   U21662 : NAND2_X1 port map( A1 => n20488, A2 => n20491, ZN => n20489);
   U21663 : XNOR2_X1 port map( A => n21027, B => n20964, ZN => n21618);
   U21664 : XNOR2_X1 port map( A => n21618, B => n20493, ZN => n20494);
   U21666 : NOR2_X1 port map( A1 => n3016, A2 => n20501, ZN => n20499);
   U21667 : INV_X1 port map( A => n21193, ZN => n20503);
   U21668 : XNOR2_X1 port map( A => n21414, B => n20503, ZN => n20505);
   U21669 : XNOR2_X1 port map( A => n21312, B => n886, ZN => n20504);
   U21670 : OAI22_X1 port map( A1 => n20511, A2 => n20510, B1 => n24327, B2 => 
                           n20508, ZN => n20512);
   U21671 : XNOR2_X1 port map( A => n21307, B => n21675, ZN => n20769);
   U21672 : XNOR2_X1 port map( A => n20769, B => n20948, ZN => n21156);
   U21673 : XNOR2_X2 port map( A => n20521, B => n21156, ZN => n22774);
   U21674 : MUX2_X1 port map( A => n22680, B => n21856, S => n22774, Z => 
                           n20608);
   U21675 : INV_X1 port map( A => n20522, ZN => n20525);
   U21676 : NAND2_X1 port map( A1 => n20525, A2 => n20523, ZN => n20527);
   U21678 : AOI21_X1 port map( B1 => n20530, B2 => n24581, A => n20528, ZN => 
                           n20531);
   U21679 : NOR2_X1 port map( A1 => n21013, A2 => n20531, ZN => n21045);
   U21680 : OAI211_X1 port map( C1 => n20533, C2 => n19018, A => n20536, B => 
                           n20532, ZN => n20542);
   U21681 : INV_X1 port map( A => n20534, ZN => n20535);
   U21682 : NAND2_X1 port map( A1 => n20539, A2 => n20535, ZN => n20541);
   U21683 : INV_X1 port map( A => n20536, ZN => n20538);
   U21684 : NAND3_X1 port map( A1 => n20539, A2 => n20538, A3 => n20537, ZN => 
                           n20540);
   U21686 : XNOR2_X1 port map( A => n21422, B => n21045, ZN => n20762);
   U21687 : NAND2_X1 port map( A1 => n20544, A2 => n20543, ZN => n20547);
   U21688 : XNOR2_X1 port map( A => n24485, B => n21158, ZN => n21593);
   U21689 : XNOR2_X1 port map( A => n20762, B => n21593, ZN => n20553);
   U21690 : XNOR2_X1 port map( A => n21751, B => n2145, ZN => n20550);
   U21691 : XNOR2_X1 port map( A => n20551, B => n20550, ZN => n20552);
   U21692 : XNOR2_X1 port map( A => n20553, B => n20552, ZN => n22769);
   U21693 : INV_X1 port map( A => n22769, ZN => n22369);
   U21694 : AND2_X1 port map( A1 => n20556, A2 => n20555, ZN => n20558);
   U21695 : AND2_X1 port map( A1 => n20561, A2 => n20560, ZN => n20565);
   U21696 : XNOR2_X1 port map( A => n21182, B => n21579, ZN => n20781);
   U21697 : XNOR2_X1 port map( A => n20781, B => n20568, ZN => n20575);
   U21698 : XNOR2_X1 port map( A => n21058, B => n24100, ZN => n21252);
   U21699 : XNOR2_X1 port map( A => n21729, B => n2100, ZN => n20573);
   U21700 : XNOR2_X1 port map( A => n21252, B => n20573, ZN => n20574);
   U21702 : NAND2_X1 port map( A1 => n22369, A2 => n22679, ZN => n20606);
   U21703 : NAND3_X1 port map( A1 => n20577, A2 => n20576, A3 => n24940, ZN => 
                           n20581);
   U21704 : NOR2_X1 port map( A1 => n24940, A2 => n5208, ZN => n20579);
   U21705 : NAND2_X1 port map( A1 => n20583, A2 => n20579, ZN => n20580);
   U21706 : XNOR2_X1 port map( A => n20914, B => n21053, ZN => n21635);
   U21707 : INV_X1 port map( A => n21738, ZN => n21478);
   U21708 : XNOR2_X1 port map( A => n21478, B => Key(149), ZN => n20584);
   U21709 : XNOR2_X1 port map( A => n21635, B => n20584, ZN => n20604);
   U21710 : INV_X1 port map( A => n20585, ZN => n20594);
   U21711 : MUX2_X1 port map( A => n20588, B => n20587, S => n20586, Z => 
                           n20592);
   U21712 : OAI21_X1 port map( B1 => n276, B2 => n20595, A => n20599, ZN => 
                           n20601);
   U21713 : NOR3_X1 port map( A1 => n24463, A2 => n20599, A3 => n20598, ZN => 
                           n20600);
   U21714 : XNOR2_X1 port map( A => n21318, B => n21734, ZN => n21433);
   U21715 : XNOR2_X1 port map( A => n21562, B => n21433, ZN => n20603);
   U21716 : MUX2_X1 port map( A => n20606, B => n20605, S => n21856, Z => 
                           n20607);
   U21718 : INV_X1 port map( A => n23859, ZN => n23839);
   U21719 : INV_X1 port map( A => n20609, ZN => n20625);
   U21720 : XNOR2_X1 port map( A => n21694, B => n2795, ZN => n20610);
   U21721 : XNOR2_X1 port map( A => n21215, B => n20610, ZN => n20613);
   U21722 : XNOR2_X1 port map( A => n24996, B => n25073, ZN => n20611);
   U21723 : XNOR2_X1 port map( A => n21132, B => n21135, ZN => n21725);
   U21724 : XNOR2_X1 port map( A => n20611, B => n21725, ZN => n20612);
   U21725 : XNOR2_X1 port map( A => n20612, B => n20613, ZN => n21908);
   U21726 : INV_X1 port map( A => n21908, ZN => n22338);
   U21727 : XNOR2_X1 port map( A => n21319, B => n21481, ZN => n21739);
   U21728 : NAND2_X1 port map( A1 => n20615, A2 => n20614, ZN => n20622);
   U21729 : MUX2_X1 port map( A => n20617, B => n20616, S => n20615, Z => 
                           n20620);
   U21730 : MUX2_X1 port map( A => n20620, B => n20619, S => n7, Z => n20621);
   U21732 : XNOR2_X1 port map( A => n24353, B => n21630, ZN => n20624);
   U21733 : XNOR2_X1 port map( A => n21739, B => n20624, ZN => n20630);
   U21734 : XNOR2_X1 port map( A => n20626, B => n20625, ZN => n20627);
   U21735 : XNOR2_X1 port map( A => n20628, B => n20627, ZN => n20629);
   U21736 : XNOR2_X1 port map( A => n20630, B => n20629, ZN => n22137);
   U21737 : NOR2_X1 port map( A1 => n22338, A2 => n22137, ZN => n22336);
   U21738 : XNOR2_X1 port map( A => n21138, B => n21743, ZN => n21457);
   U21739 : XNOR2_X1 port map( A => n21505, B => n876, ZN => n20631);
   U21740 : XNOR2_X1 port map( A => n20631, B => n21457, ZN => n20633);
   U21741 : XNOR2_X1 port map( A => n21259, B => n21300, ZN => n20632);
   U21742 : XNOR2_X1 port map( A => n20633, B => n20632, ZN => n20635);
   U21744 : XNOR2_X1 port map( A => n21639, B => n1920, ZN => n20636);
   U21745 : XNOR2_X1 port map( A => n21192, B => n20636, ZN => n20639);
   U21746 : XNOR2_X1 port map( A => n21306, B => n20870, ZN => n21716);
   U21747 : XNOR2_X1 port map( A => n21676, B => n21600, ZN => n20637);
   U21748 : XNOR2_X1 port map( A => n20637, B => n21716, ZN => n20638);
   U21749 : AND2_X1 port map( A1 => n22139, A2 => n22338, ZN => n20649);
   U21750 : XNOR2_X1 port map( A => n20882, B => n688, ZN => n20640);
   U21751 : XNOR2_X1 port map( A => n20640, B => n21541, ZN => n20641);
   U21752 : XNOR2_X1 port map( A => n20826, B => n21042, ZN => n21755);
   U21753 : XNOR2_X1 port map( A => n20641, B => n21755, ZN => n20643);
   U21754 : XNOR2_X1 port map( A => n21336, B => n21058, ZN => n21584);
   U21755 : XNOR2_X1 port map( A => n21199, B => n21584, ZN => n20647);
   U21756 : XNOR2_X1 port map( A => n21514, B => n21728, ZN => n20645);
   U21757 : XNOR2_X1 port map( A => n25387, B => n3073, ZN => n20644);
   U21758 : XNOR2_X1 port map( A => n20645, B => n20644, ZN => n20646);
   U21759 : XNOR2_X1 port map( A => n20647, B => n20646, ZN => n22138);
   U21760 : AND2_X1 port map( A1 => n22138, A2 => n22338, ZN => n20648);
   U21761 : INV_X1 port map( A => n22139, ZN => n22141);
   U21762 : NOR2_X1 port map( A1 => n22338, A2 => n22139, ZN => n20650);
   U21763 : XNOR2_X1 port map( A => n21414, B => n21678, ZN => n20651);
   U21764 : XNOR2_X1 port map( A => n21308, B => n20651, ZN => n20656);
   U21765 : XNOR2_X1 port map( A => n20948, B => n21679, ZN => n20654);
   U21766 : INV_X1 port map( A => n62, ZN => n20652);
   U21767 : XNOR2_X1 port map( A => n24936, B => n20652, ZN => n20653);
   U21768 : XNOR2_X1 port map( A => n20654, B => n20653, ZN => n20655);
   U21770 : XNOR2_X1 port map( A => n21996, B => n21511, ZN => n21333);
   U21771 : XNOR2_X1 port map( A => n21333, B => n21184, ZN => n20660);
   U21772 : XNOR2_X1 port map( A => n24100, B => n21670, ZN => n20658);
   U21773 : XNOR2_X1 port map( A => n20999, B => n2903, ZN => n20657);
   U21774 : XNOR2_X1 port map( A => n20658, B => n20657, ZN => n20659);
   U21775 : XNOR2_X1 port map( A => n20660, B => n20659, ZN => n22973);
   U21776 : AND2_X1 port map( A1 => n22977, A2 => n3213, ZN => n20684);
   U21777 : XNOR2_X1 port map( A => n20957, B => n21696, ZN => n20664);
   U21778 : XNOR2_X1 port map( A => n21492, B => n21399, ZN => n20662);
   U21779 : XNOR2_X1 port map( A => n25377, B => n912, ZN => n20661);
   U21780 : XNOR2_X1 port map( A => n20662, B => n20661, ZN => n20663);
   U21781 : INV_X1 port map( A => n20665, ZN => n20675);
   U21782 : NAND2_X1 port map( A1 => n20666, A2 => n20669, ZN => n20667);
   U21783 : OAI211_X1 port map( C1 => n20670, C2 => n20669, A => n20668, B => 
                           n20667, ZN => n20674);
   U21784 : NAND2_X1 port map( A1 => n20672, A2 => n20671, ZN => n20673);
   U21785 : NAND3_X1 port map( A1 => n20675, A2 => n20674, A3 => n20673, ZN => 
                           n20676);
   U21786 : XNOR2_X1 port map( A => n20676, B => n681, ZN => n20678);
   U21787 : XNOR2_X1 port map( A => n21734, B => n21699, ZN => n20677);
   U21788 : XNOR2_X1 port map( A => n20914, B => n21965, ZN => n20972);
   U21789 : XNOR2_X1 port map( A => n20804, B => n21665, ZN => n20680);
   U21790 : XNOR2_X1 port map( A => n21302, B => n20680, ZN => n20683);
   U21791 : XNOR2_X1 port map( A => n21205, B => n20964, ZN => n20899);
   U21792 : XNOR2_X1 port map( A => n21040, B => n1896, ZN => n20681);
   U21793 : XNOR2_X1 port map( A => n20899, B => n20681, ZN => n20682);
   U21794 : XNOR2_X2 port map( A => n20683, B => n20682, ZN => n22387);
   U21795 : XNOR2_X1 port map( A => n21689, B => n21160, ZN => n20945);
   U21796 : XNOR2_X1 port map( A => n20798, B => n21228, ZN => n20736);
   U21797 : XNOR2_X1 port map( A => n20945, B => n20736, ZN => n20687);
   U21798 : XNOR2_X1 port map( A => n21422, B => n1827, ZN => n20685);
   U21799 : XNOR2_X1 port map( A => n21343, B => n20685, ZN => n20686);
   U21800 : XNOR2_X1 port map( A => n20687, B => n20686, ZN => n22972);
   U21802 : OR2_X1 port map( A1 => n22387, A2 => n22972, ZN => n22293);
   U21803 : OAI21_X1 port map( B1 => n25365, B2 => n21891, A => n22293, ZN => 
                           n20688);
   U21804 : NOR2_X1 port map( A1 => n23218, A2 => n23220, ZN => n23215);
   U21805 : XNOR2_X1 port map( A => n21301, B => n21554, ZN => n21207);
   U21806 : XNOR2_X1 port map( A => n21975, B => n21258, ZN => n20689);
   U21807 : XNOR2_X1 port map( A => n21207, B => n20689, ZN => n20694);
   U21808 : XNOR2_X1 port map( A => n24491, B => n21138, ZN => n20692);
   U21809 : INV_X1 port map( A => n20690, ZN => n22625);
   U21810 : XNOR2_X1 port map( A => n21172, B => n22625, ZN => n20691);
   U21811 : XNOR2_X1 port map( A => n20692, B => n20691, ZN => n20693);
   U21812 : INV_X1 port map( A => n2717, ZN => n22549);
   U21813 : XNOR2_X1 port map( A => n21573, B => n22549, ZN => n20696);
   U21814 : XNOR2_X1 port map( A => n21622, B => n21324, ZN => n20695);
   U21815 : XNOR2_X1 port map( A => n20696, B => n20695, ZN => n20699);
   U21816 : XNOR2_X1 port map( A => n21694, B => n21720, ZN => n21460);
   U21817 : XNOR2_X1 port map( A => n20697, B => n21070, ZN => n21216);
   U21818 : XNOR2_X1 port map( A => n21216, B => n21460, ZN => n20698);
   U21819 : XNOR2_X1 port map( A => n20699, B => n20698, ZN => n21934);
   U21820 : INV_X1 port map( A => n21318, ZN => n20701);
   U21821 : XNOR2_X1 port map( A => n21561, B => n22702, ZN => n20702);
   U21822 : XNOR2_X1 port map( A => n20867, B => n20702, ZN => n20705);
   U21823 : XNOR2_X1 port map( A => n21735, B => n21704, ZN => n21480);
   U21824 : INV_X1 port map( A => n21480, ZN => n20703);
   U21825 : XNOR2_X1 port map( A => n20703, B => n21429, ZN => n20704);
   U21827 : XNOR2_X1 port map( A => n21445, B => n21227, ZN => n20707);
   U21828 : XNOR2_X1 port map( A => n21157, B => n1776, ZN => n20706);
   U21829 : XNOR2_X1 port map( A => n20707, B => n20706, ZN => n20710);
   U21830 : XNOR2_X1 port map( A => n21229, B => n20708, ZN => n20709);
   U21831 : INV_X1 port map( A => n21934, ZN => n22563);
   U21832 : XNOR2_X1 port map( A => n21310, B => n25265, ZN => n21153);
   U21833 : XNOR2_X1 port map( A => n20831, B => n21153, ZN => n20713);
   U21834 : INV_X1 port map( A => n24287, ZN => n22767);
   U21835 : XNOR2_X1 port map( A => n21676, B => n22767, ZN => n20711);
   U21836 : XNOR2_X1 port map( A => n21601, B => n21312, ZN => n21191);
   U21837 : XNOR2_X1 port map( A => n21191, B => n20711, ZN => n20712);
   U21838 : XNOR2_X2 port map( A => n20712, B => n20713, ZN => n22409);
   U21839 : OAI21_X1 port map( B1 => n22406, B2 => n24951, A => n20714, ZN => 
                           n20721);
   U21840 : XNOR2_X1 port map( A => n21331, B => n21578, ZN => n21198);
   U21841 : XNOR2_X1 port map( A => n21253, B => n21198, ZN => n20718);
   U21842 : XNOR2_X1 port map( A => n21582, B => n21334, ZN => n20716);
   U21843 : XNOR2_X1 port map( A => n25386, B => n1864, ZN => n20715);
   U21844 : XNOR2_X1 port map( A => n20716, B => n20715, ZN => n20717);
   U21845 : XNOR2_X1 port map( A => n20718, B => n20717, ZN => n22407);
   U21846 : NAND2_X1 port map( A1 => n24971, A2 => n22407, ZN => n20719);
   U21847 : AOI21_X1 port map( B1 => n22132, B2 => n20719, A => n22133, ZN => 
                           n20720);
   U21849 : INV_X1 port map( A => n24955, ZN => n23229);
   U21850 : XNOR2_X1 port map( A => n21454, B => n20722, ZN => n20726);
   U21851 : XNOR2_X1 port map( A => n21505, B => n1826, ZN => n20724);
   U21852 : XNOR2_X1 port map( A => n20724, B => n20723, ZN => n20725);
   U21853 : XNOR2_X1 port map( A => n20725, B => n20726, ZN => n21380);
   U21854 : XNOR2_X1 port map( A => n21399, B => n21212, ZN => n20729);
   U21855 : XNOR2_X1 port map( A => n20727, B => n2208, ZN => n20728);
   U21856 : XNOR2_X1 port map( A => n20728, B => n20729, ZN => n20731);
   U21857 : XNOR2_X1 port map( A => n21721, B => n21087, ZN => n21461);
   U21858 : XNOR2_X1 port map( A => n21461, B => n20954, ZN => n20730);
   U21859 : XNOR2_X1 port map( A => n21514, B => n21998, ZN => n20732);
   U21860 : XNOR2_X1 port map( A => n20732, B => n24985, ZN => n21110);
   U21861 : XNOR2_X1 port map( A => n20733, B => n20999, ZN => n20734);
   U21862 : XNOR2_X1 port map( A => n20734, B => n21121, ZN => n20735);
   U21863 : XNOR2_X1 port map( A => n21587, B => n21541, ZN => n20737);
   U21864 : XNOR2_X1 port map( A => n20736, B => n20737, ZN => n20740);
   U21865 : XNOR2_X1 port map( A => n22007, B => n21751, ZN => n21449);
   U21866 : XNOR2_X1 port map( A => n22006, B => n881, ZN => n20738);
   U21867 : XNOR2_X1 port map( A => n21449, B => n20738, ZN => n20739);
   U21868 : XNOR2_X1 port map( A => n20739, B => n20740, ZN => n22455);
   U21869 : XNOR2_X1 port map( A => n20741, B => n21967, ZN => n20743);
   U21870 : XNOR2_X1 port map( A => n21559, B => n20742, ZN => n20969);
   U21871 : XNOR2_X1 port map( A => n20743, B => n20969, ZN => n20746);
   U21872 : INV_X1 port map( A => n20744, ZN => n23183);
   U21873 : XNOR2_X1 port map( A => n21469, B => n21713, ZN => n22012);
   U21874 : XNOR2_X1 port map( A => n22012, B => n21116, ZN => n20750);
   U21875 : XNOR2_X1 port map( A => n21193, B => n24936, ZN => n20748);
   U21876 : XNOR2_X1 port map( A => n21639, B => Key(190), ZN => n20747);
   U21877 : XNOR2_X1 port map( A => n20748, B => n20747, ZN => n20749);
   U21878 : NOR2_X1 port map( A1 => n1352, A2 => n22453, ZN => n22326);
   U21879 : NOR2_X1 port map( A1 => n23229, A2 => n23227, ZN => n20787);
   U21880 : XNOR2_X1 port map( A => n21027, B => n21297, ZN => n21005);
   U21881 : XNOR2_X1 port map( A => n21975, B => n23750, ZN => n20751);
   U21882 : XNOR2_X1 port map( A => n21005, B => n20751, ZN => n20753);
   U21883 : XNOR2_X1 port map( A => n21616, B => n21040, ZN => n21262);
   U21884 : XNOR2_X1 port map( A => n21173, B => n21136, ZN => n20808);
   U21885 : XNOR2_X1 port map( A => n20808, B => n21262, ZN => n20752);
   U21886 : XNOR2_X1 port map( A => n20753, B => n20752, ZN => n22134);
   U21887 : XNOR2_X1 port map( A => n21133, B => n21247, ZN => n21626);
   U21888 : XNOR2_X1 port map( A => n21245, B => n21693, ZN => n20992);
   U21889 : XNOR2_X1 port map( A => n20992, B => n21626, ZN => n20757);
   U21890 : XNOR2_X1 port map( A => n21573, B => n1801, ZN => n20755);
   U21891 : XNOR2_X1 port map( A => n25377, B => n25385, ZN => n20754);
   U21892 : XNOR2_X1 port map( A => n20755, B => n20754, ZN => n20756);
   U21893 : XNOR2_X1 port map( A => n20757, B => n20756, ZN => n21888);
   U21894 : AND2_X1 port map( A1 => n22134, A2 => n22401, ZN => n20775);
   U21895 : XNOR2_X1 port map( A => n21126, B => n21273, ZN => n21632);
   U21896 : XNOR2_X1 port map( A => n21561, B => n21053, ZN => n20758);
   U21897 : XNOR2_X1 port map( A => n21632, B => n20758, ZN => n20761);
   U21898 : XNOR2_X1 port map( A => n21176, B => n20982, ZN => n21316);
   U21899 : XNOR2_X1 port map( A => n21734, B => n3344, ZN => n20759);
   U21900 : XNOR2_X1 port map( A => n20759, B => n21316, ZN => n20760);
   U21901 : XNOR2_X1 port map( A => n20761, B => n20760, ZN => n22397);
   U21902 : XNOR2_X1 port map( A => n21158, B => n21142, ZN => n20797);
   U21903 : XNOR2_X1 port map( A => n20762, B => n20797, ZN => n20766);
   U21904 : XNOR2_X1 port map( A => n21227, B => n21266, ZN => n20764);
   U21905 : XNOR2_X1 port map( A => n21267, B => n2222, ZN => n20763);
   U21906 : XNOR2_X1 port map( A => n20764, B => n20763, ZN => n20765);
   U21907 : XNOR2_X1 port map( A => n20766, B => n20765, ZN => n20776);
   U21908 : INV_X1 port map( A => n20776, ZN => n22265);
   U21909 : NOR2_X1 port map( A1 => n22265, A2 => n22401, ZN => n20774);
   U21910 : INV_X1 port map( A => n21311, ZN => n20768);
   U21911 : XNOR2_X1 port map( A => n20768, B => n20767, ZN => n21241);
   U21912 : XNOR2_X1 port map( A => n21241, B => n20769, ZN => n20773);
   U21913 : XNOR2_X1 port map( A => n21414, B => n21115, ZN => n20771);
   U21914 : XNOR2_X1 port map( A => n21596, B => n765, ZN => n20770);
   U21915 : XNOR2_X1 port map( A => n20771, B => n20770, ZN => n20772);
   U21917 : AOI22_X1 port map( A1 => n20775, A2 => n22397, B1 => n20774, B2 => 
                           n22398, ZN => n20786);
   U21918 : INV_X1 port map( A => n2049, ZN => n20777);
   U21919 : XNOR2_X1 port map( A => n20779, B => n21648, ZN => n20783);
   U21920 : XNOR2_X1 port map( A => n21332, B => n20780, ZN => n21254);
   U21921 : XNOR2_X1 port map( A => n21254, B => n20781, ZN => n20782);
   U21922 : AOI21_X1 port map( B1 => n25381, B2 => n22400, A => n22134, ZN => 
                           n20784);
   U21923 : OAI21_X1 port map( B1 => n22400, B2 => n21885, A => n20784, ZN => 
                           n20785);
   U21925 : OAI21_X1 port map( B1 => n23215, B2 => n20787, A => n23231, ZN => 
                           n20824);
   U21926 : INV_X1 port map( A => n1340, ZN => n23213);
   U21928 : XNOR2_X1 port map( A => n21108, B => n21668, ZN => n20791);
   U21929 : XNOR2_X1 port map( A => n21579, B => n25091, ZN => n20789);
   U21930 : XNOR2_X1 port map( A => n20999, B => n3798, ZN => n20788);
   U21931 : XNOR2_X1 port map( A => n20789, B => n20788, ZN => n20790);
   U21932 : XNOR2_X1 port map( A => n20791, B => n20790, ZN => n21375);
   U21934 : XNOR2_X1 port map( A => n21307, B => n24916, ZN => n20794);
   U21935 : XNOR2_X1 port map( A => n20792, B => n812, ZN => n20793);
   U21936 : INV_X1 port map( A => n21523, ZN => n20927);
   U21938 : XNOR2_X1 port map( A => n20795, B => n20927, ZN => n21683);
   U21939 : XNOR2_X1 port map( A => n22005, B => n21444, ZN => n21684);
   U21940 : XNOR2_X1 port map( A => n20797, B => n21684, ZN => n20802);
   U21941 : XNOR2_X1 port map( A => n20798, B => n21141, ZN => n20800);
   U21942 : XNOR2_X1 port map( A => n21686, B => n2726, ZN => n20799);
   U21943 : XNOR2_X1 port map( A => n20800, B => n20799, ZN => n20801);
   U21945 : NOR2_X1 port map( A1 => n1363, A2 => n22459, ZN => n20803);
   U21946 : XNOR2_X1 port map( A => n20804, B => n21979, ZN => n20807);
   U21947 : XNOR2_X1 port map( A => n21658, B => n20805, ZN => n20806);
   U21948 : XNOR2_X1 port map( A => n20807, B => n20806, ZN => n20810);
   U21949 : XNOR2_X1 port map( A => n21659, B => n21660, ZN => n21503);
   U21950 : XNOR2_X1 port map( A => n20808, B => n21503, ZN => n20809);
   U21951 : XNOR2_X1 port map( A => n21971, B => n21701, ZN => n20813);
   U21952 : XNOR2_X1 port map( A => n21567, B => n921, ZN => n20815);
   U21953 : XNOR2_X1 port map( A => n20817, B => n20816, ZN => n20819);
   U21955 : XNOR2_X2 port map( A => n20819, B => n21697, ZN => n22464);
   U21956 : AOI21_X1 port map( B1 => n22462, B2 => n22465, A => n3908, ZN => 
                           n20821);
   U21957 : NAND2_X1 port map( A1 => n21929, A2 => n24367, ZN => n20820);
   U21958 : AOI21_X1 port map( B1 => n23213, B2 => n23219, A => n20822, ZN => 
                           n20823);
   U21959 : INV_X1 port map( A => n20825, ZN => n21398);
   U21960 : XNOR2_X1 port map( A => n21449, B => n22004, ZN => n20829);
   U21961 : XNOR2_X1 port map( A => n21686, B => n1835, ZN => n20827);
   U21962 : XNOR2_X1 port map( A => n20881, B => n20827, ZN => n20828);
   U21963 : XNOR2_X1 port map( A => n20829, B => n20828, ZN => n20845);
   U21964 : INV_X1 port map( A => n20845, ZN => n22176);
   U21965 : XNOR2_X1 port map( A => n21193, B => n21469, ZN => n20830);
   U21966 : XNOR2_X1 port map( A => n20831, B => n20830, ZN => n20835);
   U21967 : XNOR2_X1 port map( A => n21520, B => n21523, ZN => n20833);
   U21968 : XNOR2_X1 port map( A => n20870, B => n859, ZN => n20832);
   U21969 : XNOR2_X1 port map( A => n20833, B => n20832, ZN => n20834);
   U21970 : XNOR2_X1 port map( A => n21087, B => n21495, ZN => n21986);
   U21971 : XNOR2_X1 port map( A => n21135, B => n21622, ZN => n20860);
   U21972 : XNOR2_X1 port map( A => n21986, B => n20860, ZN => n20838);
   U21973 : XNOR2_X1 port map( A => n25222, B => n1855, ZN => n20836);
   U21974 : XNOR2_X1 port map( A => n25442, B => n20836, ZN => n20837);
   U21975 : XNOR2_X2 port map( A => n20837, B => n20838, ZN => n22175);
   U21976 : BUF_X2 port map( A => n22175, Z => n22200);
   U21977 : XNOR2_X1 port map( A => n21200, B => n20839, ZN => n20844);
   U21978 : XNOR2_X1 port map( A => n21998, B => n20840, ZN => n20841);
   U21979 : XNOR2_X1 port map( A => n20842, B => n20841, ZN => n20843);
   U21980 : XNOR2_X1 port map( A => n20844, B => n20843, ZN => n21759);
   U21981 : MUX2_X1 port map( A => n22197, B => n4360, S => n23571, Z => n20846
                           );
   U21982 : INV_X1 port map( A => n21222, ZN => n21536);
   U21984 : XNOR2_X1 port map( A => n20847, B => n21970, ZN => n20850);
   U21985 : XNOR2_X1 port map( A => n21224, B => n20848, ZN => n20849);
   U21987 : NOR2_X1 port map( A1 => n325, A2 => n22200, ZN => n20856);
   U21988 : XNOR2_X1 port map( A => n21743, B => n2477, ZN => n20851);
   U21989 : XNOR2_X1 port map( A => n20851, B => n25498, ZN => n20852);
   U21990 : XNOR2_X1 port map( A => n21208, B => n20852, ZN => n20855);
   U21991 : XNOR2_X1 port map( A => n21980, B => n21258, ZN => n20853);
   U21992 : XNOR2_X1 port map( A => n20853, B => n21981, ZN => n20854);
   U21993 : INV_X1 port map( A => n23619, ZN => n23637);
   U21994 : XNOR2_X1 port map( A => n1326, B => n887, ZN => n20857);
   U21995 : XNOR2_X1 port map( A => n21207, B => n20857, ZN => n20859);
   U21996 : XNOR2_X1 port map( A => n21501, B => n21258, ZN => n21615);
   U21997 : XNOR2_X1 port map( A => n21551, B => n21615, ZN => n20858);
   U21998 : XNOR2_X1 port map( A => n21492, B => n21567, ZN => n21326);
   U21999 : XNOR2_X1 port map( A => n21326, B => n20860, ZN => n20863);
   U22000 : XNOR2_X1 port map( A => n24996, B => n187, ZN => n20861);
   U22001 : XNOR2_X1 port map( A => n21216, B => n20861, ZN => n20862);
   U22003 : XNOR2_X1 port map( A => n21481, B => n20864, ZN => n20865);
   U22004 : XNOR2_X1 port map( A => n20865, B => n21633, ZN => n20866);
   U22005 : XNOR2_X1 port map( A => n20866, B => n21562, ZN => n20868);
   U22006 : XNOR2_X1 port map( A => n20868, B => n20867, ZN => n22889);
   U22008 : INV_X1 port map( A => n20870, ZN => n21471);
   U22009 : XNOR2_X1 port map( A => n21471, B => n21307, ZN => n20871);
   U22010 : XNOR2_X1 port map( A => n21191, B => n20871, ZN => n20880);
   U22011 : XNOR2_X1 port map( A => n21525, B => n25065, ZN => n20878);
   U22012 : NAND3_X1 port map( A1 => n20872, A2 => n23225, A3 => n20412, ZN => 
                           n20875);
   U22013 : NAND3_X1 port map( A1 => n20873, A2 => n1754, A3 => n20876, ZN => 
                           n20874);
   U22014 : OAI211_X1 port map( C1 => n1754, C2 => n20876, A => n20875, B => 
                           n20874, ZN => n20877);
   U22015 : XNOR2_X1 port map( A => n20878, B => n20877, ZN => n20879);
   U22017 : XNOR2_X1 port map( A => n21229, B => n20881, ZN => n20886);
   U22018 : XNOR2_X1 port map( A => n24485, B => n1768, ZN => n20884);
   U22019 : XNOR2_X1 port map( A => n21158, B => n21606, ZN => n20883);
   U22020 : XNOR2_X1 port map( A => n20884, B => n20883, ZN => n20885);
   U22021 : XNOR2_X1 port map( A => n21649, B => n23620, ZN => n20888);
   U22022 : XNOR2_X1 port map( A => n21579, B => n21728, ZN => n20887);
   U22023 : XNOR2_X1 port map( A => n20887, B => n20888, ZN => n20891);
   U22024 : XNOR2_X1 port map( A => n21198, B => n20889, ZN => n20890);
   U22025 : XNOR2_X1 port map( A => n20891, B => n20890, ZN => n22728);
   U22026 : NOR2_X1 port map( A1 => n22889, A2 => n25375, ZN => n20894);
   U22027 : INV_X1 port map( A => n23634, ZN => n20896);
   U22028 : INV_X1 port map( A => n21974, ZN => n20897);
   U22029 : XNOR2_X1 port map( A => n21550, B => n20897, ZN => n21747);
   U22030 : XNOR2_X1 port map( A => n21747, B => n20898, ZN => n20902);
   U22031 : XNOR2_X1 port map( A => n25498, B => n2745, ZN => n20900);
   U22032 : XNOR2_X1 port map( A => n20900, B => n20899, ZN => n20901);
   U22033 : XNOR2_X2 port map( A => n20902, B => n20901, ZN => n22159);
   U22034 : XNOR2_X1 port map( A => n21694, B => n21212, ZN => n20903);
   U22035 : XNOR2_X1 port map( A => n20904, B => n449, ZN => n20905);
   U22036 : XNOR2_X1 port map( A => n20905, B => n25222, ZN => n20907);
   U22037 : XNOR2_X1 port map( A => n21568, B => n21621, ZN => n20906);
   U22038 : XNOR2_X1 port map( A => n20907, B => n20906, ZN => n20908);
   U22039 : NOR2_X1 port map( A1 => n22159, A2 => n25485, ZN => n22212);
   U22040 : XNOR2_X1 port map( A => n21736, B => n2991, ZN => n20916);
   U22041 : XNOR2_X1 port map( A => n20914, B => n21532, ZN => n20915);
   U22042 : XNOR2_X1 port map( A => n20916, B => n20915, ZN => n20917);
   U22043 : XNOR2_X1 port map( A => n21699, B => n21704, ZN => n21129);
   U22044 : XNOR2_X1 port map( A => n20917, B => n21129, ZN => n20918);
   U22045 : XNOR2_X1 port map( A => n21971, B => n21967, ZN => n21538);
   U22046 : XNOR2_X1 port map( A => n21445, B => n21228, ZN => n21685);
   U22047 : XNOR2_X1 port map( A => n21686, B => n21141, ZN => n21543);
   U22048 : XNOR2_X1 port map( A => n21685, B => n21543, ZN => n20922);
   U22049 : XNOR2_X1 port map( A => n21591, B => n22739, ZN => n20920);
   U22050 : XNOR2_X1 port map( A => n22006, B => n21160, ZN => n20919);
   U22051 : XNOR2_X1 port map( A => n20920, B => n20919, ZN => n20921);
   U22052 : XNOR2_X1 port map( A => n20922, B => n20921, ZN => n22209);
   U22053 : XNOR2_X1 port map( A => n20948, B => n21678, ZN => n20923);
   U22054 : XNOR2_X1 port map( A => n21114, B => n20923, ZN => n20931);
   U22055 : INV_X1 port map( A => n21713, ZN => n20924);
   U22056 : XNOR2_X1 port map( A => n21599, B => n20924, ZN => n20929);
   U22057 : AOI21_X1 port map( B1 => n20927, B2 => n3115, A => n20926, ZN => 
                           n20928);
   U22058 : XNOR2_X1 port map( A => n20929, B => n20928, ZN => n20930);
   U22059 : AOI22_X1 port map( A1 => n22212, A2 => n2315, B1 => n20932, B2 => 
                           n25018, ZN => n20942);
   U22060 : XNOR2_X1 port map( A => n21992, B => n21670, ZN => n20934);
   U22061 : XNOR2_X1 port map( A => n21997, B => n21577, ZN => n20933);
   U22062 : XNOR2_X1 port map( A => n20934, B => n20933, ZN => n20939);
   U22063 : XNOR2_X1 port map( A => n21515, B => n21439, ZN => n20937);
   U22064 : INV_X1 port map( A => n2236, ZN => n20935);
   U22065 : XNOR2_X1 port map( A => n21647, B => n20935, ZN => n20936);
   U22066 : XNOR2_X1 port map( A => n20937, B => n20936, ZN => n20938);
   U22067 : XNOR2_X1 port map( A => n20939, B => n20938, ZN => n21766);
   U22068 : INV_X1 port map( A => n22205, ZN => n22156);
   U22069 : OAI21_X1 port map( B1 => n22064, B2 => n22156, A => n22159, ZN => 
                           n20940);
   U22071 : XNOR2_X1 port map( A => n21587, B => n21267, ZN => n20944);
   U22072 : XNOR2_X1 port map( A => n22005, B => n1815, ZN => n20943);
   U22073 : XNOR2_X1 port map( A => n20944, B => n20943, ZN => n20947);
   U22074 : XNOR2_X1 port map( A => n21142, B => n21541, ZN => n21612);
   U22075 : XNOR2_X1 port map( A => n21612, B => n20945, ZN => n20946);
   U22076 : XNOR2_X1 port map( A => n20946, B => n20947, ZN => n22916);
   U22077 : XNOR2_X1 port map( A => n21115, B => n20948, ZN => n20949);
   U22078 : XNOR2_X1 port map( A => n21096, B => n20949, ZN => n20953);
   U22079 : XNOR2_X1 port map( A => n22014, B => n24962, ZN => n20951);
   U22080 : XNOR2_X1 port map( A => n21311, B => n1746, ZN => n20950);
   U22081 : XNOR2_X1 port map( A => n20951, B => n20950, ZN => n20952);
   U22082 : XNOR2_X1 port map( A => n20953, B => n20952, ZN => n22070);
   U22083 : NOR2_X1 port map( A1 => n22916, A2 => n24902, ZN => n22116);
   U22084 : XNOR2_X1 port map( A => n21084, B => n21133, ZN => n20955);
   U22085 : XNOR2_X1 port map( A => n20954, B => n20955, ZN => n20959);
   U22086 : XNOR2_X1 port map( A => n21245, B => n2990, ZN => n20956);
   U22087 : XNOR2_X1 port map( A => n20957, B => n20956, ZN => n20958);
   U22088 : XNOR2_X1 port map( A => n21658, B => n21452, ZN => n21977);
   U22089 : XNOR2_X1 port map( A => n21136, B => n21505, ZN => n21614);
   U22090 : XNOR2_X1 port map( A => n21977, B => n21614, ZN => n20968);
   U22091 : XNOR2_X1 port map( A => n20964, B => n1804, ZN => n20965);
   U22092 : XNOR2_X1 port map( A => n20965, B => n21297, ZN => n20966);
   U22093 : XNOR2_X1 port map( A => n20966, B => n24898, ZN => n20967);
   U22094 : NAND2_X1 port map( A1 => n22918, A2 => n22072, ZN => n22115);
   U22095 : XNOR2_X1 port map( A => n25202, B => n21126, ZN => n20970);
   U22096 : XNOR2_X1 port map( A => n20970, B => n20969, ZN => n20974);
   U22097 : XNOR2_X1 port map( A => n20982, B => n2989, ZN => n20971);
   U22098 : XNOR2_X1 port map( A => n20972, B => n20971, ZN => n20973);
   U22100 : NAND2_X1 port map( A1 => n22917, A2 => n22072, ZN => n22169);
   U22101 : INV_X1 port map( A => n22115, ZN => n20980);
   U22102 : INV_X1 port map( A => Key(38), ZN => n20975);
   U22103 : XNOR2_X1 port map( A => n21996, B => n21514, ZN => n20976);
   U22104 : XNOR2_X1 port map( A => n21648, B => n20976, ZN => n20977);
   U22105 : NOR2_X1 port map( A1 => n22166, A2 => n22072, ZN => n20979);
   U22106 : AOI22_X1 port map( A1 => n20981, A2 => n23637, B1 => n23648, B2 => 
                           n23649, ZN => n21078);
   U22107 : XNOR2_X1 port map( A => n20983, B => n20982, ZN => n20985);
   U22108 : XNOR2_X1 port map( A => n20985, B => n20984, ZN => n20988);
   U22109 : INV_X1 port map( A => n21053, ZN => n20986);
   U22110 : XNOR2_X1 port map( A => n21534, B => n20986, ZN => n21706);
   U22111 : XNOR2_X1 port map( A => n21706, B => n21429, ZN => n20987);
   U22112 : XNOR2_X1 port map( A => n21070, B => n21399, ZN => n20989);
   U22113 : XNOR2_X1 port map( A => n20990, B => n20989, ZN => n20994);
   U22114 : XNOR2_X1 port map( A => n20992, B => n20991, ZN => n20993);
   U22116 : XNOR2_X1 port map( A => n21415, B => n21241, ZN => n20998);
   U22117 : INV_X1 port map( A => n20995, ZN => n23945);
   U22118 : XNOR2_X1 port map( A => n24899, B => n23945, ZN => n20996);
   U22119 : XNOR2_X1 port map( A => n21023, B => n20996, ZN => n20997);
   U22121 : XNOR2_X1 port map( A => n21182, B => n21510, ZN => n21669);
   U22122 : XNOR2_X1 port map( A => n21254, B => n21669, ZN => n21002);
   U22123 : XNOR2_X1 port map( A => n21334, B => n20999, ZN => n21392);
   U22124 : XNOR2_X1 port map( A => n21578, B => n3131, ZN => n21000);
   U22125 : XNOR2_X1 port map( A => n21392, B => n21000, ZN => n21001);
   U22126 : XNOR2_X1 port map( A => n21002, B => n21001, ZN => n22923);
   U22127 : INV_X1 port map( A => n22923, ZN => n22712);
   U22129 : XNOR2_X1 port map( A => n21409, B => n21003, ZN => n21007);
   U22130 : XNOR2_X1 port map( A => n21554, B => n3164, ZN => n21004);
   U22131 : XNOR2_X1 port map( A => n21005, B => n21004, ZN => n21006);
   U22132 : INV_X1 port map( A => n22927, ZN => n22188);
   U22133 : NAND2_X1 port map( A1 => n22926, A2 => n22188, ZN => n21020);
   U22134 : NAND2_X1 port map( A1 => n21009, A2 => n21008, ZN => n21011);
   U22135 : NAND2_X1 port map( A1 => n21011, A2 => n21010, ZN => n21012);
   U22136 : XNOR2_X1 port map( A => n21043, B => n21687, ZN => n21015);
   U22137 : XNOR2_X1 port map( A => n21267, B => n2241, ZN => n21014);
   U22138 : XNOR2_X1 port map( A => n21015, B => n21014, ZN => n21018);
   U22139 : XNOR2_X1 port map( A => n25400, B => n21266, ZN => n21016);
   U22140 : XNOR2_X1 port map( A => n21420, B => n21016, ZN => n21017);
   U22141 : XNOR2_X1 port map( A => n21017, B => n21018, ZN => n22922);
   U22142 : NAND2_X1 port map( A1 => n22923, A2 => n22922, ZN => n21019);
   U22143 : OAI21_X1 port map( B1 => n22926, B2 => n22927, A => n21019, ZN => 
                           n22711);
   U22144 : XNOR2_X1 port map( A => n25265, B => n21414, ZN => n21025);
   U22145 : XNOR2_X1 port map( A => n21025, B => n21600, ZN => n21243);
   U22147 : XNOR2_X1 port map( A => n21027, B => n2882, ZN => n21028);
   U22148 : XNOR2_X1 port map( A => n21028, B => n20475, ZN => n21029);
   U22149 : OAI21_X1 port map( B1 => n21033, B2 => n24378, A => n21031, ZN => 
                           n21037);
   U22150 : AOI21_X1 port map( B1 => n21035, B2 => n21034, A => n21038, ZN => 
                           n21036);
   U22151 : AOI21_X1 port map( B1 => n21038, B2 => n21037, A => n21036, ZN => 
                           n21039);
   U22152 : XNOR2_X1 port map( A => n21041, B => n21040, ZN => n21748);
   U22153 : INV_X1 port map( A => n22245, ZN => n22240);
   U22154 : XNOR2_X1 port map( A => n22007, B => n21750, ZN => n21044);
   U22155 : XNOR2_X1 port map( A => n21043, B => n21042, ZN => n21589);
   U22156 : XNOR2_X1 port map( A => n21044, B => n21589, ZN => n21050);
   U22157 : XNOR2_X1 port map( A => n24485, B => n21045, ZN => n21048);
   U22158 : XNOR2_X1 port map( A => n21422, B => n21046, ZN => n21047);
   U22159 : XNOR2_X1 port map( A => n21048, B => n21047, ZN => n21049);
   U22160 : XNOR2_X1 port map( A => n21050, B => n21049, ZN => n22239);
   U22161 : INV_X1 port map( A => n22239, ZN => n22181);
   U22162 : XNOR2_X1 port map( A => n21477, B => n21735, ZN => n21052);
   U22163 : XNOR2_X1 port map( A => n21734, B => n3093, ZN => n21051);
   U22164 : XNOR2_X1 port map( A => n21052, B => n21051, ZN => n21057);
   U22165 : XNOR2_X1 port map( A => n24353, B => n21053, ZN => n21055);
   U22166 : INV_X1 port map( A => n21319, ZN => n21054);
   U22167 : XNOR2_X1 port map( A => n21055, B => n21564, ZN => n21056);
   U22168 : OAI22_X1 port map( A1 => n22243, A2 => n22240, B1 => n22181, B2 => 
                           n22244, ZN => n21077);
   U22169 : XNOR2_X1 port map( A => n21058, B => n21182, ZN => n21060);
   U22170 : INV_X1 port map( A => n21336, ZN => n21059);
   U22171 : XNOR2_X1 port map( A => n21059, B => n21436, ZN => n21726);
   U22172 : XNOR2_X1 port map( A => n21726, B => n21060, ZN => n21064);
   U22173 : XNOR2_X1 port map( A => n24100, B => n2137, ZN => n21062);
   U22174 : XNOR2_X1 port map( A => n21061, B => n21062, ZN => n21063);
   U22175 : XNOR2_X1 port map( A => n21064, B => n21063, ZN => n22242);
   U22176 : INV_X1 port map( A => n22242, ZN => n22180);
   U22179 : XNOR2_X1 port map( A => n21071, B => n21070, ZN => n21574);
   U22180 : XNOR2_X1 port map( A => n21574, B => n21246, ZN => n21075);
   U22181 : XNOR2_X1 port map( A => n21087, B => n21720, ZN => n21073);
   U22182 : XNOR2_X1 port map( A => n21693, B => n836, ZN => n21072);
   U22183 : XNOR2_X1 port map( A => n21073, B => n21072, ZN => n21074);
   U22184 : XNOR2_X1 port map( A => n21074, B => n21075, ZN => n22059);
   U22186 : XNOR2_X1 port map( A => n25202, B => n21630, ZN => n21080);
   U22187 : XNOR2_X1 port map( A => n21477, B => n2318, ZN => n21081);
   U22189 : XNOR2_X1 port map( A => n25073, B => n21084, ZN => n21086);
   U22190 : XNOR2_X1 port map( A => n25040, B => n21324, ZN => n21085);
   U22191 : XNOR2_X1 port map( A => n21086, B => n21085, ZN => n21090);
   U22192 : XNOR2_X1 port map( A => n21087, B => n1952, ZN => n21088);
   U22193 : XNOR2_X1 port map( A => n21496, B => n21088, ZN => n21089);
   U22194 : INV_X1 port map( A => n21157, ZN => n21091);
   U22195 : XNOR2_X1 port map( A => n21091, B => n3125, ZN => n21092);
   U22196 : XNOR2_X1 port map( A => n21612, B => n21093, ZN => n21094);
   U22198 : INV_X1 port map( A => n23998, ZN => n22373);
   U22199 : XNOR2_X1 port map( A => n22012, B => n21096, ZN => n21100);
   U22200 : XNOR2_X1 port map( A => n21310, B => n21115, ZN => n21098);
   U22201 : XNOR2_X1 port map( A => n24899, B => n2739, ZN => n21097);
   U22202 : XNOR2_X1 port map( A => n21098, B => n21097, ZN => n21099);
   U22204 : XNOR2_X1 port map( A => n21172, B => n21980, ZN => n21101);
   U22205 : XNOR2_X1 port map( A => n24898, B => n21101, ZN => n21105);
   U22206 : XNOR2_X1 port map( A => n21974, B => n763, ZN => n21102);
   U22207 : XNOR2_X1 port map( A => n21102, B => n21660, ZN => n21103);
   U22208 : XNOR2_X1 port map( A => n21614, B => n21103, ZN => n21104);
   U22209 : XNOR2_X1 port map( A => n21107, B => n21334, ZN => n21109);
   U22210 : XNOR2_X1 port map( A => n21108, B => n21109, ZN => n21111);
   U22211 : AND2_X1 port map( A1 => n24439, A2 => n25414, ZN => n21112);
   U22212 : INV_X1 port map( A => n23997, ZN => n21855);
   U22213 : OAI21_X1 port map( B1 => n22676, B2 => n21112, A => n21855, ZN => 
                           n21113);
   U22214 : XNOR2_X1 port map( A => n21114, B => n21716, ZN => n21119);
   U22215 : XNOR2_X1 port map( A => n21115, B => Key(172), ZN => n21117);
   U22216 : XNOR2_X1 port map( A => n21116, B => n21117, ZN => n21118);
   U22217 : XNOR2_X1 port map( A => n21119, B => n21118, ZN => n22667);
   U22218 : XNOR2_X1 port map( A => n21439, B => n23699, ZN => n21120);
   U22219 : XNOR2_X1 port map( A => n21120, B => n21728, ZN => n21122);
   U22220 : XNOR2_X1 port map( A => n21122, B => n21121, ZN => n21125);
   U22221 : XNOR2_X1 port map( A => n21336, B => n25091, ZN => n21123);
   U22222 : XNOR2_X1 port map( A => n21648, B => n21123, ZN => n21124);
   U22224 : OR2_X1 port map( A1 => n22667, A2 => n25023, ZN => n21147);
   U22225 : XNOR2_X1 port map( A => n21127, B => n21126, ZN => n21128);
   U22226 : XNOR2_X1 port map( A => n21739, B => n21128, ZN => n21131);
   U22227 : XNOR2_X1 port map( A => n21971, B => n21129, ZN => n21130);
   U22229 : XNOR2_X1 port map( A => n21132, B => n1726, ZN => n21134);
   U22231 : XNOR2_X1 port map( A => n21136, B => n21506, ZN => n21137);
   U22232 : XNOR2_X1 port map( A => n21452, B => n21300, ZN => n21556);
   U22233 : XNOR2_X1 port map( A => n21556, B => n21137, ZN => n21139);
   U22234 : OAI21_X1 port map( B1 => n21147, B2 => n22675, A => n22365, ZN => 
                           n21149);
   U22235 : XNOR2_X1 port map( A => n21587, B => n21141, ZN => n22003);
   U22236 : XNOR2_X1 port map( A => n21685, B => n22003, ZN => n21145);
   U22237 : XNOR2_X1 port map( A => n21142, B => n1739, ZN => n21143);
   U22238 : XNOR2_X1 port map( A => n21755, B => n21143, ZN => n21144);
   U22239 : XNOR2_X1 port map( A => n21145, B => n21144, ZN => n22670);
   U22240 : INV_X1 port map( A => n22670, ZN => n22784);
   U22241 : OAI22_X1 port map( A1 => n21147, A2 => n25462, B1 => n22784, B2 => 
                           n21146, ZN => n21148);
   U22242 : NAND2_X1 port map( A1 => n23074, A2 => n25452, ZN => n21239);
   U22243 : NOR3_X1 port map( A1 => n22462, A2 => n24367, A3 => n25450, ZN => 
                           n21150);
   U22244 : NAND2_X1 port map( A1 => n21375, A2 => n22459, ZN => n21930);
   U22246 : XNOR2_X1 port map( A => n21525, B => n173, ZN => n21152);
   U22247 : XNOR2_X1 port map( A => n21152, B => n21679, ZN => n21154);
   U22248 : XNOR2_X1 port map( A => n21154, B => n21153, ZN => n21155);
   U22249 : XNOR2_X1 port map( A => n21689, B => n21606, ZN => n21159);
   U22250 : XNOR2_X1 port map( A => n21157, B => n21158, ZN => n21342);
   U22251 : XNOR2_X1 port map( A => n21342, B => n21159, ZN => n21165);
   U22252 : INV_X1 port map( A => n1767, ZN => n21161);
   U22253 : XNOR2_X1 port map( A => n21687, B => n21161, ZN => n21162);
   U22254 : XNOR2_X1 port map( A => n21163, B => n21162, ZN => n21164);
   U22255 : XNOR2_X1 port map( A => n21084, B => n21720, ZN => n21166);
   U22256 : XNOR2_X1 port map( A => n21326, B => n21166, ZN => n21168);
   U22257 : INV_X1 port map( A => n3084, ZN => n23045);
   U22258 : XNOR2_X1 port map( A => n21501, B => n21169, ZN => n21170);
   U22259 : XNOR2_X1 port map( A => n21170, B => n24491, ZN => n21171);
   U22260 : XNOR2_X1 port map( A => n21171, B => n21618, ZN => n21175);
   U22261 : XNOR2_X1 port map( A => n21173, B => n21172, ZN => n21298);
   U22262 : XNOR2_X1 port map( A => n21298, B => n24898, ZN => n21174);
   U22263 : NOR2_X1 port map( A1 => n24042, A2 => n274, ZN => n21181);
   U22264 : XNOR2_X1 port map( A => n25202, B => n24896, ZN => n21177);
   U22265 : XNOR2_X1 port map( A => n25495, B => n21177, ZN => n21180);
   U22266 : XNOR2_X1 port map( A => n21735, B => n1869, ZN => n21178);
   U22267 : XNOR2_X1 port map( A => n21635, B => n21178, ZN => n21179);
   U22268 : AOI22_X1 port map( A1 => n21923, A2 => n274, B1 => n21181, B2 => 
                           n22448, ZN => n21190);
   U22269 : XNOR2_X1 port map( A => n21182, B => n21511, ZN => n21646);
   U22270 : XNOR2_X1 port map( A => n21436, B => n21579, ZN => n21183);
   U22271 : XNOR2_X1 port map( A => n21646, B => n21183, ZN => n21187);
   U22272 : XNOR2_X1 port map( A => n21334, B => n3183, ZN => n21185);
   U22273 : XNOR2_X1 port map( A => n21184, B => n21185, ZN => n21186);
   U22274 : XNOR2_X1 port map( A => n21191, B => n21192, ZN => n21197);
   U22275 : XNOR2_X1 port map( A => n21596, B => n21678, ZN => n21195);
   U22276 : XNOR2_X1 port map( A => n21193, B => n1797, ZN => n21194);
   U22277 : XNOR2_X1 port map( A => n21195, B => n21194, ZN => n21196);
   U22278 : XNOR2_X1 port map( A => n21199, B => n21198, ZN => n21203);
   U22279 : XNOR2_X1 port map( A => n21670, B => n3152, ZN => n21201);
   U22280 : XNOR2_X1 port map( A => n21200, B => n21201, ZN => n21202);
   U22282 : XNOR2_X1 port map( A => n24305, B => n21204, ZN => n21206);
   U22283 : XNOR2_X1 port map( A => n21207, B => n21206, ZN => n21211);
   U22284 : XNOR2_X2 port map( A => n21210, B => n21211, ZN => n22804);
   U22285 : INV_X1 port map( A => n21212, ZN => n21213);
   U22286 : XNOR2_X1 port map( A => n21213, B => n1364, ZN => n21214);
   U22287 : XNOR2_X1 port map( A => n21215, B => n21214, ZN => n21219);
   U22288 : XNOR2_X1 port map( A => n21217, B => n21216, ZN => n21218);
   U22290 : MUX2_X1 port map( A => n22798, B => n22804, S => n24559, Z => 
                           n21238);
   U22291 : XNOR2_X1 port map( A => n24434, B => n2881, ZN => n21220);
   U22292 : XNOR2_X1 port map( A => n21221, B => n21220, ZN => n21226);
   U22293 : XNOR2_X1 port map( A => n21318, B => n21222, ZN => n21223);
   U22294 : XNOR2_X1 port map( A => n21224, B => n21223, ZN => n21225);
   U22295 : XNOR2_X2 port map( A => n21225, B => n21226, ZN => n22800);
   U22296 : NOR2_X1 port map( A1 => n22804, A2 => n22800, ZN => n22583);
   U22297 : XNOR2_X1 port map( A => n21227, B => n21228, ZN => n21230);
   U22298 : XNOR2_X1 port map( A => n21229, B => n21230, ZN => n21235);
   U22299 : XNOR2_X1 port map( A => n21591, B => n923, ZN => n21232);
   U22300 : XNOR2_X1 port map( A => n21233, B => n21232, ZN => n21234);
   U22302 : INV_X1 port map( A => n22805, ZN => n21236);
   U22303 : NOR2_X1 port map( A1 => n21236, A2 => n22803, ZN => n21237);
   U22304 : INV_X1 port map( A => n24561, ZN => n22799);
   U22305 : XNOR2_X1 port map( A => n21640, B => n2970, ZN => n21240);
   U22306 : XNOR2_X1 port map( A => n21240, B => n21520, ZN => n21242);
   U22307 : XNOR2_X1 port map( A => n21241, B => n21242, ZN => n21244);
   U22308 : XNOR2_X1 port map( A => n21245, B => n21622, ZN => n21403);
   U22309 : XNOR2_X1 port map( A => n21246, B => n21403, ZN => n21251);
   U22310 : XNOR2_X1 port map( A => n21495, B => n1924, ZN => n21249);
   U22311 : XOR2_X1 port map( A => n21720, B => n21247, Z => n21248);
   U22312 : XNOR2_X1 port map( A => n21249, B => n21248, ZN => n21250);
   U22313 : XNOR2_X1 port map( A => n21251, B => n21250, ZN => n21265);
   U22314 : XNOR2_X1 port map( A => n21253, B => n21252, ZN => n21257);
   U22315 : XNOR2_X1 port map( A => n1381, B => n2005, ZN => n21255);
   U22316 : XNOR2_X1 port map( A => n21254, B => n21255, ZN => n21256);
   U22317 : XNOR2_X1 port map( A => n21297, B => n21258, ZN => n21408);
   U22318 : XNOR2_X1 port map( A => n21260, B => n21259, ZN => n21261);
   U22319 : XNOR2_X1 port map( A => n21261, B => n21408, ZN => n21264);
   U22320 : XNOR2_X1 port map( A => n21262, B => n21981, ZN => n21263);
   U22321 : XNOR2_X1 port map( A => n21264, B => n21263, ZN => n22619);
   U22323 : INV_X1 port map( A => n22792, ZN => n22313);
   U22324 : INV_X1 port map( A => n21265, ZN => n22612);
   U22325 : XNOR2_X1 port map( A => n21750, B => n21266, ZN => n21268);
   U22326 : XNOR2_X1 port map( A => n21608, B => n21267, ZN => n21421);
   U22327 : XNOR2_X1 port map( A => n21421, B => n21268, ZN => n21272);
   U22328 : XNOR2_X1 port map( A => n21422, B => n1810, ZN => n21269);
   U22329 : XNOR2_X1 port map( A => n21270, B => n21269, ZN => n21271);
   U22330 : XNOR2_X1 port map( A => n21272, B => n21271, ZN => n22791);
   U22331 : NAND3_X1 port map( A1 => n22313, A2 => n22612, A3 => n22791, ZN => 
                           n21279);
   U22332 : NAND2_X1 port map( A1 => n22619, A2 => n22614, ZN => n21370);
   U22333 : XNOR2_X1 port map( A => n24353, B => n21273, ZN => n21274);
   U22334 : XNOR2_X1 port map( A => n21430, B => n21274, ZN => n21278);
   U22335 : XNOR2_X1 port map( A => n21536, B => n21735, ZN => n21276);
   U22336 : XNOR2_X1 port map( A => n21734, B => n2743, ZN => n21275);
   U22337 : XNOR2_X1 port map( A => n21276, B => n21275, ZN => n21277);
   U22338 : XNOR2_X1 port map( A => n21278, B => n21277, ZN => n22615);
   U22341 : NAND2_X1 port map( A1 => n21282, A2 => n21281, ZN => n21284);
   U22342 : INV_X1 port map( A => n1789, ZN => n21283);
   U22343 : XNOR2_X1 port map( A => n21284, B => n21283, ZN => Ciphertext(10));
   U22344 : AND2_X1 port map( A1 => n23217, A2 => n23228, ZN => n21285);
   U22345 : AOI22_X1 port map( A1 => n23215, A2 => n23219, B1 => n21285, B2 => 
                           n1340, ZN => n21286);
   U22346 : INV_X1 port map( A => n21742, ZN => n21287);
   U22347 : XNOR2_X1 port map( A => n21288, B => n21287, ZN => Ciphertext(39));
   U22348 : INV_X1 port map( A => n21816, ZN => n22687);
   U22349 : NOR2_X1 port map( A1 => n22685, A2 => n22689, ZN => n21290);
   U22350 : OAI21_X1 port map( B1 => n21856, B2 => n22774, A => n21292, ZN => 
                           n21293);
   U22351 : INV_X1 port map( A => n22679, ZN => n22771);
   U22352 : NAND2_X1 port map( A1 => n21856, A2 => n22770, ZN => n22682);
   U22353 : OR2_X1 port map( A1 => n22682, A2 => n22370, ZN => n21294);
   U22355 : INV_X1 port map( A => n21841, ZN => n21840);
   U22356 : NOR2_X1 port map( A1 => n23828, A2 => n891, ZN => n21351);
   U22357 : XNOR2_X1 port map( A => n21297, B => n1870, ZN => n21299);
   U22358 : XNOR2_X1 port map( A => n21299, B => n21298, ZN => n21305);
   U22359 : XNOR2_X1 port map( A => n21301, B => n21300, ZN => n21303);
   U22360 : XNOR2_X1 port map( A => n21303, B => n21302, ZN => n21304);
   U22362 : INV_X1 port map( A => n22220, ZN => n22216);
   U22363 : XNOR2_X1 port map( A => n21306, B => n21307, ZN => n21598);
   U22364 : XNOR2_X1 port map( A => n21308, B => n21598, ZN => n21315);
   U22365 : XNOR2_X1 port map( A => n21310, B => n21309, ZN => n21313);
   U22366 : XNOR2_X1 port map( A => n21311, B => n25062, ZN => n21416);
   U22367 : XNOR2_X1 port map( A => n21416, B => n21313, ZN => n21314);
   U22368 : XNOR2_X1 port map( A => n21317, B => n21316, ZN => n21323);
   U22369 : XNOR2_X1 port map( A => n21318, B => n21965, ZN => n21321);
   U22370 : XNOR2_X1 port map( A => n21319, B => n2782, ZN => n21320);
   U22371 : XNOR2_X1 port map( A => n21321, B => n21320, ZN => n21322);
   U22373 : MUX2_X1 port map( A => n22216, B => n22222, S => n22214, Z => 
                           n21347);
   U22374 : XNOR2_X1 port map( A => n21325, B => n21324, ZN => n21400);
   U22375 : XNOR2_X1 port map( A => n21400, B => n21326, ZN => n21330);
   U22376 : XNOR2_X1 port map( A => n21985, B => n2761, ZN => n21327);
   U22377 : XNOR2_X1 port map( A => n21328, B => n21327, ZN => n21329);
   U22378 : XNOR2_X1 port map( A => n21332, B => n21331, ZN => n21395);
   U22379 : XNOR2_X1 port map( A => n21395, B => n21333, ZN => n21340);
   U22380 : XNOR2_X1 port map( A => n21579, B => n21334, ZN => n21338);
   U22381 : INV_X1 port map( A => n21335, ZN => n23961);
   U22382 : XNOR2_X1 port map( A => n21336, B => n23961, ZN => n21337);
   U22383 : XNOR2_X1 port map( A => n21338, B => n21337, ZN => n21339);
   U22384 : XNOR2_X1 port map( A => n21340, B => n21339, ZN => n22219);
   U22385 : NAND2_X1 port map( A1 => n22222, A2 => n22219, ZN => n21341);
   U22386 : INV_X1 port map( A => n1951, ZN => n23663);
   U22387 : OAI21_X2 port map( B1 => n21347, B2 => n2817, A => n21346, ZN => 
                           n23827);
   U22388 : AND2_X1 port map( A1 => n23827, A2 => n891, ZN => n21361);
   U22389 : INV_X1 port map( A => n21361, ZN => n21350);
   U22390 : INV_X1 port map( A => n23828, ZN => n23834);
   U22391 : NAND2_X1 port map( A1 => n23834, A2 => n891, ZN => n21362);
   U22392 : AOI22_X1 port map( A1 => n22231, A2 => n24905, B1 => n22226, B2 => 
                           n22225, ZN => n22058);
   U22393 : NOR2_X1 port map( A1 => n22058, A2 => n21794, ZN => n21354);
   U22394 : AOI211_X1 port map( C1 => n3231, C2 => n22228, A => n22226, B => 
                           n22056, ZN => n21353);
   U22395 : INV_X1 port map( A => n23817, ZN => n23811);
   U22397 : OAI22_X1 port map( A1 => n21355, A2 => n23827, B1 => n23811, B2 => 
                           n21359, ZN => n21356);
   U22398 : NAND2_X1 port map( A1 => n23810, A2 => n23827, ZN => n21358);
   U22399 : NAND2_X1 port map( A1 => n21358, A2 => n24972, ZN => n23034);
   U22400 : INV_X1 port map( A => n23034, ZN => n21360);
   U22401 : NAND3_X1 port map( A1 => n21360, A2 => n21359, A3 => n23827, ZN => 
                           n21366);
   U22402 : NAND2_X1 port map( A1 => n21364, A2 => n23034, ZN => n21365);
   U22403 : INV_X1 port map( A => n22138, ZN => n22334);
   U22404 : OAI21_X1 port map( B1 => n22337, B2 => n22334, A => n21368, ZN => 
                           n21367);
   U22406 : INV_X1 port map( A => n22137, ZN => n22274);
   U22407 : INV_X1 port map( A => n22791, ZN => n22617);
   U22408 : NOR2_X1 port map( A1 => n22789, A2 => n22614, ZN => n21374);
   U22409 : INV_X1 port map( A => n21370, ZN => n21373);
   U22410 : INV_X1 port map( A => n22615, ZN => n22790);
   U22411 : OAI211_X1 port map( C1 => n22614, C2 => n22790, A => n22313, B => 
                           n21371, ZN => n21372);
   U22413 : INV_X1 port map( A => n23153, ZN => n23138);
   U22414 : NOR2_X1 port map( A1 => n1363, A2 => n21375, ZN => n22328);
   U22415 : AND2_X1 port map( A1 => n21375, A2 => n22464, ZN => n21376);
   U22416 : INV_X1 port map( A => n22592, ZN => n21921);
   U22417 : MUX2_X1 port map( A => n21921, B => n2393, S => n25066, Z => n21378
                           );
   U22418 : INV_X1 port map( A => n23129, ZN => n23146);
   U22419 : INV_X1 port map( A => n21380, ZN => n21918);
   U22420 : INV_X1 port map( A => n22453, ZN => n21382);
   U22421 : NOR2_X1 port map( A1 => n22455, A2 => n1352, ZN => n21381);
   U22422 : AOI21_X1 port map( B1 => n21382, B2 => n22455, A => n21381, ZN => 
                           n21385);
   U22423 : INV_X1 port map( A => n24311, ZN => n21383);
   U22424 : NOR2_X1 port map( A1 => n22456, A2 => n21383, ZN => n21384);
   U22425 : AND2_X1 port map( A1 => n22799, A2 => n22803, ZN => n22806);
   U22426 : INV_X1 port map( A => n22800, ZN => n21386);
   U22427 : AOI22_X1 port map( A1 => n22806, A2 => n21386, B1 => n22803, B2 => 
                           n24992, ZN => n21390);
   U22431 : INV_X1 port map( A => n2033, ZN => n21391);
   U22432 : XNOR2_X1 port map( A => n24472, B => n2746, ZN => n21393);
   U22433 : XNOR2_X1 port map( A => n21392, B => n21393, ZN => n21397);
   U22434 : XNOR2_X1 port map( A => n24100, B => n21577, ZN => n21727);
   U22435 : XNOR2_X1 port map( A => n21395, B => n21727, ZN => n21396);
   U22436 : INV_X1 port map( A => n23334, ZN => n21413);
   U22437 : XNOR2_X1 port map( A => n21399, B => n21398, ZN => n21401);
   U22438 : XNOR2_X1 port map( A => n21400, B => n21401, ZN => n21405);
   U22439 : XNOR2_X1 port map( A => n25377, B => n21568, ZN => n21723);
   U22440 : XNOR2_X1 port map( A => n21723, B => n21403, ZN => n21404);
   U22441 : XNOR2_X1 port map( A => n21550, B => n2039, ZN => n21407);
   U22442 : XNOR2_X1 port map( A => n21407, B => n21406, ZN => n21411);
   U22443 : XNOR2_X1 port map( A => n21409, B => n21408, ZN => n21410);
   U22446 : XNOR2_X1 port map( A => n21599, B => n21414, ZN => n21717);
   U22447 : XNOR2_X1 port map( A => n21415, B => n21717, ZN => n21419);
   U22448 : XNOR2_X1 port map( A => n25065, B => n22635, ZN => n21417);
   U22449 : XNOR2_X1 port map( A => n21417, B => n21416, ZN => n21418);
   U22450 : INV_X1 port map( A => n24342, ZN => n22501);
   U22451 : XNOR2_X1 port map( A => n21420, B => n21421, ZN => n21426);
   U22452 : XNOR2_X1 port map( A => n21591, B => n21422, ZN => n21754);
   U22453 : INV_X1 port map( A => n21423, ZN => n22525);
   U22454 : XNOR2_X1 port map( A => n21754, B => n21424, ZN => n21425);
   U22456 : INV_X1 port map( A => n23336, ZN => n22499);
   U22457 : OAI21_X1 port map( B1 => n22855, B2 => n21428, A => n21427, ZN => 
                           n22431);
   U22458 : XNOR2_X1 port map( A => n21430, B => n21429, ZN => n21435);
   U22459 : XNOR2_X1 port map( A => n21433, B => n21432, ZN => n21434);
   U22460 : XNOR2_X1 port map( A => n21434, B => n21435, ZN => n22852);
   U22461 : NAND2_X1 port map( A1 => n22852, A2 => n22932, ZN => n22498);
   U22462 : NOR2_X1 port map( A1 => n24309, A2 => n22498, ZN => n22432);
   U22464 : XNOR2_X1 port map( A => n21436, B => n21510, ZN => n21438);
   U22465 : XNOR2_X1 port map( A => n21728, B => n21998, ZN => n21437);
   U22466 : XNOR2_X1 port map( A => n21437, B => n21438, ZN => n21443);
   U22467 : XNOR2_X1 port map( A => n21583, B => n25387, ZN => n21441);
   U22468 : XNOR2_X1 port map( A => n21729, B => n21942, ZN => n21440);
   U22469 : XNOR2_X1 port map( A => n21441, B => n21440, ZN => n21442);
   U22470 : XNOR2_X1 port map( A => n25400, B => n21445, ZN => n21447);
   U22471 : XNOR2_X1 port map( A => n21750, B => n2826, ZN => n21446);
   U22472 : XNOR2_X1 port map( A => n21447, B => n21446, ZN => n21451);
   U22473 : XNOR2_X1 port map( A => n21449, B => n21448, ZN => n21450);
   U22474 : XNOR2_X1 port map( A => n21452, B => n21660, ZN => n21453);
   U22475 : XNOR2_X1 port map( A => n21454, B => n21453, ZN => n21459);
   U22476 : XNOR2_X1 port map( A => n24491, B => n1724, ZN => n21456);
   U22477 : XNOR2_X1 port map( A => n21457, B => n21456, ZN => n21458);
   U22478 : XNOR2_X1 port map( A => n21459, B => n21458, ZN => n22128);
   U22479 : XNOR2_X1 port map( A => n21461, B => n21460, ZN => n21465);
   U22480 : XNOR2_X1 port map( A => n21463, B => n21462, ZN => n21464);
   U22481 : XNOR2_X1 port map( A => n21465, B => n21464, ZN => n21467);
   U22482 : NAND2_X1 port map( A1 => n22128, A2 => n21467, ZN => n21466);
   U22483 : OAI21_X1 port map( B1 => n22965, B2 => n22962, A => n21466, ZN => 
                           n22131);
   U22484 : INV_X1 port map( A => n22131, ZN => n21490);
   U22485 : INV_X1 port map( A => n21466, ZN => n21468);
   U22486 : NOR2_X1 port map( A1 => n21468, A2 => n22969, ZN => n21489);
   U22487 : XNOR2_X1 port map( A => n21676, B => n21469, ZN => n21470);
   U22488 : XNOR2_X1 port map( A => n21715, B => n21470, ZN => n21475);
   U22489 : XNOR2_X1 port map( A => n24962, B => n4233, ZN => n21473);
   U22490 : XNOR2_X1 port map( A => n21471, B => n24899, ZN => n21472);
   U22491 : XNOR2_X1 port map( A => n21472, B => n21473, ZN => n21474);
   U22492 : INV_X1 port map( A => n21959, ZN => n21487);
   U22493 : XNOR2_X1 port map( A => n21479, B => n21480, ZN => n21485);
   U22494 : XNOR2_X1 port map( A => n21534, B => n21559, ZN => n21483);
   U22495 : XNOR2_X1 port map( A => n21481, B => n2031, ZN => n21482);
   U22496 : XNOR2_X1 port map( A => n21483, B => n21482, ZN => n21484);
   U22498 : NAND2_X1 port map( A1 => n21487, A2 => n21486, ZN => n21488);
   U22499 : INV_X1 port map( A => n23369, ZN => n22741);
   U22500 : OR2_X1 port map( A1 => n24515, A2 => n22741, ZN => n21954);
   U22501 : XNOR2_X1 port map( A => n25470, B => n25073, ZN => n21627);
   U22502 : XNOR2_X1 port map( A => n21494, B => n21627, ZN => n21499);
   U22503 : XNOR2_X1 port map( A => n21495, B => n23072, ZN => n21497);
   U22504 : XNOR2_X1 port map( A => n21496, B => n21497, ZN => n21498);
   U22505 : XNOR2_X1 port map( A => n21498, B => n21499, ZN => n21540);
   U22506 : INV_X1 port map( A => n21540, ZN => n22947);
   U22507 : XNOR2_X1 port map( A => n21974, B => n21502, ZN => n21504);
   U22508 : XNOR2_X1 port map( A => n21503, B => n21504, ZN => n21509);
   U22509 : XNOR2_X1 port map( A => n21506, B => n21505, ZN => n21507);
   U22510 : XNOR2_X1 port map( A => n21981, B => n21507, ZN => n21508);
   U22511 : XNOR2_X1 port map( A => n21509, B => n21508, ZN => n21872);
   U22512 : INV_X1 port map( A => n21872, ZN => n22282);
   U22513 : XNOR2_X1 port map( A => n21510, B => n1381, ZN => n21513);
   U22514 : XNOR2_X1 port map( A => n21992, B => n21511, ZN => n21512);
   U22515 : XNOR2_X1 port map( A => n21512, B => n21513, ZN => n21519);
   U22517 : XNOR2_X1 port map( A => n21514, B => n24624, ZN => n21517);
   U22518 : XNOR2_X1 port map( A => n25091, B => n21515, ZN => n21516);
   U22519 : XNOR2_X1 port map( A => n21517, B => n21516, ZN => n21518);
   U22520 : INV_X1 port map( A => n22946, ZN => n21530);
   U22521 : XNOR2_X1 port map( A => n21521, B => n21520, ZN => n22013);
   U22522 : XNOR2_X1 port map( A => n21523, B => n21522, ZN => n21524);
   U22523 : XNOR2_X1 port map( A => n22013, B => n21524, ZN => n21529);
   U22524 : XNOR2_X1 port map( A => n21525, B => n853, ZN => n21527);
   U22525 : XNOR2_X1 port map( A => n21713, B => n21639, ZN => n21526);
   U22526 : XNOR2_X1 port map( A => n21527, B => n21526, ZN => n21528);
   U22527 : XNOR2_X1 port map( A => n21532, B => n21630, ZN => n21535);
   U22528 : XNOR2_X1 port map( A => n21536, B => n21633, ZN => n21537);
   U22529 : XNOR2_X1 port map( A => n21539, B => n21538, ZN => n22948);
   U22530 : INV_X1 port map( A => n22948, ZN => n22424);
   U22531 : XNOR2_X1 port map( A => n21541, B => n21606, ZN => n21542);
   U22532 : XNOR2_X1 port map( A => n21544, B => n21543, ZN => n21545);
   U22533 : OAI21_X1 port map( B1 => n22948, B2 => n21548, A => n21547, ZN => 
                           n22435);
   U22534 : INV_X1 port map( A => n22435, ZN => n21549);
   U22535 : XNOR2_X1 port map( A => n21550, B => n21975, ZN => n21552);
   U22536 : XNOR2_X1 port map( A => n21551, B => n21552, ZN => n21558);
   U22537 : INV_X1 port map( A => n21553, ZN => n23589);
   U22538 : XNOR2_X1 port map( A => n21554, B => n23589, ZN => n21555);
   U22539 : XNOR2_X1 port map( A => n21556, B => n21555, ZN => n21557);
   U22542 : XNOR2_X1 port map( A => n21561, B => n24306, ZN => n21963);
   U22543 : XNOR2_X1 port map( A => n21562, B => n21963, ZN => n21566);
   U22544 : XNOR2_X1 port map( A => n24434, B => n1856, ZN => n21563);
   U22545 : XNOR2_X1 port map( A => n21564, B => n21563, ZN => n21565);
   U22546 : XNOR2_X1 port map( A => n21568, B => n25385, ZN => n21571);
   U22547 : XNOR2_X1 port map( A => n24996, B => n2211, ZN => n21570);
   U22548 : XNOR2_X1 port map( A => n21571, B => n21570, ZN => n21576);
   U22549 : XNOR2_X1 port map( A => n21572, B => n21573, ZN => n21989);
   U22550 : XNOR2_X1 port map( A => n21989, B => n21574, ZN => n21575);
   U22551 : XNOR2_X1 port map( A => n21575, B => n21576, ZN => n22953);
   U22553 : XNOR2_X1 port map( A => n21577, B => n22385, ZN => n21581);
   U22554 : XNOR2_X1 port map( A => n21579, B => n21578, ZN => n21580);
   U22555 : XNOR2_X1 port map( A => n21580, B => n21581, ZN => n21586);
   U22556 : XNOR2_X1 port map( A => n21582, B => n21583, ZN => n21993);
   U22557 : XNOR2_X1 port map( A => n21993, B => n21584, ZN => n21585);
   U22558 : XNOR2_X1 port map( A => n21586, B => n21585, ZN => n22952);
   U22559 : XNOR2_X1 port map( A => n21588, B => n21587, ZN => n21590);
   U22560 : XNOR2_X1 port map( A => n21590, B => n21589, ZN => n21595);
   U22561 : XNOR2_X1 port map( A => n21591, B => n1831, ZN => n21592);
   U22562 : XNOR2_X1 port map( A => n21593, B => n21592, ZN => n21594);
   U22563 : XNOR2_X1 port map( A => n21597, B => n21596, ZN => n22016);
   U22564 : XNOR2_X1 port map( A => n22016, B => n21598, ZN => n21605);
   U22565 : XNOR2_X1 port map( A => n21599, B => n21600, ZN => n21603);
   U22566 : XNOR2_X1 port map( A => n21601, B => n21861, ZN => n21602);
   U22567 : XNOR2_X1 port map( A => n21603, B => n21602, ZN => n21604);
   U22568 : NAND2_X1 port map( A1 => n24885, A2 => n22954, ZN => n21878);
   U22569 : XNOR2_X1 port map( A => n21687, B => n21606, ZN => n21610);
   U22570 : INV_X1 port map( A => n494, ZN => n21607);
   U22571 : XNOR2_X1 port map( A => n21608, B => n21607, ZN => n21609);
   U22572 : XNOR2_X1 port map( A => n21610, B => n21609, ZN => n21613);
   U22573 : INV_X1 port map( A => n22027, ZN => n22829);
   U22574 : XNOR2_X1 port map( A => n21614, B => n21615, ZN => n21620);
   U22575 : INV_X1 port map( A => n3062, ZN => n22875);
   U22576 : XNOR2_X1 port map( A => n21616, B => n22875, ZN => n21617);
   U22577 : XNOR2_X1 port map( A => n21618, B => n21617, ZN => n21619);
   U22579 : XNOR2_X1 port map( A => n21622, B => n21621, ZN => n21625);
   U22580 : INV_X1 port map( A => n21623, ZN => n23916);
   U22581 : XNOR2_X1 port map( A => n21693, B => n23916, ZN => n21624);
   U22582 : XNOR2_X1 port map( A => n21625, B => n21624, ZN => n21629);
   U22583 : XNOR2_X1 port map( A => n21626, B => n21627, ZN => n21628);
   U22584 : XNOR2_X1 port map( A => n21632, B => n21631, ZN => n21637);
   U22585 : XNOR2_X1 port map( A => n21633, B => n23602, ZN => n21634);
   U22586 : XNOR2_X1 port map( A => n21635, B => n21634, ZN => n21636);
   U22587 : INV_X1 port map( A => n22938, ZN => n21644);
   U22588 : INV_X1 port map( A => n92, ZN => n23322);
   U22589 : XNOR2_X1 port map( A => n21525, B => n23322, ZN => n21638);
   U22590 : XNOR2_X1 port map( A => n25065, B => n21639, ZN => n21641);
   U22592 : MUX2_X1 port map( A => n21644, B => n25063, S => n24932, Z => 
                           n21656);
   U22593 : XNOR2_X1 port map( A => n21645, B => n21646, ZN => n21652);
   U22594 : XNOR2_X1 port map( A => n21647, B => n1777, ZN => n21650);
   U22595 : XNOR2_X1 port map( A => n21651, B => n21652, ZN => n22722);
   U22596 : INV_X1 port map( A => n22722, ZN => n22941);
   U22598 : NAND2_X1 port map( A1 => n22832, A2 => n22939, ZN => n21653);
   U22599 : MUX2_X1 port map( A => n21654, B => n21653, S => n22027, Z => 
                           n21655);
   U22600 : NAND2_X1 port map( A1 => n23374, A2 => n23379, ZN => n22430);
   U22601 : XNOR2_X1 port map( A => n25498, B => n21658, ZN => n21661);
   U22602 : INV_X1 port map( A => n21662, ZN => n23763);
   U22603 : XNOR2_X1 port map( A => n21027, B => n23763, ZN => n21663);
   U22604 : XNOR2_X1 port map( A => n21664, B => n24898, ZN => n21666);
   U22605 : XNOR2_X1 port map( A => n21669, B => n21668, ZN => n21674);
   U22606 : XNOR2_X1 port map( A => n21670, B => n16574, ZN => n21672);
   U22607 : XNOR2_X1 port map( A => n21671, B => n21672, ZN => n21673);
   U22609 : XNOR2_X1 port map( A => n21675, B => n1789, ZN => n21677);
   U22610 : XNOR2_X1 port map( A => n21677, B => n21676, ZN => n21681);
   U22611 : XNOR2_X1 port map( A => n21679, B => n21678, ZN => n21680);
   U22612 : XNOR2_X1 port map( A => n21681, B => n21680, ZN => n21682);
   U22613 : XNOR2_X1 port map( A => n21685, B => n21684, ZN => n21691);
   U22614 : XNOR2_X1 port map( A => n21686, B => n5433, ZN => n21688);
   U22615 : XNOR2_X1 port map( A => n21691, B => n21690, ZN => n22483);
   U22617 : OAI22_X1 port map( A1 => n21692, A2 => n22901, B1 => n22842, B2 => 
                           n25569, ZN => n21710);
   U22618 : XNOR2_X1 port map( A => n21693, B => n447, ZN => n21695);
   U22619 : NAND2_X1 port map( A1 => n25569, A2 => n22900, ZN => n21709);
   U22620 : XNOR2_X1 port map( A => n25202, B => n21699, ZN => n21702);
   U22621 : XNOR2_X1 port map( A => n21702, B => n21701, ZN => n21708);
   U22622 : INV_X1 port map( A => n21703, ZN => n23330);
   U22623 : XNOR2_X1 port map( A => n21704, B => n23330, ZN => n21705);
   U22624 : XNOR2_X1 port map( A => n21706, B => n21705, ZN => n21707);
   U22625 : XNOR2_X1 port map( A => n21708, B => n21707, ZN => n22905);
   U22626 : INV_X1 port map( A => n22905, ZN => n22907);
   U22627 : INV_X1 port map( A => n22070, ZN => n21712);
   U22629 : XNOR2_X1 port map( A => n21713, B => n3118, ZN => n21714);
   U22630 : XNOR2_X1 port map( A => n21715, B => n21714, ZN => n21719);
   U22631 : XNOR2_X1 port map( A => n21717, B => n21716, ZN => n21718);
   U22632 : XNOR2_X2 port map( A => n21718, B => n21719, ZN => n23016);
   U22633 : XNOR2_X1 port map( A => n21721, B => n21720, ZN => n21722);
   U22634 : XNOR2_X1 port map( A => n20727, B => n3901, ZN => n21724);
   U22635 : XNOR2_X1 port map( A => n21726, B => n21727, ZN => n21733);
   U22636 : XNOR2_X1 port map( A => n24985, B => n21728, ZN => n21731);
   U22637 : XNOR2_X1 port map( A => n21729, B => n22382, ZN => n21730);
   U22638 : XNOR2_X1 port map( A => n21731, B => n21730, ZN => n21732);
   U22639 : XNOR2_X1 port map( A => n21733, B => n21732, ZN => n23458);
   U22640 : NAND2_X1 port map( A1 => n23016, A2 => n23458, ZN => n21741);
   U22641 : XNOR2_X1 port map( A => n21736, B => n2747, ZN => n21737);
   U22642 : XNOR2_X1 port map( A => n21738, B => n21739, ZN => n21740);
   U22643 : MUX2_X1 port map( A => n22914, B => n21741, S => n24877, Z => 
                           n21758);
   U22644 : XNOR2_X1 port map( A => n1326, B => n21742, ZN => n21744);
   U22645 : XNOR2_X1 port map( A => n21745, B => n21744, ZN => n21746);
   U22646 : XNOR2_X1 port map( A => n21747, B => n21746, ZN => n21749);
   U22647 : XNOR2_X2 port map( A => n21749, B => n21748, ZN => n23464);
   U22648 : INV_X1 port map( A => n23016, ZN => n23460);
   U22649 : XNOR2_X1 port map( A => n21751, B => n21750, ZN => n21753);
   U22650 : XNOR2_X1 port map( A => n21753, B => n21752, ZN => n21757);
   U22651 : XNOR2_X1 port map( A => n21754, B => n21755, ZN => n21756);
   U22652 : XNOR2_X1 port map( A => n21756, B => n21757, ZN => n23015);
   U22653 : NAND2_X1 port map( A1 => n24611, A2 => n23595, ZN => n22639);
   U22654 : INV_X1 port map( A => n23575, ZN => n22079);
   U22655 : INV_X1 port map( A => n21759, ZN => n23576);
   U22656 : AOI21_X1 port map( B1 => n22079, B2 => n23576, A => n22176, ZN => 
                           n21760);
   U22657 : INV_X1 port map( A => n23566, ZN => n21763);
   U22658 : INV_X1 port map( A => n22922, ZN => n22107);
   U22659 : INV_X1 port map( A => n22209, ZN => n21767);
   U22660 : OAI21_X1 port map( B1 => n24333, B2 => n22208, A => n21767, ZN => 
                           n21764);
   U22661 : NOR2_X1 port map( A1 => n21765, A2 => n21764, ZN => n21771);
   U22662 : NOR2_X1 port map( A1 => n22159, A2 => n22206, ZN => n21768);
   U22663 : NOR2_X1 port map( A1 => n21768, A2 => n21767, ZN => n21770);
   U22664 : NAND2_X1 port map( A1 => n22159, A2 => n24333, ZN => n21769);
   U22665 : INV_X1 port map( A => n23596, ZN => n22633);
   U22666 : INV_X1 port map( A => n22889, ZN => n22496);
   U22668 : AOI22_X1 port map( A1 => n21772, A2 => n22887, B1 => n22729, B2 => 
                           n22890, ZN => n21773);
   U22669 : NAND3_X1 port map( A1 => n24390, A2 => n22633, A3 => n24901, ZN => 
                           n21776);
   U22670 : NOR2_X1 port map( A1 => n24390, A2 => n24397, ZN => n21947);
   U22671 : NAND2_X1 port map( A1 => n21947, A2 => n23596, ZN => n21775);
   U22672 : NAND4_X1 port map( A1 => n22639, A2 => n21777, A3 => n21776, A4 => 
                           n21775, ZN => n21779);
   U22673 : INV_X1 port map( A => n1801, ZN => n21778);
   U22674 : XNOR2_X1 port map( A => n21779, B => n21778, ZN => Ciphertext(114))
                           ;
   U22676 : AOI21_X1 port map( B1 => n24114, B2 => n21838, A => n21839, ZN => 
                           n21785);
   U22677 : NOR2_X1 port map( A1 => n22355, A2 => n22354, ZN => n21781);
   U22678 : NAND2_X1 port map( A1 => n21781, A2 => n22356, ZN => n21784);
   U22679 : NOR2_X1 port map( A1 => n21782, A2 => n21839, ZN => n21845);
   U22681 : NAND2_X1 port map( A1 => n21845, A2 => n25082, ZN => n21783);
   U22683 : INV_X1 port map( A => n23757, ZN => n21800);
   U22686 : INV_X1 port map( A => n22244, ZN => n21815);
   U22689 : NOR2_X1 port map( A1 => n21800, A2 => n23769, ZN => n21795);
   U22690 : MUX2_X1 port map( A => n25461, B => n22217, S => n22221, Z => 
                           n21790);
   U22691 : NAND2_X1 port map( A1 => n21829, A2 => n22222, ZN => n21789);
   U22692 : NOR2_X1 port map( A1 => n25051, A2 => n24921, ZN => n23771);
   U22693 : NAND2_X1 port map( A1 => n22231, A2 => n22226, ZN => n21792);
   U22694 : NOR2_X1 port map( A1 => n22233, A2 => n22226, ZN => n21793);
   U22695 : OAI21_X1 port map( B1 => n21795, B2 => n23771, A => n23779, ZN => 
                           n21809);
   U22696 : INV_X1 port map( A => n23752, ZN => n21798);
   U22697 : NAND2_X1 port map( A1 => n22522, A2 => n22255, ZN => n21797);
   U22699 : NAND2_X1 port map( A1 => n22521, A2 => n4373, ZN => n21796);
   U22700 : NAND3_X1 port map( A1 => n21798, A2 => n21797, A3 => n21796, ZN => 
                           n21799);
   U22701 : NAND3_X1 port map( A1 => n25051, A2 => n21800, A3 => n21799, ZN => 
                           n21808);
   U22702 : NOR2_X1 port map( A1 => n22079, A2 => n22197, ZN => n21801);
   U22703 : NOR2_X1 port map( A1 => n21802, A2 => n21801, ZN => n21805);
   U22704 : NOR2_X1 port map( A1 => n22079, A2 => n24369, ZN => n21803);
   U22705 : NAND2_X1 port map( A1 => n23768, A2 => n24921, ZN => n21806);
   U22706 : NAND3_X1 port map( A1 => n21809, A2 => n21808, A3 => n21807, ZN => 
                           n21811);
   U22707 : INV_X1 port map( A => n1777, ZN => n21810);
   U22708 : XNOR2_X1 port map( A => n21811, B => n21810, ZN => Ciphertext(146))
                           ;
   U22709 : NOR2_X1 port map( A1 => n22243, A2 => n22239, ZN => n21814);
   U22710 : INV_X1 port map( A => n22184, ZN => n21813);
   U22711 : NAND2_X1 port map( A1 => n21815, A2 => n22243, ZN => n23001);
   U22712 : NOR2_X1 port map( A1 => n21848, A2 => n21816, ZN => n22348);
   U22714 : NAND3_X1 port map( A1 => n21848, A2 => n22688, A3 => n22685, ZN => 
                           n21820);
   U22715 : NAND2_X1 port map( A1 => n21848, A2 => n21817, ZN => n21818);
   U22716 : NOR2_X1 port map( A1 => n24468, A2 => n21841, ZN => n21824);
   U22717 : NOR2_X1 port map( A1 => n332, A2 => n21825, ZN => n21823);
   U22718 : MUX2_X1 port map( A => n21824, B => n21823, S => n21822, Z => 
                           n21827);
   U22719 : NAND2_X1 port map( A1 => n24362, A2 => n21841, ZN => n21826);
   U22721 : NOR2_X1 port map( A1 => n22214, A2 => n22221, ZN => n21832);
   U22722 : NAND2_X1 port map( A1 => n22222, A2 => n24918, ZN => n21831);
   U22723 : NAND2_X1 port map( A1 => n22216, A2 => n22221, ZN => n22218);
   U22724 : OAI211_X1 port map( C1 => n21832, C2 => n21831, A => n22218, B => 
                           n21830, ZN => n23799);
   U22725 : NAND3_X1 port map( A1 => n24307, A2 => n24895, A3 => n24920, ZN => 
                           n21833);
   U22726 : NAND2_X1 port map( A1 => n22233, A2 => n22225, ZN => n21834);
   U22729 : MUX2_X1 port map( A => n21845, B => n22356, S => n21844, Z => 
                           n23893);
   U22730 : NAND2_X1 port map( A1 => n22355, A2 => n22354, ZN => n21846);
   U22731 : AND2_X1 port map( A1 => n22359, A2 => n21846, ZN => n23892);
   U22732 : NOR2_X2 port map( A1 => n23893, A2 => n23892, ZN => n23904);
   U22733 : MUX2_X1 port map( A => n22689, B => n22685, S => n22688, Z => 
                           n21849);
   U22734 : MUX2_X2 port map( A => n21850, B => n21849, S => n22687, Z => 
                           n23905);
   U22737 : INV_X1 port map( A => n21866, ZN => n21851);
   U22738 : NAND2_X1 port map( A1 => n21851, A2 => n21861, ZN => n21870);
   U22739 : NAND2_X1 port map( A1 => n22813, A2 => n4469, ZN => n21852);
   U22741 : AOI22_X1 port map( A1 => n25439, A2 => n22677, B1 => n23998, B2 => 
                           n25414, ZN => n22598);
   U22742 : INV_X1 port map( A => n23995, ZN => n22596);
   U22743 : OAI21_X1 port map( B1 => n22596, B2 => n24439, A => n23998, ZN => 
                           n21853);
   U22744 : INV_X1 port map( A => n23994, ZN => n22678);
   U22745 : NAND2_X1 port map( A1 => n21853, A2 => n22678, ZN => n21854);
   U22746 : AOI21_X1 port map( B1 => n23906, B2 => n23889, A => n23905, ZN => 
                           n21869);
   U22747 : AND2_X1 port map( A1 => n21856, A2 => n22679, ZN => n21858);
   U22748 : NOR2_X1 port map( A1 => n22769, A2 => n22770, ZN => n21857);
   U22749 : MUX2_X1 port map( A => n21858, B => n21857, S => n22774, Z => 
                           n23891);
   U22750 : NOR2_X1 port map( A1 => n23890, A2 => n16, ZN => n21860);
   U22751 : NAND2_X1 port map( A1 => n23879, A2 => n23889, ZN => n21859);
   U22752 : OAI211_X1 port map( C1 => n23905, C2 => n23879, A => n21860, B => 
                           n21859, ZN => n21868);
   U22753 : NOR2_X1 port map( A1 => n23890, A2 => n23889, ZN => n21862);
   U22754 : AOI21_X1 port map( B1 => n21862, B2 => n23879, A => n21861, ZN => 
                           n21865);
   U22756 : NAND2_X1 port map( A1 => n23909, A2 => n23903, ZN => n21864);
   U22759 : INV_X1 port map( A => n22852, ZN => n22933);
   U22761 : NAND2_X1 port map( A1 => n22426, A2 => n22947, ZN => n21874);
   U22762 : NAND3_X1 port map( A1 => n22422, A2 => n22420, A3 => n22421, ZN => 
                           n21873);
   U22763 : OAI21_X1 port map( B1 => n21874, B2 => n22948, A => n21873, ZN => 
                           n21877);
   U22765 : NAND2_X1 port map( A1 => n23317, A2 => n23326, ZN => n22629);
   U22766 : INV_X1 port map( A => n21878, ZN => n21882);
   U22767 : OAI21_X1 port map( B1 => n22954, B2 => n22953, A => n22033, ZN => 
                           n21881);
   U22768 : NOR2_X1 port map( A1 => n24885, A2 => n22033, ZN => n22394);
   U22769 : AOI21_X1 port map( B1 => n22394, B2 => n24922, A => n21879, ZN => 
                           n21880);
   U22770 : OAI21_X1 port map( B1 => n21882, B2 => n21881, A => n21880, ZN => 
                           n23324);
   U22771 : INV_X1 port map( A => n23324, ZN => n23313);
   U22772 : OR2_X1 port map( A1 => n22629, A2 => n23313, ZN => n21897);
   U22773 : INV_X1 port map( A => n22397, ZN => n21883);
   U22774 : NAND2_X1 port map( A1 => n22398, A2 => n22265, ZN => n21887);
   U22775 : INV_X1 port map( A => n25381, ZN => n21884);
   U22776 : OAI21_X1 port map( B1 => n21885, B2 => n22397, A => n21884, ZN => 
                           n21886);
   U22777 : NOR2_X1 port map( A1 => n22397, A2 => n22134, ZN => n22268);
   U22778 : INV_X1 port map( A => n21888, ZN => n22396);
   U22779 : NAND2_X1 port map( A1 => n22968, A2 => n21467, ZN => n21956);
   U22780 : NAND3_X1 port map( A1 => n22962, A2 => n21476, A3 => n22969, ZN => 
                           n21890);
   U22781 : NAND2_X1 port map( A1 => n24411, A2 => n22965, ZN => n21889);
   U22782 : NAND3_X1 port map( A1 => n23327, A2 => n23318, A3 => n4108, ZN => 
                           n21896);
   U22783 : INV_X1 port map( A => n22975, ZN => n21892);
   U22784 : NOR2_X1 port map( A1 => n21892, A2 => n24881, ZN => n21893);
   U22785 : NOR3_X1 port map( A1 => n21893, A2 => n22977, A3 => n3213, ZN => 
                           n21894);
   U22786 : INV_X1 port map( A => n2039, ZN => n21898);
   U22787 : XNOR2_X1 port map( A => n21899, B => n21898, ZN => Ciphertext(63));
   U22788 : INV_X1 port map( A => n23805, ZN => n23788);
   U22789 : NAND2_X1 port map( A1 => n23787, A2 => n21902, ZN => n21901);
   U22790 : OAI211_X1 port map( C1 => n23805, C2 => n21901, A => Key(33), B => 
                           n21900, ZN => n21906);
   U22791 : INV_X1 port map( A => Key(33), ZN => n21903);
   U22792 : NAND2_X1 port map( A1 => n21907, A2 => n21903, ZN => n21904);
   U22793 : OAI211_X1 port map( C1 => n21907, C2 => n21906, A => n21905, B => 
                           n21904, ZN => Ciphertext(153));
   U22794 : NAND2_X1 port map( A1 => n21909, A2 => n24415, ZN => n21913);
   U22795 : AND2_X1 port map( A1 => n22334, A2 => n22139, ZN => n22273);
   U22796 : NOR2_X1 port map( A1 => n22335, A2 => n21910, ZN => n22142);
   U22797 : NAND2_X1 port map( A1 => n22142, A2 => n22274, ZN => n21912);
   U22798 : NAND3_X1 port map( A1 => n22333, A2 => n22139, A3 => n21910, ZN => 
                           n21911);
   U22799 : OR2_X1 port map( A1 => n21914, A2 => n22134, ZN => n21916);
   U22800 : AND2_X1 port map( A1 => n22396, A2 => n22134, ZN => n22404);
   U22802 : NOR2_X1 port map( A1 => n21918, A2 => n24311, ZN => n21919);
   U22803 : AND2_X1 port map( A1 => n25066, A2 => n21921, ZN => n21922);
   U22805 : OAI21_X1 port map( B1 => n24043, B2 => n22448, A => n274, ZN => 
                           n21926);
   U22806 : INV_X1 port map( A => n22448, ZN => n21924);
   U22808 : OAI21_X1 port map( B1 => n21929, B2 => n22464, A => n21928, ZN => 
                           n21933);
   U22809 : INV_X1 port map( A => n22562, ZN => n22341);
   U22810 : INV_X1 port map( A => n22407, ZN => n22567);
   U22811 : NOR2_X1 port map( A1 => n22341, A2 => n22567, ZN => n21935);
   U22812 : NOR2_X1 port map( A1 => n333, A2 => n22409, ZN => n22411);
   U22813 : INV_X1 port map( A => n22411, ZN => n21937);
   U22815 : INV_X1 port map( A => n21946, ZN => n21940);
   U22816 : NAND3_X1 port map( A1 => n23595, A2 => n24390, A3 => n1328, ZN => 
                           n21939);
   U22817 : OAI211_X1 port map( C1 => n22633, C2 => n21940, A => n21942, B => 
                           n21939, ZN => n21952);
   U22818 : INV_X1 port map( A => n23592, ZN => n21941);
   U22819 : NAND2_X1 port map( A1 => n24372, A2 => n23566, ZN => n22634);
   U22820 : OR2_X1 port map( A1 => n21943, A2 => n21942, ZN => n21950);
   U22821 : AOI21_X1 port map( B1 => n22633, B2 => n21946, A => n21945, ZN => 
                           n21948);
   U22822 : INV_X1 port map( A => n21947, ZN => n22632);
   U22823 : OAI211_X1 port map( C1 => n24611, C2 => n22634, A => n21948, B => 
                           n22632, ZN => n21949);
   U22824 : INV_X1 port map( A => n23374, ZN => n23370);
   U22825 : AOI21_X1 port map( B1 => n24515, B2 => n24911, A => n24404, ZN => 
                           n21953);
   U22826 : NAND2_X1 port map( A1 => n21954, A2 => n21953, ZN => n21955);
   U22827 : NAND2_X1 port map( A1 => n24515, A2 => n22987, ZN => n22744);
   U22828 : OAI21_X1 port map( B1 => n22966, B2 => n22969, A => n21956, ZN => 
                           n21957);
   U22829 : INV_X1 port map( A => n21957, ZN => n21962);
   U22830 : NAND2_X1 port map( A1 => n22962, A2 => n24411, ZN => n21958);
   U22831 : NOR2_X1 port map( A1 => n334, A2 => n24411, ZN => n21960);
   U22832 : AOI21_X2 port map( B1 => n21962, B2 => n21961, A => n21960, ZN => 
                           n23396);
   U22833 : INV_X1 port map( A => n23396, ZN => n22032);
   U22834 : INV_X1 port map( A => n21963, ZN => n21969);
   U22835 : XNOR2_X1 port map( A => n21965, B => n21964, ZN => n21966);
   U22836 : XNOR2_X1 port map( A => n21966, B => n21967, ZN => n21968);
   U22837 : XNOR2_X1 port map( A => n21968, B => n21969, ZN => n21973);
   U22838 : XNOR2_X1 port map( A => n21971, B => n21970, ZN => n21972);
   U22839 : XNOR2_X1 port map( A => n21974, B => n924, ZN => n21976);
   U22840 : XNOR2_X1 port map( A => n21976, B => n21975, ZN => n21978);
   U22841 : XNOR2_X1 port map( A => n21977, B => n21978, ZN => n21984);
   U22842 : XNOR2_X1 port map( A => n21979, B => n21980, ZN => n21982);
   U22843 : XNOR2_X1 port map( A => n21982, B => n21981, ZN => n21983);
   U22845 : XNOR2_X1 port map( A => n21986, B => n21987, ZN => n21991);
   U22846 : XNOR2_X1 port map( A => n20727, B => n3900, ZN => n21988);
   U22847 : XNOR2_X1 port map( A => n21989, B => n21988, ZN => n21990);
   U22851 : XNOR2_X1 port map( A => n25091, B => n21996, ZN => n22000);
   U22852 : XNOR2_X1 port map( A => n21998, B => n1863, ZN => n21999);
   U22853 : XNOR2_X1 port map( A => n22000, B => n21999, ZN => n22001);
   U22854 : XNOR2_X1 port map( A => n22002, B => n22001, ZN => n22836);
   U22855 : XNOR2_X1 port map( A => n22004, B => n22003, ZN => n22011);
   U22856 : INV_X1 port map( A => n1874, ZN => n23922);
   U22857 : XNOR2_X1 port map( A => n22005, B => n23922, ZN => n22009);
   U22858 : XNOR2_X1 port map( A => n22007, B => n22006, ZN => n22008);
   U22859 : XNOR2_X1 port map( A => n22008, B => n22009, ZN => n22010);
   U22860 : XNOR2_X1 port map( A => n22011, B => n22010, ZN => n22837);
   U22861 : OAI22_X1 port map( A1 => n22838, A2 => n22893, B1 => n22836, B2 => 
                           n22837, ZN => n22896);
   U22862 : XNOR2_X1 port map( A => n22012, B => n22013, ZN => n22018);
   U22863 : INV_X1 port map( A => n2772, ZN => n23775);
   U22864 : XNOR2_X1 port map( A => n22014, B => n23775, ZN => n22015);
   U22865 : XNOR2_X1 port map( A => n22016, B => n22015, ZN => n22017);
   U22866 : INV_X1 port map( A => n22837, ZN => n22841);
   U22867 : OAI21_X1 port map( B1 => n25041, B2 => n22836, A => n22841, ZN => 
                           n22019);
   U22868 : NAND3_X1 port map( A1 => n25382, A2 => n22905, A3 => n22842, ZN => 
                           n22025);
   U22869 : INV_X1 port map( A => n22842, ZN => n22906);
   U22870 : NAND3_X1 port map( A1 => n22906, A2 => n25569, A3 => n22901, ZN => 
                           n22024);
   U22871 : NOR2_X1 port map( A1 => n22901, A2 => n22483, ZN => n22903);
   U22872 : NAND2_X1 port map( A1 => n22903, A2 => n22904, ZN => n22023);
   U22873 : NOR2_X1 port map( A1 => n25569, A2 => n22900, ZN => n22021);
   U22874 : NAND2_X1 port map( A1 => n22021, A2 => n22906, ZN => n22022);
   U22875 : INV_X1 port map( A => n22940, ZN => n22936);
   U22876 : OAI21_X1 port map( B1 => n22936, B2 => n22938, A => n22832, ZN => 
                           n22030);
   U22877 : NOR2_X1 port map( A1 => n22940, A2 => n22722, ZN => n22029);
   U22878 : NAND2_X1 port map( A1 => n22029, A2 => n22939, ZN => n22028);
   U22880 : INV_X1 port map( A => n24449, ZN => n22031);
   U22881 : AOI22_X1 port map( A1 => n24884, A2 => n22953, B1 => n22952, B2 => 
                           n22033, ZN => n22393);
   U22882 : NAND3_X1 port map( A1 => n22034, A2 => n24922, A3 => n22954, ZN => 
                           n22035);
   U22883 : INV_X1 port map( A => n23394, ZN => n22036);
   U22884 : NOR3_X1 port map( A1 => n24933, A2 => n22036, A3 => n24465, ZN => 
                           n22040);
   U22885 : MUX2_X1 port map( A => n24341, B => n22852, S => n23332, Z => 
                           n22038);
   U22886 : MUX2_X1 port map( A => n23334, B => n25081, S => n22501, Z => 
                           n22037);
   U22888 : NOR3_X1 port map( A1 => n324, A2 => n23392, A3 => n24465, ZN => 
                           n22039);
   U22889 : NOR3_X1 port map( A1 => n22041, A2 => n22040, A3 => n22039, ZN => 
                           n22042);
   U22890 : XNOR2_X1 port map( A => n22042, B => n677, ZN => Ciphertext(78));
   U22891 : NAND2_X1 port map( A1 => n22044, A2 => n23805, ZN => n22048);
   U22892 : NOR3_X1 port map( A1 => n22046, A2 => n23002, A3 => n22045, ZN => 
                           n22047);
   U22893 : OAI21_X1 port map( B1 => n21829, B2 => n22217, A => n25461, ZN => 
                           n22054);
   U22894 : NAND2_X1 port map( A1 => n22216, A2 => n22214, ZN => n22050);
   U22895 : NAND2_X1 port map( A1 => n22050, A2 => n2817, ZN => n22052);
   U22898 : NOR2_X1 port map( A1 => n22239, A2 => n22059, ZN => n22060);
   U22899 : AOI22_X1 port map( A1 => n22184, A2 => n1336, B1 => n22243, B2 => 
                           n22060, ZN => n22061);
   U22900 : OAI21_X1 port map( B1 => n22063, B2 => n22062, A => n22061, ZN => 
                           n23697);
   U22901 : INV_X1 port map( A => n22212, ZN => n22068);
   U22902 : AOI22_X2 port map( A1 => n22067, A2 => n22068, B1 => n22065, B2 => 
                           n22066, ZN => n23720);
   U22903 : INV_X1 port map( A => n22916, ZN => n22170);
   U22905 : NOR2_X1 port map( A1 => n24674, A2 => n22166, ZN => n22071);
   U22909 : NOR2_X2 port map( A1 => n22075, A2 => n22074, ZN => n23712);
   U22910 : NOR2_X1 port map( A1 => n23712, A2 => n23720, ZN => n23724);
   U22911 : INV_X1 port map( A => n3125, ZN => n22082);
   U22912 : AOI21_X1 port map( B1 => n23724, B2 => n22082, A => n23714, ZN => 
                           n22077);
   U22913 : OR2_X1 port map( A1 => n23724, A2 => n22082, ZN => n22076);
   U22914 : OAI211_X1 port map( C1 => n23696, C2 => n22148, A => n22077, B => 
                           n22076, ZN => n22085);
   U22916 : AND2_X1 port map( A1 => n23571, A2 => n22200, ZN => n22081);
   U22917 : NAND4_X1 port map( A1 => n24374, A2 => n22082, A3 => n22148, A4 => 
                           n23714, ZN => n22083);
   U22918 : INV_X1 port map( A => n23712, ZN => n23719);
   U22919 : OAI21_X1 port map( B1 => n23723, B2 => n23720, A => n23721, ZN => 
                           n22086);
   U22920 : OAI21_X1 port map( B1 => n23719, B2 => n24381, A => n22086, ZN => 
                           n22091);
   U22921 : NAND2_X1 port map( A1 => n23714, A2 => n22089, ZN => n22087);
   U22922 : AOI21_X1 port map( B1 => n23723, B2 => n24381, A => n22087, ZN => 
                           n22088);
   U22923 : OAI21_X1 port map( B1 => n24374, B2 => n23723, A => n22088, ZN => 
                           n22090);
   U22925 : NAND2_X1 port map( A1 => n22496, A2 => n22093, ZN => n22099);
   U22926 : NOR2_X1 port map( A1 => n22890, A2 => n327, ZN => n22097);
   U22927 : INV_X1 port map( A => n22887, ZN => n22494);
   U22928 : OAI21_X1 port map( B1 => n25375, B2 => n22494, A => n22095, ZN => 
                           n22096);
   U22929 : NAND2_X1 port map( A1 => n24877, A2 => n23014, ZN => n22100);
   U22931 : AND3_X1 port map( A1 => n22100, A2 => n24364, A3 => n23016, ZN => 
                           n22102);
   U22932 : AND2_X1 port map( A1 => n23015, A2 => n23458, ZN => n22862);
   U22933 : AND2_X1 port map( A1 => n23014, A2 => n22862, ZN => n22101);
   U22934 : NOR3_X2 port map( A1 => n22102, A2 => n22863, A3 => n22101, ZN => 
                           n23555);
   U22935 : INV_X1 port map( A => n22893, ZN => n22834);
   U22936 : NAND2_X1 port map( A1 => n22834, A2 => n25438, ZN => n22897);
   U22937 : NAND2_X1 port map( A1 => n22717, A2 => n25041, ZN => n22103);
   U22938 : AOI21_X1 port map( B1 => n22897, B2 => n22103, A => n22835, ZN => 
                           n22106);
   U22939 : NAND2_X1 port map( A1 => n22835, A2 => n22834, ZN => n22104);
   U22940 : AOI21_X1 port map( B1 => n22104, B2 => n22837, A => n25041, ZN => 
                           n22105);
   U22941 : NOR2_X1 port map( A1 => n22106, A2 => n22105, ZN => n23547);
   U22942 : OAI22_X1 port map( A1 => n323, A2 => n23554, B1 => n23555, B2 => 
                           n23547, ZN => n22701);
   U22943 : INV_X1 port map( A => n22926, ZN => n22929);
   U22945 : NAND2_X1 port map( A1 => n25479, A2 => n22188, ZN => n22109);
   U22946 : NAND3_X1 port map( A1 => n25070, A2 => n22107, A3 => n22927, ZN => 
                           n22108);
   U22947 : AND2_X1 port map( A1 => n24379, A2 => n22927, ZN => n22110);
   U22948 : INV_X1 port map( A => n22110, ZN => n22111);
   U22949 : AND2_X1 port map( A1 => n25071, A2 => n23555, ZN => n23551);
   U22950 : MUX2_X1 port map( A => n21712, B => n22166, S => n22916, Z => 
                           n22114);
   U22951 : INV_X1 port map( A => n22918, ZN => n22113);
   U22952 : NAND2_X1 port map( A1 => n22114, A2 => n22113, ZN => n22120);
   U22953 : OR2_X1 port map( A1 => n22115, A2 => n22917, ZN => n22119);
   U22954 : INV_X1 port map( A => n22116, ZN => n22117);
   U22955 : NAND2_X1 port map( A1 => n323, A2 => n23537, ZN => n22121);
   U22956 : AOI22_X1 port map( A1 => n22701, A2 => n23544, B1 => n23551, B2 => 
                           n22121, ZN => n22122);
   U22957 : XNOR2_X1 port map( A => n22122, B => n1767, ZN => Ciphertext(109));
   U22958 : NOR3_X1 port map( A1 => n22948, A2 => n22426, A3 => n22422, ZN => 
                           n22124);
   U22959 : NOR3_X1 port map( A1 => n22282, A2 => n22421, A3 => n22946, ZN => 
                           n22123);
   U22960 : NOR2_X1 port map( A1 => n22124, A2 => n22123, ZN => n22127);
   U22961 : AOI21_X1 port map( B1 => n22963, B2 => n22129, A => n22128, ZN => 
                           n22130);
   U22963 : NOR2_X1 port map( A1 => n22536, A2 => n24907, ZN => n22145);
   U22964 : INV_X1 port map( A => n22134, ZN => n22261);
   U22966 : NAND2_X1 port map( A1 => n22337, A2 => n22138, ZN => n22140);
   U22967 : OAI21_X1 port map( B1 => n5767, B2 => n22337, A => n22140, ZN => 
                           n22143);
   U22968 : AOI21_X1 port map( B1 => n22145, B2 => n24360, A => n22144, ZN => 
                           n22146);
   U22969 : XNOR2_X1 port map( A => n22146, B => n2145, ZN => Ciphertext(49));
   U22970 : NAND3_X1 port map( A1 => n23712, A2 => n24381, A3 => n23716, ZN => 
                           n22149);
   U22973 : OAI21_X1 port map( B1 => n22159, B2 => n22156, A => n22155, ZN => 
                           n22157);
   U22974 : INV_X1 port map( A => n25485, ZN => n22158);
   U22976 : NAND2_X1 port map( A1 => n22218, A2 => n22162, ZN => n22165);
   U22977 : OAI21_X1 port map( B1 => n22222, B2 => n22217, A => n21829, ZN => 
                           n22163);
   U22978 : AND2_X1 port map( A1 => n25461, A2 => n22163, ZN => n22164);
   U22980 : INV_X1 port map( A => n22166, ZN => n22919);
   U22981 : NOR2_X1 port map( A1 => n22919, A2 => n24902, ZN => n22168);
   U22982 : NAND2_X1 port map( A1 => n22169, A2 => n22168, ZN => n22172);
   U22983 : NAND2_X1 port map( A1 => n23576, A2 => n22175, ZN => n22173);
   U22984 : OAI21_X1 port map( B1 => n23576, B2 => n24396, A => n22173, ZN => 
                           n22174);
   U22985 : INV_X1 port map( A => n22175, ZN => n22199);
   U22986 : NAND3_X1 port map( A1 => n22199, A2 => n1323, A3 => n4360, ZN => 
                           n22177);
   U22987 : NOR2_X1 port map( A1 => n22240, A2 => n22180, ZN => n22182);
   U22988 : OR2_X1 port map( A1 => n1336, A2 => n22244, ZN => n22185);
   U22991 : OAI21_X1 port map( B1 => n23686, B2 => n22186, A => n23658, ZN => 
                           n22194);
   U22993 : INV_X1 port map( A => n25026, ZN => n23678);
   U22995 : OAI21_X1 port map( B1 => n22926, B2 => n25479, A => n22188, ZN => 
                           n22191);
   U22996 : AOI21_X2 port map( B1 => n22192, B2 => n22191, A => n22190, ZN => 
                           n23690);
   U22997 : INV_X1 port map( A => n1855, ZN => n22195);
   U22999 : NAND2_X1 port map( A1 => n24396, A2 => n22197, ZN => n22202);
   U23000 : OAI21_X1 port map( B1 => n22199, B2 => n22202, A => n22198, ZN => 
                           n22204);
   U23001 : OAI22_X1 port map( A1 => n24369, A2 => n22202, B1 => n22201, B2 => 
                           n22175, ZN => n22203);
   U23003 : NAND2_X1 port map( A1 => n22208, A2 => n22206, ZN => n22207);
   U23004 : OAI21_X1 port map( B1 => n22209, B2 => n25018, A => n22207, ZN => 
                           n22210);
   U23006 : NAND2_X1 port map( A1 => n22214, A2 => n22221, ZN => n22215);
   U23007 : OAI22_X1 port map( A1 => n22218, A2 => n24918, B1 => n22216, B2 => 
                           n22215, ZN => n22224);
   U23009 : MUX2_X1 port map( A => n23740, B => n23743, S => n24064, Z => 
                           n22259);
   U23010 : NOR2_X1 port map( A1 => n22226, A2 => n22225, ZN => n22230);
   U23011 : NOR2_X1 port map( A1 => n22228, A2 => n24905, ZN => n22229);
   U23012 : MUX2_X1 port map( A => n22230, B => n22229, S => n22231, Z => 
                           n22238);
   U23013 : INV_X1 port map( A => n22231, ZN => n22234);
   U23014 : AOI21_X1 port map( B1 => n22234, B2 => n22233, A => n22232, ZN => 
                           n22236);
   U23015 : NOR2_X1 port map( A1 => n22236, A2 => n22235, ZN => n22237);
   U23019 : NAND2_X1 port map( A1 => n22240, A2 => n22243, ZN => n22248);
   U23020 : OAI21_X1 port map( B1 => n22243, B2 => n22242, A => n22241, ZN => 
                           n22247);
   U23021 : MUX2_X1 port map( A => n24063, B => n23730, S => n23748, Z => 
                           n22258);
   U23022 : NAND2_X1 port map( A1 => n24468, A2 => n22252, ZN => n22253);
   U23023 : XNOR2_X1 port map( A => n22260, B => n1864, ZN => Ciphertext(140));
   U23024 : AOI22_X1 port map( A1 => n22456, A2 => n5224, B1 => n25487, B2 => 
                           n22324, ZN => n22272);
   U23025 : OAI21_X1 port map( B1 => n22452, B2 => n24496, A => n1352, ZN => 
                           n22271);
   U23026 : OAI21_X1 port map( B1 => n22272, B2 => n24311, A => n22271, ZN => 
                           n23242);
   U23027 : OAI21_X1 port map( B1 => n22338, B2 => n22274, A => n22273, ZN => 
                           n22277);
   U23028 : NAND2_X1 port map( A1 => n21368, A2 => n22275, ZN => n22276);
   U23030 : OAI21_X1 port map( B1 => n24377, B2 => n23242, A => n22298, ZN => 
                           n22278);
   U23031 : XNOR2_X1 port map( A => n22278, B => n4668, ZN => n22297);
   U23032 : AND2_X1 port map( A1 => n22946, A2 => n22421, ZN => n22280);
   U23033 : NOR2_X1 port map( A1 => n22426, A2 => n22947, ZN => n22279);
   U23034 : INV_X1 port map( A => n22421, ZN => n22281);
   U23035 : NAND2_X1 port map( A1 => n22341, A2 => n22409, ZN => n22285);
   U23036 : MUX2_X1 port map( A => n22566, B => n22409, S => n24971, Z => 
                           n22284);
   U23037 : AND2_X1 port map( A1 => n22411, A2 => n22567, ZN => n22286);
   U23038 : INV_X1 port map( A => n22977, ZN => n22288);
   U23039 : NAND2_X1 port map( A1 => n22387, A2 => n22288, ZN => n22291);
   U23040 : INV_X1 port map( A => n22972, ZN => n22388);
   U23041 : AOI21_X1 port map( B1 => n22977, B2 => n22974, A => n22388, ZN => 
                           n22290);
   U23042 : NOR2_X1 port map( A1 => n24881, A2 => n22975, ZN => n22289);
   U23044 : XNOR2_X1 port map( A => n23252, B => n4668, ZN => n22294);
   U23045 : XNOR2_X1 port map( A => n23251, B => n4668, ZN => n22295);
   U23046 : NAND2_X1 port map( A1 => n23256, A2 => n22295, ZN => n22296);
   U23047 : INV_X1 port map( A => n23251, ZN => n23241);
   U23048 : INV_X1 port map( A => n23242, ZN => n23249);
   U23049 : NAND3_X1 port map( A1 => n23245, A2 => n23241, A3 => n23249, ZN => 
                           n22299);
   U23050 : INV_X1 port map( A => n1870, ZN => n22301);
   U23052 : OR2_X1 port map( A1 => n24933, A2 => n23394, ZN => n23385);
   U23053 : AOI21_X1 port map( B1 => n24880, B2 => n23385, A => n23392, ZN => 
                           n22306);
   U23054 : INV_X1 port map( A => n24465, ZN => n22304);
   U23055 : NAND3_X1 port map( A1 => n23396, A2 => n23394, A3 => n23392, ZN => 
                           n22303);
   U23056 : NOR2_X1 port map( A1 => n22306, A2 => n22305, ZN => n22307);
   U23057 : XNOR2_X1 port map( A => n22307, B => n1739, ZN => Ciphertext(79));
   U23059 : NOR2_X1 port map( A1 => n22309, A2 => n23743, ZN => n22311);
   U23061 : XNOR2_X1 port map( A => n22312, B => n62, ZN => Ciphertext(142));
   U23062 : AND2_X1 port map( A1 => n22615, A2 => n22619, ZN => n22472);
   U23063 : INV_X1 port map( A => n22472, ZN => n22316);
   U23064 : NOR2_X1 port map( A1 => n22615, A2 => n22612, ZN => n22788);
   U23065 : OAI21_X1 port map( B1 => n22788, B2 => n22617, A => n22792, ZN => 
                           n22315);
   U23066 : NOR2_X1 port map( A1 => n22448, A2 => n274, ZN => n22321);
   U23067 : NAND2_X1 port map( A1 => n25066, A2 => n22592, ZN => n22320);
   U23068 : NOR2_X1 port map( A1 => n22591, A2 => n22318, ZN => n22319);
   U23069 : OAI21_X1 port map( B1 => n22321, B2 => n22320, A => n22319, ZN => 
                           n23178);
   U23070 : NOR2_X1 port map( A1 => n24496, A2 => n22323, ZN => n22325);
   U23071 : MUX2_X1 port map( A => n23164, B => n23178, S => n23177, Z => 
                           n22345);
   U23072 : INV_X1 port map( A => n23177, ZN => n23168);
   U23073 : OR3_X1 port map( A1 => n22462, A2 => n22465, A3 => n22464, ZN => 
                           n22332);
   U23074 : INV_X1 port map( A => n22328, ZN => n22330);
   U23075 : OAI21_X1 port map( B1 => n22511, B2 => n25496, A => n23165, ZN => 
                           n22340);
   U23076 : MUX2_X1 port map( A => n22338, B => n4350, S => n22337, Z => n22512
                           );
   U23077 : NOR2_X1 port map( A1 => n22512, A2 => n22511, ZN => n22339);
   U23078 : OAI22_X1 port map( A1 => n23168, A2 => n23165, B1 => n22340, B2 => 
                           n22339, ZN => n22344);
   U23079 : INV_X1 port map( A => n22566, ZN => n22412);
   U23080 : OAI21_X1 port map( B1 => n22409, B2 => n22407, A => n22341, ZN => 
                           n22342);
   U23082 : INV_X1 port map( A => n2005, ZN => n22346);
   U23083 : XNOR2_X1 port map( A => n22347, B => n22346, ZN => Ciphertext(26));
   U23085 : INV_X1 port map( A => n22348, ZN => n22351);
   U23086 : NAND2_X1 port map( A1 => n22349, A2 => n22689, ZN => n22350);
   U23088 : INV_X1 port map( A => n23933, ZN => n23918);
   U23089 : AOI21_X1 port map( B1 => n22356, B2 => n22355, A => n245, ZN => 
                           n22357);
   U23090 : INV_X1 port map( A => n22357, ZN => n22362);
   U23091 : INV_X1 port map( A => n23940, ZN => n23934);
   U23092 : INV_X1 port map( A => n22656, ZN => n22810);
   U23093 : MUX2_X1 port map( A => n23918, B => n23934, S => n23926, Z => 
                           n22381);
   U23094 : NAND2_X1 port map( A1 => n22670, A2 => n25023, ZN => n22364);
   U23095 : NAND2_X1 port map( A1 => n24963, A2 => n25023, ZN => n22366);
   U23096 : AOI21_X1 port map( B1 => n22366, B2 => n22670, A => n22779, ZN => 
                           n22367);
   U23097 : OR2_X2 port map( A1 => n22368, A2 => n22367, ZN => n23924);
   U23098 : INV_X1 port map( A => n23924, ZN => n23938);
   U23099 : MUX2_X1 port map( A => n22679, B => n22369, S => n22774, Z => 
                           n22372);
   U23101 : NAND2_X1 port map( A1 => n22376, A2 => n25439, ZN => n22375);
   U23102 : NAND2_X1 port map( A1 => n22373, A2 => n25414, ZN => n22374);
   U23103 : OAI211_X1 port map( C1 => n22376, C2 => n22677, A => n22375, B => 
                           n22374, ZN => n22378);
   U23104 : NAND3_X1 port map( A1 => n23997, A2 => n25439, A3 => n25079, ZN => 
                           n22377);
   U23105 : AOI21_X1 port map( B1 => n23939, B2 => n23926, A => n23924, ZN => 
                           n22379);
   U23106 : OAI21_X1 port map( B1 => n24948, B2 => n23937, A => n22379, ZN => 
                           n22380);
   U23107 : OAI21_X1 port map( B1 => n22381, B2 => n23938, A => n22380, ZN => 
                           n22383);
   U23108 : XNOR2_X1 port map( A => n22383, B => n22382, ZN => Ciphertext(176))
                           ;
   U23109 : XNOR2_X1 port map( A => n22386, B => n22385, ZN => Ciphertext(62));
   U23111 : NOR2_X1 port map( A1 => n22387, A2 => n22975, ZN => n22391);
   U23112 : NOR2_X1 port map( A1 => n22388, A2 => n22977, ZN => n22390);
   U23113 : NOR2_X1 port map( A1 => n22397, A2 => n22396, ZN => n22399);
   U23114 : NOR2_X1 port map( A1 => n22399, A2 => n25381, ZN => n22403);
   U23117 : NOR2_X1 port map( A1 => n1593, A2 => n22407, ZN => n22408);
   U23118 : NOR2_X1 port map( A1 => n22562, A2 => n22409, ZN => n22410);
   U23119 : AOI21_X1 port map( B1 => n22412, B2 => n22411, A => n22410, ZN => 
                           n22413);
   U23120 : NOR2_X1 port map( A1 => n23293, A2 => n23305, ZN => n22415);
   U23121 : MUX2_X1 port map( A => n22969, B => n22966, S => n21476, Z => 
                           n22419);
   U23122 : NAND2_X1 port map( A1 => n22962, A2 => n22965, ZN => n22417);
   U23124 : MUX2_X1 port map( A => n22417, B => n22416, S => n22966, Z => 
                           n22418);
   U23125 : OAI21_X1 port map( B1 => n22419, B2 => n22962, A => n22418, ZN => 
                           n23297);
   U23126 : INV_X1 port map( A => n23297, ZN => n23308);
   U23129 : INV_X1 port map( A => n23285, ZN => n22509);
   U23130 : NAND3_X1 port map( A1 => n22510, A2 => n22509, A3 => n23293, ZN => 
                           n22427);
   U23131 : OAI21_X1 port map( B1 => n23309, B2 => n23298, A => n22427, ZN => 
                           n22429);
   U23132 : INV_X1 port map( A => n2726, ZN => n22428);
   U23133 : XNOR2_X1 port map( A => n22429, B => n22428, ZN => Ciphertext(55));
   U23134 : NOR2_X1 port map( A1 => n23371, A2 => n22987, ZN => n23375);
   U23135 : INV_X1 port map( A => n22987, ZN => n23368);
   U23136 : INV_X1 port map( A => n22431, ZN => n22434);
   U23137 : INV_X1 port map( A => n22432, ZN => n22433);
   U23138 : OAI211_X1 port map( C1 => n22436, C2 => n22435, A => n22434, B => 
                           n22433, ZN => n22437);
   U23139 : OAI21_X1 port map( B1 => n24911, B2 => n24412, A => n22437, ZN => 
                           n22438);
   U23140 : NAND2_X1 port map( A1 => n22438, A2 => n4606, ZN => n22439);
   U23141 : NAND2_X1 port map( A1 => n24906, A2 => n23146, ZN => n22441);
   U23142 : OAI21_X1 port map( B1 => n24906, B2 => n22442, A => n22441, ZN => 
                           n22446);
   U23143 : NOR2_X1 port map( A1 => n23155, A2 => n24473, ZN => n22443);
   U23144 : NAND2_X1 port map( A1 => n22443, A2 => n24325, ZN => n22444);
   U23146 : XNOR2_X1 port map( A => n22447, B => n886, ZN => Ciphertext(22));
   U23148 : MUX2_X1 port map( A => n25450, B => n24367, S => n22459, Z => 
                           n22466);
   U23149 : INV_X1 port map( A => n23125, ZN => n23094);
   U23151 : INV_X1 port map( A => n25462, ZN => n22603);
   U23152 : NAND3_X1 port map( A1 => n25068, A2 => n22603, A3 => n24963, ZN => 
                           n22471);
   U23154 : NOR2_X1 port map( A1 => n24963, A2 => n24607, ZN => n22468);
   U23155 : NAND2_X1 port map( A1 => n22675, A2 => n22780, ZN => n22469);
   U23156 : AOI21_X1 port map( B1 => n24941, B2 => n23094, A => n5036, ZN => 
                           n22480);
   U23157 : NOR2_X1 port map( A1 => n22792, A2 => n22619, ZN => n22623);
   U23158 : NOR2_X1 port map( A1 => n22623, A2 => n22472, ZN => n22473);
   U23159 : INV_X1 port map( A => n23104, ZN => n23110);
   U23161 : INV_X1 port map( A => n23112, ZN => n23122);
   U23162 : MUX2_X1 port map( A => n22475, B => n22804, S => n25115, Z => 
                           n22477);
   U23164 : NOR2_X1 port map( A1 => n23122, A2 => n24059, ZN => n22478);
   U23165 : OAI21_X1 port map( B1 => n23093, B2 => n22478, A => n23125, ZN => 
                           n22479);
   U23166 : NAND2_X1 port map( A1 => n22482, A2 => n22842, ZN => n22486);
   U23167 : INV_X1 port map( A => n22900, ZN => n22847);
   U23168 : NOR2_X1 port map( A1 => n22905, A2 => n22904, ZN => n22721);
   U23169 : NAND2_X1 port map( A1 => n22906, A2 => n22721, ZN => n22485);
   U23170 : NAND3_X1 port map( A1 => n22837, A2 => n25041, A3 => n22893, ZN => 
                           n22487);
   U23171 : INV_X1 port map( A => n22835, ZN => n22894);
   U23172 : NOR2_X1 port map( A1 => n22897, A2 => n22894, ZN => n22488);
   U23173 : NOR2_X1 port map( A1 => n3176, A2 => n23458, ZN => n22490);
   U23174 : NAND2_X1 port map( A1 => n23464, A2 => n23016, ZN => n22492);
   U23175 : INV_X1 port map( A => n23015, ZN => n22864);
   U23176 : AOI21_X1 port map( B1 => n22492, B2 => n22914, A => n22864, ZN => 
                           n22493);
   U23177 : AOI21_X1 port map( B1 => n327, B2 => n22889, A => n22728, ZN => 
                           n22495);
   U23178 : AOI21_X1 port map( B1 => n22496, B2 => n22887, A => n3837, ZN => 
                           n22497);
   U23179 : NAND2_X1 port map( A1 => n23332, A2 => n22932, ZN => n22856);
   U23180 : NAND2_X1 port map( A1 => n22856, A2 => n22498, ZN => n22504);
   U23181 : AND2_X1 port map( A1 => n24342, A2 => n22499, ZN => n22500);
   U23182 : NOR2_X1 port map( A1 => n22855, A2 => n22500, ZN => n22503);
   U23183 : NAND2_X1 port map( A1 => n22501, A2 => n24356, ZN => n22502);
   U23184 : NOR2_X1 port map( A1 => n22938, A2 => n22832, ZN => n22505);
   U23185 : XNOR2_X1 port map( A => n22507, B => n16574, ZN => Ciphertext(92));
   U23186 : NOR2_X1 port map( A1 => n23292, A2 => n23305, ZN => n22763);
   U23187 : NOR2_X1 port map( A1 => n24904, A2 => n22509, ZN => n23306);
   U23188 : INV_X1 port map( A => n23181, ZN => n22513);
   U23189 : INV_X1 port map( A => n23165, ZN => n23179);
   U23190 : NAND3_X1 port map( A1 => n22513, A2 => n23166, A3 => n23179, ZN => 
                           n22517);
   U23191 : INV_X1 port map( A => n23166, ZN => n22551);
   U23192 : NAND3_X1 port map( A1 => n25488, A2 => n23164, A3 => n22551, ZN => 
                           n22516);
   U23193 : INV_X1 port map( A => n23178, ZN => n23167);
   U23194 : INV_X1 port map( A => n23164, ZN => n23176);
   U23195 : NAND3_X1 port map( A1 => n23165, A2 => n23167, A3 => n23176, ZN => 
                           n22515);
   U23196 : NAND3_X1 port map( A1 => n23168, A2 => n23164, A3 => n23165, ZN => 
                           n22514);
   U23197 : NAND4_X1 port map( A1 => n22517, A2 => n22516, A3 => n22515, A4 => 
                           n22514, ZN => n22519);
   U23198 : INV_X1 port map( A => n812, ZN => n22518);
   U23199 : XNOR2_X1 port map( A => n22519, B => n22518, ZN => Ciphertext(28));
   U23200 : INV_X1 port map( A => n23770, ZN => n23781);
   U23201 : AOI22_X1 port map( A1 => n23778, A2 => n23768, B1 => n23781, B2 => 
                           n24921, ZN => n23783);
   U23202 : NAND2_X1 port map( A1 => n25051, A2 => n23757, ZN => n23758);
   U23203 : INV_X1 port map( A => n23758, ZN => n22523);
   U23204 : XNOR2_X1 port map( A => n22526, B => n22525, ZN => Ciphertext(145))
                           ;
   U23205 : NAND2_X1 port map( A1 => n25042, A2 => n1370, ZN => n23437);
   U23206 : INV_X1 port map( A => n23865, ZN => n23853);
   U23207 : AOI21_X1 port map( B1 => n22982, B2 => n23857, A => n23853, ZN => 
                           n22533);
   U23208 : NOR3_X1 port map( A1 => n23860, A2 => n23862, A3 => n25399, ZN => 
                           n22532);
   U23209 : NOR3_X1 port map( A1 => n23858, A2 => n25399, A3 => n23865, ZN => 
                           n22531);
   U23210 : XNOR2_X1 port map( A => n22534, B => n1726, ZN => Ciphertext(162));
   U23211 : INV_X1 port map( A => n23275, ZN => n23278);
   U23212 : XNOR2_X1 port map( A => n22538, B => n2757, ZN => Ciphertext(50));
   U23213 : INV_X1 port map( A => n22539, ZN => n23813);
   U23214 : NOR2_X1 port map( A1 => n23813, A2 => n23030, ZN => n23833);
   U23215 : AND2_X1 port map( A1 => n22539, A2 => n23828, ZN => n23818);
   U23216 : NAND2_X1 port map( A1 => n23818, A2 => n25391, ZN => n22541);
   U23217 : INV_X1 port map( A => n2193, ZN => n22542);
   U23218 : XNOR2_X1 port map( A => n22543, B => n22542, ZN => Ciphertext(156))
                           ;
   U23219 : NOR2_X1 port map( A1 => n23904, A2 => n21863, ZN => n22545);
   U23220 : INV_X1 port map( A => n23906, ZN => n22544);
   U23221 : OAI21_X1 port map( B1 => n23888, B2 => n22545, A => n22544, ZN => 
                           n22548);
   U23222 : INV_X1 port map( A => n23890, ZN => n22546);
   U23223 : XNOR2_X1 port map( A => n22550, B => n22549, ZN => Ciphertext(168))
                           ;
   U23224 : NAND3_X1 port map( A1 => n23168, A2 => n23176, A3 => n23166, ZN => 
                           n22554);
   U23225 : XNOR2_X1 port map( A => n22557, B => n22556, ZN => Ciphertext(27));
   U23226 : INV_X1 port map( A => n23743, ZN => n22558);
   U23227 : OAI21_X1 port map( B1 => n23740, B2 => n24065, A => n22558, ZN => 
                           n22559);
   U23228 : OAI22_X1 port map( A1 => n23743, A2 => n23740, B1 => n24991, B2 => 
                           n23748, ZN => n23735);
   U23229 : INV_X1 port map( A => n23730, ZN => n23745);
   U23230 : AOI22_X1 port map( A1 => n23748, A2 => n22559, B1 => n23735, B2 => 
                           n23745, ZN => n22560);
   U23231 : XNOR2_X1 port map( A => n22560, B => n4164, ZN => Ciphertext(143));
   U23232 : NAND2_X1 port map( A1 => n24971, A2 => n22563, ZN => n22565);
   U23233 : OAI22_X1 port map( A1 => n22568, A2 => n22567, B1 => n24951, B2 => 
                           n22565, ZN => n22570);
   U23234 : OAI21_X1 port map( B1 => n22571, B2 => n22570, A => n22569, ZN => 
                           n22572);
   U23235 : NOR2_X1 port map( A1 => n22573, A2 => n22572, ZN => n22574);
   U23236 : NOR2_X1 port map( A1 => n23184, A2 => n22575, ZN => n23203);
   U23237 : MUX2_X1 port map( A => n22574, B => n23203, S => n24334, Z => 
                           n22576);
   U23238 : INV_X1 port map( A => n23200, ZN => n22824);
   U23239 : INV_X1 port map( A => n23201, ZN => n22820);
   U23240 : INV_X1 port map( A => n22578, ZN => n23069);
   U23242 : INV_X1 port map( A => n23064, ZN => n22580);
   U23244 : INV_X1 port map( A => n22872, ZN => n22579);
   U23245 : OAI21_X1 port map( B1 => n22580, B2 => n23077, A => n22579, ZN => 
                           n22581);
   U23246 : NOR2_X1 port map( A1 => n22803, A2 => n22805, ZN => n22582);
   U23248 : NAND2_X1 port map( A1 => n22585, A2 => n22584, ZN => n22587);
   U23249 : NAND2_X1 port map( A1 => n22798, A2 => n24561, ZN => n22586);
   U23250 : NOR2_X2 port map( A1 => n22589, A2 => n22588, ZN => n23052);
   U23251 : OAI21_X1 port map( B1 => n22591, B2 => n22590, A => n22448, ZN => 
                           n22595);
   U23252 : OAI211_X1 port map( C1 => n23997, C2 => n22677, A => n24439, B => 
                           n22596, ZN => n22597);
   U23253 : OAI21_X1 port map( B1 => n22598, B2 => n22676, A => n22597, ZN => 
                           n23047);
   U23254 : MUX2_X1 port map( A => n23052, B => n23040, S => n23047, Z => 
                           n22624);
   U23255 : NAND2_X1 port map( A1 => n24963, A2 => n22779, ZN => n22600);
   U23256 : OAI21_X1 port map( B1 => n22675, B2 => n22779, A => n22600, ZN => 
                           n22601);
   U23257 : INV_X1 port map( A => n22601, ZN => n22605);
   U23258 : MUX2_X1 port map( A => n22670, B => n25022, S => n24963, Z => 
                           n22602);
   U23259 : INV_X1 port map( A => n22602, ZN => n22604);
   U23260 : INV_X1 port map( A => n23050, ZN => n23058);
   U23261 : NOR2_X1 port map( A1 => n22813, A2 => n25241, ZN => n22608);
   U23262 : NOR3_X1 port map( A1 => n22813, A2 => n22606, A3 => n25075, ZN => 
                           n22607);
   U23263 : AOI21_X1 port map( B1 => n22656, B2 => n22608, A => n22607, ZN => 
                           n22611);
   U23265 : NAND2_X1 port map( A1 => n22792, A2 => n22612, ZN => n22613);
   U23266 : NAND2_X1 port map( A1 => n22613, A2 => n22617, ZN => n22622);
   U23267 : NOR2_X1 port map( A1 => n22615, A2 => n22614, ZN => n22616);
   U23268 : NAND2_X1 port map( A1 => n24953, A2 => n22616, ZN => n22621);
   U23269 : NAND2_X1 port map( A1 => n22619, A2 => n22618, ZN => n22620);
   U23270 : OAI211_X1 port map( C1 => n22623, C2 => n22622, A => n22620, B => 
                           n22621, ZN => n22698);
   U23271 : XNOR2_X1 port map( A => n22626, B => n22625, ZN => Ciphertext(3));
   U23272 : OAI22_X1 port map( A1 => n23318, A2 => n23326, B1 => n23327, B2 => 
                           n23320, ZN => n23325);
   U23273 : NAND2_X1 port map( A1 => n23318, A2 => n23313, ZN => n22627);
   U23274 : AOI22_X1 port map( A1 => n22629, A2 => n23325, B1 => n22628, B2 => 
                           n22627, ZN => n22630);
   U23275 : XNOR2_X1 port map( A => n22630, B => n2826, ZN => Ciphertext(61));
   U23276 : NAND2_X1 port map( A1 => n24390, A2 => n23592, ZN => n22631);
   U23277 : AOI21_X1 port map( B1 => n22632, B2 => n22631, A => n23591, ZN => 
                           n22642);
   U23278 : INV_X1 port map( A => n23594, ZN => n23565);
   U23279 : AND2_X1 port map( A1 => n23592, A2 => n23565, ZN => n22637);
   U23280 : AOI21_X1 port map( B1 => n22637, B2 => n23591, A => n22635, ZN => 
                           n22636);
   U23281 : AOI21_X1 port map( B1 => n21941, B2 => n24389, A => n2040, ZN => 
                           n22638);
   U23282 : INV_X1 port map( A => n23047, ZN => n23053);
   U23283 : NOR2_X1 port map( A1 => n23052, A2 => n23053, ZN => n23060);
   U23284 : INV_X1 port map( A => n23052, ZN => n23042);
   U23285 : INV_X1 port map( A => n23040, ZN => n23049);
   U23286 : OAI21_X1 port map( B1 => n23042, B2 => n23059, A => n23049, ZN => 
                           n22646);
   U23287 : NAND2_X1 port map( A1 => n22643, A2 => n23050, ZN => n22645);
   U23288 : OAI211_X1 port map( C1 => n23060, C2 => n22646, A => n22645, B => 
                           n22644, ZN => n22647);
   U23289 : XNOR2_X1 port map( A => n22647, B => n3073, ZN => Ciphertext(2));
   U23291 : INV_X1 port map( A => n23252, ZN => n23236);
   U23292 : AOI22_X1 port map( A1 => n22650, A2 => n22649, B1 => n22648, B2 => 
                           n23256, ZN => n22651);
   U23293 : XNOR2_X1 port map( A => n22651, B => n663, ZN => Ciphertext(46));
   U23294 : MUX2_X1 port map( A => n23227, B => n23228, S => n24955, Z => 
                           n22653);
   U23296 : XNOR2_X1 port map( A => n22654, B => n1863, ZN => Ciphertext(38));
   U23297 : NOR2_X1 port map( A1 => n22804, A2 => n22805, ZN => n22802);
   U23298 : AND2_X1 port map( A1 => n22798, A2 => n22803, ZN => n22661);
   U23300 : NOR2_X1 port map( A1 => n22800, A2 => n24559, ZN => n22663);
   U23301 : NAND2_X1 port map( A1 => n22663, A2 => n22804, ZN => n22664);
   U23302 : NAND2_X1 port map( A1 => n22779, A2 => n25462, ZN => n22674);
   U23303 : NAND2_X1 port map( A1 => n24963, A2 => n22782, ZN => n22669);
   U23304 : INV_X1 port map( A => n22667, ZN => n22783);
   U23305 : NOR2_X1 port map( A1 => n22779, A2 => n25023, ZN => n22671);
   U23306 : INV_X1 port map( A => n23958, ZN => n23952);
   U23307 : NOR2_X1 port map( A1 => n23969, A2 => n23952, ZN => n23970);
   U23308 : INV_X1 port map( A => n23970, ZN => n22696);
   U23309 : NAND3_X1 port map( A1 => n22771, A2 => n22680, A3 => n22769, ZN => 
                           n22681);
   U23313 : AOI22_X1 port map( A1 => n21848, A2 => n22687, B1 => n22686, B2 => 
                           n22685, ZN => n22692);
   U23314 : OAI21_X1 port map( B1 => n22690, B2 => n22689, A => n22688, ZN => 
                           n22691);
   U23315 : OAI21_X1 port map( B1 => n22692, B2 => n25395, A => n22691, ZN => 
                           n23966);
   U23316 : NAND2_X1 port map( A1 => n22693, A2 => n23966, ZN => n22694);
   U23317 : AND2_X1 port map( A1 => n23966, A2 => n24910, ZN => n23953);
   U23318 : AOI22_X1 port map( A1 => n25076, A2 => n22694, B1 => n23953, B2 => 
                           n25017, ZN => n22695);
   U23319 : NAND2_X1 port map( A1 => n23040, A2 => n22698, ZN => n22699);
   U23320 : INV_X1 port map( A => n23537, ZN => n23557);
   U23321 : OAI21_X1 port map( B1 => n25071, B2 => n23555, A => n24893, ZN => 
                           n22700);
   U23322 : AOI22_X1 port map( A1 => n22701, A2 => n23557, B1 => n23554, B2 => 
                           n22700, ZN => n22703);
   U23323 : XNOR2_X1 port map( A => n22703, B => n22702, ZN => Ciphertext(113))
                           ;
   U23326 : INV_X1 port map( A => n23259, ZN => n23282);
   U23327 : INV_X1 port map( A => n23281, ZN => n23267);
   U23328 : OR2_X1 port map( A1 => n23277, A2 => n24349, ZN => n22705);
   U23329 : OAI22_X1 port map( A1 => n23282, A2 => n24360, B1 => n23267, B2 => 
                           n22705, ZN => n22708);
   U23330 : NOR2_X1 port map( A1 => n23277, A2 => n23273, ZN => n22706);
   U23331 : NOR2_X1 port map( A1 => n22708, A2 => n22707, ZN => n22709);
   U23332 : XNOR2_X1 port map( A => n22709, B => n673, ZN => Ciphertext(48));
   U23333 : MUX2_X1 port map( A => n23546, B => n23537, S => n23554, Z => 
                           n22710);
   U23334 : INV_X1 port map( A => n22711, ZN => n22716);
   U23335 : NOR2_X1 port map( A1 => n22712, A2 => n22928, ZN => n22713);
   U23336 : OAI21_X1 port map( B1 => n22713, B2 => n22107, A => n22926, ZN => 
                           n22714);
   U23337 : INV_X1 port map( A => n23479, ZN => n23483);
   U23338 : MUX2_X1 port map( A => n22717, B => n22841, S => n25041, Z => 
                           n22720);
   U23339 : INV_X1 port map( A => n25041, ZN => n22718);
   U23340 : MUX2_X1 port map( A => n22718, B => n22835, S => n25438, Z => 
                           n22719);
   U23341 : NAND2_X1 port map( A1 => n24932, A2 => n22832, ZN => n22724);
   U23342 : INV_X1 port map( A => n22939, ZN => n22723);
   U23343 : NAND2_X1 port map( A1 => n22938, A2 => n22832, ZN => n22935);
   U23344 : AOI21_X1 port map( B1 => n22935, B2 => n22829, A => n22723, ZN => 
                           n22725);
   U23346 : NOR2_X1 port map( A1 => n23491, A2 => n23481, ZN => n23495);
   U23348 : MUX2_X1 port map( A => n22889, B => n22727, S => n22890, Z => 
                           n22732);
   U23349 : NOR2_X1 port map( A1 => n22729, A2 => n22890, ZN => n22731);
   U23350 : NOR2_X1 port map( A1 => n23464, A2 => n23458, ZN => n22734);
   U23351 : INV_X1 port map( A => n23464, ZN => n22733);
   U23352 : INV_X1 port map( A => n22911, ZN => n23462);
   U23353 : AND3_X1 port map( A1 => n22864, A2 => n23016, A3 => n23014, ZN => 
                           n23467);
   U23354 : AOI21_X1 port map( B1 => n22734, B2 => n23460, A => n23467, ZN => 
                           n22735);
   U23355 : NAND3_X1 port map( A1 => n22736, A2 => n23492, A3 => n24442, ZN => 
                           n22737);
   U23357 : XNOR2_X1 port map( A => n22740, B => n22739, ZN => Ciphertext(97));
   U23358 : NAND2_X1 port map( A1 => n22988, A2 => n23374, ZN => n22743);
   U23359 : NAND2_X1 port map( A1 => n22741, A2 => n24515, ZN => n22989);
   U23360 : OAI211_X1 port map( C1 => n22741, C2 => n23368, A => n23379, B => 
                           n22989, ZN => n22742);
   U23361 : XNOR2_X1 port map( A => n22746, B => n22745, ZN => Ciphertext(75));
   U23362 : INV_X1 port map( A => n23670, ZN => n22749);
   U23363 : INV_X1 port map( A => n23689, ZN => n22747);
   U23364 : NAND2_X1 port map( A1 => n22747, A2 => n23690, ZN => n23659);
   U23365 : OAI21_X1 port map( B1 => n22749, B2 => n23692, A => n23659, ZN => 
                           n22750);
   U23366 : NAND2_X1 port map( A1 => n23676, A2 => n23690, ZN => n22748);
   U23369 : INV_X1 port map( A => n22752, ZN => n23193);
   U23370 : NAND2_X1 port map( A1 => n23193, A2 => n23206, ZN => n22754);
   U23371 : NAND2_X1 port map( A1 => n23201, A2 => n23184, ZN => n22753);
   U23372 : OAI21_X1 port map( B1 => n22754, B2 => n23196, A => n22753, ZN => 
                           n22821);
   U23373 : AOI21_X1 port map( B1 => n24334, B2 => n25059, A => n5769, ZN => 
                           n22756);
   U23374 : NAND2_X1 port map( A1 => n5769, A2 => n23206, ZN => n22755);
   U23375 : OAI22_X1 port map( A1 => n22821, A2 => n22756, B1 => n22755, B2 => 
                           n23200, ZN => n22757);
   U23376 : XNOR2_X1 port map( A => n22757, B => n2222, ZN => Ciphertext(31));
   U23377 : MUX2_X1 port map( A => n23178, B => n23164, S => n25488, Z => 
                           n22759);
   U23378 : AOI21_X1 port map( B1 => n23181, B2 => n23179, A => n23166, ZN => 
                           n22758);
   U23379 : OAI22_X1 port map( A1 => n22759, A2 => n22758, B1 => n23181, B2 => 
                           n24394, ZN => n22760);
   U23380 : XNOR2_X1 port map( A => n22760, B => n1952, ZN => Ciphertext(24));
   U23381 : INV_X1 port map( A => n24904, ZN => n23299);
   U23382 : BUF_X1 port map( A => n23285, Z => n23294);
   U23383 : OAI21_X1 port map( B1 => n23293, B2 => n22762, A => n22761, ZN => 
                           n22766);
   U23384 : AND2_X1 port map( A1 => n23297, A2 => n23292, ZN => n22764);
   U23385 : AOI22_X1 port map( A1 => n22763, A2 => n23294, B1 => n22764, B2 => 
                           n23303, ZN => n22765);
   U23386 : OAI21_X1 port map( B1 => n22766, B2 => n23303, A => n22765, ZN => 
                           n22768);
   U23387 : XNOR2_X1 port map( A => n22768, B => n22767, ZN => Ciphertext(58));
   U23388 : MUX2_X1 port map( A => n25414, B => n23998, S => n24439, Z => 
                           n22776);
   U23391 : NAND2_X1 port map( A1 => n25068, A2 => n22780, ZN => n22786);
   U23392 : NAND3_X1 port map( A1 => n22784, A2 => n22783, A3 => n25462, ZN => 
                           n22785);
   U23394 : NAND2_X1 port map( A1 => n22788, A2 => n24953, ZN => n22797);
   U23395 : NAND2_X1 port map( A1 => n22790, A2 => n22789, ZN => n22796);
   U23397 : NAND2_X1 port map( A1 => n24006, A2 => n24010, ZN => n23984);
   U23399 : NOR2_X1 port map( A1 => n22800, A2 => n25115, ZN => n22801);
   U23400 : AOI22_X1 port map( A1 => n22802, A2 => n22584, B1 => n22801, B2 => 
                           n22804, ZN => n22808);
   U23401 : NOR2_X1 port map( A1 => n22804, A2 => n22803, ZN => n22807);
   U23402 : NOR2_X1 port map( A1 => n22810, A2 => n25241, ZN => n22816);
   U23403 : NOR2_X1 port map( A1 => n22812, A2 => n22811, ZN => n22815);
   U23404 : OAI21_X1 port map( B1 => n22813, B2 => n22812, A => n1477, ZN => 
                           n22814);
   U23407 : OAI21_X1 port map( B1 => n22820, B2 => n23202, A => n24889, ZN => 
                           n22823);
   U23408 : INV_X1 port map( A => n23186, ZN => n22822);
   U23409 : AOI22_X1 port map( A1 => n22824, A2 => n22823, B1 => n22822, B2 => 
                           n22821, ZN => n22825);
   U23410 : XNOR2_X1 port map( A => n22825, B => n1856, ZN => Ciphertext(35));
   U23411 : INV_X1 port map( A => n24910, ZN => n23964);
   U23412 : INV_X1 port map( A => n23967, ZN => n23947);
   U23413 : MUX2_X1 port map( A => n23964, B => n23947, S => n23966, Z => 
                           n22828);
   U23414 : NOR2_X1 port map( A1 => n22939, A2 => n22829, ZN => n22830);
   U23415 : MUX2_X1 port map( A => n22834, B => n25438, S => n25041, Z => 
                           n22840);
   U23419 : NOR2_X1 port map( A1 => n142, A2 => n25035, ZN => n22851);
   U23421 : INV_X1 port map( A => n22033, ZN => n22859);
   U23422 : OAI21_X1 port map( B1 => n22958, B2 => n22959, A => n22859, ZN => 
                           n22860);
   U23423 : AND2_X1 port map( A1 => n22860, A2 => n4128, ZN => n22861);
   U23425 : XNOR2_X1 port map( A => n22867, B => n2049, ZN => Ciphertext(86));
   U23426 : INV_X1 port map( A => n23403, ZN => n23418);
   U23427 : XNOR2_X1 port map( A => n22870, B => n1896, ZN => Ciphertext(87));
   U23429 : NOR2_X1 port map( A1 => n24075, A2 => n23064, ZN => n23076);
   U23431 : NAND3_X1 port map( A1 => n23064, A2 => n23074, A3 => n23066, ZN => 
                           n22873);
   U23434 : AOI21_X1 port map( B1 => n25179, B2 => n25452, A => n23064, ZN => 
                           n22878);
   U23435 : NAND2_X1 port map( A1 => n23074, A2 => n23066, ZN => n22877);
   U23436 : AOI22_X1 port map( A1 => n22879, A2 => n23064, B1 => n22878, B2 => 
                           n22877, ZN => n22880);
   U23437 : XNOR2_X1 port map( A => n22880, B => n2746, ZN => Ciphertext(8));
   U23438 : NAND2_X1 port map( A1 => n23394, A2 => n24933, ZN => n22881);
   U23439 : NAND2_X1 port map( A1 => n22881, A2 => n23396, ZN => n22883);
   U23440 : AND3_X1 port map( A1 => n23394, A2 => n23396, A3 => n23393, ZN => 
                           n22882);
   U23441 : NOR2_X1 port map( A1 => n25375, A2 => n22887, ZN => n22892);
   U23442 : NOR2_X1 port map( A1 => n22729, A2 => n22889, ZN => n22891);
   U23443 : MUX2_X1 port map( A => n22892, B => n22891, S => n22890, Z => 
                           n23514);
   U23444 : NAND2_X1 port map( A1 => n22894, A2 => n22893, ZN => n22899);
   U23445 : INV_X1 port map( A => n22895, ZN => n22898);
   U23446 : AOI22_X1 port map( A1 => n22899, A2 => n22898, B1 => n22897, B2 => 
                           n22896, ZN => n22915);
   U23447 : OR2_X1 port map( A1 => n24380, A2 => n23510, ZN => n23013);
   U23448 : AND2_X1 port map( A1 => n22900, A2 => n22901, ZN => n22902);
   U23449 : NOR2_X1 port map( A1 => n22903, A2 => n22902, ZN => n22910);
   U23450 : OAI21_X1 port map( B1 => n22906, B2 => n22905, A => n22904, ZN => 
                           n22909);
   U23452 : MUX2_X1 port map( A => n23016, B => n22911, S => n23464, Z => 
                           n22913);
   U23453 : NAND2_X1 port map( A1 => n23016, A2 => n3176, ZN => n22912);
   U23454 : OR2_X1 port map( A1 => n22914, A2 => n24364, ZN => n23018);
   U23455 : INV_X1 port map( A => n22915, ZN => n23530);
   U23456 : NAND2_X1 port map( A1 => n23530, A2 => n23529, ZN => n22921);
   U23458 : XNOR2_X1 port map( A => n22930, B => n2120, ZN => Ciphertext(107));
   U23459 : NOR2_X1 port map( A1 => n24309, A2 => n23334, ZN => n22931);
   U23460 : AOI21_X1 port map( B1 => n22936, B2 => n22935, A => n22934, ZN => 
                           n22943);
   U23462 : NAND2_X1 port map( A1 => n23361, A2 => n24492, ZN => n22979);
   U23464 : INV_X1 port map( A => n22945, ZN => n22950);
   U23466 : NOR2_X1 port map( A1 => n22033, A2 => n22953, ZN => n22955);
   U23467 : MUX2_X1 port map( A => n22958, B => n24922, S => n24884, Z => 
                           n22960);
   U23468 : INV_X1 port map( A => n22962, ZN => n22963);
   U23469 : OAI21_X1 port map( B1 => n22965, B2 => n21476, A => n22964, ZN => 
                           n22971);
   U23470 : OAI22_X1 port map( A1 => n22387, A2 => n22974, B1 => n22977, B2 => 
                           n22973, ZN => n22976);
   U23471 : AOI22_X2 port map( A1 => n22978, A2 => n22977, B1 => n22976, B2 => 
                           n25365, ZN => n23359);
   U23472 : XNOR2_X1 port map( A => n22980, B => n1768, ZN => Ciphertext(67));
   U23475 : INV_X1 port map( A => n22989, ZN => n22990);
   U23476 : AOI22_X1 port map( A1 => n22993, A2 => n22992, B1 => n22991, B2 => 
                           n22990, ZN => n22994);
   U23477 : XNOR2_X1 port map( A => n22994, B => n1792, ZN => Ciphertext(73));
   U23478 : INV_X1 port map( A => n23350, ZN => n23340);
   U23479 : NAND3_X1 port map( A1 => n22961, A2 => n24492, A3 => n23359, ZN => 
                           n22995);
   U23480 : NAND2_X1 port map( A1 => n23670, A2 => n23692, ZN => n22997);
   U23481 : NOR2_X1 port map( A1 => n22997, A2 => n23658, ZN => n23000);
   U23482 : NOR2_X1 port map( A1 => n22998, A2 => n23692, ZN => n22999);
   U23483 : NAND2_X1 port map( A1 => n23805, A2 => n23786, ZN => n23005);
   U23484 : INV_X1 port map( A => n24392, ZN => n23796);
   U23485 : OAI21_X1 port map( B1 => n21837, B2 => n23002, A => n23796, ZN => 
                           n23003);
   U23486 : XNOR2_X1 port map( A => n23006, B => n2782, ZN => Ciphertext(155));
   U23487 : AOI21_X1 port map( B1 => n23525, B2 => n24351, A => n23530, ZN => 
                           n23007);
   U23488 : AOI22_X1 port map( A1 => n23009, A2 => n23008, B1 => n23527, B2 => 
                           n23007, ZN => n23010);
   U23489 : XNOR2_X1 port map( A => n23010, B => n2042, ZN => Ciphertext(103));
   U23490 : INV_X1 port map( A => n23470, ZN => n23011);
   U23491 : XNOR2_X1 port map( A => n23012, B => n2050, ZN => Ciphertext(100));
   U23492 : NAND2_X1 port map( A1 => n24380, A2 => n23529, ZN => n23533);
   U23493 : OAI21_X1 port map( B1 => n25055, B2 => n23460, A => n23014, ZN => 
                           n23019);
   U23494 : NAND3_X1 port map( A1 => n23016, A2 => n23461, A3 => n3176, ZN => 
                           n23017);
   U23495 : OAI211_X1 port map( C1 => n24435, C2 => n23019, A => n23018, B => 
                           n23017, ZN => n23022);
   U23496 : NAND2_X1 port map( A1 => n23022, A2 => n23505, ZN => n23021);
   U23497 : OAI211_X1 port map( C1 => n23527, C2 => n23022, A => n24351, B => 
                           n23021, ZN => n23023);
   U23498 : NAND2_X1 port map( A1 => n23024, A2 => n23023, ZN => n23025);
   U23499 : XNOR2_X1 port map( A => n23025, B => n2100, ZN => Ciphertext(104));
   U23500 : NAND2_X1 port map( A1 => n23939, A2 => n23924, ZN => n23920);
   U23501 : NAND2_X1 port map( A1 => n25084, A2 => n23933, ZN => n23921);
   U23502 : NAND2_X1 port map( A1 => n23920, A2 => n23921, ZN => n23028);
   U23503 : INV_X1 port map( A => n24948, ZN => n23027);
   U23504 : OAI21_X1 port map( B1 => n23926, B2 => n23918, A => n25084, ZN => 
                           n23026);
   U23505 : AOI22_X1 port map( A1 => n23028, A2 => n23937, B1 => n23027, B2 => 
                           n23026, ZN => n23029);
   U23506 : XNOR2_X1 port map( A => n23029, B => n2989, ZN => Ciphertext(179));
   U23507 : NOR2_X1 port map( A1 => n23810, A2 => n23817, ZN => n23830);
   U23508 : INV_X1 port map( A => n23828, ZN => n23032);
   U23509 : AND2_X1 port map( A1 => n23828, A2 => n23030, ZN => n23031);
   U23510 : AOI21_X1 port map( B1 => n23810, B2 => n23032, A => n23031, ZN => 
                           n23033);
   U23511 : XNOR2_X1 port map( A => n23035, B => n2058, ZN => Ciphertext(158));
   U23512 : NOR3_X1 port map( A1 => n23361, A2 => n24492, A3 => n22961, ZN => 
                           n23036);
   U23513 : AOI211_X1 port map( C1 => n23361, C2 => n23037, A => n23355, B => 
                           n23036, ZN => n23038);
   U23514 : XNOR2_X1 port map( A => n23038, B => n2034, ZN => Ciphertext(66));
   U23516 : OAI21_X1 port map( B1 => n23039, B2 => n23055, A => n322, ZN => 
                           n23044);
   U23517 : OAI21_X1 port map( B1 => n322, B2 => n23040, A => n23059, ZN => 
                           n23041);
   U23518 : NAND2_X1 port map( A1 => n23042, A2 => n23041, ZN => n23043);
   U23519 : NAND2_X1 port map( A1 => n23044, A2 => n23043, ZN => n23046);
   U23520 : XNOR2_X1 port map( A => n23046, B => n23045, ZN => Ciphertext(0));
   U23521 : AOI22_X1 port map( A1 => n23050, A2 => n23049, B1 => n23048, B2 => 
                           n23047, ZN => n23062);
   U23522 : OAI21_X1 port map( B1 => n23062, B2 => n23055, A => n23054, ZN => 
                           n23057);
   U23523 : INV_X1 port map( A => n881, ZN => n23056);
   U23524 : XNOR2_X1 port map( A => n23057, B => n23056, ZN => Ciphertext(1));
   U23525 : OAI21_X1 port map( B1 => n23060, B2 => n23059, A => n23058, ZN => 
                           n23061);
   U23526 : INV_X1 port map( A => n681, ZN => n23063);
   U23527 : INV_X1 port map( A => n23074, ZN => n23079);
   U23528 : OAI21_X1 port map( B1 => n23076, B2 => n23079, A => n25179, ZN => 
                           n23071);
   U23529 : NOR2_X1 port map( A1 => n23064, A2 => n23077, ZN => n23068);
   U23530 : NOR2_X1 port map( A1 => n23077, A2 => n25452, ZN => n23067);
   U23531 : AOI22_X1 port map( A1 => n23069, A2 => n23068, B1 => n23067, B2 => 
                           n23066, ZN => n23070);
   U23533 : XNOR2_X1 port map( A => n23073, B => n23072, ZN => Ciphertext(6));
   U23534 : AOI21_X1 port map( B1 => n25179, B2 => n25024, A => n23074, ZN => 
                           n23082);
   U23535 : NAND2_X1 port map( A1 => n23076, A2 => n22578, ZN => n23081);
   U23536 : NAND3_X1 port map( A1 => n23079, A2 => n25024, A3 => n23077, ZN => 
                           n23080);
   U23537 : NOR2_X1 port map( A1 => n23119, A2 => n23120, ZN => n23085);
   U23538 : AOI21_X1 port map( B1 => n23123, B2 => n24941, A => n23085, ZN => 
                           n23126);
   U23539 : OAI211_X1 port map( C1 => n23094, C2 => n24941, A => n23112, B => 
                           n24993, ZN => n23086);
   U23540 : OAI21_X1 port map( B1 => n23126, B2 => n23093, A => n23086, ZN => 
                           n23088);
   U23541 : INV_X1 port map( A => n2241, ZN => n23087);
   U23542 : XNOR2_X1 port map( A => n23088, B => n23087, ZN => Ciphertext(13));
   U23543 : MUX2_X1 port map( A => n23112, B => n23125, S => n23104, Z => 
                           n23089);
   U23544 : NOR2_X1 port map( A1 => n24941, A2 => n5036, ZN => n23090);
   U23545 : NAND2_X1 port map( A1 => n23090, A2 => n23112, ZN => n23097);
   U23546 : NAND2_X1 port map( A1 => n24993, A2 => n23112, ZN => n23091);
   U23547 : NAND2_X1 port map( A1 => n23094, A2 => n23093, ZN => n23095);
   U23548 : NAND3_X1 port map( A1 => n23097, A2 => n23096, A3 => n23095, ZN => 
                           n23099);
   U23549 : INV_X1 port map( A => n2745, ZN => n23098);
   U23550 : XNOR2_X1 port map( A => n23099, B => n23098, ZN => Ciphertext(15));
   U23551 : NAND2_X1 port map( A1 => n23120, A2 => n859, ZN => n23102);
   U23552 : INV_X1 port map( A => n859, ZN => n23108);
   U23553 : NAND3_X1 port map( A1 => n24059, A2 => n23120, A3 => n23108, ZN => 
                           n23101);
   U23554 : NOR2_X1 port map( A1 => n23120, A2 => n859, ZN => n23113);
   U23555 : NAND2_X1 port map( A1 => n23112, A2 => n23113, ZN => n23100);
   U23556 : OAI211_X1 port map( C1 => n24059, C2 => n23102, A => n23101, B => 
                           n23100, ZN => n23106);
   U23557 : NAND3_X1 port map( A1 => n24498, A2 => n859, A3 => n5036, ZN => 
                           n23103);
   U23558 : NOR2_X1 port map( A1 => n23103, A2 => n23112, ZN => n23105);
   U23559 : OAI21_X1 port map( B1 => n23106, B2 => n23105, A => n23104, ZN => 
                           n23118);
   U23560 : XNOR2_X1 port map( A => n23125, B => n859, ZN => n23107);
   U23561 : NAND3_X1 port map( A1 => n23123, A2 => n24498, A3 => n23107, ZN => 
                           n23117);
   U23562 : NOR2_X1 port map( A1 => n24498, A2 => n23108, ZN => n23109);
   U23563 : OAI211_X1 port map( C1 => n23120, C2 => n23112, A => n23123, B => 
                           n23109, ZN => n23116);
   U23564 : NOR2_X1 port map( A1 => n23112, A2 => n24498, ZN => n23114);
   U23565 : NAND2_X1 port map( A1 => n23114, A2 => n23113, ZN => n23115);
   U23566 : NAND4_X1 port map( A1 => n23118, A2 => n23117, A3 => n23116, A4 => 
                           n23115, ZN => Ciphertext(16));
   U23567 : INV_X1 port map( A => n24993, ZN => n23121);
   U23568 : AOI21_X1 port map( B1 => n23122, B2 => n23121, A => n23120, ZN => 
                           n23124);
   U23569 : OAI22_X1 port map( A1 => n23126, A2 => n23125, B1 => n23124, B2 => 
                           n23123, ZN => n23128);
   U23570 : INV_X1 port map( A => n3093, ZN => n23127);
   U23571 : XNOR2_X1 port map( A => n23128, B => n23127, ZN => Ciphertext(17));
   U23572 : INV_X1 port map( A => n23157, ZN => n23131);
   U23573 : INV_X1 port map( A => n23154, ZN => n23139);
   U23575 : OAI21_X1 port map( B1 => n23133, B2 => n22442, A => n23132, ZN => 
                           n23134);
   U23576 : INV_X1 port map( A => n23134, ZN => n23136);
   U23577 : OAI21_X1 port map( B1 => n23160, B2 => n23155, A => n24906, ZN => 
                           n23135);
   U23578 : INV_X1 port map( A => n2761, ZN => n23137);
   U23579 : AND2_X1 port map( A1 => n24473, A2 => n23155, ZN => n23158);
   U23580 : NAND2_X1 port map( A1 => n23158, A2 => n23143, ZN => n23141);
   U23581 : OAI211_X1 port map( C1 => n23146, C2 => n1349, A => n23139, B => 
                           n23138, ZN => n23140);
   U23582 : OAI211_X1 port map( C1 => n24325, C2 => n23143, A => n23141, B => 
                           n23140, ZN => n23142);
   U23583 : XNOR2_X1 port map( A => n23142, B => n1528, ZN => Ciphertext(19));
   U23584 : OAI21_X1 port map( B1 => n22442, B2 => n1349, A => n23143, ZN => 
                           n23150);
   U23585 : NOR2_X1 port map( A1 => n24325, A2 => n24906, ZN => n23149);
   U23586 : NAND3_X1 port map( A1 => n23147, A2 => n23146, A3 => n23145, ZN => 
                           n23148);
   U23587 : OAI21_X1 port map( B1 => n23150, B2 => n23149, A => n23148, ZN => 
                           n23152);
   U23588 : XNOR2_X1 port map( A => n23152, B => n23151, ZN => Ciphertext(20));
   U23589 : NAND2_X1 port map( A1 => n23154, A2 => n24473, ZN => n23156);
   U23590 : NAND2_X1 port map( A1 => n23156, A2 => n23155, ZN => n23159);
   U23591 : AOI22_X1 port map( A1 => n24325, A2 => n23159, B1 => n23158, B2 => 
                           n1349, ZN => n23162);
   U23592 : NAND2_X1 port map( A1 => n23160, A2 => n22442, ZN => n23161);
   U23593 : NAND2_X1 port map( A1 => n23162, A2 => n23161, ZN => n23163);
   U23594 : XNOR2_X1 port map( A => n23163, B => n14879, ZN => Ciphertext(23));
   U23595 : AND2_X1 port map( A1 => n23178, A2 => n23164, ZN => n23174);
   U23596 : NOR2_X1 port map( A1 => n23165, A2 => n23166, ZN => n23175);
   U23597 : AOI21_X1 port map( B1 => n23174, B2 => n23166, A => n23175, ZN => 
                           n23171);
   U23598 : NAND2_X1 port map( A1 => n23181, A2 => n23166, ZN => n23169);
   U23599 : NAND3_X1 port map( A1 => n23169, A2 => n23168, A3 => n23167, ZN => 
                           n23170);
   U23600 : NAND2_X1 port map( A1 => n23171, A2 => n23170, ZN => n23173);
   U23601 : INV_X1 port map( A => n923, ZN => n23172);
   U23602 : XNOR2_X1 port map( A => n23173, B => n23172, ZN => Ciphertext(25));
   U23603 : NOR2_X1 port map( A1 => n23175, A2 => n23174, ZN => n23182);
   U23604 : AOI21_X1 port map( B1 => n23178, B2 => n24394, A => n23176, ZN => 
                           n23180);
   U23605 : NAND2_X1 port map( A1 => n23186, A2 => n23206, ZN => n23190);
   U23606 : NAND3_X1 port map( A1 => n23201, A2 => n23202, A3 => n25059, ZN => 
                           n23189);
   U23607 : INV_X1 port map( A => n24889, ZN => n23185);
   U23608 : OAI21_X1 port map( B1 => n25059, B2 => n24334, A => n23185, ZN => 
                           n23187);
   U23609 : NAND2_X1 port map( A1 => n23187, A2 => n23194, ZN => n23188);
   U23610 : INV_X1 port map( A => n2903, ZN => n23207);
   U23611 : XNOR2_X1 port map( A => n23186, B => n23207, ZN => n23199);
   U23612 : NAND3_X1 port map( A1 => n23194, A2 => n23207, A3 => n23193, ZN => 
                           n23195);
   U23614 : NOR2_X1 port map( A1 => n23202, A2 => n23201, ZN => n23204);
   U23616 : INV_X1 port map( A => n23208, ZN => n23205);
   U23618 : NAND3_X1 port map( A1 => n23208, A2 => n23207, A3 => n23206, ZN => 
                           n23209);
   U23619 : AND3_X1 port map( A1 => n23211, A2 => n23210, A3 => n23209, ZN => 
                           Ciphertext(32));
   U23620 : NOR2_X1 port map( A1 => n23227, A2 => n25367, ZN => n23212);
   U23621 : OAI211_X1 port map( C1 => n23213, C2 => n23219, A => n24955, B => 
                           n23227, ZN => n23214);
   U23622 : OAI21_X1 port map( B1 => n23232, B2 => n23215, A => n23214, ZN => 
                           n23216);
   U23623 : XNOR2_X1 port map( A => n23216, B => n5433, ZN => Ciphertext(37));
   U23624 : MUX2_X1 port map( A => n1340, B => n23218, S => n23217, Z => n23224
                           );
   U23626 : OAI21_X1 port map( B1 => n23224, B2 => n25367, A => n23223, ZN => 
                           n23226);
   U23627 : XNOR2_X1 port map( A => n23226, B => n23225, ZN => Ciphertext(40));
   U23628 : AOI21_X1 port map( B1 => n317, B2 => n23229, A => n25367, ZN => 
                           n23230);
   U23629 : OAI22_X1 port map( A1 => n23232, A2 => n23231, B1 => n23218, B2 => 
                           n23230, ZN => n23234);
   U23630 : INV_X1 port map( A => n2036, ZN => n23233);
   U23631 : XNOR2_X1 port map( A => n23234, B => n23233, ZN => Ciphertext(41));
   U23632 : OAI21_X1 port map( B1 => n23235, B2 => n23254, A => n24377, ZN => 
                           n23238);
   U23633 : NAND3_X1 port map( A1 => n23236, A2 => n23241, A3 => n23250, ZN => 
                           n23237);
   U23634 : AND2_X1 port map( A1 => n23242, A2 => n23250, ZN => n23253);
   U23635 : NAND2_X1 port map( A1 => n23253, A2 => n23245, ZN => n23243);
   U23636 : OAI211_X1 port map( C1 => n189, C2 => n23245, A => n23244, B => 
                           n23243, ZN => n23248);
   U23637 : INV_X1 port map( A => n1835, ZN => n23247);
   U23638 : XNOR2_X1 port map( A => n23248, B => n23247, ZN => Ciphertext(43));
   U23639 : AOI21_X1 port map( B1 => n24377, B2 => n23250, A => n23249, ZN => 
                           n23255);
   U23640 : INV_X1 port map( A => n2190, ZN => n23257);
   U23641 : MUX2_X1 port map( A => n24349, B => n23274, S => n23273, Z => 
                           n23261);
   U23642 : AND2_X1 port map( A1 => n23275, A2 => n24349, ZN => n23258);
   U23643 : AOI22_X1 port map( A1 => n23259, A2 => n23281, B1 => n23258, B2 => 
                           n24360, ZN => n23260);
   U23644 : OAI21_X1 port map( B1 => n23261, B2 => n23281, A => n23260, ZN => 
                           n23262);
   U23645 : XNOR2_X1 port map( A => n23262, B => n2964, ZN => Ciphertext(51));
   U23646 : AND2_X1 port map( A1 => n23277, A2 => n24349, ZN => n23266);
   U23647 : NOR2_X1 port map( A1 => n23275, A2 => n24349, ZN => n23264);
   U23648 : AOI22_X1 port map( A1 => n23267, A2 => n23266, B1 => n23265, B2 => 
                           n23264, ZN => n23270);
   U23649 : NAND2_X1 port map( A1 => n24907, A2 => n23275, ZN => n23268);
   U23650 : OAI211_X1 port map( C1 => n24360, C2 => n24486, A => n23281, B => 
                           n23268, ZN => n23269);
   U23651 : NAND2_X1 port map( A1 => n23270, A2 => n23269, ZN => n23272);
   U23652 : XNOR2_X1 port map( A => n23272, B => n23271, ZN => Ciphertext(52));
   U23653 : NOR2_X1 port map( A1 => n23274, A2 => n23273, ZN => n23276);
   U23654 : OAI21_X1 port map( B1 => n23276, B2 => n24486, A => n23281, ZN => 
                           n23280);
   U23655 : NAND3_X1 port map( A1 => n23278, A2 => n24907, A3 => n23277, ZN => 
                           n23279);
   U23656 : OAI211_X1 port map( C1 => n23282, C2 => n23281, A => n23280, B => 
                           n23279, ZN => n23284);
   U23657 : XNOR2_X1 port map( A => n23284, B => n23283, ZN => Ciphertext(53));
   U23658 : NOR2_X1 port map( A1 => n24903, A2 => n23294, ZN => n23286);
   U23659 : OAI21_X1 port map( B1 => n23298, B2 => n23286, A => n23308, ZN => 
                           n23289);
   U23660 : OAI21_X1 port map( B1 => n23292, B2 => n23308, A => n23305, ZN => 
                           n23287);
   U23661 : NAND2_X1 port map( A1 => n23287, A2 => n23294, ZN => n23288);
   U23663 : INV_X1 port map( A => n1924, ZN => n23290);
   U23664 : XNOR2_X1 port map( A => n23291, B => n23290, ZN => Ciphertext(54));
   U23665 : NAND2_X1 port map( A1 => n23292, A2 => n23305, ZN => n23296);
   U23666 : MUX2_X1 port map( A => n23296, B => n23295, S => n23294, Z => 
                           n23301);
   U23667 : INV_X1 port map( A => n876, ZN => n23302);
   U23668 : INV_X1 port map( A => n23303, ZN => n23304);
   U23669 : OAI21_X1 port map( B1 => n23306, B2 => n23305, A => n23304, ZN => 
                           n23307);
   U23670 : OAI21_X1 port map( B1 => n23309, B2 => n23308, A => n23307, ZN => 
                           n23310);
   U23671 : XNOR2_X1 port map( A => n23310, B => n3344, ZN => Ciphertext(59));
   U23672 : OAI21_X1 port map( B1 => n4108, B2 => n23318, A => n24316, ZN => 
                           n23312);
   U23673 : NAND3_X1 port map( A1 => n23313, A2 => n23326, A3 => n23317, ZN => 
                           n23314);
   U23674 : INV_X1 port map( A => n912, ZN => n23315);
   U23675 : XNOR2_X1 port map( A => n23316, B => n23315, ZN => Ciphertext(60));
   U23676 : OAI211_X1 port map( C1 => n23320, C2 => n5659, A => n23319, B => 
                           n23326, ZN => n23321);
   U23677 : XNOR2_X1 port map( A => n23323, B => n23322, ZN => Ciphertext(64));
   U23678 : NAND2_X1 port map( A1 => n23325, A2 => n24316, ZN => n23329);
   U23680 : XNOR2_X1 port map( A => n23331, B => n23330, ZN => Ciphertext(65));
   U23681 : AOI21_X1 port map( B1 => n25081, B2 => n24341, A => n25004, ZN => 
                           n23339);
   U23682 : NAND2_X1 port map( A1 => n24342, A2 => n5421, ZN => n23337);
   U23683 : NOR2_X1 port map( A1 => n23334, A2 => n25081, ZN => n23335);
   U23684 : AOI21_X1 port map( B1 => n23337, B2 => n25081, A => n23335, ZN => 
                           n23338);
   U23685 : OAI21_X1 port map( B1 => n23339, B2 => n23338, A => n1397, ZN => 
                           n23341);
   U23686 : AOI21_X1 port map( B1 => n24492, B2 => n23341, A => n23340, ZN => 
                           n23346);
   U23687 : AOI21_X1 port map( B1 => n24400, B2 => n24492, A => n23350, ZN => 
                           n23345);
   U23688 : NOR2_X1 port map( A1 => n23354, A2 => n22961, ZN => n23360);
   U23689 : NOR2_X1 port map( A1 => n24400, A2 => n23359, ZN => n23343);
   U23690 : OAI21_X1 port map( B1 => n23360, B2 => n23343, A => n23349, ZN => 
                           n23344);
   U23691 : OAI21_X1 port map( B1 => n23346, B2 => n23345, A => n23344, ZN => 
                           n23348);
   U23692 : XNOR2_X1 port map( A => n23348, B => n23347, ZN => Ciphertext(68));
   U23695 : INV_X1 port map( A => n23359, ZN => n23353);
   U23696 : OAI21_X1 port map( B1 => n24343, B2 => n23353, A => n23350, ZN => 
                           n23356);
   U23697 : XNOR2_X1 port map( A => n23358, B => n3115, ZN => Ciphertext(70));
   U23698 : OAI21_X1 port map( B1 => n23360, B2 => n23359, A => n23350, ZN => 
                           n23365);
   U23699 : INV_X1 port map( A => n889, ZN => n23366);
   U23700 : XNOR2_X1 port map( A => n23367, B => n23366, ZN => Ciphertext(71));
   U23701 : NAND2_X1 port map( A1 => n23370, A2 => n23368, ZN => n23378);
   U23702 : NAND3_X1 port map( A1 => n23370, A2 => n23371, A3 => n24412, ZN => 
                           n23377);
   U23703 : INV_X1 port map( A => n23371, ZN => n23373);
   U23704 : AOI22_X1 port map( A1 => n23375, A2 => n23374, B1 => n23373, B2 => 
                           n23372, ZN => n23376);
   U23705 : OAI211_X1 port map( C1 => n23379, C2 => n23378, A => n23377, B => 
                           n23376, ZN => n23381);
   U23706 : INV_X1 port map( A => n836, ZN => n23380);
   U23707 : XNOR2_X1 port map( A => n23381, B => n23380, ZN => Ciphertext(72));
   U23708 : MUX2_X1 port map( A => n23396, B => n23394, S => n23391, Z => 
                           n23383);
   U23709 : MUX2_X1 port map( A => n24933, B => n23393, S => n24880, Z => 
                           n23382);
   U23710 : MUX2_X1 port map( A => n23383, B => n23382, S => n23392, Z => 
                           n23384);
   U23711 : XNOR2_X1 port map( A => n23384, B => n5251, ZN => Ciphertext(80));
   U23712 : AOI22_X1 port map( A1 => n24880, A2 => n23386, B1 => n23392, B2 => 
                           n23394, ZN => n23388);
   U23713 : NOR3_X1 port map( A1 => n24449, A2 => n22026, A3 => n23396, ZN => 
                           n23387);
   U23714 : AOI21_X1 port map( B1 => n23388, B2 => n23389, A => n23387, ZN => 
                           n23390);
   U23715 : XNOR2_X1 port map( A => n23390, B => n1891, ZN => Ciphertext(81));
   U23716 : MUX2_X1 port map( A => n24880, B => n22026, S => n24449, Z => 
                           n23397);
   U23718 : INV_X1 port map( A => n23410, ZN => n23417);
   U23719 : NAND3_X1 port map( A1 => n906, A2 => n25035, A3 => n24426, ZN => 
                           n23399);
   U23720 : INV_X1 port map( A => n2208, ZN => n23401);
   U23721 : INV_X1 port map( A => n23416, ZN => n23402);
   U23722 : AOI22_X1 port map( A1 => n23402, A2 => n23417, B1 => n23420, B2 => 
                           n23411, ZN => n23422);
   U23723 : NAND2_X1 port map( A1 => n24977, A2 => n23398, ZN => n23404);
   U23724 : NAND3_X1 port map( A1 => n23404, A2 => n25035, A3 => n24947, ZN => 
                           n23405);
   U23725 : OAI21_X1 port map( B1 => n23422, B2 => n23406, A => n23405, ZN => 
                           n23408);
   U23726 : INV_X1 port map( A => n1776, ZN => n23407);
   U23727 : XNOR2_X1 port map( A => n23408, B => n23407, ZN => Ciphertext(85));
   U23728 : NAND2_X1 port map( A1 => n23416, A2 => n23410, ZN => n23413);
   U23729 : AOI21_X1 port map( B1 => n23418, B2 => n23417, A => n23416, ZN => 
                           n23419);
   U23730 : OAI22_X1 port map( A1 => n23422, A2 => n24426, B1 => n23420, B2 => 
                           n23419, ZN => n23424);
   U23731 : INV_X1 port map( A => n2031, ZN => n23423);
   U23732 : XNOR2_X1 port map( A => n23424, B => n23423, ZN => Ciphertext(89));
   U23733 : NAND3_X1 port map( A1 => n23449, A2 => n22528, A3 => n23443, ZN => 
                           n23429);
   U23734 : OAI21_X1 port map( B1 => n23449, B2 => n23425, A => n23442, ZN => 
                           n23433);
   U23735 : NAND2_X1 port map( A1 => n23433, A2 => n22506, ZN => n23427);
   U23736 : NOR2_X1 port map( A1 => n24989, A2 => n1370, ZN => n23426);
   U23737 : NAND2_X1 port map( A1 => n23449, A2 => n23426, ZN => n23428);
   U23738 : NAND4_X1 port map( A1 => n23429, A2 => n23427, A3 => n2211, A4 => 
                           n23428, ZN => n23436);
   U23739 : INV_X1 port map( A => n23428, ZN => n23431);
   U23740 : INV_X1 port map( A => n23429, ZN => n23430);
   U23741 : OAI21_X1 port map( B1 => n23431, B2 => n23430, A => n23432, ZN => 
                           n23435);
   U23742 : NAND3_X1 port map( A1 => n23433, A2 => n23432, A3 => n22506, ZN => 
                           n23434);
   U23743 : NAND3_X1 port map( A1 => n23436, A2 => n23435, A3 => n23434, ZN => 
                           Ciphertext(90));
   U23744 : AOI21_X1 port map( B1 => n23449, B2 => n23425, A => n23437, ZN => 
                           n23439);
   U23745 : NAND3_X1 port map( A1 => n23437, A2 => n22528, A3 => n23443, ZN => 
                           n23438);
   U23746 : OAI21_X1 port map( B1 => n23439, B2 => n23453, A => n23438, ZN => 
                           n23440);
   U23747 : XNOR2_X1 port map( A => n23440, B => n494, ZN => Ciphertext(91));
   U23748 : NAND3_X1 port map( A1 => n321, A2 => n23450, A3 => n22528, ZN => 
                           n23446);
   U23749 : NAND3_X1 port map( A1 => n23442, A2 => n1370, A3 => n22528, ZN => 
                           n23445);
   U23750 : INV_X1 port map( A => n23449, ZN => n23452);
   U23751 : OAI21_X1 port map( B1 => n23450, B2 => n1370, A => n321, ZN => 
                           n23451);
   U23752 : AOI22_X1 port map( A1 => n23453, A2 => n23452, B1 => n23451, B2 => 
                           n22528, ZN => n23454);
   U23753 : XNOR2_X1 port map( A => n23454, B => n2240, ZN => Ciphertext(95));
   U23754 : MUX2_X1 port map( A => n23491, B => n23481, S => n23480, Z => 
                           n23456);
   U23755 : OAI21_X1 port map( B1 => n23499, B2 => n23494, A => n24336, ZN => 
                           n23455);
   U23758 : AOI21_X1 port map( B1 => n23458, B2 => n23461, A => n23464, ZN => 
                           n23466);
   U23759 : NAND2_X1 port map( A1 => n23460, A2 => n24364, ZN => n23465);
   U23761 : AOI22_X1 port map( A1 => n23466, A2 => n23465, B1 => n25055, B2 => 
                           n23463, ZN => n23468);
   U23763 : NAND2_X1 port map( A1 => n23483, A2 => n23472, ZN => n23475);
   U23765 : NAND2_X1 port map( A1 => n23011, A2 => n23472, ZN => n23471);
   U23766 : OAI211_X1 port map( C1 => n24442, C2 => n23472, A => n23471, B => 
                           n24336, ZN => n23473);
   U23767 : OAI211_X1 port map( C1 => n23499, C2 => n23475, A => n23474, B => 
                           n23473, ZN => n23477);
   U23768 : XNOR2_X1 port map( A => n23477, B => n23476, ZN => Ciphertext(98));
   U23769 : AND2_X1 port map( A1 => n23479, A2 => n23478, ZN => n23490);
   U23770 : NOR2_X1 port map( A1 => n23480, A2 => n23479, ZN => n23482);
   U23771 : AOI22_X1 port map( A1 => n23490, A2 => n23499, B1 => n23482, B2 => 
                           n23481, ZN => n23488);
   U23773 : OAI211_X1 port map( C1 => n24442, C2 => n24336, A => n23485, B => 
                           n23484, ZN => n23487);
   U23774 : INV_X1 port map( A => n2882, ZN => n23489);
   U23775 : INV_X1 port map( A => n23490, ZN => n23498);
   U23776 : NAND2_X1 port map( A1 => n23493, A2 => n23499, ZN => n23497);
   U23777 : NAND2_X1 port map( A1 => n23495, A2 => n23494, ZN => n23496);
   U23778 : OAI211_X1 port map( C1 => n23499, C2 => n23498, A => n23497, B => 
                           n23496, ZN => n23501);
   U23779 : XNOR2_X1 port map( A => n23501, B => n23500, ZN => Ciphertext(101))
                           ;
   U23780 : NOR2_X1 port map( A1 => n24351, A2 => n23505, ZN => n23504);
   U23781 : INV_X1 port map( A => n23527, ZN => n23503);
   U23782 : OAI21_X1 port map( B1 => n23510, B2 => n23505, A => n24380, ZN => 
                           n23506);
   U23783 : OAI21_X1 port map( B1 => n23527, B2 => n24313, A => n23506, ZN => 
                           n23507);
   U23784 : XNOR2_X1 port map( A => n23509, B => n23508, ZN => Ciphertext(102))
                           ;
   U23785 : NOR2_X1 port map( A1 => n23527, A2 => n23530, ZN => n23512);
   U23786 : NOR2_X1 port map( A1 => n24351, A2 => n23510, ZN => n23511);
   U23787 : NAND2_X1 port map( A1 => n23513, A2 => n23531, ZN => n23521);
   U23788 : NOR2_X1 port map( A1 => n23514, A2 => n24313, ZN => n23519);
   U23789 : NOR3_X1 port map( A1 => n23517, A2 => n23516, A3 => n23515, ZN => 
                           n23518);
   U23790 : NAND2_X1 port map( A1 => n23519, A2 => n23518, ZN => n23520);
   U23791 : OAI211_X1 port map( C1 => n23522, C2 => n23531, A => n23521, B => 
                           n23520, ZN => n23524);
   U23792 : XNOR2_X1 port map( A => n23524, B => n23523, ZN => Ciphertext(105))
                           ;
   U23793 : INV_X1 port map( A => n24313, ZN => n23526);
   U23794 : NOR3_X1 port map( A1 => n23527, A2 => n23526, A3 => n24351, ZN => 
                           n23528);
   U23795 : OR2_X1 port map( A1 => n23530, A2 => n23529, ZN => n23532);
   U23796 : XNOR2_X1 port map( A => n23534, B => n2739, ZN => Ciphertext(106));
   U23797 : NOR2_X1 port map( A1 => n23546, A2 => n23547, ZN => n23563);
   U23798 : INV_X1 port map( A => n23563, ZN => n23540);
   U23799 : NAND2_X1 port map( A1 => n23537, A2 => n23554, ZN => n23535);
   U23800 : OAI21_X1 port map( B1 => n25071, B2 => n23537, A => n23535, ZN => 
                           n23536);
   U23801 : INV_X1 port map( A => n23555, ZN => n23538);
   U23802 : NAND3_X1 port map( A1 => n23538, A2 => n25071, A3 => n23537, ZN => 
                           n23539);
   U23803 : INV_X1 port map( A => n1364, ZN => n23541);
   U23804 : XNOR2_X1 port map( A => n23542, B => n23541, ZN => Ciphertext(108))
                           ;
   U23805 : INV_X1 port map( A => n23554, ZN => n23556);
   U23806 : OAI21_X1 port map( B1 => n23555, B2 => n24057, A => n23556, ZN => 
                           n23550);
   U23809 : NAND3_X1 port map( A1 => n323, A2 => n23547, A3 => n25071, ZN => 
                           n23548);
   U23810 : OAI211_X1 port map( C1 => n23551, C2 => n23550, A => n23549, B => 
                           n23548, ZN => n23553);
   U23811 : INV_X1 port map( A => n1826, ZN => n23552);
   U23812 : XNOR2_X1 port map( A => n23553, B => n23552, ZN => Ciphertext(111))
                           ;
   U23813 : OAI21_X1 port map( B1 => n24893, B2 => n23555, A => n23554, ZN => 
                           n23562);
   U23814 : NAND3_X1 port map( A1 => n23557, A2 => n23556, A3 => n323, ZN => 
                           n23561);
   U23815 : NAND2_X1 port map( A1 => n23563, A2 => n24057, ZN => n23560);
   U23816 : INV_X1 port map( A => n1920, ZN => n23564);
   U23817 : NOR2_X1 port map( A1 => n23592, A2 => n23566, ZN => n23597);
   U23818 : INV_X1 port map( A => n23597, ZN => n23569);
   U23819 : OAI211_X1 port map( C1 => n1328, C2 => n23596, A => n24389, B => 
                           n23565, ZN => n23568);
   U23820 : NAND3_X1 port map( A1 => n23595, A2 => n23566, A3 => n24901, ZN => 
                           n23567);
   U23821 : NAND3_X1 port map( A1 => n23569, A2 => n23568, A3 => n23567, ZN => 
                           n23570);
   U23822 : XNOR2_X1 port map( A => n23570, B => n4589, ZN => Ciphertext(115));
   U23823 : OR2_X1 port map( A1 => n23573, A2 => n23572, ZN => n23581);
   U23824 : AND2_X1 port map( A1 => n23576, A2 => n23577, ZN => n23582);
   U23825 : NOR4_X1 port map( A1 => n23579, A2 => n23581, A3 => n23578, A4 => 
                           n23582, ZN => n23580);
   U23826 : NAND2_X1 port map( A1 => n23580, A2 => n23591, ZN => n23588);
   U23827 : OAI21_X1 port map( B1 => n23582, B2 => n23581, A => n23594, ZN => 
                           n23583);
   U23828 : OAI21_X1 port map( B1 => n24389, B2 => n24901, A => n23583, ZN => 
                           n23585);
   U23829 : NAND2_X1 port map( A1 => n23585, A2 => n21941, ZN => n23587);
   U23830 : XNOR2_X1 port map( A => n23590, B => n23589, ZN => Ciphertext(117))
                           ;
   U23831 : NAND2_X1 port map( A1 => n23591, A2 => n23592, ZN => n23601);
   U23832 : NAND3_X1 port map( A1 => n24611, A2 => n23592, A3 => n24901, ZN => 
                           n23600);
   U23833 : NAND3_X1 port map( A1 => n23595, A2 => n23596, A3 => n24901, ZN => 
                           n23599);
   U23834 : NAND2_X1 port map( A1 => n23597, A2 => n23596, ZN => n23598);
   U23835 : NAND4_X1 port map( A1 => n23601, A2 => n23600, A3 => n23599, A4 => 
                           n23598, ZN => n23603);
   U23836 : XNOR2_X1 port map( A => n23603, B => n23602, ZN => Ciphertext(119))
                           ;
   U23837 : INV_X1 port map( A => n23650, ZN => n23627);
   U23838 : NAND3_X1 port map( A1 => n23627, A2 => n23647, A3 => n23645, ZN => 
                           n23605);
   U23839 : NAND4_X1 port map( A1 => n24320, A2 => n23650, A3 => n20896, A4 => 
                           n23637, ZN => n23604);
   U23840 : OAI211_X1 port map( C1 => n23606, C2 => n23645, A => n23605, B => 
                           n23604, ZN => n23608);
   U23841 : INV_X1 port map( A => n2805, ZN => n23607);
   U23842 : XNOR2_X1 port map( A => n23608, B => n23607, ZN => Ciphertext(121))
                           ;
   U23843 : NAND2_X1 port map( A1 => n23612, A2 => n23620, ZN => n23609);
   U23844 : INV_X1 port map( A => n23609, ZN => n23610);
   U23845 : OAI211_X1 port map( C1 => n23620, C2 => n24320, A => n23609, B => 
                           n23653, ZN => n23618);
   U23846 : INV_X1 port map( A => n23647, ZN => n23651);
   U23847 : NAND2_X1 port map( A1 => n23610, A2 => n23651, ZN => n23616);
   U23848 : NOR2_X1 port map( A1 => n23648, A2 => n23620, ZN => n23611);
   U23849 : AOI21_X1 port map( B1 => n23611, B2 => n23647, A => n23645, ZN => 
                           n23615);
   U23850 : INV_X1 port map( A => n23620, ZN => n23624);
   U23851 : XNOR2_X1 port map( A => n23650, B => n23624, ZN => n23613);
   U23852 : OR2_X1 port map( A1 => n23613, A2 => n24320, ZN => n23614);
   U23853 : NAND3_X1 port map( A1 => n23616, A2 => n23615, A3 => n23614, ZN => 
                           n23617);
   U23854 : NAND2_X1 port map( A1 => n23618, A2 => n23617, ZN => n23626);
   U23855 : NAND2_X1 port map( A1 => n23619, A2 => n23620, ZN => n23622);
   U23856 : NAND2_X1 port map( A1 => n23634, A2 => n23620, ZN => n23621);
   U23857 : NAND4_X1 port map( A1 => n23622, A2 => n23645, A3 => n23649, A4 => 
                           n23621, ZN => n23623);
   U23858 : AOI21_X1 port map( B1 => n23652, B2 => n23624, A => n23623, ZN => 
                           n23625);
   U23859 : NOR2_X1 port map( A1 => n23626, A2 => n23625, ZN => Ciphertext(122)
                           );
   U23860 : NAND2_X1 port map( A1 => n23627, A2 => n23645, ZN => n23638);
   U23861 : NOR2_X1 port map( A1 => n23647, A2 => n23648, ZN => n23628);
   U23862 : NAND2_X1 port map( A1 => n23628, A2 => n23645, ZN => n23632);
   U23863 : NAND3_X1 port map( A1 => n23629, A2 => n23637, A3 => n23649, ZN => 
                           n23630);
   U23864 : NAND4_X1 port map( A1 => n23631, A2 => n3164, A3 => n23632, A4 => 
                           n23630, ZN => n23644);
   U23866 : INV_X1 port map( A => n3164, ZN => n23639);
   U23868 : INV_X1 port map( A => n23645, ZN => n23636);
   U23869 : NOR2_X1 port map( A1 => n23634, A2 => n3164, ZN => n23635);
   U23870 : NAND4_X1 port map( A1 => n23637, A2 => n23636, A3 => n23635, A4 => 
                           n23649, ZN => n23642);
   U23871 : NAND4_X1 port map( A1 => n23644, A2 => n23643, A3 => n23642, A4 => 
                           n23641, ZN => Ciphertext(123));
   U23872 : NAND2_X1 port map( A1 => n23648, A2 => n23645, ZN => n23646);
   U23873 : OAI211_X1 port map( C1 => n23648, C2 => n23649, A => n23647, B => 
                           n23646, ZN => n23656);
   U23874 : NAND3_X1 port map( A1 => n23651, A2 => n23650, A3 => n23649, ZN => 
                           n23655);
   U23875 : NAND2_X1 port map( A1 => n23653, A2 => n23652, ZN => n23654);
   U23876 : INV_X1 port map( A => n1746, ZN => n23657);
   U23877 : AND2_X1 port map( A1 => n23658, A2 => n25026, ZN => n23662);
   U23878 : NAND2_X1 port map( A1 => n23665, A2 => n23689, ZN => n23661);
   U23879 : AND2_X1 port map( A1 => n23659, A2 => n25026, ZN => n23660);
   U23880 : XNOR2_X1 port map( A => n23664, B => n23663, ZN => Ciphertext(127))
                           ;
   U23881 : INV_X1 port map( A => n23679, ZN => n23666);
   U23882 : NOR3_X1 port map( A1 => n23669, A2 => n23668, A3 => n23678, ZN => 
                           n23685);
   U23883 : AOI21_X1 port map( B1 => n23671, B2 => n23679, A => n23670, ZN => 
                           n23675);
   U23884 : OR3_X1 port map( A1 => n23672, A2 => n23679, A3 => n23671, ZN => 
                           n23674);
   U23885 : NAND2_X1 port map( A1 => n23672, A2 => n23679, ZN => n23673);
   U23886 : NAND3_X1 port map( A1 => n23675, A2 => n23674, A3 => n23673, ZN => 
                           n23684);
   U23887 : OR2_X1 port map( A1 => n23692, A2 => n23679, ZN => n23682);
   U23888 : INV_X1 port map( A => n23690, ZN => n23677);
   U23890 : OAI21_X1 port map( B1 => n23682, B2 => n23681, A => n23680, ZN => 
                           n23683);
   U23891 : INV_X1 port map( A => n23699, ZN => n23703);
   U23892 : NOR2_X1 port map( A1 => n23714, A2 => n23703, ZN => n23705);
   U23893 : INV_X1 port map( A => n23705, ZN => n23695);
   U23894 : NAND3_X1 port map( A1 => n5284, A2 => n23716, A3 => n23703, ZN => 
                           n23694);
   U23895 : OAI21_X1 port map( B1 => n23696, B2 => n23695, A => n23694, ZN => 
                           n23711);
   U23896 : NOR2_X1 port map( A1 => n23715, A2 => n23699, ZN => n23698);
   U23897 : NAND2_X1 port map( A1 => n23714, A2 => n23703, ZN => n23701);
   U23898 : NAND2_X1 port map( A1 => n23712, A2 => n23699, ZN => n23700);
   U23899 : OAI21_X1 port map( B1 => n23712, B2 => n23701, A => n23700, ZN => 
                           n23708);
   U23900 : NAND2_X1 port map( A1 => n23720, A2 => n23703, ZN => n23702);
   U23901 : OAI21_X1 port map( B1 => n23720, B2 => n23703, A => n23702, ZN => 
                           n23704);
   U23902 : NAND3_X1 port map( A1 => n23704, A2 => n23715, A3 => n23714, ZN => 
                           n23707);
   U23903 : OAI211_X1 port map( C1 => n23709, C2 => n23708, A => n23707, B => 
                           n23706, ZN => n23710);
   U23904 : AOI21_X1 port map( B1 => n24374, B2 => n23711, A => n23710, ZN => 
                           Ciphertext(134));
   U23905 : INV_X1 port map( A => n23720, ZN => n23713);
   U23906 : MUX2_X1 port map( A => n23715, B => n23713, S => n23712, Z => 
                           n23718);
   U23907 : NAND3_X1 port map( A1 => n23719, A2 => n23715, A3 => n23714, ZN => 
                           n23717);
   U23908 : OAI21_X1 port map( B1 => n23721, B2 => n23720, A => n23719, ZN => 
                           n23722);
   U23909 : NAND2_X1 port map( A1 => n23724, A2 => n23723, ZN => n23725);
   U23910 : INV_X1 port map( A => n1869, ZN => n23729);
   U23911 : MUX2_X1 port map( A => n23743, B => n23740, S => n24065, Z => 
                           n23732);
   U23912 : AOI22_X1 port map( A1 => n23732, A2 => n23731, B1 => n24064, B2 => 
                           n23745, ZN => n23734);
   U23913 : INV_X1 port map( A => n921, ZN => n23733);
   U23914 : XNOR2_X1 port map( A => n23734, B => n23733, ZN => Ciphertext(138))
                           ;
   U23915 : OAI211_X1 port map( C1 => n23745, C2 => n997, A => n24065, B => 
                           n23740, ZN => n23736);
   U23916 : NAND2_X1 port map( A1 => n23737, A2 => n23736, ZN => n23739);
   U23917 : INV_X1 port map( A => n688, ZN => n23738);
   U23918 : XNOR2_X1 port map( A => n23739, B => n23738, ZN => Ciphertext(139))
                           ;
   U23919 : MUX2_X1 port map( A => n25460, B => n24063, S => n23740, Z => 
                           n23749);
   U23920 : NAND3_X1 port map( A1 => n23743, A2 => n24064, A3 => n25460, ZN => 
                           n23747);
   U23921 : NAND2_X1 port map( A1 => n23745, A2 => n23744, ZN => n23746);
   U23922 : OAI211_X1 port map( C1 => n23749, C2 => n23748, A => n23747, B => 
                           n23746, ZN => n23751);
   U23923 : XNOR2_X1 port map( A => n23751, B => n23750, ZN => Ciphertext(141))
                           ;
   U23924 : OAI21_X1 port map( B1 => n23779, B2 => n23769, A => n23758, ZN => 
                           n23755);
   U23925 : NAND2_X1 port map( A1 => n23779, A2 => n23768, ZN => n23753);
   U23926 : OAI21_X1 port map( B1 => n23765, B2 => n23782, A => n23753, ZN => 
                           n23754);
   U23927 : AOI21_X1 port map( B1 => n23782, B2 => n23755, A => n23754, ZN => 
                           n23756);
   U23928 : XNOR2_X1 port map( A => n23756, B => n1758, ZN => Ciphertext(144));
   U23929 : OAI21_X1 port map( B1 => n24921, B2 => n23769, A => n23781, ZN => 
                           n23761);
   U23930 : OR3_X1 port map( A1 => n23779, A2 => n23768, A3 => n24921, ZN => 
                           n23760);
   U23931 : OR2_X1 port map( A1 => n23758, A2 => n23782, ZN => n23759);
   U23932 : OAI211_X1 port map( C1 => n23762, C2 => n23761, A => n23760, B => 
                           n23759, ZN => n23764);
   U23933 : XNOR2_X1 port map( A => n23764, B => n23763, ZN => Ciphertext(147))
                           ;
   U23934 : INV_X1 port map( A => n23779, ZN => n23767);
   U23935 : INV_X1 port map( A => n23768, ZN => n23777);
   U23936 : OAI21_X1 port map( B1 => n23774, B2 => n23777, A => n23773, ZN => 
                           n23776);
   U23937 : XNOR2_X1 port map( A => n23776, B => n23775, ZN => Ciphertext(148))
                           ;
   U23938 : AOI21_X1 port map( B1 => n23779, B2 => n23778, A => n23777, ZN => 
                           n23780);
   U23939 : OAI22_X1 port map( A1 => n23783, A2 => n23782, B1 => n23781, B2 => 
                           n23780, ZN => n23785);
   U23940 : INV_X1 port map( A => n2747, ZN => n23784);
   U23941 : XNOR2_X1 port map( A => n23785, B => n23784, ZN => Ciphertext(149))
                           ;
   U23942 : OAI21_X1 port map( B1 => n21837, B2 => n23789, A => n23788, ZN => 
                           n23809);
   U23943 : AND2_X1 port map( A1 => n24895, A2 => n23798, ZN => n23793);
   U23944 : AOI21_X1 port map( B1 => n23790, B2 => n23798, A => n23793, ZN => 
                           n23791);
   U23945 : OAI21_X1 port map( B1 => n23792, B2 => n23798, A => n23791, ZN => 
                           n23808);
   U23946 : NAND3_X1 port map( A1 => n23796, A2 => n23793, A3 => n24307, ZN => 
                           n23807);
   U23947 : NAND3_X1 port map( A1 => n23796, A2 => n21837, A3 => n896, ZN => 
                           n23804);
   U23948 : OAI211_X1 port map( C1 => n24895, C2 => n23798, A => n23796, B => 
                           n24307, ZN => n23803);
   U23949 : XNOR2_X1 port map( A => n24920, B => n23798, ZN => n23801);
   U23950 : NAND2_X1 port map( A1 => n23801, A2 => n24983, ZN => n23802);
   U23951 : NAND4_X1 port map( A1 => n23805, A2 => n23804, A3 => n23803, A4 => 
                           n23802, ZN => n23806);
   U23952 : OAI211_X1 port map( C1 => n23809, C2 => n23808, A => n23807, B => 
                           n23806, ZN => Ciphertext(154));
   U23953 : AND2_X1 port map( A1 => n23810, A2 => n23817, ZN => n23824);
   U23954 : OAI21_X1 port map( B1 => n24972, B2 => n23831, A => n23824, ZN => 
                           n23815);
   U23955 : AND2_X1 port map( A1 => n23811, A2 => n23827, ZN => n23832);
   U23956 : NOR2_X1 port map( A1 => n23828, A2 => n23813, ZN => n23812);
   U23957 : AOI21_X1 port map( B1 => n23832, B2 => n23813, A => n23812, ZN => 
                           n23814);
   U23958 : INV_X1 port map( A => n641, ZN => n23816);
   U23959 : OAI21_X1 port map( B1 => n23817, B2 => n24972, A => n23032, ZN => 
                           n23823);
   U23960 : NAND2_X1 port map( A1 => n23818, A2 => n23831, ZN => n23822);
   U23961 : NOR2_X1 port map( A1 => n23827, A2 => n24972, ZN => n23820);
   U23964 : INV_X1 port map( A => n23827, ZN => n23829);
   U23965 : OAI21_X1 port map( B1 => n23830, B2 => n23829, A => n23828, ZN => 
                           n23837);
   U23966 : NAND2_X1 port map( A1 => n23832, A2 => n23831, ZN => n23836);
   U23967 : NAND2_X1 port map( A1 => n23032, A2 => n23833, ZN => n23835);
   U23968 : NAND3_X1 port map( A1 => n23837, A2 => n23836, A3 => n23835, ZN => 
                           n23838);
   U23969 : XNOR2_X1 port map( A => n23838, B => n3696, ZN => Ciphertext(161));
   U23970 : INV_X1 port map( A => n23860, ZN => n23866);
   U23971 : INV_X1 port map( A => n23857, ZN => n23864);
   U23972 : NAND3_X1 port map( A1 => n25240, A2 => n24428, A3 => n23864, ZN => 
                           n23840);
   U23973 : INV_X1 port map( A => n1810, ZN => n23841);
   U23974 : INV_X1 port map( A => n3183, ZN => n23842);
   U23975 : NOR2_X1 port map( A1 => n23857, A2 => n23842, ZN => n23844);
   U23976 : AOI21_X1 port map( B1 => n23844, B2 => n23843, A => n23865, ZN => 
                           n23850);
   U23977 : NOR2_X1 port map( A1 => n23862, A2 => n3183, ZN => n23846);
   U23978 : NAND2_X1 port map( A1 => n23857, A2 => n23846, ZN => n23849);
   U23980 : AOI21_X1 port map( B1 => n24469, B2 => n23846, A => n23853, ZN => 
                           n23847);
   U23982 : OAI21_X1 port map( B1 => n23853, B2 => n3183, A => n24428, ZN => 
                           n23852);
   U23983 : AOI211_X1 port map( C1 => n3183, C2 => n23853, A => n23866, B => 
                           n23852, ZN => n23854);
   U23984 : NOR3_X1 port map( A1 => n23856, A2 => n23855, A3 => n23854, ZN => 
                           Ciphertext(164));
   U23985 : NAND2_X1 port map( A1 => n24469, A2 => n23857, ZN => n23861);
   U23986 : NAND2_X1 port map( A1 => n24428, A2 => n23865, ZN => n23863);
   U23987 : OAI211_X1 port map( C1 => n23866, C2 => n23865, A => n23864, B => 
                           n23863, ZN => n23867);
   U23988 : INV_X1 port map( A => Key(190), ZN => n23868);
   U23990 : NOR2_X1 port map( A1 => n23904, A2 => n23890, ZN => n23907);
   U23991 : NAND2_X1 port map( A1 => n23907, A2 => n23889, ZN => n23871);
   U23992 : INV_X1 port map( A => n1827, ZN => n23873);
   U23993 : XNOR2_X1 port map( A => n23874, B => n23873, ZN => Ciphertext(169))
                           ;
   U23994 : NAND2_X1 port map( A1 => n23896, A2 => n23883, ZN => n23875);
   U23996 : XNOR2_X1 port map( A => n23890, B => n24624, ZN => n23876);
   U23997 : OAI21_X1 port map( B1 => n23876, B2 => n23879, A => n23902, ZN => 
                           n23877);
   U23998 : XNOR2_X1 port map( A => n23906, B => n24624, ZN => n23886);
   U23999 : NAND2_X1 port map( A1 => n23905, A2 => n23889, ZN => n23885);
   U24000 : NOR2_X1 port map( A1 => n23905, A2 => n23902, ZN => n23882);
   U24001 : NAND2_X1 port map( A1 => n23903, A2 => n23883, ZN => n23881);
   U24002 : NAND2_X1 port map( A1 => n23888, A2 => n23906, ZN => n23899);
   U24003 : NAND3_X1 port map( A1 => n23890, A2 => n23889, A3 => n23903, ZN => 
                           n23898);
   U24004 : NOR2_X1 port map( A1 => n23894, A2 => n23905, ZN => n23895);
   U24005 : OAI21_X1 port map( B1 => n23896, B2 => n23902, A => n23895, ZN => 
                           n23897);
   U24007 : INV_X1 port map( A => n1724, ZN => n23900);
   U24008 : XNOR2_X1 port map( A => n23901, B => n23900, ZN => Ciphertext(171))
                           ;
   U24009 : AOI21_X1 port map( B1 => n23906, B2 => n23902, A => n23905, ZN => 
                           n23908);
   U24010 : XNOR2_X1 port map( A => n23910, B => n5484, ZN => Ciphertext(173));
   U24011 : NAND2_X1 port map( A1 => n23911, A2 => n25083, ZN => n23936);
   U24012 : INV_X1 port map( A => n23937, ZN => n23912);
   U24013 : NAND3_X1 port map( A1 => n23912, A2 => n23926, A3 => n23933, ZN => 
                           n23914);
   U24014 : NAND4_X1 port map( A1 => n23915, A2 => n23936, A3 => n23914, A4 => 
                           n23913, ZN => n23917);
   U24015 : XNOR2_X1 port map( A => n23917, B => n23916, ZN => Ciphertext(174))
                           ;
   U24016 : OAI211_X1 port map( C1 => n23937, C2 => n23924, A => n23926, B => 
                           n23918, ZN => n23919);
   U24017 : OAI211_X1 port map( C1 => n23924, C2 => n23921, A => n23920, B => 
                           n23919, ZN => n23923);
   U24018 : XNOR2_X1 port map( A => n23923, B => n23922, ZN => Ciphertext(175))
                           ;
   U24019 : NAND2_X1 port map( A1 => n23937, A2 => n23924, ZN => n23930);
   U24020 : NAND3_X1 port map( A1 => n23934, A2 => n23926, A3 => n23938, ZN => 
                           n23929);
   U24021 : NAND2_X1 port map( A1 => n23924, A2 => n23933, ZN => n23925);
   U24022 : OAI21_X1 port map( B1 => n23926, B2 => n23933, A => n23925, ZN => 
                           n23927);
   U24025 : INV_X1 port map( A => n887, ZN => n23931);
   U24027 : AOI21_X1 port map( B1 => n23934, B2 => n23933, A => n23939, ZN => 
                           n23935);
   U24028 : NAND2_X1 port map( A1 => n23936, A2 => n23935, ZN => n23944);
   U24029 : NAND3_X1 port map( A1 => n24948, A2 => n23938, A3 => n23937, ZN => 
                           n23943);
   U24030 : NAND2_X1 port map( A1 => n23941, A2 => n25083, ZN => n23942);
   U24031 : NAND3_X1 port map( A1 => n23944, A2 => n23943, A3 => n23942, ZN => 
                           n23946);
   U24032 : XNOR2_X1 port map( A => n23946, B => n23945, ZN => Ciphertext(178))
                           ;
   U24033 : OAI21_X1 port map( B1 => n23970, B2 => n23966, A => n23967, ZN => 
                           n23951);
   U24034 : OR2_X1 port map( A1 => n23969, A2 => n25017, ZN => n23948);
   U24035 : INV_X1 port map( A => n23949, ZN => n23950);
   U24036 : NAND2_X1 port map( A1 => n23969, A2 => n23952, ZN => n23955);
   U24037 : OR2_X1 port map( A1 => n23967, A2 => n24910, ZN => n23963);
   U24038 : INV_X1 port map( A => n23963, ZN => n23954);
   U24039 : XNOR2_X1 port map( A => n23956, B => n4023, ZN => Ciphertext(181));
   U24040 : MUX2_X1 port map( A => n23966, B => n24910, S => n23967, Z => 
                           n23960);
   U24041 : MUX2_X1 port map( A => n23960, B => n23959, S => n23969, Z => 
                           n23962);
   U24042 : XNOR2_X1 port map( A => n23962, B => n23961, ZN => Ciphertext(182))
                           ;
   U24043 : INV_X1 port map( A => n23969, ZN => n23965);
   U24044 : NOR2_X1 port map( A1 => n23967, A2 => n23966, ZN => n23968);
   U24045 : AOI22_X1 port map( A1 => n25076, A2 => n23970, B1 => n23969, B2 => 
                           n23968, ZN => n23971);
   U24046 : INV_X1 port map( A => n2044, ZN => n23973);
   U24047 : NAND2_X1 port map( A1 => n23982, A2 => n24012, ZN => n23974);
   U24048 : INV_X1 port map( A => n24011, ZN => n23978);
   U24049 : NOR2_X1 port map( A1 => n23982, A2 => n24011, ZN => n23975);
   U24050 : AND2_X1 port map( A1 => n24011, A2 => n24012, ZN => n24015);
   U24051 : INV_X1 port map( A => n1757, ZN => n23976);
   U24052 : XNOR2_X1 port map( A => n23977, B => n23976, ZN => Ciphertext(187))
                           ;
   U24053 : OR2_X1 port map( A1 => n23978, A2 => n23984, ZN => n23988);
   U24054 : OAI21_X1 port map( B1 => n23979, B2 => n24008, A => n23988, ZN => 
                           n23992);
   U24055 : INV_X1 port map( A => n24448, ZN => n24005);
   U24056 : NAND3_X1 port map( A1 => n24005, A2 => n24012, A3 => n24954, ZN => 
                           n23980);
   U24057 : OAI211_X1 port map( C1 => n24440, C2 => n23981, A => n23983, B => 
                           n23980, ZN => n23991);
   U24058 : NOR3_X1 port map( A1 => n24440, A2 => n24448, A3 => n24954, ZN => 
                           n23985);
   U24059 : OAI21_X1 port map( B1 => n24008, B2 => n23987, A => n23986, ZN => 
                           n23990);
   U24060 : OAI211_X1 port map( C1 => n23992, C2 => n23991, A => n23990, B => 
                           n23989, ZN => Ciphertext(188));
   U24061 : INV_X1 port map( A => n23993, ZN => n24014);
   U24062 : NAND2_X1 port map( A1 => n24014, A2 => n24954, ZN => n24018);
   U24063 : NOR2_X1 port map( A1 => n22677, A2 => n25439, ZN => n24003);
   U24064 : NAND2_X1 port map( A1 => n23997, A2 => n24003, ZN => n24001);
   U24065 : NAND3_X1 port map( A1 => n22677, A2 => n24439, A3 => n23998, ZN => 
                           n24000);
   U24066 : OAI211_X1 port map( C1 => n24003, C2 => n24002, A => n24001, B => 
                           n24000, ZN => n24004);
   U24067 : OAI21_X1 port map( B1 => n24011, B2 => n24004, A => n24448, ZN => 
                           n24007);
   U24068 : INV_X1 port map( A => n860, ZN => n24009);
   U24069 : NAND2_X1 port map( A1 => n24011, A2 => n24010, ZN => n24013);
   U24070 : NAND2_X1 port map( A1 => n24013, A2 => n24012, ZN => n24016);
   U24071 : AOI22_X1 port map( A1 => n24440, A2 => n24016, B1 => n24015, B2 => 
                           n24014, ZN => n24017);
   U24072 : OAI21_X1 port map( B1 => n24440, B2 => n24018, A => n24017, ZN => 
                           n24020);
   U24073 : XNOR2_X1 port map( A => n24020, B => n3208, ZN => Ciphertext(191));
   U1497 : XNOR2_X2 port map( A => n12301, B => n12300, ZN => n13123);
   U515 : XNOR2_X2 port map( A => n11273, B => n11272, ZN => n13013);
   U2461 : MUX2_X2 port map( A => n9278, B => n9277, S => n24511, Z => n10836);
   U120 : OR2_X1 port map( A1 => n11031, A2 => n10772, ZN => n10779);
   U1453 : BUF_X1 port map( A => n14970, Z => n16448);
   U2570 : MUX2_X2 port map( A => n6285, B => n6284, S => n7801, Z => n9155);
   U7653 : NAND3_X2 port map( A1 => n2433, A2 => n9478, A3 => n9479, ZN => 
                           n12396);
   U2351 : XNOR2_X2 port map( A => n11814, B => n11815, ZN => n13234);
   U13628 : OAI211_X2 port map( C1 => n7965, C2 => n7966, A => n7964, B => 
                           n7963, ZN => n8961);
   U1505 : BUF_X1 port map( A => n10632, Z => n10819);
   U477 : NAND2_X1 port map( A1 => n4465, A2 => n4461, ZN => n11414);
   U1529 : NAND4_X2 port map( A1 => n7398, A2 => n7396, A3 => n7397, A4 => 
                           n7395, ZN => n8860);
   U1994 : NAND3_X2 port map( A1 => n16620, A2 => n2942, A3 => n16623, ZN => 
                           n17476);
   U2623 : NAND3_X2 port map( A1 => n4370, A2 => n6951, A3 => n5528, ZN => 
                           n7474);
   U157 : NOR2_X2 port map( A1 => n24341, A2 => n23334, ZN => n22855);
   U4942 : OAI211_X1 port map( C1 => n3889, C2 => n13804, A => n13803, B => 
                           n13802, ZN => n14922);
   U81 : AND4_X2 port map( A1 => n10598, A2 => n10597, A3 => n10600, A4 => 
                           n10599, ZN => n11628);
   U1816 : OAI211_X2 port map( C1 => n1662, C2 => n19293, A => n19292, B => 
                           n19291, ZN => n21670);
   U580 : XNOR2_X1 port map( A => n8110, B => n8111, ZN => n9943);
   U5199 : OAI21_X2 port map( B1 => n4512, B2 => n6937, A => n4511, ZN => n3362
                           );
   U2013 : AND2_X2 port map( A1 => n2937, A2 => n3068, ZN => n17663);
   U1943 : XNOR2_X2 port map( A => n17857, B => n17858, ZN => n19470);
   U55 : AND3_X2 port map( A1 => n13085, A2 => n13084, A3 => n13083, ZN => 
                           n15210);
   U1443 : BUF_X1 port map( A => n15873, Z => n17087);
   U22814 : NOR2_X2 port map( A1 => n23196, A2 => n22752, ZN => n23200);
   U1525 : NAND4_X2 port map( A1 => n6586, A2 => n6584, A3 => n1088, A4 => 
                           n6585, ZN => n8634);
   U1441 : BUF_X1 port map( A => n16516, Z => n17145);
   U1528 : NAND4_X2 port map( A1 => n7366, A2 => n7368, A3 => n7367, A4 => 
                           n7369, ZN => n5614);
   U1805 : NAND4_X2 port map( A1 => n1661, A2 => n1664, A3 => n19739, A4 => 
                           n1660, ZN => n21721);
   U2457 : OAI211_X2 port map( C1 => n9570, C2 => n5739, A => n9569, B => n9568
                           , ZN => n10901);
   U1053 : INV_X1 port map( A => n396, ZN => n14077);
   U1823 : NOR2_X2 port map( A1 => n20513, A2 => n20512, ZN => n21307);
   U2685 : BUF_X1 port map( A => n5915, Z => n6162);
   U5273 : INV_X1 port map( A => n8244, ZN => n8698);
   U1500 : NAND2_X2 port map( A1 => n541, A2 => n10938, ZN => n12389);
   U2698 : BUF_X2 port map( A => n6071, Z => n6658);
   U1176 : XNOR2_X1 port map( A => n8344, B => n8343, ZN => n10100);
   U2613 : NAND2_X2 port map( A1 => n1643, A2 => n3444, ZN => n7735);
   U1110 : OAI21_X2 port map( B1 => n10290, B2 => n10291, A => n4732, ZN => 
                           n11966);
   U1462 : XNOR2_X2 port map( A => n14504, B => n14503, ZN => n15857);
   U245 : XNOR2_X1 port map( A => Key(96), B => Plaintext(96), ZN => n7032);
   U1350 : CLKBUF_X1 port map( A => Key(146), Z => n23620);
   U1605 : CLKBUF_X1 port map( A => Key(4), Z => n869);
   U2752 : CLKBUF_X1 port map( A => Key(156), Z => n20825);
   U102 : CLKBUF_X1 port map( A => Key(184), Z => n92);
   U253 : CLKBUF_X1 port map( A => Key(150), Z => n1855);
   U1662 : CLKBUF_X1 port map( A => Key(93), Z => n2033);
   U2738 : CLKBUF_X1 port map( A => Key(97), Z => n923);
   U2742 : CLKBUF_X1 port map( A => Key(101), Z => n20744);
   U99 : CLKBUF_X1 port map( A => Key(168), Z => n673);
   U100 : CLKBUF_X1 port map( A => Key(74), Z => n2757);
   U2745 : XNOR2_X1 port map( A => Key(144), B => Plaintext(144), ZN => n6373);
   U101 : CLKBUF_X1 port map( A => Key(29), Z => n2747);
   U12400 : XNOR2_X1 port map( A => n5954, B => Key(172), ZN => n6490);
   U2692 : CLKBUF_X1 port map( A => n5916, Z => n7097);
   U4560 : INV_X1 port map( A => n6651, ZN => n6894);
   U447 : AND2_X1 port map( A1 => n70, A2 => n6943, ZN => n3050);
   U179 : NAND3_X1 port map( A1 => n6031, A2 => n6032, A3 => n6030, ZN => n7257
                           );
   U191 : AND2_X1 port map( A1 => n2800, A2 => n6813, ZN => n4);
   U2642 : OR2_X1 port map( A1 => n2824, A2 => n6258, ZN => n7798);
   U4853 : OAI21_X1 port map( B1 => n7513, B2 => n1690, A => n7512, ZN => n9058
                           );
   U698 : NAND3_X1 port map( A1 => n6045, A2 => n6044, A3 => n120, ZN => n9181)
                           ;
   U892 : INV_X1 port map( A => n8475, ZN => n9194);
   U8463 : XNOR2_X1 port map( A => n2785, B => n8670, ZN => n9664);
   U3190 : XNOR2_X1 port map( A => n9112, B => n9113, ZN => n10064);
   U407 : INV_X1 port map( A => n10006, ZN => n9652);
   U321 : BUF_X1 port map( A => n9550, Z => n10048);
   U826 : BUF_X1 port map( A => n8744, Z => n10070);
   U2497 : BUF_X1 port map( A => n9820, Z => n10141);
   U2481 : XNOR2_X1 port map( A => n8984, B => n8983, ZN => n9639);
   U788 : OR2_X1 port map( A1 => n2565, A2 => n2585, ZN => n9378);
   U555 : NOR2_X1 port map( A1 => n9323, A2 => n9322, ZN => n10470);
   U4346 : AND2_X1 port map( A1 => n5272, A2 => n5276, ZN => n5271);
   U543 : AND2_X1 port map( A1 => n3863, A2 => n3864, ZN => n11215);
   U14889 : OAI211_X1 port map( C1 => n9643, C2 => n24332, A => n9642, B => 
                           n9641, ZN => n11207);
   U1126 : NAND2_X1 port map( A1 => n1168, A2 => n9224, ZN => n11122);
   U6672 : INV_X1 port map( A => n11149, ZN => n4998);
   U2425 : INV_X1 port map( A => n10800, ZN => n411);
   U746 : INV_X1 port map( A => n10375, ZN => n10587);
   U7432 : NAND3_X1 port map( A1 => n4211, A2 => n8426, A3 => n4213, ZN => 
                           n11464);
   U1173 : AOI22_X1 port map( A1 => n11095, A2 => n11094, B1 => n95, B2 => 
                           n11093, ZN => n11556);
   U2360 : CLKBUF_X1 port map( A => n11776, Z => n12296);
   U16560 : XNOR2_X1 port map( A => n12265, B => n12264, ZN => n12660);
   U16306 : XNOR2_X1 port map( A => n11855, B => n11854, ZN => n11873);
   U16776 : BUF_X1 port map( A => n12594, Z => n13292);
   U2346 : XNOR2_X1 port map( A => n11250, B => n11249, ZN => n13216);
   U662 : XNOR2_X1 port map( A => n4931, B => n11979, ZN => n111);
   U405 : INV_X1 port map( A => n13291, ZN => n12910);
   U11267 : MUX2_X1 port map( A => n13064, B => n13063, S => n12440, Z => n5113
                           );
   U692 : AND2_X1 port map( A1 => n1316, A2 => n1315, ZN => n13421);
   U2250 : NAND3_X1 port map( A1 => n5544, A2 => n5543, A3 => n12502, ZN => 
                           n13533);
   U1136 : AND2_X1 port map( A1 => n1553, A2 => n1554, ZN => n13892);
   U232 : XNOR2_X1 port map( A => n14960, B => n15358, ZN => n15185);
   U2170 : XNOR2_X1 port map( A => n14583, B => n14582, ZN => n16096);
   U2140 : XNOR2_X1 port map( A => n13973, B => n13972, ZN => n16206);
   U2162 : XNOR2_X1 port map( A => n15007, B => n15008, ZN => n16226);
   U1454 : INV_X1 port map( A => n14970, ZN => n16450);
   U3394 : OAI211_X1 port map( C1 => n16424, C2 => n14433, A => n14432, B => 
                           n14431, ZN => n17229);
   U742 : AND2_X1 port map( A1 => n17158, A2 => n17156, ZN => n16260);
   U605 : AND2_X1 port map( A1 => n3424, A2 => n15785, ZN => n17130);
   U19045 : BUF_X1 port map( A => n16260, Z => n17163);
   U5008 : AND2_X1 port map( A1 => n16375, A2 => n16533, ZN => n2430);
   U20506 : XNOR2_X1 port map( A => n18545, B => n18544, ZN => n19613);
   U972 : MUX2_X1 port map( A => n18811, B => n18810, S => n3412, Z => n20913);
   U21038 : INV_X1 port map( A => n25204, ZN => n20168);
   U968 : AND3_X1 port map( A1 => n1290, A2 => n1288, A3 => n1287, ZN => n20003
                           );
   U785 : AND2_X1 port map( A1 => n1503, A2 => n1504, ZN => n1327);
   U1884 : AOI21_X1 port map( B1 => n19236, B2 => n18869, A => n18805, ZN => 
                           n20359);
   U5086 : INV_X1 port map( A => n19777, ZN => n20236);
   U7598 : NAND2_X1 port map( A1 => n2198, A2 => n18885, ZN => n20290);
   U4769 : NAND2_X1 port map( A1 => n3962, A2 => n3963, ZN => n21751);
   U151 : OAI22_X1 port map( A1 => n1627, A2 => n5227, B1 => n5226, B2 => 
                           n22159, ZN => n23543);
   U23461 : OR2_X1 port map( A1 => n22943, A2 => n22942, ZN => n23349);
   U23762 : NOR2_X1 port map( A1 => n23468, A2 => n23467, ZN => n23472);
   U23160 : NOR2_X1 port map( A1 => n23110, A2 => n24498, ZN => n23093);
   U241 : CLKBUF_X1 port map( A => Key(115), Z => n688);
   U12158 : INV_X1 port map( A => n6751, ZN => n6675);
   U1607 : INV_X1 port map( A => n6871, ZN => n314);
   U12148 : INV_X1 port map( A => n5800, ZN => n6965);
   U2606 : INV_X1 port map( A => n8511, ZN => n7250);
   U749 : AND2_X1 port map( A1 => n6160, A2 => n6159, ZN => n8475);
   U14491 : NOR2_X1 port map( A1 => n9064, A2 => n9244, ZN => n10052);
   U1494 : BUF_X1 port map( A => n11287, Z => n13246);
   U1490 : BUF_X1 port map( A => n1324, Z => n13178);
   U1085 : NAND2_X2 port map( A1 => n13538, A2 => n13535, ZN => n14022);
   U4662 : INV_X1 port map( A => n13614, ZN => n14058);
   U6155 : INV_X2 port map( A => n1516, ZN => n17629);
   U1946 : INV_X1 port map( A => n4748, ZN => n19501);
   U11312 : NOR2_X1 port map( A1 => n18734, A2 => n19477, ZN => n18971);
   U146 : INV_X1 port map( A => n22093, ZN => n22890);
   U1368 : INV_X1 port map( A => n22389, ZN => n22974);
   U1486 : BUF_X1 port map( A => n11965, Z => n12695);
   U1185 : NAND2_X2 port map( A1 => n7753, A2 => n2623, ZN => n9057);
   U5577 : AOI21_X1 port map( B1 => n16922, B2 => n3783, A => n3782, ZN => 
                           n17720);
   U10755 : NOR2_X2 port map( A1 => n9215, A2 => n9216, ZN => n4590);
   U3 : AND2_X1 port map( A1 => n3035, A2 => n21916, ZN => n24334);
   U12 : XNOR2_X1 port map( A => n15078, B => n24303, ZN => n1122);
   U95 : NAND3_X2 port map( A1 => n2512, A2 => n24099, A3 => n5586, ZN => 
                           n20125);
   U97 : BUF_X1 port map( A => n22915, Z => n23510);
   U114 : INV_X1 port map( A => n15696, ZN => n16483);
   U138 : XNOR2_X1 port map( A => n13906, B => n15103, ZN => n14973);
   U182 : INV_X1 port map( A => n15857, ZN => n16120);
   U229 : BUF_X2 port map( A => n10135, Z => n24026);
   U230 : XNOR2_X1 port map( A => n9153, B => n9152, ZN => n10135);
   U233 : OAI21_X2 port map( B1 => n20602, B2 => n20601, A => n5363, ZN => 
                           n21734);
   U288 : OAI211_X1 port map( C1 => n16074, C2 => n15802, A => n3639, B => 
                           n3637, ZN => n17107);
   U303 : NAND4_X2 port map( A1 => n5488, A2 => n6605, A3 => n6604, A4 => n6603
                           , ZN => n7418);
   U317 : AND2_X2 port map( A1 => n3977, A2 => n3976, ZN => n18693);
   U328 : XNOR2_X1 port map( A => Key(158), B => Plaintext(158), ZN => n6919);
   U334 : BUF_X1 port map( A => n18817, Z => n19103);
   U339 : AND2_X2 port map( A1 => n10004, A2 => n10003, ZN => n11012);
   U344 : OAI21_X2 port map( B1 => n3839, B2 => n6058, A => n3838, ZN => n8022)
                           ;
   U353 : XNOR2_X2 port map( A => n5895, B => Key(52), ZN => n6697);
   U381 : NOR2_X1 port map( A1 => n20721, A2 => n20720, ZN => n23217);
   U396 : OAI211_X2 port map( C1 => n9247, C2 => n10054, A => n9246, B => n5004
                           , ZN => n10858);
   U399 : XNOR2_X2 port map( A => n19342, B => n19341, ZN => n22252);
   U427 : XNOR2_X2 port map( A => n11572, B => n11573, ZN => n13041);
   U430 : XNOR2_X2 port map( A => n11480, B => n11479, ZN => n12710);
   U444 : XNOR2_X1 port map( A => n11490, B => n11491, ZN => n13077);
   U470 : XNOR2_X1 port map( A => n21175, B => n21174, ZN => n22593);
   U497 : XNOR2_X2 port map( A => n11539, B => n11540, ZN => n12470);
   U507 : AOI22_X2 port map( A1 => n12700, A2 => n12699, B1 => n12698, B2 => 
                           n25191, ZN => n14190);
   U512 : AND2_X2 port map( A1 => n5719, A2 => n5720, ZN => n7771);
   U522 : OAI211_X2 port map( C1 => n22929, C2 => n5768, A => n1396, B => n5687
                           , ZN => n23505);
   U567 : OAI21_X2 port map( B1 => n19866, B2 => n19865, A => n19864, ZN => 
                           n20964);
   U581 : OAI211_X1 port map( C1 => n6728, C2 => n6727, A => n6726, B => n6725,
                           ZN => n263);
   U614 : XNOR2_X1 port map( A => n5783, B => Key(93), ZN => n6236);
   U632 : NOR2_X1 port map( A1 => n12599, A2 => n12598, ZN => n14851);
   U644 : NAND4_X2 port map( A1 => n7275, A2 => n7274, A3 => n7273, A4 => n7272
                           , ZN => n8875);
   U676 : XNOR2_X1 port map( A => n3504, B => n3505, ZN => n9898);
   U696 : AND2_X2 port map( A1 => n18741, A2 => n18740, ZN => n20191);
   U708 : XNOR2_X2 port map( A => n3473, B => n11945, ZN => n13274);
   U744 : OAI211_X2 port map( C1 => n7898, C2 => n7233, A => n5235, B => n5236,
                           ZN => n8612);
   U748 : NOR2_X2 port map( A1 => n7921, A2 => n8078, ZN => n9189);
   U750 : BUF_X2 port map( A => n8901, Z => n24056);
   U758 : OAI22_X1 port map( A1 => n7047, A2 => n7827, B1 => n7513, B2 => n7048
                           , ZN => n8901);
   U775 : OAI21_X2 port map( B1 => n20323, B2 => n20322, A => n20321, ZN => 
                           n24485);
   U825 : NOR2_X1 port map( A1 => n22477, A2 => n22476, ZN => n23119);
   U841 : OAI21_X2 port map( B1 => n11120, B2 => n11119, A => n11118, ZN => 
                           n11715);
   U846 : XNOR2_X1 port map( A => n13606, B => n14633, ZN => n16405);
   U852 : BUF_X1 port map( A => n23742, Z => n24064);
   U854 : BUF_X1 port map( A => n23742, Z => n24065);
   U888 : BUF_X1 port map( A => n6534, Z => n24067);
   U909 : XNOR2_X1 port map( A => n5865, B => Key(26), ZN => n6534);
   U910 : XNOR2_X2 port map( A => Key(9), B => Plaintext(9), ZN => n6498);
   U958 : NAND3_X2 port map( A1 => n10857, A2 => n3502, A3 => n24251, ZN => 
                           n12391);
   U987 : OAI211_X2 port map( C1 => n11156, C2 => n11155, A => n11154, B => 
                           n11153, ZN => n11977);
   U1009 : OAI21_X2 port map( B1 => n6443, B2 => n6442, A => n6441, ZN => n2404
                           );
   U1035 : AOI22_X1 port map( A1 => n6390, A2 => n6391, B1 => n6388, B2 => 
                           n6389, ZN => n7850);
   U1050 : XNOR2_X2 port map( A => n16600, B => n16601, ZN => n19560);
   U1074 : NAND4_X2 port map( A1 => n4404, A2 => n4403, A3 => n4402, A4 => 
                           n18850, ZN => n20068);
   U1117 : OAI211_X2 port map( C1 => n7776, C2 => n7775, A => n7773, B => n7774
                           , ZN => n9106);
   U1156 : NOR2_X2 port map( A1 => n13675, A2 => n13669, ZN => n14003);
   U1170 : AOI22_X2 port map( A1 => n6085, A2 => n6767, B1 => n6084, B2 => n314
                           , ZN => n7757);
   U1174 : XNOR2_X2 port map( A => n20656, B => n20655, ZN => n22977);
   U1177 : NOR2_X2 port map( A1 => n10324, A2 => n10323, ZN => n12189);
   U1200 : BUF_X1 port map( A => n9450, Z => n24511);
   U1202 : OR2_X1 port map( A1 => n6277, A2 => n440, ZN => n24277);
   U1205 : CLKBUF_X1 port map( A => Key(82), Z => n24287);
   U1225 : INV_X1 port map( A => n23411, ZN => n24074);
   U1237 : AND2_X1 port map( A1 => n4947, A2 => n4949, ZN => n24351);
   U1241 : AND3_X1 port map( A1 => n3087, A2 => n4102, A3 => n4099, ZN => 
                           n23220);
   U1250 : INV_X1 port map( A => n23077, ZN => n24075);
   U1251 : AND3_X1 port map( A1 => n24242, A2 => n747, A3 => n3939, ZN => 
                           n23125);
   U1252 : OR2_X1 port map( A1 => n21827, A2 => n3890, ZN => n24307);
   U1257 : OR3_X1 port map( A1 => n22212, A2 => n22211, A3 => n22210, ZN => 
                           n22213);
   U1259 : AND2_X1 port map( A1 => n24115, A2 => n24113, ZN => n22046);
   U1276 : OAI211_X1 port map( C1 => n20564, C2 => n25221, A => n4009, B => 
                           n19734, ZN => n24491);
   U1285 : NOR2_X1 port map( A1 => n20078, A2 => n20077, ZN => n20912);
   U1294 : OR2_X1 port map( A1 => n19988, A2 => n24315, ZN => n24154);
   U1295 : INV_X1 port map( A => n20381, ZN => n24128);
   U1302 : AOI21_X1 port map( B1 => n20232, B2 => n25205, A => n20231, ZN => 
                           n20240);
   U1309 : INV_X1 port map( A => n20615, ZN => n24076);
   U1311 : INV_X1 port map( A => n20360, ZN => n24078);
   U1312 : BUF_X1 port map( A => n20618, Z => n24338);
   U1315 : AND3_X1 port map( A1 => n19447, A2 => n19448, A3 => n24136, ZN => 
                           n20169);
   U1325 : INV_X1 port map( A => n3989, ZN => n19036);
   U1333 : XNOR2_X1 port map( A => n18566, B => n18565, ZN => n19417);
   U1362 : INV_X1 port map( A => n19071, ZN => n24079);
   U1379 : XNOR2_X1 port map( A => n18249, B => n18250, ZN => n19546);
   U1384 : INV_X1 port map( A => n372, ZN => n16775);
   U1395 : INV_X1 port map( A => n17014, ZN => n367);
   U1422 : OR2_X1 port map( A1 => n5024, A2 => n14839, ZN => n24149);
   U1445 : INV_X1 port map( A => n1122, ZN => n16286);
   U1446 : OR2_X1 port map( A1 => n15549, A2 => n25446, ZN => n16068);
   U1452 : INV_X1 port map( A => n16352, ZN => n24080);
   U1516 : AND2_X1 port map( A1 => n1203, A2 => n1204, ZN => n24259);
   U1517 : NAND2_X1 port map( A1 => n2774, A2 => n12544, ZN => n15169);
   U1537 : NOR2_X1 port map( A1 => n24503, A2 => n14099, ZN => n24181);
   U1538 : INV_X1 port map( A => n177, ZN => n14083);
   U1539 : AND2_X1 port map( A1 => n13969, A2 => n13966, ZN => n13599);
   U1542 : AND2_X1 port map( A1 => n14065, A2 => n14064, ZN => n24135);
   U1609 : OR2_X1 port map( A1 => n13854, A2 => n13853, ZN => n177);
   U1690 : AOI21_X1 port map( B1 => n3935, B2 => n12653, A => n12724, ZN => 
                           n13670);
   U1693 : AND2_X1 port map( A1 => n13056, A2 => n12795, ZN => n12526);
   U1695 : INV_X1 port map( A => n11993, ZN => n24241);
   U1704 : XNOR2_X1 port map( A => n11313, B => n11312, ZN => n12995);
   U1710 : INV_X1 port map( A => n11263, ZN => n12225);
   U1771 : INV_X1 port map( A => n11149, ZN => n24286);
   U1811 : INV_X1 port map( A => n11209, ZN => n24082);
   U1821 : AND2_X1 port map( A1 => n11130, A2 => n10714, ZN => n24164);
   U1852 : NOR2_X1 port map( A1 => n9467, A2 => n9466, ZN => n24345);
   U1890 : OR2_X1 port map( A1 => n24534, A2 => n9991, ZN => n9659);
   U1911 : INV_X1 port map( A => n9898, ZN => n24083);
   U1915 : INV_X1 port map( A => n9934, ZN => n24084);
   U1916 : XNOR2_X1 port map( A => n6222, B => n6221, ZN => n9461);
   U1917 : INV_X1 port map( A => n9842, ZN => n24085);
   U1933 : INV_X1 port map( A => n10147, ZN => n24087);
   U1968 : OR2_X1 port map( A1 => n7721, A2 => n24072, ZN => n7727);
   U2069 : OR2_X1 port map( A1 => n6923, A2 => n1175, ZN => n24147);
   U2081 : OR2_X1 port map( A1 => n6940, A2 => n5908, ZN => n6943);
   U2085 : INV_X1 port map( A => n6969, ZN => n24089);
   U2086 : OR2_X1 port map( A1 => n6390, A2 => n6976, ZN => n24262);
   U2088 : BUF_X1 port map( A => n5795, Z => n6619);
   U2128 : OR2_X1 port map( A1 => n6373, A2 => n5824, ZN => n24177);
   U2134 : INV_X1 port map( A => n6112, ZN => n24125);
   U2139 : BUF_X1 port map( A => n6368, Z => n6997);
   U2211 : AND2_X1 port map( A1 => n6123, A2 => n6838, ZN => n24255);
   U2316 : INV_X1 port map( A => n7762, ZN => n7648);
   U2334 : OR2_X1 port map( A1 => n7899, A2 => n24103, ZN => n2758);
   U2338 : BUF_X1 port map( A => n7294, Z => n8015);
   U2341 : OR2_X1 port map( A1 => n7765, A2 => n7648, ZN => n24119);
   U2350 : XNOR2_X1 port map( A => n8333, B => n8069, ZN => n8865);
   U2376 : CLKBUF_X1 port map( A => n9496, Z => n10089);
   U2388 : INV_X1 port map( A => n11302, ZN => n95);
   U2417 : AND2_X1 port map( A1 => n24345, A2 => n10887, ZN => n24141);
   U2437 : OAI211_X1 port map( C1 => n8804, C2 => n9973, A => n8803, B => 
                           n24225, ZN => n11518);
   U2460 : OAI21_X1 port map( B1 => n1871, B2 => n9691, A => n9690, ZN => n1357
                           );
   U2473 : INV_X1 port map( A => n9367, ZN => n9825);
   U2478 : CLKBUF_X1 port map( A => n10533, Z => n11145);
   U2510 : OR2_X1 port map( A1 => n10767, A2 => n10889, ZN => n4654);
   U2539 : MUX2_X1 port map( A => n10228, B => n10227, S => n10789, Z => n10231
                           );
   U2587 : OR2_X1 port map( A1 => n13234, A2 => n12935, ZN => n148);
   U2604 : NOR2_X1 port map( A1 => n13014, A2 => n13013, ZN => n13248);
   U2656 : OR2_X1 port map( A1 => n14190, A2 => n24347, ZN => n24186);
   U2660 : XNOR2_X1 port map( A => n11994, B => n24241, ZN => n24443);
   U2686 : AND2_X1 port map( A1 => n4925, A2 => n4924, ZN => n5472);
   U2695 : AND2_X1 port map( A1 => n14252, A2 => n14251, ZN => n24301);
   U2719 : XNOR2_X1 port map( A => n3862, B => n3861, ZN => n24487);
   U2778 : OAI211_X1 port map( C1 => n12532, C2 => n12531, A => n3315, B => 
                           n3314, ZN => n14269);
   U2788 : OR2_X1 port map( A1 => n13563, A2 => n13564, ZN => n24121);
   U2809 : OR2_X1 port map( A1 => n13773, A2 => n13774, ZN => n82);
   U2821 : NAND3_X1 port map( A1 => n598, A2 => n4907, A3 => n597, ZN => n14311
                           );
   U2826 : OR2_X1 port map( A1 => n13436, A2 => n14106, ZN => n24519);
   U2841 : AOI21_X1 port map( B1 => n13849, B2 => n13848, A => n24135, ZN => 
                           n14611);
   U2855 : NAND2_X1 port map( A1 => n13816, A2 => n13817, ZN => n15094);
   U2866 : XNOR2_X1 port map( A => n15095, B => n15098, ZN => n12);
   U2875 : OAI211_X1 port map( C1 => n12703, C2 => n13785, A => n12702, B => 
                           n12701, ZN => n15358);
   U2876 : INV_X1 port map( A => n1867, ZN => n15321);
   U2886 : AND2_X1 port map( A1 => n24170, A2 => n1261, ZN => n24169);
   U2932 : OAI21_X1 port map( B1 => n24249, B2 => n15625, A => n24248, ZN => 
                           n15627);
   U2933 : OR2_X1 port map( A1 => n16064, A2 => n16060, ZN => n24227);
   U2950 : BUF_X1 port map( A => n4897, Z => n16508);
   U2958 : OR2_X1 port map( A1 => n17161, A2 => n17162, ZN => n24250);
   U3017 : AND2_X2 port map( A1 => n995, A2 => n646, ZN => n17335);
   U3021 : OAI21_X1 port map( B1 => n2233, B2 => n2234, A => n5406, ZN => n4743
                           );
   U3023 : AND2_X1 port map( A1 => n17357, A2 => n16877, ZN => n118);
   U3033 : BUF_X1 port map( A => n18832, Z => n24478);
   U3044 : XNOR2_X1 port map( A => n39, B => n16037, ZN => n17814);
   U3045 : CLKBUF_X1 port map( A => n19370, Z => n24361);
   U3090 : OR2_X1 port map( A1 => n19451, A2 => n19452, ZN => n24137);
   U3107 : AOI21_X1 port map( B1 => n4436, B2 => n18917, A => n19146, ZN => 
                           n19148);
   U3114 : OR2_X1 port map( A1 => n19522, A2 => n19523, ZN => n24252);
   U3119 : INV_X1 port map( A => n19031, ZN => n19029);
   U3125 : OR2_X1 port map( A1 => n1506, A2 => n19210, ZN => n160);
   U3129 : AOI22_X1 port map( A1 => n1307, A2 => n1306, B1 => n19423, B2 => 
                           n19167, ZN => n1305);
   U3167 : NOR2_X1 port map( A1 => n24078, A2 => n20913, ZN => n20482);
   U3191 : OR2_X1 port map( A1 => n20514, A2 => n20517, ZN => n22);
   U3202 : NOR2_X1 port map( A1 => n4287, A2 => n18938, ZN => n18940);
   U3218 : BUF_X1 port map( A => n20346, Z => n24414);
   U3223 : AOI22_X1 port map( A1 => n20569, A2 => n20617, B1 => n20614, B2 => 
                           n20618, ZN => n20327);
   U3227 : OR2_X1 port map( A1 => n20452, A2 => n20960, ZN => n24189);
   U3231 : INV_X1 port map( A => n20022, ZN => n20567);
   U3234 : AND2_X1 port map( A1 => n20341, A2 => n19709, ZN => n20665);
   U3237 : INV_X1 port map( A => n22361, ZN => n24114);
   U3246 : OR2_X1 port map( A1 => n22792, A2 => n2397, ZN => n4080);
   U3248 : OR2_X1 port map( A1 => n22946, A2 => n2674, ZN => n2673);
   U3260 : OR2_X1 port map( A1 => n24877, A2 => n23014, ZN => n23463);
   U3299 : OR2_X1 port map( A1 => n2987, A2 => n21825, ZN => n580);
   U3304 : OR2_X1 port map( A1 => n22578, A2 => n24075, ZN => n24278);
   U3327 : CLKBUF_X1 port map( A => Key(183), Z => n2745);
   U3344 : OAI211_X1 port map( C1 => n22959, C2 => n1259, A => n1258, B => 
                           n1257, ZN => n23379);
   U3347 : OR2_X1 port map( A1 => n23544, A2 => n23537, ZN => n23549);
   U3354 : CLKBUF_X1 port map( A => Key(185), Z => n22702);
   U3359 : XNOR2_X1 port map( A => Key(25), B => Plaintext(25), ZN => n6533);
   U3365 : AND2_X1 port map( A1 => n6827, A2 => n6598, ZN => n24090);
   U3371 : INV_X1 port map( A => n20578, ZN => n24194);
   U3373 : INV_X1 port map( A => n3926, ZN => n24257);
   U3410 : AND2_X1 port map( A1 => n6959, A2 => n6703, ZN => n24091);
   U3418 : INV_X1 port map( A => n3469, ZN => n24103);
   U3422 : XOR2_X1 port map( A => n9056, B => n9055, Z => n24092);
   U3425 : INV_X1 port map( A => n10406, ZN => n24118);
   U3426 : NAND3_X1 port map( A1 => n9346, A2 => n9600, A3 => n9599, ZN => 
                           n24093);
   U3427 : OR2_X1 port map( A1 => n13045, A2 => n13038, ZN => n24094);
   U3431 : INV_X1 port map( A => n12935, ZN => n24220);
   U3449 : AND2_X1 port map( A1 => n1969, A2 => n1967, ZN => n24095);
   U3460 : OR2_X1 port map( A1 => n13235, A2 => n13234, ZN => n24096);
   U3465 : AND2_X1 port map( A1 => n14419, A2 => n2863, ZN => n24097);
   U3468 : INV_X1 port map( A => n16247, ZN => n24162);
   U3485 : XNOR2_X1 port map( A => n14576, B => n14577, ZN => n16147);
   U3512 : INV_X1 port map( A => n16147, ZN => n24249);
   U3527 : XOR2_X1 port map( A => n14624, B => n14623, Z => n24098);
   U3551 : INV_X1 port map( A => n19456, ZN => n24172);
   U3587 : XNOR2_X1 port map( A => n17871, B => n17870, ZN => n17872);
   U3594 : INV_X1 port map( A => n20491, ZN => n24275);
   U3600 : AND3_X1 port map( A1 => n87, A2 => n3032, A3 => n3794, ZN => n24100)
                           ;
   U3603 : OR2_X1 port map( A1 => n20960, A2 => n24354, ZN => n24101);
   U3612 : NAND2_X1 port map( A1 => n7232, A2 => n7230, ZN => n7899);
   U3615 : OAI211_X1 port map( C1 => n421, C2 => n9836, A => n4302, B => n10098
                           , ZN => n24104);
   U3673 : NAND2_X1 port map( A1 => n356, A2 => n18927, ZN => n18928);
   U3688 : OAI22_X1 port map( A1 => n16069, A2 => n15694, B1 => n16068, B2 => 
                           n16067, ZN => n16070);
   U3697 : NAND2_X1 port map( A1 => n16063, A2 => n16062, ZN => n16069);
   U3726 : NAND3_X2 port map( A1 => n2981, A2 => n24107, A3 => n24106, ZN => 
                           n23554);
   U3727 : NAND2_X1 port map( A1 => n22096, A2 => n22890, ZN => n24106);
   U3738 : NAND2_X1 port map( A1 => n22097, A2 => n22729, ZN => n24107);
   U3739 : NAND2_X1 port map( A1 => n5291, A2 => n7054, ZN => n5294);
   U3795 : XNOR2_X1 port map( A => n15422, B => n24108, ZN => n12451);
   U3834 : XNOR2_X1 port map( A => n14892, B => n3158, ZN => n24108);
   U3853 : NAND3_X1 port map( A1 => n20567, A2 => n20094, A3 => n20560, ZN => 
                           n24109);
   U3890 : OAI21_X1 port map( B1 => n19213, B2 => n25392, A => n24110, ZN => 
                           n3811);
   U3894 : NAND3_X1 port map( A1 => n1212, A2 => n24312, A3 => n19361, ZN => 
                           n24110);
   U3928 : NAND2_X1 port map( A1 => n16133, A2 => n16074, ZN => n17159);
   U3966 : NAND2_X1 port map( A1 => n19446, A2 => n18990, ZN => n3989);
   U3967 : NAND2_X1 port map( A1 => n13628, A2 => n177, ZN => n176);
   U4003 : OR2_X1 port map( A1 => n16186, A2 => n15970, ZN => n13941);
   U4062 : XNOR2_X1 port map( A => n24112, B => n455, ZN => Ciphertext(4));
   U4084 : NAND2_X1 port map( A1 => n1925, A2 => n1926, ZN => n6614);
   U4106 : NAND2_X1 port map( A1 => n245, A2 => n24114, ZN => n24113);
   U4108 : AOI21_X1 port map( B1 => n22361, B2 => n22356, A => n21839, ZN => 
                           n24115);
   U4125 : INV_X1 port map( A => n4520, ZN => n10926);
   U4146 : NAND2_X1 port map( A1 => n10994, A2 => n10993, ZN => n4520);
   U4168 : NOR2_X1 port map( A1 => n17451, A2 => n523, ZN => n17456);
   U4169 : NOR2_X2 port map( A1 => n1900, A2 => n5335, ZN => n12404);
   U4187 : OR2_X1 port map( A1 => n9387, A2 => n9959, ZN => n2875);
   U4191 : NAND3_X1 port map( A1 => n4936, A2 => n10730, A3 => n10480, ZN => 
                           n2831);
   U4192 : NAND3_X1 port map( A1 => n16756, A2 => n16957, A3 => n17414, ZN => 
                           n16758);
   U4198 : NAND3_X2 port map( A1 => n24119, A2 => n24120, A3 => n7308, ZN => 
                           n8799);
   U4201 : NAND2_X1 port map( A1 => n2848, A2 => n7306, ZN => n24120);
   U4205 : XNOR2_X1 port map( A => n5215, B => n15174, ZN => n14494);
   U4207 : AOI22_X2 port map( A1 => n178, A2 => n14203, B1 => n14202, B2 => 
                           n14944, ZN => n15174);
   U4242 : NAND3_X1 port map( A1 => n4774, A2 => n16532, A3 => n17164, ZN => 
                           n16265);
   U4257 : AOI22_X1 port map( A1 => n16052, A2 => n16051, B1 => n16053, B2 => 
                           n16508, ZN => n16054);
   U4267 : BUF_X1 port map( A => n14100, Z => n24375);
   U4283 : BUF_X1 port map( A => n23479, Z => n24336);
   U4286 : NAND2_X1 port map( A1 => n13562, A2 => n24121, ZN => n14667);
   U4301 : NAND3_X1 port map( A1 => n23896, A2 => n23906, A3 => n23903, ZN => 
                           n23872);
   U4318 : NAND3_X1 port map( A1 => n24124, A2 => n24123, A3 => n6608, ZN => 
                           n7767);
   U4338 : NAND3_X1 port map( A1 => n6110, A2 => n6606, A3 => n6611, ZN => 
                           n24123);
   U4413 : NAND2_X1 port map( A1 => n24125, A2 => n6610, ZN => n24124);
   U4502 : NAND3_X1 port map( A1 => n14271, A2 => n14274, A3 => n13840, ZN => 
                           n13622);
   U4525 : OR2_X1 port map( A1 => n16243, A2 => n15707, ZN => n16241);
   U4545 : AND2_X1 port map( A1 => n648, A2 => n16064, ZN => n24233);
   U4551 : NAND3_X1 port map( A1 => n24326, A2 => n19395, A3 => n19393, ZN => 
                           n1458);
   U4641 : NAND3_X1 port map( A1 => n20507, A2 => n20216, A3 => n25223, ZN => 
                           n1808);
   U4747 : AND2_X1 port map( A1 => n7985, A2 => n7984, ZN => n24197);
   U4824 : NAND2_X1 port map( A1 => n24101, A2 => n24128, ZN => n24127);
   U4878 : NAND3_X1 port map( A1 => n17441, A2 => n17442, A3 => n2549, ZN => 
                           n139);
   U4884 : XNOR2_X1 port map( A => n24131, B => n24130, ZN => Ciphertext(131));
   U4898 : INV_X1 port map( A => n2228, ZN => n24130);
   U4926 : NAND2_X1 port map( A1 => n24133, A2 => n24132, ZN => n24131);
   U4953 : NAND2_X1 port map( A1 => n22748, A2 => n22749, ZN => n24132);
   U5025 : NAND2_X1 port map( A1 => n22750, A2 => n25405, ZN => n24133);
   U5087 : NAND2_X1 port map( A1 => n8023, A2 => n7531, ZN => n4708);
   U5092 : OAI21_X2 port map( B1 => n14072, B2 => n24134, A => n14070, ZN => 
                           n15497);
   U5115 : NAND2_X1 port map( A1 => n14066, A2 => n14264, ZN => n24134);
   U5130 : NAND3_X1 port map( A1 => n4106, A2 => n4053, A3 => n6925, ZN => 
                           n3311);
   U5178 : NAND2_X1 port map( A1 => n7514, A2 => n7973, ZN => n2177);
   U5196 : NAND3_X1 port map( A1 => n9133, A2 => n9132, A3 => n9951, ZN => 
                           n1092);
   U5205 : NAND2_X1 port map( A1 => n9947, A2 => n9389, ZN => n9133);
   U5213 : NAND3_X1 port map( A1 => n1879, A2 => n7854, A3 => n1880, ZN => 
                           n6419);
   U5344 : OR2_X1 port map( A1 => n20449, A2 => n20450, ZN => n24188);
   U5390 : NAND2_X1 port map( A1 => n16177, A2 => n15657, ZN => n15992);
   U5399 : NAND3_X1 port map( A1 => n19449, A2 => n25002, A3 => n24137, ZN => 
                           n24136);
   U5404 : NAND2_X1 port map( A1 => n19018, A2 => n20537, ZN => n19688);
   U5441 : NAND3_X1 port map( A1 => n2386, A2 => n10212, A3 => n10886, ZN => 
                           n10214);
   U5470 : NAND3_X2 port map( A1 => n1735, A2 => n1734, A3 => n6402, ZN => 
                           n7721);
   U5499 : NAND2_X1 port map( A1 => n19918, A2 => n19917, ZN => n24138);
   U5579 : OR2_X1 port map( A1 => n17087, A2 => n16578, ZN => n2813);
   U5605 : NAND2_X1 port map( A1 => n424, A2 => n24139, ZN => n8572);
   U5609 : AND2_X1 port map( A1 => n8571, A2 => n9782, ZN => n24139);
   U5614 : OAI21_X1 port map( B1 => n10544, B2 => n2389, A => n24140, ZN => 
                           n10545);
   U5635 : NAND2_X1 port map( A1 => n2386, A2 => n24141, ZN => n24140);
   U5722 : OAI211_X2 port map( C1 => n16782, C2 => n16859, A => n24143, B => 
                           n3002, ZN => n18103);
   U5734 : NAND2_X1 port map( A1 => n16779, A2 => n16780, ZN => n24143);
   U5757 : OAI211_X1 port map( C1 => n9600, C2 => n24084, A => n9205, B => 
                           n25217, ZN => n24144);
   U5878 : NAND3_X1 port map( A1 => n391, A2 => n14291, A3 => n13909, ZN => 
                           n24146);
   U5890 : NAND3_X1 port map( A1 => n6199, A2 => n6922, A3 => n24147, ZN => 
                           n7294);
   U5956 : NAND2_X1 port map( A1 => n9626, A2 => n10046, ZN => n24148);
   U5970 : NAND2_X2 port map( A1 => n5023, A2 => n24149, ZN => n17607);
   U6031 : NAND2_X1 port map( A1 => n24153, A2 => n24150, ZN => n13457);
   U6134 : NAND2_X1 port map( A1 => n24152, A2 => n24151, ZN => n24150);
   U6136 : NOR2_X1 port map( A1 => n13947, A2 => n14306, ZN => n24151);
   U6196 : INV_X1 port map( A => n13892, ZN => n24152);
   U6281 : NAND2_X1 port map( A1 => n12838, A2 => n12839, ZN => n3010);
   U6372 : NAND3_X1 port map( A1 => n19446, A2 => n19444, A3 => n19445, ZN => 
                           n19447);
   U6404 : NAND2_X1 port map( A1 => n883, A2 => n884, ZN => n24155);
   U6486 : INV_X1 port map( A => n7114, ZN => n5318);
   U6502 : NAND2_X1 port map( A1 => n7762, A2 => n7647, ZN => n7114);
   U6544 : NAND2_X1 port map( A1 => n23875, A2 => n24158, ZN => n23878);
   U6545 : OR2_X1 port map( A1 => n23904, A2 => n23883, ZN => n24158);
   U6556 : NAND2_X1 port map( A1 => n24159, A2 => n19465, ZN => n17890);
   U6569 : NAND2_X1 port map( A1 => n19032, A2 => n19460, ZN => n24159);
   U6575 : AOI22_X1 port map( A1 => n19814, A2 => n20507, B1 => n20510, B2 => 
                           n20218, ZN => n19815);
   U6584 : OAI21_X1 port map( B1 => n22184, B2 => n1336, A => n24160, ZN => 
                           n2296);
   U6659 : NAND2_X1 port map( A1 => n1336, A2 => n22239, ZN => n24160);
   U6706 : NAND2_X1 port map( A1 => n24161, A2 => n9575, ZN => n11845);
   U6711 : NAND3_X1 port map( A1 => n24167, A2 => n24166, A3 => n2388, ZN => 
                           n24161);
   U6728 : INV_X1 port map( A => n16252, ZN => n24163);
   U6750 : NAND2_X1 port map( A1 => n10840, A2 => n24164, ZN => n10717);
   U6787 : AND2_X2 port map( A1 => n788, A2 => n2282, ZN => n18388);
   U6818 : NAND3_X1 port map( A1 => n17366, A2 => n17363, A3 => n17364, ZN => 
                           n2452);
   U6907 : INV_X1 port map( A => n24383, ZN => n17755);
   U6914 : NAND3_X1 port map( A1 => n2790, A2 => n16259, A3 => n2789, ZN => 
                           n24383);
   U6915 : NAND2_X1 port map( A1 => n10884, A2 => n10302, ZN => n24166);
   U6930 : INV_X1 port map( A => n10884, ZN => n24168);
   U6943 : NAND2_X1 port map( A1 => n2008, A2 => n5907, ZN => n2007);
   U7002 : NAND2_X1 port map( A1 => n16122, A2 => n16155, ZN => n16158);
   U7012 : NAND2_X1 port map( A1 => n9368, A2 => n9398, ZN => n9367);
   U7037 : INV_X1 port map( A => n17277, ZN => n24300);
   U7076 : INV_X1 port map( A => n15611, ZN => n24170);
   U7134 : AOI21_X2 port map( B1 => n13442, B2 => n13443, A => n755, ZN => 
                           n15505);
   U7167 : INV_X1 port map( A => n523, ZN => n17460);
   U7170 : NAND2_X1 port map( A1 => n3451, A2 => n16359, ZN => n16361);
   U7255 : NAND2_X1 port map( A1 => n24597, A2 => n7312, ZN => n24198);
   U7260 : NAND2_X1 port map( A1 => n7582, A2 => n7584, ZN => n7312);
   U7263 : OR2_X1 port map( A1 => n17463, A2 => n16846, ZN => n17465);
   U7268 : NAND2_X1 port map( A1 => n24243, A2 => n24244, ZN => n18975);
   U7293 : NAND2_X1 port map( A1 => n508, A2 => n13953, ZN => n14159);
   U7303 : NAND2_X1 port map( A1 => n11216, A2 => n10623, ZN => n10620);
   U7368 : NAND2_X1 port map( A1 => n24178, A2 => n24177, ZN => n6790);
   U7380 : NAND2_X1 port map( A1 => n6374, A2 => n6375, ZN => n24178);
   U7513 : XNOR2_X1 port map( A => n24179, B => n18050, ZN => n18052);
   U7515 : XNOR2_X1 port map( A => n18567, B => n17663, ZN => n24179);
   U7524 : NAND2_X1 port map( A1 => n14097, A2 => n24180, ZN => n14103);
   U7553 : NAND2_X1 port map( A1 => n24182, A2 => n24181, ZN => n24180);
   U7567 : INV_X1 port map( A => n4894, ZN => n24182);
   U7585 : NAND2_X1 port map( A1 => n2909, A2 => n2907, ZN => n24183);
   U7597 : NAND2_X1 port map( A1 => n16619, A2 => n16620, ZN => n16552);
   U7601 : OAI21_X1 port map( B1 => n15694, B2 => n25446, A => n16060, ZN => 
                           n648);
   U7646 : NAND2_X1 port map( A1 => n3456, A2 => n22221, ZN => n24184);
   U7692 : NAND2_X1 port map( A1 => n15562, A2 => n24506, ZN => n24185);
   U7694 : NAND2_X1 port map( A1 => n19752, A2 => n19987, ZN => n21067);
   U7731 : NAND2_X1 port map( A1 => n16344, A2 => n24187, ZN => n16346);
   U7816 : NAND2_X1 port map( A1 => n16341, A2 => n16342, ZN => n24187);
   U7853 : AOI22_X2 port map( A1 => n10204, A2 => n10451, B1 => n9375, B2 => 
                           n4505, ZN => n12249);
   U7868 : NAND3_X1 port map( A1 => n2082, A2 => n7826, A3 => n2081, ZN => 
                           n2080);
   U7882 : NAND2_X1 port map( A1 => n249, A2 => n6848, ZN => n7028);
   U7897 : NAND2_X1 port map( A1 => n24191, A2 => n24190, ZN => n18964);
   U7899 : NAND2_X1 port map( A1 => n18957, A2 => n19471, ZN => n24190);
   U7936 : NAND2_X1 port map( A1 => n18958, A2 => n18945, ZN => n24191);
   U7965 : XNOR2_X1 port map( A => n24192, B => n18239, ZN => n18493);
   U7967 : NAND2_X1 port map( A1 => n12960, A2 => n13339, ZN => n12577);
   U8020 : OAI21_X1 port map( B1 => n20194, B2 => n24194, A => n24193, ZN => 
                           n20582);
   U8022 : NAND2_X1 port map( A1 => n20194, A2 => n20576, ZN => n24193);
   U8063 : NAND3_X1 port map( A1 => n690, A2 => n14101, A3 => n689, ZN => n672)
                           ;
   U8142 : NAND2_X1 port map( A1 => n5464, A2 => n2090, ZN => n24195);
   U8143 : NAND3_X1 port map( A1 => n17287, A2 => n17289, A3 => n17288, ZN => 
                           n24196);
   U8159 : NAND2_X1 port map( A1 => n7826, A2 => n24197, ZN => n7831);
   U8223 : NAND3_X1 port map( A1 => n7018, A2 => n24200, A3 => n24199, ZN => 
                           n7965);
   U8237 : NAND3_X1 port map( A1 => n7015, A2 => n7016, A3 => n7014, ZN => 
                           n24199);
   U8239 : NAND2_X1 port map( A1 => n24090, A2 => n6824, ZN => n24200);
   U8241 : OAI211_X1 port map( C1 => n15535, C2 => n16038, A => n1718, B => 
                           n24098, ZN => n17158);
   U8257 : NAND2_X1 port map( A1 => n9435, A2 => n9634, ZN => n10038);
   U8275 : NAND2_X1 port map( A1 => n24202, A2 => n16708, ZN => n16374);
   U8276 : NAND2_X1 port map( A1 => n16372, A2 => n16616, ZN => n24202);
   U8281 : NAND2_X1 port map( A1 => n16170, A2 => n16426, ZN => n706);
   U8298 : INV_X1 port map( A => n7926, ZN => n24203);
   U8309 : NAND2_X1 port map( A1 => n6555, A2 => n6554, ZN => n7926);
   U8336 : NOR2_X1 port map( A1 => n24012, A2 => n24011, ZN => n24204);
   U8387 : OAI21_X1 port map( B1 => n7607, B2 => n7608, A => n7606, ZN => 
                           n24205);
   U8472 : NOR2_X1 port map( A1 => n4541, A2 => n24352, ZN => n15541);
   U8488 : NAND2_X1 port map( A1 => n20125, A2 => n20547, ZN => n5638);
   U8505 : NAND2_X1 port map( A1 => n266, A2 => n4004, ZN => n16316);
   U8522 : XNOR2_X1 port map( A => n20792, B => n21713, ZN => n19955);
   U8548 : OAI22_X1 port map( A1 => n11086, A2 => n11085, B1 => n11084, B2 => 
                           n418, ZN => n1263);
   U8559 : NAND2_X1 port map( A1 => n5559, A2 => n10890, ZN => n11086);
   U8568 : OAI211_X1 port map( C1 => n9340, C2 => n10156, A => n3988, B => 
                           n10154, ZN => n10336);
   U8587 : OAI211_X1 port map( C1 => n1251, C2 => n19460, A => n24209, B => 
                           n19465, ZN => n18741);
   U8598 : NAND2_X1 port map( A1 => n1251, A2 => n18979, ZN => n24209);
   U8617 : NAND3_X1 port map( A1 => n19470, A2 => n18959, A3 => n18960, ZN => 
                           n5099);
   U8619 : XNOR2_X1 port map( A => n21572, B => n21135, ZN => n21463);
   U8625 : AND2_X2 port map( A1 => n24211, A2 => n24210, ZN => n21135);
   U8636 : NAND2_X1 port map( A1 => n18743, A2 => n20183, ZN => n24210);
   U8643 : NAND2_X1 port map( A1 => n18742, A2 => n19862, ZN => n24211);
   U8647 : OR2_X1 port map( A1 => n10148, A2 => n25207, ZN => n9522);
   U8651 : NAND3_X1 port map( A1 => n9746, A2 => n24535, A3 => n25121, ZN => 
                           n24212);
   U8652 : AND3_X2 port map( A1 => n24214, A2 => n3728, A3 => n24213, ZN => 
                           n11914);
   U8671 : INV_X1 port map( A => n8032, ZN => n24214);
   U8703 : NAND3_X1 port map( A1 => n10292, A2 => n10840, A3 => n10293, ZN => 
                           n10294);
   U8771 : NAND2_X1 port map( A1 => n11098, A2 => n11097, ZN => n24215);
   U8772 : NAND2_X1 port map( A1 => n102, A2 => n9490, ZN => n10914);
   U8809 : NAND2_X1 port map( A1 => n16485, A2 => n25238, ZN => n15698);
   U8834 : OR2_X1 port map( A1 => n6135, A2 => n1798, ZN => n2448);
   U8898 : NAND3_X1 port map( A1 => n1594, A2 => n9282, A3 => n2953, ZN => 
                           n9283);
   U8899 : NAND2_X1 port map( A1 => n2248, A2 => n2249, ZN => n19698);
   U8925 : BUF_X1 port map( A => n17421, Z => n24330);
   U8926 : AOI22_X1 port map( A1 => n23847, A2 => n24218, B1 => n23850, B2 => 
                           n23849, ZN => n23856);
   U8959 : NAND3_X1 port map( A1 => n23851, A2 => n25240, A3 => n3183, ZN => 
                           n24218);
   U8961 : NAND2_X1 port map( A1 => n24096, A2 => n24219, ZN => n34);
   U8972 : AOI21_X1 port map( B1 => n4499, B2 => n13234, A => n24220, ZN => 
                           n24219);
   U9054 : NOR2_X1 port map( A1 => n25393, A2 => n24221, ZN => n1886);
   U9055 : NAND2_X1 port map( A1 => n24222, A2 => n9772, ZN => n24221);
   U9087 : INV_X1 port map( A => n10109, ZN => n24222);
   U9108 : OAI211_X1 port map( C1 => n11122, C2 => n11123, A => n24223, B => 
                           n11121, ZN => n10462);
   U9122 : INV_X1 port map( A => n10850, ZN => n24223);
   U9153 : NOR2_X2 port map( A1 => n2994, A2 => n9230, ZN => n10850);
   U9231 : AND2_X2 port map( A1 => n24525, A2 => n3153, ZN => n7217);
   U9242 : NAND2_X1 port map( A1 => n14154, A2 => n2775, ZN => n1025);
   U9287 : NAND2_X1 port map( A1 => n7346, A2 => n7349, ZN => n24224);
   U9298 : INV_X1 port map( A => n17197, ZN => n16869);
   U9310 : NAND2_X1 port map( A1 => n17399, A2 => n17198, ZN => n17197);
   U9327 : NAND2_X1 port map( A1 => n9615, A2 => n9757, ZN => n24225);
   U9338 : INV_X1 port map( A => n6575, ZN => n443);
   U9348 : NAND2_X1 port map( A1 => n24089, A2 => n6575, ZN => n4973);
   U9357 : NAND3_X1 port map( A1 => n5596, A2 => n4054, A3 => n24226, ZN => 
                           n17341);
   U9379 : NAND3_X1 port map( A1 => n613, A2 => n16062, A3 => n24227, ZN => 
                           n24226);
   U9418 : NAND2_X1 port map( A1 => n16780, A2 => n17241, ZN => n24229);
   U9440 : NAND2_X1 port map( A1 => n3661, A2 => n3662, ZN => n3660);
   U9570 : OAI21_X1 port map( B1 => n16141, B2 => n24231, A => n24230, ZN => 
                           n16144);
   U9584 : NAND2_X1 port map( A1 => n16141, A2 => n16412, ZN => n24230);
   U9591 : INV_X1 port map( A => n16140, ZN => n24231);
   U9612 : NAND2_X1 port map( A1 => n19550, A2 => n19549, ZN => n19551);
   U9660 : OAI22_X1 port map( A1 => n19546, A2 => n19185, B1 => n24929, B2 => 
                           n19186, ZN => n19550);
   U9673 : AOI21_X2 port map( B1 => n649, B2 => n15694, A => n24233, ZN => 
                           n16550);
   U9717 : NAND2_X1 port map( A1 => n24234, A2 => n6762, ZN => n6763);
   U9738 : NAND2_X1 port map( A1 => n1454, A2 => n7460, ZN => n24234);
   U9816 : NAND2_X1 port map( A1 => n3219, A2 => n5678, ZN => n11310);
   U9818 : NAND2_X1 port map( A1 => n3220, A2 => n24168, ZN => n3219);
   U9833 : NAND2_X2 port map( A1 => n10773, A2 => n10776, ZN => n11101);
   U9836 : NAND2_X1 port map( A1 => n9494, A2 => n10020, ZN => n10773);
   U9858 : AND3_X2 port map( A1 => n22470, A2 => n22471, A3 => n22469, ZN => 
                           n23120);
   U9865 : NAND2_X1 port map( A1 => n24238, A2 => n24236, ZN => n22850);
   U9890 : NOR2_X1 port map( A1 => n22901, A2 => n22900, ZN => n24237);
   U9927 : INV_X1 port map( A => n22842, ZN => n24239);
   U9943 : INV_X1 port map( A => n16782, ZN => n16777);
   U9965 : NAND2_X1 port map( A1 => n17346, A2 => n17341, ZN => n16782);
   U9975 : NAND2_X1 port map( A1 => n3213, A2 => n22972, ZN => n21891);
   U9984 : NAND3_X1 port map( A1 => n10207, A2 => n10206, A3 => n10434, ZN => 
                           n11263);
   U10081 : NAND2_X1 port map( A1 => n24240, A2 => n10836, ZN => n547);
   U10085 : NAND2_X1 port map( A1 => n10276, A2 => n10275, ZN => n24240);
   U10141 : NAND3_X1 port map( A1 => n13065, A2 => n13162, A3 => n12736, ZN => 
                           n2859);
   U10150 : XNOR2_X1 port map( A => n1821, B => n11991, ZN => n11994);
   U10173 : OR2_X1 port map( A1 => n2464, A2 => n18809, ZN => n18166);
   U10174 : NAND2_X1 port map( A1 => n16775, A2 => n17048, ZN => n1908);
   U10197 : NAND2_X1 port map( A1 => n22466, A2 => n3938, ZN => n24242);
   U10211 : XNOR2_X2 port map( A => n20809, B => n20810, ZN => n22462);
   U10233 : NAND2_X1 port map( A1 => n16923, A2 => n16924, ZN => n16926);
   U10235 : NAND2_X1 port map( A1 => n17320, A2 => n17321, ZN => n16924);
   U10288 : NAND2_X1 port map( A1 => n7009, A2 => n7006, ZN => n5982);
   U10298 : NAND2_X1 port map( A1 => n19482, A2 => n19477, ZN => n24243);
   U10326 : NAND2_X1 port map( A1 => n19478, A2 => n24803, ZN => n24244);
   U10463 : NAND2_X2 port map( A1 => n2840, A2 => n12605, ZN => n14852);
   U10464 : NAND3_X2 port map( A1 => n3463, A2 => n5640, A3 => n5642, ZN => 
                           n14858);
   U10495 : NAND2_X1 port map( A1 => n4350, A2 => n22336, ZN => n4349);
   U10515 : MUX2_X2 port map( A => n15813, B => n15812, S => n24061, Z => 
                           n17729);
   U10517 : NAND3_X1 port map( A1 => n17001, A2 => n17002, A3 => n17003, ZN => 
                           n17004);
   U10524 : NAND2_X1 port map( A1 => n2613, A2 => n17048, ZN => n17003);
   U10530 : NAND3_X1 port map( A1 => n15949, A2 => n15948, A3 => n15947, ZN => 
                           n17050);
   U10532 : NAND3_X1 port map( A1 => n24246, A2 => n6298, A3 => n6174, ZN => 
                           n6212);
   U10562 : NAND2_X1 port map( A1 => n6209, A2 => n6296, ZN => n24246);
   U10574 : NAND2_X1 port map( A1 => n1730, A2 => n1729, ZN => n24247);
   U10578 : INV_X1 port map( A => n23235, ZN => n5081);
   U10600 : AOI22_X1 port map( A1 => n23245, A2 => n23235, B1 => n23250, B2 => 
                           n23249, ZN => n22650);
   U10606 : NAND3_X1 port map( A1 => n10840, A2 => n5101, A3 => n10470, ZN => 
                           n10472);
   U10618 : NAND2_X1 port map( A1 => n6864, A2 => n7148, ZN => n6865);
   U10619 : NAND2_X1 port map( A1 => n4365, A2 => n4366, ZN => n6864);
   U10634 : NAND2_X1 port map( A1 => n15625, A2 => n16096, ZN => n24248);
   U10639 : NAND2_X1 port map( A1 => n17160, A2 => n24250, ZN => n17169);
   U10670 : NAND3_X1 port map( A1 => n10740, A2 => n10854, A3 => n10858, ZN => 
                           n24251);
   U10696 : NAND2_X1 port map( A1 => n16777, A2 => n17342, ZN => n1883);
   U10715 : OAI22_X1 port map( A1 => n19525, A2 => n19526, B1 => n19521, B2 => 
                           n24252, ZN => n19527);
   U10737 : NAND2_X1 port map( A1 => n6533, A2 => n24253, ZN => n6264);
   U10769 : INV_X1 port map( A => n6530, ZN => n24253);
   U10778 : INV_X1 port map( A => n4199, ZN => n24254);
   U10842 : NOR2_X1 port map( A1 => n7776, A2 => n7526, ZN => n2807);
   U10859 : AOI21_X2 port map( B1 => n6125, B2 => n6124, A => n24255, ZN => 
                           n7776);
   U10882 : AND2_X1 port map( A1 => n9435, A2 => n9433, ZN => n9712);
   U10914 : OAI211_X1 port map( C1 => n6702, C2 => n6553, A => n24256, B => 
                           n6960, ZN => n7930);
   U10917 : NAND2_X1 port map( A1 => n6702, A2 => n24257, ZN => n24256);
   U10931 : NAND3_X1 port map( A1 => n10095, A2 => n10098, A3 => n10099, ZN => 
                           n10101);
   U10935 : XNOR2_X1 port map( A => n11424, B => n2989, ZN => n11425);
   U10962 : NAND2_X1 port map( A1 => n14157, A2 => n13955, ZN => n3303);
   U10969 : OR2_X1 port map( A1 => n12901, A2 => n12928, ZN => n24258);
   U10980 : NAND2_X1 port map( A1 => n10134, A2 => n24026, ZN => n10145);
   U10981 : OAI211_X2 port map( C1 => n10562, C2 => n10561, A => n10560, B => 
                           n4540, ZN => n12200);
   U11025 : NAND2_X1 port map( A1 => n806, A2 => n7962, ZN => n5163);
   U11043 : NAND2_X1 port map( A1 => n24260, A2 => n2972, ZN => n8635);
   U11088 : NAND2_X1 port map( A1 => n6924, A2 => n1176, ZN => n2355);
   U11091 : NAND2_X1 port map( A1 => n9233, A2 => n9234, ZN => n3705);
   U11100 : NAND2_X1 port map( A1 => n12827, A2 => n24476, ZN => n2915);
   U11112 : OAI211_X1 port map( C1 => n21870, C2 => n21869, A => n24261, B => 
                           n21868, ZN => Ciphertext(172));
   U11121 : OAI211_X1 port map( C1 => n21869, C2 => n21866, A => n21865, B => 
                           n21864, ZN => n24261);
   U11148 : NAND2_X1 port map( A1 => n416, A2 => n11038, ZN => n9130);
   U11155 : NAND2_X1 port map( A1 => n24262, A2 => n6067, ZN => n6068);
   U11156 : OAI22_X1 port map( A1 => n22933, A2 => n22853, B1 => n22498, B2 => 
                           n25004, ZN => n21871);
   U11157 : NAND2_X1 port map( A1 => n23336, A2 => n23334, ZN => n22853);
   U11259 : NAND2_X1 port map( A1 => n9935, A2 => n9938, ZN => n24264);
   U11260 : NAND2_X1 port map( A1 => n9936, A2 => n24511, ZN => n24265);
   U11272 : NOR2_X2 port map( A1 => n16724, A2 => n16723, ZN => n2667);
   U11290 : NAND2_X1 port map( A1 => n16721, A2 => n16931, ZN => n24267);
   U11317 : NAND3_X1 port map( A1 => n22669, A2 => n22670, A3 => n22668, ZN => 
                           n22673);
   U11437 : NAND2_X1 port map( A1 => n7590, A2 => n7464, ZN => n7460);
   U11451 : OR2_X2 port map( A1 => n5942, A2 => n5941, ZN => n7590);
   U11551 : XNOR2_X1 port map( A => n24270, B => n8761, ZN => Ciphertext(82));
   U11678 : NAND2_X1 port map( A1 => n19305, A2 => n19306, ZN => n24272);
   U11682 : NAND2_X1 port map( A1 => n19304, A2 => n19133, ZN => n19306);
   U11737 : NAND2_X1 port map( A1 => n24273, A2 => n24091, ZN => n6708);
   U11786 : NAND2_X1 port map( A1 => n6702, A2 => n6705, ZN => n24273);
   U11810 : NAND3_X1 port map( A1 => n6911, A2 => n6916, A3 => n6286, ZN => 
                           n6288);
   U11847 : OR2_X1 port map( A1 => n14052, A2 => n12821, ZN => n12822);
   U11848 : NOR2_X1 port map( A1 => n25059, A2 => n23206, ZN => n4230);
   U11958 : NAND3_X1 port map( A1 => n6064, A2 => n6061, A3 => n6731, ZN => 
                           n2401);
   U12016 : NAND2_X1 port map( A1 => n20482, A2 => n24275, ZN => n24274);
   U12084 : NAND3_X1 port map( A1 => n6028, A2 => n6278, A3 => n25398, ZN => 
                           n24276);
   U12088 : AND2_X1 port map( A1 => n25210, A2 => n16381, ZN => n692);
   U12101 : NAND2_X1 port map( A1 => n25179, A2 => n22578, ZN => n24279);
   U12122 : INV_X1 port map( A => n1797, ZN => n24280);
   U12188 : NAND2_X1 port map( A1 => n24283, A2 => n4804, ZN => n4800);
   U12251 : NAND2_X1 port map( A1 => n7057, A2 => n7738, ZN => n24283);
   U12261 : NAND2_X1 port map( A1 => n24285, A2 => n24284, ZN => n9720);
   U12272 : NAND2_X1 port map( A1 => n11149, A2 => n24479, ZN => n24284);
   U12337 : NAND2_X1 port map( A1 => n10690, A2 => n24286, ZN => n24285);
   U12448 : NAND3_X2 port map( A1 => n24291, A2 => n24288, A3 => n210, ZN => 
                           n21306);
   U12599 : NAND2_X1 port map( A1 => n1936, A2 => n20071, ZN => n24291);
   U12664 : NAND2_X1 port map( A1 => n16241, A2 => n24293, ZN => n24292);
   U12716 : INV_X1 port map( A => n16440, ZN => n24293);
   U12721 : NAND2_X1 port map( A1 => n15945, A2 => n16440, ZN => n24294);
   U12815 : INV_X1 port map( A => n6596, ZN => n6597);
   U12865 : NAND2_X1 port map( A1 => n6823, A2 => n6827, ZN => n6596);
   U12866 : NAND2_X1 port map( A1 => n9131, A2 => n9130, ZN => n24295);
   U12869 : BUF_X1 port map( A => n1363, Z => n24367);
   U12897 : XOR2_X1 port map( A => n112, B => n15075, Z => n24303);
   U12899 : NAND3_X1 port map( A1 => n6607, A2 => n6609, A3 => n6610, ZN => 
                           n4018);
   U12915 : NAND2_X1 port map( A1 => n19208, A2 => n19024, ZN => n835);
   U12952 : OAI21_X1 port map( B1 => n13356, B2 => n13993, A => n24296, ZN => 
                           n13369);
   U12953 : NAND2_X1 port map( A1 => n13993, A2 => n795, ZN => n24296);
   U13053 : NOR2_X2 port map( A1 => n635, A2 => n15559, ZN => n16974);
   U13054 : NAND2_X1 port map( A1 => n5698, A2 => n6323, ZN => n5696);
   U13136 : NAND2_X1 port map( A1 => n1577, A2 => n25064, ZN => n9815);
   U13217 : INV_X1 port map( A => n3554, ZN => n24297);
   U13305 : NAND3_X1 port map( A1 => n17252, A2 => n17254, A3 => n24300, ZN => 
                           n24299);
   U13306 : NAND2_X1 port map( A1 => n2644, A2 => n19608, ZN => n2643);
   U13448 : NAND2_X1 port map( A1 => n328, A2 => n21794, ZN => n5075);
   U13473 : NAND2_X1 port map( A1 => n148, A2 => n546, ZN => n11836);
   U13657 : NAND2_X1 port map( A1 => n17051, A2 => n372, ZN => n3643);
   U13659 : NAND2_X1 port map( A1 => n14250, A2 => n24301, ZN => n14260);
   U13674 : NAND3_X1 port map( A1 => n19388, A2 => n19389, A3 => n19390, ZN => 
                           n191);
   U13812 : NAND3_X1 port map( A1 => n1062, A2 => n14090, A3 => n13607, ZN => 
                           n1061);
   U13816 : NAND2_X1 port map( A1 => n24302, A2 => n14059, ZN => n12614);
   U13817 : NAND2_X1 port map( A1 => n14278, A2 => n14850, ZN => n24302);
   U14125 : NAND3_X1 port map( A1 => n9429, A2 => n9984, A3 => n9982, ZN => 
                           n471);
   U14397 : NAND2_X1 port map( A1 => n10427, A2 => n3100, ZN => n10430);
   U14481 : NAND2_X1 port map( A1 => n1180, A2 => n10243, ZN => n10427);
   U14583 : NAND2_X1 port map( A1 => n1859, A2 => n1860, ZN => n12639);
   U14584 : NAND3_X1 port map( A1 => n794, A2 => n10055, A3 => n10056, ZN => 
                           n11062);
   U14637 : NAND2_X1 port map( A1 => n1122, A2 => n25441, ZN => n987);
   U14660 : OAI211_X1 port map( C1 => n9927, C2 => n9346, A => n24304, B => 
                           n9604, ZN => n4730);
   U14672 : NAND2_X1 port map( A1 => n9927, A2 => n24084, ZN => n24304);
   U14692 : NAND2_X1 port map( A1 => n20388, A2 => n19345, ZN => n3165);
   U14717 : XOR2_X1 port map( A => n18098, B => n18351, Z => n18208);
   U14718 : AOI21_X1 port map( B1 => n24317, B2 => n22950, A => n22949, ZN => 
                           n24343);
   U14793 : OR2_X1 port map( A1 => n11114, A2 => n11112, ZN => n9343);
   U14807 : OR2_X1 port map( A1 => n24911, A2 => n22744, ZN => n2199);
   U14899 : AOI21_X1 port map( B1 => n20370, B2 => n19574, A => n2016, ZN => 
                           n21205);
   U15014 : NAND3_X1 port map( A1 => n3483, A2 => n3481, A3 => n3477, ZN => 
                           n24306);
   U15070 : XOR2_X1 port map( A => n21477, B => n21222, Z => n21970);
   U15071 : XNOR2_X1 port map( A => n21973, B => n21972, ZN => n22835);
   U15079 : CLKBUF_X1 port map( A => n23342, Z => n24400);
   U15081 : CLKBUF_X1 port map( A => n22395, Z => n24321);
   U15098 : XNOR2_X2 port map( A => n19870, B => n19869, ZN => n22231);
   U15131 : OAI21_X1 port map( B1 => n16531, B2 => n16530, A => n16529, ZN => 
                           n18420);
   U15182 : INV_X1 port map( A => n23332, ZN => n24309);
   U15204 : XOR2_X1 port map( A => n18418, B => n18420, Z => n18421);
   U15206 : INV_X1 port map( A => n4139, ZN => n24310);
   U15289 : INV_X1 port map( A => n4139, ZN => n19235);
   U15327 : XNOR2_X1 port map( A => n20746, B => n20745, ZN => n24311);
   U15328 : XNOR2_X1 port map( A => n18020, B => n18019, ZN => n24312);
   U15366 : AOI21_X1 port map( B1 => n22910, B2 => n22909, A => n22908, ZN => 
                           n24313);
   U15405 : XNOR2_X1 port map( A => n18019, B => n18020, ZN => n19359);
   U15458 : AOI21_X1 port map( B1 => n22910, B2 => n22909, A => n22908, ZN => 
                           n23529);
   U15580 : OR2_X1 port map( A1 => n18941, A2 => n18940, ZN => n24315);
   U15708 : OAI21_X1 port map( B1 => n21882, B2 => n21881, A => n21880, ZN => 
                           n24316);
   U15716 : XOR2_X1 port map( A => n8183, B => n8713, Z => n8186);
   U15786 : OR2_X1 port map( A1 => n22279, A2 => n22280, ZN => n24317);
   U15944 : XNOR2_X1 port map( A => n20603, B => n20604, ZN => n5378);
   U15950 : XNOR2_X1 port map( A => n8290, B => n8289, ZN => n9806);
   U16005 : OAI21_X1 port map( B1 => n25374, B2 => n18770, A => n18769, ZN => 
                           n20277);
   U16015 : XOR2_X1 port map( A => n17957, B => n17956, Z => n24318);
   U16212 : OR2_X1 port map( A1 => n19673, A2 => n19672, ZN => n24319);
   U16256 : CLKBUF_X1 port map( A => n23612, Z => n24320);
   U16275 : MUX2_X1 port map( A => n19985, B => n19986, S => n2098, Z => n19990
                           );
   U16286 : INV_X1 port map( A => n3198, ZN => n20194);
   U16397 : AND2_X1 port map( A1 => n2674, A2 => n22946, ZN => n24322);
   U16670 : XOR2_X1 port map( A => n8622, B => n8058, Z => n7042);
   U16729 : AND2_X1 port map( A1 => n5678, A2 => n3219, ZN => n24323);
   U16730 : XNOR2_X1 port map( A => n16502, B => n16503, ZN => n24324);
   U16763 : XNOR2_X1 port map( A => n16502, B => n16503, ZN => n19128);
   U16837 : AOI21_X1 port map( B1 => n15725, B2 => n16457, A => n16456, ZN => 
                           n16849);
   U16846 : XNOR2_X1 port map( A => n4810, B => n18505, ZN => n24326);
   U16882 : NAND3_X1 port map( A1 => n5501, A2 => n1458, A3 => n4363, ZN => 
                           n24327);
   U17046 : XNOR2_X1 port map( A => n18505, B => n4810, ZN => n19397);
   U17143 : XOR2_X1 port map( A => n12364, B => n12089, Z => n24328);
   U17212 : XNOR2_X1 port map( A => n17376, B => n17377, ZN => n24329);
   U17215 : XNOR2_X1 port map( A => n17376, B => n17377, ZN => n19537);
   U17225 : OAI211_X1 port map( C1 => n16196, C2 => n15901, A => n5408, B => 
                           n5407, ZN => n17421);
   U17230 : BUF_X2 port map( A => n18596, Z => n19177);
   U17235 : XNOR2_X1 port map( A => n8993, B => n8992, ZN => n24332);
   U17237 : NOR2_X1 port map( A1 => n22431, A2 => n22432, ZN => n24515);
   U17306 : BUF_X1 port map( A => n22205, Z => n24333);
   U17312 : XNOR2_X1 port map( A => n20908, B => n5503, ZN => n22205);
   U17332 : NOR2_X2 port map( A1 => n23514, A2 => n23517, ZN => n23527);
   U17344 : XNOR2_X1 port map( A => n17975, B => n5326, ZN => n24335);
   U17492 : XNOR2_X1 port map( A => n17975, B => n5326, ZN => n19092);
   U17530 : XNOR2_X1 port map( A => n18403, B => n18402, ZN => n18788);
   U17555 : OR2_X1 port map( A1 => n17886, A2 => n19471, ZN => n3749);
   U17612 : AOI21_X1 port map( B1 => n16695, B2 => n16694, A => n16693, ZN => 
                           n24337);
   U17615 : AOI21_X1 port map( B1 => n16695, B2 => n16694, A => n16693, ZN => 
                           n17664);
   U17706 : NOR2_X1 port map( A1 => n24933, A2 => n23394, ZN => n24339);
   U17956 : NAND2_X1 port map( A1 => n3863, A2 => n3864, ZN => n24340);
   U18077 : BUF_X1 port map( A => n20904, Z => n20727);
   U18109 : XNOR2_X1 port map( A => n21419, B => n21418, ZN => n24341);
   U18110 : XNOR2_X1 port map( A => n21419, B => n21418, ZN => n24342);
   U18135 : AOI21_X1 port map( B1 => n24317, B2 => n22950, A => n22949, ZN => 
                           n23354);
   U18347 : OR2_X2 port map( A1 => n4397, A2 => n4398, ZN => n23714);
   U18364 : XNOR2_X1 port map( A => n18572, B => n18571, ZN => n19166);
   U18629 : XNOR2_X1 port map( A => n14493, B => n4875, ZN => n15280);
   U18635 : OAI211_X1 port map( C1 => n12697, C2 => n13278, A => n17, B => 
                           n12696, ZN => n24347);
   U18639 : XNOR2_X1 port map( A => n11972, B => n11973, ZN => n13278);
   U18644 : OAI211_X1 port map( C1 => n12697, C2 => n13278, A => n17, B => 
                           n12696, ZN => n14189);
   U18714 : AOI21_X1 port map( B1 => n22131, B2 => n22968, A => n22130, ZN => 
                           n23263);
   U18776 : OR2_X1 port map( A1 => n24075, A2 => n23064, ZN => n24350);
   U18815 : XOR2_X1 port map( A => n15302, B => n15301, Z => n24352);
   U18962 : OR2_X1 port map( A1 => n19593, A2 => n4479, ZN => n24354);
   U18997 : INV_X2 port map( A => n23640, ZN => n23649);
   U19039 : AND2_X2 port map( A1 => n1007, A2 => n1006, ZN => n23640);
   U19073 : INV_X1 port map( A => n22933, ZN => n24356);
   U19074 : INV_X1 port map( A => n20960, ZN => n24357);
   U19083 : XNOR2_X1 port map( A => n21525, B => n22014, ZN => n21308);
   U19088 : AND2_X1 port map( A1 => n22853, A2 => n5421, ZN => n602);
   U19089 : INV_X1 port map( A => n23265, ZN => n24360);
   U19175 : XNOR2_X1 port map( A => n19624, B => n19623, ZN => n24362);
   U19189 : XNOR2_X1 port map( A => n19624, B => n19623, ZN => n21825);
   U19219 : BUF_X1 port map( A => n20102, Z => n24370);
   U19306 : XOR2_X1 port map( A => n21733, B => n21732, Z => n24364);
   U19341 : XNOR2_X1 port map( A => n1103, B => n1102, ZN => n24366);
   U19342 : XNOR2_X1 port map( A => n1103, B => n1102, ZN => n16004);
   U19373 : XNOR2_X1 port map( A => n20796, B => n21683, ZN => n1363);
   U19390 : OR2_X1 port map( A1 => n12529, A2 => n12528, ZN => n24368);
   U19406 : XNOR2_X1 port map( A => n20850, B => n20849, ZN => n24369);
   U19445 : XNOR2_X1 port map( A => n20850, B => n20849, ZN => n23574);
   U19575 : OAI21_X2 port map( B1 => n21657, B2 => n21656, A => n21655, ZN => 
                           n23374);
   U19707 : BUF_X1 port map( A => n18291, Z => n24371);
   U19726 : INV_X1 port map( A => n23592, ZN => n24372);
   U19728 : XNOR2_X1 port map( A => n10421, B => n10420, ZN => n24373);
   U19907 : XNOR2_X1 port map( A => n10421, B => n10420, ZN => n13169);
   U19950 : BUF_X1 port map( A => n23727, Z => n24374);
   U19986 : INV_X1 port map( A => n12510, ZN => n13185);
   U20069 : NAND3_X1 port map( A1 => n13106, A2 => n13105, A3 => n13104, ZN => 
                           n14100);
   U20169 : NAND2_X1 port map( A1 => n22269, A2 => n2833, ZN => n23251);
   U20194 : NAND3_X1 port map( A1 => n5099, A2 => n3749, A3 => n3747, ZN => 
                           n24378);
   U20244 : XNOR2_X2 port map( A => n21667, B => n21666, ZN => n22842);
   U20288 : XNOR2_X1 port map( A => n21002, B => n21001, ZN => n24379);
   U20293 : NOR2_X1 port map( A1 => n23514, A2 => n23517, ZN => n24380);
   U20442 : INV_X1 port map( A => n23697, ZN => n24381);
   U20607 : INV_X1 port map( A => n23697, ZN => n23721);
   U20683 : NAND3_X1 port map( A1 => n2789, A2 => n2790, A3 => n16259, ZN => 
                           n24384);
   U20687 : NAND2_X1 port map( A1 => n15633, A2 => n3592, ZN => n24385);
   U20785 : XNOR2_X1 port map( A => n16738, B => n16737, ZN => n24386);
   U20795 : XNOR2_X1 port map( A => n14796, B => n14795, ZN => n24387);
   U20811 : XNOR2_X1 port map( A => n14796, B => n14795, ZN => n2607);
   U20922 : NOR2_X1 port map( A1 => n23579, A2 => n23578, ZN => n24389);
   U21000 : NOR2_X1 port map( A1 => n23579, A2 => n23578, ZN => n24390);
   U21023 : INV_X1 port map( A => n2306, ZN => n10685);
   U21024 : OR2_X1 port map( A1 => n16256, A2 => n16255, ZN => n24391);
   U21025 : NAND2_X1 port map( A1 => n4434, A2 => n23001, ZN => n24392);
   U21026 : XNOR2_X1 port map( A => n17493, B => n17492, ZN => n24393);
   U21060 : OAI21_X1 port map( B1 => n22327, B2 => n22326, A => n3682, ZN => 
                           n24394);
   U21061 : XNOR2_X1 port map( A => n17493, B => n17492, ZN => n19270);
   U21068 : OAI21_X1 port map( B1 => n22327, B2 => n22326, A => n3682, ZN => 
                           n23177);
   U21096 : INV_X1 port map( A => n1147, ZN => n24395);
   U21152 : NOR2_X1 port map( A1 => n21761, A2 => n23573, ZN => n24397);
   U21204 : NOR2_X1 port map( A1 => n21761, A2 => n23573, ZN => n23566);
   U21237 : INV_X1 port map( A => n24386, ZN => n24399);
   U21261 : OAI211_X1 port map( C1 => n22960, C2 => n22959, A => n4127, B => 
                           n4126, ZN => n23342);
   U21263 : OAI211_X1 port map( C1 => n10958, C2 => n10699, A => n10957, B => 
                           n10956, ZN => n24401);
   U21279 : OAI211_X1 port map( C1 => n10958, C2 => n10699, A => n10957, B => 
                           n10956, ZN => n11957);
   U21303 : AOI22_X1 port map( A1 => n13354, A2 => n13353, B1 => n5588, B2 => 
                           n25430, ZN => n13996);
   U21306 : XOR2_X1 port map( A => n14925, B => n14924, Z => n24403);
   U21344 : NOR2_X1 port map( A1 => n21710, A2 => n695, ZN => n24404);
   U21372 : NOR2_X1 port map( A1 => n21710, A2 => n695, ZN => n22987);
   U21413 : XNOR2_X1 port map( A => Key(44), B => Plaintext(44), ZN => n24405);
   U21541 : XNOR2_X1 port map( A => n18411, B => n18410, ZN => n24407);
   U21578 : AND2_X2 port map( A1 => n24408, A2 => n24409, ZN => n23064);
   U21580 : NOR2_X1 port map( A1 => n21150, A2 => n570, ZN => n24408);
   U21608 : OR2_X1 port map( A1 => n21932, A2 => n22465, ZN => n24409);
   U21624 : XNOR2_X1 port map( A => n18411, B => n18410, ZN => n19395);
   U21643 : NAND2_X1 port map( A1 => n15835, A2 => n15836, ZN => n24410);
   U21644 : XNOR2_X1 port map( A => n21475, B => n21474, ZN => n24411);
   U21658 : OAI21_X1 port map( B1 => n21490, B2 => n21489, A => n21488, ZN => 
                           n24412);
   U21743 : XNOR2_X1 port map( A => n21475, B => n21474, ZN => n22967);
   U21769 : OAI21_X1 port map( B1 => n21490, B2 => n21489, A => n21488, ZN => 
                           n23369);
   U21848 : XNOR2_X1 port map( A => n20635, B => n20634, ZN => n24415);
   U21986 : XNOR2_X1 port map( A => n20635, B => n20634, ZN => n22335);
   U22203 : BUF_X1 port map( A => n18301, Z => n24416);
   U22228 : OAI211_X1 port map( C1 => n16590, C2 => n17076, A => n2374, B => 
                           n2373, ZN => n18301);
   U22289 : OAI21_X1 port map( B1 => n13404, B2 => n13403, A => n13402, ZN => 
                           n24418);
   U22445 : OAI21_X1 port map( B1 => n13404, B2 => n13403, A => n13402, ZN => 
                           n14591);
   U22463 : CLKBUF_X1 port map( A => n11005, Z => n24420);
   U22698 : XNOR2_X1 port map( A => n16570, B => n16571, ZN => n24421);
   U22720 : XNOR2_X1 port map( A => n16571, B => n16570, ZN => n19556);
   U22727 : INV_X1 port map( A => n13328, ZN => n24422);
   U22757 : NAND2_X1 port map( A1 => n13891, A2 => n1819, ZN => n24423);
   U22758 : XNOR2_X1 port map( A => n17800, B => n17799, ZN => n24424);
   U22896 : XNOR2_X1 port map( A => n17800, B => n17799, ZN => n19366);
   U22930 : AOI21_X1 port map( B1 => n22841, B2 => n22840, A => n22839, ZN => 
                           n23398);
   U22962 : XOR2_X1 port map( A => n17549, B => n17548, Z => n24427);
   U22965 : INV_X1 port map( A => n23843, ZN => n24428);
   U23005 : XNOR2_X1 port map( A => n14624, B => n14623, ZN => n24429);
   U23008 : XNOR2_X1 port map( A => n14624, B => n14623, ZN => n24430);
   U23163 : BUF_X1 port map( A => n17919, Z => n24431);
   U23290 : AOI22_X1 port map( A1 => n3306, A2 => n16546, B1 => n723, B2 => 
                           n283, ZN => n17919);
   U23368 : OAI211_X1 port map( C1 => n17275, C2 => n16690, A => n16689, B => 
                           n16688, ZN => n24433);
   U23393 : OAI211_X1 port map( C1 => n17275, C2 => n16690, A => n16689, B => 
                           n16688, ZN => n17913);
   U23405 : NAND2_X1 port map( A1 => n20912, A2 => n815, ZN => n24434);
   U23406 : NOR2_X1 port map( A1 => n23462, A2 => n22733, ZN => n24435);
   U23430 : AOI21_X2 port map( B1 => n6633, B2 => n6632, A => n6631, ZN => 
                           n7788);
   U23433 : OR2_X1 port map( A1 => n16483, A2 => n25238, ZN => n757);
   U23451 : XNOR2_X1 port map( A => n21100, B => n21099, ZN => n24439);
   U23463 : MUX2_X1 port map( A => n22777, B => n22776, S => n22677, Z => 
                           n24440);
   U23465 : XNOR2_X1 port map( A => n21099, B => n21100, ZN => n23999);
   U23717 : XNOR2_X1 port map( A => n15555, B => n15554, ZN => n24441);
   U23760 : XNOR2_X1 port map( A => n15555, B => n15554, ZN => n19302);
   U23772 : INV_X1 port map( A => n2710, ZN => n24442);
   U23807 : OAI21_X1 port map( B1 => n16395, B2 => n16394, A => n16396, ZN => 
                           n24444);
   U23808 : OAI21_X1 port map( B1 => n16395, B2 => n16394, A => n16396, ZN => 
                           n17438);
   U23979 : OAI21_X1 port map( B1 => n7936, B2 => n7935, A => n7934, ZN => 
                           n24445);
   U23981 : XNOR2_X1 port map( A => n9056, B => n9055, ZN => n24446);
   U23989 : OAI21_X1 port map( B1 => n7936, B2 => n7935, A => n7934, ZN => 
                           n9195);
   U24074 : OAI211_X1 port map( C1 => n22787, C2 => n24406, A => n22786, B => 
                           n22785, ZN => n24448);
   U24075 : OAI211_X1 port map( C1 => n22787, C2 => n24406, A => n22786, B => 
                           n22785, ZN => n24010);
   U24076 : BUF_X1 port map( A => n23391, Z => n24449);
   U24077 : OAI211_X1 port map( C1 => n22030, C2 => n22029, A => n5771, B => 
                           n22028, ZN => n23391);
   U24080 : XNOR2_X1 port map( A => n17724, B => n17725, ZN => n24451);
   U24081 : XOR2_X1 port map( A => n17964, B => n17965, Z => n24452);
   U24082 : XNOR2_X1 port map( A => n22006, B => n21444, ZN => n24453);
   U24084 : OAI21_X1 port map( B1 => n19538, B2 => n24329, A => n19536, ZN => 
                           n24454);
   U24085 : XNOR2_X1 port map( A => n17530, B => n17531, ZN => n24457);
   U24086 : XNOR2_X1 port map( A => n15108, B => n15107, ZN => n16356);
   U24087 : XNOR2_X1 port map( A => n14371, B => n14372, ZN => n24458);
   U24088 : XNOR2_X1 port map( A => n14371, B => n14372, ZN => n24459);
   U24089 : OAI211_X1 port map( C1 => n24926, C2 => n24582, A => n19356, B => 
                           n19355, ZN => n24460);
   U24090 : OAI211_X1 port map( C1 => n24926, C2 => n24582, A => n19356, B => 
                           n19355, ZN => n24461);
   U24091 : OAI211_X1 port map( C1 => n24926, C2 => n24582, A => n19356, B => 
                           n19355, ZN => n20394);
   U24092 : CLKBUF_X1 port map( A => n13488, Z => n24462);
   U24093 : INV_X1 port map( A => n20597, ZN => n24463);
   U24094 : XNOR2_X1 port map( A => n14620, B => n14721, ZN => n15170);
   U24095 : NOR2_X1 port map( A1 => n156, A2 => n18946, ZN => n24464);
   U24096 : NOR2_X1 port map( A1 => n156, A2 => n18946, ZN => n19983);
   U24097 : NAND4_X1 port map( A1 => n22024, A2 => n22022, A3 => n22023, A4 => 
                           n22025, ZN => n24465);
   U24098 : NAND4_X1 port map( A1 => n22024, A2 => n22022, A3 => n22023, A4 => 
                           n22025, ZN => n23393);
   U24099 : XOR2_X1 port map( A => Key(6), B => Plaintext(6), Z => n24466);
   U24100 : XNOR2_X1 port map( A => n12619, B => n12620, ZN => n24467);
   U24101 : XNOR2_X1 port map( A => n12619, B => n12620, ZN => n16352);
   U24102 : XNOR2_X1 port map( A => n19161, B => n19160, ZN => n24468);
   U24103 : NOR2_X1 port map( A1 => n19626, A2 => n19625, ZN => n23858);
   U24104 : NOR2_X1 port map( A1 => n2730, A2 => n8225, ZN => n24470);
   U24105 : OAI21_X1 port map( B1 => n15976, B2 => n15975, A => n15974, ZN => 
                           n24471);
   U24107 : OAI21_X1 port map( B1 => n15976, B2 => n15975, A => n15974, ZN => 
                           n17573);
   U24108 : OR2_X1 port map( A1 => n4846, A2 => n16357, ZN => n18);
   U24109 : MUX2_X2 port map( A => n22136, B => n22135, S => n22401, Z => 
                           n23281);
   U24110 : NOR2_X1 port map( A1 => n19673, A2 => n19672, ZN => n24472);
   U24112 : NOR2_X1 port map( A1 => n19673, A2 => n19672, ZN => n21649);
   U24113 : OAI21_X1 port map( B1 => n21374, B2 => n21373, A => n21372, ZN => 
                           n23153);
   U24114 : OAI21_X1 port map( B1 => n6880, B2 => n6879, A => n1888, ZN => 
                           n24474);
   U24115 : OAI21_X1 port map( B1 => n6880, B2 => n6879, A => n1888, ZN => 
                           n24475);
   U24116 : OAI21_X1 port map( B1 => n6880, B2 => n6879, A => n1888, ZN => 
                           n7948);
   U24117 : INV_X1 port map( A => n24931, ZN => n24477);
   U24118 : XNOR2_X1 port map( A => n17761, B => n17760, ZN => n19386);
   U24119 : OAI211_X1 port map( C1 => n2079, C2 => n9687, A => n9685, B => 
                           n9686, ZN => n24479);
   U24120 : OAI211_X1 port map( C1 => n2079, C2 => n9687, A => n9685, B => 
                           n9686, ZN => n24480);
   U24121 : INV_X1 port map( A => n19581, ZN => n24481);
   U24122 : OAI211_X1 port map( C1 => n2079, C2 => n9687, A => n9685, B => 
                           n9686, ZN => n11152);
   U24123 : XNOR2_X1 port map( A => n15222, B => n15221, ZN => n24482);
   U24124 : XNOR2_X1 port map( A => n18072, B => n18071, ZN => n24483);
   U24125 : XNOR2_X1 port map( A => n18072, B => n18071, ZN => n19590);
   U24126 : OR2_X1 port map( A1 => n22222, A2 => n24484, ZN => n1237);
   U24127 : OR2_X1 port map( A1 => n22220, A2 => n22219, ZN => n24484);
   U24129 : OAI21_X1 port map( B1 => n20323, B2 => n20322, A => n20321, ZN => 
                           n20882);
   U24130 : OAI211_X1 port map( C1 => n16709, C2 => n16708, A => n16707, B => 
                           n2057, ZN => n24488);
   U24132 : OAI211_X1 port map( C1 => n16709, C2 => n16708, A => n16707, B => 
                           n2057, ZN => n18678);
   U24133 : XNOR2_X1 port map( A => n11731, B => n11730, ZN => n24490);
   U24134 : XNOR2_X1 port map( A => n11731, B => n11730, ZN => n13221);
   U24135 : OAI211_X1 port map( C1 => n20564, C2 => n25221, A => n4009, B => 
                           n19734, ZN => n21455);
   U24136 : NAND2_X1 port map( A1 => n24493, A2 => n24494, ZN => n23357);
   U24137 : OR3_X1 port map( A1 => n22961, A2 => n24492, A3 => n23359, ZN => 
                           n24493);
   U24138 : OR3_X1 port map( A1 => n23361, A2 => n23350, A3 => n23349, ZN => 
                           n24494);
   U24139 : XNOR2_X1 port map( A => n15227, B => n15228, ZN => n16191);
   U24144 : XOR2_X1 port map( A => n10300, B => n10299, Z => n24499);
   U24145 : XNOR2_X1 port map( A => n5780, B => Key(95), ZN => n24500);
   U24146 : XNOR2_X1 port map( A => n5780, B => Key(95), ZN => n24501);
   U24147 : OAI211_X1 port map( C1 => n14012, C2 => n14011, A => n856, B => 
                           n855, ZN => n24502);
   U24148 : XNOR2_X1 port map( A => n5780, B => Key(95), ZN => n6715);
   U24149 : OAI211_X1 port map( C1 => n14012, C2 => n14011, A => n856, B => 
                           n855, ZN => n15138);
   U24153 : XNOR2_X1 port map( A => n8547, B => n8546, ZN => n24505);
   U24154 : XNOR2_X1 port map( A => n15014, B => n15013, ZN => n24506);
   U24155 : XNOR2_X1 port map( A => n8547, B => n8546, ZN => n9781);
   U24156 : OAI211_X1 port map( C1 => n13711, C2 => n13394, A => n11681, B => 
                           n11680, ZN => n15401);
   U24158 : BUF_X1 port map( A => n15229, Z => n24508);
   U24159 : AOI22_X2 port map( A1 => n4601, A2 => n3727, B1 => n19017, B2 => 
                           n19393, ZN => n20445);
   U24160 : XNOR2_X1 port map( A => Key(156), B => Plaintext(156), ZN => n24509
                           );
   U24161 : XNOR2_X1 port map( A => n11231, B => n11230, ZN => n24512);
   U24162 : XNOR2_X1 port map( A => n11231, B => n11230, ZN => n24513);
   U24163 : XNOR2_X1 port map( A => n8027, B => n8028, ZN => n9450);
   U24164 : AND4_X1 port map( A1 => n10442, A2 => n2766, A3 => n10440, A4 => 
                           n10441, ZN => n24514);
   U24165 : NOR2_X1 port map( A1 => n22431, A2 => n22432, ZN => n23371);
   U24166 : XNOR2_X2 port map( A => n10449, B => n10450, ZN => n4766);
   U24168 : XNOR2_X1 port map( A => n17222, B => n17221, ZN => n24516);
   U24170 : NOR2_X1 port map( A1 => n22802, A2 => n22659, ZN => n24517);
   U24171 : AND2_X1 port map( A1 => n2978, A2 => n22664, ZN => n24518);
   U24172 : NAND2_X1 port map( A1 => n23363, A2 => n23362, ZN => n23364);
   U24173 : NAND2_X1 port map( A1 => n1802, A2 => n1803, ZN => n22839);
   U24174 : NAND3_X1 port map( A1 => n24520, A2 => n13434, A3 => n24519, ZN => 
                           n14654);
   U24175 : NAND2_X1 port map( A1 => n13432, A2 => n14106, ZN => n24520);
   U24176 : NAND2_X1 port map( A1 => n24521, A2 => n10486, ZN => n9608);
   U24178 : NAND2_X1 port map( A1 => n12687, A2 => n24522, ZN => n13322);
   U24179 : NAND2_X1 port map( A1 => n12945, A2 => n12942, ZN => n24522);
   U24182 : NAND2_X1 port map( A1 => n281, A2 => n17012, ZN => n17357);
   U24183 : OR2_X1 port map( A1 => n6369, A2 => n6071, ZN => n7003);
   U24184 : NAND3_X1 port map( A1 => n5389, A2 => n5390, A3 => n7628, ZN => 
                           n5388);
   U24185 : NAND2_X1 port map( A1 => n11101, A2 => n10914, ZN => n11031);
   U24186 : NAND3_X1 port map( A1 => n5312, A2 => n5311, A3 => n5313, ZN => 
                           n5310);
   U24187 : AOI22_X1 port map( A1 => n6200, A2 => n6909, B1 => n6201, B2 => 
                           n6774, ZN => n2784);
   U24190 : NAND2_X1 port map( A1 => n6436, A2 => n25325, ZN => n24525);
   U24191 : NAND2_X1 port map( A1 => n620, A2 => n4844, ZN => n619);
   U24192 : AND2_X1 port map( A1 => n10630, A2 => n10789, ZN => n24526);
   U24193 : OR2_X1 port map( A1 => n12807, A2 => n12808, ZN => n24527);
   U24195 : OR2_X1 port map( A1 => n16128, A2 => n16154, ZN => n24528);
   U24196 : BUF_X1 port map( A => n17463, Z => n288);
   U24198 : AND2_X1 port map( A1 => n17016, A2 => n17212, ZN => n24529);
   U24199 : INV_X1 port map( A => n19357, ZN => n19037);
   U24201 : NAND3_X1 port map( A1 => n4017, A2 => n20567, A3 => n20562, ZN => 
                           n24530);
   U24202 : NOR2_X1 port map( A1 => n3428, A2 => n349, ZN => n24531);
   U8837 : XNOR2_X2 port map( A => n3506, B => n8104, ZN => n9899);
   U2447 : OAI21_X2 port map( B1 => n10157, B2 => n9854, A => n9350, ZN => 
                           n1499);
   U658 : NAND2_X2 port map( A1 => n6185, A2 => n6186, ZN => n7647);
   U1944 : AND3_X2 port map( A1 => n7117, A2 => n5689, A3 => n5691, ZN => n8616
                           );
   U2159 : XNOR2_X2 port map( A => n15372, B => n15373, ZN => n16060);
   U3222 : BUF_X2 port map( A => n19155, Z => n21038);
   U1152 : AOI21_X2 port map( B1 => n22512, B2 => n25496, A => n22511, ZN => 
                           n23181);
   U2369 : NAND4_X2 port map( A1 => n10864, A2 => n10866, A3 => n10865, A4 => 
                           n10863, ZN => n12096);
   U8717 : OR2_X2 port map( A1 => n9546, A2 => n9545, ZN => n10445);
   U1330 : XNOR2_X2 port map( A => n12014, B => n12015, ZN => n13264);
   U2047 : BUF_X1 port map( A => n16849, Z => n16985);
   U1841 : AND2_X2 port map( A1 => n5473, A2 => n5476, ZN => n20255);
   U7009 : NAND3_X2 port map( A1 => n5750, A2 => n1930, A3 => n1395, ZN => 
                           n14919);
   U15937 : BUF_X2 port map( A => n11411, Z => n13909);
   U12115 : XNOR2_X2 port map( A => Key(77), B => Plaintext(77), ZN => n6051);
   U6823 : AOI21_X2 port map( B1 => n9720, B2 => n9719, A => n204, ZN => n11967
                           );
   U3690 : AND2_X2 port map( A1 => n893, A2 => n1572, ZN => n13785);
   U80 : NAND4_X2 port map( A1 => n10797, A2 => n10796, A3 => n10795, A4 => 
                           n10794, ZN => n12401);
   U1447 : AOI22_X2 port map( A1 => n15690, A2 => n16472, B1 => n15688, B2 => 
                           n15689, ZN => n16551);
   U1521 : XNOR2_X2 port map( A => n8101, B => n8100, ZN => n2294);
   U224 : BUF_X1 port map( A => n10135, Z => n24025);
   U14020 : BUF_X2 port map( A => n9348, Z => n10162);
   U1056 : NOR2_X2 port map( A1 => n15872, A2 => n15871, ZN => n17084);
   U144 : INV_X2 port map( A => n16121, ZN => n16122);
   U2151 : BUF_X1 port map( A => n5992, Z => n6824);
   U192 : AND3_X2 port map( A1 => n2124, A2 => n3770, A3 => n3768, ZN => n2602)
                           ;
   U1684 : MUX2_X2 port map( A => n22605, B => n22604, S => n22603, Z => n23050
                           );
   U820 : BUF_X1 port map( A => n23119, Z => n24059);
   U7560 : AND2_X2 port map( A1 => n4888, A2 => n17358, ZN => n18123);
   U807 : NAND4_X2 port map( A1 => n5602, A2 => n5601, A3 => n7737, A4 => n5600
                           , ZN => n8690);
   U200 : INV_X1 port map( A => n10861, ZN => n10190);
   U2472 : NOR2_X1 port map( A1 => n307, A2 => n9692, ZN => n9880);
   U4749 : NAND2_X2 port map( A1 => n20380, A2 => n24127, ZN => n21633);
   U2297 : BUF_X1 port map( A => n12433, Z => n13137);
   U16266 : BUF_X2 port map( A => n11805, Z => n13968);
   U9360 : NAND2_X2 port map( A1 => n16190, A2 => n3222, ZN => n17185);
   U1423 : OAI211_X2 port map( C1 => n16675, C2 => n16876, A => n16674, B => 
                           n16673, ZN => n18674);
   U336 : NAND2_X2 port map( A1 => n2897, A2 => n2896, ZN => n8699);
   U988 : AND2_X2 port map( A1 => n15918, A2 => n15919, ZN => n17364);
   U1918 : BUF_X1 port map( A => n18749, Z => n19138);
   U416 : OAI21_X2 port map( B1 => n9262, B2 => n9858, A => n9261, ZN => n10737
                           );
   U2208 : NAND4_X2 port map( A1 => n870, A2 => n14248, A3 => n14247, A4 => 
                           n14246, ZN => n14907);
   U1929 : INV_X2 port map( A => n4667, ZN => n19476);
   U1503 : OAI211_X2 port map( C1 => n3575, C2 => n10905, A => n4343, B => 
                           n3574, ZN => n12159);
   U17911 : XNOR2_X2 port map( A => n14540, B => n14539, ZN => n16391);
   U14876 : AOI21_X2 port map( B1 => n20370, B2 => n19574, A => n2016, ZN => 
                           n24305);
   U2163 : XNOR2_X1 port map( A => n14991, B => n14990, ZN => n16022);
   U2512 : BUF_X2 port map( A => n9495, Z => n10090);
   U5891 : INV_X1 port map( A => n19494, ZN => n20235);
   U403 : OR2_X2 port map( A1 => n15754, A2 => n15753, ZN => n16902);
   U15697 : XNOR2_X2 port map( A => n11182, B => n11183, ZN => n12455);
   U1864 : BUF_X2 port map( A => n19851, Z => n19660);
   U19440 : AOI22_X2 port map( A1 => n16919, A2 => n16918, B1 => n16917, B2 => 
                           n16916, ZN => n17582);
   U12025 : AND2_X1 port map( A1 => n25197, A2 => n14335, ZN => n14344);
   U6931 : NAND3_X2 port map( A1 => n7343, A2 => n7344, A3 => n1999, ZN => 
                           n8964);
   U3491 : XNOR2_X1 port map( A => n15256, B => n15257, ZN => n2610);
   U10956 : NAND3_X2 port map( A1 => n4156, A2 => n10621, A3 => n3724, ZN => 
                           n11424);
   U2927 : XNOR2_X1 port map( A => n15108, B => n15107, ZN => n24456);
   U1987 : AND2_X2 port map( A1 => n567, A2 => n566, ZN => n18334);
   U13340 : OAI211_X2 port map( C1 => n7445, C2 => n7375, A => n7374, B => 
                           n7373, ZN => n9182);
   U1420 : AND2_X2 port map( A1 => n3784, A2 => n2641, ZN => n18128);
   U19856 : INV_X1 port map( A => n17653, ZN => n18601);
   U1787 : XNOR2_X2 port map( A => n20967, B => n20968, ZN => n22918);
   U22755 : NOR2_X1 port map( A1 => n25239, A2 => n23890, ZN => n23909);
   U19259 : INV_X1 port map( A => n16660, ZN => n17198);
   U18758 : OAI21_X1 port map( B1 => n15709, B2 => n15708, A => n2636, ZN => 
                           n15713);
   U12417 : XNOR2_X1 port map( A => Key(178), B => Plaintext(178), ZN => n6467)
                           ;
   U12357 : XNOR2_X1 port map( A => Key(188), B => Plaintext(188), ZN => n6452)
                           ;
   U12478 : XNOR2_X1 port map( A => Key(97), B => Plaintext(97), ZN => n6588);
   U1656 : CLKBUF_X1 port map( A => Key(3), Z => n21169);
   U2735 : XNOR2_X1 port map( A => Key(20), B => Plaintext(20), ZN => n6165);
   U1210 : CLKBUF_X1 port map( A => Key(117), Z => n1870);
   U348 : CLKBUF_X1 port map( A => Key(89), Z => n3093);
   U12472 : XNOR2_X1 port map( A => Key(115), B => Plaintext(115), ZN => n7021)
                           ;
   U4341 : XNOR2_X1 port map( A => Key(100), B => Plaintext(100), ZN => n7035);
   U1352 : CLKBUF_X1 port map( A => Key(14), Z => n21335);
   U1601 : CLKBUF_X1 port map( A => Key(161), Z => n2031);
   U2739 : XNOR2_X1 port map( A => Key(139), B => Plaintext(139), ZN => n6794);
   U12168 : XNOR2_X1 port map( A => Key(78), B => Plaintext(78), ZN => n6396);
   U1208 : CLKBUF_X1 port map( A => Key(100), Z => n16);
   U1566 : CLKBUF_X1 port map( A => Key(142), Z => n2040);
   U1583 : CLKBUF_X1 port map( A => Key(15), Z => n21742);
   U2755 : CLKBUF_X1 port map( A => Key(116), Z => n23983);
   U12146 : XNOR2_X1 port map( A => Key(62), B => Plaintext(62), ZN => n6969);
   U2724 : CLKBUF_X1 port map( A => Key(63), Z => n1896);
   U1664 : CLKBUF_X1 port map( A => Key(37), Z => n641);
   U1203 : CLKBUF_X1 port map( A => Key(137), Z => n21703);
   U1581 : CLKBUF_X1 port map( A => Key(158), Z => n23699);
   U12210 : XNOR2_X1 port map( A => Key(140), B => Plaintext(140), ZN => n6076)
                           ;
   U5902 : XNOR2_X1 port map( A => Key(148), B => Plaintext(148), ZN => n6905);
   U1600 : CLKBUF_X1 port map( A => Key(0), Z => n836);
   U1551 : BUF_X1 port map( A => n6081, Z => n6876);
   U12497 : XNOR2_X1 port map( A => n6023, B => Key(17), ZN => n6275);
   U2713 : XNOR2_X1 port map( A => n495, B => Key(65), ZN => n6570);
   U1076 : XNOR2_X1 port map( A => n5993, B => Key(103), ZN => n6827);
   U12364 : XNOR2_X1 port map( A => n5931, B => Key(191), ZN => n6187);
   U16816 : OAI211_X1 port map( C1 => n7002, C2 => n7003, A => n7001, B => 
                           n7000, ZN => n7962);
   U880 : OR2_X1 port map( A1 => n873, A2 => n6361, ZN => n8367);
   U924 : AOI22_X1 port map( A1 => n6902, A2 => n6475, B1 => n6476, B2 => n6905
                           , ZN => n8074);
   U2659 : OR2_X1 port map( A1 => n5922, A2 => n5923, ZN => n7351);
   U109 : AND3_X1 port map( A1 => n2737, A2 => n5086, A3 => n2736, ZN => n1345)
                           ;
   U2631 : OR2_X1 port map( A1 => n6831, A2 => n6830, ZN => n7984);
   U121 : NAND3_X1 port map( A1 => n4682, A2 => n4681, A3 => n6527, ZN => n7211
                           );
   U10292 : NAND3_X1 port map( A1 => n6231, A2 => n4122, A3 => n4121, ZN => 
                           n7642);
   U7185 : NAND3_X1 port map( A1 => n2032, A2 => n6914, A3 => n6913, ZN => 
                           n7942);
   U2652 : OR2_X1 port map( A1 => n6118, A2 => n6117, ZN => n7527);
   U13005 : INV_X1 port map( A => n7829, ZN => n7048);
   U3608 : NAND3_X1 port map( A1 => n6562, A2 => n6563, A3 => n6561, ZN => 
                           n7444);
   U165 : OR2_X1 port map( A1 => n4994, A2 => n436, ZN => n7669);
   U2580 : OR2_X1 port map( A1 => n7279, A2 => n8511, ZN => n7254);
   U4426 : OR2_X1 port map( A1 => n7540, A2 => n432, ZN => n7547);
   U2578 : OR2_X1 port map( A1 => n7845, A2 => n8374, ZN => n9176);
   U2564 : NAND2_X1 port map( A1 => n6863, A2 => n6862, ZN => n9167);
   U213 : NAND2_X1 port map( A1 => n6854, A2 => n6855, ZN => n8687);
   U9413 : OAI21_X1 port map( B1 => n4483, B2 => n3272, A => n3363, ZN => n8238
                           );
   U2563 : OAI21_X1 port map( B1 => n5861, B2 => n5860, A => n5859, ZN => n8666
                           );
   U2550 : AND2_X1 port map( A1 => n569, A2 => n533, ZN => n5344);
   U633 : NAND2_X1 port map( A1 => n1040, A2 => n1037, ZN => n8874);
   U2554 : OR2_X1 port map( A1 => n7712, A2 => n7711, ZN => n8468);
   U2547 : INV_X1 port map( A => n5344, ZN => n9139);
   U4439 : XNOR2_X1 port map( A => n8448, B => n8983, ZN => n9788);
   U1094 : XNOR2_X1 port map( A => n7876, B => n7875, ZN => n9939);
   U14331 : XNOR2_X1 port map( A => n8811, B => n8810, ZN => n10020);
   U2422 : XNOR2_X1 port map( A => n7744, B => n7743, ZN => n9925);
   U2530 : XNOR2_X1 port map( A => n9085, B => n1385, ZN => n4096);
   U1243 : BUF_X1 port map( A => n9859, Z => n239);
   U4583 : XNOR2_X1 port map( A => n7906, B => n7907, ZN => n9449);
   U11973 : CLKBUF_X1 port map( A => n8141, Z => n9961);
   U1044 : BUF_X1 port map( A => n9328, Z => n9774);
   U11116 : XNOR2_X1 port map( A => n8380, B => n8379, ZN => n10094);
   U14663 : INV_X1 port map( A => n9297, ZN => n10093);
   U2504 : MUX2_X1 port map( A => n9858, B => n9280, S => n239, Z => n10516);
   U2506 : NOR2_X1 port map( A1 => n9959, A2 => n9950, ZN => n9392);
   U2451 : OAI211_X1 port map( C1 => n10049, C2 => n10048, A => n4068, B => 
                           n1403, ZN => n11067);
   U10787 : NAND2_X1 port map( A1 => n10516, A2 => n10517, ZN => n10275);
   U4872 : AND2_X1 port map( A1 => n9392, A2 => n9951, ZN => n10256);
   U1097 : AND4_X1 port map( A1 => n9457, A2 => n9566, A3 => n957, A4 => n955, 
                           ZN => n10887);
   U2465 : OR2_X1 port map( A1 => n9298, A2 => n9498, ZN => n2501);
   U189 : NOR2_X1 port map( A1 => n10174, A2 => n10173, ZN => n10398);
   U9075 : MUX2_X1 port map( A => n9701, B => n9240, S => n9700, Z => n11149);
   U91 : NAND3_X1 port map( A1 => n9371, A2 => n9369, A3 => n9370, ZN => n10451
                           );
   U1509 : NAND3_X1 port map( A1 => n4207, A2 => n9508, A3 => n4210, ZN => n939
                           );
   U417 : NAND4_X1 port map( A1 => n10469, A2 => n10468, A3 => n10467, A4 => 
                           n10466, ZN => n11741);
   U8420 : NAND4_X1 port map( A1 => n2766, A2 => n10440, A3 => n10442, A4 => 
                           n10441, ZN => n11908);
   U1501 : OR2_X1 port map( A1 => n10330, A2 => n10329, ZN => n12134);
   U2556 : XNOR2_X1 port map( A => n11246, B => n11245, ZN => n13217);
   U11889 : XNOR2_X1 port map( A => n12254, B => n12253, ZN => n12272);
   U2315 : CLKBUF_X1 port map( A => n12600, Z => n12966);
   U2312 : BUF_X1 port map( A => n11755, Z => n13222);
   U402 : INV_X1 port map( A => n12674, ZN => n4923);
   U530 : AND2_X1 port map( A1 => n11350, A2 => n13213, ZN => n13208);
   U4477 : OR2_X1 port map( A1 => n13306, A2 => n13307, ZN => n13310);
   U2701 : NOR2_X1 port map( A1 => n13093, A2 => n12650, ZN => n13669);
   U645 : NAND3_X1 port map( A1 => n4867, A2 => n5012, A3 => n5010, ZN => 
                           n14112);
   U2284 : AOI22_X1 port map( A1 => n13239, A2 => n13238, B1 => n13237, B2 => 
                           n4493, ZN => n13982);
   U16926 : MUX2_X1 port map( A => n12849, B => n12848, S => n301, Z => n13504)
                           ;
   U2827 : INV_X1 port map( A => n13775, ZN => n14160);
   U2904 : AND3_X1 port map( A1 => n12567, A2 => n12566, A3 => n5747, ZN => 
                           n14076);
   U17122 : MUX2_X1 port map( A => n13287, B => n13286, S => n25191, Z => 
                           n13923);
   U2813 : NAND2_X1 port map( A1 => n13193, A2 => n13192, ZN => n14106);
   U815 : NAND2_X1 port map( A1 => n779, A2 => n12988, ZN => n14222);
   U2246 : AND2_X1 port map( A1 => n622, A2 => n624, ZN => n13895);
   U340 : OR2_X1 port map( A1 => n14126, A2 => n14129, ZN => n13826);
   U674 : NAND3_X1 port map( A1 => n2155, A2 => n985, A3 => n984, ZN => n15298)
                           ;
   U2204 : NAND2_X1 port map( A1 => n14040, A2 => n5058, ZN => n15095);
   U58 : AND3_X1 port map( A1 => n3368, A2 => n3369, A3 => n3367, ZN => n14815)
                           ;
   U337 : NAND2_X1 port map( A1 => n48, A2 => n4598, ZN => n15183);
   U10812 : AND2_X1 port map( A1 => n183, A2 => n185, ZN => n15422);
   U1510 : XNOR2_X1 port map( A => n15505, B => n24097, ZN => n14909);
   U18278 : INV_X1 port map( A => n14977, ZN => n15342);
   U2136 : BUF_X1 port map( A => n14926, Z => n16277);
   U2175 : XNOR2_X1 port map( A => n15308, B => n15307, ZN => n16048);
   U853 : XNOR2_X1 port map( A => n15101, B => n15100, ZN => n16359);
   U141 : BUF_X1 port map( A => n14664, Z => n16077);
   U2144 : BUF_X1 port map( A => n14625, Z => n15789);
   U2135 : XNOR2_X1 port map( A => n3707, B => n14918, ZN => n16030);
   U1154 : BUF_X1 port map( A => n16149, Z => n213);
   U4495 : NOR2_X1 port map( A1 => n16025, A2 => n15773, ZN => n16602);
   U2070 : AND2_X1 port map( A1 => n14974, A2 => n14975, ZN => n17409);
   U1448 : OAI211_X1 port map( C1 => n4091, C2 => n16273, A => n15771, B => 
                           n4090, ZN => n17425);
   U1439 : NOR2_X1 port map( A1 => n13943, A2 => n13942, ZN => n17419);
   U8933 : NAND3_X1 port map( A1 => n3009, A2 => n3008, A3 => n15982, ZN => 
                           n17042);
   U2056 : NAND3_X1 port map( A1 => n4939, A2 => n14666, A3 => n4938, ZN => 
                           n17276);
   U1018 : NAND2_X1 port map( A1 => n16575, A2 => n16576, ZN => n17132);
   U479 : BUF_X1 port map( A => n16561, Z => n17615);
   U21220 : BUF_X1 port map( A => n17061, Z => n24398);
   U5527 : INV_X1 port map( A => n16963, ZN => n1612);
   U73 : AND2_X1 port map( A1 => n5167, A2 => n15936, ZN => n372);
   U913 : AND2_X1 port map( A1 => n17159, A2 => n17157, ZN => n17164);
   U5526 : NOR2_X1 port map( A1 => n1612, A2 => n17438, ZN => n16830);
   U7156 : OAI22_X1 port map( A1 => n16430, A2 => n1612, B1 => n17128, B2 => 
                           n17445, ZN => n18589);
   U2828 : AND2_X1 port map( A1 => n492, A2 => n491, ZN => n18397);
   U482 : NAND3_X1 port map( A1 => n2055, A2 => n5707, A3 => n2054, ZN => 
                           n18466);
   U24079 : NAND2_X1 port map( A1 => n17004, A2 => n2614, ZN => n18695);
   U234 : NAND2_X1 port map( A1 => n16614, A2 => n16613, ZN => n18220);
   U19778 : AOI21_X1 port map( B1 => n17544, B2 => n17543, A => n17542, ZN => 
                           n18472);
   U1996 : AND4_X1 port map( A1 => n2510, A2 => n17281, A3 => n17282, A4 => 
                           n17280, ZN => n17520);
   U19532 : OR2_X1 port map( A1 => n17083, A2 => n17082, ZN => n18483);
   U1976 : XNOR2_X1 port map( A => n2041, B => n18585, ZN => n19420);
   U695 : XNOR2_X1 port map( A => n15735, B => n15736, ZN => n19307);
   U1971 : XNOR2_X1 port map( A => n18316, B => n18315, ZN => n19565);
   U9356 : XNOR2_X1 port map( A => n16092, B => n16093, ZN => n19304);
   U1965 : XNOR2_X1 port map( A => n18224, B => n18223, ZN => n19185);
   U11239 : INV_X1 port map( A => n19365, ZN => n19371);
   U35 : CLKBUF_X1 port map( A => n18830, Z => n19602);
   U23995 : BUF_X1 port map( A => n2540, Z => n24447);
   U4319 : AOI22_X1 port map( A1 => n19206, A2 => n19379, B1 => n19205, B2 => 
                           n19204, ZN => n20192);
   U7838 : OAI211_X1 port map( C1 => n19563, C2 => n19564, A => n19562, B => 
                           n19561, ZN => n20367);
   U20480 : NAND4_X1 port map( A1 => n18498, A2 => n18497, A3 => n18496, A4 => 
                           n18495, ZN => n20571);
   U11269 : INV_X1 port map( A => n20470, ZN => n5115);
   U11207 : NAND4_X1 port map( A1 => n18893, A2 => n18890, A3 => n18892, A4 => 
                           n18891, ZN => n20549);
   U21066 : OR2_X1 port map( A1 => n19542, A2 => n19541, ZN => n19544);
   U5610 : AOI21_X1 port map( B1 => n4289, B2 => n18933, A => n4288, ZN => 
                           n19155);
   U1023 : NAND2_X1 port map( A1 => n19008, A2 => n4425, ZN => n20149);
   U20909 : INV_X1 port map( A => n19155, ZN => n20101);
   U1394 : AND3_X1 port map( A1 => n19062, A2 => n1132, A3 => n1131, ZN => 
                           n20498);
   U1866 : NAND2_X1 port map( A1 => n19040, A2 => n5234, ZN => n20301);
   U8900 : NAND2_X1 port map( A1 => n24217, A2 => n17941, ZN => n1591);
   U17232 : AND3_X1 port map( A1 => n19506, A2 => n19505, A3 => n19504, ZN => 
                           n19777);
   U5651 : OR2_X1 port map( A1 => n20546, A2 => n20125, ZN => n19675);
   U664 : AND3_X1 port map( A1 => n18802, A2 => n18803, A3 => n18801, ZN => 
                           n21212);
   U21360 : AND3_X1 port map( A1 => n19931, A2 => n19930, A3 => n19929, ZN => 
                           n20999);
   U21246 : NOR3_X1 port map( A1 => n351, A2 => n19799, A3 => n19798, ZN => 
                           n19800);
   U21685 : AND3_X1 port map( A1 => n20542, A2 => n20541, A3 => n20540, ZN => 
                           n21422);
   U12080 : OAI21_X1 port map( B1 => n20548, B2 => n19677, A => n19676, ZN => 
                           n21436);
   U4331 : OAI21_X1 port map( B1 => n20131, B2 => n3833, A => n3831, ZN => 
                           n21550);
   U7110 : NAND2_X1 port map( A1 => n1995, A2 => n20201, ZN => n21445);
   U1812 : NAND2_X1 port map( A1 => n19961, A2 => n19960, ZN => n20948);
   U21618 : OAI211_X1 port map( C1 => n20398, C2 => n350, A => n20397, B => 
                           n20396, ZN => n21965);
   U11735 : OAI211_X1 port map( C1 => n20549, C2 => n20548, A => n5638, B => 
                           n5637, ZN => n21158);
   U3336 : NAND2_X1 port map( A1 => n742, A2 => n19822, ZN => n21319);
   U2999 : NAND2_X1 port map( A1 => n2104, A2 => n587, ZN => n21301);
   U1801 : NAND3_X1 port map( A1 => n20144, A2 => n5444, A3 => n5443, ZN => 
                           n21554);
   U1271 : NOR2_X1 port map( A1 => n20053, A2 => n20052, ZN => n21704);
   U598 : XNOR2_X1 port map( A => n21546, B => n21545, ZN => n22421);
   U1778 : XNOR2_X1 port map( A => n21187, B => n21186, ZN => n22592);
   U21103 : BUF_X1 port map( A => n23575, Z => n24396);
   U1263 : XNOR2_X1 port map( A => n21485, B => n21484, ZN => n22968);
   U738 : XNOR2_X1 port map( A => n21131, B => n21130, ZN => n22675);
   U584 : BUF_X1 port map( A => n21888, Z => n22401);
   U3384 : OR2_X1 port map( A1 => n772, A2 => n4371, ZN => n23265);
   U45 : AOI21_X1 port map( B1 => n21936, B2 => n21937, A => n22562, ZN => 
                           n22571);
   U23016 : NOR2_X1 port map( A1 => n22238, A2 => n22237, ZN => n23730);
   U1036 : AND2_X1 port map( A1 => n1587, A2 => n1585, ZN => n23273);
   U20246 : NAND2_X1 port map( A1 => n22213, A2 => n2314, ZN => n23743);
   U912 : AND2_X1 port map( A1 => n21113, A2 => n2595, ZN => n23074);
   U8694 : AND3_X1 port map( A1 => n2901, A2 => n3024, A3 => n3309, ZN => 
                           n23303);
   U243 : OR2_X1 port map( A1 => n22045, A2 => n22046, ZN => n22043);
   U1721 : NAND3_X1 port map( A1 => n4283, A2 => n1417, A3 => n4282, ZN => 
                           n23906);
   U1567 : CLKBUF_X1 port map( A => Key(25), Z => n21423);
   U1608 : CLKBUF_X1 port map( A => Key(189), Z => n21553);
   U12393 : XNOR2_X1 port map( A => n5950, B => Key(170), ZN => n6489);
   U2644 : NAND2_X1 port map( A1 => n4756, A2 => n5906, ZN => n8511);
   U5258 : AOI21_X1 port map( B1 => n7143, B2 => n7142, A => n2780, ZN => n8168
                           );
   U12832 : AOI22_X1 port map( A1 => n6864, A2 => n6466, B1 => n7216, B2 => 
                           n6465, ZN => n9147);
   U11965 : NOR2_X1 port map( A1 => n24944, A2 => n9463, ZN => n9351);
   U2456 : OAI211_X1 port map( C1 => n10146, C2 => n10145, A => n10144, B => 
                           n10143, ZN => n10654);
   U3368 : NAND4_X1 port map( A1 => n9030, A2 => n9031, A3 => n9029, A4 => 
                           n9032, ZN => n11039);
   U1197 : BUF_X1 port map( A => n10192, Z => n10829);
   U1239 : BUF_X1 port map( A => n11518, Z => n11525);
   U2377 : NAND2_X1 port map( A1 => n11202, A2 => n3011, ZN => n12023);
   U1495 : XNOR2_X1 port map( A => n12348, B => n12347, ZN => n13124);
   U2258 : OAI211_X1 port map( C1 => n13065, C2 => n5112, A => n3710, B => 
                           n2859, ZN => n13974);
   U1456 : INV_X1 port map( A => n16008, ZN => n3554);
   U1261 : BUF_X1 port map( A => n16428, Z => n244);
   U1467 : INV_X1 port map( A => n15706, ZN => n294);
   U2079 : INV_X1 port map( A => n16516, ZN => n17138);
   U7825 : NAND2_X1 port map( A1 => n16020, A2 => n2344, ZN => n16991);
   U2039 : OR2_X1 port map( A1 => n25200, A2 => n17208, ZN => n17017);
   U9019 : MUX2_X1 port map( A => n17318, B => n17317, S => n17316, Z => n18448
                           );
   U591 : XNOR2_X1 port map( A => n17957, B => n17956, ZN => n19380);
   U3972 : AOI22_X1 port map( A1 => n19249, A2 => n19248, B1 => n3620, B2 => 
                           n1098, ZN => n20426);
   U1846 : CLKBUF_X1 port map( A => n19494, Z => n20239);
   U4791 : INV_X1 port map( A => n23996, ZN => n22677);
   U4780 : INV_X1 port map( A => n23014, ZN => n23461);
   U207 : AND3_X2 port map( A1 => n3140, A2 => n20067, A3 => n19158, ZN => 
                           n21689);
   U24128 : BUF_X1 port map( A => n23275, Z => n24486);
   U7546 : NAND4_X2 port map( A1 => n2169, A2 => n19746, A3 => n19747, A4 => 
                           n1452, ZN => n21622);
   U7505 : OR2_X2 port map( A1 => n4123, A2 => n2153, ZN => n14221);
   U1096 : OR2_X2 port map( A1 => n16318, A2 => n16317, ZN => n18646);
   U608 : OAI21_X2 port map( B1 => n1409, B2 => n2890, A => n5384, ZN => n18429
                           );
   U19060 : NAND2_X2 port map( A1 => n16297, A2 => n16296, ZN => n17356);
   U1692 : AND2_X2 port map( A1 => n21920, A2 => n211, ZN => n23196);
   U3442 : NAND3_X2 port map( A1 => n4974, A2 => n16958, A3 => n4502, ZN => 
                           n18675);
   U6860 : BUF_X2 port map( A => n9345, Z => n9927);
   U653 : XNOR2_X2 port map( A => n7837, B => n7836, ZN => n9603);
   U1196 : AND2_X2 port map( A1 => n2392, A2 => n2390, ZN => n10302);
   U586 : NOR2_X2 port map( A1 => n5340, A2 => n10256, ZN => n10734);
   U833 : AND2_X2 port map( A1 => n4798, A2 => n4797, ZN => n14319);
   U9496 : XNOR2_X2 port map( A => n17697, B => n17696, ZN => n19445);
   U1007 : AND2_X2 port map( A1 => n4638, A2 => n4618, ZN => n13792);
   U11342 : AND3_X2 port map( A1 => n5185, A2 => n5186, A3 => n19829, ZN => 
                           n21738);
   U1046 : AND2_X2 port map( A1 => n16682, A2 => n16680, ZN => n17277);
   U176 : OAI21_X2 port map( B1 => n3818, B2 => n16606, A => n16605, ZN => 
                           n18694);
   U713 : OR2_X2 port map( A1 => n4501, A2 => n4500, ZN => n12147);
   U6328 : BUF_X2 port map( A => n18982, Z => n20014);
   U24197 : AND3_X2 port map( A1 => n1913, A2 => n963, A3 => n1911, ZN => 
                           n17293);
   U8787 : AND2_X2 port map( A1 => n15698, A2 => n16549, ZN => n2587);
   U502 : AND2_X2 port map( A1 => n4255, A2 => n4253, ZN => n11058);
   U19344 : MUX2_X2 port map( A => n16793, B => n16792, S => n1516, Z => n18602
                           );
   U401 : INV_X2 port map( A => n11084, ZN => n3119);
   U14582 : NOR2_X2 port map( A1 => n3337, A2 => n12639, ZN => n14198);
   U1029 : NAND2_X2 port map( A1 => n17036, A2 => n18925, ZN => n20336);
   U930 : OAI21_X2 port map( B1 => n20334, B2 => n20333, A => n20332, ZN => 
                           n22005);
   U980 : BUF_X2 port map( A => n15986, Z => n16141);
   U345 : OAI211_X2 port map( C1 => n8332, C2 => n10169, A => n4212, B => n2548
                           , ZN => n10596);
   U246 : NAND2_X2 port map( A1 => n21, A2 => n20, ZN => n13829);
   U10252 : OR2_X2 port map( A1 => n4089, A2 => n10636, ZN => n12167);
   U1129 : AND3_X2 port map( A1 => n867, A2 => n1857, A3 => n1858, ZN => n11045
                           );
   U2974 : NOR2_X2 port map( A1 => n575, A2 => n16580, ZN => n17881);
   U1280 : BUF_X2 port map( A => n6849, Z => n250);
   U9456 : NAND4_X2 port map( A1 => n3318, A2 => n3319, A3 => n15744, A4 => 
                           n16198, ZN => n17391);
   U570 : NAND2_X2 port map( A1 => n10231, A2 => n10230, ZN => n11704);
   U691 : NOR2_X2 port map( A1 => n14951, A2 => n14950, ZN => n15494);
   U536 : OR2_X2 port map( A1 => n5382, A2 => n5381, ZN => n12357);
   U1686 : NAND2_X2 port map( A1 => n4944, A2 => n4943, ZN => n14267);
   U1164 : XNOR2_X2 port map( A => n15400, B => n15399, ZN => n15694);
   U1277 : AND3_X2 port map( A1 => n12997, A2 => n12999, A3 => n12998, ZN => 
                           n14219);
   U643 : BUF_X2 port map( A => n18719, Z => n19497);
   U2502 : BUF_X1 port map( A => n7183, Z => n9949);
   U2666 : AND2_X2 port map( A1 => n6485, A2 => n6484, ZN => n7638);
   U511 : XNOR2_X2 port map( A => n8390, B => n8389, ZN => n10161);
   U2407 : BUF_X1 port map( A => n9769, Z => n10364);
   U963 : NOR2_X2 port map( A1 => n16421, A2 => n16420, ZN => n17445);
   U2304 : AND3_X1 port map( A1 => n2737, A2 => n5086, A3 => n2736, ZN => n1985
                           );
   U4580 : BUF_X1 port map( A => n9134, Z => n9953);
   U6054 : NOR2_X1 port map( A1 => n9461, A2 => n9459, ZN => n1470);
   U4438 : AND2_X1 port map( A1 => n9786, A2 => n10082, ZN => n9789);
   U2386 : AOI21_X1 port map( B1 => n10236, B2 => n10237, A => n10235, ZN => 
                           n11076);
   U717 : OAI211_X1 port map( C1 => n9444, C2 => n9443, A => n9442, B => n9441,
                           ZN => n12275);
   U2305 : BUF_X1 port map( A => n12625, Z => n12878);
   U323 : NAND3_X1 port map( A1 => n13557, A2 => n13556, A3 => n13555, ZN => 
                           n15444);
   U762 : XNOR2_X1 port map( A => n14531, B => n14530, ZN => n16394);
   U595 : BUF_X2 port map( A => n16765, Z => n17574);
   U21239 : OR3_X1 port map( A1 => n20244, A2 => n20241, A3 => n19937, ZN => 
                           n19789);
   U994 : OAI21_X2 port map( B1 => n20666, B2 => n19712, A => n19711, ZN => 
                           n21745);
   U3876 : OAI21_X2 port map( B1 => n20481, B2 => n20480, A => n1022, ZN => 
                           n21040);
   U1754 : BUF_X1 port map( A => n21540, Z => n22422);
   U1 : OAI21_X1 port map( B1 => n21374, B2 => n21373, A => n21372, ZN => 
                           n24473);
   U2 : NAND2_X1 port map( A1 => n1074, A2 => n21890, ZN => n23311);
   U4 : BUF_X1 port map( A => n22128, Z => n22966);
   U7 : BUF_X2 port map( A => n19953, Z => n20591);
   U13 : NOR2_X1 port map( A1 => n1014, A2 => n1010, ZN => n20338);
   U27 : XNOR2_X1 port map( A => n1387, B => n18556, ZN => n19084);
   U32 : MUX2_X1 port map( A => n15261, B => n15260, S => n24330, Z => n18074);
   U34 : NAND3_X1 port map( A1 => n14030, A2 => n14029, A3 => n76, ZN => n15506
                           );
   U37 : NAND4_X1 port map( A1 => n2302, A2 => n2303, A3 => n2301, A4 => n13723
                           , ZN => n15452);
   U43 : NOR2_X1 port map( A1 => n13625, A2 => n13624, ZN => n14678);
   U48 : NOR2_X1 port map( A1 => n8663, A2 => n8662, ZN => n25016);
   U82 : XNOR2_X2 port map( A => n21643, B => n21642, ZN => n22939);
   U105 : OR2_X2 port map( A1 => n17451, A2 => n17455, ZN => n3982);
   U122 : BUF_X2 port map( A => n16284, Z => n24540);
   U134 : AND3_X2 port map( A1 => n24647, A2 => n24646, A3 => n19357, ZN => 
                           n17714);
   U143 : AND3_X2 port map( A1 => n24767, A2 => n9663, A3 => n1943, ZN => 
                           n10630);
   U155 : BUF_X2 port map( A => n9992, Z => n24534);
   U169 : BUF_X1 port map( A => n15922, Z => n16464);
   U175 : OR2_X2 port map( A1 => n7569, A2 => n2026, ZN => n9191);
   U184 : AND2_X2 port map( A1 => n2117, A2 => n2116, ZN => n24974);
   U186 : AND2_X2 port map( A1 => n4706, A2 => n4708, ZN => n8352);
   U222 : BUF_X1 port map( A => n12226, Z => n24915);
   U250 : AND3_X2 port map( A1 => n4886, A2 => n1202, A3 => n4887, ZN => n4004)
                           ;
   U273 : NAND3_X2 port map( A1 => n24697, A2 => n1400, A3 => n4014, ZN => 
                           n2242);
   U275 : OR2_X2 port map( A1 => n18754, A2 => n18753, ZN => n19809);
   U290 : INV_X1 port map( A => n19166, ZN => n24584);
   U292 : OAI21_X1 port map( B1 => n20405, B2 => n20419, A => n20404, ZN => 
                           n20585);
   U293 : INV_X1 port map( A => n22953, ZN => n22959);
   U310 : XNOR2_X2 port map( A => n8048, B => n8047, ZN => n9864);
   U318 : OAI211_X2 port map( C1 => n12538, C2 => n1636, A => n1634, B => n1633
                           , ZN => n14268);
   U320 : OR2_X2 port map( A1 => n24259, A2 => n13516, ZN => n15476);
   U341 : XOR2_X1 port map( A => n14693, B => n14692, Z => n24532);
   U349 : NOR2_X2 port map( A1 => n16234, A2 => n1096, ZN => n17216);
   U351 : NOR2_X2 port map( A1 => n16944, A2 => n17611, ZN => n18677);
   U355 : NAND3_X1 port map( A1 => n20497, A2 => n24887, A3 => n20496, ZN => 
                           n24533);
   U367 : NOR2_X2 port map( A1 => n21827, A2 => n3890, ZN => n21837);
   U370 : BUF_X2 port map( A => n19041, Z => n19361);
   U372 : INV_X2 port map( A => n5692, ZN => n15375);
   U379 : CLKBUF_X1 port map( A => n9992, Z => n24535);
   U387 : XNOR2_X1 port map( A => n8894, B => n8895, ZN => n9992);
   U410 : XNOR2_X2 port map( A => n8284, B => n8283, ZN => n10113);
   U437 : XNOR2_X2 port map( A => n8166, B => n8165, ZN => n9564);
   U450 : OR2_X2 port map( A1 => n16071, A2 => n16070, ZN => n17165);
   U454 : NAND2_X2 port map( A1 => n20088, A2 => n20087, ZN => n21676);
   U457 : BUF_X1 port map( A => n9127, Z => n10062);
   U467 : CLKBUF_X1 port map( A => n16393, Z => n24537);
   U476 : XNOR2_X1 port map( A => n14536, B => n14535, ZN => n16393);
   U498 : XNOR2_X1 port map( A => n15050, B => n15049, ZN => n16284);
   U501 : NAND3_X2 port map( A1 => n4642, A2 => n6382, A3 => n4641, ZN => n8370
                           );
   U509 : BUF_X1 port map( A => n17313, Z => n24542);
   U517 : OAI211_X1 port map( C1 => n15660, C2 => n15659, A => n5502, B => 
                           n15658, ZN => n17313);
   U540 : XNOR2_X1 port map( A => n20314, B => n20315, ZN => n22809);
   U544 : OAI211_X2 port map( C1 => n20240, C2 => n20239, A => n20238, B => 
                           n4750, ZN => n21070);
   U554 : OAI211_X2 port map( C1 => n19861, C2 => n19860, A => n19859, B => 
                           n19858, ZN => n21136);
   U557 : XNOR2_X2 port map( A => n18048, B => n18049, ZN => n19596);
   U558 : XNOR2_X2 port map( A => n4583, B => n4581, ZN => n16334);
   U562 : BUF_X2 port map( A => n19878, Z => n20555);
   U583 : AND2_X2 port map( A1 => n5308, A2 => n5307, ZN => n16037);
   U590 : AND2_X2 port map( A1 => n5271, A2 => n5274, ZN => n11201);
   U615 : NAND2_X2 port map( A1 => n3226, A2 => n3228, ZN => n23805);
   U621 : XNOR2_X2 port map( A => n14784, B => n14783, ZN => n16246);
   U623 : AND3_X2 port map( A1 => n2144, A2 => n4817, A3 => n4818, ZN => n17816
                           );
   U626 : XNOR2_X1 port map( A => n8092, B => n8091, ZN => n9874);
   U627 : OAI21_X2 port map( B1 => n16370, B2 => n17460, A => n16369, ZN => 
                           n18610);
   U629 : BUF_X1 port map( A => n16470, Z => n24551);
   U636 : XNOR2_X1 port map( A => n15450, B => n15449, ZN => n16470);
   U638 : MUX2_X2 port map( A => n12790, B => n12789, S => n13027, Z => n13864)
                           ;
   U642 : OAI211_X2 port map( C1 => n19996, C2 => n19995, A => n19994, B => 
                           n19993, ZN => n20914);
   U657 : AND4_X2 port map( A1 => n2687, A2 => n19773, A3 => n19772, A4 => 
                           n2685, ZN => n21608);
   U673 : XNOR2_X1 port map( A => n2415, B => n2416, ZN => n21829);
   U678 : OAI21_X2 port map( B1 => n18829, B2 => n19087, A => n4194, ZN => 
                           n20353);
   U681 : NOR2_X2 port map( A1 => n19808, A2 => n19807, ZN => n20982);
   U682 : XNOR2_X2 port map( A => n8338, B => n8337, ZN => n9837);
   U683 : AND2_X2 port map( A1 => n972, A2 => n971, ZN => n23810);
   U686 : XNOR2_X2 port map( A => n14661, B => n14660, ZN => n16076);
   U741 : BUF_X1 port map( A => n13360, Z => n24554);
   U766 : XNOR2_X1 port map( A => n12126, B => n12125, ZN => n13360);
   U780 : NAND2_X2 port map( A1 => n1751, A2 => n9202, ZN => n10584);
   U783 : NOR2_X2 port map( A1 => n10653, A2 => n10652, ZN => n12146);
   U794 : XNOR2_X2 port map( A => n8196, B => n8195, ZN => n10148);
   U808 : OAI211_X2 port map( C1 => n20582, C2 => n20583, A => n20581, B => 
                           n20580, ZN => n21053);
   U816 : NOR2_X2 port map( A1 => n3800, A2 => n9667, ZN => n10789);
   U840 : NOR2_X1 port map( A1 => n12723, A2 => n12722, ZN => n14435);
   U872 : AOI22_X2 port map( A1 => n4713, A2 => n20349, B1 => n20351, B2 => 
                           n20350, ZN => n21058);
   U901 : XNOR2_X2 port map( A => n11988, B => n11989, ZN => n13267);
   U902 : NOR2_X2 port map( A1 => n1866, A2 => n12779, ZN => n14669);
   U905 : XNOR2_X2 port map( A => n8642, B => n8641, ZN => n10104);
   U911 : AND3_X2 port map( A1 => n9835, A2 => n9833, A3 => n9834, ZN => n10548
                           );
   U922 : NOR2_X2 port map( A1 => n15903, A2 => n15902, ZN => n17039);
   U923 : OAI22_X2 port map( A1 => n990, A2 => n14017, B1 => n13534, B2 => 
                           n13607, ZN => n15033);
   U926 : XNOR2_X2 port map( A => n21443, B => n21442, ZN => n22965);
   U941 : XNOR2_X2 port map( A => n20495, B => n20494, ZN => n21856);
   U955 : CLKBUF_X1 port map( A => n24510, Z => n24561);
   U956 : XNOR2_X1 port map( A => n21218, B => n21219, ZN => n24510);
   U957 : XNOR2_X2 port map( A => n15346, B => n15345, ZN => n15953);
   U962 : AND2_X2 port map( A1 => n1947, A2 => n1946, ZN => n16795);
   U966 : XNOR2_X2 port map( A => n11850, B => n1384, ZN => n12899);
   U1038 : AOI21_X2 port map( B1 => n16180, B2 => n16179, A => n16178, ZN => 
                           n17400);
   U1060 : NAND2_X2 port map( A1 => n5092, A2 => n5091, ZN => n21505);
   U1065 : INV_X1 port map( A => n12902, ZN => n4499);
   U1089 : NOR2_X1 port map( A1 => n17556, A2 => n4436, ZN => n19263);
   U1092 : OAI211_X2 port map( C1 => n7602, C2 => n7603, A => n3007, B => n3006
                           , ZN => n8446);
   U1093 : NOR2_X2 port map( A1 => n16593, A2 => n24699, ZN => n18685);
   U1095 : NOR2_X2 port map( A1 => n17448, A2 => n17447, ZN => n18456);
   U1102 : OAI211_X2 port map( C1 => n2638, C2 => n2636, A => n2637, B => n2635
                           , ZN => n5376);
   U1103 : NOR2_X1 port map( A1 => n13112, A2 => n13110, ZN => n12853);
   U1159 : AND2_X1 port map( A1 => n20941, A2 => n20942, ZN => n23612);
   U1161 : INV_X1 port map( A => n20670, ZN => n24567);
   U1167 : INV_X1 port map( A => n17364, ZN => n24569);
   U1171 : INV_X1 port map( A => n17051, ZN => n24570);
   U1181 : OR2_X1 port map( A1 => n16902, A2 => n2562, ZN => n45);
   U1187 : XNOR2_X1 port map( A => n14552, B => n14551, ZN => n15849);
   U1194 : INV_X1 port map( A => n14435, ZN => n24571);
   U1201 : XNOR2_X1 port map( A => n11882, B => n11883, ZN => n4241);
   U1204 : BUF_X2 port map( A => n13077, Z => n24573);
   U1213 : INV_X1 port map( A => n11112, ZN => n24574);
   U1217 : OR2_X1 port map( A1 => n262, A2 => n9281, ZN => n25174);
   U1224 : OAI211_X1 port map( C1 => n7152, C2 => n7217, A => n7150, B => n7149
                           , ZN => n8627);
   U1226 : INV_X1 port map( A => n7864, ZN => n24576);
   U1228 : NAND3_X1 port map( A1 => n25184, A2 => n6501, A3 => n6502, ZN => 
                           n8527);
   U1231 : INV_X1 port map( A => n7734, ZN => n24578);
   U1242 : CLKBUF_X1 port map( A => Key(113), Z => n2036);
   U1258 : CLKBUF_X1 port map( A => Key(166), Z => n62);
   U1265 : INV_X1 port map( A => n6975, ZN => n24579);
   U1267 : CLKBUF_X1 port map( A => Key(107), Z => n2228);
   U1268 : OR2_X1 port map( A1 => n23483, A2 => n23499, ZN => n24874);
   U1270 : OR2_X1 port map( A1 => n23979, A2 => n24440, ZN => n24873);
   U1282 : OR2_X1 port map( A1 => n23030, A2 => n22539, ZN => n21352);
   U1286 : AND2_X1 port map( A1 => n23052, A2 => n23047, ZN => n23039);
   U1288 : INV_X1 port map( A => n23219, ZN => n23231);
   U1290 : CLKBUF_X1 port map( A => n23799, Z => n24920);
   U1291 : AOI21_X1 port map( B1 => n25050, B2 => n22165, A => n22164, ZN => 
                           n25026);
   U1293 : OR2_X1 port map( A1 => n23297, A2 => n22395, ZN => n22510);
   U1298 : INV_X1 port map( A => n1075, ZN => n23320);
   U1299 : OR2_X1 port map( A1 => n23817, A2 => n891, ZN => n21355);
   U1317 : AND3_X1 port map( A1 => n1068, A2 => n1905, A3 => n1065, ZN => 
                           n23420);
   U1361 : OR2_X1 port map( A1 => n21894, A2 => n1076, ZN => n1075);
   U1366 : AND2_X1 port map( A1 => n25138, A2 => n2038, ZN => n23129);
   U1367 : AOI21_X1 port map( B1 => n21927, B2 => n21926, A => n21925, ZN => 
                           n24889);
   U1369 : MUX2_X1 port map( A => n22038, B => n22037, S => n603, Z => n24880);
   U1374 : MUX2_X1 port map( A => n22372, B => n22371, S => n22680, Z => n24948
                           );
   U1376 : NOR2_X1 port map( A1 => n21923, A2 => n21922, ZN => n21927);
   U1381 : AND2_X1 port map( A1 => n24673, A2 => n24672, ZN => n22074);
   U1385 : OAI211_X1 port map( C1 => n4098, C2 => n3213, A => n22977, B => 
                           n24724, ZN => n2901);
   U1391 : INV_X1 port map( A => n22282, ZN => n24631);
   U1399 : INV_X1 port map( A => n22677, ZN => n24869);
   U1400 : XNOR2_X1 port map( A => n21203, B => n21202, ZN => n22798);
   U1402 : XNOR2_X1 port map( A => n20575, B => n20574, ZN => n22679);
   U1413 : XNOR2_X1 port map( A => n20802, B => n20801, ZN => n22459);
   U1415 : BUF_X2 port map( A => n21665, Z => n24898);
   U1421 : NAND3_X1 port map( A1 => n24138, A2 => n5123, A3 => n19920, ZN => 
                           n21647);
   U1436 : AND2_X1 port map( A1 => n3903, A2 => n25028, ZN => n21273);
   U1512 : OR2_X1 port map( A1 => n19674, A2 => n20124, ZN => n5262);
   U1520 : NOR2_X1 port map( A1 => n19849, A2 => n19658, ZN => n19659);
   U1522 : NOR2_X1 port map( A1 => n20224, A2 => n20498, ZN => n24682);
   U1547 : NAND2_X1 port map( A1 => n24733, A2 => n18905, ZN => n20546);
   U1554 : AND2_X1 port map( A1 => n100, A2 => n20507, ZN => n24644);
   U1561 : AND2_X1 port map( A1 => n20557, A2 => n3480, ZN => n24749);
   U1614 : INV_X1 port map( A => n20523, ZN => n20131);
   U1681 : OR2_X1 port map( A1 => n19889, A2 => n20319, ZN => n2180);
   U1689 : INV_X1 port map( A => n20290, ZN => n24581);
   U1691 : OAI21_X1 port map( B1 => n24638, B2 => n19028, A => n24637, ZN => 
                           n4067);
   U1700 : NAND2_X1 port map( A1 => n3508, A2 => n18879, ZN => n20523);
   U1709 : OR2_X1 port map( A1 => n20169, A2 => n20173, ZN => n19958);
   U1712 : INV_X1 port map( A => n25034, ZN => n24829);
   U1727 : OR2_X1 port map( A1 => n18787, A2 => n18786, ZN => n20473);
   U1743 : AND2_X1 port map( A1 => n25158, A2 => n25157, ZN => n20510);
   U1748 : AND3_X1 port map( A1 => n17803, A2 => n17802, A3 => n17801, ZN => 
                           n20111);
   U1762 : AND2_X1 port map( A1 => n18976, A2 => n19460, ZN => n24638);
   U1763 : NAND3_X1 port map( A1 => n25105, A2 => n2304, A3 => n18716, ZN => 
                           n20042);
   U1765 : INV_X1 port map( A => n24172, ZN => n24637);
   U1768 : INV_X1 port map( A => n19037, ZN => n24582);
   U1789 : INV_X1 port map( A => n25002, ZN => n24809);
   U1807 : OR2_X1 port map( A1 => n19548, A2 => n24929, ZN => n24717);
   U1817 : INV_X1 port map( A => n16737, ZN => n24719);
   U1862 : INV_X1 port map( A => n17497, ZN => n24583);
   U1863 : XNOR2_X1 port map( A => n18555, B => n24769, ZN => n1387);
   U1875 : NAND2_X1 port map( A1 => n2829, A2 => n24615, ZN => n18523);
   U1885 : MUX2_X1 port map( A => n17301, B => n17300, S => n17299, Z => n17303
                           );
   U1914 : AND2_X1 port map( A1 => n17141, A2 => n1653, ZN => n24688);
   U1927 : NOR2_X1 port map( A1 => n16255, A2 => n16256, ZN => n17016);
   U1930 : AND2_X1 port map( A1 => n17293, A2 => n17283, ZN => n24775);
   U1937 : INV_X1 port map( A => n17249, ZN => n17252);
   U1952 : INV_X1 port map( A => n17081, ZN => n16895);
   U1967 : OAI21_X1 port map( B1 => n16280, B2 => n25180, A => n16278, ZN => 
                           n17352);
   U1970 : OR2_X1 port map( A1 => n15931, A2 => n16450, ZN => n25116);
   U1986 : NAND2_X1 port map( A1 => n16364, A2 => n16363, ZN => n523);
   U1997 : OAI21_X1 port map( B1 => n16293, B2 => n24842, A => n24841, ZN => 
                           n16297);
   U2019 : AND2_X1 port map( A1 => n257, A2 => n16447, ZN => n24774);
   U2036 : XOR2_X1 port map( A => n15092, B => n15091, Z => n24919);
   U2037 : INV_X1 port map( A => n15782, ZN => n24586);
   U2045 : INV_X1 port map( A => n15821, ZN => n24587);
   U2053 : MUX2_X2 port map( A => n14184, B => n14183, S => n14182, Z => n14642
                           );
   U2055 : OAI21_X1 port map( B1 => n13721, B2 => n13720, A => n13719, ZN => 
                           n15253);
   U2063 : XNOR2_X1 port map( A => n14703, B => n14553, ZN => n15392);
   U2077 : NAND2_X1 port map( A1 => n13698, A2 => n2741, ZN => n14690);
   U2123 : NAND3_X1 port map( A1 => n13919, A2 => n13920, A3 => n760, ZN => 
                           n15350);
   U2155 : NAND3_X1 port map( A1 => n24776, A2 => n2151, A3 => n2150, ZN => 
                           n15054);
   U2187 : OR2_X1 port map( A1 => n13675, A2 => n13674, ZN => n24691);
   U2197 : INV_X1 port map( A => n13888, ZN => n24710);
   U2201 : BUF_X1 port map( A => n12850, Z => n14335);
   U2202 : AND3_X1 port map( A1 => n2906, A2 => n24094, A3 => n2905, ZN => 
                           n13839);
   U2212 : AND3_X1 port map( A1 => n5724, A2 => n12762, A3 => n5723, ZN => 
                           n24949);
   U2220 : INV_X1 port map( A => n14059, ZN => n24785);
   U2233 : NAND2_X1 port map( A1 => n498, A2 => n24854, ZN => n14158);
   U2257 : OR3_X1 port map( A1 => n11319, A2 => n13230, A3 => n25080, ZN => 
                           n11331);
   U2319 : INV_X1 port map( A => n14166, ZN => n24773);
   U2331 : INV_X1 port map( A => n3876, ZN => n24617);
   U2364 : AND2_X1 port map( A1 => n13282, A2 => n24988, ZN => n12931);
   U2373 : XNOR2_X1 port map( A => n12115, B => n12116, ZN => n12956);
   U2423 : INV_X1 port map( A => n11689, ZN => n24778);
   U2442 : NAND3_X1 port map( A1 => n24761, A2 => n9343, A3 => n24760, ZN => 
                           n25090);
   U2486 : OR2_X1 port map( A1 => n10725, A2 => n11116, ZN => n24760);
   U2508 : INV_X1 port map( A => n10914, ZN => n24753);
   U2529 : OAI21_X1 port map( B1 => n10285, B2 => n10875, A => n11117, ZN => 
                           n24761);
   U2533 : OR2_X1 port map( A1 => n11066, A2 => n11068, ZN => n25103);
   U2544 : NOR2_X1 port map( A1 => n11518, A2 => n11519, ZN => n10918);
   U2552 : OR2_X1 port map( A1 => n10753, A2 => n10451, ZN => n25156);
   U2568 : INV_X1 port map( A => n11171, ZN => n24591);
   U2573 : NAND4_X1 port map( A1 => n8575, A2 => n8572, A3 => n8574, A4 => 
                           n8573, ZN => n24957);
   U2630 : NAND2_X1 port map( A1 => n9819, A2 => n655, ZN => n10951);
   U2634 : NOR2_X1 port map( A1 => n9624, A2 => n3674, ZN => n4871);
   U2699 : OR2_X1 port map( A1 => n7670, A2 => n7671, ZN => n25152);
   U2716 : OR2_X1 port map( A1 => n7596, A2 => n24772, ZN => n3007);
   U2720 : INV_X1 port map( A => n7688, ZN => n7148);
   U2771 : AND3_X1 port map( A1 => n25186, A2 => n6453, A3 => n6452, ZN => 
                           n7691);
   U2776 : OR2_X1 port map( A1 => n873, A2 => n6361, ZN => n24878);
   U2792 : BUF_X1 port map( A => n6577, Z => n6752);
   U2798 : CLKBUF_X1 port map( A => Key(106), Z => n173);
   U2808 : OR2_X1 port map( A1 => n6504, A2 => n6503, ZN => n25184);
   U2819 : AND3_X1 port map( A1 => n5001, A2 => n5002, A3 => n6734, ZN => n6868
                           );
   U2825 : OR2_X1 port map( A1 => n6335, A2 => n6332, ZN => n6440);
   U2836 : OR2_X1 port map( A1 => n6244, A2 => n6119, ZN => n6840);
   U2837 : AND2_X1 port map( A1 => n6069, A2 => n6971, ZN => n24810);
   U2850 : INV_X1 port map( A => n6480, ZN => n6290);
   U2864 : CLKBUF_X1 port map( A => n6845, Z => n7027);
   U2878 : CLKBUF_X1 port map( A => n6133, Z => n6543);
   U2885 : INV_X1 port map( A => n7758, ZN => n432);
   U2888 : OR2_X2 port map( A1 => n6927, A2 => n6928, ZN => n7947);
   U2891 : AND2_X1 port map( A1 => n9066, A2 => n9067, ZN => n8221);
   U2894 : MUX2_X1 port map( A => n7995, B => n7994, S => n7993, Z => n7996);
   U2911 : AOI21_X1 port map( B1 => n24599, B2 => n10169, A => n9814, ZN => 
                           n25187);
   U2928 : OR2_X1 port map( A1 => n7059, A2 => n7809, ZN => n25117);
   U2931 : XNOR2_X1 port map( A => n8632, B => n8631, ZN => n9773);
   U2934 : XNOR2_X1 port map( A => n8331, B => n8330, ZN => n10166);
   U2969 : INV_X1 port map( A => n24944, ZN => n24853);
   U3011 : XNOR2_X1 port map( A => n7571, B => n7570, ZN => n1595);
   U3018 : BUF_X1 port map( A => n9859, Z => n238);
   U3026 : OR2_X1 port map( A1 => n9961, A2 => n9468, ZN => n24804);
   U3040 : AOI22_X1 port map( A1 => n9422, A2 => n9421, B1 => n9751, B2 => 
                           n9420, ZN => n9432);
   U3055 : NOR2_X1 port map( A1 => n24575, A2 => n10082, ZN => n25163);
   U3056 : OR2_X1 port map( A1 => n9362, A2 => n9363, ZN => n25148);
   U3065 : XNOR2_X1 port map( A => n8002, B => n8001, ZN => n9905);
   U3088 : OAI21_X1 port map( B1 => n262, B2 => n24927, A => n24804, ZN => 
                           n1186);
   U3108 : OAI21_X1 port map( B1 => n9920, B2 => n24844, A => n24843, ZN => 
                           n7044);
   U3110 : OR2_X1 port map( A1 => n24526, A2 => n10477, ZN => n24799);
   U3124 : OR2_X1 port map( A1 => n10910, A2 => n24753, ZN => n24817);
   U3128 : INV_X1 port map( A => n12121, ZN => n25166);
   U3136 : OR2_X1 port map( A1 => n10958, A2 => n10703, ZN => n3244);
   U3138 : OR2_X1 port map( A1 => n10428, A2 => n10651, ZN => n10429);
   U3161 : OR2_X1 port map( A1 => n10368, A2 => n10369, ZN => n25134);
   U3178 : XNOR2_X1 port map( A => n12141, B => n12114, ZN => n24634);
   U3193 : BUF_X1 port map( A => n12611, Z => n12612);
   U3198 : OR2_X1 port map( A1 => n13108, A2 => n12674, ZN => n3829);
   U3203 : CLKBUF_X1 port map( A => n12583, Z => n13363);
   U3206 : XNOR2_X1 port map( A => n11389, B => n11956, ZN => n12786);
   U3214 : AOI22_X1 port map( A1 => n12798, A2 => n12476, B1 => n13041, B2 => 
                           n13040, ZN => n12763);
   U3215 : OR2_X1 port map( A1 => n12793, A2 => n24750, ZN => n12566);
   U3219 : NOR2_X1 port map( A1 => n12744, A2 => n13101, ZN => n13188);
   U3243 : AND2_X1 port map( A1 => n13341, A2 => n12840, ZN => n12960);
   U3261 : NAND3_X1 port map( A1 => n5724, A2 => n12762, A3 => n5723, ZN => 
                           n13795);
   U3264 : INV_X1 port map( A => n231, ZN => n12958);
   U3278 : OR2_X1 port map( A1 => n12879, A2 => n12878, ZN => n2888);
   U3285 : AND2_X1 port map( A1 => n297, A2 => n3717, ZN => n1027);
   U3287 : AND2_X1 port map( A1 => n14079, A2 => n14078, ZN => n25099);
   U3293 : INV_X1 port map( A => n13636, ZN => n24679);
   U3294 : OR2_X1 port map( A1 => n24745, A2 => n24347, ZN => n24744);
   U3310 : OR2_X1 port map( A1 => n13284, A2 => n25191, ZN => n12929);
   U3311 : AND2_X1 port map( A1 => n14083, A2 => n14073, ZN => n24815);
   U3312 : OR2_X1 port map( A1 => n13515, A2 => n297, ZN => n3536);
   U3322 : OR2_X1 port map( A1 => n14243, A2 => n4116, ZN => n13639);
   U3328 : OR2_X1 port map( A1 => n13896, A2 => n13895, ZN => n13897);
   U3330 : OR2_X1 port map( A1 => n14058, A2 => n12468, ZN => n24776);
   U3337 : XNOR2_X1 port map( A => n14919, B => n14865, ZN => n14331);
   U3351 : OR2_X1 port map( A1 => n13944, A2 => n14302, ZN => n1400);
   U3390 : OR2_X1 port map( A1 => n15612, A2 => n15611, ZN => n15860);
   U3393 : INV_X1 port map( A => n24551, ZN => n24822);
   U3395 : XNOR2_X1 port map( A => n13836, B => n13835, ZN => n16186);
   U3402 : INV_X1 port map( A => n1365, ZN => n15801);
   U3403 : OR2_X1 port map( A1 => n16390, A2 => n15977, ZN => n15852);
   U3417 : AND2_X1 port map( A1 => n24919, A2 => n16360, ZN => n24842);
   U3423 : OR2_X1 port map( A1 => n15938, A2 => n16016, ZN => n16254);
   U3436 : XNOR2_X1 port map( A => n14520, B => n14519, ZN => n15804);
   U3437 : MUX2_X1 port map( A => n15600, B => n15599, S => n16063, Z => n15601
                           );
   U3470 : OR2_X1 port map( A1 => n3406, A2 => n16230, ZN => n5023);
   U3475 : INV_X1 port map( A => n381, ZN => n24655);
   U3479 : INV_X1 port map( A => n1261, ZN => n24797);
   U3489 : OR2_X1 port map( A1 => n17276, A2 => n17273, ZN => n16746);
   U3492 : OR2_X1 port map( A1 => n15266, A2 => n2253, ZN => n2250);
   U3493 : OR2_X1 port map( A1 => n17277, A2 => n17249, ZN => n1624);
   U3494 : OR2_X1 port map( A1 => n16809, A2 => n17478, ZN => n2372);
   U3498 : OR2_X1 port map( A1 => n16702, A2 => n16618, ZN => n751);
   U3499 : AOI22_X1 port map( A1 => n17144, A2 => n16691, B1 => n16985, B2 => 
                           n24688, ZN => n16695);
   U3506 : OR2_X1 port map( A1 => n16753, A2 => n17293, ZN => n17544);
   U3523 : INV_X1 port map( A => n16902, ZN => n2561);
   U3545 : AND2_X1 port map( A1 => n17326, A2 => n17319, ZN => n1409);
   U3550 : OAI21_X1 port map( B1 => n17152, B2 => n17151, A => n17150, ZN => 
                           n18060);
   U3568 : XNOR2_X1 port map( A => n18532, B => n4023, ZN => n17835);
   U3575 : INV_X1 port map( A => n17677, ZN => n24662);
   U3577 : OR2_X1 port map( A1 => n24759, A2 => n24457, ZN => n647);
   U3578 : OR2_X1 port map( A1 => n18816, A2 => n19359, ZN => n19213);
   U3591 : AND2_X1 port map( A1 => n19057, A2 => n988, ZN => n524);
   U3599 : BUF_X1 port map( A => n19485, Z => n240);
   U3604 : BUF_X1 port map( A => n17556, Z => n18919);
   U3616 : INV_X1 port map( A => n18830, ZN => n19597);
   U3636 : INV_X1 port map( A => n19436, ZN => n19435);
   U3640 : INV_X1 port map( A => n18493, ZN => n24728);
   U3645 : INV_X1 port map( A => n20615, ZN => n24835);
   U3648 : XNOR2_X1 port map( A => n17074, B => n17073, ZN => n4291);
   U3653 : CLKBUF_X1 port map( A => n19065, Z => n19239);
   U3658 : OR2_X1 port map( A1 => n18909, A2 => n19570, ZN => n24099);
   U3676 : AND2_X1 port map( A1 => n19491, A2 => n19492, ZN => n25131);
   U3683 : OR2_X1 port map( A1 => n19094, A2 => n25067, ZN => n19378);
   U3684 : INV_X1 port map( A => n988, ZN => n280);
   U3695 : AOI22_X1 port map( A1 => n19421, A2 => n19166, B1 => n19417, B2 => 
                           n19420, ZN => n4580);
   U3773 : INV_X1 port map( A => n1155, ZN => n3016);
   U3775 : OR2_X1 port map( A1 => n19403, A2 => n19186, ZN => n18893);
   U3791 : NAND2_X1 port map( A1 => n18737, A2 => n18738, ZN => n20183);
   U3832 : INV_X1 port map( A => n19904, ZN => n24681);
   U3838 : OR2_X1 port map( A1 => n19875, A2 => n20022, ZN => n20564);
   U3855 : NAND2_X1 port map( A1 => n1613, A2 => n4176, ZN => n1326);
   U3860 : XNOR2_X1 port map( A => n22005, B => n21606, ZN => n21343);
   U3872 : AND2_X1 port map( A1 => n22483, A2 => n22901, ZN => n24718);
   U3881 : OAI21_X1 port map( B1 => n20363, B2 => n24078, A => n18825, ZN => 
                           n21572);
   U3944 : INV_X1 port map( A => n3213, ZN => n25123);
   U3945 : AND2_X1 port map( A1 => n22239, A2 => n22241, ZN => n24666);
   U3969 : AND2_X1 port map( A1 => n22454, A2 => n22323, ZN => n22452);
   U3975 : OR2_X1 port map( A1 => n24415, A2 => n22138, ZN => n2828);
   U3976 : OR2_X1 port map( A1 => n24881, A2 => n22387, ZN => n24724);
   U4034 : AOI21_X1 port map( B1 => n4062, B2 => n1679, A => n22113, ZN => 
                           n23578);
   U4036 : AND2_X1 port map( A1 => n3895, A2 => n21822, ZN => n24698);
   U4038 : NAND3_X1 port map( A1 => n22277, A2 => n22276, A3 => n1507, ZN => 
                           n23250);
   U4041 : AOI21_X1 port map( B1 => n25050, B2 => n22165, A => n22164, ZN => 
                           n23692);
   U4048 : NOR2_X1 port map( A1 => n23723, A2 => n23714, ZN => n23696);
   U4058 : OAI21_X1 port map( B1 => n24322, B2 => n22281, A => n24631, ZN => 
                           n3718);
   U4117 : CLKBUF_X1 port map( A => n23478, Z => n23494);
   U4134 : OR2_X1 port map( A1 => n22637, A2 => n23595, ZN => n24668);
   U4136 : OR2_X1 port map( A1 => n23930, A2 => n24948, ZN => n24831);
   U4139 : CLKBUF_X1 port map( A => Key(46), Z => n886);
   U4181 : CLKBUF_X1 port map( A => Key(94), Z => n3115);
   U4184 : CLKBUF_X1 port map( A => Key(79), Z => n2042);
   U4189 : CLKBUF_X1 port map( A => Key(32), Z => n2100);
   U4208 : CLKBUF_X1 port map( A => Key(149), Z => n21711);
   U4231 : OAI211_X1 port map( C1 => n21763, C2 => n22639, A => n22638, B => 
                           n24668, ZN => n4782);
   U4249 : INV_X1 port map( A => n2215, ZN => n5484);
   U4281 : OR2_X1 port map( A1 => n25572, A2 => n288, ZN => n24594);
   U4305 : AND2_X1 port map( A1 => n7865, A2 => n24576, ZN => n24595);
   U4313 : INV_X1 port map( A => n7896, ZN => n24861);
   U4317 : INV_X1 port map( A => n7600, ZN => n24772);
   U4321 : OR2_X1 port map( A1 => n7879, A2 => n7882, ZN => n24596);
   U4334 : NOR2_X1 port map( A1 => n7581, A2 => n7882, ZN => n24597);
   U4339 : AND2_X1 port map( A1 => n7313, A2 => n7883, ZN => n7881);
   U4366 : XOR2_X1 port map( A => n9035, B => n5014, Z => n24598);
   U4370 : XOR2_X1 port map( A => n8326, B => n5619, Z => n24599);
   U4402 : XOR2_X1 port map( A => n9141, B => n1869, Z => n24600);
   U4409 : INV_X1 port map( A => n11004, ZN => n24622);
   U4421 : XNOR2_X1 port map( A => n11019, B => n11018, ZN => n12656);
   U4442 : INV_X1 port map( A => n12656, ZN => n24640);
   U4464 : OAI21_X1 port map( B1 => n4061, B2 => n3343, A => n3342, ZN => 
                           n13931);
   U4468 : INV_X1 port map( A => n13931, ZN => n25128);
   U4483 : NOR2_X1 port map( A1 => n14247, A2 => n13935, ZN => n24602);
   U4494 : INV_X1 port map( A => n12995, ZN => n24750);
   U4498 : XNOR2_X1 port map( A => n11327, B => n11326, ZN => n12791);
   U4510 : INV_X1 port map( A => n13975, ZN => n24713);
   U4557 : OR2_X1 port map( A1 => n14747, A2 => n15625, ZN => n24603);
   U4595 : AND2_X1 port map( A1 => n16796, A2 => n16550, ZN => n24604);
   U4640 : INV_X1 port map( A => n16809, ZN => n24660);
   U4682 : INV_X1 port map( A => n19477, ZN => n24803);
   U4696 : OR2_X1 port map( A1 => n19478, A2 => n5070, ZN => n24605);
   U4704 : INV_X1 port map( A => n19353, ZN => n19444);
   U4716 : XOR2_X1 port map( A => n18511, B => n18510, Z => n24606);
   U4771 : INV_X1 port map( A => n20346, ZN => n20281);
   U4792 : INV_X1 port map( A => n22804, ZN => n25160);
   U4796 : XNOR2_X1 port map( A => n20974, B => n20973, ZN => n22917);
   U4822 : INV_X1 port map( A => n22917, ZN => n24674);
   U4846 : XOR2_X1 port map( A => n21125, B => n21124, Z => n24607);
   U4862 : NAND2_X1 port map( A1 => n21838, A2 => n22354, ZN => n24608);
   U4879 : AND2_X1 port map( A1 => n4112, A2 => n24334, ZN => n24609);
   U4930 : OR2_X1 port map( A1 => n2671, A2 => n22422, ZN => n24610);
   U4940 : OR2_X1 port map( A1 => n23579, A2 => n23578, ZN => n24611);
   U4951 : OR2_X1 port map( A1 => n23196, A2 => n23195, ZN => n24612);
   U4962 : OR2_X1 port map( A1 => n23904, A2 => n607, ZN => n24613);
   U5011 : NAND2_X1 port map( A1 => n16702, A2 => n16703, ZN => n16709);
   U5050 : NAND2_X1 port map( A1 => n16443, A2 => n16242, ZN => n1095);
   U5071 : XNOR2_X2 port map( A => n15519, B => n15518, ZN => n16242);
   U5123 : OR2_X1 port map( A1 => n15473, A2 => n17202, ZN => n24615);
   U5219 : NAND2_X1 port map( A1 => n7992, A2 => n7993, ZN => n7501);
   U5249 : NAND2_X1 port map( A1 => n12854, A2 => n13112, ZN => n12206);
   U5253 : AND3_X2 port map( A1 => n24618, A2 => n24848, A3 => n9924, ZN => 
                           n10799);
   U5304 : NAND2_X1 port map( A1 => n24847, A2 => n9920, ZN => n24618);
   U5384 : NOR2_X1 port map( A1 => n24604, A2 => n5375, ZN => n15703);
   U5396 : BUF_X1 port map( A => n22217, Z => n24918);
   U5398 : NAND2_X1 port map( A1 => n24729, A2 => n22729, ZN => n2364);
   U5428 : XNOR2_X2 port map( A => n20858, B => n20859, ZN => n22729);
   U5432 : NAND2_X1 port map( A1 => n15044, A2 => n15043, ZN => n14493);
   U5436 : NAND3_X1 port map( A1 => n13780, A2 => n14160, A3 => n13954, ZN => 
                           n15043);
   U5452 : NAND3_X1 port map( A1 => n19221, A2 => n5461, A3 => n25010, ZN => 
                           n5442);
   U5455 : NAND2_X1 port map( A1 => n19371, A2 => n24424, ZN => n19221);
   U5464 : XNOR2_X2 port map( A => n24619, B => n15405, ZN => n15656);
   U5471 : XNOR2_X1 port map( A => n14186, B => n4834, ZN => n24619);
   U5472 : NAND2_X1 port map( A1 => n24330, A2 => n17422, ZN => n17429);
   U5489 : NOR2_X1 port map( A1 => n595, A2 => n24620, ZN => n22870);
   U5500 : NAND2_X1 port map( A1 => n3025, A2 => n1738, ZN => n24620);
   U5508 : INV_X1 port map( A => n24621, ZN => n24174);
   U5515 : OAI21_X1 port map( B1 => n16854, B2 => n368, A => n16852, ZN => 
                           n24621);
   U5530 : NAND2_X1 port map( A1 => n113, A2 => n20041, ZN => n19866);
   U5546 : NAND3_X1 port map( A1 => n10369, A2 => n10364, A3 => n24622, ZN => 
                           n24213);
   U5564 : NAND2_X1 port map( A1 => n897, A2 => n24623, ZN => n8368);
   U5565 : NAND3_X1 port map( A1 => n3110, A2 => n3111, A3 => n3109, ZN => 
                           n24623);
   U5623 : INV_X1 port map( A => n23883, ZN => n24624);
   U5642 : NAND2_X1 port map( A1 => n23879, A2 => n24624, ZN => n107);
   U5707 : OAI21_X1 port map( B1 => n3805, B2 => n22687, A => n3804, ZN => 
                           n24625);
   U5725 : NAND3_X1 port map( A1 => n24626, A2 => n23539, A3 => n23540, ZN => 
                           n23542);
   U5750 : NAND2_X1 port map( A1 => n23536, A2 => n24057, ZN => n24626);
   U5758 : AOI21_X1 port map( B1 => n23155, B2 => n22446, A => n24627, ZN => 
                           n22447);
   U5780 : NAND2_X1 port map( A1 => n10622, A2 => n11214, ZN => n24628);
   U5786 : NAND2_X1 port map( A1 => n2018, A2 => n2017, ZN => n2016);
   U5790 : MUX2_X1 port map( A => n23410, B => n23416, S => n23403, Z => n22866
                           );
   U5795 : NOR2_X1 port map( A1 => n22849, A2 => n22850, ZN => n23403);
   U5809 : NAND2_X1 port map( A1 => n24264, A2 => n24265, ZN => n24629);
   U5873 : XNOR2_X1 port map( A => n24630, B => n23816, ZN => Ciphertext(157));
   U5887 : NAND3_X1 port map( A1 => n536, A2 => n22541, A3 => n22540, ZN => 
                           n22543);
   U5915 : AOI21_X1 port map( B1 => n19980, B2 => n19983, A => n24315, ZN => 
                           n19985);
   U5954 : NAND3_X1 port map( A1 => n19819, A2 => n19820, A3 => n19818, ZN => 
                           n742);
   U6014 : NAND2_X1 port map( A1 => n24552, A2 => n12976, ZN => n12981);
   U6048 : NAND2_X1 port map( A1 => n24865, A2 => n2581, ZN => n24632);
   U6090 : NAND3_X1 port map( A1 => n776, A2 => n22125, A3 => n22421, ZN => 
                           n22126);
   U6139 : AOI21_X2 port map( B1 => n20895, B2 => n2364, A => n20894, ZN => 
                           n23647);
   U6166 : NAND3_X1 port map( A1 => n17252, A2 => n17279, A3 => n17273, ZN => 
                           n14748);
   U6171 : NAND3_X1 port map( A1 => n24571, A2 => n14510, A3 => n24713, ZN => 
                           n24712);
   U6191 : NAND2_X1 port map( A1 => n25383, A2 => n19573, ZN => n2018);
   U6252 : NAND2_X2 port map( A1 => n24633, A2 => n12857, ZN => n14321);
   U6310 : NAND3_X2 port map( A1 => n17291, A2 => n24196, A3 => n24635, ZN => 
                           n18512);
   U6322 : NAND3_X1 port map( A1 => n3539, A2 => n4424, A3 => n24636, ZN => 
                           n3538);
   U6325 : NAND2_X1 port map( A1 => n296, A2 => n14031, ZN => n24636);
   U6331 : NAND3_X1 port map( A1 => n23787, A2 => n2476, A3 => n21902, ZN => 
                           n2475);
   U6351 : NAND2_X1 port map( A1 => n24641, A2 => n24640, ZN => n24639);
   U6353 : NAND2_X1 port map( A1 => n12742, A2 => n12740, ZN => n24641);
   U6382 : NAND2_X1 port map( A1 => n12511, A2 => n12656, ZN => n24642);
   U6389 : XNOR2_X1 port map( A => n24643, B => n22195, ZN => Ciphertext(126));
   U6402 : NAND3_X1 port map( A1 => n22194, A2 => n22193, A3 => n22998, ZN => 
                           n24643);
   U6410 : NOR2_X1 port map( A1 => n24644, A2 => n25345, ZN => n98);
   U6411 : AND2_X1 port map( A1 => n17192, A2 => n4039, ZN => n24650);
   U6479 : NAND2_X1 port map( A1 => n19449, A2 => n25002, ZN => n24646);
   U6481 : NAND2_X1 port map( A1 => n19444, A2 => n19445, ZN => n24647);
   U6555 : BUF_X2 port map( A => n22593, Z => n24043);
   U6558 : AND2_X2 port map( A1 => n22595, A2 => n22594, ZN => n23040);
   U6559 : NAND2_X1 port map( A1 => n5018, A2 => n24650, ZN => n5017);
   U6570 : NAND2_X1 port map( A1 => n17196, A2 => n17031, ZN => n5018);
   U6598 : NAND2_X1 port map( A1 => n24595, A2 => n4536, ZN => n24652);
   U6607 : NAND2_X1 port map( A1 => n16159, A2 => n24653, ZN => n17395);
   U6623 : NAND3_X1 port map( A1 => n24656, A2 => n24655, A3 => n24654, ZN => 
                           n24653);
   U6638 : NAND2_X1 port map( A1 => n16154, A2 => n24458, ZN => n24654);
   U6663 : NAND2_X1 port map( A1 => n16122, A2 => n16124, ZN => n24656);
   U6690 : NAND2_X1 port map( A1 => n5152, A2 => n24657, ZN => n20961);
   U6715 : OAI21_X1 port map( B1 => n5155, B2 => n19576, A => n24658, ZN => 
                           n24657);
   U6717 : INV_X1 port map( A => n25072, ZN => n24658);
   U6737 : OAI211_X2 port map( C1 => n5391, C2 => n3760, A => n10379, B => 
                           n24659, ZN => n12151);
   U6760 : NAND2_X1 port map( A1 => n991, A2 => n416, ZN => n24659);
   U6771 : NAND2_X1 port map( A1 => n24660, A2 => n17081, ZN => n17480);
   U6788 : NAND2_X1 port map( A1 => n3908, A2 => n22329, ZN => n3907);
   U6810 : NAND3_X1 port map( A1 => n23139, A2 => n23131, A3 => n24473, ZN => 
                           n23132);
   U6825 : AND4_X2 port map( A1 => n24790, A2 => n3660, A3 => n3772, A4 => 
                           n3665, ZN => n20415);
   U6826 : NAND2_X1 port map( A1 => n7349, A2 => n7348, ZN => n7279);
   U6837 : XNOR2_X1 port map( A => n24661, B => n23137, ZN => Ciphertext(18));
   U6846 : NAND2_X1 port map( A1 => n23136, A2 => n23135, ZN => n24661);
   U6852 : XNOR2_X1 port map( A => n797, B => n24662, ZN => n18990);
   U6881 : NAND3_X1 port map( A1 => n3165, A2 => n17674, A3 => n5280, ZN => 
                           n17675);
   U6893 : NAND2_X1 port map( A1 => n24785, A2 => n14278, ZN => n24664);
   U6895 : OR2_X2 port map( A1 => n24665, A2 => n16811, ZN => n18418);
   U6900 : AOI22_X1 port map( A1 => n16807, A2 => n16896, B1 => n16806, B2 => 
                           n17078, ZN => n24665);
   U6901 : OR2_X1 port map( A1 => n4066, A2 => n20140, ZN => n5445);
   U6903 : AOI21_X2 port map( B1 => n4550, B2 => n19589, A => n4549, ZN => 
                           n20909);
   U6909 : NAND3_X1 port map( A1 => n4434, A2 => n23799, A3 => n23001, ZN => 
                           n23786);
   U6916 : NAND2_X1 port map( A1 => n22243, A2 => n24666, ZN => n2885);
   U6925 : XNOR2_X2 port map( A => n24667, B => n5369, ZN => n18959);
   U6929 : XNOR2_X1 port map( A => n17852, B => n18225, ZN => n24667);
   U6955 : NAND2_X2 port map( A1 => n1958, A2 => n1960, ZN => n7349);
   U7024 : NAND3_X1 port map( A1 => n9952, A2 => n9953, A3 => n9951, ZN => 
                           n9954);
   U7035 : INV_X1 port map( A => n7157, ZN => n7363);
   U7038 : NAND2_X1 port map( A1 => n7629, A2 => n7155, ZN => n7157);
   U7043 : NAND3_X1 port map( A1 => n21763, A2 => n24611, A3 => n24901, ZN => 
                           n21943);
   U7052 : NAND2_X1 port map( A1 => n10364, A2 => n10369, ZN => n2751);
   U7067 : NAND2_X1 port map( A1 => n19318, A2 => n4874, ZN => n17564);
   U7082 : NAND2_X1 port map( A1 => n13107, A2 => n13661, ZN => n24669);
   U7090 : NAND2_X1 port map( A1 => n24671, A2 => n24670, ZN => n13698);
   U7091 : NAND2_X1 port map( A1 => n13932, A2 => n14241, ZN => n24670);
   U7121 : NAND2_X1 port map( A1 => n13697, A2 => n4116, ZN => n24671);
   U7129 : NAND2_X1 port map( A1 => n13633, A2 => n13935, ZN => n13697);
   U7147 : AOI21_X1 port map( B1 => n22917, B2 => n22918, A => n22072, ZN => 
                           n24672);
   U7149 : NAND2_X1 port map( A1 => n24674, A2 => n21712, ZN => n24673);
   U7155 : OAI22_X1 port map( A1 => n25240, A2 => n24675, B1 => n24428, B2 => 
                           n24469, ZN => n22983);
   U7166 : INV_X1 port map( A => n23865, ZN => n24675);
   U7176 : NOR2_X2 port map( A1 => n12647, A2 => n24677, ZN => n14988);
   U7191 : NAND2_X1 port map( A1 => n3885, A2 => n3884, ZN => n24677);
   U7192 : AOI21_X2 port map( B1 => n13639, B2 => n13638, A => n24678, ZN => 
                           n14792);
   U7194 : NOR2_X1 port map( A1 => n13697, A2 => n24679, ZN => n24678);
   U7201 : OR2_X1 port map( A1 => n25247, A2 => n14053, ZN => n2756);
   U7206 : INV_X1 port map( A => n14553, ZN => n15200);
   U7230 : NOR2_X2 port map( A1 => n24680, A2 => n24602, ZN => n14553);
   U7252 : OAI21_X1 port map( B1 => n13204, B2 => n4116, A => n13202, ZN => 
                           n24680);
   U7259 : NAND2_X1 port map( A1 => n4407, A2 => n4406, ZN => n24270);
   U7262 : NAND2_X1 port map( A1 => n23392, A2 => n24465, ZN => n4412);
   U7273 : NAND2_X1 port map( A1 => n17401, A2 => n17402, ZN => n18484);
   U7276 : AOI22_X2 port map( A1 => n19828, A2 => n19827, B1 => n24682, B2 => 
                           n24681, ZN => n21561);
   U7280 : NOR2_X1 port map( A1 => n17016, A2 => n17208, ZN => n16257);
   U7295 : NAND3_X1 port map( A1 => n16253, A2 => n24684, A3 => n24683, ZN => 
                           n2093);
   U7301 : NAND2_X1 port map( A1 => n25389, A2 => n16016, ZN => n24683);
   U7307 : OR2_X1 port map( A1 => n16016, A2 => n16247, ZN => n24684);
   U7326 : NAND2_X1 port map( A1 => n15869, A2 => n17114, ZN => n24685);
   U7328 : NAND2_X1 port map( A1 => n19093, A2 => n18877, ZN => n24721);
   U7331 : NAND2_X1 port map( A1 => n24687, A2 => n24686, ZN => n2638);
   U7344 : NAND2_X1 port map( A1 => n15945, A2 => n16443, ZN => n24686);
   U7348 : NAND2_X1 port map( A1 => n15944, A2 => n16437, ZN => n24687);
   U7373 : NAND3_X1 port map( A1 => n25154, A2 => n24596, A3 => n7584, ZN => 
                           n1779);
   U7375 : NAND3_X1 port map( A1 => n10190, A2 => n10859, A3 => n10860, ZN => 
                           n10864);
   U7376 : NAND2_X1 port map( A1 => n24689, A2 => n25189, ZN => n9342);
   U7378 : NAND2_X1 port map( A1 => n25187, A2 => n25188, ZN => n24689);
   U7384 : NAND2_X1 port map( A1 => n7688, A2 => n7217, ZN => n7216);
   U7419 : NOR2_X2 port map( A1 => n18822, A2 => n18823, ZN => n20484);
   U7434 : OAI21_X1 port map( B1 => n3563, B2 => n14000, A => n24691, ZN => 
                           n13678);
   U7445 : XNOR2_X1 port map( A => n17969, B => n2137, ZN => n17927);
   U7458 : OAI21_X1 port map( B1 => n23886, B2 => n23885, A => n24692, ZN => 
                           n23887);
   U7479 : NAND3_X1 port map( A1 => n24765, A2 => n24610, A3 => n3713, ZN => 
                           n23285);
   U7525 : OAI21_X1 port map( B1 => n22982, B2 => n23860, A => n24694, ZN => 
                           n22985);
   U7570 : NAND3_X1 port map( A1 => n24675, A2 => n23857, A3 => n23862, ZN => 
                           n24694);
   U7633 : OR2_X1 port map( A1 => n13946, A2 => n13947, ZN => n24697);
   U7635 : AOI21_X2 port map( B1 => n24698, B2 => n3896, A => n21842, ZN => 
                           n23890);
   U7642 : INV_X1 port map( A => n10918, ZN => n1940);
   U7656 : OAI21_X1 port map( B1 => n16591, B2 => n17076, A => n16892, ZN => 
                           n24699);
   U7688 : NAND2_X1 port map( A1 => n974, A2 => n975, ZN => n976);
   U7696 : OR2_X1 port map( A1 => n19075, A2 => n19076, ZN => n24700);
   U7697 : OAI21_X2 port map( B1 => n13595, B2 => n14337, A => n24701, ZN => 
                           n15347);
   U7717 : OAI211_X1 port map( C1 => n23909, C2 => n23908, A => n24613, B => 
                           n24702, ZN => n23910);
   U7718 : NAND2_X1 port map( A1 => n23907, A2 => n23906, ZN => n24702);
   U7719 : NAND2_X1 port map( A1 => n24703, A2 => n24012, ZN => n24281);
   U7723 : OAI21_X1 port map( B1 => n23982, B2 => n24008, A => n23984, ZN => 
                           n24703);
   U7794 : OAI22_X1 port map( A1 => n20469, A2 => n5115, B1 => n5114, B2 => 
                           n20473, ZN => n24704);
   U7803 : AND2_X1 port map( A1 => n21847, A2 => n21816, ZN => n22353);
   U7842 : NAND3_X1 port map( A1 => n24706, A2 => n20418, A3 => n25108, ZN => 
                           n20420);
   U7845 : NAND2_X1 port map( A1 => n4509, A2 => n20401, ZN => n24706);
   U7846 : OAI21_X1 port map( B1 => n25022, B2 => n22667, A => n24707, ZN => 
                           n22787);
   U7851 : NAND2_X1 port map( A1 => n25022, A2 => n22782, ZN => n24707);
   U7854 : NAND3_X2 port map( A1 => n15713, A2 => n15711, A3 => n15712, ZN => 
                           n17299);
   U7855 : NAND2_X1 port map( A1 => n7044, A2 => n3730, ZN => n551);
   U7864 : OAI211_X2 port map( C1 => n10705, C2 => n2754, A => n10704, B => 
                           n24709, ZN => n1568);
   U7875 : NAND2_X1 port map( A1 => n10700, A2 => n10701, ZN => n24709);
   U7889 : NAND3_X1 port map( A1 => n24711, A2 => n14306, A3 => n24710, ZN => 
                           n24153);
   U7891 : INV_X1 port map( A => n24588, ZN => n24711);
   U7907 : NAND2_X1 port map( A1 => n24714, A2 => n24712, ZN => n13980);
   U7924 : NAND2_X1 port map( A1 => n5752, A2 => n24715, ZN => n24714);
   U7934 : INV_X1 port map( A => n14510, ZN => n24715);
   U7960 : NAND2_X1 port map( A1 => n5052, A2 => n16844, ZN => n16845);
   U7969 : NAND2_X1 port map( A1 => n19479, A2 => n19480, ZN => n24716);
   U7981 : NAND2_X1 port map( A1 => n16147, A2 => n16096, ZN => n16145);
   U7988 : NAND2_X1 port map( A1 => n19719, A2 => n24717, ZN => n18774);
   U8036 : NAND2_X1 port map( A1 => n24278, A2 => n24279, ZN => n22879);
   U8044 : NAND2_X1 port map( A1 => n20546, A2 => n20127, ZN => n19674);
   U8058 : NAND2_X1 port map( A1 => n16556, A2 => n16557, ZN => n4450);
   U8097 : NAND2_X1 port map( A1 => n23714, A2 => n23723, ZN => n23728);
   U8113 : OAI21_X2 port map( B1 => n22055, B2 => n22054, A => n22053, ZN => 
                           n23723);
   U8115 : AND2_X2 port map( A1 => n19209, A2 => n3106, ZN => n20576);
   U8124 : NAND2_X1 port map( A1 => n25382, A2 => n24718, ZN => n22846);
   U8213 : NOR2_X1 port map( A1 => n24720, A2 => n17449, ZN => n17150);
   U8220 : NAND3_X1 port map( A1 => n6077, A2 => n6076, A3 => n6883, ZN => 
                           n2786);
   U8229 : NOR2_X1 port map( A1 => n17148, A2 => n17455, ZN => n24720);
   U8240 : NAND2_X1 port map( A1 => n4730, A2 => n4731, ZN => n10753);
   U8248 : NAND2_X1 port map( A1 => n24721, A2 => n24335, ZN => n18879);
   U8268 : NAND2_X1 port map( A1 => n20131, A2 => n20522, ZN => n19971);
   U8284 : NOR2_X1 port map( A1 => n22849, A2 => n22850, ZN => n25035);
   U8285 : OAI21_X1 port map( B1 => n22848, B2 => n22847, A => n22846, ZN => 
                           n22849);
   U8306 : NAND2_X1 port map( A1 => n20066, A2 => n20071, ZN => n24722);
   U8310 : NAND2_X1 port map( A1 => n5759, A2 => n16676, ZN => n16678);
   U8313 : NOR2_X1 port map( A1 => n16824, A2 => n16862, ZN => n807);
   U8314 : NOR2_X1 port map( A1 => n282, A2 => n16112, ZN => n16862);
   U8331 : AND2_X2 port map( A1 => n24723, A2 => n5997, ZN => n7609);
   U8339 : NAND2_X1 port map( A1 => n3167, A2 => n5996, ZN => n24723);
   U8343 : NAND2_X1 port map( A1 => n1978, A2 => n1977, ZN => n19875);
   U8350 : OR2_X1 port map( A1 => n10884, A2 => n10885, ZN => n24167);
   U8356 : XNOR2_X2 port map( A => n21698, B => n21697, ZN => n22904);
   U8357 : NAND3_X2 port map( A1 => n24269, A2 => n4572, A3 => n4573, ZN => 
                           n18261);
   U8369 : NAND2_X1 port map( A1 => n2660, A2 => n2708, ZN => n2710);
   U8372 : NAND2_X1 port map( A1 => n24725, A2 => n642, ZN => n12465);
   U8375 : NAND2_X1 port map( A1 => n401, A2 => n12533, ZN => n24725);
   U8376 : NAND2_X1 port map( A1 => n3046, A2 => n20211, ZN => n3045);
   U8395 : NAND2_X1 port map( A1 => n24726, A2 => n18299, ZN => n1716);
   U8418 : NAND2_X1 port map( A1 => n3752, A2 => n3751, ZN => n24726);
   U8427 : NAND2_X1 port map( A1 => n9468, A2 => n1595, ZN => n3291);
   U8440 : NAND2_X1 port map( A1 => n24442, A2 => n23481, ZN => n2997);
   U8446 : NAND2_X1 port map( A1 => n2168, A2 => n20478, ZN => n20356);
   U8454 : AND3_X2 port map( A1 => n4768, A2 => n4769, A3 => n4770, ZN => 
                           n14789);
   U8455 : OAI21_X1 port map( B1 => n24172, B2 => n19464, A => n24727, ZN => 
                           n19462);
   U8459 : NAND2_X1 port map( A1 => n19464, A2 => n19457, ZN => n24727);
   U8465 : XNOR2_X1 port map( A => n18494, B => n24728, ZN => n25072);
   U8469 : NOR2_X1 port map( A1 => n22889, A2 => n22093, ZN => n24729);
   U8477 : NAND2_X1 port map( A1 => n20136, A2 => n20134, ZN => n20016);
   U8483 : NAND2_X1 port map( A1 => n25248, A2 => n13303, ZN => n3847);
   U8487 : NAND3_X1 port map( A1 => n4714, A2 => n5428, A3 => n24730, ZN => 
                           n17592);
   U8493 : NAND3_X1 port map( A1 => n16572, A2 => n17115, A3 => n890, ZN => 
                           n24730);
   U8542 : XOR2_X1 port map( A => n24383, B => n924, Z => n24769);
   U8567 : NAND2_X1 port map( A1 => n1355, A2 => n14048, ZN => n14053);
   U8577 : NAND2_X1 port map( A1 => n14141, A2 => n14189, ZN => n14188);
   U8578 : NAND3_X1 port map( A1 => n291, A2 => n24098, A3 => n16043, ZN => 
                           n1897);
   U8580 : NAND2_X1 port map( A1 => n10399, A2 => n10659, ZN => n10315);
   U8583 : BUF_X1 port map( A => n20036, Z => n22056);
   U8600 : AOI21_X1 port map( B1 => n2253, B2 => n15789, A => n24098, ZN => 
                           n15536);
   U8618 : NAND2_X1 port map( A1 => n16706, A2 => n16705, ZN => n16707);
   U8632 : NAND2_X1 port map( A1 => n20242, A2 => n19937, ZN => n19821);
   U8648 : AOI21_X2 port map( B1 => n19338, B2 => n19337, A => n19336, ZN => 
                           n20242);
   U8663 : NAND2_X1 port map( A1 => n548, A2 => n549, ZN => n24733);
   U8687 : NAND2_X1 port map( A1 => n24184, A2 => n22052, ZN => n22053);
   U8695 : NAND2_X1 port map( A1 => n24734, A2 => n14305, ZN => n15275);
   U8726 : NOR2_X1 port map( A1 => n1526, A2 => n1450, ZN => n24734);
   U8729 : NAND2_X1 port map( A1 => n24735, A2 => n11174, ZN => n11179);
   U8731 : NAND2_X1 port map( A1 => n11170, A2 => n24736, ZN => n24735);
   U8774 : INV_X1 port map( A => n11168, ZN => n24736);
   U8776 : XNOR2_X1 port map( A => n24737, B => n11924, ZN => n861);
   U8803 : XNOR2_X1 port map( A => n11923, B => n11922, ZN => n24737);
   U8816 : NAND2_X1 port map( A1 => n4514, A2 => n1619, ZN => n4513);
   U8870 : OAI21_X1 port map( B1 => n20069, B2 => n20072, A => n24738, ZN => 
                           n19854);
   U8882 : NAND3_X1 port map( A1 => n19852, A2 => n19660, A3 => n20068, ZN => 
                           n24738);
   U8915 : INV_X1 port map( A => n10103, ZN => n24740);
   U8918 : NAND2_X1 port map( A1 => n524, A2 => n354, ZN => n1132);
   U8930 : NAND2_X1 port map( A1 => n15621, A2 => n24537, ZN => n24741);
   U8932 : NAND2_X1 port map( A1 => n19091, A2 => n19904, ZN => n2916);
   U8960 : NAND2_X2 port map( A1 => n12714, A2 => n24742, ZN => n14439);
   U8967 : OAI21_X1 port map( B1 => n12708, B2 => n12709, A => n13078, ZN => 
                           n24742);
   U8968 : NAND2_X1 port map( A1 => n24743, A2 => n16497, ZN => n17581);
   U8969 : OAI21_X1 port map( B1 => n16487, B2 => n16488, A => n368, ZN => 
                           n24743);
   U8984 : NAND2_X1 port map( A1 => n24746, A2 => n24744, ZN => n5330);
   U8988 : NAND2_X1 port map( A1 => n13785, A2 => n14190, ZN => n24745);
   U8989 : NAND2_X1 port map( A1 => n13787, A2 => n24347, ZN => n24746);
   U8992 : NAND2_X1 port map( A1 => n4946, A2 => n12539, ZN => n12984);
   U9012 : NAND2_X1 port map( A1 => n16138, A2 => n24747, ZN => n18195);
   U9018 : NAND2_X1 port map( A1 => n16780, A2 => n25256, ZN => n24747);
   U9028 : AOI21_X1 port map( B1 => n20328, B2 => n20329, A => n24749, ZN => 
                           n20334);
   U9032 : NAND2_X1 port map( A1 => n11328, A2 => n12791, ZN => n12793);
   U9037 : NAND2_X1 port map( A1 => n2883, A2 => n3257, ZN => n8506);
   U9041 : AOI22_X1 port map( A1 => n17449, A2 => n16980, B1 => n16979, B2 => 
                           n17455, ZN => n16369);
   U9076 : NAND2_X1 port map( A1 => n24751, A2 => n1806, ZN => n2198);
   U9080 : OAI21_X1 port map( B1 => n19239, B2 => n24606, A => n19614, ZN => 
                           n24751);
   U9094 : NAND2_X1 port map( A1 => n7002, A2 => n7003, ZN => n4150);
   U9097 : NAND2_X1 port map( A1 => n3860, A2 => n4788, ZN => n14059);
   U9098 : NAND2_X1 port map( A1 => n24752, A2 => n5379, ZN => n5382);
   U9099 : NAND3_X1 port map( A1 => n4281, A2 => n4143, A3 => n24753, ZN => 
                           n24752);
   U9113 : XNOR2_X1 port map( A => n24754, B => n21553, ZN => n18045);
   U9133 : NAND3_X1 port map( A1 => n2790, A2 => n16259, A3 => n2789, ZN => 
                           n24754);
   U9148 : NAND2_X2 port map( A1 => n24755, A2 => n13492, ZN => n15514);
   U9152 : NAND2_X1 port map( A1 => n24815, A2 => n25036, ZN => n24755);
   U9164 : NAND3_X1 port map( A1 => n18385, A2 => n24757, A3 => n24756, ZN => 
                           n4792);
   U9195 : NAND2_X1 port map( A1 => n25195, A2 => n19176, ZN => n24756);
   U9196 : NAND2_X1 port map( A1 => n19177, A2 => n18777, ZN => n24757);
   U9203 : INV_X1 port map( A => n19183, ZN => n24758);
   U9204 : NAND2_X1 port map( A1 => n19297, A2 => n19296, ZN => n24759);
   U9208 : XNOR2_X1 port map( A => n15238, B => n1362, ZN => n14867);
   U9211 : NOR2_X2 port map( A1 => n14323, A2 => n654, ZN => n15238);
   U9217 : NAND2_X1 port map( A1 => n17296, A2 => n1535, ZN => n17300);
   U9219 : NAND2_X1 port map( A1 => n24855, A2 => n15704, ZN => n1535);
   U9257 : NAND3_X1 port map( A1 => n6261, A2 => n6259, A3 => n6260, ZN => 
                           n6263);
   U9264 : NAND2_X1 port map( A1 => n24764, A2 => n24763, ZN => n15740);
   U9268 : NAND3_X1 port map( A1 => n2587, A2 => n16795, A3 => n16550, ZN => 
                           n24763);
   U9336 : NAND2_X1 port map( A1 => n15739, A2 => n4554, ZN => n24764);
   U9341 : NAND2_X1 port map( A1 => n22424, A2 => n22945, ZN => n24765);
   U9384 : NAND2_X1 port map( A1 => n9661, A2 => n422, ZN => n24767);
   U9385 : OR3_X1 port map( A1 => n13234, A2 => n12902, A3 => n12935, ZN => 
                           n2545);
   U9402 : OAI21_X2 port map( B1 => n16586, B2 => n16587, A => n16585, ZN => 
                           n18042);
   U9417 : NAND3_X1 port map( A1 => n21767, A2 => n25018, A3 => n22156, ZN => 
                           n24768);
   U9424 : NAND2_X1 port map( A1 => n22270, A2 => n22453, ZN => n22451);
   U9471 : NAND2_X1 port map( A1 => n2806, A2 => n2004, ZN => n2175);
   U9490 : NAND2_X1 port map( A1 => n98, A2 => n101, ZN => n1995);
   U9509 : NAND3_X1 port map( A1 => n24770, A2 => n17253, A3 => n17250, ZN => 
                           n720);
   U9513 : NAND2_X1 port map( A1 => n17247, A2 => n17248, ZN => n24770);
   U9536 : NOR2_X1 port map( A1 => n13265, A2 => n13267, ZN => n24805);
   U9567 : NAND3_X1 port map( A1 => n647, A2 => n4076, A3 => n17942, ZN => 
                           n24217);
   U9595 : OAI211_X1 port map( C1 => n7752, C2 => n2640, A => n7751, B => 
                           n24771, ZN => n7753);
   U9624 : NAND2_X1 port map( A1 => n8014, A2 => n7749, ZN => n24771);
   U9627 : NAND2_X1 port map( A1 => n24801, A2 => n24603, ZN => n17249);
   U9644 : NAND2_X1 port map( A1 => n7341, A2 => n7602, ZN => n7596);
   U9670 : NAND3_X1 port map( A1 => n6459, A2 => n6456, A3 => n6454, ZN => 
                           n6032);
   U9676 : XNOR2_X2 port map( A => n14491, B => n14492, ZN => n15611);
   U9678 : NAND3_X1 port map( A1 => n13743, A2 => n13744, A3 => n24773, ZN => 
                           n2071);
   U9682 : NAND2_X1 port map( A1 => n15726, A2 => n24774, ZN => n15727);
   U9708 : INV_X1 port map( A => n19446, ZN => n17711);
   U9720 : NAND2_X1 port map( A1 => n19645, A2 => n20027, ZN => n19649);
   U9725 : NAND2_X1 port map( A1 => n10137, A2 => n10138, ZN => n9174);
   U9726 : NAND3_X1 port map( A1 => n6812, A2 => n6367, A3 => n6815, ZN => 
                           n6813);
   U9731 : NAND2_X1 port map( A1 => n6367, A2 => n6368, ZN => n6812);
   U9739 : NAND2_X1 port map( A1 => n17230, A2 => n24775, ZN => n14588);
   U9740 : NAND2_X1 port map( A1 => n22947, A2 => n2674, ZN => n22125);
   U9751 : NAND2_X1 port map( A1 => n10584, A2 => n10583, ZN => n10370);
   U9752 : INV_X1 port map( A => n9460, ZN => n24844);
   U9756 : NAND2_X1 port map( A1 => n16299, A2 => n24506, ZN => n24777);
   U9758 : NAND3_X1 port map( A1 => n17186, A2 => n17025, A3 => n3602, ZN => 
                           n16213);
   U9774 : NAND2_X1 port map( A1 => n22888, A2 => n22887, ZN => n22727);
   U9790 : INV_X1 port map( A => n11622, ZN => n12335);
   U9793 : XNOR2_X1 port map( A => n11622, B => n24778, ZN => n11181);
   U9797 : NOR2_X2 port map( A1 => n10340, A2 => n10339, ZN => n11622);
   U9799 : NAND2_X1 port map( A1 => n24779, A2 => n6986, ZN => n5636);
   U9801 : NAND2_X1 port map( A1 => n2646, A2 => n6639, ZN => n24779);
   U9805 : XNOR2_X1 port map( A => n17806, B => n20046, ZN => n17619);
   U9806 : OAI22_X2 port map( A1 => n4414, A2 => n4413, B1 => n17176, B2 => 
                           n17177, ZN => n17806);
   U9815 : XNOR2_X1 port map( A => n24780, B => n23825, ZN => Ciphertext(159));
   U9831 : OAI211_X1 port map( C1 => n23823, C2 => n23824, A => n23822, B => 
                           n23821, ZN => n24780);
   U9832 : AND2_X2 port map( A1 => n24782, A2 => n24781, ZN => n23650);
   U9869 : OAI211_X2 port map( C1 => n16568, C2 => n17227, A => n16566, B => 
                           n24783, ZN => n18530);
   U9883 : NAND3_X1 port map( A1 => n16565, A2 => n17225, A3 => n17224, ZN => 
                           n24783);
   U9893 : NAND2_X1 port map( A1 => n939, A2 => n11032, ZN => n3467);
   U9918 : NAND3_X1 port map( A1 => n13975, A2 => n14439, A3 => n24571, ZN => 
                           n14434);
   U9919 : NAND3_X1 port map( A1 => n24784, A2 => n8512, A3 => n24224, ZN => 
                           n24851);
   U9928 : NAND2_X1 port map( A1 => n1279, A2 => n8511, ZN => n24784);
   U9976 : NAND2_X1 port map( A1 => n1108, A2 => n19786, ZN => n3214);
   U9982 : NAND2_X1 port map( A1 => n19986, A2 => n19784, ZN => n19786);
   U9989 : INV_X1 port map( A => n21352, ZN => n21363);
   U10000 : INV_X1 port map( A => n14278, ZN => n4767);
   U10004 : NAND3_X2 port map( A1 => n5156, A2 => n1970, A3 => n12609, ZN => 
                           n14278);
   U10005 : NAND3_X1 port map( A1 => n23947, A2 => n24910, A3 => n23952, ZN => 
                           n463);
   U10012 : XNOR2_X2 port map( A => n8678, B => n8679, ZN => n9981);
   U10025 : NAND2_X1 port map( A1 => n21390, A2 => n21389, ZN => n23155);
   U10056 : NAND2_X1 port map( A1 => n23065, A2 => n23066, ZN => n22872);
   U10059 : NAND2_X1 port map( A1 => n14198, A2 => n3888, ZN => n13804);
   U10063 : NAND2_X2 port map( A1 => n5402, A2 => n12631, ZN => n3888);
   U10070 : OR2_X1 port map( A1 => n18979, A2 => n19456, ZN => n19031);
   U10072 : NAND2_X1 port map( A1 => n14708, A2 => n24928, ZN => n16686);
   U10075 : OR2_X1 port map( A1 => n19097, A2 => n2216, ZN => n18726);
   U10079 : NAND2_X1 port map( A1 => n2643, A2 => n18865, ZN => n19236);
   U10082 : NAND2_X1 port map( A1 => n15859, A2 => n16120, ZN => n24786);
   U10097 : NAND2_X1 port map( A1 => n15858, A2 => n15857, ZN => n24787);
   U10098 : INV_X1 port map( A => n24864, ZN => n24788);
   U10110 : NAND2_X1 port map( A1 => n13526, A2 => n13466, ZN => n3331);
   U10133 : XNOR2_X1 port map( A => n24789, B => n4761, ZN => Ciphertext(7));
   U10224 : NAND3_X1 port map( A1 => n1210, A2 => n24087, A3 => n10148, ZN => 
                           n2732);
   U10225 : NAND3_X1 port map( A1 => n21361, A2 => n318, A3 => n23828, ZN => 
                           n1934);
   U10253 : NAND2_X1 port map( A1 => n2396, A2 => n22313, ZN => n22314);
   U10270 : NAND2_X1 port map( A1 => n279, A2 => n19541, ZN => n24790);
   U10286 : OAI211_X1 port map( C1 => n3868, C2 => n11214, A => n233, B => 
                           n24791, ZN => n543);
   U10289 : NAND2_X1 port map( A1 => n11214, A2 => n11215, ZN => n24791);
   U10296 : NAND2_X1 port map( A1 => n1340, A2 => n23219, ZN => n23222);
   U10327 : NAND2_X1 port map( A1 => n20785, A2 => n20786, ZN => n23219);
   U10333 : NAND2_X1 port map( A1 => n9943, A2 => n9945, ZN => n9287);
   U10347 : XNOR2_X2 port map( A => n8123, B => n8122, ZN => n9945);
   U10404 : NAND2_X1 port map( A1 => n18951, A2 => n3215, ZN => n19784);
   U10405 : NAND3_X1 port map( A1 => n17762, A2 => n24477, A3 => n19389, ZN => 
                           n17763);
   U10433 : XNOR2_X1 port map( A => n24794, B => n1854, ZN => Ciphertext(56));
   U10448 : NOR2_X2 port map( A1 => n17765, A2 => n17766, ZN => n20109);
   U10449 : NAND2_X1 port map( A1 => n16769, A2 => n24569, ZN => n24863);
   U10451 : NAND2_X1 port map( A1 => n22969, A2 => n22968, ZN => n22416);
   U10462 : NAND2_X1 port map( A1 => n25120, A2 => n25119, ZN => n24795);
   U10533 : OAI211_X1 port map( C1 => n16120, C2 => n15611, A => n24797, B => 
                           n24796, ZN => n5178);
   U10573 : NAND2_X1 port map( A1 => n16120, A2 => n16118, ZN => n24796);
   U10576 : NAND3_X1 port map( A1 => n366, A2 => n2566, A3 => n24798, ZN => 
                           n1035);
   U10577 : NAND2_X1 port map( A1 => n4284, A2 => n4285, ZN => n24798);
   U10582 : NAND2_X1 port map( A1 => n24800, A2 => n24799, ZN => n11892);
   U10590 : NAND2_X1 port map( A1 => n10479, A2 => n10628, ZN => n24800);
   U10602 : INV_X1 port map( A => n9990, ZN => n25121);
   U10612 : MUX2_X1 port map( A => n19132, B => n19304, S => n19133, Z => 
                           n16504);
   U10623 : NAND2_X1 port map( A1 => n2733, A2 => n7324, ZN => n1254);
   U10631 : NAND2_X1 port map( A1 => n14745, A2 => n14744, ZN => n24801);
   U10642 : OAI21_X1 port map( B1 => n19476, B2 => n24803, A => n24802, ZN => 
                           n19483);
   U10668 : NAND2_X1 port map( A1 => n19476, A2 => n18734, ZN => n24802);
   U10710 : NAND2_X1 port map( A1 => n19641, A2 => n5115, ZN => n19642);
   U10735 : NAND3_X1 port map( A1 => n3974, A2 => n10360, A3 => n12506, ZN => 
                           n3633);
   U10766 : OAI21_X1 port map( B1 => n25183, B2 => n20846, A => n1156, ZN => 
                           n23619);
   U10807 : NAND2_X1 port map( A1 => n12832, A2 => n24805, ZN => n5645);
   U10826 : NAND2_X1 port map( A1 => n4066, A2 => n20140, ZN => n4615);
   U10845 : NAND2_X2 port map( A1 => n4245, A2 => n4067, ZN => n4066);
   U10863 : NAND2_X1 port map( A1 => n13336, A2 => n231, ZN => n12839);
   U10909 : XNOR2_X2 port map( A => n10299, B => n10300, ZN => n12506);
   U10930 : XNOR2_X1 port map( A => n12303, B => n12269, ZN => n10300);
   U10936 : NAND2_X1 port map( A1 => n17284, A2 => n17288, ZN => n16753);
   U10945 : OAI21_X1 port map( B1 => n17124, B2 => n17123, A => n24806, ZN => 
                           n4661);
   U10960 : INV_X1 port map( A => n17824, ZN => n24806);
   U10963 : OAI211_X1 port map( C1 => n19352, C2 => n24809, A => n19451, B => 
                           n24808, ZN => n24807);
   U10984 : NAND2_X1 port map( A1 => n19352, A2 => n19357, ZN => n24808);
   U10986 : NOR2_X1 port map( A1 => n6068, A2 => n24810, ZN => n7278);
   U11013 : NAND3_X1 port map( A1 => n9660, A2 => n9659, A3 => n9745, ZN => 
                           n1943);
   U11021 : NAND2_X1 port map( A1 => n3737, A2 => n23851, ZN => n3739);
   U11022 : NAND2_X1 port map( A1 => n1566, A2 => n24811, ZN => n25107);
   U11027 : NAND2_X1 port map( A1 => n12612, A2 => n25248, ZN => n24811);
   U11068 : NAND2_X1 port map( A1 => n23328, A2 => n23329, ZN => n23331);
   U11115 : NAND2_X1 port map( A1 => n1261, A2 => n15612, ZN => n15861);
   U11128 : AND2_X1 port map( A1 => n1147, A2 => n6690, ZN => n1148);
   U11146 : OR2_X1 port map( A1 => n13028, A2 => n302, ZN => n2794);
   U11162 : NAND2_X1 port map( A1 => n4445, A2 => n11974, ZN => n24812);
   U11170 : NAND2_X1 port map( A1 => n19478, A2 => n4667, ZN => n17594);
   U11171 : XNOR2_X2 port map( A => n10, B => n17591, ZN => n19478);
   U11184 : OAI211_X2 port map( C1 => n16982, C2 => n16983, A => n16981, B => 
                           n3982, ZN => n18172);
   U11185 : NAND2_X1 port map( A1 => n24813, A2 => n17551, ZN => n17552);
   U11188 : OAI21_X1 port map( B1 => n18927, B2 => n18967, A => n356, ZN => 
                           n24813);
   U11198 : NAND2_X1 port map( A1 => n24169, A2 => n24171, ZN => n3122);
   U11205 : NAND2_X1 port map( A1 => n1689, A2 => n5101, ZN => n2967);
   U11208 : NAND2_X1 port map( A1 => n9231, A2 => n25457, ZN => n5688);
   U11209 : NAND2_X1 port map( A1 => n25103, A2 => n11065, ZN => n11075);
   U11215 : XNOR2_X1 port map( A => n9143, B => n24600, ZN => n1466);
   U11240 : NAND2_X1 port map( A1 => n20320, A2 => n20322, ZN => n18992);
   U11250 : OAI21_X1 port map( B1 => n10633, B2 => n11210, A => n24814, ZN => 
                           n4089);
   U11257 : NAND3_X1 port map( A1 => n11210, A2 => n11338, A3 => n24082, ZN => 
                           n24814);
   U11299 : NAND2_X1 port map( A1 => n24495, A2 => n8839, ZN => n10015);
   U11314 : NAND3_X2 port map( A1 => n4650, A2 => n13464, A3 => n13465, ZN => 
                           n14468);
   U11351 : OR2_X1 port map( A1 => n15705, A2 => n16464, ZN => n24855);
   U11352 : NAND3_X2 port map( A1 => n24817, A2 => n24816, A3 => n9509, ZN => 
                           n11396);
   U11353 : NAND3_X1 port map( A1 => n4142, A2 => n5380, A3 => n11032, ZN => 
                           n24816);
   U11376 : OAI21_X1 port map( B1 => n20243, B2 => n20244, A => n20242, ZN => 
                           n24818);
   U11385 : NAND3_X2 port map( A1 => n24819, A2 => n1113, A3 => n1114, ZN => 
                           n17086);
   U11411 : NAND2_X1 port map( A1 => n24821, A2 => n24820, ZN => n24819);
   U11462 : NAND2_X1 port map( A1 => n16469, A2 => n24551, ZN => n24820);
   U11481 : AOI21_X1 port map( B1 => n15546, B2 => n24822, A => n383, ZN => 
                           n24821);
   U11491 : NAND3_X2 port map( A1 => n9728, A2 => n24824, A3 => n24823, ZN => 
                           n11158);
   U11495 : NAND2_X1 port map( A1 => n9726, A2 => n2922, ZN => n24823);
   U11506 : NAND2_X1 port map( A1 => n9725, A2 => n25043, ZN => n24824);
   U11516 : NAND2_X1 port map( A1 => n24826, A2 => n1365, ZN => n24825);
   U11518 : XNOR2_X2 port map( A => n14632, B => n14633, ZN => n1365);
   U11529 : INV_X1 port map( A => n16073, ZN => n24826);
   U11549 : OAI22_X2 port map( A1 => n279, A2 => n19544, B1 => n19543, B2 => 
                           n19545, ZN => n20368);
   U11557 : OAI21_X1 port map( B1 => n5709, B2 => n13581, A => n14107, ZN => 
                           n24827);
   U11567 : OAI21_X1 port map( B1 => n25388, B2 => n24829, A => n24828, ZN => 
                           n19717);
   U11568 : NAND2_X1 port map( A1 => n25388, A2 => n339, ZN => n24828);
   U11587 : NAND2_X1 port map( A1 => n14150, A2 => n3717, ZN => n14154);
   U11589 : NAND3_X2 port map( A1 => n4860, A2 => n24258, A3 => n4964, ZN => 
                           n3717);
   U11593 : NAND2_X1 port map( A1 => n25480, A2 => n6480, ZN => n6926);
   U11617 : NOR2_X1 port map( A1 => n19850, A2 => n19660, ZN => n20066);
   U11665 : NAND2_X1 port map( A1 => n13188, A2 => n13187, ZN => n13189);
   U11672 : XNOR2_X1 port map( A => n24830, B => n23931, ZN => Ciphertext(177))
                           ;
   U11685 : NAND3_X1 port map( A1 => n24831, A2 => n23928, A3 => n23929, ZN => 
                           n24830);
   U11730 : NAND2_X1 port map( A1 => n24833, A2 => n4309, ZN => n22507);
   U11754 : OAI21_X1 port map( B1 => n4311, B2 => n5306, A => n23425, ZN => 
                           n24833);
   U11757 : NAND2_X1 port map( A1 => n24834, A2 => n20616, ZN => n20326);
   U11779 : NAND2_X1 port map( A1 => n20084, A2 => n24835, ZN => n24834);
   U11783 : NAND2_X1 port map( A1 => n20571, A2 => n20614, ZN => n20084);
   U11795 : NOR2_X2 port map( A1 => n4577, A2 => n24836, ZN => n11385);
   U11821 : AOI21_X1 port map( B1 => n9580, B2 => n9581, A => n11116, ZN => 
                           n24836);
   U11822 : NAND2_X1 port map( A1 => n513, A2 => n19662, ZN => n2339);
   U11826 : NAND2_X1 port map( A1 => n23469, A2 => n23499, ZN => n23474);
   U11828 : NAND2_X1 port map( A1 => n24837, A2 => n2713, ZN => n22026);
   U11833 : NAND2_X1 port map( A1 => n22019, A2 => n25438, ZN => n24837);
   U11838 : OAI21_X1 port map( B1 => n324, B2 => n4411, A => n24838, ZN => 
                           n4407);
   U11841 : NAND2_X1 port map( A1 => n4412, A2 => n324, ZN => n24838);
   U11853 : AND3_X2 port map( A1 => n5240, A2 => n5241, A3 => n16797, ZN => 
                           n16799);
   U11868 : NAND2_X1 port map( A1 => n20269, A2 => n1155, ZN => n1154);
   U11871 : OAI211_X1 port map( C1 => n9503, C2 => n10104, A => n24839, B => 
                           n8644, ZN => n9332);
   U11874 : NAND2_X1 port map( A1 => n9503, A2 => n9775, ZN => n24839);
   U11938 : INV_X1 port map( A => n16290, ZN => n24841);
   U11959 : NAND2_X1 port map( A1 => n9920, A2 => n9461, ZN => n24843);
   U11979 : OAI211_X2 port map( C1 => n20098, C2 => n20566, A => n24109, B => 
                           n24845, ZN => n21520);
   U12001 : NAND3_X1 port map( A1 => n24846, A2 => n3914, A3 => n3912, ZN => 
                           n24112);
   U12005 : NAND3_X1 port map( A1 => n3910, A2 => n3909, A3 => n23058, ZN => 
                           n24846);
   U12007 : INV_X1 port map( A => n9921, ZN => n24847);
   U12021 : OR2_X1 port map( A1 => n9922, A2 => n9920, ZN => n24848);
   U12024 : OAI21_X1 port map( B1 => n16063, B2 => n16064, A => n24849, ZN => 
                           n15602);
   U12028 : NAND2_X1 port map( A1 => n16064, A2 => n25446, ZN => n24849);
   U12033 : OAI211_X2 port map( C1 => n7107, C2 => n7250, A => n24851, B => 
                           n7106, ZN => n8280);
   U12051 : NAND2_X1 port map( A1 => n25211, A2 => n20042, ZN => n19230);
   U12083 : NOR2_X1 port map( A1 => n5800, A2 => n6964, ZN => n6672);
   U12099 : OAI211_X1 port map( C1 => n9919, C2 => n9354, A => n24852, B => 
                           n9355, ZN => n9357);
   U12100 : NAND2_X1 port map( A1 => n9919, A2 => n24853, ZN => n24852);
   U12108 : OAI21_X1 port map( B1 => n10199, B2 => n10200, A => n13092, ZN => 
                           n24854);
   U12129 : NAND2_X1 port map( A1 => n10694, A2 => n11499, ZN => n10331);
   U12147 : NAND2_X1 port map( A1 => n23905, A2 => n21863, ZN => n607);
   U12170 : NAND2_X1 port map( A1 => n14000, A2 => n12668, ZN => n14002);
   U12276 : NAND3_X1 port map( A1 => n244, A2 => n707, A3 => n16427, ZN => 
                           n17435);
   U12277 : NAND2_X1 port map( A1 => n11211, A2 => n11342, ZN => n24856);
   U12280 : NAND2_X1 port map( A1 => n2071, A2 => n24857, ZN => n14800);
   U12465 : NAND2_X1 port map( A1 => n13734, A2 => n4979, ZN => n24857);
   U12492 : NOR2_X2 port map( A1 => n24858, A2 => n13980, ZN => n15088);
   U12512 : OAI22_X1 port map( A1 => n13977, A2 => n14439, B1 => n13978, B2 => 
                           n24713, ZN => n24858);
   U12535 : OAI21_X1 port map( B1 => n10020, B2 => n9730, A => n24859, ZN => 
                           n5372);
   U12541 : NAND2_X1 port map( A1 => n9491, A2 => n10019, ZN => n24859);
   U12546 : NOR2_X1 port map( A1 => n16183, A2 => n25455, ZN => n15916);
   U12601 : NAND2_X1 port map( A1 => n15915, A2 => n15667, ZN => n16183);
   U12636 : OAI21_X1 port map( B1 => n7897, B2 => n24861, A => n24860, ZN => 
                           n7903);
   U12684 : NAND2_X1 port map( A1 => n7897, A2 => n7898, ZN => n24860);
   U12701 : NAND3_X1 port map( A1 => n22812, A2 => n22656, A3 => n22813, ZN => 
                           n2527);
   U12739 : NAND2_X1 port map( A1 => n6394, A2 => n4178, ZN => n4177);
   U12770 : NAND2_X1 port map( A1 => n24862, A2 => n24354, ZN => n2685);
   U12773 : INV_X1 port map( A => n20452, ZN => n24862);
   U12807 : NAND2_X1 port map( A1 => n1590, A2 => n20451, ZN => n20452);
   U12808 : NAND3_X2 port map( A1 => n3416, A2 => n3417, A3 => n3415, ZN => 
                           n12306);
   U12831 : AOI21_X1 port map( B1 => n15860, B2 => n15861, A => n16113, ZN => 
                           n24864);
   U12847 : NAND2_X1 port map( A1 => n9936, A2 => n2971, ZN => n2947);
   U12900 : NOR2_X1 port map( A1 => n16572, A2 => n2580, ZN => n24865);
   U12983 : OAI21_X1 port map( B1 => n20669, B2 => n24567, A => n24866, ZN => 
                           n17311);
   U12994 : NAND2_X1 port map( A1 => n20669, A2 => n20335, ZN => n24866);
   U13004 : NAND2_X1 port map( A1 => n24868, A2 => n24867, ZN => n24019);
   U13144 : NAND2_X1 port map( A1 => n22776, A2 => n22677, ZN => n24867);
   U13167 : NAND2_X1 port map( A1 => n22777, A2 => n24869, ZN => n24868);
   U13168 : NAND2_X1 port map( A1 => n2618, A2 => n2617, ZN => n22777);
   U13170 : NAND2_X1 port map( A1 => n10491, A2 => n11207, ZN => n1225);
   U13184 : OAI21_X1 port map( B1 => n20586, B2 => n3734, A => n24870, ZN => 
                           n5094);
   U13185 : NAND2_X1 port map( A1 => n20586, A2 => n20593, ZN => n24870);
   U13191 : XNOR2_X1 port map( A => n10719, B => n24871, ZN => n10745);
   U13192 : XNOR2_X1 port map( A => n24969, B => n11295, ZN => n24871);
   U13218 : XNOR2_X1 port map( A => n24872, B => n18087, ZN => n18090);
   U13245 : XNOR2_X1 port map( A => n18086, B => n18085, ZN => n24872);
   U13303 : NAND3_X1 port map( A1 => n24281, A2 => n25181, A3 => n24873, ZN => 
                           n25145);
   U13441 : NAND3_X1 port map( A1 => n24875, A2 => n22737, A3 => n24874, ZN => 
                           n22740);
   U13456 : NAND2_X1 port map( A1 => n23495, A2 => n23483, ZN => n24875);
   U13468 : NAND2_X1 port map( A1 => n5063, A2 => n3442, ZN => n12449);
   U13480 : NAND2_X1 port map( A1 => n2539, A2 => n2997, ZN => n2538);
   U13518 : BUF_X1 port map( A => n22939, Z => n25063);
   U13529 : INV_X1 port map( A => n7733, ZN => n25151);
   U13535 : OR2_X1 port map( A1 => n13047, A2 => n13046, ZN => n24876);
   U13572 : MUX2_X1 port map( A => n13043, B => n13042, S => n13041, Z => 
                           n13047);
   U13600 : OR2_X1 port map( A1 => n23632, A2 => n3164, ZN => n23643);
   U13728 : XNOR2_X1 port map( A => n801, B => n21740, ZN => n24877);
   U13839 : XNOR2_X1 port map( A => n801, B => n21740, ZN => n22911);
   U13842 : OR2_X1 port map( A1 => n15804, A2 => n15857, ZN => n24171);
   U13907 : INV_X1 port map( A => n23420, ZN => n142);
   U13937 : XNOR2_X1 port map( A => n20664, B => n20663, ZN => n24881);
   U13952 : XNOR2_X1 port map( A => n20664, B => n20663, ZN => n22389);
   U14046 : XNOR2_X1 port map( A => n24882, B => n21993, ZN => n22002);
   U14151 : XOR2_X1 port map( A => n1381, B => n24986, Z => n24882);
   U14229 : OR3_X1 port map( A1 => n25474, A2 => n19345, A3 => n5280, ZN => 
                           n5455);
   U14238 : XNOR2_X1 port map( A => n18140, B => n18141, ZN => n19107);
   U14261 : BUF_X1 port map( A => n23543, Z => n24057);
   U14367 : OR2_X1 port map( A1 => n20598, A2 => n20427, ZN => n24883);
   U14532 : XNOR2_X1 port map( A => n21558, B => n21557, ZN => n24884);
   U14540 : XNOR2_X1 port map( A => n21558, B => n21557, ZN => n24885);
   U14541 : NAND2_X1 port map( A1 => n835, A2 => n2854, ZN => n20039);
   U14561 : NAND3_X1 port map( A1 => n17458, A2 => n17459, A3 => n522, ZN => 
                           n24886);
   U14585 : CLKBUF_X1 port map( A => n3016, Z => n24887);
   U14603 : NAND3_X1 port map( A1 => n17458, A2 => n17459, A3 => n522, ZN => 
                           n18499);
   U14671 : AND2_X1 port map( A1 => n16614, A2 => n16613, ZN => n24888);
   U14683 : AOI21_X1 port map( B1 => n21927, B2 => n21926, A => n21925, ZN => 
                           n23184);
   U14686 : XNOR2_X1 port map( A => n13371, B => n13372, ZN => n24890);
   U14695 : NAND2_X2 port map( A1 => n19001, A2 => n2927, ZN => n20536);
   U14696 : NOR2_X1 port map( A1 => n24891, A2 => n24892, ZN => n5768);
   U14697 : AND2_X1 port map( A1 => n22922, A2 => n25070, ZN => n24891);
   U14704 : NOR2_X1 port map( A1 => n24379, A2 => n22922, ZN => n24892);
   U14705 : XOR2_X1 port map( A => n18458, B => n18568, Z => n18118);
   U14706 : AND2_X1 port map( A1 => n23146, A2 => n1349, ZN => n23160);
   U14707 : OR2_X1 port map( A1 => n22106, A2 => n22105, ZN => n24893);
   U14711 : NAND4_X2 port map( A1 => n21821, A2 => n21820, A3 => n21819, A4 => 
                           n21818, ZN => n24895);
   U14901 : INV_X1 port map( A => n12583, ZN => n12977);
   U14928 : NAND3_X1 port map( A1 => n2363, A2 => n2362, A3 => n2360, ZN => 
                           n24896);
   U14939 : NAND3_X1 port map( A1 => n2363, A2 => n2362, A3 => n2360, ZN => 
                           n21176);
   U14973 : OR2_X1 port map( A1 => n24897, A2 => n20395, ZN => n2425);
   U15011 : OR2_X1 port map( A1 => n1327, A2 => n20384, ZN => n24897);
   U15128 : NAND2_X1 port map( A1 => n3563, A2 => n13485, ZN => n4382);
   U15155 : NAND2_X1 port map( A1 => n24155, A2 => n24154, ZN => n21665);
   U15173 : OAI211_X1 port map( C1 => n19945, C2 => n20960, A => n19943, B => 
                           n71, ZN => n24899);
   U15195 : OAI211_X1 port map( C1 => n19945, C2 => n20960, A => n19943, B => 
                           n71, ZN => n21522);
   U15225 : XNOR2_X1 port map( A => n21083, B => n21082, ZN => n23997);
   U15248 : NOR2_X1 port map( A1 => n19626, A2 => n19625, ZN => n24469);
   U15290 : NAND2_X1 port map( A1 => n21773, A2 => n2513, ZN => n24901);
   U15296 : NAND2_X1 port map( A1 => n21773, A2 => n2513, ZN => n23594);
   U15300 : XNOR2_X1 port map( A => n20953, B => n20952, ZN => n24902);
   U15306 : NOR2_X1 port map( A1 => n22405, A2 => n22404, ZN => n24903);
   U15315 : NOR2_X1 port map( A1 => n22405, A2 => n22404, ZN => n24904);
   U15411 : XNOR2_X1 port map( A => n19903, B => n19902, ZN => n24905);
   U15429 : AND3_X1 port map( A1 => n23805, A2 => n22043, A3 => n21828, ZN => 
                           n21907);
   U15464 : NAND2_X1 port map( A1 => n21377, A2 => n3080, ZN => n24906);
   U15535 : NAND2_X1 port map( A1 => n1587, A2 => n1585, ZN => n24907);
   U15538 : XNOR2_X1 port map( A => n17754, B => n17753, ZN => n24908);
   U15546 : XNOR2_X1 port map( A => n17754, B => n17753, ZN => n24909);
   U15565 : NAND2_X1 port map( A1 => n4633, A2 => n21549, ZN => n24911);
   U15620 : NAND2_X1 port map( A1 => n4633, A2 => n21549, ZN => n23372);
   U15621 : INV_X1 port map( A => n23066, ZN => n25179);
   U15678 : XNOR2_X1 port map( A => n17035, B => n17034, ZN => n19310);
   U15690 : INV_X1 port map( A => n11191, ZN => n24913);
   U15694 : AOI22_X1 port map( A1 => n10271, A2 => n11185, B1 => n11184, B2 => 
                           n10731, ZN => n11370);
   U15695 : AND3_X1 port map( A1 => n22277, A2 => n22276, A3 => n1507, ZN => 
                           n24914);
   U15714 : NOR3_X1 port map( A1 => n20349, A2 => n19654, A3 => n20670, ZN => 
                           n19655);
   U15806 : NOR2_X1 port map( A1 => n19656, A2 => n19655, ZN => n24916);
   U15813 : NOR2_X1 port map( A1 => n19656, A2 => n19655, ZN => n21521);
   U15831 : CLKBUF_X1 port map( A => Key(98), Z => n2735);
   U15839 : XOR2_X1 port map( A => n10880, B => n11602, Z => n10882);
   U15912 : AND2_X1 port map( A1 => n22800, A2 => n22799, ZN => n25161);
   U15984 : OR2_X1 port map( A1 => n17500, A2 => n17499, ZN => n24917);
   U16147 : OAI211_X1 port map( C1 => n22356, C2 => n21785, A => n21784, B => 
                           n21783, ZN => n24921);
   U16259 : OAI211_X1 port map( C1 => n22356, C2 => n21785, A => n21784, B => 
                           n21783, ZN => n23757);
   U16297 : XOR2_X1 port map( A => n21586, B => n21585, Z => n24922);
   U16307 : AND3_X1 port map( A1 => n22679, A2 => n22774, A3 => n5377, ZN => 
                           n24923);
   U16351 : NAND2_X1 port map( A1 => n22682, A2 => n22681, ZN => n24924);
   U16502 : INV_X1 port map( A => n20264, ZN => n20410);
   U16716 : AND2_X1 port map( A1 => n19446, A2 => n19351, ZN => n24926);
   U16755 : XOR2_X1 port map( A => n7472, B => n7473, Z => n24927);
   U16762 : XNOR2_X1 port map( A => n14693, B => n14692, ZN => n24928);
   U16769 : XNOR2_X1 port map( A => n18216, B => n18217, ZN => n24929);
   U16831 : XNOR2_X1 port map( A => n18216, B => n18217, ZN => n19184);
   U16847 : BUF_X2 port map( A => n23869, Z => n23902);
   U16850 : XNOR2_X1 port map( A => n10565, B => n10566, ZN => n24930);
   U16852 : XOR2_X1 port map( A => n17761, B => n17760, Z => n24931);
   U16854 : XNOR2_X1 port map( A => n10565, B => n10566, ZN => n12719);
   U16856 : XNOR2_X1 port map( A => n21620, B => n21619, ZN => n24932);
   U16862 : BUF_X1 port map( A => n23391, Z => n24933);
   U16903 : XNOR2_X1 port map( A => n21620, B => n21619, ZN => n22940);
   U16924 : OR3_X1 port map( A1 => n24470, A2 => n10935, A3 => n10505, ZN => 
                           n10598);
   U16928 : AOI21_X1 port map( B1 => n23890, B2 => n23904, A => n25239, ZN => 
                           n21866);
   U16930 : INV_X1 port map( A => n16597, ZN => n24935);
   U16967 : NAND2_X1 port map( A1 => n3465, A2 => n3932, ZN => n24936);
   U16968 : NAND2_X1 port map( A1 => n3465, A2 => n3932, ZN => n20792);
   U16969 : NAND4_X1 port map( A1 => n13706, A2 => n13704, A3 => n13705, A4 => 
                           n13707, ZN => n24937);
   U16971 : NAND4_X1 port map( A1 => n13706, A2 => n13704, A3 => n13705, A4 => 
                           n13707, ZN => n24938);
   U17021 : NAND4_X1 port map( A1 => n13706, A2 => n13704, A3 => n13705, A4 => 
                           n13707, ZN => n15040);
   U17023 : INV_X1 port map( A => n20414, ZN => n25108);
   U17083 : AND2_X1 port map( A1 => n3810, A2 => n3809, ZN => n20578);
   U17084 : NAND2_X1 port map( A1 => n5583, A2 => n5582, ZN => n24941);
   U17101 : AND2_X1 port map( A1 => n14, A2 => n25165, ZN => n24942);
   U17106 : CLKBUF_X1 port map( A => n4052, Z => n24943);
   U17226 : XOR2_X1 port map( A => n6222, B => n6221, Z => n24944);
   U17238 : NOR2_X1 port map( A1 => n7214, A2 => n7213, ZN => n24946);
   U17239 : NOR2_X1 port map( A1 => n7214, A2 => n7213, ZN => n8781);
   U17240 : BUF_X1 port map( A => n23410, Z => n24947);
   U17260 : OR2_X1 port map( A1 => n21148, A2 => n21149, ZN => n25024);
   U17288 : MUX2_X1 port map( A => n22372, B => n22371, S => n22680, Z => 
                           n23939);
   U17336 : OAI211_X1 port map( C1 => n18726, C2 => n19376, A => n18725, B => 
                           n4317, ZN => n20181);
   U17347 : INV_X1 port map( A => n20126, ZN => n25101);
   U17355 : INV_X1 port map( A => n9874, ZN => n307);
   U17357 : NOR2_X1 port map( A1 => n20136, A2 => n20019, ZN => n24950);
   U17381 : XNOR2_X1 port map( A => n20705, B => n20704, ZN => n24951);
   U17382 : XNOR2_X1 port map( A => n20705, B => n20704, ZN => n22566);
   U17385 : INV_X1 port map( A => n23120, ZN => n24952);
   U17386 : OR2_X2 port map( A1 => n19899, A2 => n19898, ZN => n21621);
   U17391 : XOR2_X1 port map( A => n21264, B => n21263, Z => n24953);
   U17452 : NAND3_X1 port map( A1 => n22795, A2 => n22797, A3 => n22796, ZN => 
                           n24954);
   U17527 : NAND3_X1 port map( A1 => n22795, A2 => n22797, A3 => n22796, ZN => 
                           n24006);
   U17569 : NOR2_X1 port map( A1 => n20721, A2 => n20720, ZN => n24955);
   U17570 : OAI21_X1 port map( B1 => n5620, B2 => n14415, A => n13859, ZN => 
                           n24956);
   U17571 : OAI21_X1 port map( B1 => n5620, B2 => n14415, A => n13859, ZN => 
                           n15478);
   U17572 : NAND4_X1 port map( A1 => n8575, A2 => n8572, A3 => n8574, A4 => 
                           n8573, ZN => n11169);
   U17634 : INV_X1 port map( A => n14849, ZN => n24958);
   U17635 : XNOR2_X1 port map( A => n7241, B => n7240, ZN => n24959);
   U17720 : XNOR2_X1 port map( A => n7241, B => n7240, ZN => n2585);
   U17754 : XNOR2_X1 port map( A => n13641, B => n13642, ZN => n24960);
   U17872 : XNOR2_X1 port map( A => n18305, B => n24961, ZN => n18119);
   U17889 : XOR2_X1 port map( A => n18675, B => n1856, Z => n24961);
   U17890 : AOI21_X1 port map( B1 => n19671, B2 => n18887, A => n18886, ZN => 
                           n24962);
   U17963 : XNOR2_X1 port map( A => n21118, B => n21119, ZN => n24963);
   U18075 : AOI21_X1 port map( B1 => n19671, B2 => n18887, A => n18886, ZN => 
                           n21597);
   U18111 : OAI21_X2 port map( B1 => n12497, B2 => n12496, A => n12495, ZN => 
                           n14377);
   U18136 : NAND4_X1 port map( A1 => n10266, A2 => n10265, A3 => n10267, A4 => 
                           n10264, ZN => n24964);
   U18205 : XNOR2_X1 port map( A => n667, B => n11763, ZN => n24965);
   U18245 : NAND4_X1 port map( A1 => n10266, A2 => n10265, A3 => n10267, A4 => 
                           n10264, ZN => n12383);
   U18289 : XNOR2_X1 port map( A => n667, B => n11763, ZN => n12569);
   U18326 : AND2_X1 port map( A1 => n14685, A2 => n14686, ZN => n24966);
   U18365 : XNOR2_X1 port map( A => n11972, B => n11973, ZN => n24346);
   U18367 : NAND3_X1 port map( A1 => n4352, A2 => n3476, A3 => n4349, ZN => 
                           n24967);
   U18466 : XNOR2_X1 port map( A => n17793, B => n17794, ZN => n24968);
   U18634 : NOR2_X1 port map( A1 => n1169, A2 => n10723, ZN => n24969);
   U18636 : NOR2_X1 port map( A1 => n1169, A2 => n10723, ZN => n24970);
   U18645 : NOR2_X1 port map( A1 => n1169, A2 => n10723, ZN => n12138);
   U18670 : XNOR2_X1 port map( A => n20694, B => n20693, ZN => n24971);
   U18673 : XNOR2_X1 port map( A => n20694, B => n20693, ZN => n22564);
   U18675 : AND2_X1 port map( A1 => n2117, A2 => n2116, ZN => n24973);
   U18690 : NAND2_X1 port map( A1 => n4015, A2 => n1836, ZN => n24975);
   U18747 : INV_X1 port map( A => n23411, ZN => n24977);
   U18771 : INV_X1 port map( A => n23411, ZN => n24978);
   U18836 : OAI211_X1 port map( C1 => n9279, C2 => n9649, A => n9648, B => 
                           n9647, ZN => n24980);
   U18847 : INV_X1 port map( A => n15696, ZN => n24981);
   U18848 : OAI211_X1 port map( C1 => n9279, C2 => n9649, A => n9648, B => 
                           n9647, ZN => n11782);
   U18849 : XNOR2_X1 port map( A => n18488, B => n18487, ZN => n24982);
   U18868 : NAND2_X1 port map( A1 => n4434, A2 => n23001, ZN => n24983);
   U18879 : XNOR2_X1 port map( A => n18488, B => n18487, ZN => n19057);
   U18953 : XOR2_X1 port map( A => n8425, B => n8424, Z => n24984);
   U18959 : OAI21_X1 port map( B1 => n200, B2 => n19927, A => n19926, ZN => 
                           n24985);
   U18961 : OAI21_X1 port map( B1 => n200, B2 => n19927, A => n19926, ZN => 
                           n24986);
   U18986 : OAI21_X1 port map( B1 => n200, B2 => n19927, A => n19926, ZN => 
                           n21992);
   U18988 : OAI21_X1 port map( B1 => n22856, B2 => n22855, A => n22854, ZN => 
                           n23410);
   U18996 : INV_X1 port map( A => n12218, ZN => n24987);
   U19000 : AND3_X1 port map( A1 => n10214, A2 => n10213, A3 => n4327, ZN => 
                           n12261);
   U19023 : NOR2_X1 port map( A1 => n3411, A2 => n22803, ZN => n25159);
   U19040 : XNOR2_X1 port map( A => n11844, B => n11843, ZN => n24988);
   U19041 : OR2_X1 port map( A1 => n22489, A2 => n22488, ZN => n24989);
   U19049 : XNOR2_X1 port map( A => n11844, B => n11843, ZN => n13279);
   U19055 : INV_X1 port map( A => n11242, ZN => n12152);
   U19080 : XOR2_X1 port map( A => n25396, B => n11289, Z => n24990);
   U19082 : INV_X1 port map( A => n997, ZN => n24991);
   U19084 : INV_X1 port map( A => n24559, ZN => n25115);
   U19085 : CLKBUF_X1 port map( A => n22805, Z => n24992);
   U19133 : NOR2_X1 port map( A1 => n22477, A2 => n22476, ZN => n24993);
   U19184 : XNOR2_X1 port map( A => n21235, B => n21234, ZN => n22805);
   U19186 : INV_X1 port map( A => n6529, ZN => n24994);
   U19205 : INV_X1 port map( A => n13088, ZN => n24995);
   U19210 : CLKBUF_X1 port map( A => n6060, Z => n6734);
   U19277 : XOR2_X1 port map( A => n18484, B => n18356, Z => n17994);
   U19284 : NAND4_X1 port map( A1 => n20305, A2 => n5764, A3 => n20304, A4 => 
                           n20303, ZN => n24996);
   U19307 : NAND4_X1 port map( A1 => n20305, A2 => n5764, A3 => n20304, A4 => 
                           n20303, ZN => n21569);
   U19313 : OAI211_X1 port map( C1 => n22179, C2 => n24369, A => n22177, B => 
                           n22178, ZN => n2305);
   U19316 : NAND2_X1 port map( A1 => n10395, A2 => n10394, ZN => n24999);
   U19327 : NAND3_X1 port map( A1 => n1269, A2 => n15635, A3 => n15636, ZN => 
                           n25000);
   U19338 : BUF_X1 port map( A => n19595, Z => n25001);
   U19355 : XNOR2_X1 port map( A => n18029, B => n18030, ZN => n19595);
   U19363 : XNOR2_X1 port map( A => n797, B => n17677, ZN => n25002);
   U19417 : OAI21_X1 port map( B1 => n16168, B2 => n16167, A => n16166, ZN => 
                           n25003);
   U19418 : OAI21_X1 port map( B1 => n16168, B2 => n16167, A => n16166, ZN => 
                           n17195);
   U19459 : XOR2_X1 port map( A => n8844, B => n8577, Z => n8582);
   U19491 : BUF_X1 port map( A => n23332, Z => n25004);
   U19492 : XNOR2_X1 port map( A => n21410, B => n21411, ZN => n23332);
   U19564 : XOR2_X1 port map( A => n8767, B => n8768, Z => n25005);
   U19567 : XNOR2_X1 port map( A => n18660, B => n18611, ZN => n25006);
   U19568 : XNOR2_X1 port map( A => n5255, B => n8441, ZN => n7146);
   U19615 : XOR2_X1 port map( A => n8811, B => n8810, Z => n25007);
   U19641 : AOI22_X1 port map( A1 => n13570, A2 => n13571, B1 => n13572, B2 => 
                           n13573, ZN => n25008);
   U19682 : XNOR2_X1 port map( A => n15157, B => n15158, ZN => n25009);
   U19696 : AOI22_X1 port map( A1 => n13570, A2 => n13571, B1 => n13572, B2 => 
                           n13573, ZN => n14488);
   U19787 : XNOR2_X1 port map( A => n15157, B => n15158, ZN => n16267);
   U19788 : INV_X1 port map( A => n2216, ZN => n25010);
   U19793 : XNOR2_X1 port map( A => n17778, B => n2029, ZN => n4114);
   U19832 : INV_X1 port map( A => n20036, ZN => n22233);
   U19880 : BUF_X1 port map( A => n13643, Z => n25011);
   U19882 : OAI211_X1 port map( C1 => n13060, C2 => n3065, A => n13059, B => 
                           n13058, ZN => n13643);
   U19883 : XNOR2_X1 port map( A => n18511, B => n18510, ZN => n25012);
   U19888 : OAI211_X1 port map( C1 => n3889, C2 => n13804, A => n13803, B => 
                           n13802, ZN => n25013);
   U19895 : XNOR2_X1 port map( A => n14641, B => n14640, ZN => n15802);
   U19902 : XNOR2_X1 port map( A => n5864, B => Key(24), ZN => n25014);
   U19909 : CLKBUF_X1 port map( A => n12607, Z => n25015);
   U19956 : OAI211_X1 port map( C1 => n22675, C2 => n22674, A => n22673, B => 
                           n22672, ZN => n25017);
   U19957 : NOR2_X1 port map( A1 => n8663, A2 => n8662, ZN => n11840);
   U19995 : OAI211_X1 port map( C1 => n25208, C2 => n25128, A => n14240, B => 
                           n25127, ZN => n2741);
   U19997 : XNOR2_X1 port map( A => n20931, B => n20930, ZN => n25018);
   U20000 : XNOR2_X1 port map( A => n20931, B => n20930, ZN => n22208);
   U20022 : OAI211_X1 port map( C1 => n14125, C2 => n3851, A => n3849, B => 
                           n3850, ZN => n25019);
   U20097 : OAI211_X1 port map( C1 => n14125, C2 => n3851, A => n3849, B => 
                           n3850, ZN => n15480);
   U20100 : XNOR2_X1 port map( A => n9035, B => n5014, ZN => n25020);
   U20149 : INV_X1 port map( A => n15164, ZN => n2765);
   U20188 : XOR2_X1 port map( A => n8110, B => n8111, Z => n25021);
   U20225 : XNOR2_X1 port map( A => n21125, B => n21124, ZN => n25022);
   U20245 : XNOR2_X1 port map( A => n21125, B => n21124, ZN => n25023);
   U20248 : AOI21_X1 port map( B1 => n5517, B2 => n5519, A => n4871, ZN => 
                           n11209);
   U20249 : OAI211_X1 port map( C1 => n10818, C2 => n10817, A => n3594, B => 
                           n3595, ZN => n25027);
   U20496 : OAI211_X1 port map( C1 => n10818, C2 => n10817, A => n3594, B => 
                           n3595, ZN => n12112);
   U20510 : NOR2_X1 port map( A1 => n25029, A2 => n17568, ZN => n25028);
   U20588 : AND2_X1 port map( A1 => n17566, A2 => n20317, ZN => n25029);
   U20634 : OAI21_X2 port map( B1 => n18970, B2 => n17553, A => n17552, ZN => 
                           n19889);
   U20643 : XNOR2_X1 port map( A => n14700, B => n14701, ZN => n25030);
   U20657 : INV_X1 port map( A => n15631, ZN => n25031);
   U20675 : XNOR2_X1 port map( A => n14700, B => n14701, ZN => n15782);
   U20684 : NOR3_X1 port map( A1 => n14058, A2 => n13521, A3 => n14054, ZN => 
                           n13522);
   U20694 : XNOR2_X1 port map( A => n10640, B => n10639, ZN => n25033);
   U20704 : OR2_X1 port map( A1 => n17714, A2 => n17713, ZN => n25034);
   U20731 : XOR2_X1 port map( A => n11798, B => n11799, Z => n11802);
   U20738 : AOI22_X1 port map( A1 => n14074, A2 => n14078, B1 => n13852, B2 => 
                           n14077, ZN => n25036);
   U20739 : AOI22_X1 port map( A1 => n14074, A2 => n14078, B1 => n13852, B2 => 
                           n14077, ZN => n13491);
   U20747 : AND3_X1 port map( A1 => n24277, A2 => n24276, A3 => n6029, ZN => 
                           n25037);
   U20749 : INV_X1 port map( A => n16602, ZN => n25038);
   U20761 : NAND2_X1 port map( A1 => n16604, A2 => n25038, ZN => n25039);
   U20817 : OAI21_X1 port map( B1 => n19877, B2 => n25221, A => n19876, ZN => 
                           n25040);
   U20846 : OAI21_X1 port map( B1 => n19877, B2 => n25221, A => n19876, ZN => 
                           n21133);
   U20919 : NOR2_X1 port map( A1 => n22489, A2 => n22488, ZN => n25042);
   U20987 : NOR2_X1 port map( A1 => n22489, A2 => n22488, ZN => n23441);
   U20995 : XNOR2_X1 port map( A => n8608, B => n8607, ZN => n25043);
   U20996 : XNOR2_X1 port map( A => n8608, B => n8607, ZN => n10007);
   U21022 : XNOR2_X1 port map( A => n5991, B => Key(104), ZN => n25044);
   U21027 : XNOR2_X1 port map( A => n5991, B => Key(104), ZN => n25045);
   U21028 : XNOR2_X1 port map( A => n5991, B => Key(104), ZN => n6602);
   U21037 : XNOR2_X1 port map( A => n8326, B => n5619, ZN => n25046);
   U21041 : INV_X1 port map( A => n4931, ZN => n25047);
   U21048 : XOR2_X1 port map( A => n12260, B => n12221, Z => n25048);
   U21102 : XOR2_X1 port map( A => n11327, B => n11326, Z => n25049);
   U21105 : CLKBUF_X1 port map( A => n22214, Z => n25050);
   U21108 : OAI21_X1 port map( B1 => n21790, B2 => n22222, A => n2734, ZN => 
                           n25051);
   U21112 : XNOR2_X1 port map( A => n21323, B => n21322, ZN => n22214);
   U21123 : OAI21_X1 port map( B1 => n21790, B2 => n22222, A => n2734, ZN => 
                           n23770);
   U21124 : XNOR2_X1 port map( A => n17746, B => n17747, ZN => n25052);
   U21134 : XNOR2_X1 port map( A => n17746, B => n17747, ZN => n19217);
   U21149 : XNOR2_X1 port map( A => n3205, B => n3204, ZN => n25053);
   U21176 : INV_X1 port map( A => n3662, ZN => n25054);
   U21209 : XNOR2_X1 port map( A => n3205, B => n3204, ZN => n13358);
   U21223 : CLKBUF_X1 port map( A => n23441, Z => n23450);
   U21251 : CLKBUF_X1 port map( A => n23464, Z => n25055);
   U21252 : XNOR2_X1 port map( A => n13576, B => n13577, ZN => n16200);
   U21271 : XNOR2_X1 port map( A => n18231, B => n18230, ZN => n25057);
   U21280 : XNOR2_X1 port map( A => n18231, B => n18230, ZN => n19548);
   U21291 : NOR2_X1 port map( A1 => n22571, A2 => n21938, ZN => n25059);
   U21298 : NOR2_X1 port map( A1 => n22571, A2 => n21938, ZN => n23186);
   U21357 : MUX2_X1 port map( A => n19380, B => n17980, S => n19378, Z => n3518
                           );
   U21376 : XNOR2_X1 port map( A => n11656, B => n11655, ZN => n25061);
   U21388 : OAI211_X1 port map( C1 => n24077, C2 => n19941, A => n2946, B => 
                           n679, ZN => n25062);
   U21394 : OAI211_X1 port map( C1 => n24077, C2 => n19941, A => n2946, B => 
                           n679, ZN => n21312);
   U21395 : XNOR2_X2 port map( A => n11636, B => n11635, ZN => n12490);
   U21424 : XNOR2_X1 port map( A => n8300, B => n8299, ZN => n25064);
   U21467 : OAI211_X1 port map( C1 => n19639, C2 => n347, A => n19638, B => 
                           n19637, ZN => n25065);
   U21534 : OAI211_X1 port map( C1 => n19639, C2 => n347, A => n19638, B => 
                           n19637, ZN => n21640);
   U21537 : XNOR2_X1 port map( A => n21155, B => n21156, ZN => n25066);
   U21545 : XNOR2_X1 port map( A => n21155, B => n21156, ZN => n22317);
   U21546 : XOR2_X1 port map( A => n17979, B => n17978, Z => n25067);
   U21547 : XOR2_X1 port map( A => n21131, B => n21130, Z => n25068);
   U21571 : XNOR2_X1 port map( A => n8156, B => n8155, ZN => n25069);
   U21581 : XNOR2_X1 port map( A => n8156, B => n8155, ZN => n9885);
   U21582 : OR2_X1 port map( A1 => n23155, A2 => n23154, ZN => n23147);
   U21596 : XNOR2_X1 port map( A => n20998, B => n20997, ZN => n25070);
   U21615 : XNOR2_X1 port map( A => n20998, B => n20997, ZN => n22928);
   U21660 : NOR2_X1 port map( A1 => n840, A2 => n22112, ZN => n23546);
   U21826 : OAI21_X1 port map( B1 => n9840, B2 => n10099, A => n9839, ZN => 
                           n25074);
   U21924 : XNOR2_X1 port map( A => n20441, B => n20440, ZN => n25075);
   U21927 : INV_X1 port map( A => n878, ZN => n25076);
   U21937 : XNOR2_X1 port map( A => n20441, B => n20440, ZN => n22657);
   U21944 : OAI21_X1 port map( B1 => n4470, B2 => n4469, A => n481, ZN => 
                           n23972);
   U22007 : XOR2_X1 port map( A => n20891, B => n20890, Z => n25078);
   U22099 : XNOR2_X2 port map( A => n10392, B => n11284, ZN => n12652);
   U22120 : XNOR2_X1 port map( A => n21089, B => n21090, ZN => n25079);
   U22146 : XNOR2_X1 port map( A => n21089, B => n21090, ZN => n23996);
   U22185 : XOR2_X1 port map( A => n4996, B => n4995, Z => n25080);
   U22188 : XNOR2_X1 port map( A => n21426, B => n21425, ZN => n25081);
   U22197 : XNOR2_X1 port map( A => n21426, B => n21425, ZN => n23336);
   U22223 : XOR2_X1 port map( A => n20083, B => n20082, Z => n25082);
   U22245 : AOI21_X1 port map( B1 => n782, B2 => n22362, A => n1249, ZN => 
                           n25083);
   U22281 : AOI21_X1 port map( B1 => n782, B2 => n22362, A => n1249, ZN => 
                           n25084);
   U22301 : AOI21_X1 port map( B1 => n782, B2 => n22362, A => n1249, ZN => 
                           n23940);
   U22340 : INV_X1 port map( A => n18883, ZN => n25086);
   U22354 : XNOR2_X1 port map( A => n11418, B => n11417, ZN => n12795);
   U22372 : OAI211_X1 port map( C1 => n10610, C2 => n9610, A => n9609, B => 
                           n9608, ZN => n25087);
   U22396 : NOR2_X1 port map( A1 => n18787, A2 => n18786, ZN => n25088);
   U22405 : NOR2_X1 port map( A1 => n18787, A2 => n18786, ZN => n25089);
   U22412 : OAI211_X1 port map( C1 => n10610, C2 => n9610, A => n9609, B => 
                           n9608, ZN => n12143);
   U22428 : NOR2_X1 port map( A1 => n19685, A2 => n21066, ZN => n25091);
   U22429 : NOR2_X1 port map( A1 => n19685, A2 => n21066, ZN => n21997);
   U22430 : XNOR2_X1 port map( A => n13476, B => n13475, ZN => n25092);
   U22444 : NAND4_X2 port map( A1 => n4780, A2 => n19844, A3 => n25094, A4 => 
                           n25093, ZN => n21974);
   U22455 : NAND2_X1 port map( A1 => n1205, A2 => n3198, ZN => n25093);
   U22516 : NAND2_X1 port map( A1 => n1206, A2 => n24194, ZN => n25094);
   U22540 : NAND3_X1 port map( A1 => n4116, A2 => n13935, A3 => n13200, ZN => 
                           n13202);
   U22578 : NAND3_X1 port map( A1 => n10142, A2 => n9821, A3 => n24026, ZN => 
                           n9822);
   U22628 : NAND2_X1 port map( A1 => n9918, A2 => n9462, ZN => n9912);
   U22675 : AND2_X1 port map( A1 => n5376, A2 => n16795, ZN => n4553);
   U22680 : NOR2_X1 port map( A1 => n12767, A2 => n13217, ZN => n12809);
   U22682 : XNOR2_X2 port map( A => n11236, B => n11235, ZN => n12767);
   U22713 : NAND2_X1 port map( A1 => n25095, A2 => n1170, ZN => n1169);
   U22728 : NAND2_X1 port map( A1 => n1167, A2 => n1166, ZN => n25095);
   U22736 : NAND2_X1 port map( A1 => n24927, A2 => n9965, ZN => n1602);
   U22760 : AOI21_X1 port map( B1 => n6608, B2 => n6112, A => n6714, ZN => 
                           n5786);
   U22804 : NAND2_X1 port map( A1 => n6232, A2 => n6715, ZN => n6608);
   U22807 : NAND2_X1 port map( A1 => n5033, A2 => n1491, ZN => n5028);
   U22848 : NAND3_X1 port map( A1 => n5035, A2 => n24941, A3 => n5037, ZN => 
                           n5033);
   U22849 : OR2_X1 port map( A1 => n5800, A2 => n6575, ZN => n4755);
   U22850 : OAI21_X1 port map( B1 => n25097, B2 => n13266, A => n25096, ZN => 
                           n12681);
   U22879 : NAND2_X1 port map( A1 => n13266, A2 => n13264, ZN => n25096);
   U22887 : INV_X1 port map( A => n24443, ZN => n25097);
   U22908 : NAND2_X1 port map( A1 => n12705, A2 => n25098, ZN => n14960);
   U22924 : NAND2_X1 port map( A1 => n25099, A2 => n177, ZN => n25098);
   U22971 : INV_X1 port map( A => n16351, ZN => n25100);
   U22975 : NAND2_X1 port map( A1 => n16350, A2 => n25100, ZN => n25165);
   U22979 : NAND3_X1 port map( A1 => n19675, A2 => n25102, A3 => n25101, ZN => 
                           n4570);
   U23002 : NAND2_X1 port map( A1 => n20130, A2 => n20546, ZN => n25102);
   U23017 : NAND2_X1 port map( A1 => n13518, A2 => n1355, ZN => n13610);
   U23018 : NOR2_X2 port map( A1 => n2706, A2 => n25104, ZN => n20460);
   U23029 : OAI22_X1 port map( A1 => n19385, A2 => n24908, B1 => n19391, B2 => 
                           n5196, ZN => n25104);
   U23043 : XNOR2_X1 port map( A => n20700, B => n20701, ZN => n20867);
   U23058 : NAND3_X1 port map( A1 => n17735, A2 => n17730, A3 => n17486, ZN => 
                           n16815);
   U23060 : NAND3_X1 port map( A1 => n16746, A2 => n17279, A3 => n17277, ZN => 
                           n16747);
   U23084 : NAND3_X1 port map( A1 => n18714, A2 => n19351, A3 => n19451, ZN => 
                           n25105);
   U23100 : NAND2_X1 port map( A1 => n5162, A2 => n7237, ZN => n8980);
   U23110 : NAND3_X1 port map( A1 => n1984, A2 => n5163, A3 => n1345, ZN => 
                           n5162);
   U23123 : NAND2_X1 port map( A1 => n25106, A2 => n17164, ZN => n687);
   U23127 : INV_X1 port map( A => n16836, ZN => n25106);
   U23128 : NAND2_X1 port map( A1 => n4775, A2 => n17165, ZN => n16836);
   U23145 : AOI22_X2 port map( A1 => n3547, A2 => n16172, B1 => n16174, B2 => 
                           n16173, ZN => n17192);
   U23150 : NAND2_X1 port map( A1 => n25107, A2 => n13307, ZN => n1564);
   U23153 : NAND2_X1 port map( A1 => n16056, A2 => n4972, ZN => n16059);
   U23241 : NAND2_X1 port map( A1 => n25110, A2 => n25109, ZN => n11224);
   U23243 : NAND2_X1 port map( A1 => n11222, A2 => n13137, ZN => n25109);
   U23247 : NAND2_X1 port map( A1 => n25112, A2 => n25111, ZN => n25110);
   U23295 : INV_X1 port map( A => n13137, ZN => n25111);
   U23299 : NAND2_X1 port map( A1 => n11142, A2 => n12437, ZN => n25112);
   U23310 : NAND3_X1 port map( A1 => n19558, A2 => n19555, A3 => n3284, ZN => 
                           n4261);
   U23345 : NAND2_X1 port map( A1 => n25114, A2 => n25113, ZN => n22589);
   U23347 : NAND2_X1 port map( A1 => n22582, A2 => n24561, ZN => n25113);
   U23356 : NAND2_X1 port map( A1 => n22583, A2 => n25115, ZN => n25114);
   U23367 : NAND3_X1 port map( A1 => n5250, A2 => n6904, A3 => n5249, ZN => 
                           n5248);
   U23398 : NAND3_X2 port map( A1 => n7058, A2 => n25118, A3 => n25117, ZN => 
                           n9044);
   U23416 : NAND2_X1 port map( A1 => n3248, A2 => n7809, ZN => n25118);
   U23417 : NAND2_X1 port map( A1 => n21829, A2 => n22219, ZN => n22162);
   U23418 : NAND2_X1 port map( A1 => n2788, A2 => n6968, ZN => n7065);
   U23420 : NAND3_X1 port map( A1 => n13950, A2 => n3069, A3 => n13949, ZN => 
                           n1836);
   U23424 : NAND3_X1 port map( A1 => n24195, A2 => n15628, A3 => n15629, ZN => 
                           n15631);
   U23428 : NAND2_X1 port map( A1 => n25005, A2 => n9977, ZN => n9416);
   U23432 : NAND2_X1 port map( A1 => n25250, A2 => n10556, ZN => n10657);
   U23457 : NAND2_X1 port map( A1 => n9745, A2 => n9990, ZN => n25119);
   U23473 : AOI21_X1 port map( B1 => n25121, B2 => n24534, A => n9991, ZN => 
                           n25120);
   U23474 : AOI21_X1 port map( B1 => n9351, B2 => n9460, A => n1470, ZN => 
                           n9358);
   U23515 : NAND2_X1 port map( A1 => n118, A2 => n119, ZN => n18129);
   U23613 : NAND3_X1 port map( A1 => n13325, A2 => n12952, A3 => n13329, ZN => 
                           n12847);
   U23625 : AND3_X2 port map( A1 => n5501, A2 => n4363, A3 => n1458, ZN => 
                           n20507);
   U23679 : NAND2_X1 port map( A1 => n22292, A2 => n25122, ZN => n23252);
   U23693 : NAND2_X1 port map( A1 => n25124, A2 => n25123, ZN => n25122);
   U23764 : INV_X1 port map( A => n22293, ZN => n25124);
   U23865 : NAND2_X1 port map( A1 => n25126, A2 => n25125, ZN => n20283);
   U23867 : NAND2_X1 port map( A1 => n20282, A2 => n20281, ZN => n25125);
   U23962 : NAND2_X1 port map( A1 => n4460, A2 => n24414, ZN => n25126);
   U23963 : NAND2_X1 port map( A1 => n25208, A2 => n14244, ZN => n25127);
   U24024 : NAND2_X1 port map( A1 => n5760, A2 => n17122, ZN => n25129);
   U24078 : NAND2_X1 port map( A1 => n19486, A2 => n25440, ZN => n25130);
   U24111 : OAI21_X1 port map( B1 => n19806, B2 => n20235, A => n25132, ZN => 
                           n19807);
   U24131 : NAND3_X1 port map( A1 => n19804, A2 => n25205, A3 => n20170, ZN => 
                           n25132);
   U24143 : XNOR2_X1 port map( A => n22014, B => n21522, ZN => n20795);
   U24167 : NAND2_X1 port map( A1 => n14510, A2 => n14439, ZN => n13978);
   U24177 : MUX2_X1 port map( A => n4273, B => n22655, S => n25075, Z => n22658
                           );
   U24181 : NAND2_X1 port map( A1 => n7528, A2 => n7527, ZN => n25133);
   U24204 : NAND2_X1 port map( A1 => n3934, A2 => n10364, ZN => n25135);
   U24205 : NAND2_X1 port map( A1 => n9595, A2 => n10129, ZN => n7440);
   U24206 : OAI22_X1 port map( A1 => n10254, A2 => n24959, B1 => n5057, B2 => 
                           n9211, ZN => n9595);
   U24207 : OR2_X1 port map( A1 => n12433, A2 => n12455, ZN => n12730);
   U24209 : XNOR2_X1 port map( A => n8206, B => n8753, ZN => n25136);
   U24210 : XNOR2_X1 port map( A => n8204, B => n8205, ZN => n25137);
   U24211 : NAND3_X1 port map( A1 => n22233, A2 => n3231, A3 => n22235, ZN => 
                           n1164);
   U24212 : AOI22_X2 port map( A1 => n6167, A2 => n127, B1 => n6166, B2 => 
                           n6542, ZN => n7761);
   U24213 : INV_X1 port map( A => n17330, ZN => n15559);
   U24214 : NAND2_X1 port map( A1 => n3553, A2 => n16309, ZN => n17330);
   U24217 : XNOR2_X1 port map( A => n18198, B => n18476, ZN => n18109);
   U24218 : NAND3_X2 port map( A1 => n16747, A2 => n16764, A3 => n24299, ZN => 
                           n18198);
   U24219 : NAND2_X1 port map( A1 => n21367, A2 => n4350, ZN => n25138);
   U24220 : AND3_X2 port map( A1 => n3188, A2 => n5843, A3 => n5842, ZN => 
                           n7313);
   U24221 : NAND2_X1 port map( A1 => n11678, A2 => n11677, ZN => n24165);
   U24222 : NAND3_X1 port map( A1 => n15557, A2 => n24297, A3 => n16012, ZN => 
                           n634);
   U24223 : NAND2_X1 port map( A1 => n1152, A2 => n25139, ZN => n1150);
   U24225 : XNOR2_X1 port map( A => n17804, B => n17805, ZN => n25140);
   U24226 : NAND2_X1 port map( A1 => n11170, A2 => n11169, ZN => n10313);
   U24227 : NAND3_X1 port map( A1 => n17242, A2 => n17346, A3 => n17241, ZN => 
                           n16136);
   U24229 : NAND2_X1 port map( A1 => n22883, A2 => n24879, ZN => n25141);
   U24230 : INV_X1 port map( A => n22882, ZN => n25142);
   U24231 : AND3_X2 port map( A1 => n1262, A2 => n1264, A3 => n5558, ZN => 
                           n12214);
   U24232 : NAND2_X1 port map( A1 => n25143, A2 => n5478, ZN => n5477);
   U24233 : NAND2_X1 port map( A1 => n5480, A2 => n19270, ZN => n25143);
   U24234 : NAND2_X1 port map( A1 => n10616, A2 => n10412, ZN => n24521);
   U24235 : NAND3_X1 port map( A1 => n25144, A2 => n4852, A3 => n4851, ZN => 
                           n20360);
   U24236 : NAND2_X1 port map( A1 => n4314, A2 => n1212, ZN => n25144);
   U24237 : XNOR2_X1 port map( A => n25145, B => n24280, ZN => Ciphertext(190))
                           ;
   U24238 : NAND3_X1 port map( A1 => n262, A2 => n24927, A3 => n9281, ZN => 
                           n25146);
   U24239 : NAND2_X1 port map( A1 => n25147, A2 => n9505, ZN => n11032);
   U24241 : XNOR2_X1 port map( A => n15350, B => n15190, ZN => n14490);
   U24242 : NAND2_X1 port map( A1 => n9361, A2 => n25148, ZN => n10757);
   U24243 : NAND2_X1 port map( A1 => n24237, A2 => n22842, ZN => n24236);
   U24245 : OAI21_X2 port map( B1 => n15627, B2 => n16097, A => n25149, ZN => 
                           n17059);
   U24246 : NAND2_X1 port map( A1 => n15864, A2 => n15626, ZN => n25149);
   U24247 : NAND3_X1 port map( A1 => n1548, A2 => n2462, A3 => n2463, ZN => 
                           n19924);
   U24250 : OR2_X1 port map( A1 => n17439, A2 => n16962, ZN => n2550);
   U24251 : OAI21_X1 port map( B1 => n7735, B2 => n25151, A => n25150, ZN => 
                           n6251);
   U24252 : NAND2_X1 port map( A1 => n7735, A2 => n7642, ZN => n25150);
   U24253 : NAND3_X1 port map( A1 => n14381, A2 => n14382, A3 => n16154, ZN => 
                           n14396);
   U24254 : NAND3_X2 port map( A1 => n25152, A2 => n7669, A3 => n7668, ZN => 
                           n8673);
   U24255 : NOR2_X2 port map( A1 => n13457, A2 => n25153, ZN => n14477);
   U24256 : OAI22_X1 port map( A1 => n13454, A2 => n24711, B1 => n13889, B2 => 
                           n24710, ZN => n25153);
   U24257 : NAND2_X1 port map( A1 => n7222, A2 => n7474, ZN => n1531);
   U24258 : NAND2_X1 port map( A1 => n3362, A2 => n7421, ZN => n7222);
   U24259 : NAND2_X1 port map( A1 => n6050, A2 => n6630, ZN => n6750);
   U24260 : XNOR2_X2 port map( A => Key(75), B => Plaintext(75), ZN => n6630);
   U24261 : XNOR2_X1 port map( A => n18628, B => n16037, ZN => n16091);
   U24263 : NAND2_X1 port map( A1 => n20142, A2 => n4066, ZN => n20141);
   U24264 : NAND2_X1 port map( A1 => n7460, A2 => n268, ZN => n7467);
   U24265 : NAND2_X1 port map( A1 => n10903, A2 => n10445, ZN => n10443);
   U24266 : NAND2_X1 port map( A1 => n10904, A2 => n10746, ZN => n10903);
   U24267 : NAND2_X1 port map( A1 => n10654, A2 => n10660, ZN => n10399);
   U24268 : NOR2_X1 port map( A1 => n13234, A2 => n13298, ZN => n1445);
   U24269 : INV_X1 port map( A => n7881, ZN => n25154);
   U24270 : NAND2_X1 port map( A1 => n8013, A2 => n8012, ZN => n8019);
   U24271 : NAND2_X1 port map( A1 => n2376, A2 => n2679, ZN => n2394);
   U24272 : NAND2_X1 port map( A1 => n25156, A2 => n25155, ZN => n10455);
   U24273 : NAND2_X1 port map( A1 => n10756, A2 => n10451, ZN => n25155);
   U24274 : NAND2_X1 port map( A1 => n20510, A2 => n20215, ZN => n20508);
   U24275 : NAND2_X1 port map( A1 => n19188, A2 => n19187, ZN => n25157);
   U24276 : NAND2_X1 port map( A1 => n19189, A2 => n19550, ZN => n25158);
   U24277 : NAND2_X1 port map( A1 => n24051, A2 => n6232, ZN => n6607);
   U24278 : AOI21_X1 port map( B1 => n25161, B2 => n25160, A => n25159, ZN => 
                           n21389);
   U24279 : NAND2_X1 port map( A1 => n11178, A2 => n11175, ZN => n10939);
   U24280 : NAND2_X1 port map( A1 => n17040, A2 => n17364, ZN => n25162);
   U24281 : NAND2_X1 port map( A1 => n2469, A2 => n2470, ZN => n2468);
   U24283 : INV_X1 port map( A => n10088, ZN => n25164);
   U24284 : NAND2_X1 port map( A1 => n14, A2 => n25165, ZN => n16980);
   U24285 : NAND2_X1 port map( A1 => n15992, A2 => n15654, ZN => n15660);
   U24286 : XNOR2_X1 port map( A => n25166, B => n12375, ZN => n11463);
   U24287 : NAND2_X2 port map( A1 => n10765, A2 => n734, ZN => n12375);
   U24288 : NAND2_X1 port map( A1 => n11301, A2 => n11298, ZN => n10435);
   U24289 : NAND2_X1 port map( A1 => n6906, A2 => n6905, ZN => n6787);
   U24290 : OAI21_X1 port map( B1 => n1340, B2 => n25168, A => n25167, ZN => 
                           n22654);
   U24291 : NAND2_X1 port map( A1 => n22652, A2 => n1340, ZN => n25167);
   U24292 : INV_X1 port map( A => n22653, ZN => n25168);
   U24293 : NOR2_X1 port map( A1 => n22311, A2 => n25169, ZN => n22312);
   U24294 : NAND2_X1 port map( A1 => n3095, A2 => n3097, ZN => n25169);
   U24295 : NAND2_X1 port map( A1 => n25172, A2 => n25170, ZN => n20392);
   U24296 : NAND2_X1 port map( A1 => n352, A2 => n19345, ZN => n25170);
   U24297 : NAND2_X1 port map( A1 => n20387, A2 => n25440, ZN => n25172);
   U24299 : NAND2_X1 port map( A1 => n25173, A2 => n392, ZN => n599);
   U24300 : NAND2_X1 port map( A1 => n1, A2 => n3, ZN => n25173);
   U24301 : NAND2_X1 port map( A1 => n665, A2 => n25174, ZN => n608);
   U24303 : NAND3_X2 port map( A1 => n952, A2 => n951, A3 => n18857, ZN => 
                           n19849);
   U24304 : NAND2_X1 port map( A1 => n25175, A2 => n593, ZN => n22405);
   U24306 : NAND3_X1 port map( A1 => n24239, A2 => n22905, A3 => n22904, ZN => 
                           n24238);
   U24307 : OR2_X2 port map( A1 => n13668, A2 => n13670, ZN => n14000);
   U24308 : NAND3_X1 port map( A1 => n16727, A2 => n16726, A3 => n16725, ZN => 
                           n16728);
   U24309 : NAND2_X1 port map( A1 => n22464, A2 => n22462, ZN => n21932);
   U24311 : OR2_X1 port map( A1 => n14122, A2 => n13811, ZN => n3849);
   U24312 : NAND2_X1 port map( A1 => n14123, A2 => n14208, ZN => n14122);
   U24313 : NAND3_X1 port map( A1 => n1231, A2 => n5705, A3 => n5707, ZN => 
                           n24269);
   U24314 : NAND2_X1 port map( A1 => n25176, A2 => n576, ZN => n19604);
   U24315 : NAND2_X1 port map( A1 => n19600, A2 => n19601, ZN => n25176);
   U24317 : NAND3_X1 port map( A1 => n23079, A2 => n25178, A3 => n25177, ZN => 
                           n21281);
   U24318 : NAND2_X1 port map( A1 => n23066, A2 => n22578, ZN => n25177);
   U24319 : NAND2_X1 port map( A1 => n25179, A2 => n23064, ZN => n25178);
   U24320 : NAND3_X1 port map( A1 => n3037, A2 => n23188, A3 => n23189, ZN => 
                           n3036);
   U24321 : NAND2_X1 port map( A1 => n19361, A2 => n19211, ZN => n1266);
   U24322 : NOR2_X1 port map( A1 => n16273, A2 => n16274, ZN => n25180);
   U24323 : NAND2_X1 port map( A1 => n24204, A2 => n24019, ZN => n25181);
   U24324 : NAND2_X1 port map( A1 => n6538, A2 => n6530, ZN => n6130);
   U24325 : OR3_X1 port map( A1 => n10682, A2 => n2306, A3 => n9769, ZN => 
                           n8031);
   U24326 : OAI211_X1 port map( C1 => n4232, C2 => n4234, A => n25182, B => 
                           n4231, ZN => Ciphertext(34));
   U24327 : NAND2_X1 port map( A1 => n4229, A2 => n4236, ZN => n25182);
   U24328 : NAND2_X1 port map( A1 => n1158, A2 => n1146, ZN => n25183);
   U24329 : NAND2_X1 port map( A1 => n1890, A2 => n25469, ZN => n18785);
   U24331 : NAND2_X1 port map( A1 => n4694, A2 => n6051, ZN => n25185);
   U24332 : NAND2_X1 port map( A1 => n6449, A2 => n6450, ZN => n25186);
   U24333 : NAND2_X1 port map( A1 => n25, A2 => n25064, ZN => n25188);
   U24334 : NAND2_X1 port map( A1 => n10172, A2 => n9814, ZN => n25189);
   U24338 : INV_X1 port map( A => n11873, ZN => n25191);
   U24339 : NAND2_X1 port map( A1 => n12899, A2 => n24988, ZN => n13284);
   U24340 : OAI21_X1 port map( B1 => n1331, B2 => n14127, A => n25192, ZN => 
                           n14134);
   U24341 : NAND2_X1 port map( A1 => n1331, A2 => n25193, ZN => n25192);
   U24342 : INV_X1 port map( A => n14126, ZN => n25193);
   U24343 : XNOR2_X1 port map( A => n8311, B => n8312, ZN => n10168);
   U24344 : XNOR2_X2 port map( A => n7472, B => n7473, ZN => n9468);
   U10040 : NAND4_X2 port map( A1 => n3870, A2 => n3867, A3 => n10238, A4 => 
                           n3869, ZN => n11582);
   U3424 : OR2_X2 port map( A1 => n2962, A2 => n2963, ZN => n10891);
   U2253 : NAND3_X2 port map( A1 => n3524, A2 => n4992, A3 => n3523, ZN => 
                           n13614);
   U20847 : OAI211_X2 port map( C1 => n20235, C2 => n20173, A => n20172, B => 
                           n20171, ZN => n21998);
   U1019 : BUF_X2 port map( A => n7850, Z => n24072);
   U786 : NAND4_X2 port map( A1 => n2534, A2 => n2533, A3 => n5917, A4 => n7104
                           , ZN => n7350);
   U1457 : BUF_X1 port map( A => n16423, Z => n1329);
   U3043 : BUF_X2 port map( A => n9365, Z => n10146);
   U1115 : INV_X2 port map( A => n5522, ZN => n3374);
   U3445 : NAND2_X2 port map( A1 => n2136, A2 => n2135, ZN => n21332);
   U6597 : NAND3_X2 port map( A1 => n2622, A2 => n6215, A3 => n6214, ZN => 
                           n8935);
   U1209 : NAND2_X2 port map( A1 => n24183, A2 => n2399, ZN => n11301);
   U8646 : AND3_X2 port map( A1 => n4743, A2 => n1416, A3 => n4742, ZN => n3703
                           );
   U2551 : NAND2_X2 port map( A1 => n4803, A2 => n4799, ZN => n8691);
   U8824 : AND2_X2 port map( A1 => n10257, A2 => n10259, ZN => n10728);
   U3015 : NAND2_X2 port map( A1 => n594, A2 => n19617, ZN => n20448);
   U2385 : OAI211_X2 port map( C1 => n10679, C2 => n2984, A => n4815, B => 
                           n1401, ZN => n11717);
   U18822 : BUF_X1 port map( A => n19987, Z => n24979);
   U2113 : BUF_X1 port map( A => n15714, Z => n16471);
   U24194 : NAND3_X2 port map( A1 => n2250, A2 => n14627, A3 => n14626, ZN => 
                           n17273);
   U24157 : BUF_X1 port map( A => n13386, Z => n24507);
   U1819 : XNOR2_X2 port map( A => n15878, B => n15879, ZN => n19133);
   U1750 : XNOR2_X2 port map( A => n20978, B => n20977, ZN => n22166);
   U755 : AND2_X2 port map( A1 => n4415, A2 => n13489, ZN => n15191);
   U1232 : OAI211_X2 port map( C1 => n14586, C2 => n14747, A => n1675, B => 
                           n1674, ZN => n2285);
   U1647 : BUF_X2 port map( A => n14100, Z => n24376);
   U506 : XNOR2_X2 port map( A => n12329, B => n12328, ZN => n13350);
   U1004 : AND2_X2 port map( A1 => n22414, A2 => n22413, ZN => n23305);
   U1989 : NOR2_X2 port map( A1 => n17124, A2 => n17123, ZN => n17958);
   U9301 : NAND4_X2 port map( A1 => n13430, A2 => n13431, A3 => n14069, A4 => 
                           n13429, ZN => n14799);
   U1839 : CLKBUF_X3 port map( A => n17567, Z => n20322);
   U1879 : NAND2_X2 port map( A1 => n18799, A2 => n18798, ZN => n20062);
   U1953 : NOR2_X2 port map( A1 => n16979, A2 => n17450, ZN => n17449);
   U17681 : AND2_X2 port map( A1 => n1305, A2 => n1308, ZN => n20174);
   U709 : MUX2_X2 port map( A => n7979, B => n7978, S => n7977, Z => n8069);
   U1877 : AND2_X2 port map( A1 => n3683, A2 => n1476, ZN => n18310);
   U21457 : BUF_X1 port map( A => n21140, Z => n24406);
   U12294 : XNOR2_X2 port map( A => n5880, B => Key(34), ZN => n6952);
   U1215 : MUX2_X2 port map( A => n8712, B => n8711, S => n9985, Z => n11529);
   U185 : AND3_X2 port map( A1 => n3136, A2 => n3137, A3 => n3135, ZN => n22578
                           );
   U21731 : OAI21_X2 port map( B1 => n20623, B2 => n20622, A => n20621, ZN => 
                           n21630);
   U10086 : AND3_X2 port map( A1 => n8139, A2 => n8138, A3 => n8137, ZN => 
                           n10993);
   U576 : NAND4_X2 port map( A1 => n7547, A2 => n7544, A3 => n7546, A4 => n7545
                           , ZN => n9075);
   U510 : BUF_X1 port map( A => n17313, Z => n24543);
   U1191 : AND2_X2 port map( A1 => n3085, A2 => n4824, ZN => n15044);
   U675 : OR2_X2 port map( A1 => n9303, A2 => n9304, ZN => n10713);
   U1189 : XNOR2_X2 port map( A => n14862, B => n14863, ZN => n16219);
   U2404 : INV_X2 port map( A => n10952, ZN => n2754);
   U21492 : AND3_X2 port map( A1 => n20153, A2 => n20152, A3 => n20151, ZN => 
                           n21138);
   U17263 : OAI22_X2 port map( A1 => n13481, A2 => n13480, B1 => n13479, B2 => 
                           n13801, ZN => n14827);
   U6023 : NAND3_X2 port map( A1 => n16909, A2 => n24632, A3 => n2583, ZN => 
                           n18582);
   U3618 : BUF_X1 port map( A => n18761, Z => n19532);
   U824 : AND3_X2 port map( A1 => n17848, A2 => n17847, A3 => n17846, ZN => 
                           n19887);
   U149 : AND3_X2 port map( A1 => n17218, A2 => n17219, A3 => n17217, ZN => 
                           n18187);
   U160 : OAI211_X2 port map( C1 => n17609, C2 => n16564, A => n16563, B => 
                           n16562, ZN => n18269);
   U2006 : OAI211_X2 port map( C1 => n17054, C2 => n16935, A => n16934, B => 
                           n16933, ZN => n18067);
   U22322 : XNOR2_X1 port map( A => n11919, B => n11918, ZN => n12688);
   U1708 : AND2_X2 port map( A1 => n25130, A2 => n25131, ZN => n20231);
   U985 : OAI211_X2 port map( C1 => n16299, C2 => n15024, A => n15022, B => 
                           n24777, ZN => n17408);
   U721 : OR2_X2 port map( A1 => n5868, A2 => n5869, ZN => n7232);
   U2213 : OAI22_X2 port map( A1 => n13599, A2 => n5520, B1 => n13962, B2 => 
                           n13598, ZN => n15430);
   U2681 : BUF_X1 port map( A => n6770, Z => n6909);
   U2025 : AND4_X2 port map( A1 => n1701, A2 => n1703, A3 => n1702, A4 => n1705
                           , ZN => n18157);
   U488 : OR2_X2 port map( A1 => n19027, A2 => n19026, ZN => n20142);
   U3586 : BUF_X1 port map( A => n19310, Z => n24912);
   U23390 : NAND2_X2 port map( A1 => n15930, A2 => n25116, ZN => n17051);
   U593 : MUX2_X2 port map( A => n11021, B => n11020, S => n24640, Z => n13775)
                           ;
   U1988 : NAND3_X2 port map( A1 => n3396, A2 => n5225, A3 => n3395, ZN => 
                           n18375);
   U3659 : NOR2_X2 port map( A1 => n21354, A2 => n21353, ZN => n23817);
   U3582 : AND3_X2 port map( A1 => n9254, A2 => n9252, A3 => n9253, ZN => 
                           n10861);
   U1064 : AND3_X2 port map( A1 => n19892, A2 => n3541, A3 => n3540, ZN => 
                           n20697);
   U2100 : AND2_X2 port map( A1 => n15633, A2 => n3592, ZN => n17054);
   U5036 : XNOR2_X1 port map( A => n1759, B => n17815, ZN => n19457);
   U2142 : XNOR2_X2 port map( A => n14175, B => n14174, ZN => n17183);
   U9454 : NAND2_X2 port map( A1 => n2158, A2 => n12603, ZN => n14849);
   U2073 : OAI21_X2 port map( B1 => n16315, B2 => n16314, A => n16313, ZN => 
                           n17351);
   U2327 : XNOR2_X2 port map( A => n11514, B => n11513, ZN => n12774);
   U1147 : OR3_X2 port map( A1 => n20068, A2 => n19849, A3 => n19660, ZN => 
                           n210);
   U2005 : NAND2_X2 port map( A1 => n15876, A2 => n4614, ZN => n18294);
   U2058 : OR2_X2 port map( A1 => n6283, A2 => n6282, ZN => n7801);
   U851 : BUF_X1 port map( A => n23742, Z => n24063);
   U2922 : NAND2_X2 port map( A1 => n25133, A2 => n7530, ZN => n8790);
   U1434 : NOR2_X2 port map( A1 => n17437, A2 => n3000, ZN => n17439);
   U1810 : AND3_X2 port map( A1 => n2365, A2 => n2371, A3 => n2366, ZN => 
                           n21599);
   U505 : NAND3_X2 port map( A1 => n7411, A2 => n4277, A3 => n4278, ZN => n9015
                           );
   U606 : AND3_X2 port map( A1 => n19287, A2 => n19285, A3 => n19286, ZN => 
                           n20401);
   U2087 : MUX2_X2 port map( A => n16144, B => n16143, S => n16416, Z => n17399
                           );
   U2293 : BUF_X1 port map( A => n12560, Z => n13015);
   U14 : OR2_X2 port map( A1 => n19790, A2 => n5338, ZN => n21141);
   U1870 : AND2_X2 port map( A1 => n18898, A2 => n2844, ZN => n20126);
   U5897 : AND3_X2 port map( A1 => n24148, A2 => n9631, A3 => n9630, ZN => 
                           n11342);
   U12061 : BUF_X2 port map( A => n19353, Z => n19451);
   U523 : XNOR2_X1 port map( A => n4504, B => n14844, ZN => n16221);
   U2349 : XNOR2_X1 port map( A => n11663, B => n11664, ZN => n13061);
   U2161 : AOI21_X1 port map( B1 => n6735, B2 => n6736, A => n6734, ZN => n6867
                           );
   U1685 : NAND2_X2 port map( A1 => n493, A2 => n3454, ZN => n13521);
   U6643 : NAND2_X2 port map( A1 => n13471, A2 => n1770, ZN => n15488);
   U19056 : AND2_X2 port map( A1 => n19056, A2 => n19057, ZN => n19576);
   U18623 : AND2_X2 port map( A1 => n203, A2 => n530, ZN => n12122);
   U300 : BUF_X2 port map( A => n13360, Z => n24552);
   U1214 : INV_X1 port map( A => n10767, ZN => n11085);
   U7603 : NAND3_X2 port map( A1 => n5489, A2 => n7586, A3 => n5490, ZN => 
                           n8782);
   U556 : AND3_X2 port map( A1 => n15942, A2 => n3437, A3 => n2771, ZN => 
                           n17053);
   U21354 : BUF_X1 port map( A => n11519, Z => n25060);
   U7665 : NAND3_X2 port map( A1 => n2224, A2 => n7127, A3 => n3898, ZN => 
                           n8755);
   U1072 : BUF_X2 port map( A => n12510, Z => n12742);
   U495 : BUF_X1 port map( A => n16284, Z => n24539);
   U1984 : NOR2_X2 port map( A1 => n4565, A2 => n4562, ZN => n18579);
   U492 : AND2_X2 port map( A1 => n1115, A2 => n15551, ZN => n16649);
   U2538 : XNOR2_X2 port map( A => n9014, B => n9013, ZN => n10027);
   U1469 : NAND4_X2 port map( A1 => n5564, A2 => n5563, A3 => n5565, A4 => 
                           n20925, ZN => n21523);
   U2582 : NAND2_X2 port map( A1 => n2080, A2 => n7988, ZN => n9158);
   U472 : NAND4_X2 port map( A1 => n5206, A2 => n5209, A3 => n20196, A4 => 
                           n5205, ZN => n21043);
   U4779 : XNOR2_X1 port map( A => n20886, B => n20885, ZN => n22887);
   U804 : XNOR2_X1 port map( A => Key(54), B => Plaintext(54), ZN => n6975);
   U13601 : CLKBUF_X1 port map( A => Key(99), Z => n3164);
   U789 : CLKBUF_X1 port map( A => Key(35), Z => n4711);
   U1597 : CLKBUF_X1 port map( A => Key(157), Z => n1776);
   U1247 : CLKBUF_X1 port map( A => Key(28), Z => n2050);
   U1633 : CLKBUF_X1 port map( A => Key(152), Z => n2903);
   U12248 : XNOR2_X1 port map( A => Key(153), B => Plaintext(153), ZN => n6874)
                           ;
   U1063 : XNOR2_X1 port map( A => Key(114), B => Plaintext(114), ZN => n7026);
   U4226 : XNOR2_X1 port map( A => Key(165), B => Plaintext(165), ZN => n6775);
   U1240 : CLKBUF_X1 port map( A => Key(2), Z => n23883);
   U936 : XNOR2_X1 port map( A => n5968, B => Key(175), ZN => n6426);
   U12566 : INV_X1 port map( A => n6905, ZN => n6089);
   U426 : OR2_X1 port map( A1 => n6987, A2 => n6119, ZN => n6642);
   U792 : XNOR2_X1 port map( A => n5789, B => Key(88), ZN => n6622);
   U1131 : XNOR2_X1 port map( A => n5877, B => Key(30), ZN => n6529);
   U12308 : XNOR2_X1 port map( A => n5886, B => Key(40), ZN => n6683);
   U1249 : XNOR2_X1 port map( A => n5892, B => Key(48), ZN => n6556);
   U12384 : XNOR2_X1 port map( A => n5944, B => Key(181), ZN => n6297);
   U152 : XNOR2_X1 port map( A => n5962, B => Key(164), ZN => n6292);
   U354 : XNOR2_X1 port map( A => n6025, B => Key(15), ZN => n6519);
   U2680 : BUF_X1 port map( A => n5835, Z => n6793);
   U9169 : OR2_X1 port map( A1 => n4696, A2 => n5774, ZN => n6053);
   U282 : INV_X1 port map( A => n5794, ZN => n6722);
   U1235 : INV_X1 port map( A => n1698, ZN => n5451);
   U4806 : OR2_X1 port map( A1 => n6198, A2 => n6292, ZN => n6922);
   U5174 : OR2_X1 port map( A1 => n6519, A2 => n6179, ZN => n6518);
   U2632 : OAI21_X1 port map( B1 => n2496, B2 => n6578, A => n2495, ZN => n7533
                           );
   U343 : OAI211_X1 port map( C1 => n3763, C2 => n6940, A => n4826, B => n6681,
                           ZN => n7358);
   U2748 : AND3_X1 port map( A1 => n773, A2 => n6462, A3 => n6461, ZN => n7688)
                           ;
   U6515 : OR2_X1 port map( A1 => n6300, A2 => n6299, ZN => n7862);
   U2662 : NAND2_X1 port map( A1 => n5977, A2 => n5978, ZN => n7890);
   U7342 : OR2_X1 port map( A1 => n5270, A2 => n6472, ZN => n7917);
   U268 : OAI21_X1 port map( B1 => n6278, B2 => n6279, A => n791, ZN => n7166);
   U921 : NAND2_X1 port map( A1 => n2149, A2 => n2025, ZN => n8219);
   U88 : INV_X1 port map( A => n7638, ZN => n7918);
   U952 : OR2_X1 port map( A1 => n6417, A2 => n6416, ZN => n7857);
   U2031 : NAND2_X1 port map( A1 => n77, A2 => n703, ZN => n7255);
   U3087 : NAND2_X1 port map( A1 => n6981, A2 => n6980, ZN => n7477);
   U2629 : NOR2_X1 port map( A1 => n5648, A2 => n2836, ZN => n7973);
   U112 : OR2_X1 port map( A1 => n6022, A2 => n2166, ZN => n7595);
   U12707 : MUX2_X1 port map( A => n6270, B => n6269, S => n6136, Z => n7800);
   U2649 : INV_X1 port map( A => n7351, ZN => n7346);
   U1017 : INV_X1 port map( A => n7883, ZN => n7582);
   U566 : AND2_X1 port map( A1 => n6851, A2 => n6850, ZN => n7983);
   U1230 : INV_X1 port map( A => n8367, ZN => n24577);
   U1100 : AND2_X1 port map( A1 => n6149, A2 => n6148, ZN => n7619);
   U2643 : OR2_X1 port map( A1 => n2784, A2 => n6202, ZN => n8012);
   U2635 : NAND2_X1 port map( A1 => n1750, A2 => n4321, ZN => n7230);
   U480 : NAND3_X1 port map( A1 => n2786, A2 => n6079, A3 => n6080, ZN => n7292
                           );
   U1099 : OR2_X1 port map( A1 => n7087, A2 => n7211, ZN => n7663);
   U773 : BUF_X1 port map( A => n7211, Z => n8528);
   U13063 : INV_X1 port map( A => n7065, ZN => n7952);
   U5194 : OR2_X1 port map( A1 => n5468, A2 => n7349, ZN => n7107);
   U8484 : AND3_X1 port map( A1 => n5329, A2 => n7417, A3 => n7416, ZN => n8119
                           );
   U2566 : OR3_X1 port map( A1 => n3259, A2 => n4206, A3 => n7533, ZN => n2883)
                           ;
   U228 : OAI211_X1 port map( C1 => n7289, C2 => n7288, A => n7287, B => n7286,
                           ZN => n8798);
   U2559 : AND2_X1 port map( A1 => n3345, A2 => n6495, ZN => n8960);
   U4007 : OAI211_X1 port map( C1 => n1124, C2 => n199, A => n2092, B => n5050,
                           ZN => n8928);
   U13406 : AOI22_X1 port map( A1 => n7470, A2 => n7884, B1 => n7469, B2 => 
                           n7313, ZN => n9045);
   U1037 : OAI211_X1 port map( C1 => n7122, C2 => n7338, A => n1904, B => n7121
                           , ZN => n5179);
   U2639 : OAI211_X1 port map( C1 => n7903, C2 => n7902, A => n7899, B => n7900
                           , ZN => n8796);
   U6640 : OAI211_X1 port map( C1 => n6098, C2 => n7755, A => n2521, B => n1769
                           , ZN => n8674);
   U986 : AND2_X1 port map( A1 => n7407, A2 => n7408, ZN => n8476);
   U652 : OR2_X1 port map( A1 => n7270, A2 => n7269, ZN => n8989);
   U491 : AND2_X1 port map( A1 => n7679, A2 => n7678, ZN => n8116);
   U409 : OAI21_X1 port map( B1 => n7321, B2 => n7320, A => n2768, ZN => n8959)
                           ;
   U197 : OAI21_X1 port map( B1 => n5204, B2 => n2522, A => n5203, ZN => n5014)
                           ;
   U622 : BUF_X1 port map( A => n8627, Z => n24547);
   U6214 : OAI21_X1 port map( B1 => n7337, B2 => n7464, A => n6763, ZN => n9140
                           );
   U1951 : NAND3_X1 port map( A1 => n3082, A2 => n24205, A3 => n3083, ZN => 
                           n8682);
   U21801 : OAI21_X1 port map( B1 => n5116, B2 => n7952, A => n2490, ZN => 
                           n24413);
   U7618 : NAND4_X1 port map( A1 => n7871, A2 => n7872, A3 => n7870, A4 => 
                           n7869, ZN => n9179);
   U2553 : AND2_X1 port map( A1 => n5548, A2 => n5547, ZN => n9011);
   U13964 : XNOR2_X1 port map( A => n8345, B => n8970, ZN => n8725);
   U103 : AND3_X1 port map( A1 => n5053, A2 => n5055, A3 => n6010, ZN => n8951)
                           ;
   U2789 : NAND2_X1 port map( A1 => n472, A2 => n7194, ZN => n8772);
   U6484 : OAI211_X1 port map( C1 => n6319, C2 => n4536, A => n24652, B => 
                           n24648, ZN => n8945);
   U1079 : NAND2_X1 port map( A1 => n7072, A2 => n3814, ZN => n8923);
   U1118 : XNOR2_X1 port map( A => n3307, B => n8272, ZN => n9805);
   U2527 : XNOR2_X1 port map( A => n8743, B => n8742, ZN => n9231);
   U2433 : BUF_X1 port map( A => n9893, Z => n227);
   U2513 : XNOR2_X1 port map( A => n8957, B => n8958, ZN => n10044);
   U14249 : XNOR2_X1 port map( A => n8695, B => n8694, ZN => n9980);
   U625 : BUF_X1 port map( A => n9874, Z => n24549);
   U823 : BUF_X1 port map( A => n9856, Z => n9558);
   U289 : XNOR2_X1 port map( A => n1906, B => n8665, ZN => n10082);
   U534 : BUF_X1 port map( A => n9454, Z => n9887);
   U1306 : BUF_X1 port map( A => n9962, Z => n262);
   U10264 : MUX2_X1 port map( A => n9063, B => n5004, S => n10053, Z => n9088);
   U14990 : OAI21_X1 port map( B1 => n9865, B2 => n9864, A => n9863, ZN => 
                           n10971);
   U2625 : NAND2_X1 port map( A1 => n9540, A2 => n4594, ZN => n10751);
   U474 : AND2_X1 port map( A1 => n8144, A2 => n8143, ZN => n10405);
   U15059 : OAI21_X1 port map( B1 => n10076, B2 => n10075, A => n10074, ZN => 
                           n11063);
   U23311 : NAND3_X1 port map( A1 => n9283, A2 => n9284, A3 => n25146, ZN => 
                           n2243);
   U2445 : OAI211_X1 port map( C1 => n9880, C2 => n9879, A => n9878, B => n9877
                           , ZN => n10968);
   U494 : OAI21_X1 port map( B1 => n9265, B2 => n9899, A => n9264, ZN => n10736
                           );
   U2535 : BUF_X1 port map( A => n8934, Z => n11524);
   U1838 : OAI21_X1 port map( B1 => n2564, B2 => n3134, A => n9213, ZN => 
                           n10590);
   U1112 : OAI22_X1 port map( A1 => n8030, A2 => n9937, B1 => n8029, B2 => 
                           n24511, ZN => n10682);
   U787 : AND3_X1 port map( A1 => n9785, A2 => n9784, A3 => n9783, ZN => n11009
                           );
   U13694 : MUX2_X1 port map( A => n8064, B => n8063, S => n25464, Z => n10406)
                           ;
   U2450 : OAI211_X1 port map( C1 => n4586, C2 => n10120, A => n5356, B => 
                           n9340, ZN => n11113);
   U140 : NAND3_X1 port map( A1 => n24795, A2 => n4832, A3 => n24212, ZN => 
                           n10552);
   U3244 : NAND3_X1 port map( A1 => n9593, A2 => n698, A3 => n9594, ZN => 
                           n10486);
   U449 : NOR2_X1 port map( A1 => n9467, A2 => n9466, ZN => n10538);
   U553 : OAI21_X1 port map( B1 => n9235, B2 => n10070, A => n3705, ZN => 
                           n10846);
   U1165 : AND2_X1 port map( A1 => n1346, A2 => n1347, ZN => n11196);
   U307 : OR2_X1 port map( A1 => n3261, A2 => n3262, ZN => n11171);
   U24106 : NOR2_X1 port map( A1 => n2730, A2 => n8225, ZN => n10594);
   U1830 : NAND2_X1 port map( A1 => n10086, A2 => n2835, ZN => n11214);
   U89 : AND3_X1 port map( A1 => n9902, A2 => n9901, A3 => n9900, ZN => n10969)
                           ;
   U7787 : NAND2_X1 port map( A1 => n7440, A2 => n7439, ZN => n2306);
   U314 : AOI21_X1 port map( B1 => n5517, B2 => n5519, A => n4871, ZN => n25025
                           );
   U630 : INV_X1 port map( A => n11058, ZN => n11054);
   U3103 : INV_X1 port map( A => n10538, ZN => n2388);
   U516 : BUF_X1 port map( A => n9892, Z => n10606);
   U1770 : OR2_X1 port map( A1 => n10961, A2 => n10534, ZN => n10690);
   U776 : OAI211_X1 port map( C1 => n10836, C2 => n10829, A => n10194, B => 
                           n10193, ZN => n12255);
   U884 : OR2_X1 port map( A1 => n10619, A2 => n10618, ZN => n10627);
   U585 : OAI211_X1 port map( C1 => n10735, C2 => n10734, A => n10733, B => 
                           n10732, ZN => n12137);
   U2387 : OAI211_X1 port map( C1 => n10473, C2 => n10840, A => n10472, B => 
                           n10471, ZN => n12286);
   U2394 : NAND3_X1 port map( A1 => n5059, A2 => n5061, A3 => n5062, ZN => 
                           n11659);
   U10632 : AOI21_X1 port map( B1 => n11002, B2 => n11067, A => n11001, ZN => 
                           n12369);
   U3847 : OAI21_X1 port map( B1 => n991, B2 => n10946, A => n10945, ZN => 
                           n12226);
   U126 : NAND2_X1 port map( A1 => n4357, A2 => n10750, ZN => n12048);
   U15348 : OR2_X1 port map( A1 => n10511, A2 => n10510, ZN => n11672);
   U16041 : OAI211_X1 port map( C1 => n11529, C2 => n11528, A => n11527, B => 
                           n11526, ZN => n12323);
   U2476 : NAND2_X1 port map( A1 => n10377, A2 => n10376, ZN => n12324);
   U2555 : AOI22_X1 port map( A1 => n11035, A2 => n939, B1 => n11034, B2 => 
                           n11033, ZN => n11561);
   U352 : OAI211_X1 port map( C1 => n1358, C2 => n11166, A => n11165, B => 
                           n11164, ZN => n12065);
   U8576 : MUX2_X1 port map( A => n9910, B => n9911, S => n10497, Z => n12355);
   U10203 : NAND2_X1 port map( A1 => n4051, A2 => n4048, ZN => n12102);
   U2371 : NAND3_X1 port map( A1 => n2831, A2 => n10483, A3 => n2830, ZN => 
                           n12224);
   U1502 : AND2_X1 port map( A1 => n2763, A2 => n2762, ZN => n11607);
   U1735 : NAND2_X1 port map( A1 => n9243, A2 => n9242, ZN => n12089);
   U1006 : BUF_X1 port map( A => n12101, Z => n11897);
   U20691 : CLKBUF_X1 port map( A => n12150, Z => n25032);
   U6942 : NAND2_X1 port map( A1 => n3312, A2 => n10390, ZN => n12040);
   U2365 : NOR2_X1 port map( A1 => n11308, A2 => n11307, ZN => n11796);
   U9473 : AND2_X1 port map( A1 => n3447, A2 => n3446, ZN => n11295);
   U238 : BUF_X2 port map( A => n11556, Z => n24027);
   U464 : XNOR2_X1 port map( A => n9409, B => n9408, ZN => n12648);
   U965 : XNOR2_X1 port map( A => n11257, B => n11256, ZN => n13012);
   U1706 : XOR2_X1 port map( A => n11790, B => n11791, Z => n24476);
   U2401 : XNOR2_X1 port map( A => n11794, B => n24634, ZN => n12824);
   U7302 : XNOR2_X1 port map( A => n12172, B => n12171, ZN => n12976);
   U77 : INV_X1 port map( A => n11287, ZN => n13014);
   U16111 : XNOR2_X1 port map( A => n11612, B => n11611, ZN => n12535);
   U940 : XNOR2_X1 port map( A => n12100, B => n12099, ZN => n13341);
   U4623 : NOR2_X1 port map( A1 => n12478, A2 => n13041, ZN => n1646);
   U973 : OR2_X1 port map( A1 => n12597, A2 => n13291, ZN => n13289);
   U4284 : AOI22_X1 port map( A1 => n24443, A2 => n13264, B1 => n5361, B2 => 
                           n13267, ZN => n12832);
   U10365 : NOR2_X1 port map( A1 => n304, A2 => n24930, ZN => n13171);
   U2595 : OR2_X1 port map( A1 => n399, A2 => n13341, ZN => n13337);
   U8050 : OAI211_X1 port map( C1 => n2543, C2 => n13235, A => n2545, B => 
                           n1374, ZN => n13807);
   U2264 : OAI22_X1 port map( A1 => n12441, A2 => n5112, B1 => n5113, B2 => 
                           n12737, ZN => n14166);
   U359 : OR2_X1 port map( A1 => n11685, A2 => n5538, ZN => n13966);
   U16834 : MUX2_X1 port map( A => n12682, B => n12681, S => n13267, Z => 
                           n13788);
   U1055 : AND3_X1 port map( A1 => n12564, A2 => n12562, A3 => n12561, ZN => 
                           n396);
   U569 : NAND3_X1 port map( A1 => n12480, A2 => n12481, A3 => n12479, ZN => 
                           n14242);
   U5418 : AOI22_X1 port map( A1 => n12892, A2 => n11367, B1 => n11366, B2 => 
                           n13211, ZN => n11411);
   U326 : OR2_X1 port map( A1 => n4548, A2 => n4547, ZN => n13981);
   U9030 : AND3_X1 port map( A1 => n11331, A2 => n5748, A3 => n11330, ZN => 
                           n13951);
   U1481 : AND3_X1 port map( A1 => n12954, A2 => n12953, A3 => n2472, ZN => 
                           n14205);
   U330 : OR2_X1 port map( A1 => n12474, A2 => n12475, ZN => n4116);
   U64 : BUF_X1 port map( A => n13996, Z => n24402);
   U2269 : BUF_X1 port map( A => n13635, Z => n13935);
   U10615 : NAND2_X1 port map( A1 => n4448, A2 => n4443, ZN => n14301);
   U255 : OAI21_X1 port map( B1 => n4447, B2 => n4446, A => n24812, ZN => 
                           n13888);
   U4471 : NAND3_X1 port map( A1 => n1828, A2 => n2715, A3 => n1393, ZN => 
                           n14009);
   U159 : INV_X1 port map( A => n13965, ZN => n13962);
   U3420 : NAND3_X1 port map( A1 => n2888, A2 => n2889, A3 => n12880, ZN => 
                           n14320);
   U10334 : AND2_X1 port map( A1 => n12487, A2 => n12488, ZN => n14245);
   U17162 : NOR2_X1 port map( A1 => n13989, A2 => n13982, ZN => n13985);
   U119 : BUF_X2 port map( A => n14851, Z => n24572);
   U1329 : INV_X1 port map( A => n13744, ZN => n13526);
   U212 : NAND2_X1 port map( A1 => n11224, A2 => n2929, ZN => n14156);
   U2222 : AND2_X1 port map( A1 => n13444, A2 => n14060, ZN => n14419);
   U373 : AOI21_X1 port map( B1 => n4129, B2 => n4131, A => n13827, ZN => 
                           n15507);
   U3364 : NAND2_X1 port map( A1 => n5708, A2 => n24827, ZN => n15165);
   U1052 : AOI22_X1 port map( A1 => n13855, A2 => n13856, B1 => n13857, B2 => 
                           n14078, ZN => n14558);
   U1533 : NAND2_X1 port map( A1 => n1966, A2 => n24095, ZN => n15483);
   U65 : NAND2_X1 port map( A1 => n59, A2 => n684, ZN => n14993);
   U2192 : OAI211_X1 port map( C1 => n2658, C2 => n13255, A => n13254, B => 
                           n2657, ZN => n14952);
   U235 : NOR2_X1 port map( A1 => n13314, A2 => n13315, ZN => n15273);
   U6904 : NAND3_X1 port map( A1 => n2503, A2 => n2507, A3 => n2502, ZN => 
                           n15177);
   U486 : NAND3_X1 port map( A1 => n13897, A2 => n13899, A3 => n13898, ZN => 
                           n15326);
   U5467 : AND2_X1 port map( A1 => n4593, A2 => n4592, ZN => n14500);
   U2186 : AND2_X1 port map( A1 => n13992, A2 => n1112, ZN => n14788);
   U8318 : AND3_X1 port map( A1 => n13369, A2 => n13368, A3 => n13367, ZN => 
                           n15203);
   U9707 : AND2_X1 port map( A1 => n3538, A2 => n3536, ZN => n14977);
   U3879 : NAND3_X1 port map( A1 => n13751, A2 => n1026, A3 => n1025, ZN => 
                           n15464);
   U18277 : XNOR2_X1 port map( A => n14976, B => n912, ZN => n14978);
   U33 : XNOR2_X1 port map( A => n14422, B => n14421, ZN => n16427);
   U597 : XNOR2_X1 port map( A => n14771, B => n14772, ZN => n16016);
   U2164 : XNOR2_X1 port map( A => n14228, B => n14229, ZN => n16176);
   U18163 : XNOR2_X1 port map( A => n14804, B => n14803, ZN => n16491);
   U17181 : INV_X1 port map( A => n15019, ZN => n15499);
   U374 : XNOR2_X1 port map( A => n15337, B => n15336, ZN => n15697);
   U2176 : XNOR2_X1 port map( A => n15214, B => n15213, ZN => n16312);
   U9437 : XNOR2_X1 port map( A => n3308, B => n14047, ZN => n16367);
   U1461 : XNOR2_X1 port map( A => n13738, B => n13737, ZN => n15646);
   U2127 : XNOR2_X1 port map( A => n4204, B => n4205, ZN => n2253);
   U2146 : BUF_X1 port map( A => n15707, Z => n16442);
   U2173 : XNOR2_X1 port map( A => n15288, B => n15289, ZN => n16051);
   U1086 : BUF_X1 port map( A => n14350, Z => n16177);
   U283 : INV_X1 port map( A => n15545, ZN => n16469);
   U1253 : XNOR2_X1 port map( A => n14736, B => n14735, ZN => n16102);
   U11601 : XNOR2_X1 port map( A => n5494, B => n15323, ZN => n15695);
   U1450 : INV_X1 port map( A => n3779, ZN => n3544);
   U18434 : XNOR2_X1 port map( A => n15206, B => n15207, ZN => n15557);
   U446 : BUF_X1 port map( A => n15637, Z => n15972);
   U2097 : MUX2_X1 port map( A => n15475, B => n15474, S => n15950, Z => n15872
                           );
   U1961 : AND2_X1 port map( A1 => n17436, A2 => n16429, ZN => n17442);
   U1323 : AND4_X1 port map( A1 => n15598, A2 => n15597, A3 => n15595, A4 => 
                           n15596, ZN => n1139);
   U2078 : AND3_X1 port map( A1 => n16446, A2 => n16444, A3 => n16445, ZN => 
                           n1653);
   U4506 : AND2_X1 port map( A1 => n5581, A2 => n15650, ZN => n17305);
   U42 : AND2_X1 port map( A1 => n16810, A2 => n16808, ZN => n17076);
   U46 : NAND2_X1 port map( A1 => n1791, A2 => n1832, ZN => n17389);
   U8230 : AND3_X1 port map( A1 => n2648, A2 => n2649, A3 => n2650, ZN => 
                           n17336);
   U4689 : NOR2_X1 port map( A1 => n15744, A2 => n16328, ZN => n17624);
   U378 : NAND2_X1 port map( A1 => n1245, A2 => n4575, ZN => n17304);
   U10488 : AND2_X1 port map( A1 => n4420, A2 => n4416, ZN => n17114);
   U870 : OR2_X1 port map( A1 => n3576, A2 => n15589, ZN => n16731);
   U688 : NAND2_X1 port map( A1 => n15601, A2 => n1673, ZN => n16546);
   U2057 : AND2_X1 port map( A1 => n15683, A2 => n15682, ZN => n17319);
   U274 : BUF_X2 port map( A => n17062, Z => n24585);
   U19554 : MUX2_X1 port map( A => n17122, B => n17121, S => n17120, Z => 
                           n17123);
   U83 : OR2_X1 port map( A1 => n16288, A2 => n2701, ZN => n17014);
   U769 : NAND2_X1 port map( A1 => n3005, A2 => n3003, ZN => n18200);
   U2000 : NAND3_X1 port map( A1 => n1133, A2 => n17070, A3 => n1070, ZN => 
                           n18599);
   U3556 : AND3_X1 port map( A1 => n24594, A2 => n16992, A3 => n16993, ZN => 
                           n17959);
   U1163 : INV_X1 port map( A => n3706, ZN => n24568);
   U6441 : OR2_X1 port map( A1 => n1625, A2 => n1623, ZN => n17681);
   U441 : BUF_X1 port map( A => n17933, Z => n24536);
   U1383 : NAND2_X1 port map( A1 => n24174, A2 => n16853, ZN => n18669);
   U1083 : BUF_X1 port map( A => n18589, Z => n24565);
   U11658 : OAI21_X1 port map( B1 => n16615, B2 => n16514, A => n5555, ZN => 
                           n18214);
   U429 : NAND3_X1 port map( A1 => n16900, A2 => n4613, A3 => n4612, ZN => 
                           n18540);
   U19959 : XNOR2_X1 port map( A => n18098, B => n17768, ZN => n18573);
   U710 : AND2_X1 port map( A1 => n1253, A2 => n1252, ZN => n17819);
   U388 : XNOR2_X1 port map( A => n17930, B => n17929, ZN => n19499);
   U1932 : BUF_X1 port map( A => n4748, Z => n3296);
   U211 : XNOR2_X1 port map( A => n17885, B => n17884, ZN => n19466);
   U425 : XNOR2_X1 port map( A => n670, B => n18148, ZN => n19105);
   U19901 : XNOR2_X1 port map( A => n17703, B => n17702, ZN => n19357);
   U1958 : CLKBUF_X1 port map( A => n18914, Z => n17559);
   U1956 : XNOR2_X1 port map( A => n17879, B => n17878, ZN => n19472);
   U11003 : XNOR2_X1 port map( A => n18013, B => n18012, ZN => n19210);
   U1318 : BUF_X1 port map( A => n19015, Z => n19393);
   U903 : XNOR2_X1 port map( A => n4086, B => n1408, ZN => n19255);
   U154 : BUF_X1 port map( A => n18690, Z => n19412);
   U16146 : OR2_X1 port map( A1 => n19412, A2 => n19413, ZN => n18783);
   U5855 : MUX2_X1 port map( A => n18775, B => n18774, S => n19186, Z => n20470
                           );
   U1146 : AND3_X1 port map( A1 => n18167, A2 => n18168, A3 => n1426, ZN => 
                           n3480);
   U1872 : NAND4_X1 port map( A1 => n19089, A2 => n3668, A3 => n19085, A4 => 
                           n19086, ZN => n20268);
   U1878 : AND2_X1 port map( A1 => n19137, A2 => n19136, ZN => n20264);
   U11719 : NAND3_X1 port map( A1 => n19175, A2 => n19174, A3 => n5617, ZN => 
                           n20216);
   U8158 : OAI211_X1 port map( C1 => n4580, C2 => n19167, A => n4579, B => 
                           n4578, ZN => n20217);
   U25 : AND3_X1 port map( A1 => n115, A2 => n18790, A3 => n114, ZN => n20590);
   U7103 : OAI211_X1 port map( C1 => n1990, C2 => n19406, A => n18783, B => 
                           n1987, ZN => n20617);
   U24200 : NAND2_X1 port map( A1 => n1000, A2 => n1003, ZN => n20480);
   U4115 : AND2_X1 port map( A1 => n19224, A2 => n5681, ZN => n20193);
   U201 : OAI21_X1 port map( B1 => n18093, B2 => n18092, A => n18091, ZN => 
                           n20557);
   U20797 : NOR2_X1 port map( A1 => n18964, A2 => n18963, ZN => n19991);
   U6 : BUF_X1 port map( A => n20484, Z => n20486);
   U1144 : NAND2_X1 port map( A1 => n1822, A2 => n519, ZN => n20309);
   U1571 : NAND2_X1 port map( A1 => n19350, A2 => n20390, ZN => n20395);
   U1392 : OR2_X1 port map( A1 => n17940, A2 => n17939, ZN => n17943);
   U1388 : BUF_X2 port map( A => n17943, Z => n20100);
   U20958 : AOI22_X1 port map( A1 => n19740, A2 => n25397, B1 => n19259, B2 => 
                           n20425, ZN => n19260);
   U15 : AND3_X1 port map( A1 => n3430, A2 => n5541, A3 => n3429, ZN => n1381);
   U13641 : AND3_X1 port map( A1 => n3466, A2 => n3732, A3 => n19954, ZN => 
                           n3465);
   U1828 : OAI21_X1 port map( B1 => n19657, B2 => n19197, A => n19196, ZN => 
                           n20780);
   U17356 : OR2_X1 port map( A1 => n20017, A2 => n24950, ZN => n3041);
   U7106 : AND3_X1 port map( A1 => n1992, A2 => n1993, A3 => n1991, ZN => 
                           n21596);
   U1827 : OAI21_X1 port map( B1 => n1521, B2 => n200, A => n19118, ZN => 
                           n20826);
   U21385 : MUX2_X1 port map( A => n19968, B => n19967, S => n20127, Z => 
                           n19970);
   U22667 : NAND2_X1 port map( A1 => n20876, A2 => n20873, ZN => n21600);
   U20821 : NAND2_X1 port map( A1 => n18996, A2 => n18997, ZN => n21679);
   U21567 : NOR2_X1 port map( A1 => n20295, A2 => n20294, ZN => n21492);
   U1274 : BUF_X1 port map( A => n20585, Z => n24353);
   U8563 : AND3_X1 port map( A1 => n20119, A2 => n2874, A3 => n2873, ZN => 
                           n21601);
   U1806 : NOR2_X1 port map( A1 => n21013, A2 => n21012, ZN => n21687);
   U11 : AND3_X1 port map( A1 => n19824, A2 => n2916, A3 => n19090, ZN => 
                           n21587);
   U1776 : XNOR2_X1 port map( A => n20342, B => n4169, ZN => n4273);
   U1407 : XNOR2_X1 port map( A => n19935, B => n19934, ZN => n22226);
   U568 : XNOR2_X1 port map( A => n19795, B => n19796, ZN => n22689);
   U8061 : BUF_X1 port map( A => n21872, Z => n22426);
   U1755 : BUF_X1 port map( A => n20845, Z => n23571);
   U947 : BUF_X2 port map( A => n24510, Z => n24559);
   U19358 : NOR2_X1 port map( A1 => n21791, A2 => n22231, ZN => n21794);
   U5748 : NOR2_X1 port map( A1 => n22176, A2 => n24396, ZN => n21802);
   U1740 : XNOR2_X1 port map( A => n21256, B => n21257, ZN => n2397);
   U1002 : NOR2_X1 port map( A1 => n4437, A2 => n22244, ZN => n22184);
   U1715 : MUX2_X1 port map( A => n22183, B => n22182, S => n22181, Z => n23672
                           );
   U362 : OR2_X1 port map( A1 => n996, A2 => n998, ZN => n997);
   U19984 : OAI211_X1 port map( C1 => n4362, C2 => n22200, A => n4361, B => 
                           n4359, ZN => n23727);
   U7250 : MUX2_X1 port map( A => n22474, B => n22473, S => n22612, Z => n23104
                           );
   U1724 : AOI21_X1 port map( B1 => n21804, B2 => n21805, A => n21803, ZN => 
                           n23768);
   U254 : INV_X1 port map( A => n23911, ZN => n23926);
   U3335 : AND2_X1 port map( A1 => n2296, A2 => n2297, ZN => n23645);
   U1234 : BUF_X1 port map( A => n23129, Z => n23143);
   U22990 : NOR2_X1 port map( A1 => n23672, A2 => n23671, ZN => n23658);
   U1707 : BUF_X2 port map( A => n21863, Z => n23879);
   U24347 : NAND2_X1 port map( A1 => n1799, A2 => n22865, ZN => n23411);
   U976 : NOR2_X1 port map( A1 => n840, A2 => n22112, ZN => n25071);
   U8867 : NAND2_X1 port map( A1 => n23650, A2 => n23612, ZN => n1619);
   U4793 : OR2_X1 port map( A1 => n5090, A2 => n24334, ZN => n4235);
   U23081 : MUX2_X1 port map( A => n22345, B => n22344, S => n23166, Z => 
                           n22347);
   U1342 : CLKBUF_X1 port map( A => Key(182), Z => n2058);
   U2718 : BUF_X1 port map( A => Key(175), Z => n1831);
   U1346 : BUF_X1 port map( A => Key(48), Z => n768);
   U1348 : BUF_X2 port map( A => Key(136), Z => n859);
   U793 : CLKBUF_X1 port map( A => Key(40), Z => n1920);
   U1595 : BUF_X1 port map( A => Key(105), Z => n1875);
   U8283 : NAND2_X1 port map( A1 => n24203, A2 => n7930, ZN => n7445);
   U6046 : BUF_X1 port map( A => n7065, Z => n7476);
   U1335 : INV_X1 port map( A => n7662, ZN => n269);
   U8027 : INV_X1 port map( A => n7757, ZN => n2522);
   U322 : NOR2_X2 port map( A1 => n7747, A2 => n2402, ZN => n3588);
   U125 : OAI21_X1 port map( B1 => n7998, B2 => n7997, A => n7996, ZN => n8779)
                           ;
   U2565 : NAND3_X1 port map( A1 => n2554, A2 => n2553, A3 => n2551, ZN => 
                           n8818);
   U13808 : INV_X1 port map( A => n9886, ZN => n9563);
   U6161 : INV_X2 port map( A => n9694, ZN => n4993);
   U1223 : INV_X2 port map( A => n9788, ZN => n24575);
   U1221 : INV_X2 port map( A => n9786, ZN => n10088);
   U2452 : NAND4_X1 port map( A1 => n8887, A2 => n8886, A3 => n9436, A4 => 
                           n8888, ZN => n8934);
   U168 : NAND2_X1 port map( A1 => n9088, A2 => n9087, ZN => n10571);
   U533 : XNOR2_X1 port map( A => n10270, B => n10269, ZN => n12459);
   U8208 : NOR2_X1 port map( A1 => n13266, A2 => n13264, ZN => n12830);
   U1482 : AOI21_X1 port map( B1 => n13322, B2 => n13321, A => n13320, ZN => 
                           n14230);
   U1134 : OAI211_X1 port map( C1 => n13051, C2 => n25408, A => n12492, B => 
                           n12491, ZN => n14244);
   U1643 : INV_X1 port map( A => n14852, ZN => n14415);
   U2227 : CLKBUF_X1 port map( A => n12772, Z => n14179);
   U665 : OAI211_X1 port map( C1 => n13575, C2 => n13826, A => n13896, B => 
                           n13574, ZN => n15034);
   U2189 : AND2_X1 port map( A1 => n5252, A2 => n5253, ZN => n13906);
   U23574 : OR2_X1 port map( A1 => n13881, A2 => n13882, ZN => n15393);
   U53 : BUF_X1 port map( A => n14499, Z => n16118);
   U18820 : AND3_X1 port map( A1 => n15818, A2 => n16366, A3 => n15817, ZN => 
                           n17485);
   U11872 : MUX2_X1 port map( A => n16790, B => n16789, S => n17131, Z => 
                           n18098);
   U14863 : INV_X1 port map( A => n2333, ZN => n20388);
   U1920 : CLKBUF_X1 port map( A => n18762, Z => n19534);
   U3472 : NAND2_X1 port map( A1 => n19101, A2 => n19102, ZN => n20517);
   U10572 : NAND2_X1 port map( A1 => n3470, A2 => n24247, ZN => n20422);
   U1284 : NAND3_X1 port map( A1 => n171, A2 => n20229, A3 => n170, ZN => 
                           n21694);
   U299 : INV_X1 port map( A => n21467, ZN => n22969);
   U1756 : BUF_X1 port map( A => n21380, Z => n22456);
   U1296 : NAND3_X1 port map( A1 => n535, A2 => n21294, A3 => n534, ZN => 
                           n24972);
   U620 : NAND2_X1 port map( A1 => n22378, A2 => n22377, ZN => n23937);
   U4072 : NAND2_X1 port map( A1 => n3035, A2 => n21916, ZN => n23206);
   U1157 : NOR2_X1 port map( A1 => n22405, A2 => n22404, ZN => n23293);
   U1098 : AND3_X2 port map( A1 => n13511, A2 => n13510, A3 => n13509, ZN => 
                           n14880);
   U319 : MUX2_X2 port map( A => n6962, B => n6961, S => n6960, Z => n7423);
   U2494 : BUF_X2 port map( A => n9918, Z => n9355);
   U2011 : AND2_X2 port map( A1 => n6482, A2 => n839, ZN => n512);
   U518 : BUF_X2 port map( A => n7941, Z => n9276);
   U24 : BUF_X2 port map( A => n18730, Z => n19479);
   U2359 : AND3_X2 port map( A1 => n201, A2 => n9293, A3 => n547, ZN => n12365)
                           ;
   U672 : OR2_X2 port map( A1 => n7690, A2 => n7692, ZN => n8315);
   U204 : AOI21_X2 port map( B1 => n10132, B2 => n10133, A => n10131, ZN => 
                           n10559);
   U8827 : NAND2_X2 port map( A1 => n6205, A2 => n5450, ZN => n8014);
   U10047 : AND3_X2 port map( A1 => n3874, A2 => n3875, A3 => n3873, ZN => 
                           n13417);
   U684 : NAND3_X2 port map( A1 => n7394, A2 => n2893, A3 => n7393, ZN => n8375
                           );
   U360 : OR2_X2 port map( A1 => n6433, A2 => n6432, ZN => n8316);
   U1266 : XNOR2_X2 port map( A => n7780, B => n7779, ZN => n9934);
   U828 : AND3_X2 port map( A1 => n9413, A2 => n9412, A3 => n2778, ZN => n11084
                           );
   U1175 : OAI21_X2 port map( B1 => n17021, B2 => n17022, A => n17020, ZN => 
                           n18325);
   U266 : NAND2_X2 port map( A1 => n9258, A2 => n10047, ZN => n10740);
   U13297 : OR2_X2 port map( A1 => n7301, A2 => n7300, ZN => n8147);
   U2141 : BUF_X2 port map( A => n15549, Z => n16063);
   U2242 : NOR2_X2 port map( A1 => n300, A2 => n14063, ZN => n3533);
   U6701 : NAND3_X2 port map( A1 => n24276, A2 => n24277, A3 => n6029, ZN => 
                           n7602);
   U865 : NAND2_X2 port map( A1 => n3431, A2 => n3433, ZN => n18350);
   U2655 : OR2_X2 port map( A1 => n6249, A2 => n6248, ZN => n7734);
   U2590 : OR2_X2 port map( A1 => n24578, A2 => n7735, ZN => n7645);
   U3031 : AND2_X2 port map( A1 => n9762, A2 => n9620, ZN => n9760);
   U1077 : OR2_X2 port map( A1 => n16407, A2 => n802, ZN => n16962);
   U1049 : AND3_X2 port map( A1 => n5695, A2 => n2061, A3 => n6181, ZN => n7762
                           );
   U2028 : BUF_X2 port map( A => n15774, Z => n16302);
   U1995 : AND2_X2 port map( A1 => n3392, A2 => n3390, ZN => n17970);
   U607 : BUF_X2 port map( A => n6236, Z => n24051);
   U1979 : NAND2_X2 port map( A1 => n16977, A2 => n4246, ZN => n18562);
   U20750 : OR2_X2 port map( A1 => n25039, A2 => n17335, ZN => n3818);
   U12974 : OR2_X2 port map( A1 => n6761, A2 => n6760, ZN => n8427);
   U23694 : XNOR2_X2 port map( A => n11400, B => n11399, ZN => n12785);
   U1222 : OAI211_X2 port map( C1 => n1510, C2 => n1512, A => n1511, B => 
                           n16350, ZN => n17734);
   U1109 : XNOR2_X2 port map( A => n8260, B => n8259, ZN => n10176);
   U603 : BUF_X1 port map( A => n6236, Z => n24050);
   U720 : NAND4_X2 port map( A1 => n5986, A2 => n2593, A3 => n5987, A4 => n5988
                           , ZN => n7323);
   U4455 : NAND3_X2 port map( A1 => n16238, A2 => n16237, A3 => n16239, ZN => 
                           n17208);
   U1127 : BUF_X2 port map( A => n11217, Z => n233);
   U2277 : OR2_X2 port map( A1 => n3631, A2 => n3632, ZN => n14089);
   U117 : OR2_X2 port map( A1 => n5820, A2 => n5821, ZN => n7585);
   U1025 : AND4_X2 port map( A1 => n3079, A2 => n9968, A3 => n9967, A4 => n9966
                           , ZN => n11268);
   U414 : AND2_X2 port map( A1 => n6056, A2 => n6055, ZN => n8021);
   U8534 : MUX2_X2 port map( A => n18595, B => n18594, S => n19419, Z => n20618
                           );
   U23264 : NOR2_X2 port map( A1 => n23050, A2 => n23040, ZN => n23055);
   U572 : XNOR2_X2 port map( A => Key(128), B => Plaintext(128), ZN => n6072);
   U217 : AND2_X2 port map( A1 => n7249, A2 => n7248, ZN => n8460);
   U19699 : OAI211_X2 port map( C1 => n5406, C2 => n17429, A => n17428, B => 
                           n17427, ZN => n18515);
   U2463 : OR2_X2 port map( A1 => n9843, A2 => n24085, ZN => n9340);
   U386 : NAND2_X2 port map( A1 => n19143, A2 => n19144, ZN => n20411);
   U2443 : AND3_X2 port map( A1 => n9396, A2 => n9395, A3 => n9394, ZN => 
                           n10730);
   U1218 : XNOR2_X2 port map( A => Key(0), B => Plaintext(0), ZN => n6455);
   U242 : NAND2_X2 port map( A1 => n40, A2 => n1232, ZN => n17413);
   U8893 : NAND3_X2 port map( A1 => n24740, A2 => n10101, A3 => n4258, ZN => 
                           n11216);
   U1045 : NOR2_X2 port map( A1 => n14515, A2 => n14514, ZN => n15063);
   U532 : NOR2_X2 port map( A1 => n1286, A2 => n1285, ZN => n16859);
   U10626 : OR2_X2 port map( A1 => n7624, A2 => n7623, ZN => n8458);
   U707 : BUF_X2 port map( A => n6267, Z => n6164);
   U843 : BUF_X2 port map( A => n16405, Z => n24061);
   U1303 : BUF_X2 port map( A => n9255, Z => n260);
   U2291 : BUF_X2 port map( A => n12576, Z => n13336);
   U1513 : NOR2_X2 port map( A1 => n10209, A2 => n10208, ZN => n10884);
   U12150 : XNOR2_X2 port map( A => Key(60), B => Plaintext(60), ZN => n6964);
   U648 : NAND2_X2 port map( A1 => n3628, A2 => n3629, ZN => n17312);
   U2558 : AND2_X2 port map( A1 => n24629, A2 => n9940, ZN => n10800);
   U11897 : NOR2_X2 port map( A1 => n13047, A2 => n13046, ZN => n13824);
   U2736 : NAND2_X2 port map( A1 => n25185, A2 => n4697, ZN => n7573);
   U2348 : NAND2_X2 port map( A1 => n5816, A2 => n3365, ZN => n8596);
   U264 : MUX2_X2 port map( A => n16387, B => n16386, S => n15655, Z => n16963)
                           ;
   U1411 : BUF_X2 port map( A => n18812, Z => n19384);
   U15557 : MUX2_X2 port map( A => n10909, B => n10908, S => n10907, Z => 
                           n12183);
   U428 : OR2_X2 port map( A1 => n7927, A2 => n7928, ZN => n5607);
   U934 : XNOR2_X2 port map( A => n5844, B => Key(160), ZN => n6912);
   U948 : OR2_X2 port map( A1 => n7050, A2 => n7051, ZN => n8457);
   U39 : AND3_X2 port map( A1 => n16263, A2 => n16265, A3 => n16264, ZN => 
                           n17824);
   U3105 : OAI21_X2 port map( B1 => n14256, B2 => n13927, A => n13382, ZN => 
                           n14694);
   U315 : CLKBUF_X3 port map( A => n14304, Z => n24588);
   U11400 : INV_X2 port map( A => n6375, ZN => n6906);
   U5430 : OR2_X2 port map( A1 => n13984, A2 => n13922, ZN => n1899);
   U2781 : BUF_X2 port map( A => n6534, Z => n24592);
   U461 : BUF_X1 port map( A => n9481, Z => n10008);
   U1514 : INV_X1 port map( A => n10079, ZN => n9507);
   U9716 : NAND3_X1 port map( A1 => n9607, A2 => n9605, A3 => n9606, ZN => 
                           n10613);
   U1788 : OR2_X1 port map( A1 => n9826, A2 => n9825, ZN => n10952);
   U219 : BUF_X2 port map( A => n10534, Z => n11151);
   U279 : AND3_X1 port map( A1 => n31, A2 => n1893, A3 => n1894, ZN => n13569);
   U964 : NAND3_X1 port map( A1 => n13630, A2 => n13631, A3 => n176, ZN => 
                           n15436);
   U18259 : XNOR2_X1 port map( A => n14942, B => n14941, ZN => n16447);
   U8921 : AND2_X1 port map( A1 => n24741, A2 => n15623, ZN => n16932);
   U11851 : AOI21_X2 port map( B1 => n16013, B2 => n16012, A => n16011, ZN => 
                           n16021);
   U1888 : NAND2_X1 port map( A1 => n1120, A2 => n1121, ZN => n20055);
   U1861 : AND3_X1 port map( A1 => n18780, A2 => n18781, A3 => n18779, ZN => 
                           n20060);
   U9 : BUF_X2 port map( A => n14435, Z => n24556);
   U21 : MUX2_X1 port map( A => n10402, B => n10401, S => n25250, Z => n11640);
   U23 : BUF_X2 port map( A => n10147, Z => n25206);
   U29 : INV_X2 port map( A => n1629, ZN => n25242);
   U31 : XNOR2_X2 port map( A => n18430, B => n18429, ZN => n18505);
   U38 : OR2_X2 port map( A1 => n19661, A2 => n19850, ZN => n24288);
   U44 : NAND2_X2 port map( A1 => n25290, A2 => n18988, ZN => n20136);
   U47 : BUF_X2 port map( A => n20249, Z => n24077);
   U68 : AND2_X2 port map( A1 => n1556, A2 => n209, ZN => n20345);
   U71 : BUF_X2 port map( A => n10245, Z => n10648);
   U72 : OR2_X2 port map( A1 => n1983, A2 => n16219, ZN => n15925);
   U75 : OAI21_X2 port map( B1 => n8320, B2 => n2404, A => n1463, ZN => n8551);
   U79 : BUF_X2 port map( A => n22809, Z => n25241);
   U84 : OAI211_X1 port map( C1 => n20184, C2 => n20186, A => n19663, B => 
                           n2339, ZN => n21311);
   U87 : NAND3_X1 port map( A1 => n20490, A2 => n24274, A3 => n20489, ZN => 
                           n21027);
   U92 : AOI211_X1 port map( C1 => n21289, C2 => n22686, A => n5770, B => 
                           n21817, ZN => n21291);
   U113 : INV_X1 port map( A => n13643, ZN => n24589);
   U128 : NAND2_X1 port map( A1 => n16308, A2 => n16307, ZN => n17012);
   U131 : BUF_X1 port map( A => n15905, Z => n15904);
   U132 : INV_X1 port map( A => n15905, ZN => n17180);
   U136 : AOI22_X1 port map( A1 => n3127, A2 => n20562, B1 => n20093, B2 => 
                           n25221, ZN => n19876);
   U150 : OAI211_X1 port map( C1 => n13614, C2 => n25247, A => n12823, B => 
                           n12822, ZN => n14900);
   U153 : NOR2_X1 port map( A1 => n13788, A2 => n13785, ZN => n14140);
   U161 : BUF_X2 port map( A => n9931, Z => n25217);
   U173 : OAI211_X2 port map( C1 => n3119, C2 => n10222, A => n10766, B => 
                           n10221, ZN => n12313);
   U177 : BUF_X1 port map( A => n13012, Z => n25198);
   U203 : OAI21_X2 port map( B1 => n300, B2 => n12592, A => n25549, ZN => 
                           n15168);
   U206 : AOI21_X2 port map( B1 => n14103, B2 => n4877, A => n4876, ZN => 
                           n25394);
   U225 : NOR2_X2 port map( A1 => n15832, A2 => n151, ZN => n25472);
   U231 : AND3_X2 port map( A1 => n24788, A2 => n24787, A3 => n24786, ZN => 
                           n16572);
   U236 : AND3_X2 port map( A1 => n638, A2 => n16632, A3 => n16631, ZN => 
                           n25390);
   U237 : OAI211_X2 port map( C1 => n17169, C2 => n2430, A => n17168, B => n514
                           , ZN => n25380);
   U251 : XNOR2_X2 port map( A => n20642, B => n20213, ZN => n21839);
   U256 : NAND4_X2 port map( A1 => n15727, A2 => n15730, A3 => n15728, A4 => 
                           n15729, ZN => n17296);
   U258 : OAI21_X2 port map( B1 => n22732, B2 => n22731, A => n22730, ZN => 
                           n23478);
   U262 : BUF_X2 port map( A => n18396, Z => n25194);
   U271 : NAND4_X1 port map( A1 => n16880, A2 => n16881, A3 => n16882, A4 => 
                           n16879, ZN => n18396);
   U276 : OAI211_X2 port map( C1 => n1409, C2 => n16712, A => n27, B => n26, ZN
                           => n18633);
   U277 : OAI21_X2 port map( B1 => n2349, B2 => n2352, A => n2348, ZN => n5971)
                           ;
   U278 : AND4_X2 port map( A1 => n5424, A2 => n5425, A3 => n24533, A4 => n5423
                           , ZN => n21414);
   U297 : XNOR2_X2 port map( A => Key(71), B => Plaintext(71), ZN => n6578);
   U305 : NAND4_X2 port map( A1 => n3991, A2 => n3992, A3 => n15684, A4 => 
                           n15685, ZN => n18080);
   U308 : AOI21_X2 port map( B1 => n1268, B2 => n12662, A => n1267, ZN => 
                           n13488);
   U309 : BUF_X2 port map( A => n16405, Z => n24062);
   U311 : NAND3_X2 port map( A1 => n2758, A2 => n2759, A3 => n5901, ZN => n8412
                           );
   U324 : MUX2_X2 port map( A => n22170, B => n22071, S => n21712, Z => n22075)
                           ;
   U327 : NAND3_X2 port map( A1 => n6043, A2 => n6042, A3 => n6041, ZN => n7597
                           );
   U342 : OR2_X2 port map( A1 => n7632, A2 => n7631, ZN => n8706);
   U350 : XNOR2_X2 port map( A => Plaintext(64), B => Key(64), ZN => n6575);
   U358 : MUX2_X2 port map( A => n6349, B => n6348, S => n6347, Z => n7809);
   U365 : XNOR2_X2 port map( A => Key(79), B => Plaintext(79), ZN => n6732);
   U366 : XNOR2_X2 port map( A => n8254, B => n8253, ZN => n10186);
   U371 : XNOR2_X2 port map( A => n21566, B => n21565, ZN => n22958);
   U389 : OAI21_X2 port map( B1 => n6672, B2 => n6671, A => n6670, ZN => n7991)
                           ;
   U390 : NAND2_X2 port map( A1 => n2858, A2 => n3056, ZN => n8754);
   U394 : OR2_X2 port map( A1 => n28, A2 => n6786, ZN => n7977);
   U395 : XNOR2_X2 port map( A => n5862, B => Key(28), ZN => n6532);
   U397 : BUF_X2 port map( A => n13305, Z => n13307);
   U406 : XNOR2_X2 port map( A => n11697, B => n11696, ZN => n13305);
   U408 : BUF_X2 port map( A => n19762, Z => n25195);
   U424 : XNOR2_X1 port map( A => n18391, B => n18392, ZN => n19762);
   U434 : CLKBUF_X1 port map( A => n14338, Z => n25196);
   U435 : BUF_X2 port map( A => n14338, Z => n25197);
   U440 : NOR2_X1 port map( A1 => n13503, A2 => n13504, ZN => n14338);
   U448 : XNOR2_X2 port map( A => n5870, B => Key(46), ZN => n6956);
   U456 : XNOR2_X2 port map( A => n9006, B => n9005, ZN => n10026);
   U460 : AOI22_X2 port map( A1 => n11454, A2 => n24973, B1 => n14289, B2 => 
                           n11453, ZN => n14685);
   U463 : NAND2_X2 port map( A1 => n24807, A2 => n818, ZN => n20134);
   U465 : OR2_X2 port map( A1 => n9561, A2 => n25307, ZN => n10907);
   U473 : BUF_X1 port map( A => n13012, Z => n25199);
   U504 : XNOR2_X2 port map( A => n17708, B => n18493, ZN => n19452);
   U513 : BUF_X2 port map( A => n6414, Z => n6695);
   U514 : BUF_X2 port map( A => n11350, Z => n13206);
   U519 : XNOR2_X2 port map( A => n13914, B => n13913, ZN => n16397);
   U525 : XNOR2_X2 port map( A => n5872, B => Key(55), ZN => n6690);
   U526 : NAND2_X2 port map( A1 => n6614, A2 => n6613, ZN => n7781);
   U537 : XNOR2_X2 port map( A => n2408, B => n2407, ZN => n223);
   U547 : MUX2_X2 port map( A => n19096, B => n19095, S => n19380, Z => n20515)
                           ;
   U552 : OAI21_X2 port map( B1 => n4741, B2 => n13227, A => n3351, ZN => 
                           n13918);
   U563 : OAI211_X2 port map( C1 => n14298, C2 => n14297, A => n14295, B => 
                           n24146, ZN => n14634);
   U565 : BUF_X1 port map( A => n17215, Z => n25200);
   U571 : BUF_X2 port map( A => n17215, Z => n25201);
   U578 : AOI22_X1 port map( A1 => n16227, A2 => n16226, B1 => n16228, B2 => 
                           n16304, ZN => n17215);
   U579 : CLKBUF_X3 port map( A => n21700, Z => n25202);
   U582 : NOR2_X1 port map( A1 => n17494, A2 => n20665, ZN => n21700);
   U609 : BUF_X2 port map( A => n11063, Z => n25203);
   U611 : AND2_X2 port map( A1 => n25467, A2 => n25468, ZN => n18611);
   U624 : OAI211_X2 port map( C1 => n7915, C2 => n8076, A => n7160, B => n7159,
                           ZN => n9082);
   U628 : OAI211_X2 port map( C1 => n22316, C2 => n22612, A => n22315, B => 
                           n22314, ZN => n23164);
   U635 : AND2_X2 port map( A1 => n2448, A2 => n6540, ZN => n7384);
   U637 : NOR2_X2 port map( A1 => n12949, A2 => n12950, ZN => n14208);
   U639 : NAND2_X2 port map( A1 => n10629, A2 => n25306, ZN => n11735);
   U650 : AND3_X2 port map( A1 => n1435, A2 => n1378, A3 => n4609, ZN => n1370)
                           ;
   U655 : NAND4_X2 port map( A1 => n7253, A2 => n7254, A3 => n7251, A4 => n7252
                           , ZN => n8542);
   U661 : OAI22_X2 port map( A1 => n4807, A2 => n3736, B1 => n4806, B2 => n3735
                           , ZN => n17275);
   U667 : AND2_X2 port map( A1 => n683, A2 => n682, ZN => n4807);
   U669 : AOI22_X1 port map( A1 => n9385, A2 => n10185, B1 => n8262, B2 => 
                           n8261, ZN => n10505);
   U697 : OR2_X2 port map( A1 => n5491, A2 => n3834, ZN => n21981);
   U715 : AND2_X2 port map( A1 => n1665, A2 => n25318, ZN => n21573);
   U722 : OAI211_X1 port map( C1 => n23200, C2 => n23199, A => n24609, B => 
                           n24612, ZN => n23211);
   U728 : AND2_X2 port map( A1 => n473, A2 => n474, ZN => n18275);
   U731 : NAND2_X2 port map( A1 => n13961, A2 => n13960, ZN => n15109);
   U732 : XNOR2_X2 port map( A => Key(8), B => Plaintext(8), ZN => n6034);
   U734 : AND2_X2 port map( A1 => n3757, A2 => n24295, ZN => n11401);
   U736 : NOR2_X2 port map( A1 => n953, A2 => n954, ZN => n10886);
   U739 : NOR2_X2 port map( A1 => n13616, A2 => n13615, ZN => n14755);
   U740 : CLKBUF_X1 port map( A => n20233, Z => n25204);
   U752 : BUF_X2 port map( A => n20233, Z => n25205);
   U753 : OAI211_X1 port map( C1 => n19483, C2 => n19482, A => n24605, B => 
                           n24716, ZN => n20233);
   U754 : BUF_X1 port map( A => n10147, Z => n25207);
   U761 : XNOR2_X1 port map( A => n25137, B => n25136, ZN => n10147);
   U764 : AND2_X2 port map( A1 => n4673, A2 => n4674, ZN => n4672);
   U771 : AND2_X2 port map( A1 => n1318, A2 => n1317, ZN => n10870);
   U795 : NAND2_X2 port map( A1 => n22920, A2 => n23018, ZN => n23531);
   U803 : MUX2_X2 port map( A => n22913, B => n22912, S => n23461, Z => n22920)
                           ;
   U809 : NAND2_X2 port map( A1 => n10981, A2 => n10980, ZN => n12410);
   U812 : AND3_X4 port map( A1 => n5259, A2 => n5258, A3 => n5260, ZN => n23112
                           );
   U819 : XNOR2_X2 port map( A => n11963, B => n11964, ZN => n12834);
   U821 : OR2_X2 port map( A1 => n16701, A2 => n16700, ZN => n20335);
   U822 : AND2_X2 port map( A1 => n1532, A2 => n5273, ZN => n10793);
   U827 : CLKBUF_X1 port map( A => n14242, Z => n25208);
   U835 : BUF_X1 port map( A => n14242, Z => n25209);
   U836 : AOI22_X2 port map( A1 => n15578, A2 => n15577, B1 => n15576, B2 => 
                           n15575, ZN => n18240);
   U842 : BUF_X2 port map( A => n6062, Z => n6733);
   U844 : OR2_X2 port map( A1 => n18654, A2 => n18655, ZN => n20616);
   U845 : XNOR2_X2 port map( A => n16664, B => n16665, ZN => n19555);
   U847 : XNOR2_X2 port map( A => n5851, B => Key(154), ZN => n6767);
   U857 : OAI211_X2 port map( C1 => n7344, C2 => n7256, A => n7260, B => n7259,
                           ZN => n8345);
   U858 : XNOR2_X2 port map( A => Key(176), B => Plaintext(176), ZN => n5966);
   U859 : XNOR2_X2 port map( A => n5874, B => Key(58), ZN => n6976);
   U860 : NAND2_X2 port map( A1 => n3173, A2 => n6646, ZN => n7364);
   U866 : BUF_X2 port map( A => n12795, Z => n25085);
   U871 : OAI211_X2 port map( C1 => n2413, C2 => n9848, A => n9847, B => n9846,
                           ZN => n10698);
   U873 : AOI21_X2 port map( B1 => n17269, B2 => n17270, A => n17268, ZN => 
                           n18285);
   U878 : NAND3_X2 port map( A1 => n13608, A2 => n1061, A3 => n1060, ZN => 
                           n15487);
   U885 : XNOR2_X2 port map( A => Key(159), B => Plaintext(159), ZN => n6915);
   U894 : AND2_X1 port map( A1 => n13108, A2 => n12856, ZN => n13661);
   U895 : XNOR2_X2 port map( A => n12229, B => n12228, ZN => n13108);
   U897 : AND3_X2 port map( A1 => n5353, A2 => n5352, A3 => n5354, ZN => n11116
                           );
   U904 : BUF_X1 port map( A => n19105, Z => n24344);
   U914 : XNOR2_X2 port map( A => n3670, B => n3669, ZN => n16268);
   U915 : NAND2_X2 port map( A1 => n16860, A2 => n24229, ZN => n18308);
   U917 : MUX2_X2 port map( A => n10578, B => n10577, S => n11175, Z => n11638)
                           ;
   U918 : AND3_X2 port map( A1 => n3244, A2 => n5108, A3 => n3243, ZN => n11637
                           );
   U919 : OAI211_X2 port map( C1 => n15669, C2 => n16334, A => n2286, B => 
                           n1444, ZN => n16927);
   U925 : XNOR2_X2 port map( A => n15511, B => n15510, ZN => n16437);
   U927 : OAI211_X2 port map( C1 => n5630, C2 => n5628, A => n5629, B => n5627,
                           ZN => n11619);
   U928 : OAI211_X2 port map( C1 => n6754, C2 => n5808, A => n5807, B => n5806,
                           ZN => n7579);
   U931 : XNOR2_X2 port map( A => n21095, B => n21094, ZN => n23998);
   U937 : XNOR2_X2 port map( A => n11497, B => n11496, ZN => n13067);
   U938 : OR2_X2 port map( A1 => n962, A2 => n958, ZN => n3428);
   U939 : NAND3_X2 port map( A1 => n3054, A2 => n17133, A3 => n3053, ZN => 
                           n18341);
   U946 : NAND2_X2 port map( A1 => n10998, A2 => n10999, ZN => n11907);
   U951 : NAND2_X2 port map( A1 => n3918, A2 => n109, ZN => n20597);
   U960 : XNOR2_X2 port map( A => n15030, B => n15031, ZN => n16342);
   U961 : XNOR2_X2 port map( A => n5782, B => Key(94), ZN => n6233);
   U969 : XNOR2_X2 port map( A => n6004, B => Key(101), ZN => n625);
   U970 : NAND2_X2 port map( A1 => n15652, A2 => n726, ZN => n17316);
   U971 : XNOR2_X2 port map( A => n5159, B => n5160, ZN => n19446);
   U975 : NAND3_X2 port map( A1 => n25134, A2 => n25135, A3 => n10366, ZN => 
                           n11960);
   U1008 : BUF_X1 port map( A => n16176, Z => n25210);
   U1012 : MUX2_X2 port map( A => n9381, B => n10255, S => n10128, Z => n10729)
                           ;
   U1014 : BUF_X1 port map( A => n20182, Z => n25211);
   U1020 : BUF_X1 port map( A => n20182, Z => n25212);
   U1021 : OAI21_X1 port map( B1 => n358, B2 => n18723, A => n18722, ZN => 
                           n20182);
   U1026 : XNOR2_X2 port map( A => n12418, B => n12417, ZN => n13345);
   U1030 : OR2_X2 port map( A1 => n15722, A2 => n15721, ZN => n16708);
   U1033 : CLKBUF_X1 port map( A => n17361, Z => n25213);
   U1051 : BUF_X1 port map( A => n17361, Z => n25214);
   U1057 : BUF_X1 port map( A => n17361, Z => n25215);
   U1058 : OAI211_X1 port map( C1 => n3544, C2 => n16402, A => n15913, B => 
                           n24792, ZN => n17361);
   U1067 : NAND2_X2 port map( A1 => n12693, A2 => n5021, ZN => n14141);
   U1068 : NOR2_X2 port map( A1 => n17500, A2 => n17499, ZN => n18994);
   U1070 : AOI21_X2 port map( B1 => n13866, B2 => n13865, A => n2225, ZN => 
                           n14724);
   U1073 : XNOR2_X2 port map( A => n5790, B => Key(86), ZN => n5796);
   U1078 : XNOR2_X2 port map( A => n11720, B => n11721, ZN => n12555);
   U1080 : AOI22_X1 port map( A1 => n9579, A2 => n9578, B1 => n9577, B2 => 
                           n10904, ZN => n12150);
   U1081 : XNOR2_X2 port map( A => n11430, B => n12013, ZN => n13057);
   U1084 : OAI21_X2 port map( B1 => n18882, B2 => n24344, A => n1547, ZN => 
                           n20522);
   U1101 : OAI21_X2 port map( B1 => n1282, B2 => n1281, A => n1280, ZN => n8613
                           );
   U1113 : XNOR2_X2 port map( A => n21637, B => n21636, ZN => n22938);
   U1138 : BUF_X2 port map( A => n16388, Z => n15977);
   U1139 : XNOR2_X2 port map( A => n5839, B => Key(138), ZN => n6078);
   U1143 : CLKBUF_X1 port map( A => n9931, Z => n25216);
   U1148 : XNOR2_X1 port map( A => n7614, B => n7613, ZN => n9931);
   U1150 : CLKBUF_X1 port map( A => n17167, Z => n25218);
   U1158 : BUF_X2 port map( A => n17167, Z => n25219);
   U1160 : AOI22_X1 port map( A1 => n16059, A2 => n16473, B1 => n16058, B2 => 
                           n16474, ZN => n17167);
   U1162 : XNOR2_X2 port map( A => n7310, B => n7311, ZN => n9211);
   U1172 : NAND2_X2 port map( A1 => n2841, A2 => n6399, ZN => n7563);
   U1178 : CLKBUF_X1 port map( A => n20095, Z => n25220);
   U1179 : CLKBUF_X3 port map( A => n20095, Z => n25221);
   U1180 : NOR2_X1 port map( A1 => n19730, A2 => n18395, ZN => n20095);
   U1183 : XNOR2_X2 port map( A => n11625, B => n11624, ZN => n12534);
   U1184 : XNOR2_X2 port map( A => Key(157), B => Plaintext(157), ZN => n6918);
   U1186 : XNOR2_X2 port map( A => n5990, B => Key(105), ZN => n6823);
   U1192 : XNOR2_X2 port map( A => n2113, B => n14316, ZN => n16381);
   U1193 : BUF_X2 port map( A => n21493, Z => n25222);
   U1195 : OAI22_X1 port map( A1 => n18859, A2 => n19850, B1 => n20071, B2 => 
                           n18858, ZN => n21493);
   U1206 : XNOR2_X2 port map( A => n10745, B => n10744, ZN => n13150);
   U1207 : XNOR2_X2 port map( A => n20123, B => n20122, ZN => n22361);
   U1219 : XNOR2_X2 port map( A => n12374, B => n12373, ZN => n12636);
   U1220 : NAND3_X2 port map( A1 => n24215, A2 => n11103, A3 => n11104, ZN => 
                           n12212);
   U1238 : NAND2_X2 port map( A1 => n3088, A2 => n4561, ZN => n10772);
   U1245 : XNOR2_X2 port map( A => n11383, B => n11382, ZN => n13027);
   U1246 : NOR2_X2 port map( A1 => n2385, A2 => n10454, ZN => n12209);
   U1254 : AOI21_X2 port map( B1 => n9870, B2 => n9869, A => n9868, ZN => 
                           n10970);
   U1255 : OR2_X2 port map( A1 => n14024, A2 => n14023, ZN => n15097);
   U1260 : AND4_X2 port map( A1 => n10697, A2 => n10695, A3 => n10696, A4 => 
                           n3209, ZN => n11661);
   U1269 : XNOR2_X2 port map( A => n8097, B => n8096, ZN => n9027);
   U1278 : OAI21_X2 port map( B1 => n17245, B2 => n17246, A => n17244, ZN => 
                           n18621);
   U1283 : AND2_X2 port map( A1 => n14441, A2 => n1446, ZN => n15223);
   U1287 : XNOR2_X2 port map( A => Key(107), B => Plaintext(107), ZN => n5992);
   U1292 : INV_X1 port map( A => n13578, ZN => n14182);
   U1300 : NOR2_X2 port map( A1 => n13542, A2 => n13541, ZN => n15178);
   U1301 : XNOR2_X2 port map( A => n21405, B => n21404, ZN => n22932);
   U1307 : BUF_X1 port map( A => n20217, Z => n25223);
   U1308 : CLKBUF_X1 port map( A => n20217, Z => n25224);
   U1313 : XNOR2_X2 port map( A => Key(109), B => Plaintext(109), ZN => n6244);
   U1320 : BUF_X1 port map( A => n17108, Z => n25225);
   U1321 : BUF_X1 port map( A => n17108, Z => n25226);
   U1324 : CLKBUF_X1 port map( A => n17108, Z => n25227);
   U1326 : AOI21_X1 port map( B1 => n4338, B2 => n15805, A => n4337, ZN => 
                           n17108);
   U1331 : OAI211_X2 port map( C1 => n14198, C2 => n14148, A => n14147, B => 
                           n3678, ZN => n15526);
   U1339 : OAI211_X2 port map( C1 => n13484, C2 => n12678, A => n12677, B => 
                           n12676, ZN => n14845);
   U1358 : OAI21_X2 port map( B1 => n5934, B2 => n5935, A => n5933, ZN => n7464
                           );
   U1372 : BUF_X2 port map( A => n9045, Z => n25228);
   U1373 : BUF_X1 port map( A => n10736, Z => n25229);
   U1380 : BUF_X2 port map( A => n10736, Z => n25230);
   U1382 : XNOR2_X2 port map( A => n16738, B => n24719, ZN => n19264);
   U1396 : CLKBUF_X1 port map( A => n10953, Z => n25231);
   U1416 : BUF_X1 port map( A => n10953, Z => n25232);
   U1427 : CLKBUF_X1 port map( A => n10953, Z => n25233);
   U1438 : XNOR2_X2 port map( A => n11859, B => n11860, ZN => n12928);
   U1444 : XNOR2_X2 port map( A => n5961, B => Key(163), ZN => n6480);
   U1460 : XNOR2_X2 port map( A => n11871, B => n11872, ZN => n12897);
   U1470 : OAI21_X2 port map( B1 => n12832, B2 => n5644, A => n5643, ZN => 
                           n4844);
   U1479 : OAI21_X2 port map( B1 => n6994, B2 => n6995, A => n6993, ZN => n7961
                           );
   U1484 : XNOR2_X2 port map( A => n7206, B => n7207, ZN => n9388);
   U1498 : OAI21_X2 port map( B1 => n20363, B2 => n20362, A => n20361, ZN => 
                           n21996);
   U1508 : XNOR2_X2 port map( A => n25140, B => n18503, ZN => n19460);
   U1515 : OAI21_X2 port map( B1 => n4898, B2 => n4896, A => n16511, ZN => 
                           n16616);
   U1527 : AND2_X2 port map( A1 => n4900, A2 => n617, ZN => n16511);
   U1541 : XNOR2_X2 port map( A => n14872, B => n14871, ZN => n16220);
   U1544 : XNOR2_X2 port map( A => n111, B => n11980, ZN => n13265);
   U1546 : NOR2_X2 port map( A1 => n16874, A2 => n16875, ZN => n17969);
   U1553 : XNOR2_X2 port map( A => n11405, B => n11404, ZN => n13028);
   U1564 : XNOR2_X2 port map( A => n15382, B => n15381, ZN => n16067);
   U1612 : OAI211_X2 port map( C1 => n12749, C2 => n14058, A => n12748, B => 
                           n12747, ZN => n15184);
   U1621 : NOR2_X2 port map( A1 => n22943, A2 => n22942, ZN => n24492);
   U1638 : OAI21_X2 port map( B1 => n15671, B2 => n5706, A => n13375, ZN => 
                           n17414);
   U1657 : BUF_X2 port map( A => n12369, Z => n25234);
   U1688 : XNOR2_X2 port map( A => n12078, B => n12079, ZN => n231);
   U1697 : XNOR2_X2 port map( A => n6002, B => Key(118), ZN => n6848);
   U1698 : XNOR2_X2 port map( A => n5303, B => n5301, ZN => n19313);
   U1717 : OAI21_X2 port map( B1 => n9392, B2 => n1093, A => n1092, ZN => 
                           n10583);
   U1718 : BUF_X2 port map( A => n8945, Z => n25235);
   U1722 : OAI21_X2 port map( B1 => n3729, B2 => n3730, A => n551, ZN => n10369
                           );
   U1739 : XNOR2_X2 port map( A => n1576, B => Key(59), ZN => n1147);
   U1775 : BUF_X2 port map( A => n12137, Z => n25236);
   U1783 : AND3_X2 port map( A1 => n1216, A2 => n1215, A3 => n1220, ZN => 
                           n11440);
   U1804 : AOI21_X2 port map( B1 => n7245, B2 => n7186, A => n1736, ZN => n9107
                           );
   U1808 : XNOR2_X2 port map( A => n8885, B => n8884, ZN => n9433);
   U1809 : NAND2_X2 port map( A1 => n20189, A2 => n1487, ZN => n22007);
   U1813 : CLKBUF_X1 port map( A => n15697, Z => n25237);
   U1818 : BUF_X2 port map( A => n15697, Z => n25238);
   U1822 : CLKBUF_X1 port map( A => n23251, Z => n24377);
   U1848 : NAND2_X1 port map( A1 => n21758, A2 => n2690, ZN => n23595);
   U1855 : BUF_X1 port map( A => n23470, Z => n23481);
   U1874 : OAI211_X1 port map( C1 => n21913, C2 => n22273, A => n21912, B => 
                           n21911, ZN => n22575);
   U1881 : NOR2_X1 port map( A1 => n22204, A2 => n22203, ZN => n23740);
   U1882 : INV_X1 port map( A => n20561, ZN => n20562);
   U1889 : AOI22_X1 port map( A1 => n16834, A2 => n3981, B1 => n3982, B2 => 
                           n16833, ZN => n18124);
   U1910 : BUF_X1 port map( A => n17107, Z => n25245);
   U1919 : INV_X1 port map( A => n12535, ZN => n13051);
   U1959 : BUF_X1 port map( A => n9432, Z => n10890);
   U1983 : OR2_X1 port map( A1 => n434, A2 => n25251, ZN => n7675);
   U1990 : INV_X1 port map( A => n8219, ZN => n7812);
   U1991 : BUF_X1 port map( A => n8074, Z => n25253);
   U1999 : NAND3_X1 port map( A1 => n1764, A2 => n6816, A3 => n5830, ZN => 
                           n7581);
   U2007 : INV_X1 port map( A => n6699, ZN => n2008);
   U2018 : BUF_X2 port map( A => Key(45), Z => n22986);
   U2024 : AND2_X1 port map( A1 => n25550, A2 => n23277, ZN => n23259);
   U2052 : INV_X1 port map( A => n23905, ZN => n25239);
   U2054 : OAI211_X1 port map( C1 => n22179, C2 => n24369, A => n22177, B => 
                           n22178, ZN => n24998);
   U2076 : AND3_X1 port map( A1 => n22120, A2 => n22119, A3 => n22118, ZN => 
                           n23537);
   U2082 : INV_X1 port map( A => n23858, ZN => n25240);
   U2084 : OR2_X1 port map( A1 => n23201, A2 => n22575, ZN => n5769);
   U2090 : AND3_X1 port map( A1 => n22486, A2 => n4648, A3 => n22485, ZN => 
                           n22528);
   U2102 : AND2_X1 port map( A1 => n25299, A2 => n25298, ZN => n21786);
   U2111 : OR2_X1 port map( A1 => n22752, A2 => n211, ZN => n22569);
   U2120 : OR2_X1 port map( A1 => n24924, A2 => n24923, ZN => n24910);
   U2137 : AND2_X1 port map( A1 => n22689, A2 => n22685, ZN => n25275);
   U2143 : INV_X1 port map( A => n22235, ZN => n25553);
   U2152 : AND2_X1 port map( A1 => n22242, A2 => n22243, ZN => n22063);
   U2188 : AND2_X1 port map( A1 => n22208, A2 => n22064, ZN => n22066);
   U2193 : XNOR2_X1 port map( A => n25334, B => n20739, ZN => n24496);
   U2196 : INV_X1 port map( A => n20740, ZN => n25334);
   U2198 : XNOR2_X1 port map( A => n21674, B => n21673, ZN => n22900);
   U2199 : AND3_X1 port map( A1 => n25556, A2 => n20013, A3 => n25555, ZN => 
                           n21160);
   U2200 : NOR2_X1 port map( A1 => n20295, A2 => n20294, ZN => n25470);
   U2247 : NAND2_X1 port map( A1 => n5466, A2 => n19123, ZN => n21541);
   U2265 : OAI21_X1 port map( B1 => n20004, B2 => n2864, A => n1420, ZN => 
                           n25400);
   U2274 : NAND3_X1 port map( A1 => n25316, A2 => n20347, A3 => n25315, ZN => 
                           n21334);
   U2303 : OR2_X1 port map( A1 => n20328, A2 => n19878, ZN => n20091);
   U2308 : AND2_X1 port map( A1 => n19714, A2 => n20317, ZN => n19888);
   U2313 : NOR2_X1 port map( A1 => n55, A2 => n21008, ZN => n19668);
   U2323 : INV_X1 port map( A => n21068, ZN => n25579);
   U2325 : OR2_X1 port map( A1 => n20174, A2 => n20588, ZN => n19952);
   U2330 : AND2_X1 port map( A1 => n18212, A2 => n19723, ZN => n20561);
   U2332 : AND2_X1 port map( A1 => n3810, A2 => n3809, ZN => n24940);
   U2344 : OR2_X1 port map( A1 => n18845, A2 => n18844, ZN => n19851);
   U2367 : AOI21_X1 port map( B1 => n19760, B2 => n25540, A => n25539, ZN => 
                           n2662);
   U2368 : INV_X1 port map( A => n19376, ZN => n25243);
   U2411 : AND2_X1 port map( A1 => n19097, A2 => n4114, ZN => n19363);
   U2421 : INV_X1 port map( A => n19598, ZN => n25244);
   U2429 : NAND3_X1 port map( A1 => n5103, A2 => n644, A3 => n208, ZN => n18423
                           );
   U2459 : AND2_X1 port map( A1 => n5295, A2 => n16559, ZN => n18102);
   U2503 : NAND2_X1 port map( A1 => n17232, A2 => n1339, ZN => n18665);
   U2523 : OAI211_X1 port map( C1 => n3602, C2 => n16214, A => n16213, B => 
                           n16212, ZN => n18549);
   U2525 : AND2_X1 port map( A1 => n25524, A2 => n16556, ZN => n2790);
   U2549 : INV_X1 port map( A => n17464, ZN => n25572);
   U2576 : AND3_X1 port map( A1 => n15586, A2 => n25280, A3 => n25279, ZN => 
                           n17069);
   U2597 : OR2_X1 port map( A1 => n4624, A2 => n15691, ZN => n25575);
   U2645 : NOR2_X1 port map( A1 => n15693, A2 => n25259, ZN => n25576);
   U2657 : AOI22_X1 port map( A1 => n14352, A2 => n16381, B1 => n15659, B2 => 
                           n14351, ZN => n25433);
   U2675 : INV_X1 port map( A => n16303, ZN => n25272);
   U2679 : INV_X1 port map( A => n16955, ZN => n25246);
   U2683 : AND2_X1 port map( A1 => n16102, A2 => n25586, ZN => n25585);
   U2694 : CLKBUF_X1 port map( A => n15986, Z => n25492);
   U2704 : OR2_X1 port map( A1 => n4600, A2 => n14101, ZN => n2002);
   U2708 : AND2_X1 port map( A1 => n25570, A2 => n4497, ZN => n13969);
   U2747 : NAND3_X1 port map( A1 => n2436, A2 => n2438, A3 => n25592, ZN => 
                           n14150);
   U2774 : INV_X1 port map( A => n14054, ZN => n25247);
   U2785 : OAI21_X1 port map( B1 => n13661, B2 => n13663, A => n13662, ZN => 
                           n13485);
   U2787 : OR2_X1 port map( A1 => n12733, A2 => n12728, ZN => n137);
   U2801 : OR2_X1 port map( A1 => n12206, A2 => n24617, ZN => n13662);
   U2820 : XNOR2_X1 port map( A => n11656, B => n25541, ZN => n24601);
   U2830 : INV_X1 port map( A => n12914, ZN => n25248);
   U2867 : AND2_X1 port map( A1 => n24856, A2 => n5516, ZN => n25396);
   U2879 : BUF_X2 port map( A => n12368, Z => n25371);
   U2895 : AND2_X1 port map( A1 => n9333, A2 => n9332, ZN => n11112);
   U2908 : INV_X1 port map( A => n11128, ZN => n25249);
   U2909 : INV_X1 port map( A => n11117, ZN => n10868);
   U2943 : AND3_X1 port map( A1 => n711, A2 => n471, A3 => n25341, ZN => n11046
                           );
   U2956 : OAI21_X1 port map( B1 => n10043, B2 => n10042, A => n10041, ZN => 
                           n11069);
   U2976 : BUF_X2 port map( A => n10336, Z => n25250);
   U2980 : AND3_X1 port map( A1 => n24104, A2 => n5741, A3 => n5334, ZN => 
                           n11117);
   U2982 : OR2_X1 port map( A1 => n9281, A2 => n8141, ZN => n9203);
   U2987 : XNOR2_X1 port map( A => n8822, B => n8823, ZN => n9729);
   U3001 : AND2_X1 port map( A1 => n25538, A2 => n7219, ZN => n8336);
   U3012 : NAND2_X1 port map( A1 => n25319, A2 => n2217, ZN => n7813);
   U3013 : BUF_X2 port map( A => n263, Z => n25251);
   U3039 : OR2_X1 port map( A1 => n6366, A2 => n6365, ZN => n25527);
   U3041 : AOI21_X1 port map( B1 => n6879, B2 => n2976, A => n2045, ZN => n7449
                           );
   U3051 : INV_X1 port map( A => n7581, ZN => n7879);
   U3069 : INV_X1 port map( A => n7771, ZN => n25252);
   U3072 : INV_X1 port map( A => n6686, ZN => n6977);
   U3113 : BUF_X2 port map( A => n6919, Z => n24037);
   U3116 : XNOR2_X1 port map( A => n5873, B => Key(56), ZN => n6686);
   U3118 : OR2_X1 port map( A1 => n6301, A2 => n6489, ZN => n6305);
   U3126 : XNOR2_X1 port map( A => Key(35), B => Plaintext(35), ZN => n25437);
   U3137 : AND2_X1 port map( A1 => n6010, A2 => n7609, ZN => n25277);
   U3141 : OR2_X1 port map( A1 => n6398, A2 => n6730, ZN => n2841);
   U3158 : BUF_X1 port map( A => n6122, Z => n6990);
   U3211 : BUF_X1 port map( A => n7327, Z => n248);
   U3228 : OR2_X1 port map( A1 => n6551, A2 => n6860, ZN => n25305);
   U3266 : OR2_X1 port map( A1 => n7862, A2 => n7864, ZN => n25535);
   U3270 : OAI211_X1 port map( C1 => n6070, C2 => n1975, A => n1974, B => n1973
                           , ZN => n8604);
   U3315 : OR2_X1 port map( A1 => n9603, A2 => n9599, ZN => n9930);
   U3329 : BUF_X1 port map( A => n10018, Z => n24495);
   U3345 : BUF_X1 port map( A => n9997, Z => n246);
   U3350 : CLKBUF_X1 port map( A => n9898, Z => n24054);
   U3379 : INV_X1 port map( A => n714, ZN => n10306);
   U3387 : AND3_X1 port map( A1 => n9326, A2 => n10082, A3 => n10079, ZN => 
                           n10871);
   U3389 : OR2_X1 port map( A1 => n9986, A2 => n9985, ZN => n25341);
   U3392 : NAND3_X1 port map( A1 => n9552, A2 => n1399, A3 => n9551, ZN => 
                           n10746);
   U3399 : INV_X1 port map( A => n10371, ZN => n25507);
   U3400 : OAI211_X1 port map( C1 => n7839, C2 => n9346, A => n848, B => n847, 
                           ZN => n11005);
   U3411 : OR2_X1 port map( A1 => n11112, A2 => n11117, ZN => n10725);
   U3459 : INV_X1 port map( A => n10728, ZN => n10481);
   U3466 : AND2_X1 port map( A1 => n10574, A2 => n11038, ZN => n991);
   U3469 : NOR2_X1 port map( A1 => n408, A2 => n13057, ZN => n25551);
   U3482 : XNOR2_X1 port map( A => n12104, B => n25257, ZN => n4568);
   U3486 : XNOR2_X1 port map( A => n11637, B => n11638, ZN => n12132);
   U3518 : XNOR2_X1 port map( A => n11713, B => n11712, ZN => n12914);
   U3564 : OR2_X1 port map( A1 => n13056, A2 => n12795, ZN => n25336);
   U3579 : INV_X1 port map( A => n11655, ZN => n25541);
   U3590 : OAI211_X1 port map( C1 => n13365, C2 => n12980, A => n13366, B => 
                           n25301, ZN => n1316);
   U3593 : BUF_X1 port map( A => n13039, Z => n12799);
   U3605 : XNOR2_X1 port map( A => n11904, B => n11903, ZN => n12945);
   U3613 : AND2_X1 port map( A1 => n14194, A2 => n25360, ZN => n13478);
   U3620 : OR2_X1 port map( A1 => n1579, A2 => n3755, ZN => n25537);
   U3661 : OR2_X1 port map( A1 => n14082, A2 => n14083, ZN => n25504);
   U3663 : AND2_X1 port map( A1 => n14419, A2 => n628, ZN => n15451);
   U3689 : NAND2_X1 port map( A1 => n13715, A2 => n25321, ZN => n14671);
   U3705 : OR2_X1 port map( A1 => n16101, A2 => n16100, ZN => n15579);
   U3745 : CLKBUF_X1 port map( A => n16008, Z => n25410);
   U3749 : XNOR2_X1 port map( A => n25518, B => n15168, ZN => n14699);
   U3790 : AND2_X1 port map( A1 => n1365, A2 => n15802, ZN => n25294);
   U3807 : INV_X1 port map( A => n16462, ZN => n25596);
   U3808 : CLKBUF_X1 port map( A => n15470, Z => n15546);
   U3817 : BUF_X1 port map( A => n16451, Z => n257);
   U3821 : CLKBUF_X1 port map( A => n16470, Z => n24550);
   U3825 : OR2_X1 port map( A1 => n16422, A2 => n15958, ZN => n25591);
   U3846 : INV_X1 port map( A => n940, ZN => n16404);
   U3850 : AND2_X1 port map( A1 => n213, A2 => n25510, ZN => n25509);
   U3851 : OR2_X1 port map( A1 => n17207, A2 => n17015, ZN => n5510);
   U3865 : OR2_X1 port map( A1 => n15546, A2 => n383, ZN => n16056);
   U3886 : CLKBUF_X1 port map( A => n15656, Z => n15659);
   U3889 : OAI21_X1 port map( B1 => n16193, B2 => n25447, A => n25323, ZN => 
                           n5414);
   U3917 : AND2_X1 port map( A1 => n25213, A2 => n16989, ZN => n16769);
   U3930 : OAI21_X1 port map( B1 => n16280, B2 => n4092, A => n5336, ZN => 
                           n16561);
   U3935 : CLKBUF_X1 port map( A => n17352, Z => n25491);
   U3993 : OAI211_X1 port map( C1 => n4972, C2 => n16472, A => n16056, B => 
                           n25356, ZN => n17297);
   U4017 : OR2_X1 port map( A1 => n376, A2 => n16917, ZN => n15576);
   U4060 : OR2_X1 port map( A1 => n16634, A2 => n24570, ZN => n638);
   U4065 : AND2_X1 port map( A1 => n19472, A2 => n19470, ZN => n18958);
   U4112 : AND3_X1 port map( A1 => n5136, A2 => n1437, A3 => n3993, ZN => 
                           n18435);
   U4120 : INV_X1 port map( A => n4647, ZN => n19106);
   U4128 : INV_X1 port map( A => n1361, ZN => n25540);
   U4142 : BUF_X1 port map( A => n17496, Z => n19327);
   U4199 : OR2_X1 port map( A1 => n3470, A2 => n4436, ZN => n5237);
   U4204 : NOR2_X1 port map( A1 => n20317, A2 => n20319, ZN => n25309);
   U4234 : NAND2_X1 port map( A1 => n19258, A2 => n5027, ZN => n20427);
   U4243 : OR2_X1 port map( A1 => n20507, A2 => n20216, ZN => n25348);
   U4248 : OAI21_X1 port map( B1 => n17896, B2 => n17895, A => n17894, ZN => 
                           n20102);
   U4251 : AOI21_X1 port map( B1 => n19116, B2 => n19115, A => n19114, ZN => 
                           n20516);
   U4268 : OAI211_X1 port map( C1 => n18773, C2 => n353, A => n4458, B => n4459
                           , ZN => n20346);
   U4275 : BUF_X1 port map( A => n20367, Z => n24558);
   U4285 : AND2_X1 port map( A1 => n25266, A2 => n19668, ZN => n19673);
   U4289 : INV_X1 port map( A => n20309, ZN => n20130);
   U4290 : OR2_X1 port map( A1 => n20469, A2 => n20062, ZN => n25302);
   U4291 : NAND2_X1 port map( A1 => n4185, A2 => n20267, ZN => n21172);
   U4328 : XNOR2_X1 port map( A => n21583, B => n21670, ZN => n21121);
   U4340 : XNOR2_X1 port map( A => n20903, B => n2569, ZN => n5503);
   U4359 : INV_X1 port map( A => n21815, ZN => n25297);
   U4396 : XNOR2_X1 port map( A => n21244, B => n21243, ZN => n22792);
   U4400 : OR2_X1 port map( A1 => n333, A2 => n22564, ZN => n22406);
   U4417 : AND2_X1 port map( A1 => n22131, A2 => n22968, ZN => n25308);
   U4454 : BUF_X1 port map( A => n22139, Z => n22337);
   U4523 : NOR2_X1 port map( A1 => n22185, A2 => n22184, ZN => n23671);
   U4713 : AND2_X1 port map( A1 => n23492, A2 => n23494, ZN => n25517);
   U4744 : OR2_X1 port map( A1 => n23204, A2 => n23203, ZN => n23208);
   U4745 : AOI21_X1 port map( B1 => n22841, B2 => n22840, A => n22839, ZN => 
                           n24426);
   U4746 : AOI21_X1 port map( B1 => n23455, B2 => n23456, A => n25517, ZN => 
                           n25516);
   U4752 : CLKBUF_X1 port map( A => Key(176), Z => n1854);
   U4760 : CLKBUF_X1 port map( A => Key(20), Z => n16574);
   U4886 : CLKBUF_X1 port map( A => Key(68), Z => n1864);
   U4888 : CLKBUF_X1 port map( A => Key(131), Z => n2782);
   U4950 : AND2_X1 port map( A1 => n16023, A2 => n15773, ZN => n25254);
   U4983 : OR2_X1 port map( A1 => n19465, A2 => n19464, ZN => n25255);
   U4988 : AND2_X1 port map( A1 => n17242, A2 => n17241, ZN => n25256);
   U4992 : INV_X1 port map( A => n6034, ZN => n25325);
   U4998 : INV_X1 port map( A => n20217, ZN => n25345);
   U4999 : XOR2_X1 port map( A => n12102, B => n16, Z => n25257);
   U5023 : XNOR2_X1 port map( A => n11436, B => n11437, ZN => n13053);
   U5034 : INV_X1 port map( A => n13053, ZN => n25337);
   U5073 : INV_X1 port map( A => n13221, ZN => n25292);
   U5090 : INV_X1 port map( A => n13788, ZN => n25560);
   U5097 : XOR2_X1 port map( A => n15253, B => n20690, Z => n25258);
   U5104 : AND2_X1 port map( A1 => n16051, A2 => n4897, ZN => n25259);
   U5131 : INV_X1 port map( A => n25389, ZN => n25284);
   U5163 : XNOR2_X1 port map( A => n10882, B => n10883, ZN => n13102);
   U5168 : INV_X1 port map( A => n17119, ZN => n25357);
   U5211 : XOR2_X1 port map( A => n18617, B => n18618, Z => n25260);
   U5290 : OR2_X1 port map( A1 => n25260, A2 => n19441, ZN => n25261);
   U5310 : AND3_X1 port map( A1 => n17675, A2 => n5456, A3 => n5455, ZN => 
                           n25262);
   U5336 : AND2_X1 port map( A1 => n20316, A2 => n19889, ZN => n25263);
   U5355 : AND2_X1 port map( A1 => n24982, A2 => n19578, ZN => n25264);
   U5375 : NAND2_X1 port map( A1 => n19181, A2 => n4792, ZN => n20215);
   U5387 : INV_X1 port map( A => n20215, ZN => n25347);
   U5400 : AND3_X1 port map( A1 => n25303, A2 => n19642, A3 => n25302, ZN => 
                           n25265);
   U5401 : OR2_X1 port map( A1 => n20522, A2 => n20523, ZN => n25266);
   U5438 : NAND2_X1 port map( A1 => n13713, A2 => n13394, ZN => n1486);
   U5513 : XNOR2_X1 port map( A => n25267, B => n23729, ZN => Ciphertext(137));
   U5588 : NAND3_X1 port map( A1 => n23726, A2 => n23725, A3 => n786, ZN => 
                           n25267);
   U5697 : NAND2_X1 port map( A1 => n13234, A2 => n13298, ZN => n2842);
   U5716 : XNOR2_X2 port map( A => n11831, B => n11830, ZN => n13298);
   U5721 : NAND2_X1 port map( A1 => n25163, A2 => n25164, ZN => n9309);
   U5728 : XNOR2_X1 port map( A => n25268, B => n768, ZN => Ciphertext(120));
   U5732 : NAND2_X1 port map( A1 => n22153, A2 => n22152, ZN => n25268);
   U5749 : OR2_X2 port map( A1 => n25269, A2 => n6821, ZN => n7985);
   U5759 : AOI21_X1 port map( B1 => n6816, B2 => n6817, A => n6894, ZN => 
                           n25269);
   U5762 : NAND2_X1 port map( A1 => n7585, A2 => n7581, ZN => n7314);
   U5767 : OAI21_X2 port map( B1 => n13654, B2 => n1899, A => n25270, ZN => 
                           n14644);
   U5772 : NAND3_X1 port map( A1 => n13657, A2 => n13658, A3 => n13922, ZN => 
                           n25270);
   U5774 : NAND2_X1 port map( A1 => n25412, A2 => n16971, ZN => n16915);
   U5844 : NAND3_X1 port map( A1 => n535, A2 => n21294, A3 => n534, ZN => 
                           n22539);
   U5876 : NAND2_X1 port map( A1 => n6425, A2 => n5966, ZN => n6314);
   U5886 : OAI211_X2 port map( C1 => n4884, C2 => n4167, A => n18867, B => 
                           n25271, ZN => n21008);
   U5936 : NAND2_X1 port map( A1 => n18866, A2 => n19113, ZN => n25271);
   U5950 : NAND2_X1 port map( A1 => n4139, A2 => n19112, ZN => n18865);
   U6035 : NOR2_X2 port map( A1 => n17333, A2 => n16602, ZN => n16917);
   U6082 : NAND2_X1 port map( A1 => n24185, A2 => n965, ZN => n17333);
   U6168 : NAND2_X1 port map( A1 => n25272, A2 => n25254, ZN => n965);
   U6195 : NAND2_X1 port map( A1 => n25273, A2 => n16107, ZN => n969);
   U6207 : NAND2_X1 port map( A1 => n15854, A2 => n2478, ZN => n25273);
   U6216 : AND3_X2 port map( A1 => n3481, A2 => n3483, A3 => n3477, ZN => 
                           n21559);
   U6222 : NAND2_X1 port map( A1 => n3479, A2 => n3478, ZN => n3477);
   U6237 : NAND2_X1 port map( A1 => n5756, A2 => n16068, ZN => n15795);
   U6242 : NAND2_X1 port map( A1 => n365, A2 => n17633, ZN => n17475);
   U6261 : NAND2_X1 port map( A1 => n15606, A2 => n25274, ZN => n879);
   U6263 : NOR2_X1 port map( A1 => n294, A2 => n16051, ZN => n25274);
   U6274 : NAND2_X1 port map( A1 => n16838, A2 => n25219, ZN => n16839);
   U6295 : NAND4_X1 port map( A1 => n21821, A2 => n21818, A3 => n21820, A4 => 
                           n21819, ZN => n21828);
   U6308 : NAND2_X1 port map( A1 => n25395, A2 => n25275, ZN => n21819);
   U6309 : OAI21_X1 port map( B1 => n25264, B2 => n25276, A => n280, ZN => 
                           n1131);
   U6311 : NOR2_X1 port map( A1 => n19056, A2 => n19057, ZN => n25276);
   U6320 : NAND3_X1 port map( A1 => n4894, A2 => n13437, A3 => n25445, ZN => 
                           n2003);
   U6343 : INV_X1 port map( A => n1514, ZN => n22475);
   U6350 : NAND2_X1 port map( A1 => n22798, A2 => n22805, ZN => n1514);
   U6365 : NAND2_X1 port map( A1 => n20269, A2 => n20498, ZN => n61);
   U6413 : NAND2_X1 port map( A1 => n19074, A2 => n24700, ZN => n20269);
   U6425 : AOI22_X1 port map( A1 => n14099, A2 => n14211, B1 => n24376, B2 => 
                           n14101, ZN => n14217);
   U6444 : OAI211_X2 port map( C1 => n13120, C2 => n13119, A => n2097, B => 
                           n2980, ZN => n14101);
   U6455 : NAND3_X1 port map( A1 => n4927, A2 => n15061, A3 => n15679, ZN => 
                           n564);
   U6496 : OR2_X1 port map( A1 => n11109, A2 => n13144, ZN => n13141);
   U6503 : NAND2_X1 port map( A1 => n2555, A2 => n25277, ZN => n2554);
   U6507 : NAND3_X1 port map( A1 => n25278, A2 => n14101, A3 => n13552, ZN => 
                           n4891);
   U6513 : INV_X1 port map( A => n24375, ZN => n25278);
   U6514 : NAND2_X1 port map( A1 => n15585, A2 => n5100, ZN => n25279);
   U6546 : NAND2_X1 port map( A1 => n25587, A2 => n3410, ZN => n25280);
   U6554 : NAND2_X1 port map( A1 => n7760, A2 => n7761, ZN => n7392);
   U6594 : OR2_X2 port map( A1 => n6172, A2 => n5068, ZN => n7760);
   U6603 : NAND2_X1 port map( A1 => n3743, A2 => n15767, ZN => n16639);
   U6613 : NAND2_X1 port map( A1 => n10533, A2 => n11146, ZN => n714);
   U6667 : NAND2_X1 port map( A1 => n24116, A2 => n21010, ZN => n19972);
   U6668 : NAND2_X1 port map( A1 => n21008, A2 => n20290, ZN => n21010);
   U6708 : NAND2_X1 port map( A1 => n23070, A2 => n23071, ZN => n23073);
   U6786 : NAND2_X1 port map( A1 => n20089, A2 => n3480, ZN => n3479);
   U6809 : NAND3_X1 port map( A1 => n20459, A2 => n20461, A3 => n24461, ZN => 
                           n25139);
   U6819 : NAND2_X2 port map( A1 => n25281, A2 => n2885, ZN => n23748);
   U6882 : NAND3_X1 port map( A1 => n22248, A2 => n22247, A3 => n22246, ZN => 
                           n25281);
   U6883 : NAND2_X1 port map( A1 => n486, A2 => n25282, ZN => n17832);
   U6884 : NAND2_X1 port map( A1 => n25562, A2 => n4683, ZN => n25282);
   U6928 : NAND2_X1 port map( A1 => n23927, A2 => n24948, ZN => n23928);
   U6951 : NAND2_X1 port map( A1 => n2604, A2 => n2093, ZN => n14786);
   U6960 : NAND2_X1 port map( A1 => n15765, A2 => n25283, ZN => n17081);
   U7022 : OAI211_X1 port map( C1 => n16246, C2 => n16247, A => n25285, B => 
                           n25284, ZN => n25283);
   U7109 : NAND2_X1 port map( A1 => n16246, A2 => n25484, ZN => n25285);
   U7114 : XNOR2_X2 port map( A => n18672, B => n25286, ZN => n19173);
   U7115 : XNOR2_X1 port map( A => n18668, B => n18667, ZN => n25286);
   U7137 : NAND3_X1 port map( A1 => n23205, A2 => n23206, A3 => n2903, ZN => 
                           n23210);
   U7151 : NAND2_X1 port map( A1 => n10119, A2 => n10118, ZN => n11212);
   U7152 : AND3_X2 port map( A1 => n1035, A2 => n1036, A3 => n25287, ZN => 
                           n5120);
   U7171 : NAND3_X1 port map( A1 => n1032, A2 => n17475, A3 => n1033, ZN => 
                           n25287);
   U7177 : NAND2_X2 port map( A1 => n20431, A2 => n5043, ZN => n21525);
   U7195 : AOI21_X1 port map( B1 => n25289, B2 => n25288, A => n20428, ZN => 
                           n20430);
   U7261 : INV_X1 port map( A => n3047, ZN => n25288);
   U7265 : NAND2_X1 port map( A1 => n19253, A2 => n24943, ZN => n25289);
   U7320 : AND2_X1 port map( A1 => n18959, A2 => n19466, ZN => n18840);
   U7325 : OAI22_X1 port map( A1 => n3646, A2 => n3645, B1 => n17049, B2 => 
                           n17052, ZN => n17532);
   U7353 : NAND2_X1 port map( A1 => n25378, A2 => n20017, ZN => n25362);
   U7386 : NOR2_X1 port map( A1 => n20137, A2 => n19991, ZN => n20017);
   U7399 : AND2_X2 port map( A1 => n21917, A2 => n22324, ZN => n22752);
   U7409 : OAI21_X1 port map( B1 => n18986, B2 => n3296, A => n3297, ZN => 
                           n25290);
   U7416 : XNOR2_X1 port map( A => n17839, B => n17874, ZN => n24192);
   U7418 : NOR2_X2 port map( A1 => n16825, A2 => n807, ZN => n17839);
   U7446 : NAND2_X1 port map( A1 => n25291, A2 => n3098, ZN => n10653);
   U7447 : NAND2_X1 port map( A1 => n10804, A2 => n3100, ZN => n25291);
   U7448 : NAND2_X1 port map( A1 => n4340, A2 => n1544, ZN => n1539);
   U7459 : NAND3_X1 port map( A1 => n20433, A2 => n24940, A3 => n20434, ZN => 
                           n20435);
   U7472 : NAND2_X1 port map( A1 => n5208, A2 => n20576, ZN => n20433);
   U7492 : OR3_X1 port map( A1 => n23696, A2 => n22148, A3 => n22082, ZN => 
                           n3441);
   U7501 : NAND3_X1 port map( A1 => n25293, A2 => n13222, A3 => n25292, ZN => 
                           n4486);
   U7504 : INV_X1 port map( A => n12919, ZN => n25293);
   U7518 : NAND2_X1 port map( A1 => n656, A2 => n658, ZN => n6441);
   U7526 : NAND2_X1 port map( A1 => n7702, A2 => n7701, ZN => n8203);
   U7558 : NAND2_X1 port map( A1 => n4353, A2 => n25294, ZN => n15313);
   U7578 : XNOR2_X2 port map( A => n25295, B => n14994, ZN => n16225);
   U7579 : XNOR2_X1 port map( A => n14995, B => n15000, ZN => n25295);
   U7599 : NAND2_X1 port map( A1 => n17338, A2 => n17337, ZN => n645);
   U7602 : NAND2_X1 port map( A1 => n19395, A2 => n19163, ZN => n19016);
   U7662 : NAND3_X1 port map( A1 => n18, A2 => n2258, A3 => n19, ZN => n17321);
   U7668 : OAI21_X1 port map( B1 => n23311, B2 => n23327, A => n5660, ZN => 
                           n2143);
   U7682 : OAI21_X2 port map( B1 => n21788, B2 => n22063, A => n25296, ZN => 
                           n23769);
   U7689 : NAND2_X1 port map( A1 => n21786, A2 => n25297, ZN => n25296);
   U7691 : NAND2_X1 port map( A1 => n22180, A2 => n22239, ZN => n25298);
   U7695 : INV_X1 port map( A => n22241, ZN => n25299);
   U7698 : NAND2_X1 port map( A1 => n12973, A2 => n25300, ZN => n14124);
   U7715 : OR2_X1 port map( A1 => n12971, A2 => n5412, ZN => n25300);
   U7745 : NAND2_X1 port map( A1 => n17207, A2 => n17216, ZN => n17210);
   U7804 : NAND2_X1 port map( A1 => n12583, A2 => n12980, ZN => n25301);
   U7817 : OAI21_X1 port map( B1 => n19640, B2 => n20471, A => n20470, ZN => 
                           n25303);
   U7819 : XNOR2_X1 port map( A => n25304, B => n23448, ZN => Ciphertext(94));
   U7820 : NAND4_X1 port map( A1 => n23447, A2 => n23446, A3 => n23445, A4 => 
                           n23444, ZN => n25304);
   U7884 : NAND2_X1 port map( A1 => n16639, A2 => n15557, ZN => n3744);
   U7916 : NAND3_X1 port map( A1 => n1214, A2 => n15912, A3 => n3544, ZN => 
                           n24792);
   U7968 : NAND2_X1 port map( A1 => n6550, A2 => n25305, ZN => n8484);
   U7977 : NAND2_X1 port map( A1 => n10628, A2 => n44, ZN => n25306);
   U8057 : NAND2_X1 port map( A1 => n7474, A2 => n7421, ZN => n7953);
   U8069 : AOI21_X1 port map( B1 => n9557, B2 => n9556, A => n9555, ZN => 
                           n25307);
   U8092 : NAND2_X1 port map( A1 => n5529, A2 => n5530, ZN => n22144);
   U8114 : NOR2_X2 port map( A1 => n25308, A2 => n22130, ZN => n24349);
   U8171 : OAI21_X1 port map( B1 => n25263, B2 => n25309, A => n24917, ZN => 
                           n19892);
   U8183 : NAND2_X1 port map( A1 => n25311, A2 => n25310, ZN => n15976);
   U8207 : NAND2_X1 port map( A1 => n15973, A2 => n15970, ZN => n25310);
   U8226 : NAND2_X1 port map( A1 => n746, A2 => n25312, ZN => n25311);
   U8238 : INV_X1 port map( A => n15973, ZN => n25312);
   U8242 : NAND2_X1 port map( A1 => n22187, A2 => n25313, ZN => n22192);
   U8244 : OR2_X1 port map( A1 => n25070, A2 => n22922, ZN => n25313);
   U8252 : NAND2_X1 port map( A1 => n22712, A2 => n22928, ZN => n22187);
   U8255 : OAI211_X2 port map( C1 => n20248, C2 => n24077, A => n25314, B => 
                           n20247, ZN => n21087);
   U8265 : NAND2_X1 port map( A1 => n24818, A2 => n24077, ZN => n25314);
   U8269 : NAND2_X1 port map( A1 => n9236, A2 => n9757, ZN => n2268);
   U8273 : NAND2_X1 port map( A1 => n2269, A2 => n1814, ZN => n9236);
   U8305 : NAND2_X1 port map( A1 => n22959, A2 => n22958, ZN => n22034);
   U8322 : NOR2_X1 port map( A1 => n7562, A2 => n7725, ZN => n1596);
   U8348 : NAND2_X1 port map( A1 => n7246, A2 => n7563, ZN => n7562);
   U8351 : NOR2_X2 port map( A1 => n23667, A2 => n5508, ZN => n23670);
   U8366 : NAND2_X1 port map( A1 => n22161, A2 => n24768, ZN => n23667);
   U8380 : NAND2_X1 port map( A1 => n19463, A2 => n25255, ZN => n19494);
   U8391 : NAND2_X1 port map( A1 => n24414, A2 => n20343, ZN => n25315);
   U8411 : NAND2_X1 port map( A1 => n3671, A2 => n20344, ZN => n25316);
   U8419 : OAI21_X2 port map( B1 => n15703, B2 => n4552, A => n25317, ZN => 
                           n18539);
   U8447 : NAND3_X1 port map( A1 => n2338, A2 => n15701, A3 => n15700, ZN => 
                           n25317);
   U8460 : AOI22_X1 port map( A1 => n19740, A2 => n1667, B1 => n20430, B2 => 
                           n5044, ZN => n25318);
   U8462 : NAND2_X1 port map( A1 => n25324, A2 => n25327, ZN => n25319);
   U8509 : NAND3_X1 port map( A1 => n16127, A2 => n129, A3 => n24528, ZN => 
                           n17173);
   U8510 : OAI21_X1 port map( B1 => n7382, B2 => n7622, A => n7616, ZN => n6223
                           );
   U8512 : NAND2_X1 port map( A1 => n7618, A2 => n7382, ZN => n7616);
   U8515 : NAND3_X1 port map( A1 => n17287, A2 => n17284, A3 => n16951, ZN => 
                           n24635);
   U8516 : INV_X1 port map( A => n24249, ZN => n25508);
   U8519 : NAND2_X1 port map( A1 => n25320, A2 => n849, ZN => n16256);
   U8528 : NAND3_X1 port map( A1 => n15938, A2 => n25389, A3 => n24162, ZN => 
                           n25320);
   U8529 : OAI21_X1 port map( B1 => n3031, B2 => n3030, A => n13394, ZN => 
                           n25321);
   U8540 : NAND2_X1 port map( A1 => n7111, A2 => n7112, ZN => n8891);
   U8543 : NAND2_X1 port map( A1 => n22348, A2 => n25395, ZN => n21821);
   U8570 : NAND2_X1 port map( A1 => n16257, A2 => n17216, ZN => n25524);
   U8607 : NOR2_X2 port map( A1 => n25322, A2 => n13872, ZN => n15120);
   U8609 : AOI21_X1 port map( B1 => n3403, B2 => n3400, A => n5440, ZN => 
                           n25322);
   U8627 : NAND2_X1 port map( A1 => n23288, A2 => n23289, ZN => n23291);
   U8678 : NAND2_X1 port map( A1 => n1030, A2 => n25261, ZN => n19082);
   U8732 : NAND2_X1 port map( A1 => n305, A2 => n10850, ZN => n10272);
   U8749 : NAND3_X1 port map( A1 => n24669, A2 => n3826, A3 => n3829, ZN => 
                           n24633);
   U8780 : NAND3_X1 port map( A1 => n7945, A2 => n7946, A3 => n7657, ZN => 
                           n7950);
   U8795 : INV_X1 port map( A => n16191, ZN => n25323);
   U8799 : NAND2_X1 port map( A1 => n25326, A2 => n25325, ZN => n25324);
   U8801 : NAND2_X1 port map( A1 => n6499, A2 => n6434, ZN => n25326);
   U8821 : NAND2_X1 port map( A1 => n6353, A2 => n6034, ZN => n25327);
   U8831 : NAND2_X1 port map( A1 => n25328, A2 => n3410, ZN => n2076);
   U8846 : NAND2_X1 port map( A1 => n15579, A2 => n15582, ZN => n25328);
   U8851 : NAND2_X1 port map( A1 => n556, A2 => n9587, ZN => n10612);
   U8856 : OAI21_X2 port map( B1 => n138, B2 => n16242, A => n25329, ZN => 
                           n16578);
   U8878 : NAND2_X1 port map( A1 => n24294, A2 => n24292, ZN => n25329);
   U8885 : OAI22_X1 port map( A1 => n5020, A2 => n25330, B1 => n14192, B2 => 
                           n14191, ZN => n14197);
   U8886 : NAND2_X1 port map( A1 => n24186, A2 => n14191, ZN => n25330);
   U8887 : NAND2_X1 port map( A1 => n1694, A2 => n4446, ZN => n17);
   U8892 : NAND2_X1 port map( A1 => n25331, A2 => n4823, ZN => n12962);
   U8922 : NAND2_X1 port map( A1 => n4822, A2 => n399, ZN => n25331);
   U8950 : XNOR2_X1 port map( A => n15252, B => n25258, ZN => n15256);
   U8996 : NAND3_X1 port map( A1 => n1275, A2 => n1272, A3 => n1273, ZN => 
                           n25147);
   U8998 : XNOR2_X1 port map( A => n25332, B => n22301, ZN => Ciphertext(45));
   U9003 : NAND3_X1 port map( A1 => n188, A2 => n2083, A3 => n22299, ZN => 
                           n25332);
   U9025 : OAI22_X1 port map( A1 => n14270, A2 => n14271, B1 => n14273, B2 => 
                           n24368, ZN => n14277);
   U9027 : NAND2_X1 port map( A1 => n14344, A2 => n3059, ZN => n24701);
   U9036 : XNOR2_X1 port map( A => n25333, B => n17868, ZN => n17871);
   U9038 : XNOR2_X1 port map( A => n17866, B => n18601, ZN => n25333);
   U9102 : NAND2_X1 port map( A1 => n5404, A2 => n19678, ZN => n21336);
   U9135 : NAND3_X2 port map( A1 => n3801, A2 => n3802, A3 => n13967, ZN => 
                           n15153);
   U9187 : NAND3_X1 port map( A1 => n715, A2 => n973, A3 => n25335, ZN => 
                           n14324);
   U9236 : NAND3_X1 port map( A1 => n25337, A2 => n13057, A3 => n25336, ZN => 
                           n25335);
   U9238 : NAND2_X1 port map( A1 => n22941, A2 => n22940, ZN => n21654);
   U9256 : NAND2_X1 port map( A1 => n17559, A2 => n19264, ZN => n3470);
   U9259 : XNOR2_X2 port map( A => n3852, B => n3853, ZN => n19413);
   U9262 : INV_X1 port map( A => n22483, ZN => n25569);
   U9263 : NAND3_X1 port map( A1 => n10481, A2 => n10482, A3 => n10262, ZN => 
                           n10267);
   U9296 : NAND2_X1 port map( A1 => n13744, A2 => n14168, ZN => n14171);
   U9323 : NAND2_X2 port map( A1 => n1783, A2 => n12446, ZN => n13744);
   U9343 : NAND2_X1 port map( A1 => n25338, A2 => n17374, ZN => n17874);
   U9344 : NAND2_X1 port map( A1 => n3693, A2 => n5522, ZN => n25338);
   U9345 : NAND2_X1 port map( A1 => n17574, A2 => n373, ZN => n17370);
   U9380 : OAI21_X1 port map( B1 => n7615, B2 => n7382, A => n25339, ZN => 
                           n7383);
   U9382 : NAND2_X1 port map( A1 => n7382, A2 => n7380, ZN => n25339);
   U9398 : NAND3_X1 port map( A1 => n1217, A2 => n410, A3 => n1219, ZN => n1215
                           );
   U9406 : NAND3_X1 port map( A1 => n25340, A2 => n1478, A3 => n22188, ZN => 
                           n2456);
   U9410 : NAND2_X1 port map( A1 => n22107, A2 => n25070, ZN => n25340);
   U9411 : NAND2_X1 port map( A1 => n25342, A2 => n24267, ZN => n16724);
   U9526 : NAND2_X1 port map( A1 => n16720, A2 => n17059, ZN => n25342);
   U9556 : AND2_X2 port map( A1 => n25343, A2 => n24272, ZN => n19939);
   U9559 : NAND2_X1 port map( A1 => n19308, A2 => n19307, ZN => n25343);
   U9596 : NAND2_X1 port map( A1 => n4328, A2 => n25344, ZN => n20804);
   U9643 : NAND3_X1 port map( A1 => n25348, A2 => n25346, A3 => n25345, ZN => 
                           n25344);
   U9645 : NAND2_X1 port map( A1 => n25347, A2 => n20507, ZN => n25346);
   U9689 : NAND2_X1 port map( A1 => n24910, A2 => n23967, ZN => n22693);
   U9712 : NAND3_X1 port map( A1 => n2600, A2 => n6686, A3 => n24579, ZN => 
                           n5876);
   U9812 : NAND3_X1 port map( A1 => n6721, A2 => n1609, A3 => n6720, ZN => 
                           n6726);
   U9813 : NAND2_X1 port map( A1 => n16367, A2 => n16206, ZN => n16365);
   U9849 : NAND2_X1 port map( A1 => n19469, A2 => n19470, ZN => n458);
   U9854 : NAND2_X1 port map( A1 => n19466, A2 => n19321, ZN => n19469);
   U9859 : NAND2_X1 port map( A1 => n11085, A2 => n10438, ZN => n10221);
   U9873 : OR3_X1 port map( A1 => n9459, A2 => n9918, A3 => n9463, ZN => n9135)
                           ;
   U9874 : NAND3_X1 port map( A1 => n1968, A2 => n13994, A3 => n13993, ZN => 
                           n1966);
   U9889 : NAND3_X1 port map( A1 => n16998, A2 => n24471, A3 => n374, ZN => 
                           n15994);
   U9951 : NAND3_X1 port map( A1 => n19374, A2 => n19373, A3 => n25349, ZN => 
                           n19774);
   U9979 : NAND2_X1 port map( A1 => n19363, A2 => n25243, ZN => n25349);
   U10008 : NAND4_X2 port map( A1 => n2425, A2 => n19776, A3 => n2427, A4 => 
                           n2426, ZN => n21267);
   U10023 : NOR2_X2 port map( A1 => n20044, A2 => n20045, ZN => n4294);
   U10027 : BUF_X1 port map( A => n12439, Z => n13064);
   U10057 : AND2_X1 port map( A1 => n22715, A2 => n22927, ZN => n25557);
   U10069 : NAND3_X1 port map( A1 => n10694, A2 => n11057, A3 => n11053, ZN => 
                           n3209);
   U10146 : NAND2_X2 port map( A1 => n25350, A2 => n12432, ZN => n14165);
   U10147 : NAND3_X1 port map( A1 => n2192, A2 => n12429, A3 => n12430, ZN => 
                           n25350);
   U10161 : NAND3_X1 port map( A1 => n1895, A2 => n7384, A3 => n7380, ZN => 
                           n7201);
   U10196 : NAND2_X1 port map( A1 => n4181, A2 => n25351, ZN => n1268);
   U10220 : NAND2_X1 port map( A1 => n13114, A2 => n12660, ZN => n25351);
   U10239 : NAND2_X1 port map( A1 => n17172, A2 => n17522, ZN => n17176);
   U10247 : NAND2_X1 port map( A1 => n17170, A2 => n17171, ZN => n17172);
   U10267 : NAND3_X1 port map( A1 => n3283, A2 => n23716, A3 => n23723, ZN => 
                           n3280);
   U10280 : NAND2_X1 port map( A1 => n3888, A2 => n2684, ZN => n2683);
   U10348 : NAND3_X1 port map( A1 => n17353, A2 => n4840, A3 => n4004, ZN => 
                           n16673);
   U10361 : NAND2_X1 port map( A1 => n25354, A2 => n25352, ZN => n12599);
   U10395 : NAND2_X1 port map( A1 => n25353, A2 => n13292, ZN => n25352);
   U10397 : MUX2_X1 port map( A => n12911, B => n13288, S => n12593, Z => 
                           n25353);
   U10420 : NAND2_X1 port map( A1 => n25355, A2 => n12596, ZN => n25354);
   U10455 : INV_X1 port map( A => n13292, ZN => n25355);
   U10458 : NAND3_X2 port map( A1 => n24628, A2 => n10624, A3 => n10625, ZN => 
                           n12370);
   U10478 : OAI211_X1 port map( C1 => n16472, C2 => n16473, A => n16469, B => 
                           n24550, ZN => n25356);
   U10483 : AND3_X2 port map( A1 => n21279, A2 => n5765, A3 => n4079, ZN => 
                           n23066);
   U10563 : NAND3_X1 port map( A1 => n25358, A2 => n2580, A3 => n25357, ZN => 
                           n17105);
   U10581 : INV_X1 port map( A => n17100, ZN => n25358);
   U10596 : NAND3_X2 port map( A1 => n687, A2 => n16536, A3 => n686, ZN => 
                           n18451);
   U10664 : XNOR2_X1 port map( A => n25359, B => n451, ZN => Ciphertext(83));
   U10673 : NAND3_X1 port map( A1 => n25142, A2 => n25141, A3 => n22884, ZN => 
                           n25359);
   U10692 : XNOR2_X2 port map( A => n18236, B => n18235, ZN => n19186);
   U10697 : NAND2_X1 port map( A1 => n10162, A2 => n10161, ZN => n8417);
   U10712 : INV_X1 port map( A => n14189, ZN => n25360);
   U10721 : NAND2_X1 port map( A1 => n13785, A2 => n14143, ZN => n14194);
   U10723 : OAI21_X1 port map( B1 => n997, B2 => n24063, A => n25361, ZN => 
                           n22309);
   U10768 : NAND2_X1 port map( A1 => n22308, A2 => n24063, ZN => n25361);
   U10789 : OAI211_X2 port map( C1 => n19758, C2 => n19759, A => n19756, B => 
                           n25362, ZN => n21245);
   U10793 : NAND2_X1 port map( A1 => n18768, A2 => n25363, ZN => n18769);
   U10794 : NAND2_X1 port map( A1 => n25364, A2 => n18767, ZN => n25363);
   U10806 : INV_X1 port map( A => n19307, ZN => n25364);
   U10808 : NAND3_X1 port map( A1 => n12477, A2 => n13041, A3 => n12797, ZN => 
                           n12480);
   U10809 : NAND2_X1 port map( A1 => n13039, A2 => n13038, ZN => n12797);
   U10838 : NAND2_X1 port map( A1 => n24118, A2 => n4520, ZN => n25548);
   U10840 : NAND2_X1 port map( A1 => n19183, A2 => n18597, ZN => n19426);
   U10895 : NAND2_X1 port map( A1 => n4795, A2 => n4793, ZN => n654);
   U10911 : NAND3_X1 port map( A1 => n24344, A2 => n18166, A3 => n4647, ZN => 
                           n18167);
   U10949 : NAND2_X1 port map( A1 => n19199, A2 => n18809, ZN => n4647);
   U10966 : OAI21_X2 port map( B1 => n17950, B2 => n17949, A => n17948, ZN => 
                           n21532);
   U10997 : OAI21_X2 port map( B1 => n17393, B2 => n3602, A => n17392, ZN => 
                           n18531);
   U11074 : BUF_X1 port map( A => n23904, Z => n23896);
   U11106 : BUF_X1 port map( A => n22593, Z => n24042);
   U11127 : OAI21_X1 port map( B1 => n19699, B2 => n24378, A => n19698, ZN => 
                           n21300);
   U11137 : INV_X1 port map( A => n11159, ZN => n4737);
   U11159 : CLKBUF_X1 port map( A => n22975, Z => n25365);
   U11167 : XNOR2_X1 port map( A => n4101, B => n4100, ZN => n22975);
   U11169 : MUX2_X2 port map( A => n19848, B => n19847, S => n276, Z => n21660)
                           ;
   U11218 : INV_X1 port map( A => n12636, ZN => n25366);
   U11281 : OAI21_X1 port map( B1 => n5121, B2 => n20821, A => n20820, ZN => 
                           n25367);
   U11333 : OAI21_X1 port map( B1 => n5121, B2 => n20821, A => n20820, ZN => 
                           n23228);
   U11372 : OR2_X1 port map( A1 => n348, A2 => n20479, ZN => n1008);
   U11375 : OR2_X1 port map( A1 => n21885, A2 => n25368, ZN => n25175);
   U11407 : NAND2_X1 port map( A1 => n22401, A2 => n22400, ZN => n25368);
   U11433 : XNOR2_X2 port map( A => n19769, B => n19768, ZN => n21816);
   U11510 : NAND2_X1 port map( A1 => n13028, A2 => n13023, ZN => n25369);
   U11527 : XOR2_X1 port map( A => n11401, B => n12381, Z => n12385);
   U11528 : MUX2_X1 port map( A => n25214, B => n25058, S => n17039, Z => 
                           n25370);
   U11565 : AND2_X1 port map( A1 => n12934, A2 => n13267, ZN => n2632);
   U11569 : AOI21_X1 port map( B1 => n5711, B2 => n20473, A => n24704, ZN => 
                           n21173);
   U11571 : AOI22_X1 port map( A1 => n10316, A2 => n10661, B1 => n10315, B2 => 
                           n10556, ZN => n12368);
   U11575 : BUF_X1 port map( A => n20778, Z => n25372);
   U11581 : AOI21_X1 port map( B1 => n19908, B2 => n19912, A => n1755, ZN => 
                           n20778);
   U11599 : INV_X1 port map( A => n2869, ZN => n25373);
   U11600 : OR2_X1 port map( A1 => n24908, A2 => n24451, ZN => n19629);
   U11604 : BUF_X1 port map( A => n18902, Z => n19275);
   U11631 : OR2_X1 port map( A1 => n20491, A2 => n24078, ZN => n20076);
   U11641 : XOR2_X1 port map( A => n18268, B => n17110, Z => n17112);
   U11692 : MUX2_X1 port map( A => n14944, B => n14945, S => n2684, Z => n14948
                           );
   U11693 : CLKBUF_X1 port map( A => n14943, Z => n25458);
   U11784 : AND2_X1 port map( A1 => n5290, A2 => n18765, ZN => n25374);
   U11792 : XNOR2_X1 port map( A => n20880, B => n20879, ZN => n25375);
   U11793 : XNOR2_X1 port map( A => n20880, B => n20879, ZN => n22888);
   U11811 : OAI21_X1 port map( B1 => n3686, B2 => n13062, A => n24165, ZN => 
                           n14360);
   U11814 : BUF_X1 port map( A => n2375, Z => n25376);
   U11815 : OAI211_X1 port map( C1 => n20456, C2 => n24357, A => n24189, B => 
                           n24188, ZN => n25377);
   U11842 : XNOR2_X1 port map( A => n15279, B => n15278, ZN => n2375);
   U11846 : OAI211_X1 port map( C1 => n20456, C2 => n24357, A => n24189, B => 
                           n24188, ZN => n21402);
   U11888 : INV_X1 port map( A => n25242, ZN => n25378);
   U11957 : OAI211_X1 port map( C1 => n18974, C2 => n18975, A => n18973, B => 
                           n18972, ZN => n1629);
   U11975 : XNOR2_X1 port map( A => n20994, B => n20993, ZN => n22927);
   U11977 : XNOR2_X1 port map( A => n20863, B => n20862, ZN => n22093);
   U12050 : OAI211_X1 port map( C1 => n17169, C2 => n2430, A => n17168, B => 
                           n514, ZN => n25379);
   U12060 : BUF_X1 port map( A => n23697, Z => n23715);
   U12069 : XNOR2_X1 port map( A => n20773, B => n20772, ZN => n25381);
   U12096 : XNOR2_X1 port map( A => n20773, B => n20772, ZN => n22398);
   U12105 : AND2_X1 port map( A1 => n23251, A2 => n23242, ZN => n23235);
   U12127 : OR2_X1 port map( A1 => n7045, A2 => n5264, ZN => n24260);
   U12265 : OR2_X1 port map( A1 => n17300, A2 => n16708, ZN => n3775);
   U12281 : XOR2_X1 port map( A => n21698, B => n21697, Z => n25382);
   U12312 : XNOR2_X2 port map( A => n20818, B => n25222, ZN => n21697);
   U12369 : INV_X1 port map( A => n22655, ZN => n22606);
   U12482 : AND3_X2 port map( A1 => n3087, A2 => n4102, A3 => n4099, ZN => 
                           n1340);
   U12542 : CLKBUF_X1 port map( A => n20373, Z => n25383);
   U12656 : INV_X1 port map( A => n20373, ZN => n20369);
   U12675 : INV_X1 port map( A => n16360, ZN => n25546);
   U12725 : INV_X1 port map( A => n16105, ZN => n25587);
   U12756 : BUF_X1 port map( A => n22059, Z => n22241);
   U12769 : NAND3_X1 port map( A1 => n1747, A2 => n1748, A3 => n14224, ZN => 
                           n25384);
   U12822 : XOR2_X1 port map( A => n18109, B => n18218, Z => n16760);
   U12864 : NAND3_X1 port map( A1 => n1747, A2 => n1748, A3 => n14224, ZN => 
                           n15522);
   U12914 : NAND2_X1 port map( A1 => n3076, A2 => n3075, ZN => n25385);
   U13127 : NAND2_X1 port map( A1 => n3076, A2 => n3075, ZN => n21567);
   U13146 : NAND3_X1 port map( A1 => n2724, A2 => n20177, A3 => n2725, ZN => 
                           n25386);
   U13158 : NAND3_X1 port map( A1 => n2724, A2 => n20177, A3 => n2725, ZN => 
                           n25387);
   U13193 : NAND3_X1 port map( A1 => n2724, A2 => n20177, A3 => n2725, ZN => 
                           n21439);
   U13234 : NAND3_X2 port map( A1 => n17675, A2 => n5456, A3 => n5455, ZN => 
                           n25388);
   U13268 : OAI211_X1 port map( C1 => n20423, C2 => n20422, A => n20421, B => 
                           n20420, ZN => n21310);
   U13346 : OAI211_X1 port map( C1 => n22847, C2 => n22901, A => n25568, B => 
                           n22904, ZN => n4648);
   U13347 : OR2_X1 port map( A1 => n23147, A2 => n23146, ZN => n4627);
   U13547 : NAND2_X1 port map( A1 => n21190, A2 => n2781, ZN => n23077);
   U13597 : CLKBUF_X1 port map( A => n9237, Z => n10031);
   U13651 : XNOR2_X1 port map( A => n14766, B => n14767, ZN => n25389);
   U13983 : AND3_X1 port map( A1 => n638, A2 => n16632, A3 => n16631, ZN => 
                           n17873);
   U13993 : NOR2_X1 port map( A1 => n21291, A2 => n24625, ZN => n25391);
   U14016 : NOR2_X1 port map( A1 => n21291, A2 => n24625, ZN => n23030);
   U14021 : XNOR2_X1 port map( A => n18008, B => n18007, ZN => n25392);
   U14147 : XNOR2_X1 port map( A => n18008, B => n18007, ZN => n19360);
   U14386 : XNOR2_X1 port map( A => n8656, B => n8655, ZN => n25393);
   U14537 : XOR2_X1 port map( A => n11561, B => n11646, Z => n12246);
   U14560 : XNOR2_X1 port map( A => n8656, B => n8655, ZN => n10108);
   U14577 : OR2_X1 port map( A1 => n19257, A2 => n18831, ZN => n18055);
   U14588 : OAI211_X1 port map( C1 => n12846, C2 => n4241, A => n2769, B => 
                           n2770, ZN => n14336);
   U14691 : OR2_X1 port map( A1 => n21140, A2 => n22667, ZN => n22668);
   U14710 : AOI21_X1 port map( B1 => n14103, B2 => n4877, A => n4876, ZN => 
                           n3462);
   U14764 : OR2_X1 port map( A1 => n20216, A2 => n20510, ZN => n20200);
   U14808 : XOR2_X1 port map( A => n19832, B => n19833, Z => n25395);
   U14842 : AND2_X1 port map( A1 => n24856, A2 => n5516, ZN => n12003);
   U14921 : BUF_X1 port map( A => n20428, Z => n25397);
   U15030 : AOI22_X1 port map( A1 => n19236, A2 => n19237, B1 => n24310, B2 => 
                           n19234, ZN => n20428);
   U15121 : XNOR2_X1 port map( A => Key(14), B => Plaintext(14), ZN => n25398);
   U15162 : XNOR2_X1 port map( A => Key(14), B => Plaintext(14), ZN => n6521);
   U15215 : OAI211_X1 port map( C1 => n19010, C2 => n19171, A => n3821, B => 
                           n3820, ZN => n20145);
   U15269 : OAI21_X1 port map( B1 => n20608, B2 => n22369, A => n20607, ZN => 
                           n25399);
   U15301 : OAI21_X1 port map( B1 => n20608, B2 => n22369, A => n20607, ZN => 
                           n23859);
   U15308 : OR2_X1 port map( A1 => n22187, A2 => n25557, ZN => n24782);
   U15462 : OAI21_X1 port map( B1 => n20004, B2 => n2864, A => n1420, ZN => 
                           n21444);
   U15498 : XNOR2_X1 port map( A => n5951, B => Key(171), ZN => n25401);
   U15511 : OR2_X2 port map( A1 => n25402, A2 => n25403, ZN => n7537);
   U15586 : AND3_X1 port map( A1 => n6305, A2 => n6303, A3 => n6493, ZN => 
                           n25402);
   U15638 : NOR2_X1 port map( A1 => n1561, A2 => n4727, ZN => n25403);
   U15656 : XNOR2_X1 port map( A => n5951, B => Key(171), ZN => n6427);
   U15983 : OR2_X1 port map( A1 => n20248, A2 => n174, ZN => n679);
   U16070 : OAI21_X1 port map( B1 => n22393, B2 => n22858, A => n22035, ZN => 
                           n23394);
   U16071 : AOI22_X2 port map( A1 => n10204, A2 => n4507, B1 => n3443, B2 => 
                           n10203, ZN => n12314);
   U16126 : XOR2_X1 port map( A => n5968, B => Key(175), Z => n25404);
   U16186 : OR2_X1 port map( A1 => n23672, A2 => n23671, ZN => n25405);
   U16195 : AND2_X1 port map( A1 => n19875, A2 => n20022, ZN => n20093);
   U16251 : AOI21_X1 port map( B1 => n16013, B2 => n16012, A => n16011, ZN => 
                           n25406);
   U16469 : OAI21_X1 port map( B1 => n7199, B2 => n7198, A => n7197, ZN => 
                           n25407);
   U16586 : OAI21_X1 port map( B1 => n7199, B2 => n7198, A => n7197, ZN => 
                           n8633);
   U16621 : XNOR2_X1 port map( A => n11631, B => n11630, ZN => n25408);
   U16628 : XNOR2_X1 port map( A => n14728, B => n14727, ZN => n25409);
   U16641 : XNOR2_X1 port map( A => n11631, B => n11630, ZN => n13050);
   U16692 : BUF_X1 port map( A => n15657, Z => n16383);
   U16701 : NAND2_X1 port map( A1 => n892, A2 => n539, ZN => n25411);
   U16705 : NAND2_X1 port map( A1 => n892, A2 => n539, ZN => n18283);
   U16754 : BUF_X1 port map( A => n20475, Z => n21259);
   U16774 : NAND2_X1 port map( A1 => n17662, A2 => n17661, ZN => n18559);
   U16777 : OAI211_X1 port map( C1 => n24370, C2 => n20101, A => n20100, B => 
                           n20099, ZN => n2010);
   U16786 : BUF_X1 port map( A => n17334, Z => n25412);
   U16792 : OAI211_X1 port map( C1 => n22353, C2 => n22352, A => n22351, B => 
                           n22350, ZN => n23933);
   U16796 : OAI211_X1 port map( C1 => n13591, C2 => n13864, A => n2417, B => 
                           n5150, ZN => n25413);
   U16798 : XNOR2_X1 port map( A => n21111, B => n21110, ZN => n25414);
   U16812 : XNOR2_X1 port map( A => n21110, B => n21111, ZN => n23995);
   U16838 : XNOR2_X1 port map( A => n12394, B => n12395, ZN => n25415);
   U16896 : NOR3_X1 port map( A1 => n12883, A2 => n12882, A3 => n13600, ZN => 
                           n25416);
   U16918 : NOR3_X1 port map( A1 => n12883, A2 => n12882, A3 => n13600, ZN => 
                           n25417);
   U16927 : XNOR2_X1 port map( A => n12394, B => n12395, ZN => n13344);
   U16947 : NOR3_X1 port map( A1 => n12883, A2 => n12882, A3 => n13600, ZN => 
                           n14992);
   U16978 : XOR2_X1 port map( A => n12413, B => n12207, Z => n25418);
   U16992 : AND2_X1 port map( A1 => n13844, A2 => n13843, ZN => n1579);
   U17047 : XNOR2_X1 port map( A => n17788, B => n25419, ZN => n17794);
   U17059 : XOR2_X1 port map( A => n24488, B => n2318, Z => n25419);
   U17075 : NAND2_X1 port map( A1 => n4430, A2 => n4429, ZN => n25420);
   U17178 : NAND2_X1 port map( A1 => n4430, A2 => n4429, ZN => n25421);
   U17227 : NAND2_X1 port map( A1 => n4430, A2 => n4429, ZN => n20413);
   U17236 : XNOR2_X1 port map( A => n18617, B => n18618, ZN => n25422);
   U17257 : XNOR2_X1 port map( A => n18617, B => n18618, ZN => n25423);
   U17301 : XOR2_X1 port map( A => Key(98), B => Plaintext(98), Z => n25424);
   U17334 : INV_X1 port map( A => n301, ZN => n25425);
   U17564 : NAND2_X1 port map( A1 => n24734, A2 => n14305, ZN => n25426);
   U17617 : XNOR2_X1 port map( A => n5936, B => Key(3), ZN => n25427);
   U17659 : XNOR2_X1 port map( A => n5936, B => Key(3), ZN => n25428);
   U17691 : INV_X1 port map( A => n16895, ZN => n25429);
   U17730 : XNOR2_X1 port map( A => n5936, B => Key(3), ZN => n6513);
   U17807 : XNOR2_X1 port map( A => n12310, B => n12309, ZN => n25430);
   U17957 : OAI21_X1 port map( B1 => n13604, B2 => n14319, A => n13603, ZN => 
                           n25431);
   U18144 : XNOR2_X1 port map( A => n12310, B => n12309, ZN => n13352);
   U18261 : OAI21_X1 port map( B1 => n13604, B2 => n14319, A => n13603, ZN => 
                           n15521);
   U18333 : XOR2_X1 port map( A => n12783, B => n12782, Z => n25432);
   U18334 : AOI22_X1 port map( A1 => n14352, A2 => n16381, B1 => n15659, B2 => 
                           n14351, ZN => n16955);
   U18406 : BUF_X1 port map( A => n13998, Z => n25434);
   U18464 : BUF_X1 port map( A => n13998, Z => n25435);
   U18465 : AOI21_X1 port map( B1 => n13342, B2 => n13341, A => n3126, ZN => 
                           n13998);
   U18467 : OAI211_X1 port map( C1 => n13780, C2 => n13779, A => n4354, B => 
                           n13778, ZN => n25436);
   U18492 : OAI211_X1 port map( C1 => n13780, C2 => n13779, A => n4354, B => 
                           n13778, ZN => n14384);
   U18495 : XNOR2_X1 port map( A => n21984, B => n21983, ZN => n25438);
   U18648 : XNOR2_X1 port map( A => Key(35), B => Plaintext(35), ZN => n5904);
   U18676 : XNOR2_X1 port map( A => n21984, B => n21983, ZN => n22838);
   U18677 : XNOR2_X1 port map( A => n21104, B => n21105, ZN => n25439);
   U18678 : XNOR2_X1 port map( A => n21104, B => n21105, ZN => n23994);
   U18695 : OR2_X1 port map( A1 => n10104, A2 => n9773, ZN => n8643);
   U18706 : CLKBUF_X1 port map( A => n20386, Z => n25440);
   U18716 : XNOR2_X1 port map( A => n17668, B => n17667, ZN => n20386);
   U18763 : XNOR2_X1 port map( A => n15060, B => n15059, ZN => n25441);
   U18788 : XNOR2_X1 port map( A => n21573, B => n21721, ZN => n25442);
   U18789 : XNOR2_X1 port map( A => n15060, B => n15059, ZN => n15746);
   U18790 : XNOR2_X2 port map( A => n15182, B => n15181, ZN => n16311);
   U18818 : OAI21_X1 port map( B1 => n13885, B2 => n4293, A => n790, ZN => 
                           n25443);
   U18819 : OAI21_X1 port map( B1 => n13885, B2 => n4293, A => n790, ZN => 
                           n15316);
   U18910 : CLKBUF_X1 port map( A => n9423, Z => n25444);
   U18923 : OR2_X1 port map( A1 => n21008, A2 => n20290, ZN => n25558);
   U18955 : NOR2_X1 port map( A1 => n13099, A2 => n13100, ZN => n25445);
   U18966 : XNOR2_X1 port map( A => n15414, B => n15413, ZN => n25446);
   U18983 : NOR2_X1 port map( A1 => n13099, A2 => n13100, ZN => n24503);
   U19042 : AOI22_X2 port map( A1 => n20357, A2 => n20356, B1 => n20355, B2 => 
                           n2168, ZN => n21511);
   U19071 : XNOR2_X1 port map( A => n15256, B => n15257, ZN => n25447);
   U19072 : OAI21_X1 port map( B1 => n18873, B2 => n18874, A => n18872, ZN => 
                           n20291);
   U19108 : INV_X1 port map( A => n19554, ZN => n25448);
   U19109 : XNOR2_X1 port map( A => n16698, B => n16697, ZN => n19290);
   U19122 : XNOR2_X2 port map( A => n14855, B => n14856, ZN => n16465);
   U19191 : XNOR2_X1 port map( A => n14380, B => n14379, ZN => n25449);
   U19300 : XOR2_X1 port map( A => n20791, B => n20790, Z => n25450);
   U19329 : INV_X1 port map( A => n2624, ZN => n25451);
   U19330 : NOR2_X1 port map( A1 => n21148, A2 => n21149, ZN => n25452);
   U19383 : NOR2_X1 port map( A1 => n21148, A2 => n21149, ZN => n23065);
   U19541 : XNOR2_X1 port map( A => n8474, B => n8473, ZN => n25453);
   U19542 : AND3_X2 port map( A1 => n4005, A2 => n5599, A3 => n4003, ZN => 
                           n17817);
   U19546 : INV_X1 port map( A => n20428, ZN => n276);
   U19549 : XOR2_X1 port map( A => n2797, B => n8570, Z => n25454);
   U19578 : XNOR2_X1 port map( A => n2812, B => n13544, ZN => n25455);
   U19593 : XNOR2_X1 port map( A => n2812, B => n13544, ZN => n16331);
   U19601 : NOR2_X1 port map( A1 => n20319, A2 => n25456, ZN => n17568);
   U19629 : NAND2_X1 port map( A1 => n19889, A2 => n19714, ZN => n25456);
   U19635 : OR2_X1 port map( A1 => n6866, A2 => n2404, ZN => n2965);
   U19677 : XNOR2_X1 port map( A => n8723, B => n8724, ZN => n25457);
   U19714 : AOI22_X1 port map( A1 => n12644, A2 => n12643, B1 => n12641, B2 => 
                           n12642, ZN => n14943);
   U19729 : XNOR2_X1 port map( A => n17937, B => n17936, ZN => n25459);
   U19730 : INV_X1 port map( A => n997, ZN => n25460);
   U19868 : BUF_X1 port map( A => n22220, Z => n25461);
   U19876 : XNOR2_X1 port map( A => n21305, B => n21304, ZN => n22220);
   U19976 : INV_X1 port map( A => n14721, ZN => n25518);
   U19985 : XNOR2_X1 port map( A => n2577, B => n5503, ZN => n25462);
   U20052 : XNOR2_X1 port map( A => n5503, B => n2577, ZN => n22782);
   U20053 : XNOR2_X1 port map( A => n9173, B => n9172, ZN => n25463);
   U20070 : XNOR2_X1 port map( A => n9173, B => n9172, ZN => n10137);
   U20317 : CLKBUF_X1 port map( A => n9554, Z => n25464);
   U20402 : OAI211_X1 port map( C1 => n16199, C2 => n3143, A => n16201, B => 
                           n3542, ZN => n25465);
   U20446 : XOR2_X1 port map( A => n11786, B => n11785, Z => n25466);
   U20566 : AND2_X1 port map( A1 => n24863, A2 => n25162, ZN => n25467);
   U20581 : OR2_X1 port map( A1 => n16771, A2 => n17039, ZN => n25468);
   U20594 : XOR2_X1 port map( A => n18699, B => n18698, Z => n25469);
   U20609 : CLKBUF_X1 port map( A => n22449, Z => n25471);
   U20628 : XNOR2_X1 port map( A => n17658, B => n17659, ZN => n25473);
   U20630 : XNOR2_X1 port map( A => n17658, B => n17659, ZN => n25474);
   U20707 : NOR2_X1 port map( A1 => n15832, A2 => n151, ZN => n17728);
   U20727 : XNOR2_X1 port map( A => n17658, B => n17659, ZN => n19487);
   U20729 : INV_X1 port map( A => n19326, ZN => n25566);
   U20788 : XNOR2_X1 port map( A => n8838, B => n8837, ZN => n25475);
   U20793 : AOI21_X1 port map( B1 => n19253, B2 => n24943, A => n3047, ZN => 
                           n25476);
   U20800 : AOI21_X1 port map( B1 => n19253, B2 => n24943, A => n3047, ZN => 
                           n25477);
   U20829 : XNOR2_X1 port map( A => n8838, B => n8837, ZN => n9491);
   U20834 : OAI211_X1 port map( C1 => n18726, C2 => n19376, A => n18725, B => 
                           n4317, ZN => n25478);
   U20857 : XOR2_X1 port map( A => n20988, B => n20987, Z => n25479);
   U20858 : NAND3_X2 port map( A1 => n2468, A2 => n2467, A3 => n2466, ZN => 
                           n21699);
   U20873 : XOR2_X1 port map( A => Key(165), B => Plaintext(165), Z => n25480);
   U20904 : NOR2_X1 port map( A1 => n4969, A2 => n4528, ZN => n25481);
   U20929 : NOR2_X1 port map( A1 => n4969, A2 => n4528, ZN => n25482);
   U20942 : NOR2_X1 port map( A1 => n4969, A2 => n4528, ZN => n18628);
   U20972 : BUF_X1 port map( A => n21477, Z => n25483);
   U20980 : OAI211_X1 port map( C1 => n20070, C2 => n20071, A => n1469, B => 
                           n24722, ZN => n21477);
   U21001 : XOR2_X1 port map( A => n14779, B => n14778, Z => n25484);
   U21031 : XNOR2_X1 port map( A => n20908, B => n5503, ZN => n25485);
   U21047 : XNOR2_X1 port map( A => n8190, B => n8189, ZN => n25486);
   U21097 : CLKBUF_X1 port map( A => n22453, Z => n25487);
   U21107 : OAI21_X1 port map( B1 => n22327, B2 => n22326, A => n3682, ZN => 
                           n25488);
   U21109 : XOR2_X1 port map( A => n18427, B => n18426, Z => n25489);
   U21110 : NOR2_X1 port map( A1 => n18791, A2 => n18792, ZN => n25490);
   U21132 : NOR2_X1 port map( A1 => n18791, A2 => n18792, ZN => n20054);
   U21133 : XNOR2_X2 port map( A => n14717, B => n14718, ZN => n16101);
   U21161 : AOI21_X2 port map( B1 => n10380, B2 => n4928, A => n1418, ZN => 
                           n12207);
   U21175 : XNOR2_X2 port map( A => n861, B => n11926, ZN => n13318);
   U21191 : OAI21_X2 port map( B1 => n3964, B2 => n13729, A => n3298, ZN => 
                           n15071);
   U21208 : OAI211_X1 port map( C1 => n15870, C2 => n16802, A => n25129, B => 
                           n24685, ZN => n25493);
   U21216 : OAI211_X1 port map( C1 => n15870, C2 => n16802, A => n25129, B => 
                           n24685, ZN => n18636);
   U21253 : XOR2_X1 port map( A => n11605, B => n11606, Z => n25494);
   U21310 : XNOR2_X1 port map( A => n21429, B => n21633, ZN => n25495);
   U21319 : OR3_X1 port map( A1 => n25253, A2 => n7449, A3 => n7917, ZN => 
                           n3346);
   U21320 : CLKBUF_X1 port map( A => n21368, Z => n25496);
   U21321 : INV_X1 port map( A => n13151, ZN => n13148);
   U21422 : OAI21_X1 port map( B1 => n9865, B2 => n9864, A => n9863, ZN => 
                           n25497);
   U21465 : NOR2_X1 port map( A1 => n19509, A2 => n19508, ZN => n25498);
   U21469 : NOR2_X1 port map( A1 => n19509, A2 => n19508, ZN => n21659);
   U21470 : XNOR2_X1 port map( A => n11919, B => n11918, ZN => n25499);
   U21482 : XNOR2_X1 port map( A => n13576, B => n13577, ZN => n25500);
   U21524 : BUF_X1 port map( A => n15515, Z => n25501);
   U21525 : XOR2_X1 port map( A => n13939, B => n13938, Z => n25502);
   U21561 : NAND2_X1 port map( A1 => n1054, A2 => n10895, ZN => n10898);
   U21591 : NAND2_X1 port map( A1 => n14077, A2 => n14075, ZN => n769);
   U21593 : NAND3_X1 port map( A1 => n25505, A2 => n25504, A3 => n25503, ZN => 
                           n15274);
   U21597 : NAND2_X1 port map( A1 => n2122, A2 => n14079, ZN => n25503);
   U21601 : NAND2_X1 port map( A1 => n14080, A2 => n12704, ZN => n25505);
   U21630 : OAI21_X1 port map( B1 => n10585, B2 => n25507, A => n25506, ZN => 
                           n9444);
   U21665 : NAND2_X1 port map( A1 => n10585, A2 => n10375, ZN => n25506);
   U21677 : NAND2_X1 port map( A1 => n25509, A2 => n25508, ZN => n1674);
   U21701 : INV_X1 port map( A => n15625, ZN => n25510);
   U21717 : NAND4_X2 port map( A1 => n5076, A2 => n5075, A3 => n1163, A4 => 
                           n1164, ZN => n23779);
   U21916 : NAND3_X1 port map( A1 => n13282, A2 => n24988, A3 => n25191, ZN => 
                           n12610);
   U21933 : NAND2_X1 port map( A1 => n23814, A2 => n23815, ZN => n24630);
   U21954 : NAND2_X1 port map( A1 => n18134, A2 => n18135, ZN => n20328);
   U21983 : NAND2_X1 port map( A1 => n25512, A2 => n25511, ZN => n24879);
   U22002 : NAND2_X1 port map( A1 => n5421, A2 => n22038, ZN => n25511);
   U22016 : NAND2_X1 port map( A1 => n22037, A2 => n603, ZN => n25512);
   U22070 : NAND4_X2 port map( A1 => n15313, A2 => n4440, A3 => n15311, A4 => 
                           n15312, ZN => n15314);
   U22115 : OR2_X1 port map( A1 => n9851, A2 => n9853, ZN => n8419);
   U22128 : NOR2_X1 port map( A1 => n9592, A2 => n10158, ZN => n9853);
   U22177 : OAI21_X1 port map( B1 => n19883, B2 => n25514, A => n25513, ZN => 
                           n19120);
   U22178 : NAND2_X1 port map( A1 => n19883, A2 => n20111, ZN => n25513);
   U22230 : INV_X1 port map( A => n20109, ZN => n25514);
   U22339 : NAND2_X1 port map( A1 => n5409, A2 => n17425, ZN => n16644);
   U22361 : NOR2_X2 port map( A1 => n1887, A2 => n25515, ZN => n12241);
   U22497 : NAND2_X1 port map( A1 => n4999, A2 => n5000, ZN => n25515);
   U22541 : NAND2_X1 port map( A1 => n22711, A2 => n21020, ZN => n24781);
   U22552 : XNOR2_X1 port map( A => n25516, B => n452, ZN => Ciphertext(96));
   U22591 : OAI21_X2 port map( B1 => n20275, B2 => n20276, A => n25519, ZN => 
                           n21658);
   U22597 : NAND2_X1 port map( A1 => n3520, A2 => n3521, ZN => n25519);
   U22608 : NAND2_X1 port map( A1 => n16138, A2 => n24747, ZN => n25077);
   U22616 : NAND2_X1 port map( A1 => n1836, A2 => n4015, ZN => n24976);
   U22684 : NAND2_X1 port map( A1 => n25523, A2 => n25520, ZN => n8383);
   U22685 : NAND2_X1 port map( A1 => n25522, A2 => n25521, ZN => n25520);
   U22687 : INV_X1 port map( A => n9837, ZN => n25521);
   U22688 : NAND2_X1 port map( A1 => n421, A2 => n10099, ZN => n25522);
   U22735 : NAND2_X1 port map( A1 => n8381, A2 => n9837, ZN => n25523);
   U22740 : OR2_X1 port map( A1 => n20290, A2 => n20291, ZN => n24116);
   U22764 : XNOR2_X2 port map( A => n21026, B => n21243, ZN => n22243);
   U22801 : AOI22_X1 port map( A1 => n23805, A2 => n23003, B1 => n25525, B2 => 
                           n23005, ZN => n23006);
   U22844 : NOR2_X1 port map( A1 => n2411, A2 => n23790, ZN => n25525);
   U22897 : NAND3_X1 port map( A1 => n10286, A2 => n11112, A3 => n11113, ZN => 
                           n2752);
   U22904 : NAND3_X1 port map( A1 => n23681, A2 => n23678, A3 => n23679, ZN => 
                           n23680);
   U22906 : NAND2_X1 port map( A1 => n25526, A2 => n15957, ZN => n18557);
   U22907 : NAND3_X1 port map( A1 => n1909, A2 => n284, A3 => n1908, ZN => 
                           n25526);
   U22915 : NAND2_X1 port map( A1 => n6364, A2 => n25527, ZN => n7713);
   U22944 : NAND2_X1 port map( A1 => n16461, A2 => n16466, ZN => n3271);
   U22972 : NAND2_X1 port map( A1 => n25529, A2 => n25528, ZN => n12948);
   U22989 : NAND2_X1 port map( A1 => n13317, A2 => n12945, ZN => n25528);
   U22992 : NAND2_X1 port map( A1 => n12946, A2 => n25530, ZN => n25529);
   U22994 : INV_X1 port map( A => n13317, ZN => n25530);
   U22998 : NAND3_X1 port map( A1 => n13619, A2 => n4771, A3 => n14852, ZN => 
                           n4768);
   U23051 : NAND3_X1 port map( A1 => n13054, A2 => n408, A3 => n13055, ZN => 
                           n715);
   U23087 : AND3_X2 port map( A1 => n25532, A2 => n22172, A3 => n25531, ZN => 
                           n23689);
   U23115 : NAND2_X1 port map( A1 => n4064, A2 => n22918, ZN => n25531);
   U23116 : NAND2_X1 port map( A1 => n4063, A2 => n22170, ZN => n25532);
   U23147 : NAND2_X1 port map( A1 => n20103, A2 => n20102, ZN => n20099);
   U23312 : NAND2_X1 port map( A1 => n746, A2 => n25533, ZN => n2419);
   U23324 : NOR2_X1 port map( A1 => n25502, A2 => n16397, ZN => n25533);
   U23325 : NAND3_X1 port map( A1 => n22454, A2 => n24496, A3 => n22453, ZN => 
                           n2188);
   U23389 : NAND3_X1 port map( A1 => n25534, A2 => n3404, A3 => n5256, ZN => 
                           n3369);
   U23396 : NAND2_X1 port map( A1 => n14458, A2 => n14317, ZN => n25534);
   U23532 : NAND3_X1 port map( A1 => n4537, A2 => n4534, A3 => n25535, ZN => 
                           n24648);
   U23615 : NAND3_X1 port map( A1 => n1238, A2 => n22222, A3 => n1728, ZN => 
                           n24832);
   U23617 : NAND2_X1 port map( A1 => n2918, A2 => n12580, ZN => n12581);
   U23662 : NAND3_X1 port map( A1 => n23452, A2 => n23425, A3 => n3242, ZN => 
                           n23447);
   U23756 : NAND2_X1 port map( A1 => n5703, A2 => n6984, ZN => n8499);
   U23757 : NAND3_X2 port map( A1 => n25537, A2 => n2955, A3 => n25536, ZN => 
                           n15486);
   U23889 : NAND2_X1 port map( A1 => n3533, A2 => n13426, ZN => n25536);
   U24006 : NAND2_X1 port map( A1 => n1744, A2 => n1742, ZN => n25538);
   U24023 : NAND2_X1 port map( A1 => n24144, A2 => n9208, ZN => n135);
   U24026 : NAND2_X1 port map( A1 => n2068, A2 => n19106, ZN => n2463);
   U24083 : OAI21_X1 port map( B1 => n19760, B2 => n18385, A => n25195, ZN => 
                           n25539);
   U24140 : OAI21_X1 port map( B1 => n10453, B2 => n10756, A => n10452, ZN => 
                           n10454);
   U24141 : NAND2_X1 port map( A1 => n10756, A2 => n3324, ZN => n10452);
   U24142 : NAND2_X1 port map( A1 => n24639, A2 => n24642, ZN => n13538);
   U24150 : NAND3_X2 port map( A1 => n4388, A2 => n4387, A3 => n13276, ZN => 
                           n14251);
   U24151 : NAND2_X1 port map( A1 => n5047, A2 => n25542, ZN => n24325);
   U24152 : NAND2_X1 port map( A1 => n21379, A2 => n25543, ZN => n25542);
   U24169 : INV_X1 port map( A => n274, ZN => n25543);
   U24180 : NAND2_X1 port map( A1 => n2394, A2 => n2395, ZN => n21379);
   U24188 : OAI211_X2 port map( C1 => n3642, C2 => n22678, A => n3640, B => 
                           n25544, ZN => n23967);
   U24189 : NAND2_X1 port map( A1 => n22676, A2 => n23997, ZN => n25544);
   U24203 : NAND3_X2 port map( A1 => n3029, A2 => n5492, A3 => n3028, ZN => 
                           n11302);
   U24208 : NAND2_X1 port map( A1 => n5049, A2 => n22444, ZN => n24627);
   U24215 : NAND2_X1 port map( A1 => n20093, A2 => n25545, ZN => n24845);
   U24216 : INV_X1 port map( A => n25220, ZN => n25545);
   U24224 : NAND2_X1 port map( A1 => n23319, A2 => n23317, ZN => n2668);
   U24228 : NAND3_X1 port map( A1 => n1682, A2 => n1684, A3 => n23311, ZN => 
                           n23319);
   U24240 : AND3_X2 port map( A1 => n5178, A2 => n5176, A3 => n5177, ZN => 
                           n17171);
   U24244 : NAND3_X1 port map( A1 => n3625, A2 => n3624, A3 => n2861, ZN => 
                           n25561);
   U24248 : NAND2_X1 port map( A1 => n6730, A2 => n6733, ZN => n5001);
   U24249 : AND2_X2 port map( A1 => n24518, A2 => n24517, ZN => n23969);
   U24262 : NAND2_X1 port map( A1 => n20417, A2 => n20419, ZN => n20418);
   U24282 : NAND3_X1 port map( A1 => n24919, A2 => n24456, A3 => n25546, ZN => 
                           n19);
   U24298 : NAND2_X1 port map( A1 => n19006, A2 => n19007, ZN => n19008);
   U24302 : NAND3_X1 port map( A1 => n24664, A2 => n24572, A3 => n14060, ZN => 
                           n4222);
   U24305 : NAND2_X1 port map( A1 => n14059, A2 => n14850, ZN => n14060);
   U24310 : NAND3_X2 port map( A1 => n25547, A2 => n10843, A3 => n10842, ZN => 
                           n12381);
   U24316 : NAND3_X1 port map( A1 => n2967, A2 => n11135, A3 => n10839, ZN => 
                           n25547);
   U24330 : NAND3_X1 port map( A1 => n13307, A2 => n13304, A3 => n12613, ZN => 
                           n4791);
   U24335 : NAND3_X2 port map( A1 => n5248, A2 => n5247, A3 => n5825, ZN => 
                           n7882);
   U24336 : NAND2_X1 port map( A1 => n6351, A2 => n24466, ZN => n6504);
   U24337 : NOR2_X1 port map( A1 => n25548, A2 => n10925, ZN => n8180);
   U24345 : NAND2_X1 port map( A1 => n14265, A2 => n13426, ZN => n25549);
   U24346 : NAND2_X1 port map( A1 => n22127, A2 => n22126, ZN => n23277);
   U24348 : INV_X1 port map( A => n23263, ZN => n25550);
   U24349 : AND2_X2 port map( A1 => n3567, A2 => n3618, ZN => n4400);
   U24350 : NAND3_X1 port map( A1 => n6765, A2 => n6766, A3 => n6764, ZN => 
                           n3567);
   U24351 : NAND2_X1 port map( A1 => n23069, A2 => n21239, ZN => n1304);
   U24352 : OAI21_X1 port map( B1 => n25552, B2 => n25551, A => n3065, ZN => 
                           n3064);
   U24353 : INV_X1 port map( A => n12752, ZN => n25552);
   U24354 : NAND2_X1 port map( A1 => n10919, A2 => n10918, ZN => n10921);
   U24355 : OAI21_X1 port map( B1 => n17040, B2 => n25058, A => n3949, ZN => 
                           n3955);
   U24356 : OAI211_X2 port map( C1 => n15893, C2 => n24587, A => n15892, B => 
                           n15891, ZN => n25058);
   U24357 : NAND2_X1 port map( A1 => n20185, A2 => n20191, ZN => n19662);
   U24358 : OR2_X1 port map( A1 => n25485, A2 => n21766, ZN => n22155);
   U24359 : AOI21_X1 port map( B1 => n25554, B2 => n25553, A => n22231, ZN => 
                           n4397);
   U24360 : NAND2_X1 port map( A1 => n22056, A2 => n22226, ZN => n25554);
   U24361 : NAND2_X1 port map( A1 => n20296, A2 => n20142, ZN => n25555);
   U24362 : NAND2_X1 port map( A1 => n20011, A2 => n20301, ZN => n25556);
   U24363 : NAND3_X1 port map( A1 => n20528, A2 => n20525, A3 => n55, ZN => 
                           n20526);
   U24364 : OAI21_X1 port map( B1 => n55, B2 => n20528, A => n25558, ZN => 
                           n3833);
   U24365 : NAND2_X1 port map( A1 => n7556, A2 => n25559, ZN => n9016);
   U24366 : NAND2_X1 port map( A1 => n3572, A2 => n3569, ZN => n25559);
   U24367 : NAND3_X1 port map( A1 => n14194, A2 => n13785, A3 => n25560, ZN => 
                           n4202);
   U24368 : XNOR2_X1 port map( A => n17782, B => n17781, ZN => n19097);
   U24369 : OR2_X2 port map( A1 => n3449, A2 => n15749, ZN => n2562);
   U24370 : NAND3_X1 port map( A1 => n3268, A2 => n7757, A3 => n432, ZN => 
                           n7544);
   U24371 : NAND2_X1 port map( A1 => n19522, A2 => n19523, ZN => n18796);
   U24372 : NAND2_X1 port map( A1 => n17028, A2 => n25003, ZN => n17398);
   U24373 : NAND2_X1 port map( A1 => n1069, A2 => n5324, ZN => n4332);
   U24374 : NAND2_X1 port map( A1 => n11112, A2 => n11117, ZN => n9581);
   U24375 : NAND2_X1 port map( A1 => n244, A2 => n16426, ZN => n15649);
   U24376 : AOI22_X1 port map( A1 => n1550, A2 => n20486, B1 => n20485, B2 => 
                           n20913, ZN => n20490);
   U24377 : AND3_X2 port map( A1 => n3311, A2 => n6778, A3 => n6779, ZN => 
                           n7972);
   U24378 : NAND2_X1 port map( A1 => n25561, A2 => n3622, ZN => n24794);
   U24379 : NAND2_X1 port map( A1 => n4686, A2 => n17109, ZN => n25562);
   U24380 : NAND2_X1 port map( A1 => n19332, A2 => n25563, ZN => n19937);
   U24381 : NAND2_X1 port map( A1 => n25565, A2 => n25564, ZN => n25563);
   U24382 : AOI21_X1 port map( B1 => n24516, B2 => n19326, A => n4291, ZN => 
                           n25564);
   U24383 : NAND2_X1 port map( A1 => n19327, A2 => n25566, ZN => n25565);
   U24384 : NAND2_X1 port map( A1 => n25249, A2 => n10714, ZN => n10293);
   U24385 : NAND3_X2 port map( A1 => n9311, A2 => n25567, A3 => n9312, ZN => 
                           n10714);
   U24386 : OR2_X1 port map( A1 => n9313, A2 => n9314, ZN => n25567);
   U24387 : NAND2_X1 port map( A1 => n16100, A2 => n16101, ZN => n5458);
   U24388 : XNOR2_X2 port map( A => n14713, B => n14712, ZN => n16100);
   U24389 : NAND3_X1 port map( A1 => n23881, A2 => n107, A3 => n23882, ZN => 
                           n24692);
   U24390 : NAND3_X1 port map( A1 => n23897, A2 => n23899, A3 => n23898, ZN => 
                           n23901);
   U24391 : NAND2_X1 port map( A1 => n24825, A2 => n16072, ZN => n16133);
   U24392 : NAND3_X1 port map( A1 => n4487, A2 => n17255, A3 => n16942, ZN => 
                           n3189);
   U24393 : NAND2_X1 port map( A1 => n22901, A2 => n25569, ZN => n25568);
   U24394 : NAND2_X1 port map( A1 => n11837, A2 => n4499, ZN => n25570);
   U24395 : XNOR2_X1 port map( A => n25571, B => n21391, ZN => Ciphertext(21));
   U24396 : NAND3_X1 port map( A1 => n4627, A2 => n4628, A3 => n4626, ZN => 
                           n25571);
   U24397 : MUX2_X1 port map( A => n20567, B => n20560, S => n20561, Z => 
                           n20098);
   U24398 : NAND3_X1 port map( A1 => n25573, A2 => n2062, A3 => n25572, ZN => 
                           n3993);
   U24399 : NAND2_X1 port map( A1 => n2064, A2 => n287, ZN => n25573);
   U24400 : OAI21_X1 port map( B1 => n22426, B2 => n22125, A => n25574, ZN => 
                           n21876);
   U24401 : NAND2_X1 port map( A1 => n24322, A2 => n22422, ZN => n25574);
   U24402 : OR2_X1 port map( A1 => n16365, A2 => n17183, ZN => n15817);
   U24403 : AND2_X2 port map( A1 => n25576, A2 => n25575, ZN => n16796);
   U24404 : NAND2_X2 port map( A1 => n25577, A2 => n2802, ZN => n19986);
   U24405 : NAND3_X1 port map( A1 => n19149, A2 => n19150, A3 => n19266, ZN => 
                           n25577);
   U24406 : NAND3_X1 port map( A1 => n5285, A2 => n5287, A3 => n22090, ZN => 
                           Ciphertext(132));
   U24407 : NAND2_X1 port map( A1 => n25578, A2 => n21067, ZN => n21071);
   U24408 : OAI21_X1 port map( B1 => n21066, B2 => n21065, A => n25579, ZN => 
                           n25578);
   U24409 : NAND3_X1 port map( A1 => n22581, A2 => n4989, A3 => n4990, ZN => 
                           n24789);
   U24410 : NAND2_X1 port map( A1 => n21825, A2 => n21822, ZN => n3856);
   U24411 : XNOR2_X2 port map( A => n18861, B => n18860, ZN => n21822);
   U24412 : NAND3_X2 port map( A1 => n14238, A2 => n1342, A3 => n1343, ZN => 
                           n15369);
   U24413 : NAND2_X1 port map( A1 => n25580, A2 => n24198, ZN => n8853);
   U24414 : NAND2_X1 port map( A1 => n7470, A2 => n25154, ZN => n25580);
   U24415 : NAND2_X1 port map( A1 => n2718, A2 => n15811, ZN => n42);
   U24416 : NAND2_X1 port map( A1 => n24061, A2 => n16403, ZN => n2718);
   U24417 : NAND2_X1 port map( A1 => n10960, A2 => n4998, ZN => n10963);
   U24418 : NAND2_X1 port map( A1 => n25583, A2 => n25581, ZN => n12628);
   U24419 : NAND2_X1 port map( A1 => n13364, A2 => n25582, ZN => n25581);
   U24420 : NOR2_X1 port map( A1 => n12977, A2 => n12980, ZN => n25582);
   U24421 : NAND2_X1 port map( A1 => n25584, A2 => n12624, ZN => n25583);
   U24422 : INV_X1 port map( A => n13364, ZN => n25584);
   U24423 : NAND2_X1 port map( A1 => n25587, A2 => n25585, ZN => n16088);
   U24424 : INV_X1 port map( A => n16080, ZN => n25586);
   U24425 : NOR2_X1 port map( A1 => n1737, A2 => n7721, ZN => n1736);
   U24426 : NAND3_X1 port map( A1 => n269, A2 => n8531, A3 => n7087, ZN => 
                           n7089);
   U24427 : OAI211_X1 port map( C1 => n16340, C2 => n16339, A => n25589, B => 
                           n25588, ZN => n16527);
   U24428 : NAND2_X1 port map( A1 => n16337, A2 => n16336, ZN => n25588);
   U24429 : NAND2_X1 port map( A1 => n16335, A2 => n16334, ZN => n25589);
   U24430 : NAND2_X1 port map( A1 => n25590, A2 => n6525, ZN => n7662);
   U24431 : NAND3_X1 port map( A1 => n1321, A2 => n1320, A3 => n6520, ZN => 
                           n25590);
   U24432 : OAI211_X1 port map( C1 => n15961, C2 => n1329, A => n16424, B => 
                           n25591, ZN => n17436);
   U24433 : NAND3_X1 port map( A1 => n3847, A2 => n3848, A3 => n24487, ZN => 
                           n25592);
   U24434 : NAND2_X1 port map( A1 => n4973, A2 => n4755, ZN => n4751);
   U24435 : XNOR2_X1 port map( A => n25593, B => n15319, ZN => n5494);
   U24436 : XNOR2_X1 port map( A => n15317, B => n15318, ZN => n25593);
   U24437 : NAND3_X1 port map( A1 => n22548, A2 => n25595, A3 => n25594, ZN => 
                           n22550);
   U24438 : NAND2_X1 port map( A1 => n22547, A2 => n23906, ZN => n25594);
   U24439 : NAND2_X1 port map( A1 => n22546, A2 => n23879, ZN => n25595);
   U24440 : NOR2_X1 port map( A1 => n19012, A2 => n19689, ZN => n19020);
   U24441 : NAND3_X1 port map( A1 => n16458, A2 => n16459, A3 => n25596, ZN => 
                           n4724);
   U24442 : NOR2_X1 port map( A1 => n22224, A2 => n25597, ZN => n23742);
   U24443 : NAND2_X1 port map( A1 => n24832, A2 => n1237, ZN => n25597);
   U24444 : AND2_X2 port map( A1 => n16055, A2 => n16054, ZN => n16375);
   U24445 : NAND2_X1 port map( A1 => n2322, A2 => n20533, ZN => n3076);
   U24446 : NAND2_X1 port map( A1 => n19687, A2 => n19688, ZN => n2322);
   U24447 : OAI211_X2 port map( C1 => n5360, C2 => n12830, A => n2631, B => 
                           n12608, ZN => n14850);
   U24448 : NAND3_X2 port map( A1 => n14396, A2 => n14395, A3 => n14394, ZN => 
                           n17283);
   U24449 : AOI22_X2 port map( A1 => n5244, A2 => n20477, B1 => n999, B2 => 
                           n18839, ZN => n25073);
   U24450 : XNOR2_X2 port map( A => n22018, B => n22017, ZN => n25041);
   U24451 : AND2_X2 port map( A1 => n5583, A2 => n5582, ZN => n24498);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Top is

   port( clk : in std_logic;  Plaintext, Key : in std_logic_vector (191 downto 
         0);  Ciphertext : out std_logic_vector (191 downto 0));

end SPEEDY_Top;

architecture SYN_Behavioral of SPEEDY_Top is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFRS_X1
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SPEEDY_Rounds6_0
      port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : 
            out std_logic_vector (191 downto 0));
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal reg_in_191_port, reg_in_190_port, reg_in_189_port, reg_in_188_port, 
      reg_in_187_port, reg_in_186_port, reg_in_185_port, reg_in_184_port, 
      reg_in_183_port, reg_in_182_port, reg_in_181_port, reg_in_180_port, 
      reg_in_179_port, reg_in_178_port, reg_in_177_port, reg_in_176_port, 
      reg_in_175_port, reg_in_174_port, reg_in_173_port, reg_in_172_port, 
      reg_in_171_port, reg_in_170_port, reg_in_169_port, reg_in_168_port, 
      reg_in_167_port, reg_in_166_port, reg_in_165_port, reg_in_164_port, 
      reg_in_163_port, reg_in_162_port, reg_in_161_port, reg_in_160_port, 
      reg_in_159_port, reg_in_158_port, reg_in_157_port, reg_in_156_port, 
      reg_in_155_port, reg_in_154_port, reg_in_153_port, reg_in_152_port, 
      reg_in_151_port, reg_in_150_port, reg_in_149_port, reg_in_148_port, 
      reg_in_147_port, reg_in_146_port, reg_in_145_port, reg_in_144_port, 
      reg_in_143_port, reg_in_142_port, reg_in_141_port, reg_in_140_port, 
      reg_in_139_port, reg_in_138_port, reg_in_137_port, reg_in_136_port, 
      reg_in_135_port, reg_in_134_port, reg_in_133_port, reg_in_132_port, 
      reg_in_131_port, reg_in_130_port, reg_in_129_port, reg_in_128_port, 
      reg_in_127_port, reg_in_126_port, reg_in_125_port, reg_in_124_port, 
      reg_in_123_port, reg_in_122_port, reg_in_121_port, reg_in_120_port, 
      reg_in_119_port, reg_in_118_port, reg_in_117_port, reg_in_116_port, 
      reg_in_115_port, reg_in_114_port, reg_in_113_port, reg_in_112_port, 
      reg_in_111_port, reg_in_110_port, reg_in_109_port, reg_in_108_port, 
      reg_in_107_port, reg_in_106_port, reg_in_105_port, reg_in_104_port, 
      reg_in_103_port, reg_in_102_port, reg_in_101_port, reg_in_100_port, 
      reg_in_99_port, reg_in_98_port, reg_in_97_port, reg_in_96_port, 
      reg_in_95_port, reg_in_94_port, reg_in_93_port, reg_in_92_port, 
      reg_in_91_port, reg_in_90_port, reg_in_89_port, reg_in_88_port, 
      reg_in_87_port, reg_in_86_port, reg_in_85_port, reg_in_84_port, 
      reg_in_83_port, reg_in_82_port, reg_in_81_port, reg_in_80_port, 
      reg_in_79_port, reg_in_78_port, reg_in_77_port, reg_in_76_port, 
      reg_in_75_port, reg_in_74_port, reg_in_73_port, reg_in_72_port, 
      reg_in_71_port, reg_in_70_port, reg_in_69_port, reg_in_68_port, 
      reg_in_67_port, reg_in_66_port, reg_in_65_port, reg_in_64_port, 
      reg_in_63_port, reg_in_62_port, reg_in_61_port, reg_in_60_port, 
      reg_in_59_port, reg_in_58_port, reg_in_57_port, reg_in_56_port, 
      reg_in_55_port, reg_in_54_port, reg_in_53_port, reg_in_52_port, 
      reg_in_51_port, reg_in_50_port, reg_in_49_port, reg_in_48_port, 
      reg_in_47_port, reg_in_46_port, reg_in_45_port, reg_in_44_port, 
      reg_in_43_port, reg_in_42_port, reg_in_41_port, reg_in_40_port, 
      reg_in_39_port, reg_in_38_port, reg_in_37_port, reg_in_36_port, 
      reg_in_35_port, reg_in_34_port, reg_in_33_port, reg_in_32_port, 
      reg_in_31_port, reg_in_30_port, reg_in_29_port, reg_in_28_port, 
      reg_in_27_port, reg_in_26_port, reg_in_25_port, reg_in_24_port, 
      reg_in_23_port, reg_in_22_port, reg_in_21_port, reg_in_20_port, 
      reg_in_19_port, reg_in_18_port, reg_in_17_port, reg_in_16_port, 
      reg_in_15_port, reg_in_14_port, reg_in_13_port, reg_in_12_port, 
      reg_in_11_port, reg_in_10_port, reg_in_9_port, reg_in_8_port, 
      reg_in_7_port, reg_in_6_port, reg_in_5_port, reg_in_4_port, reg_in_3_port
      , reg_in_2_port, reg_in_1_port, reg_in_0_port, reg_key_191_port, 
      reg_key_190_port, reg_key_189_port, reg_key_188_port, reg_key_187_port, 
      reg_key_186_port, reg_key_185_port, reg_key_184_port, reg_key_183_port, 
      reg_key_182_port, reg_key_181_port, reg_key_180_port, reg_key_179_port, 
      reg_key_178_port, reg_key_177_port, reg_key_176_port, reg_key_175_port, 
      reg_key_174_port, reg_key_173_port, reg_key_172_port, reg_key_171_port, 
      reg_key_170_port, reg_key_169_port, reg_key_168_port, reg_key_167_port, 
      reg_key_166_port, reg_key_165_port, reg_key_164_port, reg_key_163_port, 
      reg_key_162_port, reg_key_161_port, reg_key_160_port, reg_key_159_port, 
      reg_key_158_port, reg_key_157_port, reg_key_156_port, reg_key_155_port, 
      reg_key_154_port, reg_key_153_port, reg_key_152_port, reg_key_151_port, 
      reg_key_150_port, reg_key_149_port, reg_key_148_port, reg_key_147_port, 
      reg_key_146_port, reg_key_145_port, reg_key_144_port, reg_key_143_port, 
      reg_key_142_port, reg_key_141_port, reg_key_140_port, reg_key_139_port, 
      reg_key_138_port, reg_key_137_port, reg_key_136_port, reg_key_135_port, 
      reg_key_134_port, reg_key_133_port, reg_key_132_port, reg_key_131_port, 
      reg_key_130_port, reg_key_129_port, reg_key_128_port, reg_key_127_port, 
      reg_key_126_port, reg_key_125_port, reg_key_124_port, reg_key_123_port, 
      reg_key_122_port, reg_key_121_port, reg_key_120_port, reg_key_119_port, 
      reg_key_118_port, reg_key_117_port, reg_key_116_port, reg_key_115_port, 
      reg_key_114_port, reg_key_113_port, reg_key_112_port, reg_key_111_port, 
      reg_key_110_port, reg_key_109_port, reg_key_108_port, reg_key_107_port, 
      reg_key_106_port, reg_key_105_port, reg_key_104_port, reg_key_103_port, 
      reg_key_102_port, reg_key_101_port, reg_key_100_port, reg_key_99_port, 
      reg_key_98_port, reg_key_97_port, reg_key_96_port, reg_key_95_port, 
      reg_key_94_port, reg_key_93_port, reg_key_92_port, reg_key_91_port, 
      reg_key_90_port, reg_key_89_port, reg_key_88_port, reg_key_87_port, 
      reg_key_86_port, reg_key_85_port, reg_key_84_port, reg_key_83_port, 
      reg_key_82_port, reg_key_81_port, reg_key_80_port, reg_key_79_port, 
      reg_key_78_port, reg_key_77_port, reg_key_76_port, reg_key_75_port, 
      reg_key_74_port, reg_key_73_port, reg_key_72_port, reg_key_71_port, 
      reg_key_70_port, reg_key_69_port, reg_key_68_port, reg_key_67_port, 
      reg_key_66_port, reg_key_65_port, reg_key_64_port, reg_key_63_port, 
      reg_key_62_port, reg_key_61_port, reg_key_60_port, reg_key_59_port, 
      reg_key_58_port, reg_key_57_port, reg_key_56_port, reg_key_55_port, 
      reg_key_54_port, reg_key_53_port, reg_key_52_port, reg_key_51_port, 
      reg_key_50_port, reg_key_49_port, reg_key_48_port, reg_key_47_port, 
      reg_key_46_port, reg_key_45_port, reg_key_44_port, reg_key_43_port, 
      reg_key_42_port, reg_key_41_port, reg_key_40_port, reg_key_39_port, 
      reg_key_38_port, reg_key_37_port, reg_key_36_port, reg_key_35_port, 
      reg_key_34_port, reg_key_33_port, reg_key_32_port, reg_key_31_port, 
      reg_key_30_port, reg_key_29_port, reg_key_28_port, reg_key_27_port, 
      reg_key_26_port, reg_key_25_port, reg_key_24_port, reg_key_23_port, 
      reg_key_22_port, reg_key_21_port, reg_key_20_port, reg_key_19_port, 
      reg_key_18_port, reg_key_17_port, reg_key_16_port, reg_key_15_port, 
      reg_key_14_port, reg_key_13_port, reg_key_12_port, reg_key_11_port, 
      reg_key_10_port, reg_key_9_port, reg_key_8_port, reg_key_7_port, 
      reg_key_6_port, reg_key_5_port, reg_key_4_port, reg_key_3_port, 
      reg_key_2_port, reg_key_1_port, reg_key_0_port, reg_out_191_port, 
      reg_out_190_port, reg_out_189_port, reg_out_188_port, reg_out_187_port, 
      reg_out_186_port, reg_out_185_port, reg_out_184_port, reg_out_183_port, 
      reg_out_182_port, reg_out_181_port, reg_out_180_port, reg_out_179_port, 
      reg_out_178_port, reg_out_177_port, reg_out_176_port, reg_out_175_port, 
      reg_out_174_port, reg_out_173_port, reg_out_172_port, reg_out_171_port, 
      reg_out_170_port, reg_out_169_port, reg_out_168_port, reg_out_167_port, 
      reg_out_166_port, reg_out_165_port, reg_out_164_port, reg_out_163_port, 
      reg_out_162_port, reg_out_161_port, reg_out_160_port, reg_out_159_port, 
      reg_out_158_port, reg_out_157_port, reg_out_156_port, reg_out_155_port, 
      reg_out_154_port, reg_out_153_port, reg_out_152_port, reg_out_151_port, 
      reg_out_150_port, reg_out_149_port, reg_out_148_port, reg_out_147_port, 
      reg_out_146_port, reg_out_145_port, reg_out_144_port, reg_out_143_port, 
      reg_out_142_port, reg_out_141_port, reg_out_140_port, reg_out_139_port, 
      reg_out_138_port, reg_out_137_port, reg_out_136_port, reg_out_135_port, 
      reg_out_134_port, reg_out_133_port, reg_out_132_port, reg_out_131_port, 
      reg_out_130_port, reg_out_129_port, reg_out_128_port, reg_out_127_port, 
      reg_out_126_port, reg_out_125_port, reg_out_124_port, reg_out_123_port, 
      reg_out_122_port, reg_out_121_port, reg_out_120_port, reg_out_119_port, 
      reg_out_118_port, reg_out_117_port, reg_out_116_port, reg_out_115_port, 
      reg_out_114_port, reg_out_113_port, reg_out_112_port, reg_out_111_port, 
      reg_out_110_port, reg_out_109_port, reg_out_108_port, reg_out_107_port, 
      reg_out_106_port, reg_out_105_port, reg_out_104_port, reg_out_103_port, 
      reg_out_102_port, reg_out_101_port, reg_out_100_port, reg_out_99_port, 
      reg_out_98_port, reg_out_97_port, reg_out_96_port, reg_out_95_port, 
      reg_out_94_port, reg_out_93_port, reg_out_92_port, reg_out_91_port, 
      reg_out_90_port, reg_out_89_port, reg_out_88_port, reg_out_87_port, 
      reg_out_86_port, reg_out_85_port, reg_out_84_port, reg_out_83_port, 
      reg_out_82_port, reg_out_81_port, reg_out_80_port, reg_out_79_port, 
      reg_out_78_port, reg_out_77_port, reg_out_76_port, reg_out_75_port, 
      reg_out_74_port, reg_out_73_port, reg_out_72_port, reg_out_71_port, 
      reg_out_70_port, reg_out_69_port, reg_out_68_port, reg_out_67_port, 
      reg_out_66_port, reg_out_65_port, reg_out_64_port, reg_out_63_port, 
      reg_out_62_port, reg_out_61_port, reg_out_60_port, reg_out_59_port, 
      reg_out_58_port, reg_out_57_port, reg_out_56_port, reg_out_55_port, 
      reg_out_54_port, reg_out_53_port, reg_out_52_port, reg_out_51_port, 
      reg_out_50_port, reg_out_49_port, reg_out_48_port, reg_out_47_port, 
      reg_out_46_port, reg_out_45_port, reg_out_44_port, reg_out_43_port, 
      reg_out_42_port, reg_out_41_port, reg_out_40_port, reg_out_39_port, 
      reg_out_38_port, reg_out_37_port, reg_out_36_port, reg_out_35_port, 
      reg_out_34_port, reg_out_33_port, reg_out_32_port, reg_out_31_port, 
      reg_out_30_port, reg_out_29_port, reg_out_28_port, reg_out_27_port, 
      reg_out_26_port, reg_out_25_port, reg_out_24_port, reg_out_23_port, 
      reg_out_22_port, reg_out_21_port, reg_out_20_port, reg_out_19_port, 
      reg_out_18_port, reg_out_17_port, reg_out_16_port, reg_out_15_port, 
      reg_out_14_port, reg_out_13_port, reg_out_12_port, reg_out_11_port, 
      reg_out_10_port, reg_out_9_port, reg_out_8_port, reg_out_7_port, 
      reg_out_6_port, reg_out_5_port, reg_out_4_port, reg_out_3_port, 
      reg_out_2_port, reg_out_1_port, reg_out_0_port, n9, n14, n15, n_1000, 
      n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, 
      n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, 
      n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, 
      n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, 
      n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, 
      n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, 
      n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, 
      n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, 
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, 
      n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, 
      n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, 
      n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, 
      n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, 
      n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, 
      n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, 
      n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, 
      n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, 
      n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, 
      n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, 
      n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, 
      n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, 
      n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, 
      n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, 
      n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, 
      n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, 
      n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, 
      n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, 
      n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, 
      n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, 
      n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, 
      n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, 
      n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, 
      n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, 
      n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, 
      n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, 
      n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, 
      n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, 
      n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, 
      n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, 
      n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, 
      n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, 
      n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, 
      n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575 : 
      std_logic;

begin
   
   reg_in_regx191x : DFF_X1 port map( D => Plaintext(191), CK => clk, Q => 
                           reg_in_191_port, QN => n_1000);
   reg_in_regx190x : DFF_X1 port map( D => Plaintext(190), CK => clk, Q => 
                           reg_in_190_port, QN => n_1001);
   reg_in_regx189x : DFF_X1 port map( D => Plaintext(189), CK => clk, Q => 
                           reg_in_189_port, QN => n_1002);
   reg_in_regx188x : DFF_X1 port map( D => Plaintext(188), CK => clk, Q => 
                           reg_in_188_port, QN => n_1003);
   reg_in_regx187x : DFF_X1 port map( D => Plaintext(187), CK => clk, Q => 
                           reg_in_187_port, QN => n_1004);
   reg_in_regx186x : DFF_X1 port map( D => Plaintext(186), CK => clk, Q => 
                           reg_in_186_port, QN => n_1005);
   reg_in_regx185x : DFF_X1 port map( D => Plaintext(185), CK => clk, Q => 
                           reg_in_185_port, QN => n_1006);
   reg_in_regx184x : DFF_X1 port map( D => Plaintext(184), CK => clk, Q => 
                           reg_in_184_port, QN => n_1007);
   reg_in_regx183x : DFF_X1 port map( D => Plaintext(183), CK => clk, Q => 
                           reg_in_183_port, QN => n_1008);
   reg_in_regx182x : DFF_X1 port map( D => Plaintext(182), CK => clk, Q => 
                           reg_in_182_port, QN => n_1009);
   reg_in_regx181x : DFF_X1 port map( D => Plaintext(181), CK => clk, Q => 
                           reg_in_181_port, QN => n_1010);
   reg_in_regx180x : DFF_X1 port map( D => Plaintext(180), CK => clk, Q => 
                           reg_in_180_port, QN => n_1011);
   reg_in_regx179x : DFF_X1 port map( D => Plaintext(179), CK => clk, Q => 
                           reg_in_179_port, QN => n_1012);
   reg_in_regx178x : DFF_X1 port map( D => Plaintext(178), CK => clk, Q => 
                           reg_in_178_port, QN => n_1013);
   reg_in_regx177x : DFF_X1 port map( D => Plaintext(177), CK => clk, Q => 
                           reg_in_177_port, QN => n_1014);
   reg_in_regx176x : DFF_X1 port map( D => Plaintext(176), CK => clk, Q => 
                           reg_in_176_port, QN => n_1015);
   reg_in_regx175x : DFF_X1 port map( D => Plaintext(175), CK => clk, Q => 
                           reg_in_175_port, QN => n_1016);
   reg_in_regx174x : DFF_X1 port map( D => Plaintext(174), CK => clk, Q => 
                           reg_in_174_port, QN => n_1017);
   reg_in_regx173x : DFF_X1 port map( D => Plaintext(173), CK => clk, Q => 
                           reg_in_173_port, QN => n_1018);
   reg_in_regx172x : DFF_X1 port map( D => Plaintext(172), CK => clk, Q => 
                           reg_in_172_port, QN => n_1019);
   reg_in_regx171x : DFF_X1 port map( D => Plaintext(171), CK => clk, Q => 
                           reg_in_171_port, QN => n_1020);
   reg_in_regx170x : DFF_X1 port map( D => Plaintext(170), CK => clk, Q => 
                           reg_in_170_port, QN => n_1021);
   reg_in_regx169x : DFF_X1 port map( D => Plaintext(169), CK => clk, Q => 
                           reg_in_169_port, QN => n_1022);
   reg_in_regx168x : DFF_X1 port map( D => Plaintext(168), CK => clk, Q => 
                           reg_in_168_port, QN => n_1023);
   reg_in_regx167x : DFF_X1 port map( D => Plaintext(167), CK => clk, Q => 
                           reg_in_167_port, QN => n_1024);
   reg_in_regx166x : DFF_X1 port map( D => Plaintext(166), CK => clk, Q => 
                           reg_in_166_port, QN => n_1025);
   reg_in_regx165x : DFF_X1 port map( D => Plaintext(165), CK => clk, Q => 
                           reg_in_165_port, QN => n_1026);
   reg_in_regx164x : DFF_X1 port map( D => Plaintext(164), CK => clk, Q => 
                           reg_in_164_port, QN => n_1027);
   reg_in_regx163x : DFF_X1 port map( D => Plaintext(163), CK => clk, Q => 
                           reg_in_163_port, QN => n_1028);
   reg_in_regx162x : DFF_X1 port map( D => Plaintext(162), CK => clk, Q => 
                           reg_in_162_port, QN => n_1029);
   reg_in_regx161x : DFF_X1 port map( D => Plaintext(161), CK => clk, Q => 
                           reg_in_161_port, QN => n_1030);
   reg_in_regx160x : DFF_X1 port map( D => Plaintext(160), CK => clk, Q => 
                           reg_in_160_port, QN => n_1031);
   reg_in_regx159x : DFF_X1 port map( D => Plaintext(159), CK => clk, Q => 
                           reg_in_159_port, QN => n_1032);
   reg_in_regx158x : DFF_X1 port map( D => Plaintext(158), CK => clk, Q => 
                           reg_in_158_port, QN => n_1033);
   reg_in_regx157x : DFF_X1 port map( D => Plaintext(157), CK => clk, Q => 
                           reg_in_157_port, QN => n_1034);
   reg_in_regx156x : DFF_X1 port map( D => Plaintext(156), CK => clk, Q => 
                           reg_in_156_port, QN => n_1035);
   reg_in_regx155x : DFF_X1 port map( D => Plaintext(155), CK => clk, Q => 
                           reg_in_155_port, QN => n_1036);
   reg_in_regx154x : DFF_X1 port map( D => Plaintext(154), CK => clk, Q => 
                           reg_in_154_port, QN => n_1037);
   reg_in_regx153x : DFF_X1 port map( D => Plaintext(153), CK => clk, Q => 
                           reg_in_153_port, QN => n_1038);
   reg_in_regx152x : DFF_X1 port map( D => Plaintext(152), CK => clk, Q => 
                           reg_in_152_port, QN => n_1039);
   reg_in_regx151x : DFF_X1 port map( D => Plaintext(151), CK => clk, Q => 
                           reg_in_151_port, QN => n_1040);
   reg_in_regx150x : DFF_X1 port map( D => Plaintext(150), CK => clk, Q => 
                           reg_in_150_port, QN => n_1041);
   reg_in_regx149x : DFF_X1 port map( D => Plaintext(149), CK => clk, Q => 
                           reg_in_149_port, QN => n_1042);
   reg_in_regx148x : DFF_X1 port map( D => Plaintext(148), CK => clk, Q => 
                           reg_in_148_port, QN => n_1043);
   reg_in_regx147x : DFF_X1 port map( D => Plaintext(147), CK => clk, Q => 
                           reg_in_147_port, QN => n_1044);
   reg_in_regx146x : DFF_X1 port map( D => Plaintext(146), CK => clk, Q => 
                           reg_in_146_port, QN => n_1045);
   reg_in_regx145x : DFF_X1 port map( D => Plaintext(145), CK => clk, Q => 
                           reg_in_145_port, QN => n_1046);
   reg_in_regx144x : DFF_X1 port map( D => Plaintext(144), CK => clk, Q => 
                           reg_in_144_port, QN => n_1047);
   reg_in_regx143x : DFF_X1 port map( D => Plaintext(143), CK => clk, Q => 
                           reg_in_143_port, QN => n_1048);
   reg_in_regx142x : DFF_X1 port map( D => Plaintext(142), CK => clk, Q => 
                           reg_in_142_port, QN => n_1049);
   reg_in_regx141x : DFF_X1 port map( D => Plaintext(141), CK => clk, Q => 
                           reg_in_141_port, QN => n_1050);
   reg_in_regx140x : DFF_X1 port map( D => Plaintext(140), CK => clk, Q => 
                           reg_in_140_port, QN => n_1051);
   reg_in_regx139x : DFF_X1 port map( D => Plaintext(139), CK => clk, Q => 
                           reg_in_139_port, QN => n_1052);
   reg_in_regx138x : DFF_X1 port map( D => Plaintext(138), CK => clk, Q => 
                           reg_in_138_port, QN => n_1053);
   reg_in_regx137x : DFF_X1 port map( D => Plaintext(137), CK => clk, Q => 
                           reg_in_137_port, QN => n_1054);
   reg_in_regx136x : DFF_X1 port map( D => Plaintext(136), CK => clk, Q => 
                           reg_in_136_port, QN => n_1055);
   reg_in_regx135x : DFF_X1 port map( D => Plaintext(135), CK => clk, Q => 
                           reg_in_135_port, QN => n_1056);
   reg_in_regx134x : DFF_X1 port map( D => Plaintext(134), CK => clk, Q => 
                           reg_in_134_port, QN => n_1057);
   reg_in_regx133x : DFF_X1 port map( D => Plaintext(133), CK => clk, Q => 
                           reg_in_133_port, QN => n_1058);
   reg_in_regx132x : DFF_X1 port map( D => Plaintext(132), CK => clk, Q => 
                           reg_in_132_port, QN => n_1059);
   reg_in_regx131x : DFF_X1 port map( D => Plaintext(131), CK => clk, Q => 
                           reg_in_131_port, QN => n_1060);
   reg_in_regx130x : DFF_X1 port map( D => Plaintext(130), CK => clk, Q => 
                           reg_in_130_port, QN => n_1061);
   reg_in_regx129x : DFF_X1 port map( D => Plaintext(129), CK => clk, Q => 
                           reg_in_129_port, QN => n_1062);
   reg_in_regx128x : DFF_X1 port map( D => Plaintext(128), CK => clk, Q => 
                           reg_in_128_port, QN => n_1063);
   reg_in_regx127x : DFF_X1 port map( D => Plaintext(127), CK => clk, Q => 
                           reg_in_127_port, QN => n_1064);
   reg_in_regx126x : DFF_X1 port map( D => Plaintext(126), CK => clk, Q => 
                           reg_in_126_port, QN => n_1065);
   reg_in_regx125x : DFF_X1 port map( D => Plaintext(125), CK => clk, Q => 
                           reg_in_125_port, QN => n_1066);
   reg_in_regx124x : DFF_X1 port map( D => Plaintext(124), CK => clk, Q => 
                           reg_in_124_port, QN => n_1067);
   reg_in_regx123x : DFF_X1 port map( D => Plaintext(123), CK => clk, Q => 
                           reg_in_123_port, QN => n_1068);
   reg_in_regx122x : DFF_X1 port map( D => Plaintext(122), CK => clk, Q => 
                           reg_in_122_port, QN => n_1069);
   reg_in_regx121x : DFF_X1 port map( D => Plaintext(121), CK => clk, Q => 
                           reg_in_121_port, QN => n_1070);
   reg_in_regx120x : DFF_X1 port map( D => Plaintext(120), CK => clk, Q => 
                           reg_in_120_port, QN => n_1071);
   reg_in_regx119x : DFF_X1 port map( D => Plaintext(119), CK => clk, Q => 
                           reg_in_119_port, QN => n_1072);
   reg_in_regx118x : DFF_X1 port map( D => Plaintext(118), CK => clk, Q => 
                           reg_in_118_port, QN => n_1073);
   reg_in_regx117x : DFF_X1 port map( D => Plaintext(117), CK => clk, Q => 
                           reg_in_117_port, QN => n_1074);
   reg_in_regx116x : DFF_X1 port map( D => Plaintext(116), CK => clk, Q => 
                           reg_in_116_port, QN => n_1075);
   reg_in_regx115x : DFF_X1 port map( D => Plaintext(115), CK => clk, Q => 
                           reg_in_115_port, QN => n_1076);
   reg_in_regx114x : DFF_X1 port map( D => Plaintext(114), CK => clk, Q => 
                           reg_in_114_port, QN => n_1077);
   reg_in_regx113x : DFF_X1 port map( D => Plaintext(113), CK => clk, Q => 
                           reg_in_113_port, QN => n_1078);
   reg_in_regx112x : DFF_X1 port map( D => Plaintext(112), CK => clk, Q => 
                           reg_in_112_port, QN => n_1079);
   reg_in_regx111x : DFF_X1 port map( D => Plaintext(111), CK => clk, Q => 
                           reg_in_111_port, QN => n_1080);
   reg_in_regx110x : DFF_X1 port map( D => Plaintext(110), CK => clk, Q => 
                           reg_in_110_port, QN => n_1081);
   reg_in_regx109x : DFF_X1 port map( D => Plaintext(109), CK => clk, Q => 
                           reg_in_109_port, QN => n_1082);
   reg_in_regx108x : DFF_X1 port map( D => Plaintext(108), CK => clk, Q => 
                           reg_in_108_port, QN => n_1083);
   reg_in_regx107x : DFF_X1 port map( D => Plaintext(107), CK => clk, Q => 
                           reg_in_107_port, QN => n_1084);
   reg_in_regx106x : DFF_X1 port map( D => Plaintext(106), CK => clk, Q => 
                           reg_in_106_port, QN => n_1085);
   reg_in_regx105x : DFF_X1 port map( D => Plaintext(105), CK => clk, Q => 
                           reg_in_105_port, QN => n_1086);
   reg_in_regx104x : DFF_X1 port map( D => Plaintext(104), CK => clk, Q => 
                           reg_in_104_port, QN => n_1087);
   reg_in_regx103x : DFF_X1 port map( D => Plaintext(103), CK => clk, Q => 
                           reg_in_103_port, QN => n_1088);
   reg_in_regx102x : DFF_X1 port map( D => Plaintext(102), CK => clk, Q => 
                           reg_in_102_port, QN => n_1089);
   reg_in_regx101x : DFF_X1 port map( D => Plaintext(101), CK => clk, Q => 
                           reg_in_101_port, QN => n_1090);
   reg_in_regx100x : DFF_X1 port map( D => Plaintext(100), CK => clk, Q => 
                           reg_in_100_port, QN => n_1091);
   reg_in_regx99x : DFF_X1 port map( D => Plaintext(99), CK => clk, Q => 
                           reg_in_99_port, QN => n_1092);
   reg_in_regx98x : DFF_X1 port map( D => Plaintext(98), CK => clk, Q => 
                           reg_in_98_port, QN => n_1093);
   reg_in_regx97x : DFF_X1 port map( D => Plaintext(97), CK => clk, Q => 
                           reg_in_97_port, QN => n_1094);
   reg_in_regx96x : DFF_X1 port map( D => Plaintext(96), CK => clk, Q => 
                           reg_in_96_port, QN => n_1095);
   reg_in_regx95x : DFF_X1 port map( D => Plaintext(95), CK => clk, Q => 
                           reg_in_95_port, QN => n_1096);
   reg_in_regx94x : DFF_X1 port map( D => Plaintext(94), CK => clk, Q => 
                           reg_in_94_port, QN => n_1097);
   reg_in_regx93x : DFF_X1 port map( D => Plaintext(93), CK => clk, Q => 
                           reg_in_93_port, QN => n_1098);
   reg_in_regx92x : DFF_X1 port map( D => Plaintext(92), CK => clk, Q => 
                           reg_in_92_port, QN => n_1099);
   reg_in_regx91x : DFF_X1 port map( D => Plaintext(91), CK => clk, Q => 
                           reg_in_91_port, QN => n_1100);
   reg_in_regx90x : DFF_X1 port map( D => Plaintext(90), CK => clk, Q => 
                           reg_in_90_port, QN => n_1101);
   reg_in_regx89x : DFF_X1 port map( D => Plaintext(89), CK => clk, Q => 
                           reg_in_89_port, QN => n_1102);
   reg_in_regx88x : DFF_X1 port map( D => Plaintext(88), CK => clk, Q => 
                           reg_in_88_port, QN => n_1103);
   reg_in_regx87x : DFF_X1 port map( D => Plaintext(87), CK => clk, Q => 
                           reg_in_87_port, QN => n_1104);
   reg_in_regx86x : DFF_X1 port map( D => Plaintext(86), CK => clk, Q => 
                           reg_in_86_port, QN => n_1105);
   reg_in_regx85x : DFF_X1 port map( D => Plaintext(85), CK => clk, Q => 
                           reg_in_85_port, QN => n_1106);
   reg_in_regx84x : DFF_X1 port map( D => Plaintext(84), CK => clk, Q => 
                           reg_in_84_port, QN => n_1107);
   reg_in_regx83x : DFF_X1 port map( D => Plaintext(83), CK => clk, Q => 
                           reg_in_83_port, QN => n_1108);
   reg_in_regx82x : DFF_X1 port map( D => Plaintext(82), CK => clk, Q => 
                           reg_in_82_port, QN => n_1109);
   reg_in_regx81x : DFF_X1 port map( D => Plaintext(81), CK => clk, Q => 
                           reg_in_81_port, QN => n_1110);
   reg_in_regx80x : DFF_X1 port map( D => Plaintext(80), CK => clk, Q => 
                           reg_in_80_port, QN => n_1111);
   reg_in_regx79x : DFF_X1 port map( D => Plaintext(79), CK => clk, Q => 
                           reg_in_79_port, QN => n_1112);
   reg_in_regx78x : DFF_X1 port map( D => Plaintext(78), CK => clk, Q => 
                           reg_in_78_port, QN => n_1113);
   reg_in_regx77x : DFF_X1 port map( D => Plaintext(77), CK => clk, Q => 
                           reg_in_77_port, QN => n_1114);
   reg_in_regx76x : DFF_X1 port map( D => Plaintext(76), CK => clk, Q => 
                           reg_in_76_port, QN => n_1115);
   reg_in_regx75x : DFF_X1 port map( D => Plaintext(75), CK => clk, Q => 
                           reg_in_75_port, QN => n_1116);
   reg_in_regx74x : DFF_X1 port map( D => Plaintext(74), CK => clk, Q => 
                           reg_in_74_port, QN => n_1117);
   reg_in_regx73x : DFF_X1 port map( D => Plaintext(73), CK => clk, Q => 
                           reg_in_73_port, QN => n_1118);
   reg_in_regx72x : DFF_X1 port map( D => Plaintext(72), CK => clk, Q => 
                           reg_in_72_port, QN => n_1119);
   reg_in_regx71x : DFF_X1 port map( D => Plaintext(71), CK => clk, Q => 
                           reg_in_71_port, QN => n_1120);
   reg_in_regx70x : DFF_X1 port map( D => Plaintext(70), CK => clk, Q => 
                           reg_in_70_port, QN => n_1121);
   reg_in_regx69x : DFF_X1 port map( D => Plaintext(69), CK => clk, Q => 
                           reg_in_69_port, QN => n_1122);
   reg_in_regx68x : DFF_X1 port map( D => Plaintext(68), CK => clk, Q => 
                           reg_in_68_port, QN => n_1123);
   reg_in_regx67x : DFF_X1 port map( D => Plaintext(67), CK => clk, Q => 
                           reg_in_67_port, QN => n_1124);
   reg_in_regx66x : DFF_X1 port map( D => Plaintext(66), CK => clk, Q => 
                           reg_in_66_port, QN => n_1125);
   reg_in_regx65x : DFF_X1 port map( D => Plaintext(65), CK => clk, Q => 
                           reg_in_65_port, QN => n_1126);
   reg_in_regx64x : DFF_X1 port map( D => Plaintext(64), CK => clk, Q => 
                           reg_in_64_port, QN => n_1127);
   reg_in_regx63x : DFF_X1 port map( D => Plaintext(63), CK => clk, Q => 
                           reg_in_63_port, QN => n_1128);
   reg_in_regx62x : DFF_X1 port map( D => Plaintext(62), CK => clk, Q => 
                           reg_in_62_port, QN => n_1129);
   reg_in_regx61x : DFF_X1 port map( D => Plaintext(61), CK => clk, Q => 
                           reg_in_61_port, QN => n_1130);
   reg_in_regx60x : DFF_X1 port map( D => Plaintext(60), CK => clk, Q => 
                           reg_in_60_port, QN => n_1131);
   reg_in_regx59x : DFF_X1 port map( D => Plaintext(59), CK => clk, Q => 
                           reg_in_59_port, QN => n_1132);
   reg_in_regx58x : DFF_X1 port map( D => Plaintext(58), CK => clk, Q => 
                           reg_in_58_port, QN => n_1133);
   reg_in_regx57x : DFF_X1 port map( D => Plaintext(57), CK => clk, Q => 
                           reg_in_57_port, QN => n_1134);
   reg_in_regx56x : DFF_X1 port map( D => Plaintext(56), CK => clk, Q => 
                           reg_in_56_port, QN => n_1135);
   reg_in_regx55x : DFF_X1 port map( D => Plaintext(55), CK => clk, Q => 
                           reg_in_55_port, QN => n_1136);
   reg_in_regx54x : DFF_X1 port map( D => Plaintext(54), CK => clk, Q => 
                           reg_in_54_port, QN => n_1137);
   reg_in_regx53x : DFF_X1 port map( D => Plaintext(53), CK => clk, Q => 
                           reg_in_53_port, QN => n_1138);
   reg_in_regx52x : DFF_X1 port map( D => Plaintext(52), CK => clk, Q => 
                           reg_in_52_port, QN => n_1139);
   reg_in_regx51x : DFF_X1 port map( D => Plaintext(51), CK => clk, Q => 
                           reg_in_51_port, QN => n_1140);
   reg_in_regx50x : DFF_X1 port map( D => Plaintext(50), CK => clk, Q => 
                           reg_in_50_port, QN => n_1141);
   reg_in_regx49x : DFF_X1 port map( D => Plaintext(49), CK => clk, Q => 
                           reg_in_49_port, QN => n_1142);
   reg_in_regx48x : DFF_X1 port map( D => Plaintext(48), CK => clk, Q => 
                           reg_in_48_port, QN => n_1143);
   reg_in_regx47x : DFF_X1 port map( D => Plaintext(47), CK => clk, Q => 
                           reg_in_47_port, QN => n_1144);
   reg_in_regx46x : DFF_X1 port map( D => Plaintext(46), CK => clk, Q => 
                           reg_in_46_port, QN => n_1145);
   reg_in_regx45x : DFF_X1 port map( D => Plaintext(45), CK => clk, Q => 
                           reg_in_45_port, QN => n_1146);
   reg_in_regx44x : DFF_X1 port map( D => Plaintext(44), CK => clk, Q => 
                           reg_in_44_port, QN => n_1147);
   reg_in_regx43x : DFF_X1 port map( D => Plaintext(43), CK => clk, Q => 
                           reg_in_43_port, QN => n_1148);
   reg_in_regx42x : DFF_X1 port map( D => Plaintext(42), CK => clk, Q => 
                           reg_in_42_port, QN => n_1149);
   reg_in_regx41x : DFF_X1 port map( D => Plaintext(41), CK => clk, Q => 
                           reg_in_41_port, QN => n_1150);
   reg_in_regx40x : DFF_X1 port map( D => Plaintext(40), CK => clk, Q => 
                           reg_in_40_port, QN => n_1151);
   reg_in_regx39x : DFF_X1 port map( D => Plaintext(39), CK => clk, Q => 
                           reg_in_39_port, QN => n_1152);
   reg_in_regx38x : DFF_X1 port map( D => Plaintext(38), CK => clk, Q => 
                           reg_in_38_port, QN => n_1153);
   reg_in_regx37x : DFF_X1 port map( D => Plaintext(37), CK => clk, Q => 
                           reg_in_37_port, QN => n_1154);
   reg_in_regx36x : DFF_X1 port map( D => Plaintext(36), CK => clk, Q => 
                           reg_in_36_port, QN => n_1155);
   reg_in_regx35x : DFF_X1 port map( D => Plaintext(35), CK => clk, Q => 
                           reg_in_35_port, QN => n_1156);
   reg_in_regx34x : DFF_X1 port map( D => Plaintext(34), CK => clk, Q => 
                           reg_in_34_port, QN => n_1157);
   reg_in_regx33x : DFF_X1 port map( D => Plaintext(33), CK => clk, Q => 
                           reg_in_33_port, QN => n_1158);
   reg_in_regx32x : DFF_X1 port map( D => Plaintext(32), CK => clk, Q => 
                           reg_in_32_port, QN => n_1159);
   reg_in_regx31x : DFF_X1 port map( D => Plaintext(31), CK => clk, Q => 
                           reg_in_31_port, QN => n_1160);
   reg_in_regx30x : DFF_X1 port map( D => Plaintext(30), CK => clk, Q => 
                           reg_in_30_port, QN => n_1161);
   reg_in_regx29x : DFF_X1 port map( D => Plaintext(29), CK => clk, Q => 
                           reg_in_29_port, QN => n_1162);
   reg_in_regx28x : DFF_X1 port map( D => Plaintext(28), CK => clk, Q => 
                           reg_in_28_port, QN => n_1163);
   reg_in_regx27x : DFF_X1 port map( D => Plaintext(27), CK => clk, Q => 
                           reg_in_27_port, QN => n_1164);
   reg_in_regx26x : DFF_X1 port map( D => Plaintext(26), CK => clk, Q => 
                           reg_in_26_port, QN => n_1165);
   reg_in_regx25x : DFF_X1 port map( D => Plaintext(25), CK => clk, Q => 
                           reg_in_25_port, QN => n_1166);
   reg_in_regx24x : DFF_X1 port map( D => Plaintext(24), CK => clk, Q => 
                           reg_in_24_port, QN => n_1167);
   reg_in_regx23x : DFF_X1 port map( D => Plaintext(23), CK => clk, Q => 
                           reg_in_23_port, QN => n_1168);
   reg_in_regx22x : DFF_X1 port map( D => Plaintext(22), CK => clk, Q => 
                           reg_in_22_port, QN => n_1169);
   reg_in_regx21x : DFF_X1 port map( D => Plaintext(21), CK => clk, Q => 
                           reg_in_21_port, QN => n_1170);
   reg_in_regx20x : DFF_X1 port map( D => Plaintext(20), CK => clk, Q => 
                           reg_in_20_port, QN => n_1171);
   reg_in_regx19x : DFF_X1 port map( D => Plaintext(19), CK => clk, Q => 
                           reg_in_19_port, QN => n_1172);
   reg_in_regx18x : DFF_X1 port map( D => Plaintext(18), CK => clk, Q => 
                           reg_in_18_port, QN => n_1173);
   reg_in_regx17x : DFF_X1 port map( D => Plaintext(17), CK => clk, Q => 
                           reg_in_17_port, QN => n_1174);
   reg_in_regx16x : DFF_X1 port map( D => Plaintext(16), CK => clk, Q => 
                           reg_in_16_port, QN => n_1175);
   reg_in_regx15x : DFF_X1 port map( D => Plaintext(15), CK => clk, Q => 
                           reg_in_15_port, QN => n_1176);
   reg_in_regx14x : DFF_X1 port map( D => Plaintext(14), CK => clk, Q => 
                           reg_in_14_port, QN => n_1177);
   reg_in_regx13x : DFF_X1 port map( D => Plaintext(13), CK => clk, Q => 
                           reg_in_13_port, QN => n_1178);
   reg_in_regx12x : DFF_X1 port map( D => Plaintext(12), CK => clk, Q => 
                           reg_in_12_port, QN => n_1179);
   reg_in_regx11x : DFF_X1 port map( D => Plaintext(11), CK => clk, Q => 
                           reg_in_11_port, QN => n_1180);
   reg_in_regx10x : DFF_X1 port map( D => Plaintext(10), CK => clk, Q => 
                           reg_in_10_port, QN => n_1181);
   reg_in_regx9x : DFF_X1 port map( D => Plaintext(9), CK => clk, Q => 
                           reg_in_9_port, QN => n_1182);
   reg_in_regx8x : DFF_X1 port map( D => Plaintext(8), CK => clk, Q => 
                           reg_in_8_port, QN => n_1183);
   reg_in_regx7x : DFF_X1 port map( D => Plaintext(7), CK => clk, Q => 
                           reg_in_7_port, QN => n_1184);
   reg_in_regx6x : DFF_X1 port map( D => Plaintext(6), CK => clk, Q => 
                           reg_in_6_port, QN => n_1185);
   reg_in_regx5x : DFF_X1 port map( D => Plaintext(5), CK => clk, Q => 
                           reg_in_5_port, QN => n_1186);
   reg_in_regx4x : DFF_X1 port map( D => Plaintext(4), CK => clk, Q => 
                           reg_in_4_port, QN => n_1187);
   reg_in_regx3x : DFF_X1 port map( D => Plaintext(3), CK => clk, Q => 
                           reg_in_3_port, QN => n_1188);
   reg_in_regx2x : DFF_X1 port map( D => Plaintext(2), CK => clk, Q => 
                           reg_in_2_port, QN => n_1189);
   reg_in_regx1x : DFF_X1 port map( D => Plaintext(1), CK => clk, Q => 
                           reg_in_1_port, QN => n_1190);
   reg_in_regx0x : DFF_X1 port map( D => Plaintext(0), CK => clk, Q => 
                           reg_in_0_port, QN => n_1191);
   reg_key_regx191x : DFF_X1 port map( D => Key(191), CK => clk, Q => 
                           reg_key_191_port, QN => n_1192);
   reg_key_regx190x : DFF_X1 port map( D => Key(190), CK => clk, Q => 
                           reg_key_190_port, QN => n_1193);
   reg_key_regx189x : DFF_X1 port map( D => Key(189), CK => clk, Q => 
                           reg_key_189_port, QN => n_1194);
   reg_key_regx188x : DFF_X1 port map( D => Key(188), CK => clk, Q => 
                           reg_key_188_port, QN => n_1195);
   reg_key_regx187x : DFF_X1 port map( D => Key(187), CK => clk, Q => 
                           reg_key_187_port, QN => n_1196);
   reg_key_regx184x : DFF_X1 port map( D => Key(184), CK => clk, Q => 
                           reg_key_184_port, QN => n_1197);
   reg_key_regx179x : DFF_X1 port map( D => Key(179), CK => clk, Q => 
                           reg_key_179_port, QN => n_1198);
   reg_key_regx178x : DFF_X1 port map( D => Key(178), CK => clk, Q => 
                           reg_key_178_port, QN => n_1199);
   reg_key_regx177x : DFF_X1 port map( D => Key(177), CK => clk, Q => 
                           reg_key_177_port, QN => n_1200);
   reg_key_regx173x : DFF_X1 port map( D => Key(173), CK => clk, Q => 
                           reg_key_173_port, QN => n_1201);
   reg_key_regx171x : DFF_X1 port map( D => Key(171), CK => clk, Q => 
                           reg_key_171_port, QN => n_1202);
   reg_key_regx169x : DFF_X1 port map( D => Key(169), CK => clk, Q => 
                           reg_key_169_port, QN => n_1203);
   reg_key_regx165x : DFF_X1 port map( D => Key(165), CK => clk, Q => 
                           reg_key_165_port, QN => n_1204);
   reg_key_regx160x : DFF_X1 port map( D => Key(160), CK => clk, Q => 
                           reg_key_160_port, QN => n_1205);
   reg_key_regx156x : DFF_X1 port map( D => Key(156), CK => clk, Q => 
                           reg_key_156_port, QN => n_1206);
   reg_key_regx151x : DFF_X1 port map( D => Key(151), CK => clk, Q => 
                           reg_key_151_port, QN => n_1207);
   reg_key_regx149x : DFF_X1 port map( D => Key(149), CK => clk, Q => 
                           reg_key_149_port, QN => n_1208);
   reg_key_regx143x : DFF_X1 port map( D => Key(143), CK => clk, Q => 
                           reg_key_143_port, QN => n_1209);
   reg_key_regx140x : DFF_X1 port map( D => Key(140), CK => clk, Q => 
                           reg_key_140_port, QN => n_1210);
   reg_key_regx137x : DFF_X1 port map( D => Key(137), CK => clk, Q => 
                           reg_key_137_port, QN => n_1211);
   reg_key_regx135x : DFF_X1 port map( D => Key(135), CK => clk, Q => 
                           reg_key_135_port, QN => n_1212);
   reg_key_regx132x : DFF_X1 port map( D => Key(132), CK => clk, Q => 
                           reg_key_132_port, QN => n_1213);
   reg_key_regx125x : DFF_X1 port map( D => Key(125), CK => clk, Q => 
                           reg_key_125_port, QN => n_1214);
   reg_key_regx123x : DFF_X1 port map( D => Key(123), CK => clk, Q => 
                           reg_key_123_port, QN => n_1215);
   reg_key_regx120x : DFF_X1 port map( D => Key(120), CK => clk, Q => 
                           reg_key_120_port, QN => n_1216);
   reg_key_regx119x : DFF_X1 port map( D => Key(119), CK => clk, Q => 
                           reg_key_119_port, QN => n_1217);
   reg_key_regx118x : DFF_X1 port map( D => Key(118), CK => clk, Q => 
                           reg_key_118_port, QN => n_1218);
   reg_key_regx109x : DFF_X1 port map( D => Key(109), CK => clk, Q => 
                           reg_key_109_port, QN => n_1219);
   reg_key_regx108x : DFF_X1 port map( D => Key(108), CK => clk, Q => 
                           reg_key_108_port, QN => n_1220);
   reg_key_regx105x : DFF_X1 port map( D => Key(105), CK => clk, Q => 
                           reg_key_105_port, QN => n_1221);
   reg_key_regx104x : DFF_X1 port map( D => Key(104), CK => clk, Q => 
                           reg_key_104_port, QN => n_1222);
   reg_key_regx103x : DFF_X1 port map( D => Key(103), CK => clk, Q => 
                           reg_key_103_port, QN => n_1223);
   reg_key_regx101x : DFF_X1 port map( D => Key(101), CK => clk, Q => 
                           reg_key_101_port, QN => n_1224);
   reg_key_regx100x : DFF_X1 port map( D => Key(100), CK => clk, Q => 
                           reg_key_100_port, QN => n_1225);
   reg_key_regx96x : DFF_X1 port map( D => Key(96), CK => clk, Q => 
                           reg_key_96_port, QN => n_1226);
   reg_key_regx95x : DFF_X1 port map( D => Key(95), CK => clk, Q => 
                           reg_key_95_port, QN => n_1227);
   reg_key_regx82x : DFF_X1 port map( D => Key(82), CK => clk, Q => 
                           reg_key_82_port, QN => n_1228);
   reg_key_regx81x : DFF_X1 port map( D => Key(81), CK => clk, Q => 
                           reg_key_81_port, QN => n_1229);
   reg_key_regx80x : DFF_X1 port map( D => Key(80), CK => clk, Q => 
                           reg_key_80_port, QN => n_1230);
   reg_key_regx76x : DFF_X1 port map( D => Key(76), CK => clk, Q => 
                           reg_key_76_port, QN => n_1231);
   reg_key_regx71x : DFF_X1 port map( D => Key(71), CK => clk, Q => 
                           reg_key_71_port, QN => n_1232);
   reg_key_regx66x : DFF_X1 port map( D => Key(66), CK => clk, Q => 
                           reg_key_66_port, QN => n_1233);
   reg_key_regx65x : DFF_X1 port map( D => Key(65), CK => clk, Q => 
                           reg_key_65_port, QN => n_1234);
   reg_key_regx60x : DFF_X1 port map( D => Key(60), CK => clk, Q => 
                           reg_key_60_port, QN => n_1235);
   reg_key_regx59x : DFF_X1 port map( D => Key(59), CK => clk, Q => 
                           reg_key_59_port, QN => n_1236);
   reg_key_regx58x : DFF_X1 port map( D => Key(58), CK => clk, Q => 
                           reg_key_58_port, QN => n_1237);
   reg_key_regx51x : DFF_X1 port map( D => Key(51), CK => clk, Q => 
                           reg_key_51_port, QN => n_1238);
   reg_key_regx48x : DFF_X1 port map( D => Key(48), CK => clk, Q => 
                           reg_key_48_port, QN => n_1239);
   reg_key_regx45x : DFF_X1 port map( D => Key(45), CK => clk, Q => 
                           reg_key_45_port, QN => n_1240);
   reg_key_regx44x : DFF_X1 port map( D => Key(44), CK => clk, Q => 
                           reg_key_44_port, QN => n_1241);
   reg_key_regx38x : DFF_X1 port map( D => Key(38), CK => clk, Q => 
                           reg_key_38_port, QN => n_1242);
   reg_key_regx36x : DFF_X1 port map( D => Key(36), CK => clk, Q => 
                           reg_key_36_port, QN => n_1243);
   reg_key_regx30x : DFF_X1 port map( D => Key(30), CK => clk, Q => 
                           reg_key_30_port, QN => n_1244);
   reg_key_regx28x : DFF_X1 port map( D => Key(28), CK => clk, Q => 
                           reg_key_28_port, QN => n_1245);
   reg_key_regx25x : DFF_X1 port map( D => Key(25), CK => clk, Q => 
                           reg_key_25_port, QN => n_1246);
   reg_key_regx24x : DFF_X1 port map( D => Key(24), CK => clk, Q => 
                           reg_key_24_port, QN => n_1247);
   reg_key_regx21x : DFF_X1 port map( D => Key(21), CK => clk, Q => 
                           reg_key_21_port, QN => n_1248);
   reg_key_regx20x : DFF_X1 port map( D => Key(20), CK => clk, Q => 
                           reg_key_20_port, QN => n_1249);
   reg_key_regx18x : DFF_X1 port map( D => Key(18), CK => clk, Q => 
                           reg_key_18_port, QN => n_1250);
   reg_key_regx10x : DFF_X1 port map( D => Key(10), CK => clk, Q => 
                           reg_key_10_port, QN => n_1251);
   reg_key_regx9x : DFF_X1 port map( D => Key(9), CK => clk, Q => 
                           reg_key_9_port, QN => n_1252);
   reg_key_regx6x : DFF_X1 port map( D => Key(6), CK => clk, Q => 
                           reg_key_6_port, QN => n_1253);
   reg_key_regx5x : DFF_X1 port map( D => Key(5), CK => clk, Q => 
                           reg_key_5_port, QN => n_1254);
   reg_key_regx4x : DFF_X1 port map( D => Key(4), CK => clk, Q => 
                           reg_key_4_port, QN => n_1255);
   reg_key_regx3x : DFF_X1 port map( D => Key(3), CK => clk, Q => 
                           reg_key_3_port, QN => n_1256);
   Ciphertext_regx190x : DFF_X1 port map( D => reg_out_190_port, CK => clk, Q 
                           => Ciphertext(190), QN => n_1257);
   Ciphertext_regx188x : DFF_X1 port map( D => reg_out_188_port, CK => clk, Q 
                           => Ciphertext(188), QN => n_1258);
   Ciphertext_regx187x : DFF_X1 port map( D => reg_out_187_port, CK => clk, Q 
                           => Ciphertext(187), QN => n_1259);
   Ciphertext_regx185x : DFF_X1 port map( D => reg_out_185_port, CK => clk, Q 
                           => Ciphertext(185), QN => n_1260);
   Ciphertext_regx183x : DFF_X1 port map( D => reg_out_183_port, CK => clk, Q 
                           => Ciphertext(183), QN => n_1261);
   Ciphertext_regx177x : DFF_X1 port map( D => reg_out_177_port, CK => clk, Q 
                           => Ciphertext(177), QN => n_1262);
   Ciphertext_regx171x : DFF_X1 port map( D => reg_out_171_port, CK => clk, Q 
                           => Ciphertext(171), QN => n_1263);
   Ciphertext_regx170x : DFF_X1 port map( D => reg_out_170_port, CK => clk, Q 
                           => Ciphertext(170), QN => n_1264);
   Ciphertext_regx169x : DFF_X1 port map( D => reg_out_169_port, CK => clk, Q 
                           => Ciphertext(169), QN => n_1265);
   Ciphertext_regx168x : DFF_X1 port map( D => reg_out_168_port, CK => clk, Q 
                           => Ciphertext(168), QN => n_1266);
   Ciphertext_regx167x : DFF_X1 port map( D => reg_out_167_port, CK => clk, Q 
                           => Ciphertext(167), QN => n_1267);
   Ciphertext_regx165x : DFF_X1 port map( D => reg_out_165_port, CK => clk, Q 
                           => Ciphertext(165), QN => n_1268);
   Ciphertext_regx164x : DFF_X1 port map( D => reg_out_164_port, CK => clk, Q 
                           => Ciphertext(164), QN => n_1269);
   Ciphertext_regx163x : DFF_X1 port map( D => reg_out_163_port, CK => clk, Q 
                           => Ciphertext(163), QN => n_1270);
   Ciphertext_regx160x : DFF_X1 port map( D => reg_out_160_port, CK => clk, Q 
                           => Ciphertext(160), QN => n_1271);
   Ciphertext_regx159x : DFF_X1 port map( D => reg_out_159_port, CK => clk, Q 
                           => Ciphertext(159), QN => n_1272);
   Ciphertext_regx158x : DFF_X1 port map( D => reg_out_158_port, CK => clk, Q 
                           => Ciphertext(158), QN => n_1273);
   Ciphertext_regx155x : DFF_X1 port map( D => reg_out_155_port, CK => clk, Q 
                           => Ciphertext(155), QN => n_1274);
   Ciphertext_regx152x : DFF_X1 port map( D => reg_out_152_port, CK => clk, Q 
                           => Ciphertext(152), QN => n_1275);
   Ciphertext_regx149x : DFF_X1 port map( D => reg_out_149_port, CK => clk, Q 
                           => Ciphertext(149), QN => n_1276);
   Ciphertext_regx148x : DFF_X1 port map( D => reg_out_148_port, CK => clk, Q 
                           => Ciphertext(148), QN => n_1277);
   Ciphertext_regx147x : DFF_X1 port map( D => reg_out_147_port, CK => clk, Q 
                           => Ciphertext(147), QN => n_1278);
   Ciphertext_regx145x : DFF_X1 port map( D => reg_out_145_port, CK => clk, Q 
                           => Ciphertext(145), QN => n_1279);
   Ciphertext_regx143x : DFF_X1 port map( D => reg_out_143_port, CK => clk, Q 
                           => Ciphertext(143), QN => n_1280);
   Ciphertext_regx142x : DFF_X1 port map( D => reg_out_142_port, CK => clk, Q 
                           => Ciphertext(142), QN => n_1281);
   Ciphertext_regx141x : DFF_X1 port map( D => reg_out_141_port, CK => clk, Q 
                           => Ciphertext(141), QN => n_1282);
   Ciphertext_regx140x : DFF_X1 port map( D => reg_out_140_port, CK => clk, Q 
                           => Ciphertext(140), QN => n_1283);
   Ciphertext_regx139x : DFF_X1 port map( D => reg_out_139_port, CK => clk, Q 
                           => Ciphertext(139), QN => n_1284);
   Ciphertext_regx138x : DFF_X1 port map( D => reg_out_138_port, CK => clk, Q 
                           => Ciphertext(138), QN => n_1285);
   Ciphertext_regx137x : DFF_X1 port map( D => reg_out_137_port, CK => clk, Q 
                           => Ciphertext(137), QN => n_1286);
   Ciphertext_regx136x : DFF_X1 port map( D => reg_out_136_port, CK => clk, Q 
                           => Ciphertext(136), QN => n_1287);
   Ciphertext_regx135x : DFF_X1 port map( D => reg_out_135_port, CK => clk, Q 
                           => Ciphertext(135), QN => n_1288);
   Ciphertext_regx131x : DFF_X1 port map( D => reg_out_131_port, CK => clk, Q 
                           => Ciphertext(131), QN => n_1289);
   Ciphertext_regx130x : DFF_X1 port map( D => reg_out_130_port, CK => clk, Q 
                           => Ciphertext(130), QN => n_1290);
   Ciphertext_regx129x : DFF_X1 port map( D => reg_out_129_port, CK => clk, Q 
                           => Ciphertext(129), QN => n_1291);
   Ciphertext_regx128x : DFF_X1 port map( D => reg_out_128_port, CK => clk, Q 
                           => Ciphertext(128), QN => n_1292);
   Ciphertext_regx126x : DFF_X1 port map( D => reg_out_126_port, CK => clk, Q 
                           => Ciphertext(126), QN => n_1293);
   Ciphertext_regx125x : DFF_X1 port map( D => reg_out_125_port, CK => clk, Q 
                           => Ciphertext(125), QN => n_1294);
   Ciphertext_regx122x : DFF_X1 port map( D => reg_out_122_port, CK => clk, Q 
                           => Ciphertext(122), QN => n_1295);
   Ciphertext_regx120x : DFF_X1 port map( D => reg_out_120_port, CK => clk, Q 
                           => Ciphertext(120), QN => n_1296);
   Ciphertext_regx118x : DFF_X1 port map( D => reg_out_118_port, CK => clk, Q 
                           => Ciphertext(118), QN => n_1297);
   Ciphertext_regx116x : DFF_X1 port map( D => reg_out_116_port, CK => clk, Q 
                           => Ciphertext(116), QN => n_1298);
   Ciphertext_regx112x : DFF_X1 port map( D => reg_out_112_port, CK => clk, Q 
                           => Ciphertext(112), QN => n_1299);
   Ciphertext_regx108x : DFF_X1 port map( D => reg_out_108_port, CK => clk, Q 
                           => Ciphertext(108), QN => n_1300);
   Ciphertext_regx106x : DFF_X1 port map( D => reg_out_106_port, CK => clk, Q 
                           => Ciphertext(106), QN => n_1301);
   Ciphertext_regx101x : DFF_X1 port map( D => reg_out_101_port, CK => clk, Q 
                           => Ciphertext(101), QN => n_1302);
   Ciphertext_regx98x : DFF_X1 port map( D => reg_out_98_port, CK => clk, Q => 
                           Ciphertext(98), QN => n_1303);
   Ciphertext_regx92x : DFF_X1 port map( D => reg_out_92_port, CK => clk, Q => 
                           Ciphertext(92), QN => n_1304);
   Ciphertext_regx91x : DFF_X1 port map( D => reg_out_91_port, CK => clk, Q => 
                           Ciphertext(91), QN => n_1305);
   Ciphertext_regx89x : DFF_X1 port map( D => reg_out_89_port, CK => clk, Q => 
                           Ciphertext(89), QN => n_1306);
   Ciphertext_regx88x : DFF_X1 port map( D => reg_out_88_port, CK => clk, Q => 
                           Ciphertext(88), QN => n_1307);
   Ciphertext_regx87x : DFF_X1 port map( D => reg_out_87_port, CK => clk, Q => 
                           Ciphertext(87), QN => n_1308);
   Ciphertext_regx86x : DFF_X1 port map( D => reg_out_86_port, CK => clk, Q => 
                           Ciphertext(86), QN => n_1309);
   Ciphertext_regx84x : DFF_X1 port map( D => reg_out_84_port, CK => clk, Q => 
                           Ciphertext(84), QN => n_1310);
   Ciphertext_regx83x : DFF_X1 port map( D => reg_out_83_port, CK => clk, Q => 
                           Ciphertext(83), QN => n_1311);
   Ciphertext_regx82x : DFF_X1 port map( D => reg_out_82_port, CK => clk, Q => 
                           Ciphertext(82), QN => n_1312);
   Ciphertext_regx77x : DFF_X1 port map( D => reg_out_77_port, CK => clk, Q => 
                           Ciphertext(77), QN => n_1313);
   Ciphertext_regx74x : DFF_X1 port map( D => reg_out_74_port, CK => clk, Q => 
                           Ciphertext(74), QN => n_1314);
   Ciphertext_regx72x : DFF_X1 port map( D => reg_out_72_port, CK => clk, Q => 
                           Ciphertext(72), QN => n_1315);
   Ciphertext_regx64x : DFF_X1 port map( D => reg_out_64_port, CK => clk, Q => 
                           Ciphertext(64), QN => n_1316);
   Ciphertext_regx62x : DFF_X1 port map( D => reg_out_62_port, CK => clk, Q => 
                           Ciphertext(62), QN => n_1317);
   Ciphertext_regx57x : DFF_X1 port map( D => reg_out_57_port, CK => clk, Q => 
                           Ciphertext(57), QN => n_1318);
   Ciphertext_regx56x : DFF_X1 port map( D => reg_out_56_port, CK => clk, Q => 
                           Ciphertext(56), QN => n_1319);
   Ciphertext_regx54x : DFF_X1 port map( D => reg_out_54_port, CK => clk, Q => 
                           Ciphertext(54), QN => n_1320);
   Ciphertext_regx49x : DFF_X1 port map( D => reg_out_49_port, CK => clk, Q => 
                           Ciphertext(49), QN => n_1321);
   Ciphertext_regx46x : DFF_X1 port map( D => reg_out_46_port, CK => clk, Q => 
                           Ciphertext(46), QN => n_1322);
   Ciphertext_regx41x : DFF_X1 port map( D => reg_out_41_port, CK => clk, Q => 
                           Ciphertext(41), QN => n_1323);
   Ciphertext_regx37x : DFF_X1 port map( D => reg_out_37_port, CK => clk, Q => 
                           Ciphertext(37), QN => n_1324);
   Ciphertext_regx35x : DFF_X1 port map( D => reg_out_35_port, CK => clk, Q => 
                           Ciphertext(35), QN => n_1325);
   Ciphertext_regx34x : DFF_X1 port map( D => reg_out_34_port, CK => clk, Q => 
                           Ciphertext(34), QN => n_1326);
   Ciphertext_regx33x : DFF_X1 port map( D => reg_out_33_port, CK => clk, Q => 
                           Ciphertext(33), QN => n_1327);
   Ciphertext_regx32x : DFF_X1 port map( D => reg_out_32_port, CK => clk, Q => 
                           Ciphertext(32), QN => n_1328);
   Ciphertext_regx31x : DFF_X1 port map( D => reg_out_31_port, CK => clk, Q => 
                           Ciphertext(31), QN => n_1329);
   Ciphertext_regx30x : DFF_X1 port map( D => reg_out_30_port, CK => clk, Q => 
                           Ciphertext(30), QN => n_1330);
   Ciphertext_regx29x : DFF_X1 port map( D => reg_out_29_port, CK => clk, Q => 
                           Ciphertext(29), QN => n_1331);
   Ciphertext_regx28x : DFF_X1 port map( D => reg_out_28_port, CK => clk, Q => 
                           Ciphertext(28), QN => n_1332);
   Ciphertext_regx26x : DFF_X1 port map( D => reg_out_26_port, CK => clk, Q => 
                           Ciphertext(26), QN => n_1333);
   Ciphertext_regx23x : DFF_X1 port map( D => reg_out_23_port, CK => clk, Q => 
                           Ciphertext(23), QN => n_1334);
   Ciphertext_regx18x : DFF_X1 port map( D => reg_out_18_port, CK => clk, Q => 
                           Ciphertext(18), QN => n_1335);
   Ciphertext_regx17x : DFF_X1 port map( D => reg_out_17_port, CK => clk, Q => 
                           Ciphertext(17), QN => n_1336);
   Ciphertext_regx15x : DFF_X1 port map( D => reg_out_15_port, CK => clk, Q => 
                           Ciphertext(15), QN => n_1337);
   Ciphertext_regx14x : DFF_X1 port map( D => reg_out_14_port, CK => clk, Q => 
                           Ciphertext(14), QN => n_1338);
   Ciphertext_regx13x : DFF_X1 port map( D => reg_out_13_port, CK => clk, Q => 
                           Ciphertext(13), QN => n_1339);
   Ciphertext_regx11x : DFF_X1 port map( D => reg_out_11_port, CK => clk, Q => 
                           Ciphertext(11), QN => n_1340);
   Ciphertext_regx10x : DFF_X1 port map( D => reg_out_10_port, CK => clk, Q => 
                           Ciphertext(10), QN => n_1341);
   Ciphertext_regx8x : DFF_X1 port map( D => reg_out_8_port, CK => clk, Q => 
                           Ciphertext(8), QN => n_1342);
   Ciphertext_regx6x : DFF_X1 port map( D => reg_out_6_port, CK => clk, Q => 
                           Ciphertext(6), QN => n_1343);
   Ciphertext_regx5x : DFF_X1 port map( D => reg_out_5_port, CK => clk, Q => 
                           Ciphertext(5), QN => n_1344);
   Ciphertext_regx4x : DFF_X1 port map( D => reg_out_4_port, CK => clk, Q => 
                           Ciphertext(4), QN => n_1345);
   Ciphertext_regx2x : DFF_X1 port map( D => reg_out_2_port, CK => clk, Q => 
                           Ciphertext(2), QN => n_1346);
   Ciphertext_regx0x : DFF_X1 port map( D => reg_out_0_port, CK => clk, Q => 
                           Ciphertext(0), QN => n_1347);
   reg_key_regx14x : DFF_X1 port map( D => Key(14), CK => clk, Q => 
                           reg_key_14_port, QN => n_1348);
   reg_key_regx122x : DFF_X1 port map( D => Key(122), CK => clk, Q => 
                           reg_key_122_port, QN => n_1349);
   reg_key_regx86x : DFF_X1 port map( D => Key(86), CK => clk, Q => 
                           reg_key_86_port, QN => n_1350);
   Ciphertext_regx100x : DFF_X1 port map( D => reg_out_100_port, CK => clk, Q 
                           => Ciphertext(100), QN => n_1351);
   reg_key_regx111x : DFF_X1 port map( D => Key(111), CK => clk, Q => 
                           reg_key_111_port, QN => n_1352);
   reg_key_regx54x : DFF_X1 port map( D => Key(54), CK => clk, Q => 
                           reg_key_54_port, QN => n_1353);
   reg_key_regx61x : DFF_X1 port map( D => Key(61), CK => clk, Q => 
                           reg_key_61_port, QN => n_1354);
   reg_key_regx116x : DFF_X1 port map( D => Key(116), CK => clk, Q => 
                           reg_key_116_port, QN => n_1355);
   reg_key_regx158x : DFF_X1 port map( D => Key(158), CK => clk, Q => 
                           reg_key_158_port, QN => n_1356);
   reg_key_regx15x : DFF_X1 port map( D => Key(15), CK => clk, Q => 
                           reg_key_15_port, QN => n_1357);
   reg_key_regx185x : DFF_X1 port map( D => Key(185), CK => clk, Q => 
                           reg_key_185_port, QN => n_1358);
   reg_key_regx13x : DFF_X1 port map( D => Key(13), CK => clk, Q => 
                           reg_key_13_port, QN => n_1359);
   reg_key_regx8x : DFF_X1 port map( D => Key(8), CK => clk, Q => 
                           reg_key_8_port, QN => n_1360);
   reg_key_regx2x : DFF_X1 port map( D => Key(2), CK => clk, Q => 
                           reg_key_2_port, QN => n_1361);
   reg_key_regx29x : DFF_X1 port map( D => Key(29), CK => clk, Q => 
                           reg_key_29_port, QN => n_1362);
   reg_key_regx74x : DFF_X1 port map( D => Key(74), CK => clk, Q => 
                           reg_key_74_port, QN => n_1363);
   reg_key_regx98x : DFF_X1 port map( D => Key(98), CK => clk, Q => 
                           reg_key_98_port, QN => n_1364);
   reg_key_regx83x : DFF_X1 port map( D => Key(83), CK => clk, Q => 
                           reg_key_83_port, QN => n_1365);
   reg_key_regx183x : DFF_X1 port map( D => Key(183), CK => clk, Q => 
                           reg_key_183_port, QN => n_1366);
   reg_key_regx107x : DFF_X1 port map( D => Key(107), CK => clk, Q => 
                           reg_key_107_port, QN => n_1367);
   reg_key_regx146x : DFF_X1 port map( D => Key(146), CK => clk, Q => 
                           reg_key_146_port, QN => n_1368);
   reg_key_regx56x : DFF_X1 port map( D => Key(56), CK => clk, Q => 
                           reg_key_56_port, QN => n_1369);
   reg_key_regx152x : DFF_X1 port map( D => Key(152), CK => clk, Q => 
                           reg_key_152_port, QN => n_1370);
   reg_key_regx63x : DFF_X1 port map( D => Key(63), CK => clk, Q => 
                           reg_key_63_port, QN => n_1371);
   reg_key_regx134x : DFF_X1 port map( D => Key(134), CK => clk, Q => 
                           reg_key_134_port, QN => n_1372);
   reg_key_regx106x : DFF_X1 port map( D => Key(106), CK => clk, Q => 
                           reg_key_106_port, QN => n_1373);
   reg_key_regx41x : DFF_X1 port map( D => Key(41), CK => clk, Q => 
                           reg_key_41_port, QN => n_1374);
   reg_key_regx16x : DFF_X1 port map( D => Key(16), CK => clk, Q => 
                           reg_key_16_port, QN => n_1375);
   reg_key_regx35x : DFF_X1 port map( D => Key(35), CK => clk, Q => 
                           reg_key_35_port, QN => n_1376);
   reg_key_regx102x : DFF_X1 port map( D => Key(102), CK => clk, Q => 
                           reg_key_102_port, QN => n_1377);
   reg_key_regx27x : DFF_X1 port map( D => Key(27), CK => clk, Q => 
                           reg_key_27_port, QN => n_1378);
   Ciphertext_regx124x : DFF_X1 port map( D => reg_out_124_port, CK => clk, Q 
                           => Ciphertext(124), QN => n_1379);
   reg_key_regx22x : DFF_X1 port map( D => Key(22), CK => clk, Q => 
                           reg_key_22_port, QN => n_1380);
   reg_key_regx163x : DFF_X1 port map( D => Key(163), CK => clk, Q => 
                           reg_key_163_port, QN => n_1381);
   reg_key_regx159x : DFF_X1 port map( D => Key(159), CK => clk, Q => 
                           reg_key_159_port, QN => n_1382);
   reg_key_regx155x : DFF_X1 port map( D => Key(155), CK => clk, Q => 
                           reg_key_155_port, QN => n_1383);
   reg_key_regx147x : DFF_X1 port map( D => Key(147), CK => clk, Q => 
                           reg_key_147_port, QN => n_1384);
   reg_key_regx49x : DFF_X1 port map( D => Key(49), CK => clk, Q => 
                           reg_key_49_port, QN => n_1385);
   reg_key_regx92x : DFF_X1 port map( D => Key(92), CK => clk, Q => 
                           reg_key_92_port, QN => n_1386);
   reg_key_regx186x : DFF_X1 port map( D => Key(186), CK => clk, Q => 
                           reg_key_186_port, QN => n_1387);
   reg_key_regx182x : DFF_X1 port map( D => Key(182), CK => clk, Q => 
                           reg_key_182_port, QN => n_1388);
   reg_key_regx84x : DFF_X1 port map( D => Key(84), CK => clk, Q => 
                           reg_key_84_port, QN => n_1389);
   reg_key_regx131x : DFF_X1 port map( D => Key(131), CK => clk, Q => 
                           reg_key_131_port, QN => n_1390);
   reg_key_regx170x : DFF_X1 port map( D => Key(170), CK => clk, Q => 
                           reg_key_170_port, QN => n_1391);
   reg_key_regx72x : DFF_X1 port map( D => Key(72), CK => clk, Q => 
                           reg_key_72_port, QN => n_1392);
   reg_key_regx68x : DFF_X1 port map( D => Key(68), CK => clk, Q => 
                           reg_key_68_port, QN => n_1393);
   reg_key_regx17x : DFF_X1 port map( D => Key(17), CK => clk, Q => 
                           reg_key_17_port, QN => n_1394);
   reg_key_regx154x : DFF_X1 port map( D => Key(154), CK => clk, Q => 
                           reg_key_154_port, QN => n_1395);
   reg_key_regx150x : DFF_X1 port map( D => Key(150), CK => clk, Q => 
                           reg_key_150_port, QN => n_1396);
   reg_key_regx99x : DFF_X1 port map( D => Key(99), CK => clk, Q => 
                           reg_key_99_port, QN => n_1397);
   reg_key_regx1x : DFF_X1 port map( D => Key(1), CK => clk, Q => 
                           reg_key_1_port, QN => n_1398);
   reg_key_regx138x : DFF_X1 port map( D => Key(138), CK => clk, Q => 
                           reg_key_138_port, QN => n_1399);
   reg_key_regx40x : DFF_X1 port map( D => Key(40), CK => clk, Q => 
                           reg_key_40_port, QN => n_1400);
   reg_key_regx87x : DFF_X1 port map( D => Key(87), CK => clk, Q => 
                           reg_key_87_port, QN => n_1401);
   reg_key_regx181x : DFF_X1 port map( D => Key(181), CK => clk, Q => 
                           reg_key_181_port, QN => n_1402);
   reg_key_regx130x : DFF_X1 port map( D => Key(130), CK => clk, Q => 
                           reg_key_130_port, QN => n_1403);
   reg_key_regx32x : DFF_X1 port map( D => Key(32), CK => clk, Q => 
                           reg_key_32_port, QN => n_1404);
   reg_key_regx79x : DFF_X1 port map( D => Key(79), CK => clk, Q => 
                           reg_key_79_port, QN => n_1405);
   reg_key_regx75x : DFF_X1 port map( D => Key(75), CK => clk, Q => 
                           reg_key_75_port, QN => n_1406);
   reg_key_regx114x : DFF_X1 port map( D => Key(114), CK => clk, Q => 
                           reg_key_114_port, QN => n_1407);
   reg_key_regx161x : DFF_X1 port map( D => Key(161), CK => clk, Q => 
                           reg_key_161_port, QN => n_1408);
   reg_key_regx157x : DFF_X1 port map( D => Key(157), CK => clk, Q => 
                           reg_key_157_port, QN => n_1409);
   reg_key_regx12x : DFF_X1 port map( D => Key(12), CK => clk, Q => 
                           reg_key_12_port, QN => n_1410);
   reg_key_regx153x : DFF_X1 port map( D => Key(153), CK => clk, Q => 
                           reg_key_153_port, QN => n_1411);
   reg_key_regx55x : DFF_X1 port map( D => Key(55), CK => clk, Q => 
                           reg_key_55_port, QN => n_1412);
   reg_key_regx145x : DFF_X1 port map( D => Key(145), CK => clk, Q => 
                           reg_key_145_port, QN => n_1413);
   reg_key_regx94x : DFF_X1 port map( D => Key(94), CK => clk, Q => 
                           reg_key_94_port, QN => n_1414);
   reg_key_regx141x : DFF_X1 port map( D => Key(141), CK => clk, Q => 
                           reg_key_141_port, QN => n_1415);
   reg_key_regx43x : DFF_X1 port map( D => Key(43), CK => clk, Q => 
                           reg_key_43_port, QN => n_1416);
   reg_key_regx39x : DFF_X1 port map( D => Key(39), CK => clk, Q => 
                           reg_key_39_port, QN => n_1417);
   reg_key_regx133x : DFF_X1 port map( D => Key(133), CK => clk, Q => 
                           reg_key_133_port, QN => n_1418);
   reg_key_regx176x : DFF_X1 port map( D => Key(176), CK => clk, Q => 
                           reg_key_176_port, QN => n_1419);
   reg_key_regx31x : DFF_X1 port map( D => Key(31), CK => clk, Q => 
                           reg_key_31_port, QN => n_1420);
   reg_key_regx78x : DFF_X1 port map( D => Key(78), CK => clk, Q => 
                           reg_key_78_port, QN => n_1421);
   reg_key_regx121x : DFF_X1 port map( D => Key(121), CK => clk, Q => 
                           reg_key_121_port, QN => n_1422);
   reg_key_regx23x : DFF_X1 port map( D => Key(23), CK => clk, Q => 
                           reg_key_23_port, QN => n_1423);
   reg_key_regx117x : DFF_X1 port map( D => Key(117), CK => clk, Q => 
                           reg_key_117_port, QN => n_1424);
   reg_key_regx19x : DFF_X1 port map( D => Key(19), CK => clk, Q => 
                           reg_key_19_port, QN => n_1425);
   reg_key_regx113x : DFF_X1 port map( D => Key(113), CK => clk, Q => 
                           reg_key_113_port, QN => n_1426);
   reg_key_regx11x : DFF_X1 port map( D => Key(11), CK => clk, Q => 
                           reg_key_11_port, QN => n_1427);
   reg_key_regx7x : DFF_X1 port map( D => Key(7), CK => clk, Q => 
                           reg_key_7_port, QN => n_1428);
   reg_key_regx50x : DFF_X1 port map( D => Key(50), CK => clk, Q => 
                           reg_key_50_port, QN => n_1429);
   reg_key_regx144x : DFF_X1 port map( D => Key(144), CK => clk, Q => 
                           reg_key_144_port, QN => n_1430);
   reg_key_regx42x : DFF_X1 port map( D => Key(42), CK => clk, Q => 
                           reg_key_42_port, QN => n_1431);
   reg_key_regx89x : DFF_X1 port map( D => Key(89), CK => clk, Q => 
                           reg_key_89_port, QN => n_1432);
   reg_key_regx85x : DFF_X1 port map( D => Key(85), CK => clk, Q => 
                           reg_key_85_port, QN => n_1433);
   reg_key_regx34x : DFF_X1 port map( D => Key(34), CK => clk, Q => 
                           reg_key_34_port, QN => n_1434);
   reg_key_regx128x : DFF_X1 port map( D => Key(128), CK => clk, Q => 
                           reg_key_128_port, QN => n_1435);
   reg_key_regx26x : DFF_X1 port map( D => Key(26), CK => clk, Q => 
                           reg_key_26_port, QN => n_1436);
   reg_key_regx90x : DFF_X1 port map( D => Key(90), CK => clk, Q => 
                           reg_key_90_port, QN => n_1437);
   reg_key_regx93x : DFF_X1 port map( D => Key(93), CK => clk, Q => 
                           reg_key_93_port, QN => n_1438);
   reg_key_regx52x : DFF_X1 port map( D => Key(52), CK => clk, Q => 
                           reg_key_52_port, QN => n_1439);
   reg_key_regx167x : DFF_X1 port map( D => Key(167), CK => clk, Q => 
                           reg_key_167_port, QN => n_1440);
   reg_key_regx53x : DFF_X1 port map( D => Key(53), CK => clk, Q => 
                           reg_key_53_port, QN => n_1441);
   reg_key_regx64x : DFF_X1 port map( D => Key(64), CK => clk, Q => 
                           reg_key_64_port, QN => n_1442);
   reg_key_regx91x : DFF_X1 port map( D => Key(91), CK => clk, Q => 
                           reg_key_91_port, QN => n_1443);
   reg_key_regx126x : DFF_X1 port map( D => Key(126), CK => clk, Q => 
                           reg_key_126_port, QN => n_1444);
   reg_key_regx175x : DFF_X1 port map( D => Key(175), CK => clk, Q => 
                           reg_key_175_port, QN => n_1445);
   reg_key_regx33x : DFF_X1 port map( D => Key(33), CK => clk, Q => 
                           reg_key_33_port, QN => n_1446);
   reg_key_regx112x : DFF_X1 port map( D => Key(112), CK => clk, Q => 
                           reg_key_112_port, QN => n_1447);
   reg_key_regx139x : DFF_X1 port map( D => Key(139), CK => clk, Q => 
                           reg_key_139_port, QN => n_1448);
   reg_key_regx127x : DFF_X1 port map( D => Key(127), CK => clk, Q => 
                           reg_key_127_port, QN => n_1449);
   reg_key_regx142x : DFF_X1 port map( D => Key(142), CK => clk, Q => 
                           reg_key_142_port, QN => n_1450);
   reg_key_regx110x : DFF_X1 port map( D => Key(110), CK => clk, Q => 
                           reg_key_110_port, QN => n_1451);
   reg_key_regx62x : DFF_X1 port map( D => Key(62), CK => clk, Q => 
                           reg_key_62_port, QN => n_1452);
   reg_key_regx164x : DFF_X1 port map( D => Key(164), CK => clk, Q => 
                           reg_key_164_port, QN => n_1453);
   reg_key_regx97x : DFF_X1 port map( D => Key(97), CK => clk, Q => 
                           reg_key_97_port, QN => n_1454);
   reg_key_regx168x : DFF_X1 port map( D => Key(168), CK => clk, Q => 
                           reg_key_168_port, QN => n_1455);
   reg_key_regx115x : DFF_X1 port map( D => Key(115), CK => clk, Q => 
                           reg_key_115_port, QN => n_1456);
   reg_key_regx162x : DFF_X1 port map( D => Key(162), CK => clk, Q => 
                           reg_key_162_port, QN => n_1457);
   reg_key_regx37x : DFF_X1 port map( D => Key(37), CK => clk, Q => 
                           reg_key_37_port, QN => n_1458);
   reg_key_regx129x : DFF_X1 port map( D => Key(129), CK => clk, Q => 
                           reg_key_129_port, QN => n_1459);
   reg_key_regx124x : DFF_X1 port map( D => Key(124), CK => clk, Q => 
                           reg_key_124_port, QN => n_1460);
   reg_key_regx69x : DFF_X1 port map( D => Key(69), CK => clk, Q => 
                           reg_key_69_port, QN => n_1461);
   reg_key_regx73x : DFF_X1 port map( D => Key(73), CK => clk, Q => 
                           reg_key_73_port, QN => n_1462);
   reg_key_regx46x : DFF_X1 port map( D => Key(46), CK => clk, Q => 
                           reg_key_46_port, QN => n_1463);
   reg_key_regx57x : DFF_X1 port map( D => Key(57), CK => clk, Q => 
                           reg_key_57_port, QN => n_1464);
   reg_key_regx180x : DFF_X1 port map( D => Key(180), CK => clk, Q => 
                           reg_key_180_port, QN => n_1465);
   reg_key_regx77x : DFF_X1 port map( D => Key(77), CK => clk, Q => 
                           reg_key_77_port, QN => n_1466);
   reg_key_regx47x : DFF_X1 port map( D => Key(47), CK => clk, Q => 
                           reg_key_47_port, QN => n_1467);
   reg_key_regx0x : DFF_X1 port map( D => Key(0), CK => clk, Q => 
                           reg_key_0_port, QN => n_1468);
   reg_key_regx67x : DFF_X1 port map( D => Key(67), CK => clk, Q => 
                           reg_key_67_port, QN => n_1469);
   reg_key_regx166x : DFF_X1 port map( D => Key(166), CK => clk, Q => 
                           reg_key_166_port, QN => n_1470);
   reg_key_regx136x : DFF_X1 port map( D => Key(136), CK => clk, Q => 
                           reg_key_136_port, QN => n_1471);
   reg_key_regx70x : DFF_X1 port map( D => Key(70), CK => clk, Q => 
                           reg_key_70_port, QN => n_1472);
   reg_key_regx148x : DFF_X1 port map( D => Key(148), CK => clk, Q => 
                           reg_key_148_port, QN => n_1473);
   reg_key_regx88x : DFF_X1 port map( D => Key(88), CK => clk, Q => 
                           reg_key_88_port, QN => n_1474);
   reg_key_regx174x : DFF_X1 port map( D => Key(174), CK => clk, Q => 
                           reg_key_174_port, QN => n_1475);
   Ciphertext_regx42x : DFFRS_X1 port map( D => reg_out_42_port, CK => clk, RN 
                           => n9, SN => n9, Q => Ciphertext(42), QN => n_1476);
   Ciphertext_regx21x : DFF_X1 port map( D => reg_out_21_port, CK => clk, Q => 
                           Ciphertext(21), QN => n_1477);
   Ciphertext_regx65x : DFF_X1 port map( D => reg_out_65_port, CK => clk, Q => 
                           Ciphertext(65), QN => n_1478);
   n9 <= '1';
   Ciphertext_regx105x : DFF_X1 port map( D => reg_out_105_port, CK => clk, Q 
                           => Ciphertext(105), QN => n_1479);
   Ciphertext_regx27x : DFF_X1 port map( D => reg_out_27_port, CK => clk, Q => 
                           Ciphertext(27), QN => n_1480);
   Ciphertext_regx133x : DFF_X1 port map( D => reg_out_133_port, CK => clk, Q 
                           => Ciphertext(133), QN => n_1481);
   Ciphertext_regx154x : DFF_X1 port map( D => reg_out_154_port, CK => clk, Q 
                           => Ciphertext(154), QN => n_1482);
   Ciphertext_regx103x : DFF_X1 port map( D => reg_out_103_port, CK => clk, Q 
                           => Ciphertext(103), QN => n_1483);
   Ciphertext_regx73x : DFF_X1 port map( D => reg_out_73_port, CK => clk, Q => 
                           Ciphertext(73), QN => n_1484);
   Ciphertext_regx90x : DFF_X1 port map( D => reg_out_90_port, CK => clk, Q => 
                           Ciphertext(90), QN => n_1485);
   Ciphertext_regx39x : DFF_X1 port map( D => reg_out_39_port, CK => clk, Q => 
                           Ciphertext(39), QN => n_1486);
   Ciphertext_regx132x : DFF_X1 port map( D => reg_out_132_port, CK => clk, Q 
                           => Ciphertext(132), QN => n_1487);
   Ciphertext_regx79x : DFF_X1 port map( D => reg_out_79_port, CK => clk, Q => 
                           Ciphertext(79), QN => n_1488);
   Ciphertext_regx3x : DFF_X1 port map( D => reg_out_3_port, CK => clk, Q => 
                           Ciphertext(3), QN => n_1489);
   Ciphertext_regx50x : DFF_X1 port map( D => reg_out_50_port, CK => clk, Q => 
                           Ciphertext(50), QN => n_1490);
   Ciphertext_regx24x : DFF_X1 port map( D => reg_out_24_port, CK => clk, Q => 
                           Ciphertext(24), QN => n_1491);
   Ciphertext_regx80x : DFF_X1 port map( D => reg_out_80_port, CK => clk, Q => 
                           Ciphertext(80), QN => n_1492);
   Ciphertext_regx157x : DFF_X1 port map( D => reg_out_157_port, CK => clk, Q 
                           => Ciphertext(157), QN => n_1493);
   Ciphertext_regx114x : DFF_X1 port map( D => reg_out_114_port, CK => clk, Q 
                           => Ciphertext(114), QN => n_1494);
   Ciphertext_regx94x : DFF_X1 port map( D => reg_out_94_port, CK => clk, Q => 
                           Ciphertext(94), QN => n_1495);
   Ciphertext_regx38x : DFF_X1 port map( D => reg_out_38_port, CK => clk, Q => 
                           Ciphertext(38), QN => n_1496);
   Ciphertext_regx68x : DFF_X1 port map( D => reg_out_68_port, CK => clk, Q => 
                           Ciphertext(68), QN => n_1497);
   Ciphertext_regx70x : DFF_X1 port map( D => reg_out_70_port, CK => clk, Q => 
                           Ciphertext(70), QN => n_1498);
   Ciphertext_regx45x : DFF_X1 port map( D => reg_out_45_port, CK => clk, Q => 
                           Ciphertext(45), QN => n_1499);
   Ciphertext_regx7x : DFF_X1 port map( D => reg_out_7_port, CK => clk, Q => 
                           Ciphertext(7), QN => n_1500);
   Ciphertext_regx191x : DFF_X1 port map( D => reg_out_191_port, CK => clk, Q 
                           => Ciphertext(191), QN => n_1501);
   Ciphertext_regx180x : DFF_X1 port map( D => reg_out_180_port, CK => clk, Q 
                           => Ciphertext(180), QN => n_1502);
   reg_key_regx172x : DFF_X2 port map( D => Key(172), CK => clk, Q => 
                           reg_key_172_port, QN => n_1503);
   Ciphertext_regx176x : DFF_X2 port map( D => reg_out_176_port, CK => clk, Q 
                           => Ciphertext(176), QN => n_1504);
   Ciphertext_regx172x : DFF_X1 port map( D => reg_out_172_port, CK => clk, Q 
                           => Ciphertext(172), QN => n_1505);
   SPEEDY_instance : SPEEDY_Rounds6_0 port map( Plaintext(191) => 
                           reg_in_191_port, Plaintext(190) => reg_in_190_port, 
                           Plaintext(189) => reg_in_189_port, Plaintext(188) =>
                           reg_in_188_port, Plaintext(187) => reg_in_187_port, 
                           Plaintext(186) => reg_in_186_port, Plaintext(185) =>
                           reg_in_185_port, Plaintext(184) => reg_in_184_port, 
                           Plaintext(183) => reg_in_183_port, Plaintext(182) =>
                           reg_in_182_port, Plaintext(181) => reg_in_181_port, 
                           Plaintext(180) => reg_in_180_port, Plaintext(179) =>
                           reg_in_179_port, Plaintext(178) => reg_in_178_port, 
                           Plaintext(177) => reg_in_177_port, Plaintext(176) =>
                           reg_in_176_port, Plaintext(175) => reg_in_175_port, 
                           Plaintext(174) => reg_in_174_port, Plaintext(173) =>
                           reg_in_173_port, Plaintext(172) => reg_in_172_port, 
                           Plaintext(171) => reg_in_171_port, Plaintext(170) =>
                           reg_in_170_port, Plaintext(169) => reg_in_169_port, 
                           Plaintext(168) => reg_in_168_port, Plaintext(167) =>
                           reg_in_167_port, Plaintext(166) => reg_in_166_port, 
                           Plaintext(165) => reg_in_165_port, Plaintext(164) =>
                           reg_in_164_port, Plaintext(163) => reg_in_163_port, 
                           Plaintext(162) => reg_in_162_port, Plaintext(161) =>
                           reg_in_161_port, Plaintext(160) => reg_in_160_port, 
                           Plaintext(159) => reg_in_159_port, Plaintext(158) =>
                           reg_in_158_port, Plaintext(157) => reg_in_157_port, 
                           Plaintext(156) => reg_in_156_port, Plaintext(155) =>
                           reg_in_155_port, Plaintext(154) => reg_in_154_port, 
                           Plaintext(153) => reg_in_153_port, Plaintext(152) =>
                           reg_in_152_port, Plaintext(151) => reg_in_151_port, 
                           Plaintext(150) => reg_in_150_port, Plaintext(149) =>
                           reg_in_149_port, Plaintext(148) => reg_in_148_port, 
                           Plaintext(147) => reg_in_147_port, Plaintext(146) =>
                           reg_in_146_port, Plaintext(145) => reg_in_145_port, 
                           Plaintext(144) => reg_in_144_port, Plaintext(143) =>
                           reg_in_143_port, Plaintext(142) => reg_in_142_port, 
                           Plaintext(141) => reg_in_141_port, Plaintext(140) =>
                           reg_in_140_port, Plaintext(139) => reg_in_139_port, 
                           Plaintext(138) => reg_in_138_port, Plaintext(137) =>
                           reg_in_137_port, Plaintext(136) => reg_in_136_port, 
                           Plaintext(135) => reg_in_135_port, Plaintext(134) =>
                           reg_in_134_port, Plaintext(133) => reg_in_133_port, 
                           Plaintext(132) => reg_in_132_port, Plaintext(131) =>
                           reg_in_131_port, Plaintext(130) => reg_in_130_port, 
                           Plaintext(129) => reg_in_129_port, Plaintext(128) =>
                           reg_in_128_port, Plaintext(127) => reg_in_127_port, 
                           Plaintext(126) => reg_in_126_port, Plaintext(125) =>
                           reg_in_125_port, Plaintext(124) => reg_in_124_port, 
                           Plaintext(123) => reg_in_123_port, Plaintext(122) =>
                           reg_in_122_port, Plaintext(121) => reg_in_121_port, 
                           Plaintext(120) => reg_in_120_port, Plaintext(119) =>
                           reg_in_119_port, Plaintext(118) => reg_in_118_port, 
                           Plaintext(117) => reg_in_117_port, Plaintext(116) =>
                           reg_in_116_port, Plaintext(115) => reg_in_115_port, 
                           Plaintext(114) => reg_in_114_port, Plaintext(113) =>
                           reg_in_113_port, Plaintext(112) => reg_in_112_port, 
                           Plaintext(111) => reg_in_111_port, Plaintext(110) =>
                           reg_in_110_port, Plaintext(109) => reg_in_109_port, 
                           Plaintext(108) => reg_in_108_port, Plaintext(107) =>
                           reg_in_107_port, Plaintext(106) => reg_in_106_port, 
                           Plaintext(105) => reg_in_105_port, Plaintext(104) =>
                           reg_in_104_port, Plaintext(103) => reg_in_103_port, 
                           Plaintext(102) => reg_in_102_port, Plaintext(101) =>
                           reg_in_101_port, Plaintext(100) => reg_in_100_port, 
                           Plaintext(99) => reg_in_99_port, Plaintext(98) => 
                           reg_in_98_port, Plaintext(97) => reg_in_97_port, 
                           Plaintext(96) => reg_in_96_port, Plaintext(95) => 
                           reg_in_95_port, Plaintext(94) => reg_in_94_port, 
                           Plaintext(93) => reg_in_93_port, Plaintext(92) => 
                           reg_in_92_port, Plaintext(91) => reg_in_91_port, 
                           Plaintext(90) => reg_in_90_port, Plaintext(89) => 
                           reg_in_89_port, Plaintext(88) => reg_in_88_port, 
                           Plaintext(87) => reg_in_87_port, Plaintext(86) => 
                           reg_in_86_port, Plaintext(85) => reg_in_85_port, 
                           Plaintext(84) => reg_in_84_port, Plaintext(83) => 
                           reg_in_83_port, Plaintext(82) => reg_in_82_port, 
                           Plaintext(81) => reg_in_81_port, Plaintext(80) => 
                           reg_in_80_port, Plaintext(79) => reg_in_79_port, 
                           Plaintext(78) => reg_in_78_port, Plaintext(77) => 
                           reg_in_77_port, Plaintext(76) => reg_in_76_port, 
                           Plaintext(75) => reg_in_75_port, Plaintext(74) => 
                           reg_in_74_port, Plaintext(73) => reg_in_73_port, 
                           Plaintext(72) => reg_in_72_port, Plaintext(71) => 
                           reg_in_71_port, Plaintext(70) => reg_in_70_port, 
                           Plaintext(69) => reg_in_69_port, Plaintext(68) => 
                           reg_in_68_port, Plaintext(67) => reg_in_67_port, 
                           Plaintext(66) => reg_in_66_port, Plaintext(65) => 
                           reg_in_65_port, Plaintext(64) => reg_in_64_port, 
                           Plaintext(63) => reg_in_63_port, Plaintext(62) => 
                           reg_in_62_port, Plaintext(61) => reg_in_61_port, 
                           Plaintext(60) => reg_in_60_port, Plaintext(59) => 
                           reg_in_59_port, Plaintext(58) => reg_in_58_port, 
                           Plaintext(57) => reg_in_57_port, Plaintext(56) => 
                           reg_in_56_port, Plaintext(55) => reg_in_55_port, 
                           Plaintext(54) => reg_in_54_port, Plaintext(53) => 
                           reg_in_53_port, Plaintext(52) => reg_in_52_port, 
                           Plaintext(51) => reg_in_51_port, Plaintext(50) => 
                           reg_in_50_port, Plaintext(49) => reg_in_49_port, 
                           Plaintext(48) => reg_in_48_port, Plaintext(47) => 
                           reg_in_47_port, Plaintext(46) => reg_in_46_port, 
                           Plaintext(45) => reg_in_45_port, Plaintext(44) => 
                           reg_in_44_port, Plaintext(43) => reg_in_43_port, 
                           Plaintext(42) => reg_in_42_port, Plaintext(41) => 
                           reg_in_41_port, Plaintext(40) => reg_in_40_port, 
                           Plaintext(39) => reg_in_39_port, Plaintext(38) => 
                           reg_in_38_port, Plaintext(37) => reg_in_37_port, 
                           Plaintext(36) => reg_in_36_port, Plaintext(35) => 
                           reg_in_35_port, Plaintext(34) => reg_in_34_port, 
                           Plaintext(33) => reg_in_33_port, Plaintext(32) => 
                           reg_in_32_port, Plaintext(31) => reg_in_31_port, 
                           Plaintext(30) => reg_in_30_port, Plaintext(29) => 
                           reg_in_29_port, Plaintext(28) => reg_in_28_port, 
                           Plaintext(27) => reg_in_27_port, Plaintext(26) => 
                           reg_in_26_port, Plaintext(25) => reg_in_25_port, 
                           Plaintext(24) => reg_in_24_port, Plaintext(23) => 
                           reg_in_23_port, Plaintext(22) => reg_in_22_port, 
                           Plaintext(21) => reg_in_21_port, Plaintext(20) => 
                           reg_in_20_port, Plaintext(19) => reg_in_19_port, 
                           Plaintext(18) => reg_in_18_port, Plaintext(17) => 
                           reg_in_17_port, Plaintext(16) => reg_in_16_port, 
                           Plaintext(15) => reg_in_15_port, Plaintext(14) => 
                           reg_in_14_port, Plaintext(13) => reg_in_13_port, 
                           Plaintext(12) => reg_in_12_port, Plaintext(11) => 
                           reg_in_11_port, Plaintext(10) => reg_in_10_port, 
                           Plaintext(9) => reg_in_9_port, Plaintext(8) => 
                           reg_in_8_port, Plaintext(7) => reg_in_7_port, 
                           Plaintext(6) => reg_in_6_port, Plaintext(5) => 
                           reg_in_5_port, Plaintext(4) => reg_in_4_port, 
                           Plaintext(3) => reg_in_3_port, Plaintext(2) => 
                           reg_in_2_port, Plaintext(1) => reg_in_1_port, 
                           Plaintext(0) => reg_in_0_port, Key(191) => 
                           reg_key_191_port, Key(190) => reg_key_190_port, 
                           Key(189) => reg_key_189_port, Key(188) => 
                           reg_key_188_port, Key(187) => reg_key_187_port, 
                           Key(186) => reg_key_186_port, Key(185) => 
                           reg_key_185_port, Key(184) => reg_key_184_port, 
                           Key(183) => reg_key_183_port, Key(182) => 
                           reg_key_182_port, Key(181) => reg_key_181_port, 
                           Key(180) => reg_key_180_port, Key(179) => 
                           reg_key_179_port, Key(178) => reg_key_178_port, 
                           Key(177) => reg_key_177_port, Key(176) => 
                           reg_key_176_port, Key(175) => reg_key_175_port, 
                           Key(174) => reg_key_174_port, Key(173) => 
                           reg_key_173_port, Key(172) => reg_key_172_port, 
                           Key(171) => reg_key_171_port, Key(170) => 
                           reg_key_170_port, Key(169) => reg_key_169_port, 
                           Key(168) => reg_key_168_port, Key(167) => 
                           reg_key_167_port, Key(166) => reg_key_166_port, 
                           Key(165) => reg_key_165_port, Key(164) => 
                           reg_key_164_port, Key(163) => reg_key_163_port, 
                           Key(162) => reg_key_162_port, Key(161) => 
                           reg_key_161_port, Key(160) => reg_key_160_port, 
                           Key(159) => reg_key_159_port, Key(158) => 
                           reg_key_158_port, Key(157) => reg_key_157_port, 
                           Key(156) => reg_key_156_port, Key(155) => 
                           reg_key_155_port, Key(154) => reg_key_154_port, 
                           Key(153) => reg_key_153_port, Key(152) => 
                           reg_key_152_port, Key(151) => reg_key_151_port, 
                           Key(150) => reg_key_150_port, Key(149) => 
                           reg_key_149_port, Key(148) => reg_key_148_port, 
                           Key(147) => reg_key_147_port, Key(146) => 
                           reg_key_146_port, Key(145) => reg_key_145_port, 
                           Key(144) => reg_key_144_port, Key(143) => 
                           reg_key_143_port, Key(142) => reg_key_142_port, 
                           Key(141) => reg_key_141_port, Key(140) => 
                           reg_key_140_port, Key(139) => reg_key_139_port, 
                           Key(138) => reg_key_138_port, Key(137) => 
                           reg_key_137_port, Key(136) => reg_key_136_port, 
                           Key(135) => reg_key_135_port, Key(134) => 
                           reg_key_134_port, Key(133) => reg_key_133_port, 
                           Key(132) => reg_key_132_port, Key(131) => 
                           reg_key_131_port, Key(130) => reg_key_130_port, 
                           Key(129) => reg_key_129_port, Key(128) => 
                           reg_key_128_port, Key(127) => reg_key_127_port, 
                           Key(126) => reg_key_126_port, Key(125) => 
                           reg_key_125_port, Key(124) => reg_key_124_port, 
                           Key(123) => reg_key_123_port, Key(122) => 
                           reg_key_122_port, Key(121) => reg_key_121_port, 
                           Key(120) => reg_key_120_port, Key(119) => 
                           reg_key_119_port, Key(118) => reg_key_118_port, 
                           Key(117) => reg_key_117_port, Key(116) => 
                           reg_key_116_port, Key(115) => reg_key_115_port, 
                           Key(114) => reg_key_114_port, Key(113) => 
                           reg_key_113_port, Key(112) => reg_key_112_port, 
                           Key(111) => reg_key_111_port, Key(110) => 
                           reg_key_110_port, Key(109) => reg_key_109_port, 
                           Key(108) => reg_key_108_port, Key(107) => 
                           reg_key_107_port, Key(106) => reg_key_106_port, 
                           Key(105) => reg_key_105_port, Key(104) => 
                           reg_key_104_port, Key(103) => reg_key_103_port, 
                           Key(102) => reg_key_102_port, Key(101) => 
                           reg_key_101_port, Key(100) => reg_key_100_port, 
                           Key(99) => reg_key_99_port, Key(98) => 
                           reg_key_98_port, Key(97) => reg_key_97_port, Key(96)
                           => reg_key_96_port, Key(95) => reg_key_95_port, 
                           Key(94) => reg_key_94_port, Key(93) => 
                           reg_key_93_port, Key(92) => reg_key_92_port, Key(91)
                           => reg_key_91_port, Key(90) => reg_key_90_port, 
                           Key(89) => reg_key_89_port, Key(88) => 
                           reg_key_88_port, Key(87) => reg_key_87_port, Key(86)
                           => reg_key_86_port, Key(85) => reg_key_85_port, 
                           Key(84) => reg_key_84_port, Key(83) => 
                           reg_key_83_port, Key(82) => reg_key_82_port, Key(81)
                           => reg_key_81_port, Key(80) => reg_key_80_port, 
                           Key(79) => reg_key_79_port, Key(78) => 
                           reg_key_78_port, Key(77) => reg_key_77_port, Key(76)
                           => reg_key_76_port, Key(75) => reg_key_75_port, 
                           Key(74) => reg_key_74_port, Key(73) => 
                           reg_key_73_port, Key(72) => reg_key_72_port, Key(71)
                           => reg_key_71_port, Key(70) => reg_key_70_port, 
                           Key(69) => reg_key_69_port, Key(68) => 
                           reg_key_68_port, Key(67) => reg_key_67_port, Key(66)
                           => reg_key_66_port, Key(65) => reg_key_65_port, 
                           Key(64) => reg_key_64_port, Key(63) => 
                           reg_key_63_port, Key(62) => reg_key_62_port, Key(61)
                           => reg_key_61_port, Key(60) => reg_key_60_port, 
                           Key(59) => reg_key_59_port, Key(58) => 
                           reg_key_58_port, Key(57) => reg_key_57_port, Key(56)
                           => reg_key_56_port, Key(55) => reg_key_55_port, 
                           Key(54) => reg_key_54_port, Key(53) => 
                           reg_key_53_port, Key(52) => reg_key_52_port, Key(51)
                           => reg_key_51_port, Key(50) => reg_key_50_port, 
                           Key(49) => reg_key_49_port, Key(48) => 
                           reg_key_48_port, Key(47) => reg_key_47_port, Key(46)
                           => reg_key_46_port, Key(45) => reg_key_45_port, 
                           Key(44) => reg_key_44_port, Key(43) => 
                           reg_key_43_port, Key(42) => reg_key_42_port, Key(41)
                           => reg_key_41_port, Key(40) => reg_key_40_port, 
                           Key(39) => reg_key_39_port, Key(38) => 
                           reg_key_38_port, Key(37) => reg_key_37_port, Key(36)
                           => reg_key_36_port, Key(35) => reg_key_35_port, 
                           Key(34) => reg_key_34_port, Key(33) => 
                           reg_key_33_port, Key(32) => reg_key_32_port, Key(31)
                           => reg_key_31_port, Key(30) => reg_key_30_port, 
                           Key(29) => reg_key_29_port, Key(28) => 
                           reg_key_28_port, Key(27) => reg_key_27_port, Key(26)
                           => reg_key_26_port, Key(25) => reg_key_25_port, 
                           Key(24) => reg_key_24_port, Key(23) => 
                           reg_key_23_port, Key(22) => reg_key_22_port, Key(21)
                           => reg_key_21_port, Key(20) => reg_key_20_port, 
                           Key(19) => reg_key_19_port, Key(18) => 
                           reg_key_18_port, Key(17) => reg_key_17_port, Key(16)
                           => reg_key_16_port, Key(15) => reg_key_15_port, 
                           Key(14) => reg_key_14_port, Key(13) => 
                           reg_key_13_port, Key(12) => reg_key_12_port, Key(11)
                           => reg_key_11_port, Key(10) => reg_key_10_port, 
                           Key(9) => reg_key_9_port, Key(8) => reg_key_8_port, 
                           Key(7) => reg_key_7_port, Key(6) => reg_key_6_port, 
                           Key(5) => reg_key_5_port, Key(4) => reg_key_4_port, 
                           Key(3) => reg_key_3_port, Key(2) => reg_key_2_port, 
                           Key(1) => reg_key_1_port, Key(0) => reg_key_0_port, 
                           Ciphertext(191) => reg_out_191_port, Ciphertext(190)
                           => reg_out_190_port, Ciphertext(189) => 
                           reg_out_189_port, Ciphertext(188) => 
                           reg_out_188_port, Ciphertext(187) => 
                           reg_out_187_port, Ciphertext(186) => 
                           reg_out_186_port, Ciphertext(185) => 
                           reg_out_185_port, Ciphertext(184) => 
                           reg_out_184_port, Ciphertext(183) => 
                           reg_out_183_port, Ciphertext(182) => 
                           reg_out_182_port, Ciphertext(181) => 
                           reg_out_181_port, Ciphertext(180) => 
                           reg_out_180_port, Ciphertext(179) => 
                           reg_out_179_port, Ciphertext(178) => 
                           reg_out_178_port, Ciphertext(177) => 
                           reg_out_177_port, Ciphertext(176) => 
                           reg_out_176_port, Ciphertext(175) => 
                           reg_out_175_port, Ciphertext(174) => 
                           reg_out_174_port, Ciphertext(173) => 
                           reg_out_173_port, Ciphertext(172) => 
                           reg_out_172_port, Ciphertext(171) => 
                           reg_out_171_port, Ciphertext(170) => 
                           reg_out_170_port, Ciphertext(169) => 
                           reg_out_169_port, Ciphertext(168) => 
                           reg_out_168_port, Ciphertext(167) => 
                           reg_out_167_port, Ciphertext(166) => 
                           reg_out_166_port, Ciphertext(165) => 
                           reg_out_165_port, Ciphertext(164) => 
                           reg_out_164_port, Ciphertext(163) => 
                           reg_out_163_port, Ciphertext(162) => 
                           reg_out_162_port, Ciphertext(161) => 
                           reg_out_161_port, Ciphertext(160) => 
                           reg_out_160_port, Ciphertext(159) => 
                           reg_out_159_port, Ciphertext(158) => 
                           reg_out_158_port, Ciphertext(157) => 
                           reg_out_157_port, Ciphertext(156) => 
                           reg_out_156_port, Ciphertext(155) => 
                           reg_out_155_port, Ciphertext(154) => 
                           reg_out_154_port, Ciphertext(153) => 
                           reg_out_153_port, Ciphertext(152) => 
                           reg_out_152_port, Ciphertext(151) => 
                           reg_out_151_port, Ciphertext(150) => 
                           reg_out_150_port, Ciphertext(149) => 
                           reg_out_149_port, Ciphertext(148) => 
                           reg_out_148_port, Ciphertext(147) => 
                           reg_out_147_port, Ciphertext(146) => 
                           reg_out_146_port, Ciphertext(145) => 
                           reg_out_145_port, Ciphertext(144) => 
                           reg_out_144_port, Ciphertext(143) => 
                           reg_out_143_port, Ciphertext(142) => 
                           reg_out_142_port, Ciphertext(141) => 
                           reg_out_141_port, Ciphertext(140) => 
                           reg_out_140_port, Ciphertext(139) => 
                           reg_out_139_port, Ciphertext(138) => 
                           reg_out_138_port, Ciphertext(137) => 
                           reg_out_137_port, Ciphertext(136) => 
                           reg_out_136_port, Ciphertext(135) => 
                           reg_out_135_port, Ciphertext(134) => 
                           reg_out_134_port, Ciphertext(133) => 
                           reg_out_133_port, Ciphertext(132) => 
                           reg_out_132_port, Ciphertext(131) => 
                           reg_out_131_port, Ciphertext(130) => 
                           reg_out_130_port, Ciphertext(129) => 
                           reg_out_129_port, Ciphertext(128) => 
                           reg_out_128_port, Ciphertext(127) => 
                           reg_out_127_port, Ciphertext(126) => 
                           reg_out_126_port, Ciphertext(125) => 
                           reg_out_125_port, Ciphertext(124) => 
                           reg_out_124_port, Ciphertext(123) => 
                           reg_out_123_port, Ciphertext(122) => 
                           reg_out_122_port, Ciphertext(121) => 
                           reg_out_121_port, Ciphertext(120) => 
                           reg_out_120_port, Ciphertext(119) => 
                           reg_out_119_port, Ciphertext(118) => 
                           reg_out_118_port, Ciphertext(117) => 
                           reg_out_117_port, Ciphertext(116) => 
                           reg_out_116_port, Ciphertext(115) => 
                           reg_out_115_port, Ciphertext(114) => 
                           reg_out_114_port, Ciphertext(113) => 
                           reg_out_113_port, Ciphertext(112) => 
                           reg_out_112_port, Ciphertext(111) => 
                           reg_out_111_port, Ciphertext(110) => 
                           reg_out_110_port, Ciphertext(109) => 
                           reg_out_109_port, Ciphertext(108) => 
                           reg_out_108_port, Ciphertext(107) => 
                           reg_out_107_port, Ciphertext(106) => 
                           reg_out_106_port, Ciphertext(105) => 
                           reg_out_105_port, Ciphertext(104) => 
                           reg_out_104_port, Ciphertext(103) => 
                           reg_out_103_port, Ciphertext(102) => 
                           reg_out_102_port, Ciphertext(101) => 
                           reg_out_101_port, Ciphertext(100) => 
                           reg_out_100_port, Ciphertext(99) => reg_out_99_port,
                           Ciphertext(98) => reg_out_98_port, Ciphertext(97) =>
                           reg_out_97_port, Ciphertext(96) => reg_out_96_port, 
                           Ciphertext(95) => reg_out_95_port, Ciphertext(94) =>
                           reg_out_94_port, Ciphertext(93) => reg_out_93_port, 
                           Ciphertext(92) => reg_out_92_port, Ciphertext(91) =>
                           reg_out_91_port, Ciphertext(90) => reg_out_90_port, 
                           Ciphertext(89) => reg_out_89_port, Ciphertext(88) =>
                           reg_out_88_port, Ciphertext(87) => reg_out_87_port, 
                           Ciphertext(86) => reg_out_86_port, Ciphertext(85) =>
                           reg_out_85_port, Ciphertext(84) => reg_out_84_port, 
                           Ciphertext(83) => reg_out_83_port, Ciphertext(82) =>
                           reg_out_82_port, Ciphertext(81) => reg_out_81_port, 
                           Ciphertext(80) => reg_out_80_port, Ciphertext(79) =>
                           reg_out_79_port, Ciphertext(78) => reg_out_78_port, 
                           Ciphertext(77) => reg_out_77_port, Ciphertext(76) =>
                           reg_out_76_port, Ciphertext(75) => reg_out_75_port, 
                           Ciphertext(74) => reg_out_74_port, Ciphertext(73) =>
                           reg_out_73_port, Ciphertext(72) => reg_out_72_port, 
                           Ciphertext(71) => reg_out_71_port, Ciphertext(70) =>
                           reg_out_70_port, Ciphertext(69) => reg_out_69_port, 
                           Ciphertext(68) => reg_out_68_port, Ciphertext(67) =>
                           reg_out_67_port, Ciphertext(66) => reg_out_66_port, 
                           Ciphertext(65) => reg_out_65_port, Ciphertext(64) =>
                           reg_out_64_port, Ciphertext(63) => reg_out_63_port, 
                           Ciphertext(62) => reg_out_62_port, Ciphertext(61) =>
                           reg_out_61_port, Ciphertext(60) => reg_out_60_port, 
                           Ciphertext(59) => reg_out_59_port, Ciphertext(58) =>
                           reg_out_58_port, Ciphertext(57) => reg_out_57_port, 
                           Ciphertext(56) => reg_out_56_port, Ciphertext(55) =>
                           reg_out_55_port, Ciphertext(54) => reg_out_54_port, 
                           Ciphertext(53) => reg_out_53_port, Ciphertext(52) =>
                           reg_out_52_port, Ciphertext(51) => reg_out_51_port, 
                           Ciphertext(50) => reg_out_50_port, Ciphertext(49) =>
                           reg_out_49_port, Ciphertext(48) => reg_out_48_port, 
                           Ciphertext(47) => reg_out_47_port, Ciphertext(46) =>
                           reg_out_46_port, Ciphertext(45) => reg_out_45_port, 
                           Ciphertext(44) => reg_out_44_port, Ciphertext(43) =>
                           reg_out_43_port, Ciphertext(42) => reg_out_42_port, 
                           Ciphertext(41) => reg_out_41_port, Ciphertext(40) =>
                           reg_out_40_port, Ciphertext(39) => reg_out_39_port, 
                           Ciphertext(38) => reg_out_38_port, Ciphertext(37) =>
                           reg_out_37_port, Ciphertext(36) => reg_out_36_port, 
                           Ciphertext(35) => reg_out_35_port, Ciphertext(34) =>
                           reg_out_34_port, Ciphertext(33) => reg_out_33_port, 
                           Ciphertext(32) => reg_out_32_port, Ciphertext(31) =>
                           reg_out_31_port, Ciphertext(30) => reg_out_30_port, 
                           Ciphertext(29) => reg_out_29_port, Ciphertext(28) =>
                           reg_out_28_port, Ciphertext(27) => reg_out_27_port, 
                           Ciphertext(26) => reg_out_26_port, Ciphertext(25) =>
                           reg_out_25_port, Ciphertext(24) => reg_out_24_port, 
                           Ciphertext(23) => reg_out_23_port, Ciphertext(22) =>
                           reg_out_22_port, Ciphertext(21) => reg_out_21_port, 
                           Ciphertext(20) => reg_out_20_port, Ciphertext(19) =>
                           reg_out_19_port, Ciphertext(18) => reg_out_18_port, 
                           Ciphertext(17) => reg_out_17_port, Ciphertext(16) =>
                           reg_out_16_port, Ciphertext(15) => reg_out_15_port, 
                           Ciphertext(14) => reg_out_14_port, Ciphertext(13) =>
                           reg_out_13_port, Ciphertext(12) => reg_out_12_port, 
                           Ciphertext(11) => reg_out_11_port, Ciphertext(10) =>
                           reg_out_10_port, Ciphertext(9) => reg_out_9_port, 
                           Ciphertext(8) => reg_out_8_port, Ciphertext(7) => 
                           reg_out_7_port, Ciphertext(6) => reg_out_6_port, 
                           Ciphertext(5) => reg_out_5_port, Ciphertext(4) => 
                           reg_out_4_port, Ciphertext(3) => reg_out_3_port, 
                           Ciphertext(2) => reg_out_2_port, Ciphertext(1) => 
                           reg_out_1_port, Ciphertext(0) => reg_out_0_port);
   Ciphertext_regx53x : DFFRS_X1 port map( D => reg_out_53_port, CK => clk, RN 
                           => n15, SN => n15, Q => Ciphertext(53), QN => n_1506
                           );
   Ciphertext_regx96x : DFFS_X1 port map( D => reg_out_96_port, CK => clk, SN 
                           => n14, Q => Ciphertext(96), QN => n_1507);
   Ciphertext_regx1x : DFF_X1 port map( D => reg_out_1_port, CK => clk, Q => 
                           Ciphertext(1), QN => n_1508);
   Ciphertext_regx69x : DFF_X1 port map( D => reg_out_69_port, CK => clk, Q => 
                           Ciphertext(69), QN => n_1509);
   Ciphertext_regx63x : DFF_X1 port map( D => reg_out_63_port, CK => clk, Q => 
                           Ciphertext(63), QN => n_1510);
   Ciphertext_regx19x : DFF_X1 port map( D => reg_out_19_port, CK => clk, Q => 
                           Ciphertext(19), QN => n_1511);
   Ciphertext_regx175x : DFF_X1 port map( D => reg_out_175_port, CK => clk, Q 
                           => Ciphertext(175), QN => n_1512);
   Ciphertext_regx104x : DFF_X1 port map( D => reg_out_104_port, CK => clk, Q 
                           => Ciphertext(104), QN => n_1513);
   Ciphertext_regx117x : DFF_X1 port map( D => reg_out_117_port, CK => clk, Q 
                           => Ciphertext(117), QN => n_1514);
   Ciphertext_regx67x : DFF_X1 port map( D => reg_out_67_port, CK => clk, Q => 
                           Ciphertext(67), QN => n_1515);
   Ciphertext_regx115x : DFF_X1 port map( D => reg_out_115_port, CK => clk, Q 
                           => Ciphertext(115), QN => n_1516);
   Ciphertext_regx151x : DFF_X1 port map( D => reg_out_151_port, CK => clk, Q 
                           => Ciphertext(151), QN => n_1517);
   Ciphertext_regx44x : DFF_X1 port map( D => reg_out_44_port, CK => clk, Q => 
                           Ciphertext(44), QN => n_1518);
   Ciphertext_regx109x : DFF_X1 port map( D => reg_out_109_port, CK => clk, Q 
                           => Ciphertext(109), QN => n_1519);
   Ciphertext_regx43x : DFF_X1 port map( D => reg_out_43_port, CK => clk, Q => 
                           Ciphertext(43), QN => n_1520);
   Ciphertext_regx20x : DFF_X1 port map( D => reg_out_20_port, CK => clk, Q => 
                           Ciphertext(20), QN => n_1521);
   Ciphertext_regx178x : DFF_X1 port map( D => reg_out_178_port, CK => clk, Q 
                           => Ciphertext(178), QN => n_1522);
   Ciphertext_regx81x : DFF_X1 port map( D => reg_out_81_port, CK => clk, Q => 
                           Ciphertext(81), QN => n_1523);
   Ciphertext_regx127x : DFF_X1 port map( D => reg_out_127_port, CK => clk, Q 
                           => Ciphertext(127), QN => n_1524);
   Ciphertext_regx99x : DFF_X1 port map( D => reg_out_99_port, CK => clk, Q => 
                           Ciphertext(99), QN => n_1525);
   Ciphertext_regx85x : DFF_X1 port map( D => reg_out_85_port, CK => clk, Q => 
                           Ciphertext(85), QN => n_1526);
   Ciphertext_regx97x : DFF_X1 port map( D => reg_out_97_port, CK => clk, Q => 
                           Ciphertext(97), QN => n_1527);
   Ciphertext_regx36x : DFF_X1 port map( D => reg_out_36_port, CK => clk, Q => 
                           Ciphertext(36), QN => n_1528);
   Ciphertext_regx166x : DFF_X1 port map( D => reg_out_166_port, CK => clk, Q 
                           => Ciphertext(166), QN => n_1529);
   Ciphertext_regx60x : DFF_X1 port map( D => reg_out_60_port, CK => clk, Q => 
                           Ciphertext(60), QN => n_1530);
   Ciphertext_regx119x : DFF_X1 port map( D => reg_out_119_port, CK => clk, Q 
                           => Ciphertext(119), QN => n_1531);
   Ciphertext_regx150x : DFF_X1 port map( D => reg_out_150_port, CK => clk, Q 
                           => Ciphertext(150), QN => n_1532);
   Ciphertext_regx111x : DFF_X1 port map( D => reg_out_111_port, CK => clk, Q 
                           => Ciphertext(111), QN => n_1533);
   Ciphertext_regx102x : DFF_X1 port map( D => reg_out_102_port, CK => clk, Q 
                           => Ciphertext(102), QN => n_1534);
   Ciphertext_regx134x : DFF_X1 port map( D => reg_out_134_port, CK => clk, Q 
                           => Ciphertext(134), QN => n_1535);
   Ciphertext_regx144x : DFF_X1 port map( D => reg_out_144_port, CK => clk, Q 
                           => Ciphertext(144), QN => n_1536);
   Ciphertext_regx182x : DFF_X1 port map( D => reg_out_182_port, CK => clk, Q 
                           => Ciphertext(182), QN => n_1537);
   Ciphertext_regx52x : DFF_X1 port map( D => reg_out_52_port, CK => clk, Q => 
                           Ciphertext(52), QN => n_1538);
   Ciphertext_regx16x : DFF_X1 port map( D => reg_out_16_port, CK => clk, Q => 
                           Ciphertext(16), QN => n_1539);
   Ciphertext_regx161x : DFF_X1 port map( D => reg_out_161_port, CK => clk, Q 
                           => Ciphertext(161), QN => n_1540);
   Ciphertext_regx186x : DFF_X1 port map( D => reg_out_186_port, CK => clk, Q 
                           => Ciphertext(186), QN => n_1541);
   Ciphertext_regx179x : DFF_X1 port map( D => reg_out_179_port, CK => clk, Q 
                           => Ciphertext(179), QN => n_1542);
   Ciphertext_regx61x : DFF_X1 port map( D => reg_out_61_port, CK => clk, Q => 
                           Ciphertext(61), QN => n_1543);
   Ciphertext_regx95x : DFF_X1 port map( D => reg_out_95_port, CK => clk, Q => 
                           Ciphertext(95), QN => n_1544);
   Ciphertext_regx107x : DFF_X1 port map( D => reg_out_107_port, CK => clk, Q 
                           => Ciphertext(107), QN => n_1545);
   Ciphertext_regx75x : DFF_X1 port map( D => reg_out_75_port, CK => clk, Q => 
                           Ciphertext(75), QN => n_1546);
   Ciphertext_regx110x : DFF_X1 port map( D => reg_out_110_port, CK => clk, Q 
                           => Ciphertext(110), QN => n_1547);
   Ciphertext_regx51x : DFF_X1 port map( D => reg_out_51_port, CK => clk, Q => 
                           Ciphertext(51), QN => n_1548);
   Ciphertext_regx184x : DFF_X1 port map( D => reg_out_184_port, CK => clk, Q 
                           => Ciphertext(184), QN => n_1549);
   Ciphertext_regx71x : DFF_X1 port map( D => reg_out_71_port, CK => clk, Q => 
                           Ciphertext(71), QN => n_1550);
   Ciphertext_regx123x : DFF_X1 port map( D => reg_out_123_port, CK => clk, Q 
                           => Ciphertext(123), QN => n_1551);
   Ciphertext_regx58x : DFF_X1 port map( D => reg_out_58_port, CK => clk, Q => 
                           Ciphertext(58), QN => n_1552);
   Ciphertext_regx93x : DFF_X1 port map( D => reg_out_93_port, CK => clk, Q => 
                           Ciphertext(93), QN => n_1553);
   Ciphertext_regx66x : DFF_X1 port map( D => reg_out_66_port, CK => clk, Q => 
                           Ciphertext(66), QN => n_1554);
   Ciphertext_regx76x : DFF_X1 port map( D => reg_out_76_port, CK => clk, Q => 
                           Ciphertext(76), QN => n_1555);
   Ciphertext_regx25x : DFF_X1 port map( D => reg_out_25_port, CK => clk, Q => 
                           Ciphertext(25), QN => n_1556);
   Ciphertext_regx113x : DFF_X1 port map( D => reg_out_113_port, CK => clk, Q 
                           => Ciphertext(113), QN => n_1557);
   Ciphertext_regx59x : DFF_X1 port map( D => reg_out_59_port, CK => clk, Q => 
                           Ciphertext(59), QN => n_1558);
   Ciphertext_regx48x : DFF_X1 port map( D => reg_out_48_port, CK => clk, Q => 
                           Ciphertext(48), QN => n_1559);
   Ciphertext_regx156x : DFF_X1 port map( D => reg_out_156_port, CK => clk, Q 
                           => Ciphertext(156), QN => n_1560);
   Ciphertext_regx174x : DFF_X1 port map( D => reg_out_174_port, CK => clk, Q 
                           => Ciphertext(174), QN => n_1561);
   Ciphertext_regx9x : DFF_X1 port map( D => reg_out_9_port, CK => clk, Q => 
                           Ciphertext(9), QN => n_1562);
   Ciphertext_regx153x : DFF_X1 port map( D => reg_out_153_port, CK => clk, Q 
                           => Ciphertext(153), QN => n_1563);
   Ciphertext_regx47x : DFF_X1 port map( D => reg_out_47_port, CK => clk, Q => 
                           Ciphertext(47), QN => n_1564);
   Ciphertext_regx173x : DFF_X1 port map( D => reg_out_173_port, CK => clk, Q 
                           => Ciphertext(173), QN => n_1565);
   Ciphertext_regx146x : DFF_X1 port map( D => reg_out_146_port, CK => clk, Q 
                           => Ciphertext(146), QN => n_1566);
   Ciphertext_regx55x : DFF_X1 port map( D => reg_out_55_port, CK => clk, Q => 
                           Ciphertext(55), QN => n_1567);
   Ciphertext_regx162x : DFF_X1 port map( D => reg_out_162_port, CK => clk, Q 
                           => Ciphertext(162), QN => n_1568);
   Ciphertext_regx78x : DFF_X1 port map( D => reg_out_78_port, CK => clk, Q => 
                           Ciphertext(78), QN => n_1569);
   Ciphertext_regx121x : DFF_X1 port map( D => reg_out_121_port, CK => clk, Q 
                           => Ciphertext(121), QN => n_1570);
   Ciphertext_regx181x : DFF_X1 port map( D => reg_out_181_port, CK => clk, Q 
                           => Ciphertext(181), QN => n_1571);
   Ciphertext_regx22x : DFF_X1 port map( D => reg_out_22_port, CK => clk, Q => 
                           Ciphertext(22), QN => n_1572);
   Ciphertext_regx40x : DFF_X1 port map( D => reg_out_40_port, CK => clk, Q => 
                           Ciphertext(40), QN => n_1573);
   Ciphertext_regx189x : DFF_X1 port map( D => reg_out_189_port, CK => clk, Q 
                           => Ciphertext(189), QN => n_1574);
   Ciphertext_regx12x : DFF_X1 port map( D => reg_out_12_port, CK => clk, Q => 
                           Ciphertext(12), QN => n_1575);
   n14 <= '1';
   n15 <= '1';

end SYN_Behavioral;
